`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
D5iQGM8ohyaKc+++vSoHdD9O+aFyQU9vU1I4OVN8kwaXg4DvIsa45TJbFXcEAgSB
xLS2NGqVjUJkmqtNmiw8/8ZE8EHsWcRLeGKgF398GccvxYwcVk5QYiVaZ3ZQ/EJd
AxG8qLEizpihKnKbXc+8+6OUrlJF4BqZKfXjIAbN3Qk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10528)
7Iui6og1/6fjvCj+yE8xMay72BcP2329h4tjmK0FdVMJKnv/9fvvLTCDD0WRSgGe
eZTzieLvQo5rsvHJLDBICSl8dtUW4tDJF8XjKSa5sAlXAB/nZmNoz9b6Xt12Ttz6
VjwWe8pdBNze7ZPu0vthzeBiqEcigrP7zEfKbif8a1SGAeCg43VBWlNQF4/ocVr3
vJdkuinUR8+RVYUa1pV+OITOYvM/EHe/835URia8p+jzGDwg7OyxKyhU3Q3NkK+w
dgVpYYHFLuTTt9rz139s/e+KWm202shnb8VUYrPsYq/mO7UABwVJZLryTrP8685+
cFx36iuBqvQZR9noB0LAIPAtTDaq3TJhKBo9uF1foFX+S4Kekwdellj2Xff2a9aY
JacK6nUPRi/eU26tB3jsbjr0IykHefO3q2U7dJ6DK+2aUHapjersDqkL4QXz0d23
ueozfXB6+crCi9/nNaYyubOo5zJqipbtToutpUFlV2QTJFi8YTxH4LE/T2jXnLFD
C6ShQprMtI4fMEQtpEYk4VwrVWmtNCfJzqDZdt4fZsJ9vKbd6+ucWfjBHzKOFoBp
j8NqUFV/OAefx9C9UVbP8IKInUffVXhwQViIMemZ3QitDgHsxWOrtJpDokuCisYa
L9gNxQmFqQBZUi7JROLefBz/hQMG/HVfv2H9oL4y9zZ4zFleonQjWqHaGWP3Gaob
ixenL1QCdX7uGP1tmHx9bNjRqsN8M4ArsssHaZfNdXavPspbe8uXLecBpMtdtXqQ
7ooeR5CM4s0xxR3S/U9pbLntkEyK12/zaqDtJAJZZgRYCEnRoYzEkovtybgwBYMR
+Az7bVNEfF08HADUBsDfw0gH9+/ymBdwhXvh2RyAzzz0lXM4dC6Gh8EWYb0fPo6K
4XLY8bvyY5wsl4VISar/54ljg0i/DQ+qQeniajq7fsTnIRsjPngHFJEbwNvFazdG
DBegEXJYaALxS0cYMXhXppVta9d81/kmGvFGmiESgHt12WlqgoL1i3mKEiojCmIt
Z3cH6/WsUmEidCWx24Qu4CSXxhCvvtbO3QORYD6gs5fD+zJba2BDqqJvRkchoeS0
rEyxsDqcAJL6C0X2E+HeK06Xe+FO3uYyekHRGDf4c6I9Oyi4PGCNCoyvLRis/UpP
eI30i+teZKBktq/wcoGJ2rf6oJPXoCuAtYJnyff75JvEnaNMWyzpKAmLxwZH0JIj
1VyAnSorbOonv9liq8+YumYUL7Pviik1DzRIUCQdvHO7J/lbEPykKKM2L4Gdlh1P
0/9BTfMonr6JliFqd2J4SNweUH0nwqN/AiiSs8Q5chPEbmZRJ3AWf/yW0Y592WYX
W4MomSI5GZKACHL+khLyygS8ujkpWmkhrZLbApbw+dePxyoAqdn2TgjibjhxpEex
lALh8VBJT4n75ZaLlH190/uLzNIAM2M6eixjNpOuvE/PoG4RBNV3Mo1gNtTGHBCK
c0VQeBOp+0Y3jNixZa3DmGxq+yAsdASBFkp1sF5vNCvZQZo+QRaNBAUcCtL6d0Gf
xjBZzdYQ0RYVbSanKDTMT+KqqkhmFtAv76Krv5MhqK0/PQaD4rk3dk6+cIoi/Uqy
wyKwLcnt2jRU1Gx6z6DB+o/bv8Ae9pPMvGZ08BYYIKNeyyDP5VcilAdS1G7h3fQL
d0KZnvsveBaZr6H7rrfWwcUo0JDQJEsCIYWUk8Y2HZdKLkmFIocgmJkBzpd/ec+G
6gdK53HbMoPBBdfAqH2XHuAZcobVB31EycY3M+XwiweLcGVdj1noqyFry1Xhg4sy
tKrpy8UEWFdy/h7aIIDYqOgebtmNscHDBD0jAGY+hXQkQsTh8NuhA1h/KB+SFL0l
OemRX66re2I1/qqv13d60taikDagqhXPmqMyQu61T5N9XGrocx1IKZAKqQyKSclM
jZkeKCy+BYnsYWTK4PG+8bWfXnI4EKIgxPiXTEV5M9rRlOb0FlAByTf7zYzhFqiS
9Y6Bjmh72zsBUYrSBdgvnH53dTcRuuk1ThT86LFtDOLFJt/kk2U9dPq0DKmT5DEo
ysrIYjDlStS5QAJi+t7zHX7eiDxAuZ7FEKMSFabgYhH53+9EC9i29LQ4bI8/6rpI
Qjm/R6xP72xMqqxn7k57p/gRuPoZG1d5NNDX8kcm0vPt8D7ZrV/LUtTJ9UJK9fAh
koREn0kpIyIJlDY4IEXtGf7o4dyxrmfSe9RqBW7rPPz4He3xgPcy6cH//3BUgWI/
LF/q6RUWtB6yx/rHkedIufYI1AYf1h7IT5pDJ2qoD7OgrM2fODrOC86Bn9Sx/pVv
F2OZmL1M5hry+68C9xOIdXe+rA6to+WNYwdb3/sZKY8xMtNKQVplxmgYbG4UmHLF
lWQF3CXqk2nUyLhgm99VQ4VrOSVnKntEvPkziAvTFPIf9mY90dQOXV7H+dInaak/
u72JWDrOAnyGZXG/IT6UYV4NJ4UPUsSn0ab9c8Ww/hCS4Ux9IqTp0no9wqpCJamJ
bAAhpieLPkzWtLwJZHz8p+TJi4VTWijdR5u9y036Qc0SjJEI5RoLFekC9vBIq35t
uvWqd5oPvKUDsHQt1gO6kL8ClHA1CMKYP2B9EavWnZClQ2akRoG/Q7epx7ePP+tv
md+1hSdba5iyRUfJ4WtpGQlfPYSyT5u9Tjj/3mIEEtN65ruW79ILB/kMeTPZXIc1
ZVfrQYeCJ6CK2TjJwxDROLzNGuAdyqTf/y5GH4xV8ThGMhmECvusl16mNIf715W4
bddGIF00rpkjhnkuUI3QOobsoZlwrvqkCHtlriKnHDAUKVRJtBgQy8m/RyJRv7r2
App0wj2y/9P05oeMhpgk74I6aWCdz4Kjn0j1ArimO9ac9vY5AvVJxWW05PzvcqQm
pPe51FPQ6h76TnzLd1X2HuGyMuOPLJ8FogO2W52ZwrkwaA3ABfDyTN1pfczwGQ6Q
Z1MFKscncQlDE3SK9muUpfPRmhFcWjIQA6dZOqyqsQlxaE9cVLX1inGHW/QNKv91
ahS+9j1oXWaO37IQWV5DRxS4u2Xxl544IBr1UjIFBXTPAbsagcpHSuvmvydGoh+U
iGFrl71mJebxUUDaG7fMKO+F+Z0tMXbdk48Jzt/ZgMoG4yZSwZ7anj+0FgZBgTfG
kIHApOGRwtxtxwYOu8bhX/C8DwPi4VdeWQI4Pd+0ygEVl1iin2l5ZOmi/mlb4Jf/
orFMvwyEn9NH2UIj2IfxeZg3uPJ3pvY5kYxY588o/v4yVHTXQVljbXVSCc4ElJxj
mvf+se6TVIz/kN86RgobIJ3DEXxUrlCQy0yVyp05v8eOcLSbgZrzaFKaxzkksCsK
0HnEDnzU9rAGadKVi/7cbzTWVkOzoa6otY3IIfuVJsIycsf34/2+PD1a4F2TmgfM
ly3rYbiN86fRG0tj6XqgffmvzIbiTvHQo2To8mnzau62w5h03PVZMe+LyoJBoEZR
iFypcLKffWwsXuwT3CC/IiidE4vU9S6bvbR+He41w0z5WMGOrxPwBfiacLcuXWCF
Pj0HWl/MvocW37Ta2aIqsPSe0nlbVepAJM9WbGzWVQPE94sRIvzF+jg7gMLRVi8K
0g1wwZeIgVDadCCTSoislfOLKFm4SM9SUTj2DaqqQSl6ebkezGtw7vOxn2NNo1g9
jrD8P35Cc1wKatQdHZq4Kc2N/njyEkAl1BpBTG/zY2oemqfFlTXX3hZPVo5BCo97
dDfJD9wlTMZcicUK9+CSTjEQS4epslgpFwJpTpzrVwzRutdXe+2J/omlf+oXfBwy
TWy2ITn8lVDLK+rFBMNFqyv29CX47e6gqyzanjzlk5yS1jAd7JFKsmJeg0BpKzt6
BBgPk9O15IrtTTUwg6q7i+YrG8fL2FT4OEM+3u9+UdqwwanIq1VFX4xwXYtQUs+z
f/j6k/mNM9E0s5+G8TDjJ9obc3tuZlHibEzpRE83/BVQoKSY/CmZhWij+dkItICk
q+sSzv9sM+AoJDp1VNfJNvsCKKe6WmafuFcbxiiOEAW21fL/noUh6da/23pEHtKF
9aTpwmiQEGsHD3CoQi9oGfpHkO95jZeALGDlTLtaMGCTiKl0aMz4McJjI1SDNeUV
DJV0LLjHTU4kN7YwSfUsOiy8o6zxcmbTJsmRCqaHGrFlga1wAJQreCDZTHbs7Ymy
9kvpB1IcNO+fpEWvlWK2Et7hb6eoKEnvpIzVMhCTIx5Zf6okxkDTYaoNTxPbAs1T
ueQcBTVivjUp1ajKaMC8FoxzzlONBz+iIWZJFyuIDPS5OPtmdOCCHWyyvnB0gW9A
Tx5w5pWH/Etfrl9jZVXqvWw+hejb6TAsXYWV/SfS2uxTWCMbP4hXW7+m3Htll35H
wO4UvgviDrBAVoEaz5jYLQeekZl8rQ3mLuSwSKHe9qOtNaRWw/2cZa2GFwFjmze7
9l5U/h7GS8DsCkT08lW8LewuKx8br95Bb7b2YQltNsvqJJHkqM2TD3QlViQEp4qZ
RBuo4lzjuIZDtXpQhUlOZ2S8YdbToWNesoWJfIep0zlKZWdK2greV5hqilDjZzWf
vIGJyS3fxzVItQDTp3MCIxpWHYsIW44mgprUPh10I2LO7NkiXail8M77tXR2ZXrS
wLO3nSN7GoHlynuycncalbo1mHaW7aOCLuIpHokC3+j1tl+Gapl9dCK37RnU9HWT
OSW+HARjYjYSwc/jXoUxIWOeaMa3qDOzccInjmRqEoS0tPU9Rhv2KMkN5XlITD1G
qZiTLTOx0un7TVIWT6OWaAaTcQJyd1c6PcCRecmZWdChwCnP+Z7FrIP/e2BOJY5O
+cTJbHITOW220D3k/Mwgs5hzzx9uwC0QEXIAUBcf/2+n1S7A0tJAV97tBAsuASDX
HoNywH+bru84/tmeCd2imwAJ0cMSUPOn9AjZ1UL993cgwLKLLF6s32mnLa6o8Kii
/jFiWDKGzEufWOQ72Hqh8XwiQUOZGCMAbWBjLi2ECB28CEzSOHwYTJkQ1RnjKVWd
pBybWSAuOMijOsYLW5Y6A8otJIgnMpIWsCDT75KPwqsuzGkCODM2U/zNeNGOu9Tm
U5yprZzxpwj3XWQAhKoxJjLo8P58KtV41OjL6xVHZVS+xCIUig5G3Dbg3yOzT37G
F/ROEms0SIzqrt8QLmqBJHMpdxeVUJVvE0rAmILWnmgriPdBdFRuldJiZrOLlzjX
hjc8BcAYqUTI0+BIP/yzyydZMiltET2qV7P9gxA5LXXKSn07+0V3hMU4B67EIi83
SvJa3tiRwmbeEYgff/+GwRZyossOljbfqYbwS+XIsbsx0zHyz7vdEXbRQHD+Yior
PxVmhBBJJ8bliKqH1bk8F1CTAzAANOF3tLkQ10QS3bVY7z0H5zB+RXVE8iTjBGwI
hrtvxP7ULQhrpAct6KiXoZcPzeAiHY/8JoBN81B79u8BY52WTubVgg4GCzlpSNZZ
+zpoLjQvXRn8E8DWtKvtt8zsrWgZLVAts7//ltznhtgOAjCeHg2YzCDn+dCM4Irf
8Ul6eibYjPaVeX4B2jAeW21MiNBsFMe1BBvoODsEM++h1G14zlrh6WykoAUpEpKg
ZiSzcZAjhH7H7krxS///Hh3BsW3XctXrkuW8UnW5oxinqtc7STcGVFfGdc/nE5jo
YO/lgA2PL3ZJvFKKW/GDI4as815k0bfKpKn96xD1XBA+3OGichatiNI6ieLsecQA
GyhGHspaczaSpzuekC3eyF4YBFKU/FBONyZBJghM2ChtPpWeH0gFjLxtN32Cmviu
JS+bn2jQKpCCDaGT9dv70Cy0Wqmj8pmtq5lS3sZRAJzE3hK5s6EAntasnuPvkBDI
jcgXkctH8QaoCu/n1PWUNqTh08EYCABt+0HANUZW5ZbAfS4iK0VL5z7GWAUt2Gj6
ulVcuJK65h2HE3cmkyQUpw9vIiumPr9DBknzK6d7e9fRxUFYNv1/TtbbvoZbmn+3
xCm8yR7RSjmIQZMGQMNAicoa1ogRegf+u8qHzpcKbOQKH+fAAUENuhAOQNMBGZYZ
LSWrWIQLc6/BCiC7FAPyF4PNIImLErcAX381H2TE15LGByCiE8Va8Dh3F3GJv30E
PcczeTcDIAiAznetQuty52+DNgPcIRptrbaH59KltfZ3RLffjRnG1n7Or/dL8C3c
hh4aeusGq+kPSjybUq96yFF3zKNue0W8ti1VZIW3v0uCrpJJR68r+G2/c+kK+u4x
V+KDaMRxv3SjuVVHWExWGmCMm0j2hGdIugqZA+qY8DX7Hy6OsMV4EL2PTr4PYpIF
it7YtxWuuM7t38r1Cd/dkrLlQCWEBeFxnLJSv3GMOyp+JQt1R8PPrEjYfX+2xB3m
CFpx7JSpARVEAv3hdsnZIWah9+EmXf5g7a1XHpactjFmMosunRKJb/l/tSDUzZru
M4MvCnYepctRmXQYAaRG6tq8KzqJJw9fwqbRRm0BBunuSbC4FxC5fSjssUlwXfJ/
VK8GYvO3RT2qYLaVfFf7k8MJWDwTc+1Z/0T0nNDgnTWbLlv2avDgeHDsSH1f3KLG
Teo6f1INQB5LqDSUw9SxMQyBURjAc51z4tAyBw9RT7EoKU2EHyQGwqEwqfGnDkcf
5+NHfKP/I86Z082dZ3hMk6wDgfosUWk8tUAh0ZDHl8Xo2vo8p9vUWzpAnbPPzoWb
yXn+A6z8g7qV175WJvYEZavLYUYfbupx2wFVtXOC1W0bzmVL61hsPgnOLjR9BjxG
RyLrmYNurj++3RGpZOfUYF7F/NLg2OobDnabjE1+b22Z1MguLtBMmrPn+XNppH22
QQ7n01RXPxwNqhi+o5TaT/FA4ynyZaSAIN9u8amJlpL3vfzQM5H5AI0BtbJr0Pm3
772w/Cpl7lHhTDGyvvuxfLcMp7j/sO74O+D1nzufnvhK6Fgcsl0R3pOkB2HWqB7l
9YlqY7q04tpvkUwFvdvD/HbvJ6XseyYl+pHSW1FMI3bYxttclndOkneupJ58LhN9
g2dA7jvE8DK63LU0JBk2thn8xS1xUviUYAP5Vejh+B5DSKsg3t80N3rYre8Cwr0d
nLCkJC10sDzZMpHJfDmmD8YxvjF1YzboSLden6WYv5IoLlCeONZDRwpzh5ZWdvU/
q7oH4L0how2C4AnCx5naCfzn3E7EKVWQLxqseKjXKAzbRJf3sRMZbVjSUJBoVVo4
eKeV8Jv2fhxZTY2MOjabqQdjsgH7OIOXFO/c/k/vsE5qs6ydTsNDqB3iDK3tgZhu
kV0U6Fdax/StT2YrPfOaQ2X4qirSoSnPJKtMJTpRRGyrbJHkptMPGyAXXpb1u1fT
MCSu1UShvH70kTgQTuOGrOMw0zM7inH1Cof7CfNwWBKwP2RmeKBB3p7Q0lbWgPBc
ZoOMNR/yxTfLXLn6b+kseBNEAW3EQo7Vr+NpWIv613Sa62rmun6raK0fISVzk23I
2ZlM+qwsLuyobIlGnV74dIm5HNNHDv0nMtkrDxjdzz0H3D5wIGWf4qZ5IP/vR/gJ
jeF22JemNxRp8bvAxrXzxX7oIUZ2ZuhnQ+V6adHKAHqnCcFtQhFGQZiYzJesaxdn
WGCG6lObAXuIKU3E/DUBoF9FZuVcuxPixFaqyzYp33Fqdfjkd2AbMDlOy0cwokP5
2MCtiUOtlVAfvRXdN0jlplNebRIGhQRWouxK4+7DgJTjR3Si7qj0sqebV4qKUzE0
6YsPHuNU2ENPKhYOSrUeAypxvYYDwRufLWZLQioDrzI95QyzXO6YHJ5i2GmyquxN
nM7fNm/QNHutfe8YYmvN++pd9zuG3tSVN28mQ/B/Ib+ThL9rrvw7+Mp1y/T3Yztd
BEncksaJ4m85CPVM7DgHr+5heGeJNwx0HxfR2PaxLkIsGVE2LmPSVKUOw2pxFy6T
VRXIUah42OXxIBih6QJtULRK6ZUElwmnuaxeHz/jo05e8D673WlM3lFblBdQ1Sau
Xo5W27BgTBM0v3UC8rg9AwhRsldkUoyouRxW5zacWyl1zMsjEuRhTsPbqoOyQoES
2gCMXtgN6vHuCFWL3qL/CZ0HDMbulIZv7P2bAxMmkmY6f0CGlB9KLgO5pqPUVWCi
aeOtNu9romLKV5lLKlwiToscJsIp3NtpeuLgr7gDkacPekvu1iJ7iyOTbkNpc6Ds
cEjaSHdIeZj1x0x1F6q3QnjeBBVZQXaAKsRIVcOmeq7LHDXWkp+Y58cXhOTlYN6c
rvc6JyCeSgtq8+GC9R9Nb0O+jmd5lmug3IdMsLc76KVu0a47wGcbxqtNhrtjGFYQ
00W+pEBve2+sPsjz6JLE44N/3VpwAFTl6sKtq8JHFSUw+gE2qnPvgUoRtrjubJ9Q
noYgtLOqROBcGKUAeMjjRkcsRtRfygYtyU0kjKIb+0Ct/dvEuZLdmkRazKOY4a/m
/cl5uCTtxSM/UT/arbjnEIwliKpKOToLaiB4dTkMV9zh8+coUK/el75tNNG8YF5T
YY2Zqj5SLb8h1i5++0uTBgfqhsfAucgmmwjUyUgnG/gY6cSRpa1hzuGqOrbmfkTG
SyXfzKqR3pCwMkODhH1hwgA1Yx0cM9OiLQjUQ7SsJgO6derOPBfs8yyoYMsDekcL
p3euMIwiBnNgOGvDx2aUzpUltMhW8L8zy0kQwH7cmIWmquFokc9oOAkDSzPlMjV2
k4M2D886d8HSf0xShbKMrlgUvnQwPIJo4/iwBNKrH0WKksbr5DZg9JO8nyrhcT0x
W5mrTHBPacgGq8JIxI+aE1SvNfxpj8csG0OK1LUgbXj4W9WogLeM4vH3KW3irn7G
73BmxB43QN7JCLWMKAOlUrT1u3/bYuHzsWEBi/DNpZksgV8hByFOImyuQi/H+FbY
FT0zcjSgFhCXbq43rsyxl0e8XdeRZ1v01b/6rzV1JAfUI/1/e7o7mPyQ6EpyLeV1
8UJfbSoxnqkxtcETsrUwbFE8uOU+rIL7b1wo06/UjnLY16pPioAFLKFTgfhK27oR
LXSn1zCQL5rYyU/Cyjag9m4dAsFVRg79yJUvZfCOfNmGrXcRf/dVcn4L0YL+ik/1
mJiBDkQv38xsTcq12qjmsFBeyVz+NPawAc4aQ6Kft09StqPYg1z9vxyQNWk8fkFK
PI0tlgAIvvmCdxXtJ2yqpV40V9QTSdFxEWQ4yzvjkV8992kml+AgeWahKuEp1u8w
ynBYfBvw+6cmNE4c5IMiEL15SWRlf2b/elvJK3gAD9IK5HyFOSclXsLStvQjYMx0
MtCFmX8aiMdZzJALb/qnGZ/Dgu53VIHRUXRboC4qDuCCr7qLPPeh4mFRFxCY3BHx
nHSBND/o1fdCPBCAXWe/mK/eQ2dr39r/+KGsD1uIAaKml45lJXcr9zbLHqdOW3m/
wLHqp3m3ScIITRRxFIFH3x8lJ615WsNrshE3nKAIkOhFAFRzRPbvxjjtKlq3oLEV
9SPQPW2hA7Q8x/xv72B9oUbtzOaIba1HO+rnJFO2ARH3q/XNzaWg4XsKLJ1QedOi
9OcmdBhsioACfiOZOhZgnhCPOZ3ITC47iskuzCyR0owUGADGBt1clMF+LrhRPEl4
QLtCvhOBjghk0vlz1FjD8dzchcIy0GJxt+MyaKnbNOJYEy7CwmwmLyfgaPaycg+T
LJszdcyH74GhvXzYG+swpM8aCnBKEYT1KRVqL7EwnY2MF82iKx+PM9wDWE4ZmN3O
R3l0p6P0H12fYVikAA30VV+UrKhI/SHMuxp14f6TV9Pel+zsNPSvvJM3oP07of8Q
30tedvFaGtAYzC/ZAdizqxCk98FZ5lmblIWaWGeKbbKfzKJHjoS2JHeDnEgM5T68
TI0ypmMAZlaUwwMJ8le+mkwp42DR2+edHze/wK3ILcFkQyBqMS8sMJ2VR2UyK1Wl
04Z3YmBrVeEjBqTpI+lk+OOnMWRj8m+t2P5E2pgcfmVf5XBNAplqEOiap3MjJgkv
WaVyfNJVBLNqUVFstUlbMMw9BxK8aLETeLkGqfynfviXsgKR8JXE8jXopGqYaEKP
i9/JEnxjSi+9UDL77BYnX22REEHeDrXjGue/DDXw22Zj+IrmYy510ijTYy8O38Rw
egAWXP9eB+5EP8NOKkECGSLb+a0tEfQlDF/cF4KZp84Fcvb6IGkSJYq6ZT5YJqXq
vwZ6FxRtMAfRctDtYUx+GO6GXBegQf4NNEFyYcHjCbb+AG4YDcWAeAqunBd6Xl/G
oe4UArdukn9hJUCnqGNKi0siyZ39UQMvlviPerH7DMr3q7WFkwx60z9LJPlozYT3
Na+INlLW6Zuc3vI5nbCXhshMPPfHaf9+ZT2JAZGc9zaZ6dcPZnfndQMq9uqSErPn
yA/A2+fhYFyP6XTzbeC5fzR0xUFY6ezD4SssQaxUOYZnFmZNGeIyOoC8a022FCSU
DvgSOyi8EQWHPQ+yHVb8m6K8qXg8zSFvZBQ+hc2kyKLRYrahQ54rjEMUL2woLtK2
lLpHNjZAeEZeUY5PltiBYJnLiVT5FPRDn+vow6sG0obglr99KB0Iy+0O/Ombyu3X
FrXnU+eq7agAAfyyQDhW9d5wau/qApUW7pcW4vDKgcc+gUNTVeJxGm37FGiw5v8l
InF0J/Pt4WToXkurxgbdegaH1qK4CsNUk9xfH2mITswZyHk7t5sWBCenetbAbWPI
6nTi6ppxybSd6z3g9jUfAgjpr/0j5sH+imzewQNOjcxKYkznF5c+OjFrQ4IW/Ykn
mXtp6lWbAbMhDsGlN3v59Jyx0JyuiGfKIUsDY0QjU7xKhxyQyvRNDZSxdIjoMp9B
A77klQmq5Y76PHU02gql7ALV1cd18uEMX9z6WqfTz57xSt0Hl8gonAyFgnvz2JXR
mR36kP7unpK8Fknbqf6JBGm2G3H1A7C1CvVxOH4OJODaZ+XXAVvdNAn0yuHRl/T0
1CNySYxg4mBnEmF4MBfYCD6q6sgpxIEchNewXet1dLxkJayNF8jHnl5RcWWdqdzn
6CV0PNaFLoAxK3Wp+HRDsKt0vnf4yN197jBVtYG2buduD63lSxtMOWUdJXip1nEN
phJ59Jox2GoZ+ehpNZhxl/tZDiCvZ/1yt5oUYc5/J6nOSeXx17T337ZuPnpY2ia/
an0s4EjEAU4S2bD9M/UlU8wu6Lf67AuHnn11jOPPN8XAYPHQAYYQvi1ceUY02VxO
ooS4bcofsZsBdWCZkLnvCmpCf5ox3/HSAaFqjUqxHyG6ZgMigScnwXVv9QCDPzf4
wNtQvudW+taxUO20Td/CMznYD5QiVOLBCv2lbNNcIbexxMt8Jp9v28gyXLkcNoi6
cCn/mJbiOKwVCK02jQzTev5wuQkYpdO4p3IPlsq7Lz8DPUXiQ9US2+eP/xRz3iDm
8eGi5MODa8LcjQ4P9NrBOD1a57slnwegj8F1RPC85Eoncazc9WpOz6pkC5JAL1LM
bflv2uHbotqNKuIDRe0XvBiOLFyLn+ftKksQmcZH44jhgVpvArfjMuQShN3OIQSB
aUfQw3SAhiZYiTBt74Pm4Dk7J3tcDP3ELiAOP3Hmkrh1klIFYdhHBtFq4Ppx9DRK
+EsyKohNxUIt3jRBoEyqno3dWyH04rpr2AtuMPTHmk4kaxmv4c0oiFzvWaUsqGx6
8VHE1sMxh7CMlQYIDX5UnUbQ82OpGUPA/MBnC9ZzMJRcB+I7xMC6nLruApQxE5Up
K+d0hZ84baEinek1E2dBRJOL/5qxvkLdAtQomdVYcW9/n2+F4syfovSy56magBrv
js9sP8vNX80FZ9BFhjQbR/bKR/f+hwaxOan6NMpND4f1OufVsEZKLr6lvfe/vVA0
uXB0GAXw4iTh/hFYsqbGv13VdeDO39PeNEgG+OsmM3yR8O9EjgeUIhh3cy7GzWhv
b+r2BZhjdJ8ZlUmZLL/2RsBLFFrOUcIu8uvdwvwF2suos4TRdrHYQwkxWL2DVhjk
lCAEi2jCJgh4/QAVezgjWV7os7LqyoBRBmLkSE4WUEtMV7+er01P2wV7g7rEJgq2
vNiIPmVw3O6a0L+lhJIGfjD1MEbeGWEdWE3rGMFNVmw0ssIpWymefYCbz9MmBsc6
x5qpgAa7bxEkG0oItBGkeFaqWe2/HvMGjl+1w8SFaOoxDx/DOcQuJsuoXAMR+Ycd
85rIXcHY8yZuNUGHl4C4tRCpRs/rEiTd9EGF7F8iVnQu1LfbVMCH7//shYaKoMV/
+rXQ6Dz+T4elI6JqHdbkOy61Swjy7UNwMsWcaiF7DXV7eDfKBO/0iq5OMjXJYor9
lz3opLRGySiYUL3ghADZ9YC3mJuOJ50hgPnvNV3mdZ6SJkIccSupo0qUASzctyKh
pPMM4cGPM60hziKpRb2Cy2cbKSRHGfkAY60rCSh0RuLRVbSRTaQk1VJsJndTYy/L
Efy0KkBlnisOfh2iCUXy0gJ3qZEAEkMTDZ65CwTQdOYeTxmdoenec0qWE1avSn5I
TfgH9tgAcrMtSbI2Atkgq7ABV1/ojTi0F353N8eNaaxe7Os/P3QrvzpWu5E6j6+I
e7UwXQ7cJ4gMRD57jFsO3QwuB8x+lMpWOFTGW7uOIduK1Xu9YBxSks7erkeuTyIS
MhnNZP5+j/EyMHKjMnyJfiZ9AzbFPTHcPi7Nl/KbVmla3fJBKQ7aaXRUd7bQRY3n
RPwY1osSsBoaXgtXkEeAhWpTmWZTh0/aykiDtQ53ZrmOVrpYsOHl3QwtDp2k/ugs
aQso9w7FG3EmNkHTFjH4//LUvew3BdRjznfoM/LcDGGAAXy8v+PL+U7itK/rJEUp
FFvkhUi1Sfu7TWYn5h+PeCPN1rDcz97zATNNhFKaw8gMnqx3XCl1bzEBCx/UKjqn
zdfCIMTwytQPt+4zFLVFb5+cLcK4Y74gE8OymsPowFaBxJzOMkX0m5kiM4NAvE33
NMF4t0NlgmwP5goF1SbIp1A82u0Rvl6BgO+d6cN7/PPd6PZjZN0ojR3DkPEjnRkk
EeO5aRvFKEpb++thSUJFY0kwEYP+1ReVDG7pySgLD+q+ONWAfTJmVCOvunx92KWH
UjP5GouBSlMVL6eDy6nd+QskAtAU+HKrV0jZa6DGpqxFY7bzyNpoEwBMcMga0FRT
nLkO5jmj2UtK2HMEc2rudSJ1OQx0tmO5oWSgysD3jcp1ciTLAKhlU0gC+06BxoEk
DDn0i6hLG678tyE2vH0oHzAAS3aDPM8d0/cBk/PFLHM/W7XXjSuCisK3FSLwv3vM
Z478BWY8YcRU14ddY0Zh+1oBLAmaldwT5W18BmAJzZ+4Or77CLV3L/oLIl0ehnnY
ExHVi0RsgN647SJzLzbR968JOpah9Qx27LpoeliqrLKtvfkJ4u/+9JjHiBhKG27Z
CzBLiAE1BHKHtk3JJYX7rU0Gey+OF1muXGGFDACReXHT/tqV0P6+BnLdten1bpf5
CCwcsDd7JV3idezxnutX4oh11fVS4nPce6B5mt4d0WdW5J22/KLHjMPko+UjjbDV
qCdOK1F+ZHCW7fu6HNtLkaxW/wjO0tjKYcQaogFOgdk5CehawVifeN9kSMzheVkS
JMvUXzZXXiboQ0lePcQiRlGqPC97sb8NiiBZ02BY121GeVoWnwI+NkdzFbCfA+KN
xLGw+X65GcHFZdO/O9qWFWAKl3ktZGNa+Hk8JZ+4GibDb/jI9INLqJb2kn2lU9pp
so5LBQVe68cyRukfxTnJyEXsg2fxj7O2OszTUf1xgTU11QCagXfdg5IksJqn1lim
QvERbhEga7tE8xD/debAsgzHgft0dzDpL7rVhIXIBTN8L1esrxLM6EF/+OA6umjS
zCd0vh9kePNUX84Uug8nrfH7wS7AVezKkFB9dXoD0tyeMVNsGVmsYX7G2P+7pzL+
FSlHDJI8XDG9QhmUQ7V8u5rm+BcQ/DuVx7Fh4BKxsMOltXYPzFe3wwqdr6Pb6rns
TwFpfp0HAeeP/atlVq+iyx/9O5x1vYwqYhrShzm+v8xfzvAT+RVNIEtSLdLnYusp
qM/FCPETIytSoVRgv1sTBPbko+1/owGMrH4/XSLxLFgHtSykopVl5dW3GowKkX1u
RHieAjZYLuYcYX9fOa4z9w==
`pragma protect end_protected
