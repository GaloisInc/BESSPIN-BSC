////////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2018  Bluespec, Inc.  ALL RIGHTS RESERVED.
// $Revision$
// $Date$
////////////////////////////////////////////////////////////////////////////////
//  Filename      : XilinxDDR4.bsv
//  Description   :
////////////////////////////////////////////////////////////////////////////////
package XilinxDDR4;

// Notes :

////////////////////////////////////////////////////////////////////////////////
/// Imports
////////////////////////////////////////////////////////////////////////////////
import DDR4                ::*;
import XilinxKCU105DDR4    ::*;

////////////////////////////////////////////////////////////////////////////////
/// Exports
////////////////////////////////////////////////////////////////////////////////
export DDR4                ::*;
export XilinxKCU105DDR4    ::*;

endpackage: XilinxDDR4
