-- Copyright 2000--2003 Bluespec, Inc.  All rights reserved.

-- $Id$

package FlexBitArith((+), (-)) where

(+) :: (Add kd k m, Add ld l m) => Bit k -> Bit l -> Bit m
(+) x y = (Prelude.+) (zeroExtend x) (zeroExtend y)

(-) :: (Add kd k m, Add ld l m) => Bit k -> Bit l -> Bit m
(-) x y = (Prelude.-) (zeroExtend x) (zeroExtend y)
