// Copyright (c) 2008- 2009 Bluespec, Inc.  All rights reserved.
// $Revision$
// $Date$

package SceMiPCIE;

// This package brings together the various FPGA-specific Sce-Mi over
// PCIe packages.

import SceMiVirtex5PCIE :: *;
import SceMiVirtex6PCIE :: *;
import SceMiKintex7PCIE :: *;
import SceMiVirtex7PCIE :: *;
import SceMiVirtexUltraScalePCIE :: *;
import SceMiDiniPCIE    :: *;
import SceMiArria10PCIE :: *;

export SceMiVirtex5PCIE :: *;
export SceMiVirtex6PCIE :: *;
export SceMiKintex7PCIE :: *;
export SceMiVirtex7PCIE :: *;
export SceMiVirtexUltraScalePCIE :: *;
export SceMiDiniPCIE    :: *;
export SceMiArria10PCIE :: *;

endpackage: SceMiPCIE
