// ddr2_v12_1.v

// Generated using ACDS version 12.1 177 at 2013.04.19.15:18:38

`timescale 1 ps / 1 ps
module ddr2_v12_1 (
		input  wire         pll_ref_clk,       //  pll_ref_clk.clk
		input  wire         global_reset_n,    // global_reset.reset_n
		input  wire         soft_reset_n,      //   soft_reset.reset_n
		output wire         afi_clk,           //      afi_clk.clk
		output wire         afi_half_clk,      // afi_half_clk.clk
		output wire         afi_reset_n,       //    afi_reset.reset_n
		output wire [15:0]  mem_a,             //       memory.mem_a
		output wire [2:0]   mem_ba,            //             .mem_ba
		output wire [1:0]   mem_ck,            //             .mem_ck
		output wire [1:0]   mem_ck_n,          //             .mem_ck_n
		output wire [1:0]   mem_cke,           //             .mem_cke
		output wire [1:0]   mem_cs_n,          //             .mem_cs_n
		output wire [7:0]   mem_dm,            //             .mem_dm
		output wire [0:0]   mem_ras_n,         //             .mem_ras_n
		output wire [0:0]   mem_cas_n,         //             .mem_cas_n
		output wire [0:0]   mem_we_n,          //             .mem_we_n
		inout  wire [63:0]  mem_dq,            //             .mem_dq
		inout  wire [7:0]   mem_dqs,           //             .mem_dqs
		inout  wire [7:0]   mem_dqs_n,         //             .mem_dqs_n
		output wire [1:0]   mem_odt,           //             .mem_odt
		output wire         avl_ready,         //          avl.waitrequest_n
		input  wire         avl_burstbegin,    //             .beginbursttransfer
		input  wire [29:0]  avl_addr,          //             .address
		output wire         avl_rdata_valid,   //             .readdatavalid
		output wire [255:0] avl_rdata,         //             .readdata
		input  wire [255:0] avl_wdata,         //             .writedata
		input  wire [31:0]  avl_be,            //             .byteenable
		input  wire         avl_read_req,      //             .read
		input  wire         avl_write_req,     //             .write
		input  wire [2:0]   avl_size,          //             .burstcount
		output wire         local_init_done,   //       status.local_init_done
		output wire         local_cal_success, //             .local_cal_success
		output wire         local_cal_fail,    //             .local_cal_fail
		input  wire         oct_rdn,           //          oct.rdn
		input  wire         oct_rup,           //             .rup
		input  wire [15:0]  csr_addr,          //          csr.address
		input  wire         csr_read_req,      //             .read
		output wire [31:0]  csr_rdata,         //             .readdata
		input  wire         csr_write_req,     //             .write
		input  wire [31:0]  csr_wdata,         //             .writedata
		output wire         csr_waitrequest,   //             .waitrequest
		input  wire [3:0]   csr_be,            //             .byteenable
		output wire         csr_rdata_valid    //             .readdatavalid
	);

	ddr2_v12_1_0002 ddr2_v12_1_inst (
		.pll_ref_clk       (pll_ref_clk),       //  pll_ref_clk.clk
		.global_reset_n    (global_reset_n),    // global_reset.reset_n
		.soft_reset_n      (soft_reset_n),      //   soft_reset.reset_n
		.afi_clk           (afi_clk),           //      afi_clk.clk
		.afi_half_clk      (afi_half_clk),      // afi_half_clk.clk
		.afi_reset_n       (afi_reset_n),       //    afi_reset.reset_n
		.mem_a             (mem_a),             //       memory.mem_a
		.mem_ba            (mem_ba),            //             .mem_ba
		.mem_ck            (mem_ck),            //             .mem_ck
		.mem_ck_n          (mem_ck_n),          //             .mem_ck_n
		.mem_cke           (mem_cke),           //             .mem_cke
		.mem_cs_n          (mem_cs_n),          //             .mem_cs_n
		.mem_dm            (mem_dm),            //             .mem_dm
		.mem_ras_n         (mem_ras_n),         //             .mem_ras_n
		.mem_cas_n         (mem_cas_n),         //             .mem_cas_n
		.mem_we_n          (mem_we_n),          //             .mem_we_n
		.mem_dq            (mem_dq),            //             .mem_dq
		.mem_dqs           (mem_dqs),           //             .mem_dqs
		.mem_dqs_n         (mem_dqs_n),         //             .mem_dqs_n
		.mem_odt           (mem_odt),           //             .mem_odt
		.avl_ready         (avl_ready),         //          avl.waitrequest_n
		.avl_burstbegin    (avl_burstbegin),    //             .beginbursttransfer
		.avl_addr          (avl_addr),          //             .address
		.avl_rdata_valid   (avl_rdata_valid),   //             .readdatavalid
		.avl_rdata         (avl_rdata),         //             .readdata
		.avl_wdata         (avl_wdata),         //             .writedata
		.avl_be            (avl_be),            //             .byteenable
		.avl_read_req      (avl_read_req),      //             .read
		.avl_write_req     (avl_write_req),     //             .write
		.avl_size          (avl_size),          //             .burstcount
		.local_init_done   (local_init_done),   //       status.local_init_done
		.local_cal_success (local_cal_success), //             .local_cal_success
		.local_cal_fail    (local_cal_fail),    //             .local_cal_fail
		.oct_rdn           (oct_rdn),           //          oct.rdn
		.oct_rup           (oct_rup),           //             .rup
		.csr_addr          (csr_addr),          //          csr.address
		.csr_read_req      (csr_read_req),      //             .read
		.csr_rdata         (csr_rdata),         //             .readdata
		.csr_write_req     (csr_write_req),     //             .write
		.csr_wdata         (csr_wdata),         //             .writedata
		.csr_waitrequest   (csr_waitrequest),   //             .waitrequest
		.csr_be            (csr_be),            //             .byteenable
		.csr_rdata_valid   (csr_rdata_valid)    //             .readdatavalid
	);

endmodule
