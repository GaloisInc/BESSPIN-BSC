// Copyright 2009-2010 Bluespec, Inc.  All rights reserved.
// $Revision$
// $Date$

package Contexts;

import ModuleContext::*;
import ModuleCollect::*;

import CBus::*;
import LBus::*;



export ModuleContext::*;
export ModuleCollect::*;

endpackage
