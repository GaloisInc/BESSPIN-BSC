`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZukkqP08OWu8JRwgjUM14HeLOIShXA+i3pF9tlOGRCPGSvLMUSgIS+I3pCAt7TKt
ZUpZ0hWqoCh98uj4fFRv6hdKG8srtz6U4P9tZUZd5fjvj9pc8/d573uPGRFlVIMc
4DiIj7B/iZ3ZlAroISc6rfGoVxob7OtLksZI7ebZIm8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31712)
LLilicl25T43svM1APOI7eWuK0f4iROE8QZBEEz2oP8ELdTBlTrKapDCt6TNEkqH
IM4K2qxTuthpAqj312Uw8U5pXt+KlELpjnDWIOJ5F6eFM//6WXUFL6arq3kifpsR
9Zve1az/ICJZW86T/a9ytb+MaJYWCfsTpJL/T4i2f/joGsqKUZJhj3Qm3DMsgfCC
ZoMMjZXQ0bBTQioKgwsuLTaOm3o6V2PFX7ctqgaaY4/iow9H5aNDDzSH/AkLlj6B
uHP2n01s+ISKDJboA8cUbgjrbbK52SJSyd4D2mGCoXy6LaG3pDbkpZ0BSm/rTJK5
xWIKeOHOm09uLTlNm1tuFSdavOtyxYIgyMyer9IQfcKbiypmaKjlOOcvCpuNZUQ0
qc2AVaRfRV9ak6sgvFe2Z88Gd1rLF9MJrw5QvHIhV7Hwn5b3VwWBEHvYpfSpxRKm
XI8s722Os7tUXEa5JugEbDayYD9OxK8vMEggHvr/Gmn9K4AzeCKRknDyBjmWPK6c
JaFHLYkto/yZvhg9oVzqRj7L2kZIXu6i230e7zTAOAvPy8sT5KXdllFvsinHb/3E
q/omP7VTqZljWAQz8F4q4LGUhCNueTJ5y/UBeP0KSYH/vM6NEc5X4kTaPGU3jk54
9x1XJi2I6pXuqi7MPD5PdEF2BhRvqkF7ZSeNM9r+7TNSTYbdjQRJIZzIkammLJTM
w+Xh+6mPcmHbple/JTngnDGzwuEAYHhY8Z818u5btK/HiC1cE1oHuoAgUJZGhI2Q
QpWtOtN9CwJwIHKTfIz/vryYk9LaqEemHCgOqik66bUoCbccGIfIgJBm4PSKCKUr
0JuH5futI/d1THdkRGfCoIihGjvHX6oe9AxNYUwUAAnVQTUs2CJpSSTOfbGcZ/Qe
/zdo/UFocMe5+8SMq3hbx1Qa23wqL8Nx4kv3D88kP/pxSnyZ8qrduX/cAHZ+Kige
KuFFdwHjjyMsio4tc0tl71bynkuxZeMXqWNB5MQnJOA4dpaHBcf5M5BRC1JDpaV3
PFIcX6BnXC1jPDUL2fOHvzbBEewGKlcFKoHKK94H1ds5DcJ+KdgVkKPWXwgCarb8
YUKSSviHOKAgoISQmWZUouqUg0UaH6gkB2TT29f14PdD/AbY8H4PNOC5R6pvjrsb
W5RB1kElAj7k4z/apJCOY8PK2L1yZGC84GRv1pPGCa1L1BnGgYtJshuGHsUuqq73
o92Nxy7kDuXh38E6XDgRkJC+byNXD+t2FA4Gtl3rBZzvV8PV1Qch5p9ZjJn0xtgn
lquDEaw+C8CRTK7+1dmU03R/X7niEMzGHEdDDeXg/VIqIsnj1h1JGSnEAA6XcP/L
f3hExgc22YJjwy4Gf7rsjwh8q5155Nmv6Z+8fOasSAO5AvHjX45V6B3JS+z7cvZx
d0VljpY1Fm8p/4Y6oSP2kHQ82GKIIfF72aZDJaOk82/VRPqpAICf52b5wjmS1Rfg
7XlJ10pNZWlpSsJ07ui6DsiirSgia+RFOElf7zaAA1tjuEMa+VGsnyVUXn23LLJf
grPwR9ISVOxB705Apt5BbZhMTsxyE5GxWjTX0rA++V4X8fxum8c+xQawW+1eVr2H
vsbDD9Vs0c4JlODr/wThEQ6AYu0ZayQHhjpjI6gQ1hRHPIsnMlV0do0jwgmQJ8jw
upNC78/pstmsKw8GAN6ENrdnwN7c0qdFjLvFd5axc/fjguNqRp8uSvg+Yc9h8TAL
g0G5kspo3cmhwdWXRrkky15QLCQhCOVWVPHoCHgs4Kl9juQThLk1h0VOQ4Nedqaq
RHZhMGVO416YOkcRhoNbk0dk0Z0ruXySCA5FIiQgOdwHzHcOcjeUSTGTzP7TZ9ZU
jzpcwvYFt0g+a+7YVVHCMuostnUgHY480bsbO7fpfwusnpm2HDyARQ3vhWksBeUb
pJ7mFdedNBWUFTNjTgnoNMkZgxKK/0WqAmS/ACEG/Y5wHuYtvC/hTgQpdcp51e84
CrrpBDEt3u4J1Ymdf8JEe+R4119P9EWlGKv04KrqTqtseAoXEO6eDgmrvaHPAqtQ
lnMka0da3Irfy3LY9L27zTjPA+GhpTrs3RX4J75arqsDQFVTitpt3znbEKfhvUwl
Eg375sow62+Xj97lUNJO5vMcjOogBV9vCSgmh9zQNRzatqCzhGzGLpyH23yFomv+
O/qGHAhAuUWODgsThNoflO/6jjwXQO80HEU3Nvq/isbuhzXvdN4iCek/JFtBPR2s
jJteQRzt+RXSVGjbGKC79wILE9mWHfsZN72iafA4eovmU0zUKOw/6ugCJaVq5YtL
rpeMCBzYuVn6hfs4oT6ksGGIaCu1mjA91pTlOzQEHkRtD1jeIP5vREFAozQ/eOIP
IUH3IVOV11U+I4RGQ9fh42uRWSnQPwluxTSZzrEBAxYVbQZyYE3aiAxpGxngbkZl
R4YtFMUuZRLa0Onhwi1rTeVubCtES2oC4SpNv7fczFzNzfls8qYDzvGUsybZu0LE
HCmi/M6QhlCPsOyM00BZUzytMInrzeUFaAbf1NUju1SyJWeOQ2h5iRn5je0YoGfB
FGtnq6JWYvHrMNHPKAX2fWJ2L4RAm2mMl1pBTtRj6Stq1Ugz7yxMiMS+Ksxho6IZ
198ateRkVxVZNpYhGH6FfnApco7FbwIx1SaCzXPhzP9TSHYrBFDIGm/BedbgFDqD
18KLACaqjzJm8KombKPuSFmvE2w0fTQTNOPxQJdta9SJ1AFFIGa/FPazn9/zlnds
c+0QXurnXuNeXmMGOXOoaXULj1Y7IP7Mn/pqWJwkU/onKkXNJuDSTOBGwuKOihUG
kLQSO8n636ffwP/WW11UYfUUJxDNxPzDyPaNeuRaZYYR0WUc29+3IceUW7G4H3O4
Uv4eEKt+BXPdijt/yApEoJKXGHyVwGH9S/3qn+gl9UE5A+LyC3wHcaJhTz4jCG1S
3chVzyAjIkZVSz1OkPgi76RZQao/l4jB6WsNhgUUWbgvh6m29ixNIpuQG2+kVQh3
OzEYRIxTQPpdvBH24h77kKDbMiBG9ktMDfDMnvYMNIHdXRbB6IL0G3XfgKGBYdq9
RFb9Q8vb78eROhiZBNvOnYmJeGzLkbCZ4G4wds/YhaAQ73XrkTStkTmw3VXmTBkC
hKicbX+JEDtxEJID9ce5t6R4O2Jekrjgcvskyc+nA26Ht54+96NHxFq/RuOccNlt
dpaBqvoqXQI+3g0GflLhIMpKZ6TGHTMC1BaEPrHnSR9NfSw1y7VOhVBOTyld+1h/
R0aPMs7mXoSgZXu813YfydGO7UFIoFwOVuqs8LxFtBw9L6BVjRA/RLuwSew0baMe
Domyo1+WNI14t7ykXKdUE9QSIxDUSZclHsQj919jpoN33xWex4uYUBRSEwNbd21i
yZK3hlvGdXAp86eqs2JLZpTjFs6Vtd23iM7B1tmAR7WFTVCyfwYH2ZJbc002RhD2
x5YPn3uL7owOun5E1raCb3g7ndXm4YH+KTSLM15fA2zVis0iQbUvfNHVgCIV3ea3
EqhisZP8W6TalnGkX4FypVUvD8hEKSXsYyk2FjVF2Hk+a/xhcfGF6GuYPDAvt9F7
AXheVMc+Jj8evvxxy1VjGEMT9N2qJc3AeFsF3FzXmQbRZS3nnYLhhcaMT0oh0NoW
mr1sU3ACMrCR4oxIpgmD3yMNaMhI2KdF1OBnqyOWUcqbNdDptF6U1fWgzREXPRvQ
1ivkPlIbBFZ5zO+Ukbip+6BRe5lUWq8HZGST9RK5AFBAAdYN1Olop55K4+3/VT7J
5A+daNMQxUr48LecrVYwu88tBaN7a/Qo7LnXoHdnCjfWW6EBccuLuyWNnwrHr1of
DVOUKVifBlwK7iT2dkBYRVsIPhuWespmnlAOz4w+UBHBOLRlKI3aTs2NZulZFbX4
YA1+eAaX004uhVM1n2zeaunRVIHGUbyc4WHJ4+LkPVjfRRKJ6Y453824S40KUopq
/9TKzsfHZVUav75RsLZRorIRU7rEXvQeDnbfCMGv6C0FtNRMkERPM9tSR9qNZiGp
MQiaN/l4XdiFbQNlcQ1yZtBhAUbmSFowQSd9dRzXSMSAJZF5Qpozy80zRSNdlXT1
ASR8Y/xIyrgrW0xJgwAUiLpFvMqcK/uYqhaykva8EEypevOkOrdrzUBn5Mjvl+Zd
Pe0BAFyqKBd4KGkUqKObDDBZYeqUy/yK+ePJxgzgpVsLojZv/sCTdsQan00M8wPh
3CeDm3ZYCd5BNMAjz9jDyu7hNd14kY9/NlgBSSwfYafeV0NnSAOgcWsydZ5vBakh
k6ngaEVUP+9EAowW08YKvhe/j87ZbtjHG0GFxPcyjwxS4VDzmKZDT0FlFGMUiIXn
WSKoUyU/hvvKRpF/5qIcTQ6BGD08NTrSoukGaM2Rfba5kdh7CMOAj98ipzvCLf+5
YVkfNfjT9RnACwgfE0s1JAOrZfEhA2fXZaziWQ17CEGBrPlrHZ16aodEkqXmNybL
H5uJH5rc+y/25ROFzQxs6/jbWTxI1kMj9dRLn6B6NiZdP9jACUUsL6yu1/NZ50+e
ZVxdsheZnYPWJz1wfEa5dD4BLRUToLjl6YguLb4CMBU1VY6aF7LtLWHoq7xKdAf6
yB+PcqzU4ioPkXqAlYdkwpQXgQOjtXGni+qCFC1ruDwBG22MyFxSb9u7CP0kXUrK
QgW+5J4zwONCps+UCrNoeIFc6iGNZRCSwfB+oti8y1/9ivxXjcB3zl/lPy/e3rWc
Rab11+ZwCIq8CfxUfcqHA21WUqwYSaP/TGPduB2k4AnQNBDgf6PTgOzK8U26kbCS
VF2FrHanrhY/BFturOdUWk/lzhnqxZvaQ0fdmnqSWzp/4ZfHQtPCyOsLwxXpVyb7
vnjM41PN1uLtBs8NX0qDJAzH5+LL1Mi7hw8izkl7vM5Bf75J1ZhAzEhcMHkzUtJ5
mVO3ociioZZOizMHsVUmLobHTK4GxUnUZYpWlKKgGHVwN8+rwXW7n7kqTFUuuU6O
s5yAelIox48NPDwzsygkmfVHpWgHot1Uvfs0KMtu9+M7Er3POkQ4nZLD6w4PbMUt
ZQEGIaOON3lCRj5DQa7kerx41bNr0gSSqt46JHIBzhxtwRGuEdkGhxdqfWD0p1bt
Byjx5P2GdwsXdmzzvw2EmCtJ/KOA+Sg/F5AO1Oh38dD8XcqS4p32n6uxrBt/qsqd
J751rMsgrn/BAevQnRhZB3NVRqz7CfKkrKPlbxplLElqZXq8rXL6bCMukru/TeZH
wHamF4lU+OqV/suL59LkpjqkYaFa9Oid0X4DQ//u8YznkSNC9cHh9tOyiwApM3yh
kJNaHhmLikVvCArmGfBOWgjgcq4GPnw2BdHyFzglc7QYFGRDXcKEGtvo+2oF4epa
EadcoHtx54VZ2oFpFO1W0e/14w3zG+qvy1Bmywxbqbd4jBf9aRT/FpQwclbjwIRl
UEWJZ8SP9a9Z8PI3pKacfGGIaQ/oUX7z9X9j7EZwfp8vJqLjMcE8YjtVpSsDTYov
t8a7jeKde9aroomY/w3RDw6n/rmIiPuQu0fU0KlhErAQQDITSRD2dWQCwdSmBxdl
rj1q2XY0dQH73xLTDu6ATtC6tG/3yycaTDYdZG7EgqsH4aDxvHup7DS9gohhJGa3
G7UlzH6u8IYX03bddYmpxE82vPNXIprEDg1btoJcXtqOYYBcIAo1nvUAyvICE5yl
h311iYp3SdElkxuctfL4A7CW5Cj1TJvoOqOuO58SDcOl2LTV0pLWACQgxvZ4Es9y
AhNiPAuMn4BNqYNIDoux8bbnn2OyPhujc2hqFlqiUsgwDMu/aBmNbekOME9EHjIZ
0L2Qa3CD/QLXESCQ9TkQa9J5w55QV9A/eRHdswTGXz4rVrj2Kgrh2LKV+C8k1AsX
dXVfQR16SRektxPqeKlx7M6A20oPaGumM/OrOZy3HfR3aYlvspAb1Xlxy0ocSmxZ
8ZX4EPpNxXjKO5tUlnp1Q9LNX3RfVl9DOMpJ/gqPsCqI1Vwd/202J3q4XBLYlFdt
Vnyrq1izFjvu/nq3GjLBA7oc5qdx/VIuhg+gl5l0M9017oueR9ozUQIgx9aQkHl5
2uxBnFu68mKcCfstcmI9ACqCdXpZ/n+spgRvnsp/7oHgQEWu17rzQ4xVcw4mbwH7
lyvnQNXIh+E0hprQouWIHPhdKx6siEZONwqc8yIPeEBfuL8CpU79CASRwCmJTBtu
4g0ye2B3B36zo/9CotglctPxpbQTiJv5S2bfomNfXdd4h5O33egBkJOmsiYWouV9
+WA4I3iRDA1SKWxI9t7j+ollaLbb6hR1nOEnZRrqRG+LqiKDFiy2UM7yiKNWy9Tb
VWkyu3BGXSz6RBa662RDjJpxsrNguXKuQiryndgjZO3/IVhJr97PauozV2o/qBgV
w1SexeSzBRJoxmt9lNKL7PwCsQaiQQOqkU/frv5LCwFwnb6fRu7lNTL7i4t1mK3Z
0dq5vDYOwwbYoJ00UhwGxI+cdouc3VqcB+Y3rDSO0J6TECLhhvfTk/To0vJX9ljT
tvqZ9RxsMof8NlEw2HM7Je1VCnjdRetYMI9yWUvzoqiIoLxKdaerHgaSupidjzHY
cbOwg82L0qIAYOrWK9r1Ufc/FuG5UUhvg5B5Jeq8RgOqjF/lTHMWbfFC01Wt2Bzv
KA6Gnz0TPU5YbpEH9gHtuAyKQw027CqvPxVNPqjlmrWKbVUPW004H/6P1H0Bm7ej
9RmpTeMHjfHLqS6pPCSiCdBuesSIYY9brH7GWQvR7VqAMTMSSq1RJffVu+ed1JRb
QFzgnhdUQWbOqs+1O1Z47+arcGmZThbM7qs/lu+wTglvEyBVWYxBldMlNxMV8Y+u
AP5XbpDmqcbDta7Lhf9nrmnTtE9JvX3VvNe6fTXJ9ViQEOl0z+CA5U5Kn8mxz5PW
BC862ojE/iJEJ7NHIfFrc3gfjnrOCcx7uVUfyLIPdMwhJ7Q4mNyG/BKQuP7mq1ER
8eAN+K4u3mCoWs345MwZeyQdXDsmJ6eRMxrZzIZiND/aNWdwiE6mQz0r1pzjDZm6
PmWVRZY8vT66qjjnKhbdgFgKQ7AXD4xk2a150QA7YWoyyBqtqJgeugIeVEnZEPWn
hJEl0HW4hKJFMNceuspwidLRJu1AMnYzxUOUhCm62CiZ3oFrv1JctXhZjHySsBMy
Z0i5otUlQWOPbCgHZ5ZrE21v+VBxlSCINNS3BJlTwUU1QXfbovhSk1XBMiESso2m
zHgcp2zqG09F4KIQoFs/GF1Iifti247AV8iCUxgOvlml1ETIf/lXZe4GkP4Sv8CH
OJXlqvvKgUt8+DrxPhy84YBL1NomM46G9PqG8sOOwRYo0zSMuPLK/bzhGLzL7OxM
NIm7wLHjAiHga7A81OXC/JN0AGEYUq8cbiNEw5ZcHvMuxAbBKSsZ9qtkoFVAkVKg
IY7ZpCp1oENbLnE7Q9no5oCsVC+r1SN1iV53wcd1iWfowO8thaLexHfusk3mHZTb
E+1BrbUP3sSFF0vjOXviOO+7Zi8274aTvUooOZY2mswj/UQtQbGn7ump7EhCTW72
fzdj0RQwmnJ+2BnyCufZqZYDHXsjbsXigNvhRohjlhZ5YKAZP7jMlaSf3tP9Juio
0uNIM5zkptnREkbCdWdmuBpZcxAvmYYUWMLEhROdgC4hUbvSLHMJmsmSIBJadhEb
ya8uq1M0Gha+riqN0HyL3GaTbiEaVaEct89APA95lF79o5m7Iwl1G0tFPo214MTw
QYWp2s0p4LftLL5zPT+MCYf+bgPXK+pCMIz97ZMAybufx+2Hoefnjyrk3VZYhFxb
cvYcVPxl0T5R+BhZIxPOdV4/+SsI8NvGpw+6y1SfN2mEG8tAvyRaiAj1qlJNpByx
zIuCc0CJ+TtQfvmlljFl617kdWFeQ6HBwW2wH9cS5xsOvYa4r/1wG/SgxKQoVl2E
B8ES9MhyPCQA9XdrZ+9Xws2HSHIm3pnDzgi1LKoOpab+v/ril6+11wMp97OFtRGf
cgtI/VSnt5KCgG1ZP4lAMux0fJKN2CEQf9nMsiLsULhmcR20i55PetUgY9GS27Yk
nrv4dzS9wflK8I18agBpgsuFa0zd3oym+z3q+9LszAzGyvIPrywGY/h6ITB3zU35
nrb0PNenkZT8tfJjcSc7F+1S5nVhiiZLk9s6i/7bFir8X+/0ff/XHuRaeAfKuwsm
mgBkjozATlf7pH8m0UYL9Hu8mv7CXZRK1NW4sR3o4tCghaTC5LjTuWUov3AIyaqC
Gmpf665cCyM2n+WKfAZ/LPy929RmwIGAF+Xbm/r/nNkOcL34DEq507NVSaRAJy69
zzeSRFKdqXztfcuAz6A+8rfAyf5ylmVmGbXE0ypz+GdZoaH2hwafZXUYMr+rxHE6
5QZGJudFhLHw+Eq8nepoo9SyzGjfh0tZtprAvBSi0bdq4q/ys2+DRGbN6Yauku75
i5yUlMZ1NnlGbvp44iByt3SNOgN4CopK/a7LJGrIP4jMLYjpyRuPBmwVJAjrAbNi
+9TBSvwa4F1i5OBg4dBLIlvQHJSxZbfAGFK7Igdc0VPqiAlF/7LIPirBEJHFa9RF
V17TNBR41CzceUYp/3dMQId9O/ZkNR6z84i7nny7KztdS7sl2dblwEV4Tc7wsBwH
0qn3bvVG3llib0UbEa9jovutdj+IVHfkMFmdqAvU5q47ripIeOvAczf9yPLloZUt
zH4wRHycJcI8M6yYXscwhiqQ2wPKMCPCXcK1RxKOrgfqSdb7PfLkNFIE7vPdGD0I
k8N3+TK2mBxdY+hcz3lA0HeDdZk2U93kJIKn7Et2sM6atpiYdss2rL2Mdpe8Anlt
/U7XZ9WdrSLKOkdRwjqlA9HRHXBvLMgH5NCkKnKb4uxUWKrtI5C6D2nAW6jqNku5
djm40hQ1dvd4f1uTuxBd3NJmh02yBkfqk+faSNklA54jyqydceEF64XpZwdeBnRB
PNuabH4aPb9pyViSSM2oxtBYEH61wXImYXaLMY5ZMkRazhgItr1oqml8qQC+AvaZ
eYPiREbnFzkBjxpu/8EGbBCAAhe6kAj9vuwNCIKqyICu4DKf+rAA+xoiFgUpGQba
nDY04HuCno4uScTwY1fK/MywYZLgtRdW2NfEcEOPHFR6qqFHD2FRUk+lSl0c85hz
Yl41VTZ7QQb5KLSCtzPwHHDjuh0YeLkbyZmeULpP8M/Zp1YNtlEINua7R+zzLmW2
Lhbp383pRpP5fUaudTxWJnDtlu/bAFctVjJvYjQyafy7BZkRomb+Zjpyi+e+9F5d
rAS54Op6T6azSAFtoyQOT8KJWbw6cn8pFKHXNzp5QMhDivi4jx4It+f3SGn/ZdIr
0TTQbhxjhOQqQbroSS51FYwrSwDSI7JL6EQArod+8oi/W5qqpZgngxTbDlBTytlU
so2NuNH0YGcq0nq2lHMmimMShLcP9o4030Hg8mrkvmW/6ehrifF84rEB+iJXlUQH
Ss2jC0cwAfOsLQYtIiBFJmYgpMBi+1l39FCjxMjCIPB8bj+A8LjRnfY53A57b8ru
X70NpaUbIvd7harU24miV450T4feqJ/Rr0QWs2+Wqdfy+/xSYO3Mjv60g85R3Z87
lK7jn9h+Cv6tukk5DHR9f3q9KgRvnRXL+FD+2JsxWTE8ZXgyYo5XU3aJPRHBKe4H
TWNaDP5LYePDS1OxrgpSjcqj97Jut+XK67LXVKGWv/N8L+iEJp0ihpL4XPBKpdEt
V17j9UjqMnktiNHbnfJP56mf2G+qI8Y4jbwdZEqP6qRzZ2S62R/Ty46vcqSDa5Ea
iv2P27d0gnLF207/JMEYlKqk4Y1D0VuB3VmEuDz9ZKDDvWrmyTKQ9lUiiLtz/QEp
fuZS5wYdLAJhn+76xbquT1CTu0d9vKeVOkykvx4GJ1Kipg2J3ojZMUInBLVB0RNO
x7f5FljEwOrd6iwnuYz7X7baFaOVmn4jjfjdMzSvD0klwOKDLWVcSSBmIyF+Hkq9
d/RtsxuH83Y+9m38R1zSUgBJ1DybTjgSf0EdglfzGI8Dl1oR55/UmP5pRQj+NHra
UZI6L3xutk7OUY9ftXlUWvoXdT6Gmfz6g3uy6rU9+AIfvxQJbvj9w0GnG5fDhzrO
+93Dn3MWOX9uPIfCgq4Jq/9VE6DfSJZ07C6HA+oOGVmO9J4UdnRmT9yi8aGctaqi
ixhNNcvutdfdWDD8O8NyHLa+o9Yd8aYpQ26Lhla5B3fadBqmXVmnU48Oms6Zbcr5
Fgwvbq+k/XJ/wnmgZPraA/lPPsqIVbwZvFsoMRC97TiobgNYw8Z+zPAJwcXzzXz3
SXHn4pyigRjYRzol4dXflRAcFvcvZPZZOCf9BgVw48h/sF55ahRIqTOsfSIFxPLz
SCIRizLAgBCmj9FQKswiixKt2RUOespS1RMkm5znzL0ZV+boGkqGMdLCqVovoscg
ktLaEF8ezKjvVP24AqF2HfQ4lE2jt0jA/nKgiX+j9t3bNORt8qWnNvvUFQHZPfv3
OqPIxp3a6nOCZbL59JJhByLimpaN+Spb6NpXdQTH55SjgCziJms61VYYYQyRFLaD
6VgB7siAoo0cAb/om2aJFTqFFmbn//IujAHvoVyPvUzABUTlT9wkiw4h0dYWSi4x
Mv5Jt6WFw1+Wre389tfvQXf6vj0KGR1RYI5ls7rJqWDQkMmGlL4GDvfICyQ8oMnZ
bCD5vAdw9RQ+vW7eMnaXYCjjkLkUGC1MHM00Xd/KXZQ+9r+4uDBVRk/K9ocBwYU7
EvRddx5tsg47r3GQ1WUcVt9qD3h15DaHd9nHEozxusmFiyUOm5LLLQptxawD51WB
OIKpzkcc0x8dxc88fiUqOJuoTgnAWCSjUG0mYWz8wDGeavav99Bb90FrSkYDIsGi
0l1dBtd0PkkBW69s4fFz/tGCg7QY9L1X0l9UQvj65xxmU05CTYSq+1LE8FHF72Sy
45882GEJ/f9OI7r26BSTCBKZcwoGhEGoB+LMZNIr1i3u6Pm9vwnnfVoDxkObQEPn
80XQb+5UTobYkcfXsb573JEdh2JV3IAR30i8cgtFdHctIjE77AgfrZLMzkKKTsaA
/pBrwkoKHQiyLGECcbYkj+qJWCwdDSuYYsCmcdJmWoOYrO9+Jx7vM4fBF4QP7fmR
Z9zX6wa7LYTQAAWF4Y7yTwWV2KgygLT66Wz6CFZsGVXjhpg+GLB3GlO79Bq8+UJc
bJAhoXWDmYcPVOGGsp43ULCphEWFo1qF158/ta280PE6ZYUtkLV2zf7aHFFQp+Aw
TKs/+hM6zv0jk5v/6o4fyrWLN+SgJAGw2tod04Y3npDE1do85jHMJC47JTm8B8iE
W5eOfRre60zLsSOdtjzwVfOhADJjoEkBijf/wsfRQNhIx5YKbZe3DDqgJvBZzLGt
DgeIo85uFQbh4ct5eESOstU0x/9Wgdz8M3NTu9UXilexe5p8ERyoA+CZ3uybXBKm
Nws+Ndgkr9iAtOw/FV94wc41KQe2jayMe+weWKUkg0xoCgQaa8+acuLyhjlbmtpk
Tw+gDuvhjKuLcjKXDQmUWdkq/Ngdb1ZUvo6i4+mnV5RsXA16QQ8fh9cLpHwrqMB5
Hoxc/XUlorFG1Lc3YRu/sfeutHovC8PMtfz04Va4wsUKJkbkdZ5wITVjq3v2lG7i
Fj3SoqZVHo2uyDmx66QVp1WNtmDUISfr5y+AJBN2MO4FOgOlVyO/0Cp9lYdjHAZF
wSpnDLesftrA5862jvsZzwDdBwEXlG4HJe5xaexq+4oAo+0EA/hvOGvR6/ynJAVd
fguDTyGK0xgSQlq/rtL1JneqCr6Q4d2Ek0Oidj6a08BYmA1QsomPelpgyQrYAuuc
5qTzrSFjo9tnalb2u4H65iY0gXRnBqtzT91WAd3YfqtSl+FhNNKBHHDNhPK+8kyg
+FfHqqhk+xhX5EqEfcfUe78KtWb/EzFkTM0hnpsG+hCUO/zPSCdVqUp5bJr4DjyN
c8rTmxSSlJuKF76uPM0bL3xJ3+sSEkc6j0PJXBTz6sFkMUmj4JjbCkE31P4pYbSk
tzU55uFegnf6ce83yMP7U+KrBiOhUozuF7KPtGoH6uqviIF5UJyqkG/iug3qlmD1
ikpJgdz+SXX+cp7ROo4238emYs0bUDVxgI3cgxRr5Etl6629Hpdrn8FwsyDelxPX
fA+ZdAlxdzW8/MgYTWrWQBu47Dsnvn8iU8n1yT/H9YnREIXdLlJs96b5cmB5Ac1q
66FEWNNWcT3+UIxrDQD1delKNmbwDyf56Co9JsvFAwyewfR84rgWW2znnaNNgD9z
f34PAVP1DQaakoltEcMB7uXO0Yd3Z47XqKt5TjZjdvhfNOCRrRXWNGNH5vkDbypq
v72qlCFY8vvI33Y47KzZxYZPdA+Li1yqmgXsmAHh5LvhgPOCvBv7DTUoMaauN5Ac
viDQYhMdp7DhExHoW4esk+FhFuaOJr/gE1lWrOGc4fvWXzahb/CopNu4eMWO/0W1
xdF5JCBtsW9ADZIOUhUYrfZYz1KMIMlLbxc+5FAydWAPCeTEQUgvc5RrdHLFRkdH
SKFc1N/7MYFLg9y143WMZ/Rcna5JfmoPo3nGnNDxxEWfZZi+T3T+WF619mR+sUTx
KvTvBIXiiktdq+E+8/CDa1Yb/cJ7wmWWJZt+Dq9onRgiZd03SuAmp9p/x2qYz9sP
mBrq1K6/AKTio7Gg+Uv/a3N9LSn34PrS41UOPxIyV2whiUMTK5z52wGaRWlkkHF0
BvZTf3d0emp6kL7zzO8wVpUiHM/u7aMvFUZ5ANzZgzoFxjvEYIxUjoOhBDtj2RGz
v4CfAFl1uZlwxNSCoJep4iUiGKhoG4xKKsfH6YaHBaYg2TWz3W0RwLz5OCdLnwIa
qwKJFHa9N3/Do4SJn7DofzIrQq8Dw9QkkRFINsjpdypoqIHWBgrXwmEtnVPa9qtt
xaYUQYkWawdISGvXRuXgCAjJMflxUDHAs0Usc1jOpuGCGF4eL/xCE+nVt/HZs0S7
evE871B/xjgKl6+/kDCNfK20vJYCd5zhlrbeSSJirzvcx9dPU14I0ntrFv3Zqitg
WnZ7IZfUH/s3CVQBZosyWcohL5Ig7RTjIwI56SOjRAgkkI0VjPtiaKDXACXaYuuN
pvxAtXElLYT+iSa5cB8ujY2tkpI+qGpmIoOEgzSkSoAO8IutbMeDhG3NZkqhJyQg
tRKNA9mLzSudq5LU04gbRKVh1YePgY4i6vQx3QsYe0stkftAUGJ/ACo32Gs8ErE8
ArNeVra9Y0KITB4R3j192Ya9SKsdykS7fb3So8dKw8ZC8DnG/sx6wsPJRkzuTLg2
z1MWTr3R5o9BYgY1SBzOsJJJxY21LRZvQCRF38kswA8HutNBC+Cg0YFfZc4LDYi9
1WehlKSbgYWjZbCmRlMHGLV8eRuVjsMVR5gw1Dvns/GSjb09X1SRe09S7fQ3KGnr
KOeD2vpgtohBn5ml6X112LGgdTG9qOrGgrUtX69WRzoHYUEzDLeawM2XmoaV5ZWv
iFJ4uzz8KotNemX4uPFUZBJcsCLkLGD1v8qtOAvHpxtkBBCvsgf4CjNhnnbplZ5p
cgo0k5zWCe3cVIHwbX1Y+8/lAgOkiMY6bpnPpOu4sXpCSAX+QL6pebmPla2a47Uv
5y1Xs2KL3ibWsYHk82WHge/vc2b/6K9lWH7r93Mmra9YPTWslSI3IjznnFUyg9kF
iAGUigk0+OzZG4DI0Uj9d6Yl5AO7Muw5hlCDN7ergJPfruhEq7MbkBF4AZA6pRWb
Fo65KxwT5XhU3HgV6B5y+D2WfSvXMH8h0ZLthFdvFhKDVioaNTX5AJ2ZiZIzOqe1
96imu9tKljfGgYKGa3lr1dMpwfuBrDgA11hI3OsXAVCSNmlCPjT34/4c5KtFltGe
R0Ki2M7Kn0PMG9ppWE1eJdX6YJNa8xVLn6IWICiRQCm3fpx4u+gtYa8NsPniC8NU
FR1/s/4U/9dBaupHJcyhrGtnFjbNZWw/8D7dYh6QWkwsxlcbaZIbpXFCnMPKJvMI
1yBMTVwutqG9j3XUaqOhHH8z8Huf/uL2UF04mrAe6LfcePXF7qarDkYhpbhqHtvP
Vd+Wnv0SZWee7ESLrwyzsQa6oBY+yDrJBZSu/IKM5XFI6+Tqu7mAW4suAJrSiysd
m/fLJ7Lz7J1UtVoQEmF/BdW9Tepnl9fZQ7BRaMJSOc2p/USjjQ/9iI5iToSHrtco
5j0LijKObrvgdNta31zzW9FRr8Ap3sgTkM85AfPxE0BARukIEsMdeTXByFFxKwWj
8nyN9NMR+SqQxRZdxAujKmsSZ3x6IMgxWrckG0VPaccf0mP2CnR+lb3xAoy7f6xh
DWyAaNIuzx6itoQHED4UkfPX8xDoafHy1Gay1rZe91D75Odx5H6WGQSWLn2KYXpz
/Byb2fPu7znVARdWcNvPEVu2J4pdomDqxmOVKhfRUMYtzXC+nMjVQ3VavkC0VpUl
AJxawPN5kfVdxWHu+6Hy9ljJ7ybLuY2tOe4+hTaG6YyTVCYYP94U8tJYNVMBMnM6
Fm86VycpSMlBCJPJ76eBzDcgYZWlQO3jV19gdmLmQjkR7Y/Z8fIeM1Na9N801Frg
p1NtRpXd7FLjrFqY1lJQEFP/CzyR2mYgTqAYwTR/tM8qaxHkaAc5wLKZv5vaWqlv
R0s6QHKZaxtMRdsF4KocubYiMtfFE+9TXWi40Fex3q6MU9bU4uWE29DF7wKbfMfu
6JFw9LYhMLJghC5oPWdGbbScb3eyhKPK3/X5BvCBInCe+FSldkfyNA2Y4ro4rpeI
jdvKi5ILflPxzHV4Xc63Gm9LSnA+6Sh9GDT9GDP8cYPp4MQoAstpmAyRuXpbHq1a
1pe6RnrabQcdbQwZWlHdAe9XifzccdLs08b0Kxcsne0h42mG1kJe6r+80P/9pEdm
C7S1Ymxxj123kUXr/q7zu75zYjo5LZT/Lmdho3JIxPgW0GhhIB4CGyY+Rutn6mwj
sLpHymGyGtV/6goVO+ccXdnxPQt7oDIX5f+kUti4ByTB6EgkJDQbjNgWFSd4VTKn
EXGkPOua9g3GYAZoMoQfAn6KFKyU/zVJirYip6H4zf2YHvgCtgazh+9o+NGzTcr5
qkbWdnHLJt1J92+s/qgH4+4cygv/RvoMISQfyKihfLCJgCEvG2XidGsEDqXoyito
P1C4GlYDjEqpU5d4JrCy13+Tl5ZExLwyJs+fiqNeV62Qttto6JGyTXSzq9FXy91y
+FD91r34WsAbyYkn1Sk40KfG4mVbxYjoz6+mtNbW5Ar61RNgy2MDDR9Ivx7XZ479
ZbGfWK3fuJEMj80DgW2EWQ6MyYWRlkFh+OPRTK2vFy8v3icOYsEbTdV+jKz2uZI6
xtwaE6439Hadoqcndlpt/hh3Pfy5/dCe3kPZtVciaW+GUluoxhQe8JMHtzyp8UaZ
m5I7FBLlA+K+cDNM/rXuIVaFU2v3X9BJr1rMG+W4YowK3r0AZih9lUfUc8YBJjrT
yTZoypjaaLGYoP2jVxC6LL4BeFv9luT3qE2IxrVUBbycCBcLOVeMGEP27smz13eT
9dzpvCO590o9THoy3oQPiOKDg5I44PQ6tGeGfdaLEqZOR5ZxAfGx7k10c132HXo0
JLPlX4GsE7VPi1wyc8z74QlNNqeT/tfRy8oUIy2b7ja8j8jCDC7L9iCt8ykJ2yyv
FpLDjrvdzpFrHhwNmxquU766B6Zundo/8NvMqnPbtT8ecESp5OIi50TKb1k2SrlK
jmby/f4WdGK0Xryage1uLrDgrSqi/OInRJ9Rdqgj/f5++3YmCtsdBFkud1m/cJFo
mG89fZFetEJqu9vire0BgmQs07A8rDhf6NPKXMqC92VaX2HbyZRZV5ws3GChbNSC
UvdY8HbycXfJI34ukAqOH3dRcau+k1iNBEwm7dU48e3LCaNppLokYI/n55qpA0PT
cAeVjrgD7LFzjWRt4V3cnUVaiW8rKPMAeZr5ICwcet8cyB1E1ZcYMA95LE7FaaxR
yzkq/LtO3gv5C/6Qf7m5lbGvOjLI8pI0v04EqSu4vBzwx42z+S/wcmaNfUEPLq0C
EsfYNLCW/HreuK7fJ+UXVkqjsC+k/fZbAhKfKFnDuEJRpPKwac92rhIvdgarZjbN
jczVR/cMItDajYkw8h9eJYP38X2rpMQFq/2FeiLxfeiYiCFZfBQNxpFIdAVmktRn
m86EknfM43Mx7NSHwu95LVpv5PYtPN9rT4i5PTjlpypxBrut+7nYqapgykVAUvAU
y+2BquUAoAlAk4KuBlOSvJtgIZplidzmVrrCIdkFYp8dvxPFNzeY+5e7yl5bT+RU
rPYiOPSb54UVJiKkMRaclohYIj88bUQodIZOATbL9o4m9lSaEYUczaT4OCI+ePKq
JH6aEOl7XzECEOIy1BSFWvcCg0IOK4nW8KXSKKFdM6uuyZGPq9aY5l09RvXwuaUe
7h7CwFu/sJMTiFTmCAQOBePnO9nulryZkwvoIZpeFGsVwcg62ZCHXfuEXM376J6P
N0f1CxkXD4ZF9xrY+cmbGztgUlCirQPXARDuTIAtkBGRIppUTFk3gs7nvvsUHQI0
NQjBKEaMYhaAOyqHYFJnYvRK83bK9rGF30M+LIzM1pVBzwkmJIYOFJPTQcxYprrH
I2rYSak839RDQ9UfGoOER2HRAs2qxn2Evowd0xEjbBJUy91qs+1v5RR9Whr1t1+6
AUdfvhK0CSz/srAfo6B7lSk7YzPMJJM3IlDEisIpxTPxhP5pCaaYIVr+zBofUNkO
fxi32b10SF/mP/7wd8XmJMmoYJzSaY0ky2LFS03c1fZpp8T/WqUMiXj3HC748ZDh
rw8/ZHKdQ5blL8vsnLAjBsZr2AkIs8g1SCr8ymT2Ydz9IYTjOk1fLnF71Frqk86O
wwvNDs/rSUzPD8DpU1zt9oagtMMAHOQMIfhYczkyO/bYrjRSdM8TeO9WJW5PG41x
hffHa7vZzAX5/Sf8tEtydSwqppmT0ErtlRrd5If4xiPLbAuPlTvngPzFIvBt1D1r
hfQFtf2pCCVO8BxzxxCl/FCkOquxZ18OO/Q+0+Y0FwpYKHan3x9f8sCSXg2PeIEs
kGy0dWsZQ+d1sw4ae/xqRjKHPtpPQTND4GOYem5/uWkQix25Ttc2MIisTS1/bY9w
WSwuhYYSFqjaS1rZU0kSCELDIiUShwFwRcT+dh4pkM1hj3UOYutBmQoCx0tL3mHk
VsxrdIR3/RIEeBzskQpJiL+OMMtSH9vTkTdW5tRlzfr3CYxU6tI5DWsTcG+Pwjv4
UMsYgq8S4pk6qArF/9Z8wls9Kcppu8lOSmueZpMjLTHwsDteYZL2J5pfUOlM+B4o
jN+/Za8+/SBTWs+OhC7OiTSlmEWjtjbQRMu/A9Xg7NJ+zTBA2rjevmNCBhkJhodv
cJRHpMU3A3yXonccw+D865WNQB3p2WWhCnwSuQhrXiJAri2zTF38KcMQZjsXAh3m
2CmnZU1JxA9R0OJbsMmygaEKW7Q08eeaYdbqi/4fFAE5vUHvnqcL0XrdPns3vNyy
4T7v2tT3KFyAZn6nxpVi0/uBmvOSAOx3Q+ZtllD6OpbjRkVBesoxrrTwBmpQQTS5
dbedAs5KGdMOl59jCf1YNrJQPY/E5I1IU6DAC1452AsgfynLQmzf7WOmM8hF1U5N
/ic7BIWOd4fXC6J2HkEwfmIZ/npFy9NuNo4lGXppGPwPI+4ds6c5UFTexz4m9fBn
muqWoJG9MelMPCIu0+FpMFeh6E7nvo1SEzgt+Stob20ab3MX5K5C/BgJoG6vzvim
WfJh6H3MD5/zbmmNGY/qrAYolRa7AKN2OFNF4zW7FVHD51ZntjO/7Yotjjm6qMIi
lHJnup49Evfct0WW994R2u4baSBmVUkIka3o9Ngfv/cKgX5jwoQjFnaSuGtu53GF
i4tYL6OEHPJq/6BizbgTrl9fcvgkFkHIhiJ5GTsN+e7c+AHYYf2Eq+MR5G6iNDbz
TK+V64LwzkEU+2RqULQD6ULdutzZI68tFEf6wzOfsumbPAz9JrHRG0Vw2a8wL3oP
R36vexvI3i5zbIdGS3SIyfMAdZ0RU4NV3iKOdLGO3rnvdPmOcE32JAb4QG/uhiB5
XNEiChrWuLuVX1g1r0AAf6oMCngcqsMitxR9nd0RAgAJUUZIxAzryFt0XV7F5mf6
N2OQVmN82HHWSL56t/wli8h/lZv5GegUL5ma5rnr0A8OI+up5CDtqubIHmR3Ub4Z
kiR+hvM1ClHNlwZ/mJz9nxqzVy+68/21X7ZWKwUw8GgM8lINGyaG37kvQG4bPwuL
+wh+e0t4D5lFyxsAJ7bQJrN8Yftf9FRoFU2G6kIP+uQzni6qm+eqr7G0IyOKOQt3
5tma8CYoYpxsybss9KA74Q7+BLadflEPcevTAUSpfreGSU8OMMK2lEo+7IMNt8lH
Qn/4dPkCh9KSMF9aFv9wxKngtnmSS/1+7FbR0GjV5o4GI0GvtXj+s4xQzlEdFglO
da3QnA5P027wtHqyA4ZmMHK/Q1dejGUcCOcY6cXwED6VrodJW1viRKXM7xGckinZ
snTlq4u8w9NA/BpzLETXcvRiGWEGvKBnzSEpsLAlJXV8XFFdkX9i78m6A0LLy1WQ
TNx3LwFTOKGOJ5s94LYfn4AJFmndZMSoculb9p/a/mYmZicfn5c9ICE51a1lyXWM
vnd9dZasGLnM4G4zU41WslH1x9ZVXBY8qWuB2vrXHQDMJzAKi61Q6a9cxFP7fiox
C3BQzWgYgHFxpazVkY3LzCs0CTLqqXk+79qABpzNWpGMB65psomPeE/QpE2Tay0u
8duroE/RDhbjkzzkC3rcK8lXjK/8t2WLA3uCtNbWglpUZsziHGhgESuG+iDvKCFU
jIeqbPyRz5C7oORURgqApGFwNCD/Zon6oEire2hIhax3sXVcUaWKDMfS+BOMfHCw
RB/zGl+2DQFXj8Sauc687L45vGzFnBgt9W5zMH/eUegKjBCFHnC698398BTjG9OD
StGndIKHj0HYYgZQxxLWwQEXK01Zp9iDonkf0o472VoroYj0xffZLCajIPn/Nqrt
iagJFYdqQmatwQrjLxBZ+Hj669UyKUetPWvh9Gadh+lATpagwoJ1/Xc3dicc7REI
nXEdS5wv+4SooWukGsrMtjB7S5+5LQr8/KuKHzayDe4lmushi1/UeggI3UaulzFg
0Xde9jW7fMBt1q5iWvB6GsNs5Mf4eDRGQwsYeDDoIRIhlZCbTCmv5gGz9XXjarux
ZzOa7YPaPfJQi1HBYX1sXU/a9ST6ru64g+HpCwwDC87l7XJHcmSlLVU22zQAzmll
dmK2qWfZghdGkq31y9VNcEzlcTzws2gg5rTBoC686qHNfTh7QV9Vqi2d2gdKO80N
PdknXxw2EwRHy81/8EzBAgipQcjU3+vYhtsLSEVg7jcM/omwK95kDEa8gPAitARf
J8NNCYnfwH0/QM7JANyOOBFUtagHoqgFTyezsy3sLoAJVlgdyNV9Vvyzruj8Q9/B
UvoyhlLQ+AAYxlRnySZAR76Rj3BhoWonZPtM3HvyEsU9lae+rW4X/MTOsc3sKix6
3rftxgLrwKTOoUJRwMC8jFmdCGVOH167FyWOWkjquqDzIbTZ5nY/0vjlM3fLx6mn
SGzqWwHA6ltwYoYOQO0t2GZqqKNRg8fcv0biVHiPtMLqUTnRo15MYw4LYcM/SgN3
FeGLo2ZJqRdgGY/IP8R0d20krFFvMVRlTJGi1BNCQzw4NHgZA8sktTlCPxTjjF6p
JgetSiSkZ7WfkGUMj0B6JJgMfS+M5nFIWxoM25cmrgWoqwS+VUW4KhvY8q/8+oAs
LwY2ToEHFmc58jZwKy74xxiAFCpt+4VoIWuUc8NB5X9MKA1XNsc+0zKbCGtGPj9E
rDdc6sGYOXlYAtx6wDVNVlGy2/UqpbynRCvwTbJbsPSRWmwXF2/j+Oh20GLSW5Z8
1xLsbGEz68JQ/F+B3yQ+Qr6qn1Hlf9McOKjYNsZRv45TT29/d0HNzho4ptja7+d6
lTkdHdT3PR/kNYY6WVWjzp7xLFmBIuNlY31o7EQxlJGlwEXMfnGk6fC4W5ZW23UX
KxSNaRueVoOEeqbPdDvr88ZWcG7Pg3grzG8TdLBvpiouncn3ZQAc2zh/rkSqGM2h
J6OoAZRxyJl83cxlvOC+6RQuEJdAINu8Dle3fua7sMu9Rr5zonhFxEcfNuWuys04
3WD5MWY5imBXGmSbhCO1C662t2ZV8uigmwL8GgcHT5VPnQRbMmiMHQ/Zfj85gPLl
u0hSB5JeLwg1Mi3vznGL40W/i36NPgmohTzG83wHYwIpniW+RE4tHWZAOOtxb/FH
dXPbFoLquVCfmzcIXxg/vQv4kapwZaUHQrkqV3o6h08lGfi35qXWNx8ivezD4SJI
y9HNbGr2bH5pi81s/txKxmAh2ScdT4hi3rjJpov+xTWb7K7NIhVvPlXW1mtQraEW
eWx9CR4kdXTMbV1BmRgY+xcj+rsA0C6O6QXI4YUMqFQ9xqA3gbLqyeDlkhNb1dGw
+wNUFnkPm20FGO+QQo9dDf8KC4r6/RmZEgyhhvOCU5XhAeLUwXAPYpnVEigA8Hkk
Z2+pU5g1w3ulVwlb10tcdXbEWGKEdksSpYojuPK5Sz0h8plftIfhLJlCqGaEXVni
2+gQyhGpGinyyXhipfMAe0icIVwvSdFZOiqljMYVcouut0Owq9JvD/yvLsyy0k5Y
Kg51KbnfbQ1mBoaQUGUsypvN0jfCj5iYKx9038yjRk8ppQ2IslRSwYZwRz7b2xlX
O35TQrM+o3Kc+NdgjSXfyLC/m8d6k9koIiGVRIGKP8iiRkqm1Gw/jM2l++w4Kosx
Oaz0d6BuQHyvosfVnyOg4Xyd84kZDGwHoLU+jfB34R0p2HRNtz7LGD7hNnYHmuaI
QcsrK3rtGw8F8n/jjFFPTTvMKH9TaKt2BcQ2btV0XpLUNoiTCIMTEGj0DqeEgWpP
JuCBFxNCfcQkHhdyczrCmbi7TJpb4Dab3e1ceqGvrFu2/5AplBuUHPHM/mH9CqpP
bkeCGYaTwfQGpO8aR6siJR3DJ7BzTJGUGgxE760uPFLT4xeeXhNeJV8cXeouX+5n
4ds52AOdmyjhmGckon7Pqnfsdky67r/kD/13KS6G/aXMhHKNeQO6FSN3xFihs9fr
z7XC1fFdIqnjiCZblt0XG+6Ps2IYL6zIB77SywCyPsnYcFh0noxGm9S/psfBk1QP
ETDFT/R/Xz5utMqhMx/vXOO2T9JrhjO29tUQQEVkjlzADFhrBMO58Bnd/CdaiXfQ
YsKrIN+GKpz5xIIUGif3jPQd7dh7s5iRTTPrS0yVPyHg55NknUhIZyDyMUmkuuwG
qaL+GhBgpqdIfs4QVWAFp2HU+rlx4dCHhUqWjyYd0M0HADdET0N+ndjVOOwiBpo0
et57fWkgy6yOWSFDDRVJ+SBZ2hA+NQTsyCSN+AF/AA3WBeZAorD34dElC8lc7m2G
e5+GaBd1KZU2X2RVwFtYjXz+0agcdAgO9ZKr8I6ETGL6gTxQ/CfIi8b7mfehh9KC
PPv+6bvE4jrtCSEklBzhlPvEhIEg233I9pCr16hMkr+ZYvY1bxdImO+DB03ea+6L
UilyC51UZB3UazsQJKp0ULkPnMqAMeddIMTZv9Cr6yVldauGWnQ5hR5gDnPyD00T
v3fwnelyfSDTPZ2vzi988qeixn8FMYKHaoksoU8U9sz5dCTKUIBTM76dFtIKcYlN
KtA7n1qxf/awCQ/eVLZw3s9z19dtMBS4eBgULZI4ufW+2RCL3YPuvEXjTYN73cQv
KQQR2fQvynkso8oq/9SBHf6esxbgeipI9v1srMjAiGkpeHN5u5noZ++2noENhq1S
geB1Lvv6kKoXD7qhKVBViquwbLJBR0t9X6X2NsXo42MlRHN83XVKZetHH6jOXof+
9+NJrZhHVRfBCK53u9c+qlZZCWXKJS97Y/qC37Hw9FkuM9gYzwqMTiYmNV16vGa7
ATALaNgyJBEB/qevaeXQqW65Q6hfia+uBs8h7V8bYkBuaMhpE8NUffwjvAKoO6A6
xNR2+9Dcxgvtnp74fCewUAy2o7dMWBENZ3AYorI/IpH+KH6PE1rDbSxikwsjXmnF
z9ABgfyU5IiljvE2kXeOH/HLcWFannAuocGdwBYUsJNZXchhFGrjlC7fWYCNt/Py
HUe9jUbBYHGP6IBgbw11mZpUHufvS17Nx/MQeQMSFO1E+CX4Dzsb9JOscBERPkZE
VF0wzE/69tlNWQfJMMl2ZwA0pUy2XZZqh8SivXdw2qzS2y0tZAefMpiKH4QwVwWc
LLk0TWqGLBV9GenkMjIaLazRIK5e+jDPs/jhLySKPJmRSW4/82XkZbr4c3iKrIPh
2HLhshxCSW6BgzMyRdaKvNYhih/dJe3e5WpZB7bLPISrTLJ1OWt5M+40cA/arZwM
ynXbf+L5S40UMGM8Of/7w96OWVa2O5HjpJRVQR+VLcnoaki7xb0JJ8Bbv9QPR4yH
V2WsI6+eTbIrKmSOMiYW2ZmMboe7YK8/dd/276dyd5v1quN3mXP+ahFoLOtZn/cV
FJf84iMFUCo7DL9+rM6gXtWNXQGYk8CZlt85F/lZECK68Ny+iQ+B5j7PBeEBjGeW
hWWggGvOjLOBIIwWWfLysC3TrfxoHpE5L1TYZMugMIxbOl/LkLBgg7uA6QDwetyq
ztaLpvr9oETHLttUIvF6H80hHZYHu7nWwmphOT9AeA9SLDkV90D34GDmjw1rKpr3
pxnQCfpXkKomMUK5j9tZ2j5aBgvfhRPb84QjrdVLvboye28KgMTYlg7X2Hkt2AcH
X3SR2Ts0zu4W1X9ypqaC18DZipafsHmiV/csFujgsOrXLr84dK9nJut+KxSYn2xk
qTBtGnKmKrqTgqDnHhJwIjzllhkrIMQ4/RN2EAmSabf+GwUerHsqMCwWjygabX3T
HAHgpC5ls3kcCVsCdtgAdALXl/8xBEijFnQImPyI6mzfOyLsSIElBf3QNcPwZFlp
NX3+JX3gm/uuSXQIbS/cthfT8Csw1zPS6CnqCDuD27rR/PBUdwfqLPxYSOQOioGt
HztV1wh/mQxU9RuTuZPz87LyV1CRz08F+X018Ezp6y/PzRx1jJ2kmVCbAfAV0AuS
zsXf+FlhvirvHLDhvgXOnp5M0VOxkheifwsR24tQ1ZZLIpMSfUVuFLJjef3Kt2lF
5UKcNzJ1WD4P9EBHgaRBIImvhMDJ77OpINCB3wzBsAE/0YM+U1iU7WHjhPJfZGzY
y4qO40y7a/DCVzAOTKu8TOQwderZrUyOah7tBoqaB+1hlQmejkaw0BYvedyANAaW
dnLaIKOcr8DLySYFtpNxkZ+gCpTyf89e3ZGSV/QwNxddjf9ljGT8bzzXV7ecQO9z
2c4vsZay8/BWkVr+eg6MttgygFLSzaVqN7y/srczgSHOBD+ye+AR2C6GjgkuLIEG
EYDWaOONLqSL8NCUFCHHZ4MhpF317cCXR+bf49Q+iy/QJFhhrlq7BXK0qnbxqiT3
w4bz5oictnb+8dCXm+W6fSOrwAr9K6SksPXLoYjULuhTGS9bU8BZl0fDkFimB23s
yP2e+UkyWFYpT6z5+gTkg/Pday05kIbQjAjiZcytIc09S8ZsZQwXxbokK/GtdwpP
MQpIbUTlHmYc2OFxQMMIcGTQ4qjdee9u44PRCrG47VPlt6+S0TBcbJRWiUX16wob
d8p9WyvvT9uljQgSvOJMIPKuOBcAdlKfeN5fpst7BP8bYLvAuKIuvsAK8GCGf1db
x72UvXFIhBOAXNKJBNHOGHW6fvZ8bIvCEMkLeNycIFUk13BfUpufk92M5tcFLcgD
fYeUDLYkrJ6+rnr2XGjZH+2w//lS862mGelQuBU8HYBkMPfwmUE+ipBX2j5javXP
PosecEC9KifsBmgeMdRyAznJ0SUXNp83j8gQHtRRBWd3jIzcGcuKY9uLKiEcXHiD
yl6BC494TPh5bm1cIy7LdZtUNoqVYnX13i5FIWVGMe0EkNYApYI/NEwZbCl6ED0i
2pEMPoQpOFSXWNSSO/+5orJ3jMTQ3XC+iUulyoz3HTs7xvNpB/emMB8Z+G5KNcP1
v0R+Hc17hHKr3NV8myn45OyxHQ1aaq8eyMmzNod3MWmtFxcEIC0TntVBZyyEc4Fn
ffWPJMDrFVMJXcdr1okOj7NA2In4k8xZOLrGxYZ5CMDFasFCcCHWe2l37yRh3eyb
7MQwlXySOzDhfqG3GU5CCgnsBi4F8ti8J6qaiVIiHPIf4q4M+x9tn4qYz20G29T7
Zu5BYy4x2CpFvYnlEOeVGDl5sIbWum+cZQad9EETsbNnTUs9IBYAjXoYSRwZhtJy
a+lKdXk09jTKTEn/lByg4AvYRwFD1vjpvldMuGisXhWsIclHlqIkdUKnqwroXDSI
cnIanSxwZw1rejEItS9hqww04UZS0ZekTf124QE6ZIgW2eCFyyf7xZi9NMAMH3lZ
S8fmObjtZmnGt1e/W4tCJEe4FuS4jXFayDjH1DuBeGnn7F3Blwa5UPHwr87jdeU8
gZHTHDXsXqY48gXylZZWduk1LYF0P6X0cOpuafnmMbHi0MaynBRAyV0s2GZ+LVsq
tOS1PUcOQrG4pcFjYrfPYHefF6eYZ73nFsHzVpFaGizMQlhKh7uJ0MSJfcMMrm3h
0c8U28eMRS9Uz+o3XWm4B1bAuPPme5+aAArUkUKOfAFz5wZDgctBgMFNhJ/KiFSx
9duBZ9PO3DPV1BkVq6u9lYviN5bHzc9X2qvmLQIZGY3UM78rsRUr+sH9NGiDBFj4
cGNdu1sHNtCQW5fpiwFY6CHFv0gH7DCuIuhkudRZ2RAyJ+f6Zt6ulJ0jEM2k7xTF
r6XoJhqQ3sKFU1g70HhqB0TPuEP9xMqzHxSnBWHfLlqH4QJYm//t7c1I/v1W7eMy
7Yn5fj3+G25IeiFYF4Ja0ziGBZ//Mzjk7XvB01T+Xsm9WHpdMzRKqlFqzUkY5NSF
KN0sxS1g89Za5Wu0cmsDZZojNeYzOYGrMAq+OvZmRe0WtXozGvb5EA8XljdV/Aob
DSCtn+01y1q1KgREDBsHPp71XjwaqtZ4/20iNfftbltoOiGTjhDYP3zomEURPtrK
VFuvwYMO+spaTMgEA+WZ8izZc1RllojcUK58oDPpTbqqW/hWe6mQVjRGel1cUs82
yY0pqUvvX5kX9RMXwBJWSt6i6MuBLjAMJ1sik7W3gUotK0CDW6V3wI02b+yTA299
FEukiNKvSl7VN6yOjOiCUHXisw+Wt+Tm23wEdeb4EAQWTtHkQCwItfPN1Ah5cfv/
PbRKQx6QU+lJeFKPdDdkecg+7bL+rWn9niP+Z98IYe4rOWR4S4MQSqVhFhZP64MM
hGQQE2/4qZOx6GWkemRrZLYwK8ggYK38K8HfPWSFdIPjlRRi6rE+XP0vJhzPWl+F
ayPSesNnLXGmT8muSrdPSFG815kCPv9phHNGdRpj9C5cgi+R9j8oCmKUVR+CturM
A0VFz+awS5fMUTLfQZ1TB/bDZTVm6jXLM2YVQyEjnFV9Y37U+2icQyg/Gc+wyx5Y
VvcdFayXZt5Vyfg6jgsQXfxFf4oAY5HmC42+AXTZj0T84gyFhUtDO8fOud+qwVaY
EtolxS7Moo+PKXPeJxLLuNRTg58CwuUCCMOs+koSGS8KNSlXm8JM2ebkm4pOdosY
bm8pYSCOCmZ3tDPA0un7gUHM2ZbdIZ+Gu1SkKLW0urfgdqevCrtrVAmCeqvkc8O3
6CEpk6ZtlsrBqCttMgZcikzu+SYoMX7HR8kY7rez3I6jLLhwNAn47cLOCRKTRQ6z
SNXS+r2afQtdMzmV+S8WAw3OzgU+bJBvNEA/SMseRHF0eQOOPCIYEsq2BlZa2+/F
h0jrKheFjG7YcyAxBdAa7A05EnS2HrQmP3Lm80LYVUgEZ+rSR+MmxH4/vu1xiZJP
xK8Tfnc1HJ+QJW/i8v1RDshg+3ZBDgRn0qSRYq8sXQQfD+aI+bL8y54TqkF+aEP8
bPl6XAu0UNdI+d+QEf8vmOwS6N9uTlFzz0tkkbhQRtjmv957+1i99zRMyfOj0KBS
8NZ+HljSzQHe9qDHTBovHALqZWZQZjD/R984vDohc6dXlpeAwjGDJjQpmJzp18Gl
V9pbmqr6GVHsmH/Wj0WixvwiKvFr47lt6DElPquDW3pwJqVuAL67vzl4vygdOpdx
d3BRRxvGRvF0fwxKcK/CSIPhZw5TI++cr3Wepn0C/YbqKjMmEOg3/OjFgjYbEfDO
Ex27AkaGb70g1kAd3WPlE5U7hZLxgJeFQZz+C0S+vn/CU6u7YW0Wh3D7ksGjcLa0
ovK7KhASPp3rPpFa+wKt43V6QzPlWZoKk/UiO0/RUk/gkIcpPxURuiWEyh1DvV4G
j3Gz/a8qc8a5E0GU7AmidGi5ppyNVY4EameBIamU3+sXNJIRNi6huyK906bD7ipP
V3rupgOJmU8PCHlO9RJvDm0VcOOOaGTsIqOgFAzwik5pXMmh0HCgSWK1Sz+PiNts
4W3wc429joqAQHgrPYE7Hr8EyLkP7aEdZiOFwQ82TbI1tRCWkffBDXtlmkzqcLvq
baWgSPYXUjMf1KtCPHWW3epMxqjnP45qxUzVuOkSpmlValjUhhSwtDQqco6ZCo0V
PoiSXAOiVJtU3BbEEQu7hyRUTA/3ZhIgxp8kkBUnBCZexlkqJcN4r6RfHxhSZL7N
GL6HAZBDMo7af/J0VriPquqSi6Alj3NuNB7AjVJUyHJqDDWLQSOjnLLrE0qGAM6w
drYF/RUIYn3Z8UM1TJfkiMKwVt+2aOzw0UHB2qtwxf1LLmh+KJUiXK2Vtspx1zUU
kIK02dUPSUTLIbeMn7XYEajhSwbsM3r/1vty6ordWnKB6+ZJOOlUlcr90aSFLQAT
gTrPfWY0FiAP0w6tWEE+YDOQeIVkE6sZXASQGPOyRCuN0T1RJLpxyXTbWM9pgdBK
RUbDCRbw3qxCSoiK2rftNlB8KymfhcUquM02aZWd6fnKxm2LXJYGznP9sv3KDB0N
ADCAk4k7UNaCppJQyroBCpSTWaSw/YQe0XlNSHcihylLD0QkZLz40Ml9ivum6aQG
HJJcTEskQUXyv4xy3LLXWz2w5YC70/GJ/7uHTS5LeCbmAws0yj3aJvROtP197fj+
4IsaamSF/vvNkR0R5gA4hwBCcx7B7Ls5L2uPzrcEq+OtAAZjvJ5qfp63LRamPcM5
iR2MhP7LQ+ZqwpSMsJ5CEPMMgGendDW++Rn6m3mIAp5gX0bPwBHs7iKdNCaRXjvT
csLh99fmgDJaKQztPmXyqHh9dxw50AWHkF7fTtVAxEWBZLzrk0dggyiDKERhp1n0
5VBEYKE4qY8gdkywYcAOrNeOq7BN2LB6tV3eHV1gmgDQp3nYPxpHgDyyxVDZmFld
lXg+CPZoPoP6wTe02/saP3NShKcKz+h1bpjJVtpJp5SsLyO3DQnyc2Qs73hIMojl
hTHpADxMoAKyYbH2o8z7ESg/6NZGLcuGIJxooBPnBPWUxnDKnqedq8mxHwy1qfK/
WWHo9xNrrZUXGQAeM7NVQg+hpOn9jYhzdMbrDYazM3pWk/hgga6bvprl7mTQG1qe
5Cd7j1z2npkFpNaBkeHHCnkM7m5ok+YLrZqCPhuTHX61pytP0flZycTIYP2M9uCy
D4tBaGNmervnR0aZpQovZpVvz9PxGg9tLK64OAslBhFKSWD+GqNYWrmTSFyWzejL
l7KlkRDDGGwEFRPIS/ZYmnWvy22MH05fX8G3o8IBI2UcnXB83lnBMN5g/uAlswXc
2ev9ExYb8jRosiLNWWQhLN/ApZtQJxOLE0HCqJalInR5rfvBIH4yK1ssm6MR35ae
7OmS8NyDkARwKDI9YqG9lULh1LBp3JeWNNh8kuuut2SFtuafL+om+myvschXlxmH
X6UbUT1/NGKWLjxm9PMEEE7gt0/ei5QuHIXiKz3GuKnB84TgFs/yTgWHVcikSbtM
+Phv9ymK+MFxsKn9nRDiy3bboXNvhzw+BbfdEjj+4mBWEVeylO3IX0z8Ur0yrtO8
f4klZY/vK4Wd1ANQB+5ASDqxDpIwGJ1EAYj57D9qowgkgR7HZzD5GslW7d1a35wu
MV2hQtVKwyloy0+b8nUlvBymV814ZwbN38pWKtjaqbYjkokVmyjFzPOHhqEUc3UD
1zf9Y5/ynMDl7kZA4VT6UnlvSGKrw4YZRwI/HKe1piXwjYHYm/WKgOmN1Pwr1p3g
jlO6yKtZZvEDz34cqZguREcMPo5/N7NirHLoDAcw5vZmlIqMoUPSahNoHbbGqeJT
o1zTCxeiLhQcKZw3B9Sf7Yeux22Gbz4/ACTtjABQeAh38bAhZCGxudC7slMpWey2
sEluGwPVP3K0h3Becj3+ov8P7KAqscDUw6gn0RczG2lLSCkpm5gslMzKRMaTacx6
BU0xww6JY/KvWtL+L5lIYg1LqzW75eDFdOu45JuXCgEw7HPbBXkNArdiZwtcajde
6S5tfBYplbiSLYZaU62peGW+NFi1IWw7MNLuvRxDNXxH7F/Dct9sHEgZ0dRdPFnq
U3PvXOG25+RItaBRLHkWhKH5QQu7PV55M0rWmU+BQVew1dVa9N2Blf23wDfBJPK5
onnL/U98kuG9xuDznFP5q53hyUYD/MA4PxDK1CFRnQCHJL1Xs16AI5pj8+Sl1xXx
1zf4YCpdQxkRLDtRfeIYLPNKsPAoJkRm2W/3Q1idmg5Q0en4DjynP63YlhujGDFe
63ox38mY2FJgrhm5yBLKtcRS5tdYKqiVCa9y3o1DyXYIXR9jbuye27IiA7HDU3ME
ZIlX4ak9yRPdhOjy4ifCJfTf3iDBQQ9sY9V/LAMoR5oPSyhl/mVA8RnpJfVU2LN9
2p+4VidJldAsBQRmgkrFJhS9c/kLM7JAaghCvwJ3qAvoAWzMbFz+/ArkjJXWluV0
RwETItONIKmoagl0Nh8AhbqXiKmznhBen5ifzOFTpR6eF4CGpXgpse4F7sYEydwF
Q5LneYUFo5bFc25UmBCyik9YuFOqDUcOgdw6yAAwGpkCOAXQUhBPxX6QQigs1j33
Fv9DEEJ6koPgvGvoKgvg18zXmFyxQQcW2uoeHMGlrzS2wAxNHMJyxR9akyfageqN
vqJNx0Rx2OR7DvbKMbljhhsvNCWgNH/G/m1JNA+OedvUKp+MiJPJUeFO/B1tpCOI
Hm3/KgfS4ktIcih0Y9uq/Gx9qm4kZReIYA/hKv1QYFzu2lAea2Xk7pZO6QMqebYQ
DuGLQBEfW2d95VOgIExDcX0YhMX0d7fxeQmhN4srb68UnuWsuF5nr76Mq8VFq3BP
yD/O3PxDR9HmN52Z8iLlmowkOnD8nkfiimpIga5DfGZt2tz7QYYV2TDdn3tc/ZtX
qPVvNoBoP6Vm8IkwWL2mPmnOcRnWcNhfNc9XaoetSeQv+7F3ur+eobegp4TAJJ4Y
fYYgKSRj6ZNOW6szOedzCb7zWT1PBmaH1i4bxPonqF5klSxI6EnvZwGCpOsJv00f
ONylkmEN4nK2zcnTB9XfGDkQPW6K6pZzRxyAMp7DrpNq4KCHrrB5EXsNj4a3aKlc
/HvA48g92LwcsNnH9q6KvcsUXC5/W2cZSmDQGZrNCV0EO+gc96kOcAnswXEZHaYC
ccyzfV865ppkcxyLfVSi0itQ8V/5+6rz5cPBaI7iTNJ6fY+e+enoFxJVn6NRwTpd
IOurmQMlSKTBaJ67Na9EsR9K6SE11JV5UW3J8HpTruA49ycVjJvxYkr7SuP9KYKt
9F11/5pjr8PdBpmfLUR5vkajHFGtw53XS/8w+wKlMoiUqv72xKZaePSRcxkRH8Nz
EvQtscY0SfZD4c4Rlxx9g7IfwrbWKevZMIlBwHGWHyiRpOZC15ugRjhOqeUBwm2f
YnE4c8UzOjNzC2ZGbZwtrM4712oSgGHCtENljYo0BGOTGO/kpD3YyzgvoZHakJyS
J+vnUpjaS/39sk6H7LPxiiz2iFiHTG214e+jiDufvsi00RBbrJcgxR6/X/91vbnC
yIJUBKNEcY89/k5PnF1iPaYqPpg/dNqmsDXR3NonCIFFTOUSFdjY65oTbqfRzOiU
9kw0oO4x4C31zcvKBc4CEdZbemZUcjVilDaG69/isfnfs8W/JTjUSSZ+nNT1Ol0E
XPGxu0owKYEM1pFz2qVpKUU6GRShz/ioD59FQiRLZVBHJpoJTTiP8K5w5pXEWyVz
iK98BKhjnAJxl0sry4eQAazKTQi95RwoKW2Lm+kcIDSs4K9CslbMuNGapQy6LP2F
jqO/hriWlYptXNF0VXbkjJjolxh+Gr71nHXX/VVpc3IW4ql6IbffMbg0ftgfRgHy
NBqHWOUmfNJrNyFE05WKl40jM0wN7HmrhF22dGjyGkNXLzDhE5p0cjkn3Rbw3GV2
zQYUCAgJDBCapNjCQZwSN+W1tffLKxV2SkEUlQcPbcIlmplivfZg4VvEoT5hLj5x
4GNlSjIaUnDl8fgNOw4sSzExN7D5xDzZF0rpnSOtds8l6/4disFie7fkOq2dYQwl
VXswySOInHCos0uDyz+SX1Y8Ze7FPpR+cGPaCtKVcNGit+m9s6MZ1bT0vRRN3L5W
MpiICav+QV77nfIiuRK2/u5+tnobFmMj3l5K/mVXo8B6pYn12g9dLgAyQBf5xYkT
JfPEAsScuXNx3ckm8XMzB+/WCpSkbTMJPNRowO/ZkwrIibISRviyPHmPimo+OpSP
se5kdbyALrtf8RNkMpAG9kROxuMoZpmaKEDw9fMB5xGpImwJSoM74lCsslndhBWV
YbJqaNC6/CL9iO6iNpn71UGWJeey0IoMxllYceToSYBNh2Tddc4YrdpHm30FWDFq
TnIw7VSCW6j5kHMy2YzBs8Kjx9HmHZb9MTLzjNu6P9I4/iodNjwekruQHT08NIFh
2zItAJ8JMCGAthEGi4VOL16yrqSvpE73ugvZTJg0XHwE7vsn/m4KiaIRNMDA3YiJ
wrkZbqHFSnlJrktm5ixLqHEDwGQeRLPDAvkDigY7JjAlDbmVs7xJcgK/8G8hJsXM
sI49Ag7ixI1pDQHdQ9EvfjA2KqXbabK3GwOMQwZzdxkCScq2KN2y98uhkUKUpjUa
2g3ANajnH2vej77ssgr1lMvdfpEPtLdNE3thvYxMfx+AWSXN7jCpLfSBsf39lXf6
KnlN+VyQ7L2apHvIB48/MycBh0JAVrJgFacINjFSX91duzOELsZP3Ob6t+12Ghsz
Ogc3zCeXmZIClrFiJG7dG5h1XDRj7ZXsvQ+Elcz7TxNJ2CmZxJI5SILDvZpqr3WF
WyNXRDnycJ9n31WVGGwG0btx7lhv74sFHYM3v75Fbrvt8iWAq/TVEl2It6+qxvYE
lha3zRdHkRxyFDTmY3/MH8pOwrT5WF+PXi/aaQgduQoLe9Bew75hANoisnItyk9d
7tF3fAKUDZOM1oZqtPtgZyxrstqNVZz9XuqLkhF0KuxyL861BzDCG/TBvvv55Qvf
fSDZF4U9crbshmPE+megJEbk6qj2HdSvhqvqzgAUVOnQ9SZDYM+OavQjnn0ZYnq4
+NoqnBkDNKmoAiHpMrTsC5mhSy6r88/kF57eAS7evVXWjso1YNDHidlTftXEMZst
C+C5PxMFrXkMtZjE5xhuxZnNtuhpKXsrDV6dOY4zv4LlV7eKMbfG+ugrCGHiynFH
qKAQI13lm78Yn01ZrITaeAMnJn1VZRAKLufBesGEMtPqZUbsbykltsUxAKAtNuyr
NwasoQV6NNtkmPrI6SJZO7MSdkhPOP8UMLAtiLWuaTTxTq3liUyQyEvu/4wEfyx2
eLqUUqrtgzFlRnuABzzBypAsISoa/ua8DV75DJp5cV2pQTtQiBqCUmEL+bgIUiKb
DqLI/z5herYJFWSlenMltxyxmaA55DqyDEfshm1l6qLPwGf9SIZLIFpebsNwFUih
2HMCpJQkmhQxns33udrD/lmDqq2IZ4WJC4Vjns2TY9OPcK6doPb7sGi/jo7Ijv5Y
VocHKK81KPaDDwzdhtSk54IgbUNGSJbnV3B39paGC1WlgGOkyulJ1womDYBP1ZLX
xeKUp8965UsEMzCmADtAfhYI7P3kEvc3BMtJsGzxTVdtyJlUPOUuO0q4mhgFPhED
oCGeWwsz9m0JvmXCbBL9QnrhrjpH1LA5qTbRGK0wDmNZGz4rsh4bUCNBc5ISnnzS
Nz6mOEoimB/0yJohASS4owHfl/B+hla5ghybS69fO80w8NVB6AxXxJyJPcr6LK6e
Og51As9HnvvmplHiH04ziH70l0x2pIWo7OK+C+6TShNrinDcK3QGVfuB5jK40CdT
ddH0FT43OseoLRjZcEwm85NN7kG738kVZckLo5ulINvMKbSLckeFZU5grd4Bi1iA
LCyEeqIOOC9wCz46WDWvC/nzC3C4+SYfOazw/Cp4/LMq9ou3tuidRvFO7liGn6y4
bA/5OYInqVVe0inoikKgk4xpNJ3zbCFlNmIDoxBswv4Gmemk2VE/7IZJxgM0RwHm
+xQScYPuslk7AWssnvScj/TeH6eY5M/bvWdIY5R22IAC8tYhjt3jC8h54FWeZIZu
ux+3zvDTzbliCGU5iWxIi0xl0WTtIko0XryykaIqKuD3Bt0DV3VY48clrOIAlc/J
CZPHsZ18SVA+jxtoAwnrLhIR5RgMEEMGSlfl6x2hE0K4cp98CQZKTdCm1YrFQAQ0
9C4uARglIs7FueXUz64Vc6meCZhIa6VvfFKKAxn2HrjSOqrzHFkNdR1czj3UbAE9
om90eqaZY29z0WMnnpkVU6FAlZcDxkUY8VQmH237jpf6oQZwj/z9yK/dt9eauFnA
iToI3OW5wM3mNImIHrTZMHA1CLPI/s2peZ6mUAlJAl4RNAyk4zGaAYI4evdPV3N3
CZSD+tAEYmp5t1ffygJAwwKAVvJG8coxWQZMcHYxH98oMOCdoN9764UTPdUp9ofD
YWE7LER/mY7MXdzoeUT1Yh4Na9JzGvWROeghhhREHkYW2O8nWcjeI0SfTcUcK78E
iBJIGqil1hrsUGHfblQLUD3Cs3kxIBTyDnNFCS5FN59oQQRZYOp5hVvrQjlIeTEw
3DMQTcFvg9avhD1IrgR1gJ/omLJMFl0uH2HfINcmO+bium/M3yEy81aU2YCc+nMX
cmJOVfJaZjsv7sidwjdAkly/umE/dOC87zL9VHtRzOzDFGHqHUT/B3G97wpCfyGY
QZZJ35uTGwdwkOp8OGgXn9mVu6lQ+s9uUbPU6OPbG92sSZr+zBFRqUSJbnFknwwU
7rxJF/hEdxYtUDVRfFPij/LQ5uUM9kuvZbDvluzyzhJgO6Ufipa4mSZfc5atCGxw
tZReGE96fx+9brGijlwIbA835swY8csGrtNdUoh/8cajk9fRf+7I4TgPmTm/zsoF
2A2sAwgf23V5OEqE54IWSHqyipsZ4S4MZInqxrxKubDUD9WdLfNJAJIAqxx9GAgo
W4454Yu+UfoloqJsD2qpL9Ewsy9HMWUekk0qfoBJ0vjuUCYHOSQ5xDOk0NJHX/wL
GJexIyq43CYvGGfCKbQ7k8Xp8+CoRUiB3vjiAKc2VTi0aImGxYMUkdHTYl0pWcj1
vSbVEG1klzODFXWNV2plNeQI/Hq514QL9JG+9Gw925BJ+qgpsjHKQoNqXReThZRL
eKcd3x7NG6cebi0x7u4tE1QizKEkArzz24ZSYx19LNcPbEr8cP3YQ7oDKGszSG3T
/y2aXc9yl/Jw4yOIREFXdp/0s+2OP03THEWwmJXd1TloRuvGxo2Ugq6dEouT8Ggg
NVD9wT0ZdxCEOyqTsfUba0eVKdr049uJukqTpRyet1tTjEu3gqlAXMUhzvGKNS/7
L/0S01TVwZ0MbEc+6ElL6coCyqLta+Gwx7s46rxIoe16oJS6WxzSnvwv8EMD9981
/rG/PAmllnUZaDbKtmXecuVN3vF0orowiAP+sEI1FyC634pbVx1djy/HYGXfyGqr
uhJHnvGjRXFl+dpN1OvjqZRi3CTqhyvmdkGmbzU5ORDoxxU174Npfc2GmRC/qbH6
U7TVx4qr7QdK7oTVEiiGc9TyM3Q0xsiO/jMTRypA9u/o06V2ePyRAA/Xllq6Uw0M
cJXnEk70QxOMEiQWePaF7eL1ur5ISVYfO1ILDj5lnA4VaQdRBQNzrK4kxYCf4s42
yvexumnKhDRkmNI5miDcUtU5I9HMbNzDovehIJSu0Zfh7qNP0ye0IzyJpBnU9mg/
wAxCGXuUwWu3xVqOWwosIuPLOYnHqoOJhAvyayg/Ht/7fVrjEmHNS60ZvXt9A7vZ
F2xE2zbJsMie++fFFOOsVWXYMW+Hl4fIAmW+FYg0s6vZ6s3sgVDDNQhaUM01xmmn
bEuIsoIIQyXy2QnVPIYDyCHtwOrMhhbIjbNoUeUdVq/O26OGmAccbOdV3fOkWNZo
mnCowv4WBfD0g/GjU8T+XAVVqPM6S/8Ri3uKlkXzeNCTIAhCTAV3nXL8by4liNQG
IybsF10vRf9QS/eRPbruLyqHl55J7+FrDITcKrFZ4x8J8td8gVIewzCuRKKDPrGV
sETC/YoQS3BjFI4q5UMlvAaBDidVjyBfr6WZ6VgflI3Jo1GTMNu0p5quTVqSnMlp
moDb5pz61UjUqidUvan/xhVcI9iYdEFw0oejdxu2a5oTfg0YvO5IikDUtNfgGwIc
zYM9fQdE1RgfKTRa9e/yc3WuUE8Ad7nFC4aRHCNPVE3PRXMNyE2TIm9itOgmXUJ/
TJUt7wBXnTs5Ug7tsbRat8nIJ+SrHbCBMqhQ3bxuh+56ekLbwGHAWQAdCyhZrC0N
17iHJw+og2YT4QkomDGwjBYKjIv2uM67Kr+UzKuKg9BeEhgQFpXNyWgX2m7p6Fef
4TwySAaPn9P5d++qOWqfcRJuL5wAhR5IlXVApN7HQaFTGwddB0HdZC3QWznZw5Z1
bNC7TMuVQsrCpb5Qit4jDZc4S8e+hiN4FJ6l5FhWJWYn0AvcDT2r0F5/pz4P6Utf
ACkT+MUasfZUtLNwF6W2ODCmZ2JFvjr7CPM2s1jIJqF6FpBiexn7UsGGAJYzLrwO
LdcyFliFDXTOk86STE2+JSbhdSjZNkkoqHJT1y2yMKUQ5D9XTpihJjJLcYJ2LFNc
TQFL4Me0Zelngf2m0aM0oN6w+A1cJDYVN8gfo+8c0nRssP7MJL13sjZaxgKfGPf7
aV+VqzDMv7SjkUfIyAahmUY6RXQs2Sb0pYNj+bX1vtZJhimaz6FSpcyjhl7sI7D7
5cqjg0Qy+yJGWBW3v/zRLMvnQS2MzhtJwwFhdRx0Yekim54upNLglpPI86q6J25a
eZwxFKazRJHJl4reNSBVIuaXFqLUoc5ltrCk8QheXrHaZBQ+sXi6i5+3tXZrNWk0
ZOy4atj1gtAuPiaJ8xZ3c/s0tDzScVd6yiAJOrsCTP38gkYEAerlMQMvS1vc47rL
JeVx+SpvbpVjqbgL7C99VcAcr+owMP7D7k+56UnlKNzYIw9gWiQDPlsXWJG9ZB6w
EVilpuzekrIJ3lKHiJbZviYEIZezedZeTaPKlsGl80FcJvWrNyVpvDX83DxWFXbH
BdZtS02JqfMBVEv1ZjaSM7uSdEJOJrlGZjEcif+SRSr/Hm5wNm3a4/fBokT82MSs
tKvkuj4gOwmc7Kb4CjXdZuWeuEVS6Q0rKmudDi4gssxclRX3NrLx6J4sAjr1Upar
ndG/yROasQAgb9I8PGx4DZpA2SQ7XSIAIr5UZ+N4h/vpLhI3dxT9gPMkNisVJEZ6
4gX42+2dRd51G+/GHkCfVQXWhodJ8HV2xi2A5acdNRqipJGMzLdTasRS2f0W1WTL
LeAgkwah7+IE4F1pEvMhhfU1t+o7i5OrxeBFRSdPjprLkwhVh+RoH9wbRW60jyhq
jKo4lhSjr9mfR2p3A5PwBZ4lVNNTrLIUqXc1MybKllMPSHna1qODZnDDjAmxyFRX
IwDsAEU17dyKmy0riTqFG56wPf4sqKsZ7wyM780Wec3DTQDvgHB05Vxbu2CQ1MZ+
mTF3HbrbR27TvIxR9DbSSE6c4zCfnIzMC0gVePMPpi7bULC9wruxgEAZ/SwbiBXW
jsgdZg4K/Ni/7qZHGLqyk9SJYukgjKOmHdffSSEuEc5EWy24le4u00wd+BJm1zbn
5uOX19s6a266HIv39KeuTiOe3R6iZFiHvp+FSyn5XeUz0J3sDsnNwHciJlLEVqsZ
Y3D0HBmdHFDA0Y/Q1tYfVvH6oF63y7s28Kgfv48IWtCSqYsT7oS5pSLMYCSO/FqT
mWimWs8tHkiyCEsLQUFyqE0oi2/gcvQwd4oskfiPa336q/Of1XNgwEleDgYMOjtC
x/zia3GLvVKCEg7PH5loIdTOlbFNF5dOPsZ3JflBjXyS2VEoxbRHtGZjHr6O5+m7
RYPKHu+9D4dlmbktpSmrDyt2b4Nxg9eMI1ERkX72rF+2fDwa/5DFxqUC7s9CBj+K
RYV4uPfTVjvQ1zHiorSJ6CkhowG58kCRaJNw6GsaOVJknwNpG5rHvbw3iGaS2LeL
sDXUuwe5blar1PRR2C4TlBp9J7xi3iZuBD1Kz6aOOI8gkd3Re/4mMNRoLnjkQnxm
qYF/d1x6VGg/JfzKpgVImOkzxEzpUTiQ2naT5OCh/CnLiyvU+wGmOwTzNhzqNTkW
BSugHUF/tLtwXcvb9BQnTAIxl/6HjoCvBtrmTNpICF3q9o6yyK5zOttW4qoVbTKV
zLgG6Xio5R7V/BFnQ8bSVuuG9rAxZX8TvnIO2NEfaS9GeXSUHraPo7vvTU3zgYZQ
RSff2Z6MK1jdJ9lZ57eTEG//q4AtxluLfV4S6V8g4h4kZhKwfI6EA9JA7alDYSBp
GHQi0LlqjFVPWRPeQPg4eMFxT2KRKF7ra1qUpxClVUs7FhHy4jN13Lko0652SPxV
6M1iSVYXFznWj8ta9d4i70SIw2kZ7HfYsL2+zleIvqxA5mn+7wmBpqcZg9bVQyYX
n6ELASCLEGYBxsEeofJbwdzW+BUbn5GbPtuoACGiqaxRVsQSrz8P4SRO0/BHYRyZ
9YNRtidSublMxrfynZ2R80chj3nrQLef0j9NmDxfzAsN2xjuASTxMLD5Hs5N4uR0
HtvOhoCZ5oZtXiATO27BuWJou3RkjLe3p0/qw0uwJ2TqN5NeNdfvbjGjlWNSwfJ3
29psr4dEUBchpy8UomYGzlfkpS7+mqnVFFgQwvlgkSAx8fUrO4I9P7II3+hsuCSB
b+uYFUVYl++CYL3epuuMI1IktMhbF8pvvget3nKGE2O5J4j+4y1DN+IwDq6X0lz0
9dlUqUz9SPoBCdNEVGxfaDCG9Xz0yHPY04tutNWpx1tYPaU2kJ5C3RQlFnqzUej+
fGV1xnN2W5bI/owXe0R0dVaWBe94mrPLWkzEVoBJWE6UCiDlWli19LoVz2hF230C
EdY7U29biWTaGl+uQKrVtkZqBU18ZPQPo0Xhwyn00DpJ15CkD2fqoJIKMWZJ3gfJ
xRqfNbFQHQ8JN8GDKzgJFLkLSvIJihLx5eBlxdeSVcS9Iuy1mlDBGeMd4o8MOXKT
4iOOSWuansdkMyEG7dl5RcuML4TYdpe1o77lbaZifxPxOP8foB2ZyA7SN1iJMwuU
n0c+NgsOnb2ajuMh0FMvtdP5OLsZs6K3kbhmdoK5kt0xT4qvGBk2Ah4iDHXI6Nct
5nMUJOKoEMVLr/lYmCEwVk8wTDeMIxZpjykbfiiZ0fUiavP8DefgQdFIsT9NAoe1
YL8Ole6Q1Iy/4FmoJXhH8Fz54CVEIrbBU4liCqcdcHjgdYAqZI0YRn3zr9k4SJyB
Wm6n9X8IN8OqCXJIbqkGKAJ/mjgReIQz/EXyx7FmtJUvo276euj5XP0GhonBNTQp
b/E1m8Z70kPneunnkunuK3Rq4IEiYO0jj+Ml3lfwu1wbt4pS7dWGF6M7a0sAIIFY
2Hwm2vX/hoMoBFtE5mzedw6VaPI8J+6WVIEAN1zXoRorHHQ4LOAbos8wQeJE8g+W
TUoq9FdfdB3+aWO+UioYxeMlA6q8YNmTGkAmB112UWv6nO2rJW3AB3VCJx9HOemd
3sF15zhwHaI394z0czTIrdt3I2ituGTh9AAN98VpyPuX3rkzSHHvXUyx1+CcR/z/
ixCcYp7y8GCYEkYheYTBrwdjIecQPmM6tXzafdUwSSbDkmJ2n5Aj+/CqHAW0Al9b
sS3ydHQ+SAlDMr9dQJl+8f2sWRKNd/ePvG8bXuGoc4MJkdcj/Bnh6WrEXl14Shga
IlBYuOzst4ppogjOB7isMq1xRQ1ettiHhnLlEGuLA2ECjaTvaMvO71/cn+Dq8Sk3
H3wvo1yniE/nuaCNvqh3kszHU/4xXTF9JRI2sbeWc718kh/ms8bAyG0kp7EkLh3C
WntuGtEQTR0dmakPnPUYQy4CFVqFmxaqIw9073JvUWHdW1P6G8VN1Ozt68zRpCdO
cPXqDaqRqonJNEUxNABNDmJMHUEMP9rwzL952pVHW/J4piYQfRybC9NIZMk3QbDW
/7hcsY9vlKgYMZQmEegeoFreQ2OMHyCh/kg083gWrNsj+LVIQIxENx7neArvQohK
T5y0RpyVnLBDRdB5cy5ak6LZwl2NxOBY0N/BEjgJWpzBJRrZ8y5ovtQp4XGFjIof
dw2csdEK6To1FcqyxUA9cOHmzr3J+DhUfYLAJlV4PHM4dcEezeuQPX2g0qgotS8I
1jwPf7vYbCSxA1ekvo+FmD+Fftzo6jyy2scZdJn3D+2iTF17Z/MRUJIePaJRwKfm
N5FUGCILquepqdj4xuX/FITRnQRqBKEu2auci9PHft3qIcQ+j0mL/Gzn/KiOUnos
MwmqrqiDBkKOvW4Lf/hVNLAnBj3zE1qsyOXDldHUPYZTAxi8M2mGAW8RPN9jFC0l
sMRNpLQsrKsxrrGfWc695OC/+HD5KFUtaaPFKHHZb3oY2jee4h8fO0u5Rm6I4AP9
nGUBBd2Nq93p5jDKkfgNjiF7fMEpkO8vTRDs38XX2/D2n3jjIPrRCcfP5bDe+6kj
CcuK8bIN+8lD+LpyFBAUK2u3BQxCa6GGT7Zb8b+sWY8tRqnNe9i6nTsjS+GcbQF8
I5hkYRd53x9nsMgC+RrfZXk6qUaGxRC1VIe0c0fuaz/+U0JTXjU9OOXmrny6vSLB
6HoLmTo7kw1tBxjyvfH1DtWcgbMIhj1y73KTmINeukCjstuAto3IvX6P89Vfno5E
IOJ3qcdFKkpnQZX3fNQ9PUigYnJt3HJZzp89RP6JHFqaU4YKE8+xEk5ePiaHPjSb
T3xXkuCKLbF0JrLpkESuebVEIrkip9T3CbU9JIpfGlyXFvXUcdvBhF8uF14Yq/Tc
HSEndfjtkKrVLLZi3SNIqnKlJb6jQXhRK7iuoBQFydaaD8vgequbfsV2oh3OtxZL
73QX+POnWFit9gLKjmhnIwR2TNU6TLZPFEXbYbC9VADbMfHNo2h2rq/EMQhJtynZ
5ELrRno/gqMMh7KsAI83syvdM7Xy2NKgPbMRW1zXZ9s69Zg7JivMtt5OnhjRhvLv
iizlyewe+E2u/yE3oWsZZdbN9xpV0cSKoQHi+9bn3yAttBtKr9gmaDxrwd5UdLaT
r9sBRJzOHwavwskS0sTXcNPNkFPfucKu5yBzEspmgJM22DU7AaCulsII5xclP1i0
s6uCMXfaE4+jedQAW1lHQwpVTd4syb89vtCWfKznOXh1P25ioC4gx+QXem+FTS2J
UAEV9OYOX0zTjLUEJO9el+NBpTyDMhL4VyKT3rBQL5rC6Anq8EyRwAOHDY6Bw0PS
HgGUirqleUhpJrx620fAWxUxD9Mv+lbCNIbxU4zkrq+8Ea11Fb14Qecgsi8CPvAn
j/7qPxsraNSDwaHNaMq84kjTQLquXSXa8tYocp2QXApi9/S26cywJtZe1Ke3Buyd
4DevSy3snwFVVCzM9AuYSaQV2nNjFmttfCBw1+IuKT6gK/QRDwcCcxIZHi5ExrSe
yIALDQjbkOLpJ6xsVErgWe1e0bxzIvUOwHSWgkmyq9/VoLWiBq+ikhcE0hecpWmu
0ynXUU7XVwWZVTU7wmTDvExXXsDjw2cKwgwY0Fire6wIO2954e1e0EzdVTWXjL30
0uHbJoVDIzNuz9c2ZltDXmW2ndORbsF/HEDqmDro3m/FWiGUr7CQj3okdrWyYSAQ
kOeU5+mL0g0xIx8vfWdPcIQvFb2kyAbA8yrWbI2j5lwdH17fXclC/I3CCKlHNJAl
7XwQwmD/dWBNHFDm5T6PHVZX/MNWk0GfH0VbR7/6GePSdbnSlX9cGwLJmMrNeUTR
+YBfdkXmgKy0ifo2Es4bKyLirzm4NghU6v1TOIpOhU6dXI4RM/hAnr7VnyNu4mSp
2FNN2sCq7GA9sEQUhf3DVLue0DvT62Nh0s1IryXheeIXs04JASZUTU3IP/sXqCY6
gpsSww9G+BeJ1tSIKS71ZREFYHmjaHAHUdZncG9tcB8x3oRD6+An5ilC6FIRNRAq
Vdj8di4I7S9SrbNIbTt+0JEBQtr0KURUbqXYg32UUKyxv/GEzwewSuCKglzEoGKM
+kar1yk3Ko5T7Besyb4n1Tf+CaA4xSGPgfnV//EDgsIWWvpjEvGmA1MQhxdoWozO
Xpd0dBIGqnM4ZkBH9DDYdxOuil+j9rPTeaZpWSooMUZIbEA0ijn/FHSvluTW3M0l
3BgcytxAaCdBbNDEc3r0xdPkZpmQfRxFTmwNDJLR8K4HBJ7t6D3R6wklcRc9VuF8
agpdc+mYnYhnV2eQyjuvXQApu5hrEcmdXmd4aozFbPjfwCMNDV4BsR5G8aS6Goqj
0ylgm2cNW+1AyhlJTybPcW/WuyjxdxDCfj4UMWo9rnTflt+2DadbtK7Xu0AG59A4
WWvf7caqGfcCehMqpGiE5tD/75+pakXM34ux87xRyrZafjOo1K3qkdU/1zFxU7h8
cNGjVatemRvp3j39hzTEpQAvTkv4Mte2IXgr1o2SyFO4uR+0BocCcIdta/OEi0iK
UBDCH5xckgiUDjyHpFMLrvdJ4wI+894vFu0lYNpdJh6Ed5yqHr04tm0RqHL9D3Sf
6lUhKjP2Dmgr472WfBcvZu9w9vGPdTBeZA1qFRVHXUA3cEQ9PIj8bdMO+O+1U1l7
u5zQx1iyu7Ky3JYlRbUBbHUQb+KJJDLSTdT+sWAKEFqNJiEM73xANJzRj7iDIKN0
rpyhjqk5X9Y3fx6TBWYq/ynNpJvDmQFK6f+/VHyONC7pJpS1VLMO/OTJ1/wo71Pm
zonPMGJZyQ84ukN0GT1LMThQUi4Z+5MoJumOEXJoee+6eu6a7FR+Zgbtd/Tuo+ei
f+Oeb4QHRzyjRlM9ReCp/Xls0QOIrqPcC7bhKfA7Y4XbxeHpH5NvXjblew0+TdHD
8xYZSsYQkDXel1b32e0hOP6c2EegD4L+pkCN7eBnUBWIjM6slueh27CPYcW0cdjQ
Bl1s5YA+qB5UgvcF7yjGw6L2v3PrqrXqTPqEdN114wG3jHE+7OL01mPKxysnhTpP
FdtNHl+AItP5OOJGsOKyqR4eNS2AGRA6nOoHy1nxTO4stkg+cl27eFq/rkRBXRj9
Hrkq7JuzWLk6KlkIKmR+FSr5LwPdooiZVhyu6ycHiihwYUspfwzh1XacqoeLZkTp
9EzUV9YwT1Zanhz/0E32J9o4ApWE+xm4vDQSfrdhS5rJ5wYXLFeAFzW69nr1U8zU
1rIle0dum6tY1NYiZCl1SdvZ0dK4G/NaDnZmg0Asa4rprXF3n319eg2JjH59qdYG
pTb2GgsnxgjmbKX7cX+5EfMGhav3dkRJ/WgK3V/+Kwx3/AuEQoeO1DsHg/7VV8Aj
YsItrcxGfzJ5nXc+Vyz5InDbGrf7naX8qQ9Ce+rZSBlZ3sGyruz83fq5/hMpEp8b
UhBpbmEgwoZ8zttzFamG6bjpaOJk6s6w0zidlY/MP3G23SWqk+QcBR2K1WytmujY
R37CJs5YRN1RmJkvSJ/oadkhsm6JN5BWTBd89NDi8phH3J04yj8dD8ImAme1JA7x
SBo4+EaRc5ki3E1Ar/vqmI4ZepGREeSVZyVRWzStB+KRkPRHQlegjmRfy9bgZZyM
0umHfDVshxrJwtzvQsSP5vYS51gNXyQob70MAajWnzFuyTBSWKt1R0b7Fng2Yvlf
upq5GKoAjrrP5Tb1g04kKaAXP7NzWZ4gUGqu/F2x0YA=
`pragma protect end_protected
