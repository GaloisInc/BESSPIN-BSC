// Copyright 2009-2010 Bluespec, Inc.  All rights reserved.
// $Revision$
// $Date$

////////////////////////////////////////////////////////////////////////////////
//  Filename      : XilinxDDR2.bsv
//  Description   :
////////////////////////////////////////////////////////////////////////////////
package XilinxDDR2;

// Notes :

////////////////////////////////////////////////////////////////////////////////
/// Imports
////////////////////////////////////////////////////////////////////////////////
import XilinxVirtex5DDR2 ::*;
import XilinxVirtex7DDR2 ::*;

////////////////////////////////////////////////////////////////////////////////
/// Exports
////////////////////////////////////////////////////////////////////////////////
export XilinxVirtex5DDR2 ::*;
export XilinxVirtex7DDR2 ::*;

endpackage: XilinxDDR2
