// Copyright 2011 Bluespec, Inc.  All rights reserved.
// $Revision$
// $Date$
package AhbArbiter;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

import AhbArbiterSupport::*;
import Arbiter::*;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

export AhbArbiterSupport::*;
export Arbiter::*;
endpackage
