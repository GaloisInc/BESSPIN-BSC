// Copyright 2011 Bluespec, Inc.  All rights reserved.
// $Revision$
// $Date$
package AhbSource;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

import AhbDefines::*;
import FIFO::*;
import FShow::*;
import GetPut::*;
import Randomizable::*;
import TLM3::*;

////////////////////////////////////////////////////////////////////////////////
/// mkAHBSource provides a TLMSend interface. It provides a random stream
/// of AHBAXtorRequest objects and consumes the associated AHBXtorResponse
/// objects.
///
/// If the "m_command" argument is Invalid, it randomly selects READ and WRITE
/// transfers. If" m_command" is either tagged Valid READ or tagged Valid WRITE,
/// the stream includes only READ or WRITE commands.
///
/// The "verbose" argument specifies whether or not $display output is provided
/// for each request and response.
///
/// The "num" argument provides an identifier to the module that is used in
//  the $display output.
////////////////////////////////////////////////////////////////////////////////

module mkAhbSource#(Maybe#(AhbWrite) m_command, Bit#(8) num, Bool verbose) (TLMSendAHB);

   Reg#(Bool)                 initialized   <- mkReg(False);
   FIFO#(AHBXtorResponse)     response_fifo <- mkFIFO;
   Randomize#(AHBXtorRequest) gen           <- mkAHBRandomizer(m_command);
   Reg#(Bit#(2))              count         <- mkReg(0);

   // Limiting when responses can be consumed (using the count == 0
   // constraint) creates back pressure. For instance, if you uncomment the
   // count update rule below, the grab_responses rule will only be able to
   // fire every 4th cycle (since count is 2 bits). By changing the size of
   // count you can change the back pressure. With the update commented out,
   // count always == 0 and grab_responses can fire whenever a response is
   // available.
//   rule every;
//      count <= count + 1;
//   endrule

   rule start (!initialized);
      gen.cntrl.init;
      initialized <= True;
   endrule

   rule grab_responses (count == 0);
      let value = toTLMResponse(response_fifo.first);
      response_fifo.deq;
      if (verbose) $display("(%0d) Response (%0d) is: ", $time, num, fshow(value));
   endrule

   interface Get tx;
      method ActionValue#(AHBXtorRequest) get;
	 let value <- gen.next;
	 let tlm = toTLMRequest(value);
	 if (tlm matches tagged Descriptor .d)
	    if (verbose) $display("(%0d) Request (%0d) is: ", $time, num, fshow(d));
	 return value;
      endmethod
   endinterface

   interface Put rx = toPut(response_fifo);

endmodule

////////////////////////////////////////////////////////////////////////////////
/// mkAHBRandomizer provides a random stream of AHBAXtorRequest objects.
///
/// If the "m_command" argument is Invalid, it randomly selects READ and WRITE
/// transfers. If" m_command" is either tagged Valid READ or tagged Valid WRITE,
/// the stream includes only READ or WRITE commands.
////////////////////////////////////////////////////////////////////////////////

module mkAHBRandomizer#(Maybe#(AhbWrite) m_command) (Randomize#(AHBXtorRequest));

   Reg#(AHBUInt)         count       <- mkReg(0);

   Randomize#(AhbWrite)  command_gen <- mkGenericRandomizer;
   Randomize#(AhbBurst)  burst_gen   <- mkGenericRandomizer;
   // pick INCR burst lengths between 1 and 16.
   Randomize#(AHBUInt)   length_gen  <- mkConstrainedRandomizer(1,16);
   Randomize#(AHBAddr)   addr_gen    <- mkGenericRandomizer;
   Randomize#(AHBData)   data_gen    <- mkGenericRandomizer;

   interface Control cntrl;
      method Action init;
	 command_gen.cntrl.init;
	 burst_gen.cntrl.init;
	 length_gen.cntrl.init;
	 addr_gen.cntrl.init;
	 data_gen.cntrl.init;
      endmethod
   endinterface

   method ActionValue#(AHBXtorRequest) next ();

      if (count == 0) // needs to be a "Descriptor"
	 begin
	    AHBTbCtrl ctrl = ?;

	    ctrl.command <- command_gen.next;
	    ctrl.command =  case (m_command) matches
			       tagged Just .x: x;
			       default       : ctrl.command;
			    endcase;

	    ctrl.size     =  BITS32;
	    ctrl.burst    <- burst_gen.next;
	    ctrl.transfer = IDLE; // generated by XActor.
	    ctrl.length   = 0;

	    if (ctrl.burst == INCR) ctrl.length <- length_gen.next;

	    ctrl.prot     = 0;

	    ctrl.addr     <- addr_gen.next;

	    // align address to burst_size
	    let log_size = pack(ctrl.size); // BITS8 => 0, BITS16 => 1 etc.
	    let addr = ctrl.addr;
	    addr = addr >> log_size;
	    addr = addr << log_size;
	    ctrl.addr = addr;

	    let data <- data_gen.next;
	    if (ctrl.command == READ) data = 0;

	    let tb_request = AhbTbRequest { ctrl: ctrl, data: data};

	    AHBXtorRequest request = tagged Descriptor tb_request;
	    let remaining = fromInteger(getAhbCycleCount(ctrl.burst) - 1);
	    if (ctrl.burst == INCR) remaining = ctrl.length - 1;
	    if (ctrl.command == READ) remaining = 0;
	    count <= remaining;
	    return request;
	 end
      else
	 begin
	    let data <- data_gen.next();
	    AHBXtorRequest request = tagged Data data;
	    count <= count - 1;
	    return request;
	 end

      endmethod

endmodule

endpackage

