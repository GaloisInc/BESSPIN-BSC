// Copyright (c) 2007--2009 Bluespec, Inc.  All rights reserved.
// $Revision$
// $Date$

package Axi;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

import AxiDefines::*;
import AxiMaster::*;
import AxiSlave::*;
import AxiRdBus::*;
import AxiWrBus::*;
import AxiPC::*;
import AxiMonitor::*;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

export AxiDefines::*;
export AxiMaster::*;
export AxiSlave::*;
export AxiRdBus::*;
export AxiWrBus::*;
export AxiPC::*;
export AxiMonitor::*;

endpackage
