// Copyright (c) 2007 - 2015 Bluespec, Inc.  All rights reserved.
// $Revision$
// $Date$

package XilinxVC709;

import XilinxPCIE::*;
import XilinxDDR3::*;

export VC709_FPGA(..);
export VC709_FPGA_DDR3(..);

interface VC709_FPGA;
   (* prefix="PCIE" *)
   interface PCIE_EXP#(8) pcie;
   (* always_ready *)
   method Bit#(8) leds();
endinterface

interface VC709_FPGA_DDR3;
   (* prefix="PCIE" *)
   interface PCIE_EXP#(8) pcie;
   (* prefix="DDR3" *)
   interface DDR3_Pins_VC709 ddr3;
   (* always_ready *)
   method Bit#(8) leds();
endinterface

endpackage: XilinxVC709
