`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Jgsw7YULCtwwga3T2U6c82c/CcpDUvecYqw79Nc0liGIczx3DhaK2lWS/SgDtt2g
YujDp+/Me+RMXfquCQ1PQWDG9t0mZXFL8IfABYeQomjZWSwLxnGnKbH+KdkrZpGf
63CW9CN50udPkkYwqrxFUT+pIx7drr5xFnpNXf1GV/U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2809888)
A1J1GaX80zaqnOhjQBnePSGsprybGrr6Tv+CbIPAEMyVL7MI3BzHnugqXjo4ctAy
DIoTOpJbkUUtQGuZyAV4sOVCQPWV3IY5GfsmCCo8L8g94cgDqXLwJz0ln2D3wbY8
NM5DSmYtylp6j+qiucYWFIlrXgw7b8IlJv6D1UjVIvwTxaT4+fde+Z/pnTBNu5Sj
jNPaLTOZBXK5ddeXlzSJ0oops1JLwx5/fA4CP2mXN+tgS+ZNvpi5PCgdSThMfFCd
dRTt4BsCAvs+MWJqOxDbV6L8ZE9gXfwz+al1hi1ZvfzCkspcwo0KsBVRlokM/uWY
E/7aGt79n8P1ooO4KGHU+VTlzQ+UZveB7CUkXZghBvUyyosAluC9FcpTLKLC56X+
nsqaZiIoV0k8Z8VX1hS7CvdtiNvhDKjjRzR/t9WXKOI5Ccqz/iHti8SPc9naR0ig
n/vJL1YL049EBEPH8GYQY/jTFNBBLrIyDqpvMPwJhCP6iB6gMf4qeoKR1YhYWZn1
PWPnmz9VFRUkTrBxyeiPFdnOMapnZLTP+/H/6qoMu32f7uy0DieSFRJbXtMcQE0/
rMqMvUQZaxVI85jXO2ltSmt6gNQBq1sMMde3ZhgtB8ct11rvUCxa7I5r/O+IqEl5
qagoXJbWxbeA5uTXSCloIWbVwrV4vbnyR3ijsQECKy6layZLZ4RnZd9OqJszGaE2
7YV/YIY4RTTSAP1vRSWP2QAl5SbJMduuiELGuy5xoqGabCWfVDVDinmqPhB4I5S7
paVl2ocK78HU6x1DQ2zzDEvkQ5fsGzPpmwvVVVOIRIseBPGQAdOWP5o6rJuhGY2Q
YEiffrFySaLHJr19eb0X9VMzbXAV4GleeFsoPIDlIGlZBZpEQt4nwL/MZRELdqV8
PlEAqSVMz+NZ09ARcg2tWjojRQVXQwpGqIj+fJqRhAgtCR0XWdUvTFtZ5Qj1BK4S
ThkkY/uvkIffVl0IH5N84ne7TdCMQzghHaZrvIjopjFqEg/i4P9bdeH0MBbD2vlk
ilICyDKAMm4cHXcWWGgHutVCZ0K7W8RAM/+cDEXKF+OtwXSAuIJMpzfhS7vnNhxo
OBcE2TCB4EEBHJcLSGYRMMhxnPF0EhC+LtKYkpuDlOW6YNayYfbGeKbvE80N4i/J
kByOVWxeY4eXMzcRTXyHbrpBSbQdxOlalrKRlI7niCP7HS3zO5OBPi1AtHsawcYJ
9sr+rlb6OcJPzkLvTFHDJeFmEywV1js9PjksNm1fHnJJhs37OHG5w9f9WGB/1W2N
fFQmm526A8/GdbL/ObqJCT2EUmXe7dL/bh2o3aRf8aSRv0NBWcQZT2p+pvD4Rbmr
DPpqZWaNaWKL75a7a87z1CFZzMG+fU/2lVEoJb3mbdTylhvadIsyxEYJxmirxvhD
JOWQqv+iHehORTJMNp9Tzp/gmrzG0kjX3Xlf70f0dgeb+Nhml4HRbZbkEzgy2nrL
ENS1Yzl+KU61UYdF6E5IN+JmxVuybhCUCKMi9CsHvILTQsd5Ql3BUxaxXwqZCixB
sf0Xb8/1bod7h4HTAxU7eBuMdWqXW8aiFORqvuZA2Glq5hSb4ynpI8jhnMykP/TH
m28aQgv68leA9ZVzxakwQrrkGRpAO9CbPlr6TNdDyjTBq1957ClVMpGi5lkEkqIE
ZuBFYUqg8JmSu1u0QjIO0garqvqKDaecnly3n9UOxCUP1iGCtAV1IzUaZ/EzM8H/
Y4MB4UHaRtR+0ueolb1wM0etyFSC6+T1fy6BaardMjqhPMQtMEbVpNh56N5g4Bqh
nM2BA8MU41flVPrn35iDFbLZnifrngmUt3bZygddEy/ay2ISoMpD6lZepB9aikrf
qEo+gssoWU/WzcY+sl0Jxiw6l4HVxtqBGPcUqOknkXBGF+G8xIAObtOd4phxHzDy
ZkH1XePwEEQ5Rlj4leO7xkXJPxZQAH+YdZEfz4Ffqhuba7KvWFFRNwZyWj3Q5hQN
wInU1CPT446bkJAFZz9YHAVVwk/LAPA0XjxMuyarQgiaIfoX6zc4BOvAEnF0Nj1k
MmbQdSNFZU6lGG+bsepeEUk2piqciZcpKHXbAy7F5tMTabUhX36atl1q0wQHQjAs
SvLxpnGbEIbm0gkv+PYTQkL2A/CXbQPWF0mOBXzmmhFqCYazM3hsF/em1YTsLRqy
0W6RUcgZxPpBBloOOkPgupMBxJfZFsZfs+E6y6spb/UcK/RdTmfc0O+6U8lRKJ7G
5oOwtrFB+ZB3KTe+P+tPlmTiNoCjc0JEO+T98TVTt8KexLmseWLEv/cbIJYtOFHx
yJ9XWWYIUI3MGJdyZxVBPdv/CkasMGB/wckRgdBrD0PNHwT7WS8zyTR2HFs7r5rM
Q9G0YaLEcLTZxWQGFwyBVRCtjk/WcXRGK3N1wWqnvdGp9ZqJQNyH6st78M2kxk64
oPHL/Rh7mekK/jiNBJUjWmtQmfwxjbDL1e5MGDbyrwR4YZYccuZDs7M46AAYXoXn
QYGxXnfD2nBW7DeS76cWUfbYHqexC7InXgeIlksBoKn/Pv0rhkxWUT7hKqArCv+e
ZIh1J+reICYGHa2sOwothvcjD0RuIoKaR10LQGZ6k5S21fARLLM7soUME3TPahRL
cpVswepGF76TCc6YuMYQvWx2l15UHyisxArBe/+ITDEuN9jp2em095N+wxb+I0gB
BcC2USPgrO30lrLZ2rN5a1TWYn3SxA60JXHSbXG9EHjqE7ndXQGu5eIZapNW5CCr
gkR3YKnsKYyPmvspKbMumbqoCEvupGEWCycl4KcsF4qUis0hWyt5l4LBHC/KO8Qv
Mfd6vlshGHRzYvS8YdI6uzZ31WFzXSOPkdyznXVviLp6Fsu7+Z5X9URiGNYk0k30
X7tR8cqeODDSiYNmuxEWZa2IPwaYHi7caEQGDINU5BnzKSoMoXGf/2IKqMdtkefG
q4Qp7UH7f8ToDzkGDFR0xpzQZTynlNT+upBN2D5hPA6ElxelPOgac6aOlih7xhB2
pmBayJndYQG6/ir0yuu4sKLT3sgBnxyvmuho7R1EjYtmM9iisVvMQYb2Z+iCdzd1
KZFB9anHuoTihsSJ5QvLLLv67H0iHZ1G2zOPYhlsxhUpWLPapm7xA/hSz0rwkrFq
IoRY5gi4JCGmXirsQvPpIQO+GectUFA31i3uRrukh3Qxt5MNf+RtZ77N9dRmW+SU
NJB/9UdHBZKV/R7CWs3ku+NBQxx58Y5LWoX8uhK062D6d1wC4dPH9GW2CJv/JtBo
YYZZxtnVF2EQrFimh7ATig6c9W6rTj4sCvMUUn21z0gYw8GpaxE7KX0HYJ5fHH1+
BDDWDTc+v/snVGNQVRYZoI6LtYXaKvJ3bv2O48UO0dUaXb9xm4gmvgyWaIOso4/s
+0wYcGMJeHz1k+8kjApvvGilvZSYIIjg1vdzM0JXkqmBiOiJU3S8nFh/ndjczf8O
8TCH1NO00KJpUzh4oIRS/coFObHgL8WPLgjtFk9r9OsByDt2RoAnsAcedhYhd/12
NhhoVBqb0sS06IpMIBeL5OJak2WAff+rWrnkLMIKDLk3eTDB3XLlyHng1WG6zn6g
NvpqLZlevpSsB3fZ8Cf1YZOs8Ixs/kE/VY/aZwDKlmdRgZ5upLJTpiTEhjt4dJNr
BWzLe4M7T2P8WmhvFaDgz8/CUjDzyfBM/Qz01qp/TkNIclmFe0gxdBQuta1vlLxx
RQ39nIYsGRZL+onMy5fwzeEf7X4RAD9CROu1Ht4bKc/lRF1d/VGetAF2ThPHWRI4
I7O7aIv0hM+0LMOtAScE8B87PeRSgUCsCR/I7IRgEt/a0FciY/5E03XzUfk+d27p
RzBPYfhhjUVvcP+8hq+/44w9PvqIhjci5apAGT8apSddZZ05NXMSs+ExCUSIoX6T
LPfem1dqQr8eeOIi4t+dZ+pY8tVASZWAVav37N+g1c0mDlUn2rQ9CCtNCRS5PEt/
uWQkN1FRbYUEoyObHgy6DS1zRtBMWDtq6gFzh364FhPgmpK4uI4yHVRF3Sz1u1Qr
wNnj2VPvFLNC+/4F4XFXgpkMSJrzUVaWygdrTLFfd50kiA+SoGwbwypdGNQT4gnI
13SGsylDV5NXc81Dcdce6gLmEyv56DQ2EBwYYnKy+CmWar/PY+M5/poNVcx1jmPI
3JWL2ZtmtgLKOYdDttLF4Q7CREj+EPqyJX/ObBC1L/c5PdQrih+Ou0k6/Rvewu6g
RZSpxphI2+l9QPlNzI6JhYUJ82pBo+coH/+XmDc6e9KlUMCnlciS16QPRt8H0P3x
MSrBBiIyk3HpJ6my7ULm1jdcFy0r80DfA8mPc7skmZbXm/E1Ou1TIxMGE/I0O7T7
MKHI3H/DzmNcOSwa611xIuXYFSCgybdEng0XqARMrsv5vSlfJv9FgEX0J4+hfdlL
0I92SBZJ1xvGbdd093UU7o9kCXHBb72Ah85mQmlHKy4+fbQYBsfVIuTX7NBKZX13
uLVlAEia57K557R1piGI1uz6b19ZUGbAH76peu0bIQmS5RPSCy2Kv/y3UWGV0BXM
L9x/WC3RRGQlejGpLZq+ZQ9vS1g67kep7Kpo/Dljrp3SMvdCe4lMs1qJrogvtF6F
H0dHa6DYW1hX/bTDTpMLW8YrrNTVb01h1F6vJ6Me7Rn7sqbraiB3pGJCKdMwQ7OZ
uS6EAth1N2LXVkPfPBMNPS6lrW5cC+BNnWOVS6nTjB/bfJuEi+txjwFfZHtg2Gvo
PNdUO5CGRbYSBQ37UVNMaD9vOqZkizlUGuA3J1hxlbVA9S7pGMTOtzol8GXeHsHQ
ZAe+L7fESoAdS/1Lgb10iHE8BVGgDKwGQDnkuhMx6NdmRywam9OjCqL7dI2dcCbF
gx/5eN0UZkLyRbv4Y28YmtX8zjLXnp35V8STnxAu/XBEOQyzXoe9TEmsnh2JrKsR
ppjfPWdMVkNtIP7GohkoJe1Vi6TIFWzKcVzqRR+ORcHEPM5BSdFHZQ+/VKS248Ov
Lwpqa8TUC3uXIHYmUPtvsPQmJ9E15CfYxGnhgbEW1AdpmYt5z63eUdzo62EQfs5r
tPMxqf6v79dZBa6EJluxGtUiZI7tXA4vN11PNemaksjg1rEN8mut/hkiu3aap7Jm
pMBJdmPe9Y+sqk5cv3o0A2eXjxIajvrx06IwgUbnQDsWf22tZx5RIeLrTCgRAEur
dI676FGQqh+xSk5HsbJj41HnWt8hdT4VVJaUqIvDZMwHaV6by78aU9jqSxIW4SMQ
QtMRqKzsVxnlnq9JJsOen6sw2JYb67iAuBGBVW9QFCnKOSIGcnN2TJ9PYxb+euOx
xUdxU300+fyo2uhFj2Nu1K+S+oRGEngz9mrORzeQ7dHovYyH2sm/idWD7YvfPT7z
F5L896nX6mvP4vbvb1JnHtWnp0AbtOC+Jo6e6TZj4vzVzDbFsYycJXPVYX3it9ws
1YqIh/Pg6I5XiUEEr2a3KFY13iEm6WdoRJqctTVtJjHqDF/5bAnwWiOJFNYk25sb
pWP93wGdL4o8JeK3PKT+rXq9P8ha1uc8MZHMDV/ehPzEWUKdZTHdW2OReTO3l15r
X1tb1ZdwjSR49kYuHh1bUQ41ZtwbB2AFOJ3lC4G3mpDGppYr9Y5h2R6RuRbSXXTu
qID6vrEKuCn5Rhnf93V+0dGZK0Txagr2JAgUDNQl8hxMFDklf9pvb+TLlUxwD02Y
m/mQzrZlvqrfUBySmcfj3XdNWqbvFinYEKCIDDGicJheM+ICuxstwjQiVf0X7feE
pPfTYeSrw0DManKU85xAVx7pR46QPMmtS7q0uvJnu8FPWeh5zjr82kVHuZ3/9ie9
KR3CTwkdtt8euAL0DrEQa+4m/Ye0sBBS0jaNqo3Ph5hut2ozrQWBVSKSdbTpwbtQ
QRJkFuB5ZUWqG5mKkfpHv+2kl0zfzaLlWOMtFfcLN2i5fiIKINLSHDb6X4mcEB9w
ac01jw5vo4TxWBQVJSi7iYMXb66sjF+3N+2oHctcdHiGSJJUJtYtad7ejk7bpAra
RQEVJ1O19bT9CcBBF0HEgERZ9notWIwFTFMhQfbiRabaLye9hoWeo66XhVsk1kmJ
pmdbsWHHS2VXERU6+kklkby1Gw2lakwGujYvDChrQ/2Od+PvlrDGeAt5Bw4jWHhO
ijmLQ3LyFBYQyUogBhT2Ce1HUzEcCadEegmXC4bgsxvO7OWZbe65GMPoaOR4rM+f
DepVuqcZz8qDRJlYF2to7tMWewDj67kSA2f1jNRC52zrWxThheWoYyrnKFlIcB0p
AciGewF+dRGjQmj+Nz4rzz4NsP4/RL8kbKDtD15xBQGl/MgpYP0oMIbCx10jiPJb
5Avr95ANmcALGXNF6zfKa8g9X90WZmdE6AVekdEncPyZoe07U321wlSEcYFCzOhz
LFJzAg5Tvk1IHRViVoZbx+j5912XyD+RR0vK7MR51NYzKyxuMkb0ZdfY6Rukyqls
8c/1m1enKhuwYz7CVBdx5OEE8ad4PoIBHwKsafmmh5QWrSULSk+CPhdb0YhGg3pI
aIXF7j1y4xUVjjdkad5vpB4jC3tgPp5tQiau505zeXuENHZ8hhxDw8eDS/Ao8e8R
EYu1IZhzdUx/677ktrcUlilPzSjcNDJgQdlZXzrNZZR5gZ4eILJdU8T3+qlzJUrD
9keYTSCNtCuED+TaiM9owC5Gs0fZDDA89D0wa5G+0cIvTsNwHtGy3mTxOMstN2Yx
jOKMPt9f8NMj7vsPx0y7hjdojGKwyImdkJvIapsnh1kUI+YGdpqkcqeDK1M2jISJ
q+gT1rSKEowCXXnzt64K1LUECXc4RPxO5Q4s0YhDzejkI2IdoyqDhj2IE0B8EOOr
OkVr+fqQ6ZRgYymKDW0et3Sf9q9HkXl5rIXxGWM+BGf12+4xhkIaMApVi/C40qfi
GQl2OeW88ffBdaIVUV8W5B7TSYdn6AFoL0JVYW6yCrdhjY1O6i2BuBq3ig6hL9vR
B8DPdjBg0THEY9+TMovD/IW+yBTBfoj1AvfN+1q8iMATatgXRaay//z7yN9oUL05
mguEM0eKbyrs+g9ueoVIwIWJaiU4JwjlOL3Mh8eYd8igpU9iiZsagpe6Vv+e1LJn
QvXmhICO0zEmV1UULkYntP0FTsDu6nbp2RPEJOY6vQLWTMJiBjBF3OH9Xhkz2LQw
EdjtZE3S4+nzE7fvqqtWccW8oQdwI+i3t08kJub+u+rWSXflTpTKlDxhs1pxQ5Er
uB35keu8oynTBj0ZI9E+x/yJ5jNbQqrDFWHG1ChmLhIIojXM7pOm+r3IK0RkUw4M
ORCEkRctbg0S7Bz4TRd6cDw+LhcSN6XLi7ifmK8m2FwQxDwuQk+/KLnQ1YZA9U03
u9xJzOqv+TfRrLaa/fZMfS0k0bY3daR4KvAxoUbNBdYZ3Sd4eOOBLEZXf3StqSV5
wCf9m6e/h3JGJqGJF0uFDfANyjLLO6mhch8RkbeJuJDn3Jgw3/aPbgBXJR6A5GnV
gpNtAkDBBSD90154RK0K1guD95uyC2zh5bWZxOGBgw/yfzeIknOaYxKh6EAuD0E/
J605bdfYEm/TwoXCJh+VZS0ioKD1ZELVdccA17bpn18sZOKJytt0+NP6+tlAB5HJ
hY7R/RRDGM77Fgg7S2X7I8iDLqpsyzsT9Ouy8CpT+WVjsmFjopJr38wcIptp9N6V
DVNf+vJrN1mHnPDCFhVfCCMnQ/TttMebR6rHGNXku+Tl8G+ksakIMVhw5AAyIuyZ
6wxZqufgyfpT1FNa/ThWGvHElFWAWTkmkCUvbWKndEeix4K8Fmzhw0Ii8ydmKTZb
E96ghflp9SjbgpYOZA3eN/JsVVAZxkuKxk3vpiYf0A7VkOxQ4zx6qBSu8UkXoO04
oEU8TPkMwzaOLeEe5njPZ+/TiFPR1Kg3JOKrktGkrb2CiWS3cCVyXio7rzdsgHqz
B+DJERlMsdgCF1huZARNktPZi9vH+SWaUikgoadyL5o+lUoRhm/SygKr/pIDGyMr
mU3/GJ6pr/lPB2nV9Bilxv/5HOd5fZeitWyZd07OvlyAvULrFColVahpj6RVWzKK
gazMewOYM/WPfyjCUX0QqZLtq07TyWrgwcZnYYRVuXuyaV9DYO2mGrYSz3au3e/n
6G7/O3Z3Ypsa9N+EjeYp4KLDeRQnc5ZiGyT8aHDoVhG/UKc0DF7uA/r6hCNXHAGc
/rXzYymuXmMfMO04RR82XYjjxmgJDdjv32nw+bQ63rTPQ2P6RqxKBsBb56MeEgKj
Y99spr4xvitk2Yl7g3OzWt272FXq1XmV5NfwOPUzg8etkcAsuoXZSRR0DdIhouLE
NRfX8msFU9XX0gIwPA6FEFXvufrD+ORqXJef7Wa9NaeMSgQYzka2vtN6LH+AnZ+v
vdHmkVgS7d/Lrw1LH9l+l+CCyvTE8Piqwbj66L1lcyFsRH/AcY4vkiYsC2bjSeyo
mWJD9yFVkod/oKVqpUe0KrdeZfIy1AyOkYEUywP/bZYukedCe/rF0hS+iGpNuAr6
/vpilG4XZq7LBwAGLgaDpWwVs9XPJsPQzEvvvCKldd/tilclGafJGAMfC5Ext8Zj
Cjln1VTCpwvCkflzhLlbKHvu+Dm3Gawq3uISUI0Ld//VkDjrII2j2FTUmBQf23Nw
ceRVmSof0f14pOLZ/OsjtNIRbw6cCdjb6W3slHtIip7LcDNDT7ZkvRPmE5bj3fKU
CJzINq8qJQWiNuLlva+ZM1DGfVM1pcbq3y6FcxELG0lykbYN8LDuJBHsALrA6hQf
/euacL1uXusEyoqNvoni8ocixFE+9kaIbk37KmT08JQJnArI7gu2moWKz/8rsm7L
TLRilrG2gF4EGnFfWsKKRNNxvEZTiV8HMpgyeuF1b3Z2G3EvrsHHFUGA74o7hpv+
axK1ttKVcLcvG96R5+v0NCdHnuP3DVw5KhBnSPSu1OsJPZZcl2gWPnqGpvCrmXJ/
sS8P8AY/FoNPUWBLdzB+ubhY6zx7WqXkkoAD2SeWLzNQKa03ofZPTwYGwXas2jfw
y2B4yRp72zOv798Z8CKo0uY8vMf69yD4VBhjMZxh/eUAD3zobSVJ5vEW3IxITcS1
3JvMi5fP1yIoIDiqaTqmUu8yc6uGWDgDJHYhSUG0jc+c8d1lkUPh97K9lmkDQ6XO
OGOMeSDerQ4l86y1MSSqzP++4NF8sXsZGarfAtJJz2VknyoV1pcjK0jYM71DTvom
IzOFkg0H+EMzvX5Esl2OiWP4uGCIDNxnYHbBuFs2DgyNSZjg9br2asKqizC6tC+d
v5CUbeC7cZeJzwnQ32GSm4/17yZ0hJhGf/JS0ClBnsrJ7t9k2F4PaIKN9IynShOA
UT0hCLXcOFc+AuZ+cg8nndohSYLhM7iSTig3XHL5twQI+uojUxNr4G3PiJ28JNV6
9tlduwDn8cLKPJHn0M7LCwejMrpUnmLVLhpgz0GyO3zr4IHoW2ikH80zxhVhSrE6
vsv7csqs6kSzbC4kl7ugO0CEL1m9EEK06+vKAu2N7RJlGlj8lr33PNB9fiF37P2f
N79dfUmddcrHLPE/I99lEuSMVs8nB9Jqmh26wq6mAr8u73QrNStie4smmSnrqKnY
uP+IB2+LAz5bBS3bMD/Jejaft0gs/UJ8GgQFcJVaYOxcbRX8xHgmg9OvFwxlid/a
JCNAs6aNre8AOrfr7yIm09BX7kXK6SUF1UJpVmInqudVlnjKcAs7akbEXPF4Gfhl
Bp9ptYxHeQ6Fj4UswCyQxJKKmxjpb+k6sxBT5Q2dSzEaghJs8aI9UHbqHrqb4prn
MHcuGU2eOh2gED9kx8ACT0++ighd4CkpSgIZPuL1HN/KILiODI23t+BKLPvP6rXe
jR77dSX+axfvczP6PLKbr3c+eCippu6QEj9ODmjWO7HHBqThPfjk4fyQ8UYB9B8u
vdlheOiXw4dGKVOEVh91MAtdjJ1xWSaXjoqX77mi0I80DBUG1P2eIQJYYwWgTuHr
wBpCWl5SdEzMeyjOiBRCS6V5BbmvjwVhoVP0cwjvPxvgCTM2FyZNAqZtwVHjaqw+
otcIxSjx4fs+/JOZpasJrqDsEZeT5roTf+6IY2giOdATRg6bmK/de/iYGCTzZoJS
5RzNlusod9ODXU2/tRB1H6Leh2RKntpoQ/kKDw2FCxX1t1X9XGLjz1rwA28J6xx3
MY2SP0qXMNL+WMi8IzzxxoTSeo6ZfiSZgTWuqYNoElh7fmhNW6hiu37prp0rw/Xy
cZcjPEb+/UnJj85hos+s6yrqsXu3D6y0ws9f0Ng5KwIlsKBncrhogoxAIzZEqvGk
+J0wwMbdFgbFDfTbKP9E2D0SPbHPLyKUqTO3GR0YwYv3RPfTO8jr18BvtIWrYDoI
eiRFN03fRR0eh1Yb29KmJGShvOCCRSgSBIadRSDO8h7bwwUA9HnF+90SoucGfH00
jL/bqJNQepKGSH3I5sG5Qoifn3P0u5eKNYKQIUbezjORKrh8mqNqBC9Oolkir9xS
COXFKeHYHiDakn21dPh/+S6b6MTlZ0UcvI829yZx7wrmvkVJNK3QutGUKycpWSWR
M6U3BJdXMGC3RPnzl80PgoBisnAr/qK2ji1XwueZvY3uNTfyUBLgzlXMumj0ETXC
w2F1YxA3UPgHh+oyM1qKiVMFOAAbofJ/YORlpiXbvjC2NCvfUuEyJrZ43DwHbRrz
7BuPwhYTv82ikgQMHVadvwRq14Vw4TJf6yRf6J12D01H5haGzl2PO80VYHc87J7R
oKQpldpb5HVS8q86xQGf75TUxIOVL/h2oIa9+d6jj6t3NGDuJqPg7RlvzqSFOfO1
uy0nsGD/SBkm6DXW1lZbhmqF3u+RaBtFuoIU7q2Y5Wg5hRV8qvQazqGpHnKTPmDh
vRPrrryUjBwQKAzlb8ByIELT+0QnhDQ4OiRikE6TmpRl8MpJveMCAGntBiaJqGgv
tpo6oLbcWynqw2zHOqCMZLWOLgAMq22GXWQ48b1M/1D8fravm4il52znePnoxaE4
r1vcOYz0xdZVEAoM2bMRRPFnB3aZY8uVATwyqHxwDFsghL9vDUi1H248fOq8WNfR
RVq7x6Is6M9WBqaRPH2I1w+MkFudpVH6J/som0LTESqfX/zwxyEf88DmBSrmHUBH
axBomNCy6Ywd2r21Hk2cvu8mCaFYgrmb/yHmnCgoZ9ubgu1PX44T/zHpjHyZFBS8
sZM98mrV1ugEjC6YOKqdHtSyDRnMh2jSF5kSy+C15v/JLHT2Gr4kegM5O74UkFSv
bsF4oN+tOx/x0DOopV25JZxiqYm6Gq0JCONXBKJyjJrQ2R1K62aP5hAqhJwbdXzX
HjNM3rNRooprt/RJnS4SHcjs9a5DGuyHkgPIIp3D89HIQblISxaOpdaUOlt1DTdD
019ZC36GAyI0GuHHZC7eEKkVf66ZO3eVgM+0j3HILW1IF2aia0J1ATg8lSqYOUSL
2+O/FII7yQdGAz0boLJAVCLFC3IlkbCKyeqduB90+CgD56NCY68f5slAGgUiekRD
nqJEB18sQV5/fW+fDpJ+Zqi5d+dEQqie5p8uJjGfX38H7oVzwS34f0Ae457UdfHn
FAF1z8Ed1/QKxvtS5BJKVpDVwgMBHZBElHigE+NY4tR0H7SXD9e/NqeAxDGdwfQO
ZWN2VU+uRo6UrUqMU2xRl/Aip0HjI4Rk633DPRtscpctG01rDcl2XYuvSyJPbjf8
Fu1qgnhUjw7g7hAXF7EczdEV8UpZWYzvs3DHUOLRlSSYebO9OV7dfQorQqJhiML9
Dg5c64NxQuFpJfbT3ENGhE8a0qBzhRWaqhEHQbG8YfwyMqFR+UIR9aHo3oDYbHwU
gSs8FTICB59AKvhLy5lojeHdnhx0qDcZzXiMZD14bgS2xDXVePO43x+3ec6nACD/
LCCMDXdUDa6jdlPvjjT4jjHO33S+0Aw9x72k172akZDLT2EAHiLXl3Ob3cbHmRMq
4U2MdkUCfUdEkr6bQmXcqaHfDja514eFehCSRtCU78GLNFp9WbzqGUmU+4lbx1vc
EBgnG8wlNG8CNVGMrEL2yMkl4QZq7mVHjDl6xC8aFtgC1y+FCydlhwAK0fJjI+LH
TWWy+8UuwvmPfef/52zrL4FdzpLqrDhE27Lb/4KJ5Sq5Pt4X00nFindYkvDNv4bc
FpO6zezTHtkpQJo2nAEFqIAh0yOGdLcLWl3LjRIarxmZHRBSxtNdZ2USKJKP6TPo
2X5hKuEgX6TwM9wE8dJhAPgTlNbiwTv+i1cmFiuRN/AN48kI1IVRXMAYK+lhkfO0
uz338Kug6eA4ZXYD2uvA1f2+X/H/d/aBiKtoXqbYMDqfcXbYURiZtXX3RkZB1/b0
7aQR7ozhfBJkzG3Vng4ecvXHJi4AKgVfXk1OOIZ4BnsEygmOFEh4mtv3UFC/5rEv
6LJ8YmXdsWA7a5IWpjofEPqkwae64SRmAUhi5fM/ewbDP+QRhQTBO2nROdqwKQNS
Ycodis4L8ha2LQFV7yh3kR1Db11Us0jj0zU+uwRRs9bF7kt7SKo78KGL+L+tDo66
je+6N6omJLuTkqMfZePd9M7NslE7U/bcM3KOQi4lUSoc+hHKYDAhcZa0tGOzhlqA
pwOiHhIhSmglQB4aARa233GAO4wtT/+cesShAQuolaQO2rHZzk6AkH7FMunfBOZq
h7YyDMTGev0RwBD12f0mkA6LgupIf//4YhSNoGhOUyOsg00e158JQvceZnWHhBn+
Kj08J5Yrk+akt04pAG8kDKU+vbE5QPXyl8vZ7UiSlO2NG4cHLBG11ZpVbTvewa6h
CE0InMM9XwVGH3ed9J5IoCNOQip7Drq2yrC2sr2v1BHNplomGKnfi1NhKSL03Gm9
Ku1rI5u3WfLdDoZG1U/+/LuvETM3tDW8NuIZWlFv1qqD395LAqYsVfc8R0JDSycb
9X9BqyrIEPJGFRmxPi7nbJmRW/wYMwMFERwrtoe05Zd66dmYFV0//dBK5g+RwsIl
BAIOahgGFo53uqnkNnyxCRW3r8M0aoCK1IG/364I3keChir3P6QGS4m8m1idT9CW
6LK2X2TCIJcEUNLI0ozb3FtlxKE1F+J25mQ9eruz1MHN6F0f1WgFsX3zWBtOpV0E
d7xntHePhZF+ZngkBcTANFUHieZXLTQU4GAA9YFMC2hICLYaccNtmisJ8qaCNUvS
fue4FNlgTrXla5irUU0HP9dAx/MeF124Tqvo9ZKGsQRjH82JHJpICYE9W5dz9G4N
V6VB26ufKv+bh3wdeWd42NfaJuaRwJ5OLVhskNeglypDlzVPCz8+m76qvCJ3ITya
6kxz+IaXlmxrsOiJD4p2xy39ekbbTPNJev7RMQwouANk1xeq2tsn1fPIia9V5ean
m5tthgxUaAl5jZ04LYXxTX90u32OVYBDNxkwQkJJ64ZZKaGgje66kE3KyYEnnGg1
JSsy9EI28PqH1quiyiSnHxEwnn7TfYHiF6fWmCfYOps7JRAmH8yEgApK7OcsJuVt
6rzGxJ/QEpeJHjwm6+qgpt0QbZKc1nuKK+vuVLsarVslN3awQ0ZY+mlpiYuWSiAx
YbTwwq1rpf+YffEniSSv7rIRxiH/KLVox1L+QS1Vu8DiG9mQckq7oJu/pWtBlEs7
2bty+59uPLUlnhMMOZUYVLdrAhLVyehjtyJqeKzBD6G5y35Hqo9qYayqeIj9dH5z
AiZdDr/i+9KHMSZ13pilsVk63KgV3ulFIypnTbOqcdD7DNA2uCNUVTwYWhjU9m8I
+u4OpamQmmDQqPUsEobmhkynrnPL57eMlD8OFcjBw93RFvSTafjolyO+84f9Saxm
zvL9YFIAZByAz4qspE+5jradMeRon8Kkh8jpmAgcG/ki7mPLati1uMqPp8zY5KM5
Ay3i7v3IiGcN2ZKV9s83YWm/9GQHNw7hMFjk275s2RU4FSQsVf7i1a0ynpHLs5QW
u0Awu++SeKhjBXeggP9pWTaNdGDOx94QyQe5nbYmKuIqkcQ+r7RzCVEF53o5+5mV
qQQ0PZthk5aXytAIApiSYywimU7X5gCMElLfiUiOLhdpI3ZVW/AGcjTynAysjCzX
CKtod3bNlYjcC00ADdlFguZF4faFcJYGwLVtbmzQuhlDA/2UTpJjo/L+MADIwYws
aHylho69mCCkBiyV5H3oneo89gKedCb2S2F2DkG8hOsjc53q8ckUIbyoLmWbd/jx
pYW8b3lI/fz4Ugv9prMn8Ku4SM6cQgmqRyxTBxODxdzd1QZc0/E+L+9+djvvY229
cjqvHEOPGGqhjie0uDC7QgLMA5ZlxCFjGpuB5QFHNUFfRf1k7sZ5feO5+8ycYzZE
qKlAzoARba2iPbNazx4Kh9SDlXL1JbRvdzUdgUGj4idHNQl0KYFJ77CgGQZk+QBT
bzHRUHjtXrFZ5uIUkHIyima57+lbIZji2vr0P2X5D6Krt8+BJV2TVTfhs5Mu+np3
3cUrCE0NhzakrqjJxsC09YcVur92dEjBoILmOX2BjyVB/sHlRZXi3HT/oqbnAE0h
V7EOPu37NNVG0c67Mf3ubkCGm/AeCftnPF39ybf5mWJuUuo6b0T+bZNyZ3bZbxiE
7T/0cuWDOC1MOzbIMWex3lN9zn8QUG7V6aQBwyaITQjhmhUC29t5Fa7SqvecUXzO
ZeU+cUvpRV7DV/1LoUr2si36/NMDBYqcpyft+WT2YqWwx3z6RwYAhWVnzcN1tYzX
D2Co5xnJk9EzsNY2mwwV/XH2hUEwseOmpCtUvAqvsgZBOjA8Z9hsJWQlpamQ4R5C
1TpiEsQRvGwXWhM6pAL13gWWn18qEq7AFf0j/vdfHMW+3HjS62B/OyhnS1ryatcY
nUfN6UC1JwuGbeMBM0O5xDWxFmFqPNpqChlNaDUJcP2qzZR4uza/uAffUM8uDkfu
bssjToNTnViTwZ/snwHuJcQx3R4GEZpCH2i4dWLruUv3ekbCVfxc5tTS6Q3zkJAF
eTkw4xhWHuIgwAcpaPi79PC6RYBMyii7rwcs6UUwlbKOZDy377V371aDJlJz14Ja
7n5kU6MVZPizwh4udrE/1rjTJu8efMqPw5OgPF80TffPRq6VuiUNJPosVPIoBGTb
WpMMJAs1/rn3+oKoLSS8jNIKzMDN5jevTu5mvS92wMSL3QANloUeP8iYBj2xBu6B
QfNdVow7ZZ4IJLYcr1qCSm6e35m9Ms1mXrmY+XyBcDES/3Z4o+e27lwg55zSrEWL
MKyczHOwASMn3r1Okt1zTfB+STAFF3gT6WLMCatr3cl+NorQAVDJgH0pGVme8rQJ
TQ9Gp1H7R/GZW5dBBF4Wd6Tp/HyOygwsKwUV7SjN9uL5+rnCrPEIatc7CmdsBd8w
JWT36Sf7/hnUlgrrXjlDrBa51yCwXF/U3R0IMYgHqMYwDOw9ou4Z/oDeneYlWvtT
dmb7o89ByGtjW0pRn5BJspMK6hvjj0v7LSYDJDndXMKxK7lzNiWibY6vhbVlY+Wv
oArKmP0yPnLOwQtqM+Am+gndSZf6KfpYwVbQ1SkPx4Hk2S0kgJJupDc2Ln57BJdy
6Os2P6Vu3PESOt/M+JsfZ4gn0yWLPYTfjMvXUgZocPGnRuPnN1NcsxuJKmjldvGu
ygliyi6R+gTThYL8Zm4w51ONoRyfPKXt/1Yo45PZE+hlOYWJmwf26cg/RT0+5pJt
JmET7I0wRqgJxGCdgJctMHjD76sP9gUsxVbrUOy04lHlmUvd7Ut3qSovrCAYObMO
ccqi3WPbyV4yo9O1Ylxt8vHGS8GrRwmrsNynSweH/Yzvx1GIrKo+qgOR2WiCiwgh
dPMtk/UrA3GBsYckwaAiav+Uw0gKjikW26SlLjazGyafzuL85AADUjeHaaaZNoz2
uI45UNSzrGtHpL4KIiOBifol3skgRW64iqIuEy4no/0sCxJ1k0+ChnxxQtN8Tz/L
zWhcw5Bcrl1YmP/hIXbUIb59CCGxJfmeaZbWTDdUmD1ukhpltqUsG/ucB4QqY4n7
c0FMnY+mvY1aRnY4hi8ifwI3nh3kHAcTRDSLpYImjPIZFlhVQD7GcUfJKORQh0/4
41O5AirwwUCxp+H4MeXe6qMrGlhTRal0DEzvbl+7vfzlkS+GJPu6F7ZCpsmoTn7z
QWMh6WPaoLO7dqqqTEJZ3A24nsdya7YU/6x3Aj2EF/Yr+xh1AL/EBliW3juFxr3i
FPjeV8qpCJJga4SfAWMQ+vgjcaxv9kVdSbVocKQIrbKVsk1aPpYqvyQMmo0AmbeE
XHzmyJUlT8T9MVQi68rspR1yr2zPz/JOSNkhoSVxZj06cG8co17zsM9tOFTzXrEF
DOKuLDS++crshsmYO0bLyBAUlAHaY7UTkDCnBxsB1aSq4FBueFzwGw6NBfwD2Bai
AhaJS1opDarkieJhIXxo3Ltu2LK9FAlSEX/oXZorhnD1TT1DqkMJ3RYs4qsmzouO
FMH+qmfLPRQCfbdTwBeFxMaUxL5HnK7osfoL4qi/pf17j8ZRd6DuYpaRBbdPxgXV
kKjW7t2eojHRPW6q4UAiUVhezdWPxJFputXoPj5Xxo4WfSHMU7Y04k7OAhHT0JMk
Oj5qEuVOllYX/bp4A0xvVOteMWJwI38U8z6QQUk1CrMWfOeqeF6rc3LwRezB7pbI
c5SScxx4E5hINe0eqfNww/XsgHD6OVkaMvo/SpisZNni3YG8Lsx8X1P9HtMpF9cW
VIisjIdOG2mYvyUCEuo24YPz8Lmw0gjJz7MaROAt93qdQFae+VokZsOjz0rk0nwz
inpJcqD7/JG4am/Nqe+U9obPgrLWds7Q4ehCkSo0UzCK7SWmgvGCWV+AsyhWiqF3
lkl57j/9uj2A6I1U4dsYy8bFlGMl+BCt5ZuIYNoPCP+QcEJE8d3mVJJNPmE0YF9K
hLttnxYbXzSU1eCRPoVGhA8uMsPu1VQzWh4VSuMHd6Ar5ewKvd4CAQBQq5wr9hwo
/06t6mgxvWwmGieGCW/5rtsWX4zYcr/X/wBiWGUkrixDE8TaPFECzv344YKcrWbc
ShvCck0qGRX9GTtqgDvfRqc4NV1lioHpc8k1F+c3HHeUIh3E3eb9HKm456lcmsO9
bcu0pxAKdsolabOSEW17fZzxiIk6NM9QWkG6z+8+fz0Jdipkbnw8nGPuj1sFQgBi
rspDs7EQ+PMalLwTbbd+snen6R6MDcts9uXJKRvevo3ZP5HrXQOoZFnX/OIKOxEZ
ojcEK9nBl9YK/ZHTgFWf+WE4KH8SnqLhNQhjwQVT05fBenDah3h9MBJna65lbg4s
sS3DannnzfqJgTqmDQC+88FF0evEO/07OvRm46Rs75REexVlSzupjtCoagwmx7eA
z4cfFQTAMxB5MlZO+sZiSToqM6foRWa0r4DKVOrHwXeMfqD+aF315tRN8VKTESXd
sX7wVMFi1lV4fEbw+6A+5GKVpAE53oiObDqqvsCO1rMRPjd80hMY7iMTB+xh3NDD
vaoZyTM1JPG13ijjdvNmaqXxUazo4G8l0ImCbnjqD9V7w5ngoFAIFdSGUAKkoW/5
lUQf9vcwHmJxGdMMwgczhvjgNJe2cZnfCV3XqSeqNp9XxELmyD3NcKZ3beg+ZRJK
13P4iwjwDRo6BzGfE3dLt3miyljKzd+iZjKv+Ix3yLfjsl5gPi3ymcLtsXYhuXPd
1GYBpNYVVggIFHUMHsN8KRj3QLIO/fQU8wR05Q0DduTeIQMJbeyI1qLiVd6flDcY
8yHJCjaimtEFY+HXH/F6xpLK2HKaWBhoUMZfd1MjYs2B7b9nMxKg94ViVFBTz7jI
BQqAE9g7TICJicDPXzX5C7q4ODOgrG1BYYmvakqe6VFMxltP/rJH+yUNL8oHZs+P
5afdUMBrKnf7rv8KOI40l26xMMcep/bAMGZuphqESc9VwPkUxdVuJ/S6hm0o5JaI
PoivZF/sOoXD1/N8rW7OSLo52vLTcZV8wT/AC7MdPV/P3t9ULLcr8qcUKBYC/Zzy
exwF5qwKQI5qpk1G5+a7zYZ1cNgrus3uRt2eYzZI5m3awG3ZEhjAg51yeNLhcTSR
ZF0nFiVG6k4QaDetlJ6E1qLJ2FsfWZylxPkftucqadagYUfwlFTBDGIliQjrilxP
nfPWa83IOk4XhXCMmIhF/8Gxo91L/16uY1keshP8HKWcLGyUOdDhz3ENUEC0UBnu
giclEjg0UEqHaOdfvCmtS4J5i5mQyDw2gSY0gen5mUyo7EZL6h7xK785+uzNq6/x
xn193Ozkpfvc4PIIwxvd68csD/hNzqpSpycibPyKOfaX3fSOy8nEeIO98aO1zDYE
KRQnu+mqmBVraZxHOKs8vR7O7/mNlBdaxwPgb2blVdLe5IAi0z9CjchjX9VFAyiP
+HUt8iguf3PqTXW0SZgQbxEaJl6QGIPGlq02fcUQXRKtKlSajI0p0Ck/ejtkPmkR
VJ6zTwXqvUg/6Pr4PfTnJGyMFyBMee/HPOpP0iugn7t86yYl1zbKIz9cQmod7r5D
vCtk4jfddFvVT4TVkBxICMO5MvOJ6oxi9pCGZEOOwVzvY6b5FE/E0qU0XsHmb0CO
o18+vBBA7UaQ8FKVRrPoV3z7nF+FhubDxjoEOPp2JppxQ0creJnj7BW47qbBDQQP
tdLMXELHrqHVwVgcWXgIKLwY30w7OrMm83yn4Aa6/xoAw/tehW+0OR1cLGe2h+fe
iy3HccSPhPtuQENtF0cmwaMR4bS9TZvCWcHkSfXTBcQcg92r5bpeLcQEF8P4rAor
fjqGlbzRrmn9hN2X6XSjSYIoGavE9mHeWNxyKa/XNpYyDB0C+fgwDfRNxB6+h0FP
Y5S3IFMh85CfNTlE288hB1GccpUSDiUp+6QqOgREFHjKyLNXCc/ISfQG/Pwpwpdr
UOTfihrvIMPqI6l50Ph8fo+XSrqxXZcf8hMxKpoa14mJujy1Gmkx5ar27Wrarbl1
XwQYI2GAju0XDGeAKyonISK1rIsfgEhixxQFbQsg6d94m23Xcx4HfGPBCReNF0YS
KrbOPvP/NPRVj29drSA4pX6XZEYxYOq6XllwpFiYR87POWR9zfq0H837taJzZKo/
OW5YSAA+Ni3H1Dbv69GrCERC7SZtsBLGpbdNYuseRuzMEZ+s1+DLjkxyJYkI9Rap
X7bnHm6nebN8qiABHrYSGgV2D8YzMg4jSHj4nhnrwa9nm+kWcHPgOVI0F87BnEGy
CPyki9jjtkecx6l+Tyl0+sGL5f1mTA8+rrfcYiGgOpVvjMT8iEyI2TJZ/EZOK6S/
R5xr1lpf/4uTnCcKrAnMQEQ8PCvMBiIaJlP4de7mnNw07kwtNjj5m/lHCqjyMZNK
Ylasd2lRrBhXodVRyDC0sb7WgGvyzNj6n19rvniHH8jpfHMLso1n3xjIz7HQN0BJ
wVG/C5SwCRyVLGQAejWSLTM5Pzh1Frd2Qm4x5Uyyaqh2SCg4o7GUZ48nccFbnIEc
xJi8tUpmy+iHjpvjlBVo+3JeWluM8z6Rz96A5uzWuCHTY4iPPzROrlY82M3fdO6e
qLCf3l/0e3JyqnoheIceHRIADP8MZdLeWpAZwUADUfktZr8CcR8hrFk6tb5lmAOh
H4tFhsWz8NYlcqWcI5lje63F4xqWM3PCZXdhvDHb4b2H4jNMG8+njIpf47L98bnA
jXGT83DOyFDid7HkB4L97hYVgDkzwHsC8uneWkERHvaKtvjfTIH6e/9sp0c2RRCa
KbOalv/6ep1EFVOWxQpUT1bP6SEGEyKALcKp4YGFNJVZjir9avHCHb0FDTrWtELQ
MYstu0D1ISCS59o2m9vsd1uJBkaE9qEhnhduGoTiUxedv24BRmXPqgXBYIH4noiV
gJPUoXsmyl0L0CXZZTPJ75HW2fqIbvEBSB2uPJbCMB/gw+5xeUitMzbcupk2wVlj
jGCVOdgkVBBNvJbT9sUThmbdTLi5HKRYZu0SFV8OEPIKCi6+uRU2EUL4DPuduK/d
inouuBo8OFhD2kgOOSx4MpgWbsifkYJIUSlZ421cOfL3rO81/RIBhFevZmUKSEHa
yFJJAsaOrT2z7Y35wiC7aSt0TpT2vOinNMR8prOhjsYbQKXgnv2oUGThssWNwpVu
MzsMNaMOf8JZ0IpEomUvKgTVufCZrpORc6rEyYVyIvNkvZOa5w9dTpPjqQ+6k7Ug
8L02MC/lu0+R2peXf8qUQ56sCEVdkyF3yEty86d2R7YJpP+bD0PXFoe78Vm6r4N4
fw8lPbh6wRzD6ELLELFbGwsdRCRYw2m2YWDvI2PH9WJFJRTS5k658D2uR0HFhtg9
4QL/jvzFPoZE5MoOc7cnSYAMjrhgfL4QUZDCA1tHsSenPOogkDdWilO0odQ6FhI6
spRnrzkCKaWHtx62JujHPfHmazZL1r6RLZJ0FMGtwcMq4oTyhenmqgWF1itq/Yyv
sG69EllyrYmrqdDZZ6AFb0ybDtT6N4M2M49d5rHoo/1STDMJXfgfGCrk2kUlUcrI
NfmhpydscfkNA+rv3EL9e6kyGzrZuG/yAWAsTmwA27zitKfXGqGxsGVnVQMTg7Mn
mwSMgfqMhiAlb1zUDne4PWSyI0urf6bhKbxH+XsFZkk4p4paVtYKPL2fJiE/Nxzj
etk3MqEs0witRDmzp7Rh0gZ2hziiNTK0yEafV6RKebaUNvDUsoCpba9HslxjnGWU
FQFHWxpUrNB7fjS7yBSNPr/yYKQQlnygXDXnKNOnDTbl8gMhp9M7KUx/CMH0Jazk
dBfZaVFJdJVd3HcQ4dPwHI95pnInpU1tNfFWxqbJyDjU92xwRDbxaUNG4CmmEgLP
em9lcU4F/cFZumbR0gktcz340+Pk5XGslFHm++USs7u5/OzZCp72cpBCov1akHFH
yY7UooYc3//BuTOpTJSISja/NF81PRuj1f/EYy4YEj4FglWXsO/RXAO8naeCDQa3
ZgAFZ3GaOegDg8C9kMBhtWoL0aELTi9rP1nxSyi4ZpRxUQ+gU8902OHS/8YI8x1G
5/19Gyszfas3KjlD1A1ONvWm7geE155bAp+2416GnQkJ+zWFQkCJU2ZM42fRt/Yx
TKygFwDAG6tOwmCRWaxa6sbzUBmDZxCbm9GlshgtopgatoCweX5bHsVbPcTtotWR
uRjGJhZCMsDA1AgjlLMkPz0shX4/hLfTGcaFbYNl9MdzI9WTDgR6FxNN8YNItsdj
nxJHKTKiIeZOMStSz5M0j9XcYQCkJCneVUaixFYSqoFfoZACR40PMxR5sXcbyRUQ
mWOsc7+exrj3+PrBXspjRXaycQmyvLQnkz37HGjFSRyxVJMl/KUbl9X3ypIh8hOj
vn3hmVZwQfmVHUAxBjuQBmR9BJhJUYmz11GvEAHj4qqGWN+c4k6TFd9bEo/Yd7Rv
KnVPrV+VPIR9GFCqXYkP0B+HJOVgHhwk0RtaXFu7QYj5wnzGNh89oLU+ecjp3amI
c+K4lUemW9KH+IsbsqE/0vQNXcR4zn7Fwsnh/4f+tQ8clzw684OzkgsFIo309IPU
qd8z+zQqI/YWlBWkp04EvHW1uX8Cgx4fxrl/7hNAEgvTl+1xvRc0x0XIzODTEb7k
dDDS2X0TX1jmLvhFDCR856+8T3PJFrQbtOBPxd/xgg7/qxIhYgTSyIY1siraAdhN
OOBeLB2bW1jPliS+n9s2XjG6DiiNUpsqK7T4VAhmIbxy4uZK7UASE6H7HlL8B2L2
/cAOJWTTNz8pEI3ArCTFCFE/07Znn1ribrd11aYGwsuhupcpew9xA/FOqwJ7itNH
a6IAuNRPMiPWyYbzlruv6VwQYvyeaDZYqJCawdj7lCeXDsesnZ1E6BAOmkI54wl5
ol7/OaRj3ykoknGzmoDOkUEhPwQ1lqZxEOOowYi/+qxy+Zg+0r4qm9AVWidlQ6AI
/RVnexuWOY6RBbYA2arEtYjbwoDgfPqvXdw8FE269ptwRQuiKoTRN6kohTnwwk7A
JVUe/v2hHBtGpgSUBjIu0NN+6ihLYhWwFvfGq1g5uq48eSc7rAZpwUUqMM8R3I4f
OufEmp0P7q1I/WNt2ylZ3xF3ANrB+mLd7yDWvm/4ROc/NRxhSoXogJVPb966NZto
G1zLIvYzczJxCrSAOXPwZm+5Dzj1PGIBzIadEVKVJO0lfiQDMNtSgAwo0/q53Hrw
g6GZSLix27QR/YQoR0PV06ZrAM6D9uKuGTczby78FNxhZXR1+gONIz+EhZ8g0nC2
idBOMbgoR/R5o0YYx1+A9o7OcJeWviTB22g+NYaCegA7CFhwYjaKbZgQBsBqVB7K
wadxNCGbNXxE26tKlJejE2XW5s1KWnSnSvg3MTsJ2/QDT1uXoxLrVP+4kNkGb1q5
61BIOtr2DRH/hNttKallcSBItr0ltBqYwKXaugAPM3pj9XLYTStsbDgOcs1mergy
nx43on5GhKfDvBuRNwAOb/qSJ3ViZ/cPVDRfBWCZ06/vzKCm5mBC2JtrR4nj8oDd
qsnUCsrZLNIBFhbAyIBQ8A2UzLbDkthgbFeEpmcTs/jpV1k46mzNoTvTn2hotrBL
SqlHqIGSYb+3ZISWGTHwcT6ssRMJv3oML9IhEo0CZ8ZyH2hkEaNC+dHQh9OY6zA+
a7QZTuBD/9q7gdxsysnqPogP74U07SZf6fm1S/k23V1lANyUmY4JWWZjMm3Nsxx7
mZlVgSEgLZrd1Oi0sao+HBzmLdF/kO9A9VDjpiAhJc80+q/kNTiCqv/pc7NKve/d
wcACz7HrjQk8xgOTN8Gm51ipPc9Cx3//J2+Bv3YyVI6dHiNJ1SdBIL0sXUpd5Z3f
CILYCDb7il3qdskTYzgpG4okTcy49yNSEJanuOnBsV2qLBcmhdeAJspJp/WEMqEr
/zREqBzAQoztn0Q08iEIOYT9QKfaAHyRM9X7Wm98Rr3arT4Bw/rjs1S/n6PDe+Ga
w4dqV61UA4nyR19oSwERmsYxcKAdihRyC75ha1k/dWg3P2gTPOl0jWFD4fozYLGe
VEoeYTN6vyMadC/7yQtPJdnGDlFJs4bXy4AIINH/l2UiUMYxKSc5rCXFSL7LZg8W
cGh6yhTlCua5RK5qAGPSs/gSB6+vEYfvdOqBS9Wsn7gcR+Xh03WkNVfx6hcdwtdK
pEDYokD8Z5HF2rKtjRkRU/PvnfADPRvJedpJgukuPM7CGqpSa0HuGQaUcEzaNyHZ
cUJrtOGhs+fB2lV/0RwGh8IxOPGwen/sCOB0GVwQ05G1bUok3tzxRMSAHDPkMd3B
4faVclL3bYht1N9HJhHiHLRTuv1FOiv5AAvSGertxLUxjqJZNIcrwEjKcqAShrcH
G492A2SjViaHEzhH0rmDxrHzAFPo9d6GuiOImp1/9lTB5lfv/j5tnhlKDhMebmNA
6U/fF18liFpI/QP3PKyiy3Dq2d0X7R/95ROabqfQnW9gWEx4OVoUCn+anaGIT4qE
m/RsX+cHYD0PSDyZTRYj29IgFboDzZsqjkN2gUlXQLKlQgRBiSmR/uErH7Mz04vc
XkEQ75x18HbIUkrVA68+sFXpbC2dh+SLfqXedjwJoWK9PCxctvx6NWedbXPsWLOv
bu44ZyS3DP/NUXvvo9ixOMtloLzbnL5Sf4XyivcMPkf5zaBPmSOB0oAv1vv8NKCQ
qU4RDdZkpgJeZT9wTh/XAYCBBNCRO64NJU85qP+aCPUHmLVaEyRC5VnmjV0gZiZn
wRCBPsX9Bi2LdU3sFi7H9tvFC8w/kgZIZvtvWD3qvCB8E8200546U2HV6CsnDK4v
fnLOEJQKHc22Km9cwjEfHgaOYRVhu+3cx92U81Fr5e6BqFqjc4m1Bgpz0vhCf9LH
b7TCB43oNeJFKkTtlVAhXPIlQvQMnrSOHVLhDsOUqIE/Lkk7ZTZUhab/gYNBurob
Wwqv2aR4UG/OrwpIWyYndTqFUXGouaclCR/1/z6QaCULDH39YldLvkhs9Pty/CxR
H+ZBJXtrGtNJ6UxghefTe09YiYj5oRVroAPHnlCaVH897Yiepmxf0rseu27Q75hQ
JK4a9mU+t2c8FMQD96Pr5JLn+JQy1DI8e6MyJziENaxbIJ8wPYSZT8VBSrrycdK3
8Fm0PiAL6ovgcBlCIhWB8bLw6n86W/pp6YP00J2Ijmll4qOHvp7hwxpkTiCwKN+A
U9jNfX9ENhLA0y41wi1TH4Cwk+ltOXiowc/Xnh2pBPX250o9P6QOr7rXqm1MVtEU
mtSlivpKv8yOcndblaVkck0ZK2FMrLoBAda7UFTLfsLMj+PBnTPVMq9Jej+tyJ3e
2tHVUeX99POhVAltL9e6q7TiFDicf5qTJEb133LT2gUOud/q6xfZM5TSOcdDK/ty
+1n5ByVVd5eShmD5YtVEBvJAyT4+ZCkJrDqdGEJv0ukHwY7h0HqoFjMdJUMeB57V
F//V2NBSJY20wH7bUkbZeciDux5irzqqezQ5O8w2umA3diVXUAjYUNL/khNFQALu
Jo0MhFe+8L4nWbWS46mqYbhZLTrfTUqLNUTmcm7Hrm4cj4IF+H2q4saam8eZVgn/
w2vsaQIBqWzBA1EK4OhO3JiwgzXBrScwBNS9BWRIrVO0kuZQnlX5yOmi4ksKVHWx
FOZgMblpB9qOxMM5IA0cbn3gO/tAUZFHHYoobcvoXfk06OGKTTbuMFDBpfKhu9z0
xtzMEmIoOhMJz7/yGOzV8mUQjSfpSw+q2P0PYEJCfFymD5Kjh40KUFR7V+Vtlu/7
KZFzL6dM8GEh38C2Ky1ohTNIt/XmDl3HNsCjKtZmq/TxdKTNzNSpMQY5tzgFoGcs
TlpojGOW6KB32rPqnUTqoYmWwwgSntm37tJ1IJnOV7PjvlSIXNrw1hOTYlYMJxec
VXW98c8rtB56w9JUIMGmUZQsKn3BCs8SkEpVw+u2vnVwwFuoaDZe7JjdFIrLv0tV
TMfFOOGAS+GAjCOUmjtqXpBzUd3Ig+NPiWsYwBzi3Hs/6RsgsRceVGx27aHxUE7w
hoHLpvq0zQW2gDu8I5GS9RiYxeAvNZ4Fgpv5OzNdsRBXGq+ZjPhC+KHf21BlAwW9
YgIhsKyXc3OIPIXvpKlPS3nmgSYBr10PIqz8nztK7xWNhNwhwDLjJd0F3sz64Sav
hSIWKsjck9ZdkRwyPe/a9pL73m9eweblAp4zsYY9TrPrTiSOU5BQXJQ/qzaDhhn6
p5xY8JmmJOtdNuom8WDzzCFqrLClyoqTebhWTAPB2bFpSu3odz47V6VVPCBerBhY
+atxCPfNlO15lBlm+4FA1M6eyetzYmrOU7l/lvjZeepNnxfIvwAWg8U31yUK2sYu
bQCMC4e3eGkCuFQwoHg+Gsj4xMJUVsnWxVwxl3gftvA/m825AFHrDW9xesFFAq5/
FMzNX1B1F5HYm1k0HI7hlhPYgiEzkn1zbkr/YB525NlCChIr1BuwXagZqQzI9z5y
DVqM3Xr475vjWJWTICE+ZvJKk0tWMqXTKme09q129zuaKh6NhbgUjTKplQEmU9Cg
em0+HZ8Q9IwjCxOoYxBtvIU91EvGEMiOJvJx0UVDzis/LJGsTCDvABuXfKC2slWX
qZjlddTHf3Nzqe9kGcGm2l+WEeszh5s4hoFy6jFjGhIYd/WpiFsyeCvT0WCm93CX
rQsSjDib7008cJNPjb+3Vh4YywZKMgZ5TCHexOLwRnU/VusvGnIrLHdqrigHJV4c
7+UFcWajjgv8e04VdQH6agAwhcnlo3hrsuBEKEvUI+b0xe99YVDvlbi83qmlVWV/
WYwI8OPgoFDZcWM1bRdzcvho9bMoUNPqEXta5Hj6Nz0F0Tec5oZ3q61AMtq9pzIf
6XcTiXIo5SztKyaBHnBMRpFBC6DSN9xULuF41sE7D0sQFF61VlEeUbqsJ/Tz+Jyz
/604xcECRheUomeRErh2QUe0RgsqFclESzS9cpbNbcvXp8cIrtrcu7WWCox8seuQ
r5l+gAnEZkoA97R2/ZlxNK/tN8tZO2JGo99O5IWKFp8OSZfx58jMLaDgOh+8on4s
AwGWW7PZdwCj/4n49mM+XPNuUZ6wj7jWg1kFyvllgcijqWi39aDfS2L9bBjsw5Es
udtY64g7KAgpYoUQxMA5aHa/MjleRHX7MaBkUDNdPlu1SU/YRwwoLd4BVFA5961r
BUz/UaEimfki1K70Da/PscdjSwTiocKepzeKgGq3OszMxyZCUU88PMj7cpm07sqc
4D+QtGmawKxsM9k6z/nJmuXK1jBnw9HoCBCLIFbmlycbmtBB179KoSOPZaQ3S5vk
oetA4fmCTp9Olqknnvg85adExg5vaxf5p/gqpC5tdmSuJPwVP+wC4F40U8sb5K7i
AXg6S1c/Gmw3LdHHDCixW880ss665KJvASvUscrfnzyUscXrhFtSf/G++JpQtRZM
XpzG+j8f4c1g5Ujx4J0vfPqdbVFOiQzrOh1YZsNs7SGrTNlgAxxI1sctIlt1AfL9
KEwXwOsy2f1w4+PtnonUD5hg6zCivwbLky/7I/cUhKXDFk8y4n44kHo+3CKqL5W7
Ino2nu4z2tOANjY4vsUXYr+umEiRfci4gwRd4TpYvaRzxPlzBVE/Ohu/BrMg78LV
mJUfyTShkcRCBO1dZuCX0hAfmEur1WJAbmignrqhPNR1ZTC7hZlg/kaWdV9xVVXz
icIAviGk6f6jc+xliYeq9WWvYfcuG2Hlt6aXOzOb8mt0gohPuggoL2YhjIwPHIR5
792ZR4dKXsB0w/PmzTrcYONe/mnCC1hpnC3rwklKHZXGrbQWr/6EBkkxFsVWpwvx
AgdzipZDfxO1uMXzXT5rgVCKNhjNUibTNDdHmzBS5Pi+jOtqVMfCUrWcqerzakJb
JkCmcd9iQOBRmvFp0NwUm/AyDgcJdSSkdXra7x+GOfq8No76dqvzQuq8Tgm6Eeu2
AkPSCxt6LQOipn81dvQcS3Or1w1mqPzRYCPv++O02FIQkYjXsAun8Q6HR8Tv9HOS
ojtoe1JoflVLlCKoqwyX0IMi7xHcVaF9hGErousUVVDbNA9vhACJULNx/u/SV5Xm
KHR8SJgZJomViIYAPcHethe0L9X7MFxBvt6K9VcE4SmRe08lC43g84NPmV3tsA+e
mF5cP/DXZaXdYPAiAO9h+JGZ9SBzlCJgFH0A+xdhdqzRXREVHZY22zqCG5HJRrj6
aAiOYjQnW/JchscXLDo664b9iOmTWb3N4Cer8Q6zEYxytIKDVc+mIMpuUDlhCb6/
noEO0Ayl+eomqCVhdRQteDKqmv/diPpyuqPL4sDx4xJLcwSlVNRTfbzUN11GzSGy
mAVbdPoAdQfpWvmxgGELTvYNGA9FU6nOua3u02Vl+LviRFH2rlMym69Ne3m0x/L/
HsXPv6QB480IQDJkrvknG22l2PJpmHoZaE4UKDKNWp5vSgM0ITx4bvSpqRKDT+Jc
BQZ68ySyDq5zlSz0q7Hs60qLs6z50H2F0op1UYdPRBErcfINsBPIOy7eH5vh0ElR
y3rj0k+F/jn6y7rQPnJwvqgR8M1RNnCjEONX3zY1HKjLqOLJw/4L9rw72fBdnrr8
6FzJjrPCzf3K1OYtEG6UbRphwzoMgbQzCvHiW/Hb5xTkR786kikakZ6scFs7mrPI
m+hnUdhcXxLGOE+pUhNZW/nqIQhUKdG5z8xx+Jiu/2TBORjVhwZkaQ8tnJ5Kyr6Y
Y37R+1Iac1AgT/IZKOZ4F8juRGfoxq2HwII3SEh5/fvYIKntQOPa2uxcILJK/IvC
6+d1/Mu2XM6cW5huFELjsx1HFCzS6hXo1IZcM8eJdgFG8j8/gy3kLfUe3MOYDLIk
66DtHPydInlYuiF6tBHi1NAdAarN9BfNov3g85KE235rCoh8vFhoWQ4PjUEGfzag
S3aOp9w9mIzgqya3+S6zAKFdAC9gkhTCJXY6m2ZC2EdhVBBroWZjqiuYCUUduBrQ
o17zER8LvJ98EvaIY+rM0DtTiVQGfB2+js8aBZI3eqNs8FENgSjih78Yoqzs7FTj
rLrCl7dAdPFNhn7BAKFRb/2k6sHDNmKODnq5IJNDGe2z7kaD1WOW2A1IbQR66YvD
4SC/V1gvw3H9p46MHVOKdshbKFr38ujNUYHfcgELzkPnY9juOMoVJ8pRS19r33/h
cfZs0uDaOoU1EAjW6AWB+2ycEdEQGwrpnNP7PnnqjKAWqHggIA/jxVZYUY0YOcjI
44eEcy1JwPEZA6CUCIHuNgo19p6diVsBJKXT2/y089x3FDcglT1zGFk3ac9JlC4r
dnuPJFcM1g2gM7f0Zet/3raeUvffUYjLsy6/Vfr4I/lkUGAVL4F4zNTkLSu6euna
4cveuu7engkmbSpL0Hgi/h0719o3RIV6LzF4tr9sI/UM2dH8R8CDG/SaotDeJfmP
vnhwB58J1UFETdtXUmouH5PMdBFFoqEZ/aT90mai5/mBfyAlA6jubVup7qdTtj7I
hRBgUQUdPwJQx7a2fiSMqzrmSStqi/DbKqdGpvscS/o8S+Ql7fmkE0il/9LLhFU6
SCc73F7smKAoqjH/7m2KHteXlzGV0IVvaVPHzKu5aOEtkVub79rCFH22ytqp4s/d
6c3eMJZ9S8DfVMsVob4k6cP2e+nncyI4Fg2I8k1KHOzZxZE27L/IhswMpUgIhjyf
OLrToa3WgupJwtyOGBC9ZAZuaWSg9ImxtDM7YbkOLXZclSUEFZrH8vfoYjz6c2q4
oamCt2EsVkVABTbm02t2lodjxwkUqw/iRjeLvrdy0fZJL0nYcTXx2FXw5YTr6F1y
+VAgwfNtObFdEAUfAPZNCDOApy8hxH+21P9dhY1Mrv855btdUQsaCfcWeueuTsAn
LN0qVxtMWKKwqJTYCVhJ/5zg7cnd6sESTPovl5k6hfPpYlZ5hWdiMlzF4xV1CTQh
eYnDV+0JHNusTbNt6UoDDLPtey9iJ6V63W5dyVbgCp5ZMc8nW6I6Vo8FCmz0I9Dd
FKnK6XBltFpptcbuohjQYd+aNpVyOyMgsi+Il2u0j4jSR3anXPlyfmEk1QNvsDao
Yfs1iBdSrjsRTHd8aWirww8HVB/EoewMng8+f1eCCcXWnv/sptq+5968V9+4MCRG
EpR4HGSpSrfhVvFEFrfCH2/rD4HoNknf9F3hicFvNR4xlK5qrSY/Na2ftSMaEbBj
Zzhds03keEMArMYpyh1WXCjU12O39atTxp5umyyhx2vTwViQ1kCkD5M8p084D2aX
qoiI0iMfoNgM3Q+rJor1tQRbmgQ1+/6YWBd+WLCVk2sNaBfg1sLs5rtECeuZg7ER
Jxxo4/hhJ63Z2JzmPTyrG95qJr/P8D9vEAj3okCjGBE5LcseRI2Sw8JKj4tsMunA
WB/0COvfwNO+bKKALdLQbqNPpFGMUysJFk2DNmVqk3vLvLutjkVkLBigNP0GR7eR
EdcZkcEIWl7WuRB9crT2fOxpQNIPdSyzj45PS20Z3Jg/VPwVHY7mGWBPZPgmGhjm
jhM8Rsxj4yVj/7pLLWhQcCPTRRvLtMMNE2qLnC8AxP/ATTfsvm4V4NNXcU7c/mdK
0FpxVpmn6G3LA4h5H0gia44L9uAyfu2cIJS2AYSsze+ZlnJcA3ZV9EZfwF4ggOmt
C1VpoLllZRRSkOjRpYkq0gDD0tY+fxt5yCeGrOIokTjowMWYOvc3dzMN64FKFP1B
RTFL2eOzRGreUOf9XsmjxGpQB6Tx04BeVMZq7ocL0ozKsrG2yeJqd9JdRJJ6ADXN
71GX+g7aKDbdcrW2eY5Ldr7M5qTcSY89XQMSqiDJEnIzGEHKmwFerFslB+5obp41
04rCxut57Je1sRy4hmzm8d+uzNmWywlb2Ra8mPmalbeiYs9+UphUh/Vt47oE2+5/
3DdO3yv68KPCfxUVNGng0Ia7slqUZWywAWDP5I2w10+tmOa+MjPpZCf0YOMvest7
YQVqhML87YDb9Un5H+jY6/ZxX53DqkguY+TYsRC70A3XZUDfCbHKVYgKjWkSOc8X
2d9Jn0T9/JrR2WNTF2fpJHhen29TAgAJN/BWDJ3f/XSZHhHVX0ZWlUY4JBHwX4kj
bpfC6tycre/O1Fzc6wu94jcmiQRZtMZBR0HAywVsk1+eekm1t1GqOUN+jV3peuEY
Q2eSXegYuJ0DHMIXB2+Qpcvs43ZJsmK0IuPIsFDnlM6VV9Vjc02/cPkNZ9Nm/Tut
iM3Bs8f+ubgC4sQtPCPBSLQ5BbvY0PnOcRXjNQ4yFUeVKERcPDOnOel91typEtZz
yv6LZyE3HIOM4kdeIZhXcvcVCL9bAtxVnQbXJYkjaKAYBB5YgqDuKUuXoN4TKL6P
e9eL+LfQG103xLmeSe+HNu6LSuqaAJope+qh3FfkbTvh3lk6kwmuX0lV81kds5B6
9SpWfEpPyFYlt/ZrXJU0VuJ88AQD6DqfiOL094VbxN6AvgDguCj0mEoyGjiUBQPg
POZGQrKAjBQEoqm93/md7d5oYyjsAdu0741TepiKBpu2seVBkgikp1LVrVyjGA7Z
oFixqARLGbmjQr/O12yoqw9D8OtqyG0gA76sF6K9OQ8TTa/6m3aDUF4nTVBgCfST
F6v3DGHC8CBiLlw7d79z47M2UfBF8rUZbjUBWlgdbJojVXccXyCRwHmHNqFtuyoG
Ysin1qY886mfJ2zNAWH7TWbraheEfn9/iWQpJF3vTIgQRVWyxmvL5aHTliVnPnwx
Hs7sQREFuRWDoQGltrbW2QkltC+jzKDv/w5Sx61dvDT56op+UbFf6lVhDknsXOye
gKC2GxBanBZmeci5B/7Fp0JTuRLf12olWs9CzMw0sbjDTmD4flgfu6a2dzLyO2NA
y1dPuLwM5frigm6uqS23f4g7roVhnH+qoM4abTAjHwUWllnnVf9awuqqBRsT/+hG
iBRzq9X3XYX1UcrhxSewzC7T3guQ4sX/rSoMmpSIoSBj17I+E9NdIuew82kuTGUH
i+FUsjvlpEkV4B9wPrB9WCNi2ZXqSYuNsGdEbNtCU1KIvj/c8CNZMcZ3PcqVCHdG
/y5zNiDqWhF00QuJdfbeXoJIhIt/fyT/Qt/YFVesUHEQkUZtoAo+wreALISPQqvI
Dsnz3mQOUMH2lEohutSp//yfmX/e3/jqjwmGyTIG6wRmBwyR6aZgvsrLfZyX0mYH
3lMkjP2Q4b7WmHiT7tNJBKV3gnOu2Q4x8ggKt1GyeVRh72PcEJmc93jzfkVxCTje
Ca1KtnuwT+w7Whris7GbmOhMtpJYFOhQJwOxPYDUKCueefbu6ClN170d/3J5hcdS
VyEPHoK+uPC+NoLGW13HjPpHN9Wxr/1xLKK7/EPVgCcP0erQHaSWsjOpYYJKjhvk
RX2Yx1v7ctwUwcBnBDkxUW6cj9W28v5ZmMXzp1AFY/9uwiJ6ndFtqKwUgRIgy6DB
UbjqMB8WX0vO4y+eOb8wjkcrwKnTONTmH53v1CksElYltJrAwbEYahZJeo765dFp
bKBuKihDn6LMTEW4LlVTiEklXKTQGb9ulVfqaD8LOqgKdBX3T316WfNAGWY0t95D
MLxBrURUE7qcGxd1DArKH42/OrxeC3AbM9yu1wM/oFHAwqohjHsF/dtLfn8Azmhr
afwjp9XTjjOSMNoZpOZOd81HktH3fYLuFGY+Jn+9PWLfVxpZnCloTxxHXLZ14SPm
y6ml0q7xa5sOBiFMmcTM5zciVBQYc4RDTU+3f7jLnERFS0q2m5WNFhEVx3acbxM4
VMfbIbEEwMzBVU8OuN3eHX9ovRfx9n02+U46OpOyyMwcgYP9FsYo0tKPIk2unbpp
oqYKcACpNKuA4Ap1CNRZxwvkAa3awymEccM6dpbQgdb9s57qlOyBW32b0iDtVxjr
YjNCuVEReGr2NPylHA+JtIuPJGv+n3YiTPal3JRY7WtLcvBlH+fHpRZLP0GmjJ/H
THE6+r3ABix7q3cDmi4Qb+AgCJWXUL2N0hRk5fux2KaeTOKePocxCd2vEakIswzx
6xel8cAkahCzeIVMDTPp9RDPDQv4/SCNzVAqNESRcQmB7xd93m0Zg+En/5X+Md95
qwqaoaMGFJnVL3AKrh2HPyFgEWV283rPcqMhliIuFKapmjgkJX3l9Yj7IaC/mUQT
acl+QPjI/I2wBn7YjfW9KffZvUsBkk3Wxh3ALJQIEUvQtcLB2tWSRbmN+6DSvQZv
iTjRbGXeBi8v6pq9rYY580sofkTOWqcY01+5vEsqtpKOGRsEMHuqpMTaeEt+AWit
0Z7Gw/r2yu8gsmCx85zTar2arhIlnDJKRo+sWNDhDjIrnYkoPWo3DD8Bc6VesbOm
ec+rQC2jUXnvN/64q8YQER91yc3t1sgO/uL2p7KsZ5vFQ4GxcTlGDhL5F6VUpDJJ
QDpAHvEJI/SM/7i8oxZ/zmtXiHQzhJ9GlP7ix3Q0JhCrPWcCvvO99Gr/a17zuEqM
iSZkbluPtrROsqbxQlVWzW9QgruzuBQlN50AeV4KO3TZvtTE/VZu16SoaX73VlDl
nW30PB7jmO5XOeshHU1WyE9XuJMHJmjlb56/G3RcHBiq31Kt2uDI5n+mzcoDkXcD
ix0jg0iZ2PIFLJnf42p75ifyx3bcLXCGaqonx/b/vEBMlltu65wisDctFjodbf/C
neYoBzaW44uA15M2WbUBGOQSkccEPq3BmE6Qwg54ciZw3lck5f+wjx9y6WvICJ7V
zACBHa+musu/TEvgXyU/TO8oYRKAGmYV2oFZgKQhTkrMdF89c6XLF4cVniKffUFg
GK1VAtups0fowUaA3zCFD8EVWPma6GEyAsiwo2qvgJyq9YdONgc1jP/4G/38q8IQ
3oMbLPG1wQ5ZBtB44HISYql+7pQfPAN/qk287vgtvsh3LxoJ9G6//CspqamA9eUl
K4WfSf22aR3X4Mqw3AJ6kyGh89S36RaRUOJ4znyDXwEUEy80zg1Thfem5UJtD1+5
YpdBwqQPWxk8tEIZ23jgeEHUgwUWOvrM+Fb22lw8mcL5pYJ6H9kFskYSLMp+R+Ys
j1b7sJqfzRuQTR+Bp84nI8HgpqBX+5hL5PylpDuGCbZd5PntfNdzp6/fiW+vnGVK
DDQhQAoS8i6E1L8eL+hynPk2M08VB1F6tg7j4gDEjG2YTjiTxYYjFGmGQpFh0Xnp
DuwlULLkZeSCu4e4hoUFwnx7VBnCs0/sSAM6UBX8shNl9lVYjvsohfsLz7KsKL/g
tMPn3yyZNORbhwF6McNVdSW9J404GkfkdI/NJYp0VGn2EiJq825Bkx4kgk9SmYo8
Y6Igt5ZtWL+adBhF3aBRx4SocawqonpT8MBk6FE4SNUCCmAse9K+O9KgmJCOLcIR
ZdQq4ToHpwRSKW2d8DVnBVbKyHVLkfpn60dpFNxMkZH+Ww9cWU9Okel2gQuK4bvc
ueV0QgSSPpBTN2WvC7WpeXmBsJ4LWVKj7ePQx7KNxrE7PLdOwO95eToWfhyw6Lv6
OWDoQ/+tUO6MB+KkBypZLj4AY26e1VHH8uutoQm5ewmoq2ovkvgXAF5Or7nmQ15Y
VbNvsPlN9knFFEuN8gEtW4W+xWK1vhM6sRqIiTfkQJ5mzmfNp9hW5jxTlgmrftgd
eGrklQO1pbcU/QHsVYrkpuLSs1R2j15drcOtrO0lOeLhYZn+iu6OD1eCthp9mfay
/eUizgDPjuy/fD4q2Y9/lT/HdtM2ZkflwjfQiLGR40IKlRwwT9ILAV50XpNXM3s4
PeiMAZFsReSr6jBhym3BnVD6gWxwU3vz7bIIfUW3MSeIa1h4r4qXBkseuqFK0VZ+
GQGCtX4IUpq/VE9v3nwsq+Wa45bU+Uwz8rfvvdCaqs0qCwfP0DzG9EhW/PoBtxTJ
Vskm9VefcUhZ3MJsLjow6Mt1KN9Jlibj/lByQBs7REY4IbJT+abfmW8bMyygrTVQ
7GVWYm33QllzW+pLVE0ijF3k4G4X+1uJb54WJFPCkZw9fNkhG5T54XRxW4t8fX6y
VD5eE+JxUn0M6h25mInjmEiP9FvmlYvIhlQaYdfuDoKLGNq1ozDiNRrCZ+dzsHUe
cCssWklpn2OYLy248HQ1kiXNjo3n/OPx+Rzel6SJq1C736cW/7Lw3Z+SIdgaWuDG
3pt7Nms5UjapZNjNz8nh47Tlpmby1O04AWnx5RxShyuOwiHSY+6oiPDMuGuoA+8d
bfROdC1Qf38hZijdkeeMlIuTWxLO9Lm2ZatDzdt8vwFoQFsmH2/2sFJE8yfu+t07
SpgUxC/cPDQirjh9F3XWta0BW6C0JC+nsLwf8KK2X1p8aPv+GHbPx/Z5J6hK7udd
xxKdrzDJcFF8ikdVVpy7uhObIgA/FqulWRYEpzOdlM5Js50oMIhCoafm3sJsCSsK
9MrxepC40pwY+22sdyIaV/XapnZQhGH9tennwBoIQrtGE1X6G+TTYuxFonwSyNxh
lDYsoWKL91l4cTNqVINLRGSPCeaKbKVQGSZF0p0UrNtpN0dYarBXrpgUum/r4iqM
LwM/fozVV/6/wof4+/Pl+HwGmqo+OWSCLZqhtzvIqGFKIF4S/0G2BpuoHUEr2tC8
9o6owKsB/qyF0JuDy8+bGezSHaI6iAoHwYsIOTXAgjOkxijSM/xEUhLbUr5XERI7
rqeSR2ock4pcrAKswtsvnqcVX1nz52eFdeveehmtJ5AeOOPRpFU9/8Og76CblGOW
+0YXHSYf6K2l07hrx62PVcmIj8wVBisolVVA5FFzk4cl4Mf6DtpZ5+BcqgElEpZW
YIbo/qeAgKffgA33vCD0zCAQoKLiuXQqM+aWzCE74M/YQmSvEPC4w/4TtSEFVZ0I
4erzqLvbJq6RPb6VVYLgIn0JpovpZXt+3EdJnCdOu669aBkYyR6aoNlsh3jTWgYf
sAcmlsKD5NTyZVydu7wwQc2fpP5dVGEuKbf8XifcjdUX1JpxIE37cxq+fWIJUiht
G33HelwaP7DKk3KX9tnNh42HkoyJGywgrdo45oUczIgZ+2AWwKQohRQqbPPktFYe
k8LzHx/l0MbIlTs700abwwiHYZo4aFWffPe5owW7wauL0cap+arDmbdw6OKd/yhn
NimKz0tUkukjxiMIo9Ong9uj7u7C/XFsyMwVqb/ktkVTvw0p7956EbN6AaBseumS
fBx3dncyvvUVzP2VW0P7qn6j6kbElokcpAAYr/hpmg7uR5O4q79YS8ecjWAnc7Ei
/MRnudPwJ7eBWOOdrExQJpdnY5EyBfX/gNyd4YrEHGQq32GfRXX//w5NYMRjRK7A
DqjF0EQ3rD5zd+Nlq1nQqB+7dbXvWog61D0WNEsYfTAxk16wWXVmPIgsLCxetsPz
pZMgzzARhS5WgNXnvVFc/+KMwDgORO9qAzCoAez0UNgHAIQC3zP2nKYrrUq+3OoL
Yw+h1dmYjdgmurxdP4AYWA6/stlQVam7sOgtswSqhY7BqezSe49IRsZnuWePDvGG
iYe46OEf6GQtfX8nEH1asEBsp/+d3QKnTMsxMQeVbWN5IDHxOr0SdtNEaTusSZRB
mXXBuGexsFo3UnrPB9/uOZT+gwLvDuJcIvQBZz+d5R6RYOwvX2mPPeFtT1kVGxGt
CXadwjxsGLgg8mo2Q4mhkW2RI8O25/3+jMgCQrJ3m9IAZTZ9hiozPnnsDUrmA0rH
xRPDEsk2iWa/oj1duIpAGFJemXuCV5z5JC4xnRpa+5bxnr9wsX40vgw0p8Axqbix
TrkuzXyJ44Q/vgznF0NiZ7fq1yArgGD2jszWHDMlOkPkvXheMmlSFz8gMgI7y6pE
iWsatLX7y9YJhbRhidhTs0HnfpfcG2ks3VER8NLMbysJvJPJKfB8jgSikvJrMIeO
VHnyQFG5Hd38hrhpZ3GtQeaLwihHNM3YUG4xBH2lA2ET4D6pxiwrNZpHMDkqK7nK
zIO+X24zUQDs1Yd1eF/2olhD7v29p3VEyl4e+JdOl3OsRJKeJ5Kh2RxiuaGH5RlO
gBE/flH6JF7BRY94UhRF1jLKCb2fCR9sbnffpjlDOErYAHpN2usNyDMPDvcEncQ9
xk33yiH9z9+Ki7UYkEkfB+nKOQRVOHw2rtBy4J942eOvSfLdJLaBw/BrbS9ne1lx
+LsjPA3FB6ycDlx79aF3weX7q3/7FujdmQhBla6aNqqzWYJGfZY9flbnCsiKdlj7
y/CPLn2VJF4Cl/lf8Z0J3nhIJcC0ZSwemCfEdAnGgKEWwmU8WXrbDwXDICNPy5xQ
Ayqr0lMG5zU6ajWndagz3jhsc/MXwIDCPCZIeBDz/aU0XkxXLcSaXTLXmX1+1uF4
dPy6NV/wWGxm12rtccYTFu7T7Tn1QNZJQ4j9ixDzIZAztUl8LDxsADvCzHOXWjPo
7W2GwvdxB1SVhk9Ce3mbIBq0kP+gRtUufpvZK9xAOTz5/UCKPbyeYLAkdWJtn213
aGlPqWuMkdfnGcPC7lbo1tutLPdujDW8xxPBD+l10jVTLn/UVCYjvmtcwkVBpuvU
VOKuwu4Qi1jgje5MIo5RxkDrKjGXXuEVzBz+cwReF6QwNdvgzHiff8Ern8EZNkKh
Jk2Va08jRtbdAwpGwj0u6hEoybAMFotoFEcKJHlhNXFGWgyzQ8Ez6jrZDmRmmB4h
ud7b344dlfXOAZnZ1c9E/fwH86ym8idMo9rrXNIOlt9ILGZTjkkwftpHNFIbN/eA
LKHdcxgc5hACebBU/8DbyiIxLBVZW0RKrA94EkOu3LN/JjHOxcIG5FUhd1cSwJaM
wiL5bm9UhqjXm9gxvmeeigfgGOrIlB7jUls69awN2+iw8sboifBgGPxnKXXhZAM5
YtFWuEWDXZZBqwfEKeTdRNkJkSVhI/6n0Mir1USyC4R0goVq4/6XTobo5v87F46d
1WPxvVtO5PZ64SnKZE4YdwyPrhHWAuSXNwe6By2URGx0hVcWjg0DqfqDQGOIgQFm
J4ujD2JvBS7w2UkMZQgZ28zynLCn68alFDjznt1Ig71ru9WzummzmAgr52UlakbP
PYLuE7zZOr7LZ4LJB8khdxRNel8jeg4MhJwMojLXTfUMLoExRf40uNtQEgnWVGuQ
ESD07I6V22ZrJLFHRCKvZ6YNeYblk/6MAy37mMe4efGFYMMv1mCoMiC0hS1Y1w7b
/h2/oNtdzok+JaMpJID1bCnRff3hSXAr7vDCxw5quQKKDkotnKoJCahz3w1Yodai
wiGa3wzVqx9smqgOCxsSb17uHoj7bjXbrmJE4F7OE18wrKELgUouSV1Ge7it0mWx
tfg8+wnsQ3lmMgl6gxlJkHvnY9TFfNo52FUrFkFgF9CP6k65Hy/rf/XxErabkRCS
GgDTghwGkitZ0rTFtBNsjE3R0cp6nuQhtN+SwXRlYblv+3gpUv6Kcy2/tXLUPw3Q
7XbF0y2oR5wKBAmGKAqURXg0kCGZsPGpgfLKp8eM+VTvyk1BEZ7+04ILdMj+/a0J
722hLAc2FYp9i+vj/V+ZpOO8fQ3kgC2ZHz/74vRDAg6oEN2wpEBlbEdt37HRRab8
auQUMRACs+VaILEcWid6tgVXMbhLBZMZw9P3l3nY/s++njX6dJ29zMf29tHoT7/E
a88uBBwNPdMUxBueDabz2cbkc6BjaEkIEhYINwjbzaMa0eb2aEpuazVd7xdew/pq
1LEig5gZ8MoXuo/v+XpNzpBnkgDDqZ91OCgfuddR1c2IDac3RAqb3MRd/0ZFOkik
P5XBe5YME2qOjaG0pPnLZ7LVxtXdwoOPJJQ8UjFu5nU9BS/SyWdZlVAqcsAqbKVy
nh7Bq1tX9DYH1DdcqEGQAH3eWNaXKvZ0drvfUwM4fm0EPhqaahTzb4lw0Fa8lEwr
Ll6GQ9QB3MRtowmf+9XcHP4qsXYWYjby7i7GWInx689DxOy9cb33rEbNWspz2pNe
z9WrE4pZPZWMbDfbxn6ffBQa8xKOtSncBXFLoUXXdQjjMt5y6cjt7pNrJ3RT87tL
qngIrptUy2medjQxRzbc8PpZNgaZVLSvy/+GTRZ1QXt2sQZlCA05zMhsl9KTJNOQ
+InDFc94nXpS9W4N6w/A6yiJN9WI2xXv8T0gJPzlRSyQqGbS0BNbt+0pc9ng2oU0
1qtBqBVLnn4ax0e/9SdiloOKXdadXpe/75/eJlVPSNvKnhafSWUpqW9lGA5caFdO
LjbwpasM6nqosCbAhKI6z4qhl0mH7Rc7wwMxE8a+yYuUy/EFX28AiRHgdI1I9YId
6bVIkR/I1olC5SAIQm4lzVs354Kjkw5o67l4C3OoIaj5Z6EF1GCvYtIZzCpPYiLi
PbR794Af6Um/29DpSQKTcZLIGHlL4GVq/Z2nIgO8by8DQvK7oIn2zFsPAYgS05H5
Li3vOVOhxIVNvTOVyJuBxikDYLQ3L0qSSGbW+b5TDIadT5HApUjEp9l4HgHxUDun
7yXL8X9G6Fz30aA/unfPgBrSSzMQUUwtNOcLIwq8e19K7S/HN6y1LCC+xtP4RWZx
gJeQR48l/wJYBKumaiwObztFzYP5y0JpnopvdqvWqpgw9IuFEbd1xPVhGMENKUGv
KrmeJfYE6m62bfaHYrVFnfBeyXmftPfEnnU4YyCUwqhwK1EFTU4YL1pFyyEM2YdG
PYEiql72URkwLCqqb/kVUofdAvIZxCKGheNJ8DgbaD7uNe/5wQxQlJ7pHHIsHmj2
YhkgE0djcVo33kd9zLllGsi2W91i+z7icowv9kQWcdkXvDSBvDIdoVYLonzoz1PC
2nCFRrVKC+5tUaVkUAIIjjA2gE7UG70uzXxYBxaVT2VwZD3yQI0ROD2ksnuLgvs7
dcMw2aAFuQdu9l8XMaLHXgPJxV1MfFN27T3viUYCg16zxlbiW7zk9dvTQr3WTZuH
/xnfkQ+LcV/iGju01EvW5n/T17/Zl4bjoq9b6r8lUMXdHpmGllQFsUjvojE+VPc8
y4LRjfHPvqjH+62SH9i/n3tHcCRJo4B2yRTDisyTGzRknQusv5yIBwbuPeGwsvmO
NvYFfKlAY++Z1CsoAx14EI6Vs5jnTAkj7jDJkCs24L1uos+mOg0d8KV7wDQ7VlDE
AUJF6whzhdOHPStaUH0BsqZAE8HhSf8EFRwUSzfAo1RjQ1UMD7XEdX7dSl8vZTDZ
jYTLezcnM0+dzG7o1udSK3SBnY6cLKshES8+aM0qN2cb2IKSyge1nHWzyzJIX1pw
zw+L/VMl06ihzxOIJOOU0Rws33YTLi0xpO08SEKDf5KKSvzfSJHIg0IsbRKv9zaE
v8p1kfQFOhj4/HCFwNUDhjaJlfPPaZsrAyyT0JEvwV3U62o5SYVkne2w3p4brBpG
94S2/4Vfzj+2xGsmbksdgcV/idliJ5MudAQiWJWB68sOAy5qqPlgOk5gypVSaMBN
a3tXMkgHuM0fxziDScUBoKPoNOwusEoNM+eSjSq0rLrEC4qszPQjO+Umpbe7C+BJ
xUBJF6cNTqL5waHlZqgXj+AR+yz9+AmLoiqMPMsF4s59IITDJM1MXKVWU4ABuU1g
Ibd+m9aPexqqXHRk5xCTg1K0jgxRD/alezMk9ZoY1/EIb/fRt9iRrmAK99CH4Cw0
hO92Bx53alShbcIOc3tMCwq1Vu9czLMyUEHyngdUmJCIAfbIbDdKPsioD8qMKt35
xI5Dwh8MFpjS+yvyfRj/SE/FPEe93bTsZIAGdU8o2GJRacBDU/wDeqWaB7IVbil6
PR1x8E9WcsE+qRlPF+QmpGHMnsgNneK73BHNAX0gYR7863ijXv3E8exEAxV4x9yR
ZmMoBPBouTlygGjfs+iY7lTeoG2io7Ntb1Uq++fzACwIyCuRZbmkh8bgYfXubLaA
Jpog1IDwr6b0C0gAeifFP5vh94V5M9M4AGI2Cv9wQ5c/bKkUR9UgjBt0uYbwW+Ly
D6sP5obv1Z/r/J3LvoXBm0SmVoZtxDEK0NEyfQLBdczPgesH6VFtb8oY46GuCj4c
qm/6q5KwIzFBasY1/s/AnV79pzymznohryoKw/SRdv9VyG6bYS4g/2z0oIe7I4Jn
Rd7VXyS7H9ExYuerZT2XvE/nyU6RYdogt+Dou4SaahRMQ+C9uFjCWR2ZowPWmUX+
xsQBtK4hX7hYyb80xKIekdvqHbxDtLaymveTtBMMqf5PvU+MMVoIfui+DPXBEIF0
YYAjtRQ8ahcdxB6uCEsq0UNNoaKCOK10R4GXP9+9VGdTVv0j8iSFUXxZgxnnta1l
VbxdfcGVg/sM1HwKG/t3pe0xMA2m99d3HiyP8YuIUmu0UFaY1OMmX8gaFYFhpiJo
IOfLZSNCQOWakSNmCb9Vupz82755bbgUqaz6AeeW5cOOuE455LBE6KnNaNlYtwG+
qgkXGtPAZo/8z0Var4tFeNUoDAHHl+/w9sx2geH0kj2SCkABXRfSDIhY3SKWkSyn
u2QufD2Gw5Su925YxpP2L89JdSzyGp7ltAtstq5ZJ2NIbfTGzdFiVUjmWj4rnEP1
HQcVYJdr5BbfGpT9JDg6LDwtWoRwRltPv/QqET+PNrRD63BoNDiPNEv8RO0qPpu6
71a+nINZhShJ6GEj8zKYk/UYt+dQ+aFEpCZnP/M4JsiIS2F+uT5xk3oz19d3t2mZ
3IQ9xwSpQ4EFMnoR5VV1V2LYRba0MtFw7IbI9VjDStCdUhmse7gadcXQf5agQ3Gd
FC+LFVJTV13QOTzNoLOiP4TpemdzHGa/1sLtxBJR0E9XqMog25zI32vh5YKNyXyK
0pMG7E3NPYEdgb3DzY69I+02Rkdww4STzDKeuGc0EiMWBJDg2jbKUKkY+wxmTnyQ
MuymdK6w9/yYG1Q3Xim2IfVFzR+O2Hp+Ex7DEo+61vonHc40l4PUHNPDrVLFTUeI
un17n3inZX7gNVF7XhZNZR0L/ih9bvR8ubcWasfGXYd6BJb5UgrX3LtPCQUGjOFh
dMbXwbFlvzlc134xDYFL06LJuAzZN9Pom3eQZkFFkBPQ6mjedJ2Xq1a1fAomRjdP
Exl2XXojczBZSUXsBiDbm4zJv8Zp+5BteOBTHudUZ+KMgiuuTvY4XQ+zrvF45rq2
G2/Dqf94o4NhCsIQulRYoqt75F52BPu1+BdRtCdfrWebehwFU4CQn08GJhAAfAsH
jWsu6RYDsOUrL4RAOKXcPgcMwGfgaFCnAN2pv9Xs0eurhtQAXWMySCzIfKPrMv/M
mF6DfVSu6rpAFmpox8mxGXHAM5GwGsDnpwhqLHowliq4itl6bDQydHh1y354eUjO
emCpDhVbsemxh6nO1iXTrqBkzYo0DUOhs0eLRN1amMOYIsfSBxU9xYquXxvekqnP
Cax+CzDTnJ6ucXgW4jLidaAhSlEwa6bodkt/Mv/oMhV/KNn/1JOiGHHmz3+eJowP
NqDx2rK1U0sFU9xuDchdym4AdjHJmXym7Y3dimVPINsXNfwmFb8jRN92fI7cddsS
Slx9gg74SLao5UsgHFOWTL6xAp8Whi8KgPJvgHhe55pBMVODaEFzbaRNabS4R0VT
Kg2uamALSJoRSJRVu1C9vso3V0ABCFigFYXpBmXzowj2EmtFwDVfRPKHvjIlivu1
547y1ela0jn0yIoy9LE9vuQO3lBUkie4WuYoh0y/k8EFzNlSJbYQJzD1JnbqrboX
H9SZRfq9EfSoG1mGygz+9+kT3XzrA8OGAXD/im7VL4NMu4ltMmZO+4H3PIAqdapp
WTcT224fNpg6BTagpLlyaaEMWuNhQiOqqGaYIGT2bbQtcO1Xwtp0xn1tMq8EWRI4
bXueqgobLVi+z9G8xE+PQmlDq/OzIy5h5YevCuRZl6FibU9ZHgvT+XW3KsVYR1Po
AyGVZSxrwlHKtX3O6RPtU9XsftopcDBNtiVFynGrnL1EiGasgLzIit9ocYKtm8n3
QFKitubZoDfO7DzcnDYTbfn1FTcxuLfC2UM+QEGCBggzWAY4RyHtAZ0gjP7IiKsa
yxjs2aCFMpbSX2b302Uonnzzo28+gnDwuSFh9sFHqbs8uCZY7Q2qde52PzVnWdAq
HL7VtCal010hcry0JzcGAXWQJvkL7FR5fbJOWGWKB312nY9WGr3dgnp6IUaGKy3+
mRnOhuVKQMtoD8csX5sNnwSOpI37+dTN9N84eLe/MEPVE66wwhxnWQN4WdN/Bucz
waXlaeoFNf5l27rpOf3nSBxMfi4mGNzxr+TdODxt7pWwBjcF8+llC8RfdcFNKKvu
QJnAlUhop3FTgAf/6cOanmMwCxnKgEEFG6p4sY0LcANChxNql+2I5DxqBfJul1ze
0AxGvR8USPEiZSs+I7OvRXN9IVrVht6//+qWScOx1YMZH74YHLmWYRVN8B3JAOxS
08MztoWGAVW75ozL2SpMJcbytMMwWTECd7NP4ICIGeZlrayxhUJo2VPDStdRWuig
nCorOAeImJ5MuXGQmvp2ZkGuN11GzUhgL1UUakwuiKGfd9R1vuyJGaxG+CqDGzf9
AF3cbLdu28CyuaLvKQTtZOTsRvoJ5ZrA4JmEuw8o7p5HTP7kpQ6aAo2egb/fnRFk
L6fd4YPM7koWhKSVAxZm3D5aVVKMcG1QVMl4o/j8CAx8YxyoyEU/DxLcL3E07TIM
zS3qod9+wffly8PtL93qAAdzQ93AU+1LewyDsQW5p6piJB80c9cRaKTxLiluxHa3
mRR8L9sWqQtnG1b6gkuzBHaFfamGrXtLns2dP9mehRMglS6KlkCx/DgZ+/7lXFCN
wE77jmlraagkpLlWcPXAOYgN2/8j+ho4VW8a16ATvjK6wpwtSKMU+vL1DJpXVOmH
7Jg3hlND1lbJJ0xHj8cxez+S4ou9gBkMhGXxmj+kjUG2p3+hY2LQgScxvxqs0m9t
SF5bn7fcgvMN4A5BnBGtSsgMbBUthU0DLoxRunDEdl8MARKenCwH8syMIZ+8DKGC
bqp104EUdLqo72fac52c0ILMm6KiPmVgBu0cujLudba/tq7ZfygJi29jb7L98jja
rRywaH76Iq/kGijral/2bW4dQcyYPoAloSPh7tAHXfa6/fU7dvgZ0IwOXc8E3hAP
wOjTZtxWnzfHP4Iba4B4GNfNktSBgl22v4YOdC7fcIgZ+1Y7f8wEpLcLNHQmTBjG
ztt+hGwgtsdZDFA3odHmpfRpZIPA+IQ5pthUItJURiMkYDTZMFn5G2R+FC9AYgQZ
Omm+31Y3j18y5PCHh0TRvzgWHAT0+cSZjwQmqUZmxnTsI4xuhNInf90g6qKGEc4f
SnJ3RCSLMCMYarJlhRo50c7ZUqrbDnCP4lyikUpJZ6xMJsZl3opXbZArbIjIanef
+ql4J0LCRFTpO45goiqPMZoXTD/i0x4TJW9iLphyYZoAV/wN2hi6zVskcorqS/iX
6ThluHzHOTE2A10eEf8M6qsBPzO8BuuoB8G63Rqti+Q2RQ4rkJJY4STboTfXEXWx
SaEAN1YccZlJnXyo0rXAC0ImuXCprtBPDt9NicCDhjZbE5nwi1JBRSe3QkdL9ffl
To9PJvY4s4fTbKRI3o/lDhLMTGCBNNDgv+upo9E5EEOcg3IdsY5nqi0VbaDe+t16
ww9Jz26al6wgGUyBpX1PqEk6E8C2WBhsDFjLzrTLkNlvFMD0PppngBp8p1IMhFOe
mTgP7iNFtba22bUHoVwyfpd3h5Hm/icK/iqC4tST+E+GRep7KTng6FxrUcZE9flY
wjuYbNQQ8UDErmTUcu34Ld5uS3g8tmMaeBDLUetZNDBZwH/lv7rmx9yezrIC8q2E
rdZYyd6/V2A2B6LHsQlOBph7HAf+jxzYWZwcTeeai7NiP/48b3eaYkJTg0a3EOMv
/42iMGjVgBP6UXFu5FvLcZgx89jvUfOV2AAW26QolAnqbVfW1/9SUzILC9OlEvY5
bPo/MMdME/Wp+amsX2+wVk0jWEf6Pc2iTk/PmQmoy7z8XYa2aZo8dNDEjisMRtwS
Erpx0AinpN710hcnMwJP2A0Krhd//A6lLUUJfCI0O0oJNUKVeIlIrjZnreW0N1aX
s55SKlsUXWn7nSOAIEJfm5NqC31YXEwQSrisynV5iTqdJ8BX3RXwltQC6/V0v3dQ
2Ant9Ty+wnBcqZ3u1imURW7uyqouOgtWcvFrAk+h2oOJ1JzR3vj2ugmti6ZAhn6l
FtjgXbVU2CFM5MoZBaYChTZwZW0jFFOzrXWZvI8UjnHMbOczm+qWRDIFcb6xuAPF
8B3tXuW1h8uUNB2m6fdnsBU7gxji/ABMkiQMOgiIN98DMBzTUCgo96jyCCWCTb8y
1mK+Py3AUBM51zlne8P16QF1PVqLxt839kND9CEBQfEnoEcdWhRwn0SaWQ9h/xmD
qWC8dHfIYsXr/vBkUhL9MqQWVQ+bJ+Gx3EkO/XUXxcDWyxhEgj0PrP1IGH3bFJxj
6GgjRfaDUTn3g5pIrPBBaSfolZUBjNeYRItMd3Pzc6ddZgs6+pmqK/mf6omXonOa
MH/NeXlwIUK0eZq0XnNtD2vrybiyNU80Fo+S9S6cv/BvG5lj67yfWticmXeUym3X
2h6kYR5UtoPEfoF3oHi7dz2J1PHLyTK7WNzgMWBIsmLJS5ktrpqZELAYlSOa4QJb
9+Fl8SDa48c7BQs5rqiSpgztc6C9NvuaT79ZQZOmb+gZqlRvbMWepiE7tTgeaRxz
QFrj10ZZrfbT9MkjmWyyYvRDYWY/CbGCuKF4T/YX8j+OLfTTTtnfKASPGYDGhltZ
EWD1TSuSjGr6ALftBnFtAZWcWQ1mE/h2DJxB3sJEt9TdMSovTE6zvjsgxGezCQS5
eRVtygo1yME8Mj4Njehoq0bWIdtUMyHmPhBXf2NNY87CuEfWrtlziRAJ14M7cvMa
DwAuxC9tAFRB9u5C7wiacUH0rg3JOcXTuY9djI7g3VfTccx9qmONSD5vUY9i0ulh
o1cSrrp3pspm6ZvbfEsdDi3SxwYa1LWHDRmO9Hivaf91WwyNjU1ClfBfm0+aRMdx
IrP0z6igOM1eharKSQNPcwEyJFLqgcI/THCoXyWMUUGC5UDTw9IUKe1LpCn8yq5K
wecYwR+WxKCqwMxNbCazPSrJLPEzuK5/1Atc1L8Pksuab97/jb2tzS4ESmuMdIfi
wwo9s22zapq1TWaTM+6FH3VGcNp85rapfMc/fkyUvbxx1syy1wMyS7h+VpiofKR7
r/OYJnMWvOO/RE9yLGa8lIgeeM4VXXj7R7XxiNAW5CWTuDxmL4SjEOtmw656OYI5
laecLAewjVfng7HttfDQX4iJMlAhtKQFsqqMT2fRXpc+ex5qVxilp/+t7tjGpAFQ
tzm8FghaON81D8lClrAuyFh1jLg4N7JtMdqaGDwzVxYiliDZUSWtsG554ri6FrQP
CUF5wDHE15jUhvGfJlUoBTfhBlcQ9FzfdMDgJ0JT8MtgPfxGWmLHvtHeIss4o9io
M2qY2u4OKEUAaMsUkOezFVNyL4d/SJROyMKCq0N2r9HaCqwob+dqroRKXkctHpwU
gLAWi1fGIQyU6KyiV7b1fC/UxExSfRNT+f3qRIXDW4NxSfaxPG5hTjwe313KWkyE
m/MzvmyBBKj7JCESp4yjgYO5ImTWmJgkvq94KSQSWY4Alj+PT1CirYL0fg9fx3Cc
sB2n2zj0/DMdJy0IDf2M2b3bfIu9GgepscpkfmC0LsOxlGYorWynkOVFi1S8wjDE
p6O2I5Ax5fi2YhwVkISv81PbZ1v/II6Yr39F3toOGZPZwrT6YNReikICm0M9mD1G
RTP2rfQmq8pjWFeevjbOd2rVV18+d73Ba2Ox3f/M7irBxqLXF183bo5r1HwvhiT3
Gj57OYj/ajNTW6ZdJTvOYLukDq6B+1DaFXFn3DzDOvuFuynIg3rH9P2LQD5Ef7Fr
vJNVYDl88ZaEm57S/zZUZRvq8TZVUuCJsHJbDi7kyydFgYgGWK3mdXmXtRVdw558
tki+3O3uSQfgEiB9acWRB3uvSnymVgHFz0QTpfvYU2cpJge9fCsTeVrZCKGaBxVo
zY0khWpMXLsdHeiqW5sc1/MRuSK4gLpC/MWMCfiI16dbLSW+Qt9rSC4Nns7TiaYz
qrx0mTnWdg3qYP0g1jDulNKyqL8Ni7b27EsTJTD6gurG1edxkzwhk91HqCs/n8Jq
y5uDng1cuFIA8Qh+w8+JhmX78eMp+gafJGFazQRFI+4IyfrG/b71rfRlL96eNK1O
CHyTk8bL1/6YaXWtU14+jb6oC66m/3DvOhLvB9guDZsq3RWNLoPPWkXLOrM0jXFD
4VoQfv7zIZfFG8FDGQ04LrfL7+9e1JhZygyQAx4bFS/0f/Docs2flvH1WH5RdQw+
RQV/3UJHWw19rjkQlw/guR4qmOFRGezYXPpKSlxoJQa/RPxe4sOFhCHJRoCtLLL3
BmuSXiUQhQ9wuvUNJk2HlD+IHt3+ejL430g4tiy0b07nvwt9mZ/oErk4AxHE+xO3
G82U2YWqjxvz0/WEaDEKYAFg7ws3Z9nJbY2pFP+ydOr+refPCLTkjexL18IwgKll
yzQxhi9TOW7HbOeAGkjYiMQg0GmcR4To8naaBWrraIpDAPKmXqH1Tdz6EdZbEH1S
DIMRX8Sfqpc/HwitmlNNNxCR8jk3w6fnGwZtNi2T4gBPL2QW3mEF6jEzvhFPhy1Y
ctqTmz2JXqpR9DoRAMIzC5kiIvb+QXsxqrsEtsG2IaAFfD8hdk8JDJKRzY2AP9rl
ettkH3BijDUNTSL/zdokOXT5hTkTURnTHYg2uAaKNKiZzyhjXWedyzDfLrrnz4yQ
WNv8m2Ph1DfpHn+UkmsAUnAeexGyr3OS//az/8vSUvJtS7FOSYATUJQj30SVk3IZ
mVWxFfNm9c7JRqWol4JNgI/PbRtQWpof/TXKzBkp6DPE1p7BZYYHodUWqQCglH2W
OSbGF1V3MpEvUAIkLsXAC2zoS4h9sT1urPE2hlTyOjgEc7TTTFhbEySkD0X9dQnA
6t127Rkp9LjuqTicbjIR60jWkKVgHN4QF+e0zHdejOKRAv4QxNKJ8cHXSu4YgIR7
6WCbR1h30Hxi3J4B88oYv91hv3T71I6cpeoZFnmQBp5Y8raUjDPUebWGQWDZDL9a
ups7JOiX71sWzkvNnmkEaycX0SMXguJaaPfNh0G4uW4/9SkjFQR/4YkUs85n7gJg
6frfe+4P1He1x1DiAQDxgym7X6rlK+JvbqQAeeEa9Ri3d/WvpxLrQjqO49X/oeG1
Eq9NKxoH8JwULxL4eLK8E0hSfkyXDqaa2iycScCoMqvPRV47HsIZipcRAnPw+bgV
FAorarsYxrrIIAvLwsQXadDQzvm5NDLJQWGFPgYvrP6MMooxXsfL3BoZrW8BKYWq
BduuZ0eAPf8+tWVOoGhp4/2Blmn5wDodlXVFj51f23LgV/eX97hXPnlSltjfYhX4
rsNmS04/sBeTeFIthjuCLVRttOKQkEfTH9NX5YI8DDrHINMO6z8pqsfxPLrlLdXk
2zXx49NNpWz3T5uhw6OFhuC2PLRHxYY75xVgEmC6RF+dmMMB2NePjASAI0aJ8JzZ
N4ZirU+PFOJFz4KKLPbtRBcF71e0Zx+8PlpO/R5ktWvrRrqz5UUvWCxRmC4vmbYZ
VAavKs46Fhl4UVuXUuuDbMuU52gIKSOQTSK4KjZFDZXVInWmmD//FwP7yFlRY4Rj
q+3OyOU6Bd/R4ppmvWyEQ5tN7tuwo8ihxcqHk0RhHiW3uozcddC/qQaizyLfAaLT
QZh6yRAFD/W6o1fcznhhOGQYrZLixrb7HvGsj5jw5lI1Yr1NCevSAitBYWvoPnTU
UD17x99gy877PEx+9WnMIl3isbnCNMheEvCmCrocGd4T4KzgiDCm8mWrnUeiteUk
hV+eDSq3FAIOBOvYxQt+BHEUoT3TlyEvdKOhM0V+Jmm6M9AI0pK1Bi+k+z6yFbWK
o0FHxpC2s5QDan6pM5qg68I5O56RIvlWs7F4DDATAUeVxTbOu8t9CaBIVhhW5PAw
3ZxZPD9ATW5wB0zmlIF8LmUndOCQySsrdUr7W7M1Hpk1ka4qOhiGjbJT0IPm5n+Z
T76RCys/I8EiwGDsgnjjAd/OiMcQBgyKIIFf4Q7ldgqOdaRBP/09IXTzKEuaFBxt
MXq59KSFecnXn11Sb/wJsLtPGIEyuz60Z3Zx7yfumY9ZYX2fKC2LTynsiLhC4Ddm
FabHLcoihacQsBJMfj9Q7IP4NWABqkMmZLMqucl/kEngWC22knflSZAcZIK1p0wT
QoXHeLdm4MxN+9yv1RKOXC9kV8WR7/LsAZFjj3L8yN/bEExThnOnEaU0aUgO3v7D
Hu5dnxonUo7zxz5IEV9gNHmzaJApn6lZQ644qEzCSb+RKvnyrMMh7yWu3W1dkH2g
rU0YI3LMOYbXiW2jaVC3tMkbjwYBoEiOu6NN8zSv37p+/qa4vEmKO3eoV5lXoKS6
0mPJ4+uzt71O9mREuQw3LBTnbeSZssZMhSzEq/mWDxwmYpiSR4bles7EcQbAVea3
HsPFoijZopGFyq/pOT8QNBJarLT/nwZLLWo41hSUD03jiqPKK4fHd0r4A6DvSsvL
A32AHTG/on3gio/+7GsvT2AeR902glQInUg65BUyLxP7U5eqcri107e61CbijswA
RzT/OhJbFjeerm/Qtj4Nis1ZtttrCrn9iIN9cmcc3B3RidhJ0MypRnNnKjuEFunt
JzCFMq8dBau5IOp31o+RUYCoDjZRVHEQ7CCqsN0uGO/0yrKthGk1N87PNCdBQ15b
gZ6bdICI38w7WQMX2p0ApWDTYSrNrhldUGqlts8K2wOBhZHoUb+SYjrsVq1wnft/
HUtqmuw9NuRsa/+Ov6orC2s4Bo7/JRhPxxJEf2egZT1NuhPl5Hpcn6htQDDsf2Ky
9yg11EzRCyYd+hIF3CnTqPTSH745jyR2y+WDfJsG0gJxFnpSFaeEFFPAEhhTlvOg
K/biYQMe0U/iEBX2GJAyQuBPNFQPaV54hIRkOS5B2bvS8dUsJRUJsNf+L3ZhZtfX
KCMxJJ3E5E2M140NBmGpFnGhDP0bII5GrLdxUp7FD8gW111rIKQKQ4lLO2qA3wOP
AYZF7xPOQuI+eA21tg9cK3EnNC6WltuRataox6Xha5xz6s4+gy2bjn1NhfMKH7PY
I1Tzedytgzm6VoruEVIu36yU7WQ0/YDq1J1HIyX4ff138bnF1+Gc0u0KxC2c7wMN
Ggh+TcLalTJ4pBeNJNla3kstq9KJtI56vGA/zSumADXLm7SGWQlHF1gdGdvSV5pq
WEyJUlyIxGAxpoHyLJhF7rwIcSMWq/2+vrj+uLTgVTeNeEvTfjUklpf0wpAtZO8M
4elNTTf1PoLQqI09IGyBviD9Q5H7QiKyaORTHq0NYPXMkozv6AZBVs1jWxH8iX2G
krlxhs4ACJMah5MBU5io6iSRzvMMxkWpy1AL+2tB19iDPkPiXJzgERMSZOeP3gLq
Jntl2devn2iBiHTo1H+pXpGxauwGTCJHzWRMMRYVL+bCZa+C9pNbTptYdba0vAKq
F7E6y21CBhzH7kmFCfXyeT1vDZBtR6XIhA9cKeQDI5RO6HyuefOoEDu3DlcLdL3Q
/y4rA/4g9vH3lFxxJ5MQil2JlS9QcqxljVwiE1AJLpUwlVnl0tRgZw35mOq9BSvD
h9oS7zccZCLhYSt18dBcmEdb/8ZAzSIIkHXGBR4qTMkmOZHgsmll5o5ffePSULky
VZ5do/QW1KDvimhjvGP1k7Yy5c7Cqv8kV6fK8XNPaOghVBVFyULywKXE+t4fK7MQ
MG+F9pPP46DCnQl4GpuHBYBxE77/+5TTPDcKwRKa+Wc+eXnZ28SmCl50jMcf5+gO
6E74as5x8WiqZ7I2U1FsP2OGrv9zq2WbvAByb59A7nm6/9a1RWZsqrmJbRHJu8kE
p8qcO+/jy9xOR7nyQp8y6uCPC1pff96FFQ4lBH55jVChdc+7DljTQTy5hO9q5rlF
WMZAI+EczW6vQOx3UlO4sZOlcpvpf1cTS6c3gJeGG78Ox6FbLQ/fxBVCvrwsvd3y
VPxjrKxyczuZj/SClHKnY5gJWmW0mBEDt/mPxFpiNcurEX46rigyRIbl+fD8AA9N
Rc89wtosvx0TEwK+pu8jXSvN3gsQ4ofmDZDYD9fbdEc7VoaR/zl51+4XY9891nWW
2zR+UA30R66pDidG0FYGGxkDJNjJ6mL4wPLiH4Tn1dx+H5nddE1Ellip6PC4pEFv
IZ7cwZ0XDcxcXngq2OT43Vk6tF58h8NNyREbVJMDQkGce5ntIaFcrYH9efbOSrDj
SYGAJurahYYLUhxYStDsRbxHkKgmq/Vyi3gyVtC+lBOkCzmkrIOpQxfIwTXB3Dnj
UJgQZu6MngfttUtTe13f/ahRFnWcLi8emzKMQJdVY6p2ey3LAUXCefVpD8oiIffr
fqRx+XrsLgIS1wj7itxBaAoQ2OV8/viih/bJviRjoHGlQtdLHshVLUO9pfckqDPO
78RodG6kABexu/54Z7P71eRJ6DXAMS0H4R/izrZdO9JXslxWHHFCegbSk+cUlQRD
vJbHvAKSE5RBQdCH+YkhwvfGQtKLsT0t79XbluHo/Iz0saDWkjX/+/NLzfZPQash
kSm/xWIxLjUpun0rsrY9GrWMzeiVI7JgTZaL3eyj+h+QI9BQO7S+Ty5SsTHQr7T2
WRjUIvkP5ES+KfL9pJs/nVOHCQT72HAgqO3RbmyDtVGOB25MJQBXBZMIA+/9H5b6
UAADXTv4Mg2vAFXAhbTm7HuR1J2LiTpnX5D8RGuGK2c6lI4g0n1VQc3cm4G0KUI5
2nZ9Asp6YAHrofVJiSMrKZVPyhkPT/sUtRQI6ZKxXrsJCchZghERmCMVSOgogPVb
HyPC72GGFTcJ8IOSCgWIb/xffTXEchK9ONY90sbMT9T6w9Dp1eKLlf/CKJl9Ut0t
pjfmHsrAER+dpWaecD8C4RFY24JF82JEM3yF7kbpeU1ARsprBaY9XRlRDp1Vc5mS
XuM15dNJTmlx1y4iItnlbAHsxjKzCNmPsBrfF+uS7aFWkLvOmlCDBWO5bmMO+URS
NAmBGuXH6qnhTdr+srCUqjh4O66GuZgARS4IzJt0ipXs4EyoCMVn8whFO3j+TmoI
s+TySFhsI5SkaUlY0fK8ijbtKVZG84gscKsnQ9wOTpkvwhf6m34P0pcD2RHfE0W7
yCu2aXRvwFJw1VqFqJsBg/uDccY7wfJwx2ZfPEsSMC1CM162U0mRAXSTKKSRsaQx
3rVjjYbErRXY+x6TEX+2tgSbNXZorCke83iQY0BRzdqpOWFZxJuDj8/+S3ipQ8WY
r3F0MrbnYouFwIb369looxzcLAYJEcEKNhJEFvPneLWkcBjLLX2ZtFn5qOwohkcN
gpf1SLdIzRI0qHJNYjysDfoIGAzZoANSBXWcSkpbGW3aSLTcJUBQBd/zWwfv2g/s
WjqqC+SrRx5v4+SLGIAK2/mod3Aa6AxkjlgoiVdDu1x+YRiXvoG5AP3TqWpf2DNO
tSkq2Pqks1emmP7cSenvGrgkmdFSbiPyktQY6OsGITtE8BOlSKBXeVO0+7ghgTmX
0eh6o65f+/CiOKVM8tfAt2YpfaWTEiqY3MKUf98QqQox3W8mcZZnsqutz8MJldh/
HGdwcmCgjZJmzRvo+vLnLYjfDxWDIF1PVHTPduEctNJOM7/iLH38sLTTnluUQrpp
8wJMmkoBpqiP3hxVtePFPM7YPENPHSzgjdOZz1Yp7aYYphNRPAP353Q4TFTtGkcx
U/h1JXR3c/YDQzM6yAKhgeTV+JFGawL4zlyoAxLPsd/lA6itgc4TwJmM8gXFTQDh
k3YoK8tgihK1D/tZ8frodPiDwtkUGPtrBNbIEbwWZg5U0wFfZPmur1x0Cg6fQWn7
aixoUcsT3nU/ePu7Ptis3gqDFhqK0y2WsKPUZB3vJxXAJ3Pg75OQtjBGA8M2APw4
M0aIK0UcsLSrAtU3HnVUdquRxLM8QniX65YpuvAn7VpghPhWkwcy+CcYXZja8SFa
Mb1uZSnlsG4chtRO5dz7vNVBaIKlkRjg+D1PlWbAqiekwra+qmHH8iem2kTQ+Vg9
Q+8nvfjL6rpij5vQIhm5Ymk51wn5VSlaCF0nes5QDUeRDlJ8V1YR1lZld0hAtg1+
3kADDk/4ZodvTxl+TxXZ+cwGN6A0trTTdkEibNoOIKOQqG7OAcgWw0jgGydLBb4w
nKllo3m3z3Lp+K4Fq9rlao0h6TdQrs3TAG1U7s2bRjqrTMcMPPScL2+/Z9LmMb0h
bjLwdbyaGoTIMnjTCzqxLdgDUAocAY0L8x4hYMtJesax9TXLcSMMzEt2d5k5Hux/
zevhCsTMmAj+b5vydYGz3/veimg1nNlEe+yUnYL0xToZDjUejwTG7DMlZO/Cc86F
5tR1hMf9tl6W2NX0fjWb4bRXNlYYaUw9V1kNCcH1iq5lmHpJRo7Dta7zoSk1nYKd
95fo+k6oqS9PrDWeDyVd1c7LWOGAP9226dMvNM4VzrypKN8H9BaCK59rmwS0fk4S
XcmalWznPKgzRmaJkyvDu8CoDaXQM9BwP4Pdyzq46gPoE74SPP/K+IbkC0vMQ4oK
NBm3/08ORLcO3JJKXwXAWE1VzQ9jFP0VW6FGEN8+WWojlr0VX2hDLyif1V/PFgsr
0TL1/8fWaOOUwylxSsIk+kduee+QjFPwmdOAPvR8dbUK28alltpBu83kGuPONuNA
M8AIN64yxgty0JnUrpMlMr7ZrM2RidgQbq7GH97DZV+uHj4RmAgqZhc+1Q14VPLp
6KVXyUtb2SZVgPBatlTLbeQnff7uOxSVrSehagpuZZIZyvAEw4M2VvS7sUvufxb5
oM3hl1Fuv15pJeunyENDkMqRDmNn7/7LCp3BKZXfrKzJJiRqu5XYAgVreFCJ1yaO
4NOgeWBEqYHph74njAv5ugdMkmtVWJiu1vRxpiGA9wxTr74rSagxVlRq4TATsi9d
jlCRih7KR8n5banhhqQUauEUFZo/6XugF5yBNkNbGLSSMe0+sEe4Lo21xGeN7geo
SRmuwp2YrDf+X7XKYm4qgHgWxpVAsfIV6jecWSHzDMbiMsDSWCd1IzcMPktavFaK
KorGmukm4aQ8/d5nbgCf80BUut6gheOp08gvZKwiNs4h0Wy+BiUNdAhLip3gyrl8
MJkw6QOJm3rDQRe4NppJSdUiU4pceeu/6GnU1DJkz0wpc2RvimNi4abYaHjtOn/1
EjbNDAVrWUmjTD9da/7EkPB15ht1FEQHySmr1pV2VdwEDsy+1Qwo5WHTrPObb06u
8hAEY1C7pqqIO5BfYlJoqwUILFmMpiUswQGr7NEWWfdLrR5Y81Q3uSeO4HXVfcoj
6uOgWYcvqz2zZUExoPGna8WkMyCpGzuIRec/ct833++cM7t83y+kJzo+t+2U/J/R
QmK8JhDBrQOac/o54rf3ZTzFHd8cc/TLrmiGFj9lbvtCKUM6xV2vzK/6E4QxEmm2
YTTdHBvHVslwLYvAvggfZfrkoIU9x5PDlo+5480d0JdEQH/T0dOKRCgWrryf1jEN
I+9mw7lue/DU749UZUo5Jk/ukRaaOvWH+wTJbeguRQLzBmzaDhMpDX+l96Reaw7F
DLeGEpu1UtcHzi+ywYLgMhfXjAXGqMP7C66CUg6DOXDzLQOEIQvndfwB6X43ifTj
PG0nSHay7H5NN5DXKgPI2l8mUnFiyq+REB/HQXPNYvWylB5eLtx1O4bDftoGVrnV
KYeGwZUYc8Z5fS1u5Rm/PXMRzrsumxv83vSKnNeefR4lB94KNFvgWTWiCHrmFjsX
2rdul5ymeYuy/7+vPNBD8+Vq55zSMERtBnEydBImOZihT1uamO/1UW752MrXIAqM
aI9R9tZX1AgodaBF7Uu3gOcxK40lJYcRRG6YOdF47luifBukNmjvUtJU/Eqo5Bnm
ys6YcknjB55BJpx6CHww6k9yoFZT1o6AYNQBTb+azXK+rqD3FDlm5JSr6n/EIxOT
ev4GvA0+NXJLO7l/XY05hvho7pkHIIjbXIu4ltYkn+JHWpIRlL5T5i/ZMPp6lL33
YkzKNKROnjOqEPaelMyQ8XTaaQuiAOyufZxUHoOMmgqXzdd9c0gefhhzbVlejiSk
y7sQMGLy9/gUWQqgQjrOic1syAxpKQkSVUxbxuGyaiJDzawyrKQ6dpWvQFMeH+XB
OE+f/KB7JgXix7V8ZdydD2IMbNiW8BKsuzLEGqs0NrHzaIrlKLjcVFKIISgxemRb
LTddlFdWkEhdViYwON8gy1YqZugx8qUwaCw4iBpQFwUg89zs7PlYtJs89TJpsLUo
wHbEKF4/mROwkCBWeheTRL9nsED1rH7llchNx5EJBQPbdcKQHruU1lqRMSasZTeP
9Uxlto0lE4nsTDb9rRuUI3++BR6EHH+njcoPZfNJNARJoeDVYGKSJTs6/VcE0npJ
OxNV7Qm1SAKZPLNra1gW0gzusGCuljUOOrsocr9J5EUX0s4gid4IPA/SO80DlPEg
iYuMQuWPU2KPrjd92GmA/nQlPjC82mWunNAkcmPT7+Cb17lZ/ohZ3LPDFRvo+wzA
lJ5i1RqT4qX7oZ8YeNIzvYJxQZ6+mhnKntj3YQQpLAid63r5ou+MOUylV/9SsNsA
wziMl1BwF4sBtrqcA34tIbq+SDSqgu4h7fjECQLQuvUH4RyIcWjCSlbIYY2ZDRWG
NOo/Sc4rBleYMZ8dBp8GULjgnR8cfcmbNwrp3E/aQHJcjxLyAqMxMcOHHYPAb7Ay
gnGpGw2NzOe6QPnt9hFNgB3Uf10B8EahdCgrpWRf/8QQdxPYPyvdzgKzCTC/PmZB
VZhAO4G4A/WcASHMQY/D2MXEPSjJgI6m8VCrRO8fohPDFRgIWs6sF1ZTS8KnwGnr
1BbE72WtbtkpHDe5o47fAXE1vPORBVxdNcKmwVHx1VHaSsHhutx4wYD2QNJ1kLt1
kFvCGW87fuyYRF5GvPhimL+Zf/v5/FtCQ3NXzhAa9hF2F4T9WBC4xXJqLjqxUjvB
8am9J7/n01Eeik1gF9rGGZN+nxikG3JRsuBoaOwcqLfeuWokV3AFp66O4PdHgmjJ
tJclUKsMh9qVBweRuLOvsX8WL8THJ9xsKVSmOLYMCrU3qYi0V+Vmqq4lrkSgRYC5
ZZOy7qCen+RvowqB7JPE+hxuKZrpKR839nCbPISS0WF01B998NOlzuhB62xl/Yiv
s7JorcFb3+acrH7dG6KXuT4OaEigtYDqsR7n7POU5nLu9ISyqYWkgW2ivt4vUmXO
lUcF4bFUhyRHMzlrQDImyut9BkReb/lSiakKZh6rxkJQyqeMv+P6AkTD6hWmvYAq
cAw9ub+ALVoCoO8+d7Oabxt+tg6trbyHGfSig6ebjXOv7sgRX48YfwDCqgljvjnU
ooF0creN+ULYDeAYnuATlcARit6MLK9zTwtPmpdL7JE1Pg53xbgqPcb+ujhrLJdP
MhOcQ2v/updL06bi3Cf0TaEnn/4uuV9ApFBS7p8PUl45HtXFcxCYlSjfSEIwfBwB
OlTgao6FkP9ROn9uXoTPjp3Ie7eF7wodh8PBR37rHM9sSmS/CGOJCG2zxO1hLfU4
+PN+GIDHsaT7jeerKA17kVeCMS+oofCSt/N323XjW+XsnGxKYoipH59dWrY0Ol4B
D0ne66kQr9H4Cw/po1gGNWQeRTRMMAY5A9Z5jk9JjL93V6hLueJMOcdYYOZIo48t
bx77ZK24hwRC3KGo8iLjbLBsRAHWS1zhvI4Vl11V+yXwRYgCwmrm/byS64OAyEQJ
bZiCTge/omv4mAGiRz1Ud64NqQErwUSsoe7bcWrN69/PIdu+NbzqMSh1uZ7CNZmG
yyN6J0XD3yRMfCm6smra+expB0w4Zz+VjZPEOYAPn8CKlvJJRA1O+K4RQ7fA8EJA
blHvMX6qI7z1CT2k4jQzKHKzoSfQjT6NEP4qCfVKWanc1SzMOfRtAo7GmBTnDHLq
WGbF5LZTBhgl6wArqFr+A2pjqalOZn3Oq+XR+bah/9cDr/U7tzzjMPEr3ugoaaod
2TEiBizUQkQauPcpSH3eFCMY3483rJSC0oRR21t1n0R6s3K6p5jdMabUdSMt+Hmu
KbFa49MMMKlpckD2q61KY9hZnxI4fRil8dYO/E6HpPbU5I+4aM/4x0gAruKFPAd8
U+AdbJTYetSxyRzxtOKKl0PbubGg2yxwHrBEGNYvyjWUXrFoCAyWPRS2gqPOBdik
V2W4fzxlq9LZWUk0hPA+QPIAJ69jY1VbfZkMaNlZ5hXY579a5QdiVSb4YITzI1RX
CyclSUkMVtgHldYE/6NIIxs5yte1rih9QSvgq2NtHY3VjO40K12hzuldlRI3eZ4O
W8babPd3MoRuYzo//XX0rzGbiZngQb4494/9Iw1grUun4SE+dcxke0biwXhPe7ru
s+jjH23Qo9lqrMxbznZKsGcDoOvWZb0xY5RnT4MWjbtOo5O4n70nKTFWeMDg7cMT
YwqvWtsESrNR8L3DwPbP7bFz3Nl1/qjnZ8rtgVljWpfaHef5Zu2M4q3fxIMzpP6P
e6vbJ/YPLdrlA9iObUSs1KdB6bnwh9yifu0BRW38SniHZIhKW8c4TAp4OuNrfWuz
5dtLGg3zaT0gDzwmoaYbYYB1sCuUOhmGj1izb/B81ArYqi+EpdFHp0l4xFf+S6Xn
iS6u8K1N67CMe+PBeb/fE/vYJqZPoNLDXScfMNsGvKvSwQQhBEKYeXVi42zzKYvY
I5XHa4EeWDBMbHLKtZdfHViBy+D5fe99Ubmfs7pwjtFAzWilB/wbX9PoBB8fuJYi
u3MSVSpQ+MEd7r+T2oNE6EmbnXyOIE9g/s1SaHRLI1VDbOAfasmTdbqVObOGOLwK
FhgQPgsA6dHGAj4BRrq6zB+LtUjSwzJU25uWluzb3Nu+pudb7+FLD8X3pe1cfBJJ
pQBhGl2BbTsvdIT5s9rYEgFDvPNR3znZN4jAXJ5gMvscPV3/E0hlA5ncfdnwvtXk
ZSkr+kt9LnuALubudLW+ZeZvdpdgpFmhZwHYS5Gpa08hRBz8OTTOeZurBwuneNxP
qDeTdiAEKQkCf+qoyXKxcczdkozvwJIAJ7aH7behPA7qQ8HtG/1HMhXKj+HwMsT2
x1zzSgnykjYc5CrKX3DYqaLlzfm58UjUnLORPO22ZD1GRE5GfjbvFZkx8Hl7VWNW
NjlPkA1s8/qIXzhDVgmNpytd7oIux+60MQumD+GblHUl7sEFNTQCKQwAZIT9+aOH
KAlqmyIAk79TTJkxnWNqKNXu2uhjJZKdaWjfFlBsVpwtzJ+onhwlebYdZiasg4x8
8OBDuQCfiyrKk5hi/IbjQ469HxSXUGXhGl3XTT3BtMwHDSnyvtEwUmzGHYNjUT5s
rMpyY3OBBhYWIL4XrpccuyvIJ+bCmcZHMKzcBvpC0dbcJEUsjpwrhhrVOK+gv8wI
/7ORsOa2aTn8UBskNPpPEBjdShiWvlcEua0z/EpPrS7jI/8bx+P5SpqPkyiVUnRk
aFXwmzO5oSu1kpcBsUOx2aZUreWdaGn4YnJtk2eI13nMRm+CGT2WB93bh5LpOZqK
FIFTI/C0F5V6I8Q8dLzr1dWDXiSJi5GZ0LU+IFY3abD1aCyhuNNbcX3To+6MupL+
KSxShxWqzui/K8OnrJyfF6qBGyU/uZqVyDAh7ZxW9kh/RkDEIDIfIy3p/n4pEFz2
cDnUegInQYbpgdRObxNbZhQGPuzVOnCTFnqtXdFIJxg1nxbjyoJb4lopzjrPYT/j
t2CHtx04gWVhWF717Ncq9AGLhG8QmdB8slv6+0Q2kCujsUjiiGwV/0AR2ZUfovdA
19EVCmD20Wyv26/07ZA9K/iDIESDafY6Y+C8VoJ5/0XHgIqC1D/nkWy6Wk5gOiKJ
5K4g5SsvIUmwOHs9Bef5lmmACnECytRrq81awN/LxScjw3pbciGV2HZcJnwACWzl
iXvAx25YRDlhvWW/wsZ9BlJN1TCNsgnup5B4Ri13o6Al30Gu+oHYYifOFW6GcD/X
4NfZtPE3m7S374QHuGjlNUxBkLMk3ovXi1jSX7TWDAHT9TZghhSVQZ0DDesUVXhn
zMhSUUlSmvMR6YsNIz/WFcH6oc6FLcKoGHnUO044jWQwp9p3yiTKL5bRRgaexEKz
eYnBEbS2yihXWh4MXBTXAiOSbhVb3ynvutUlbsTp9aLLbn5oeuzSCu1Xo6eQJAAa
UVWP1+z4ohXTIFgaIqw/o+YZEF/YM8EvjvhNpf1+54tsVr6PnkW12bLad8I7JWy8
C1ofShwToj/COw7XSeIQr67iBmUdAd36W79UfUumrrfyltd0uHtFjl4hOdj/u4T7
ZE7gpKTnMZX6lZ8y9UOmnj7nzXuPFH1tIlGIHfP/T/DK7t4gHX88iKL8HFJO8pye
kQeigmQKc4AVJqw5+XQph6bdPaYUMgD13B/kQUWgbC2VyuSFmipT1f+plS3KMd9P
yJEZVhUZYvKqzVKE5knMcTzdcjWz+GwP8VQ0+KS/sb3xLy4HvalbE/cdsTyV1xCS
hKDiMI2VlUmCJDhs9VHQCUcu8hwdayNPu/WpfVevK89dtOt/s1gwtNyGMJra9bFi
hjEXziEVTlWwDVcBH2e41+Ny8M+DydRTlDC0DvNZEMPISXHhPsX+a+T8Ax84thKe
MMks288i58F8FNUbhHbi+5/q3O8layTqQBjwKtIu4l2VGPqCzMIuKM7cpJ6P5hX3
CRjfOkxBQnk4Kd/V8zaqojdFn3BT3QCKBGE2exEt4KDe3pK080pXQw6Lo5WMACQi
xsGl20jWuk03CHnhovr7gRTbovdbAFtHUXPsN+K8Fxvme174Q+i2SE2pvCcaq9nq
5FX6d9MU/sUXZzp/GH8bhjxDEkVebEshgdJ7oyz4csREy2OSKJ62MoKDqkKcmn9A
KBXu5odpETblqClNh+CZ+aSoj0/MJxzhRM3SB6uLQ6MoiIy5knFyf7LRcRhYaMAo
wEAo1yrY/ITBSWkBRrK0x5klbJqFMvaMBe3jj0aZ8tubsqXa1gP3kA8yu/veXYRZ
gU/BvtCxg7VeOi3dz12KXayoGHluiaem6sjXP7nzwAjCcDKgiLCpNsYFGo3afoKc
6B/8qmaMhQo92INattXThzdTV+8dMBt1qUtz0lH+IJfALFhChZKYkibCk23UozOb
tpgx9jzcIZ7+eaLe0RV8oR9iGXMMssb8d10Rcm5tABX/qd6sL+CBaXlOv+ZnY9oO
z3BhS9Jfu/yDjauZPC0jva3BU9GQgVfm16OKiVbUG93zOhUOYS+7wxIe6/eR8hvA
lx1Sv8RySsSAQhjjGWPtfl1ST3BDC0CSfVZEpzvYG/hJFlWHYa9E4ty5uD8WcoSP
W4NjQyaPgGdZv/Wux5OJj8fVpSndsxBXeCLXniSOdyOA6n1147LMfe1bbQFDvUnw
hHEVHXIDoWmAUkV0fPWX3EwohMy5cGclTFspJbukyib+8rcXdm6w2tBxEvKdaBj/
2cIRCx8miCH7wsLRwIYlkOiF4tyQgIrMQ1VwdbaRxIyV+sf+f3F/eE2B0w45XJ8O
iziS6gXAtR+N2knK8aihl41A2PNgr+JNQCfcLkWhgcb562RV8gOucSmRkKA24LK/
VsOSTz4O4zEyOw9rN/lFio7zRQG1v+zUlFwrLme/zBbAPOKI+jFViTyxOgHa/yLk
N1HuuD3PNZ1vpO46xh6t/nd511c0CDna7bBMp7HRRY3qMt9JLM/f/T9KNT8sRV1s
5l+qoVpzNyBb9mxj2FY1lyyPOF8YuDtuYIHdatSIUz1R+sutqF9CqhrkP0B/skJZ
djyphH5+gktjfKWWfw9Uh2k1kSW913CspptLeRR+aNi2JYp8Lgj7biwwn9nzC8FB
NGNoyelFIX4aOuTPo41p9G5+BjulCuMW6UpT0naqP6Ru983NOgkhpKGJ+klmpXIt
arAiwa6YulZ8VCUJWASUuJvdP413dTAjIyl5mCjhZPg16f227oR9TuTI6UQwrZGW
wSSqN/oZZ5a3jEuxlPxtAC5/6yQrLQI37H3b/ex0UZLftnITL3nVMEmlG9W4Dicw
ThnjNyeTJs2vBQkSP2LbQc3NM8H7pKLEZbbcqcO9IqDyNnl5nBEyrZ4KUbl+xa+k
g4UiLDGgMXbInMYbptC9sO03p5kI8A2S9sBB/JLT6lg4MhodUXac5JqNYMPIfRdv
VIjER2ZuuCAhus9PWWxdsfFUe0taodgfBavYCRr5FwUVOsxAyRbdN1ah3m51/4qf
6+uai8US8eQnOba6ZXiouAZk3Xff10y8xb2k+wqfwbNbCPMIHh9nLLOC9V37L+FN
1doVyoPrZ0KRirfITTgq9bseGP/W54omdh/5PdppoTzxSCfnwoHJd9jXbqLg4VLZ
/OP7KbVGcqcO3B+qbRJM4tBFdlLyCbwOLxq83Rjmi4mqgxlBPoU6/lDxdlCSv60r
qj0b5RvdiLmM8pp39W+9MFS+xuaHHwgnCuPrfVXZb/Mf27KtHpf8viblKYRhXQLs
NzdIonmEUgXgQsBnBAYnGJJDfOXMGEgMo+OOK117vnrLHx0gRPMv4scnvmMsQwNP
S5scHq0RSSUe/PUg54QTNUXyDuKIVdickpdBUU3EBcY2x9RA8O0eJ9Rhsz/j95Yd
d3d/TPiqjKnjtb8LiGi31lQxs0pArN3YI07ejHU84ClLMYyc3xnQE7yRQNgMjsu7
0gok1jzgZA394qtr3qxCZMbk0BUKLXHpfuXJlxER6IIs2zDHht3FJ/sAqyfPBAfd
LY/5HOFk2xZhEpLhyI3A3J2Y7B8ulhqPSl17lvip1c2rndkCzmsydmhrN2mEwZp7
igY+EoonGAzXjH3sinTEqxrj3a20jd4HtP0tERajEmNW7GUXruW4VNbhc5DTMJ6O
iOfFgAKyysm9Ha8+/YcVWsyRhrcXNw44UTxpmnsapxG2KalW2C3Johyb2HXOlncI
uBtB4+loGrDtrTMQ+fx/k19n0xZjMZMUmh5oWFp7bP+SHDyeiZGfXMruihlCA8IZ
mShq+WijuU73nUbZPAWmSFL/ELoknr4AumpPH9q7i3azuXAhqLml3NXV/eBNn4tj
42DZTWju9mpjhvnfZG84EscWA2BAzvOAq8Nk6P7wBQ68bEXkqN/KJ0J8cOAa1J3J
/9UAj96Akt6MSfMyX6jXzaiIbkiqWz/illdzhr7HEYszKPs7ZSZEYPw/KYgDm8an
uhw7tT3zOZLIa9GDdsBBnKQvPWUllHESIevMcYRbTfrFZYud/mvjDr5Zh8M/8Nwj
xoQbSr9D4G8QvzR+mizpZLlMnRi1FISX+Ln9W3SakbjevC0Dvi0dGgbiyyHOv28W
RAM0BmXI9hskx3YyT+KQCiFOewZVrq88UwhSK/zx+kQl0UpvCOx6OyrPy+Uc9CAU
ULXGUJA2xZR7v22Mw86h/jSkwTnweumKqb8th3unW9Vrc5RQMENeojDXjByGVXCE
2veZ7v5zlJ/2xWgkgqo+Cz9mcrVlflAT/PJq2rTt9Z8yULiHcnMzsQeiKSeQi9U8
X3AAzkryDf30fJZ45xUZzm8qjunLQ+HOMUC1W3vz13S2xDMULvnwABHE5Lk41pSn
j1sRnP66Z2nD0mVdoXvWqLlR984Q2ZCPRtUU8hzm5tQkKE9VAQe/S2o2pJnd6Sfn
r6Cp5pSlWef6krr4c/loyacye2vyl5suEi28Es9OqG4oTcsPl0Ur00FDScGIhD84
qzrHPEgwmWIyhE26B9PA2a1b6xwXml27ItBUayhVPKO1sWdJa999U/OBuAe4NtTE
Vvp7aLcEZQXsCZK6sYJdzcF6YeioduhcFJpAXRM4w0kFXQIJYsuiWre8fVVu1Dyt
jLmP/8Qj0/vnJH5dclRbep0C7QRFJDCvhJWxapsVJuxBUaZK5BTO7q7X/KrE6/AK
hhw7bgc7nvAc7k5vwDTWUTKxwHBkU8hy/xCCQZmwRFZ2+F93MUFr15XSsrLZZqy9
9EwDAlpcIzmI6RocFkpeMMOBrGjdd/w8ccMkjhzWDCYvLd+XbUvzp1tDHMELcwhf
KwWmRKIi4BPR5OUZ+Q+DEkBELiRo+DMYqy0IlLBdfg9V8/96TQKTW7f2VjxcZ2Je
GgjiUf0BFEurcnruCI/YcnpcfdtBNFiEPuMR458ZqnqB9v1iSZoF+oRhM3YAFLnd
/fg8ljlLBHqbWJ0FM5KlzhbOmSoJ+lzGoyN49/9waSuSAADZ2pPJcx93GMgkNgFA
Zgfux9aPncUj07wDrriV9LaaESofBb5trwrRu7xHXdrPbdl5FoS7DJbTBRanQRD2
sus4KXXs2OMHAR20jWQB2TsfA5PIYTvd5Twq0MbDia/D1aaQs8haVBh2vyMe4FD9
HEtX1cpBISkgUtUfE60EaOm2h4Mc3LuKad8HYCOxYZWLu36bgaDexk0aLJtn0SXN
839uBvbAhuifFYsLrujST7VTrDa2O7yCNZooZfDGLOo2vg1/7wJxFlgs1ENH/MW5
B3cObVKIFJrjBhcYyfXYinGCOy4xTnYY0g3R33wwH6E6duq5VebbBlhtLXF+v0Vi
U+c/6mdw4CkPRcehZpKU1TOaGPJbggXU8zRTMTN+nRlXiASPkU0VVMq+mSQp3ba2
E6+1L0bG6TBm1DNioZAEBYH7ntwbj+Ps1/7cNVINLfpfjsMSPskoO+NBEdf4OnOs
hWwGkUbE/pF07ZROztm1NG33BdAm8Pfmt7lcAtRsE+lij3CMbCo9tOUfRJLfZrYv
8Ja5WpSji/frJLnV2D/0qeJ6xWI9j28owbShEscyrvNgx4kB4xWVKX13Qef2+wF5
CAWzRiNhdOmv5TKRwO/UGaI27iAMeHbWdPTtBlaWgxqvg34qR+G20HEF2C6TVsF0
TOWl7EBhh3Jc+dE8nbDNhMCvna+u3gHX94aOFNhSiRkL/KB25jBVKGGj2idtGxtQ
DeDrHh9Fdbfqfc0mv0f5VdCtU3iDf7u+6Vg2K29QuH3mddRoDHt4HQq8eMNsolxx
c10+tWUX+11PEfIomOTLfoKvQ5c53rTottzHo7rc1m17qHrlEHKcCc9muT6+hGOp
1q27LUb2o/QeLB1pvQ5Nd6bXIhGG91wtfsev9YuDTBJ0nYjEQtgHMefw3Nzgcxaa
OhwGGNaEzscUeZXnIJBA0hoMpzMFRFUknTSTtJfnM0AEudrk6sd3q2KSapUah0/H
6r7lVH26htpV+ydj7azxTZlkhPl9oTMwx2o1qX6iJalPCBh5ZxR+1dKsEoLd0WKQ
tZACpnN2E89ittSNKNTbxQI1wdedzZ+DAUsTYEramqPTRburO2yYyFd0C0cYWVfn
q2Brj+E+BWfVsO2b7Lkrhd9KUk08LSS0a/UNa+El4dujCIcAKneNwu4d45yKsqNo
jF0I+yBnX2PVNCh2iAS4GUdsgW+anoXV8Qz8Px9Vl544PwzeYlhdsy29l+21n3Pr
L20nkRXVzCwCjXt6n7Zghf7qHdKKbJN/hWGsEe7MyQ7GptHUAf1bAcD0+IL4FO/N
K6n5GCWPcl0zmceVeHgBwdTC7KkvKgT7twa+E6f8gE3hlrSgcFTbLRuEdmv0AxNi
Y/oSk8hhi7EHeeV/TvHQXnUWhVxs8hJRQGEQ9T8rY7bR30a44gx65bXRM5mhQuYV
TZpKZl9q4MAmkhUmA50zrEFHzVP1zpRVfqqKt18AjpLjWBAru7gxxuPh6GZwD48O
9t8FG9TiBs7mhWSiYUbfuWSTcm3GX9PXQMItlJUBiLmf69pocZcvt2sWAgZkqbYp
68WDHBejUoDuri6CvN2d3vv5M6r2byr6haYSM/H99Fm4+u7cKlTKJ8SXbEllnHY0
i+hov80TCMDdLmtq/9ykqas/QEMgi/p9SdzGlzM8b0E0o1/ZTYTi64t3cFQ6rUfN
D571vzyyMmCLgs1pDJkRr917Ux+i8xXPKXoG0NYy9VVBPQppjprewexoZbt3xOfb
r/DGEOUf7OADYs3bddri6cMxFgTKuflXRsQ5u7MomQ9wxT1OVirwp01n7/z2cOIc
6A//Aunuwx53fwqu7UVxbEfeeDk1kGbuj2QqjJRDkmg4xv5/zkyTRDkZy3lSf9Sx
a8/c5fpZcXh36qDD7zEo2SU0E8Vvs+3a9HKE2vgaTYEz0xI9cUnAikZ/jVnuD2g6
IIjLZo1+Ccv7/tGG/ZoCJAs/hjlJRu8kSxS3yl8yoC81oXmicVkM4iUE5lxmAzbM
0tkRKVAMQfqyytipfao6amaeEK82QjfWiGfo6Lh1nSHDtG1u75C3xSdrezxjMgzA
liQ6FqDKSkqdgxneoTrmhcJyViJuG9dXbgL+NJSn6hTr0HfwWNVOl0LfC9WTNhTg
JxdY9BY+Zgxad2GyrTSRi/11RJRLfgPl5Uum32HTiR2GzRQIz8efKneMW61NGvRw
MYCXX3UFDmaSwmkVbMrg90ZvpVvXdP7All7SNl3PxuiGYLZVzAKu0wyDZfB1/diu
5SpcFiPkaswHmOnuc5MtBZg1+xI/G4jWTNFXOYGi/QYHBQ17nc5nQyEkyCLsz7WB
7l9FdObLjf2hdlYJrlyYNuBD36RabO+s3gjQ/CxlIOxNWNyY6hLRJ1TvQ93HZbqj
4xxye4JbGjZRer/g2n07yoc6tMkQbMMXaziDF+LnnN7ce2XOt7atRGdTr0qiguxJ
Gap4bcL90Godq1P1+tupakZfkZzb0Pv0GB0YADb502xvqpkS5YrbX6mFWtOyfh2r
q1LsGPRCx864xwO8+uXWHZ7HUd8lKA1Fyh1aTGYYz8AibevLSioASAjCwX28CIhx
RqwnN0xW7/tiDryl20WIW+gH3nwFhfgjFEAUHhX8gfApU2lbPwfspHk+LUllEM2B
vXVAXh326ZyUss78YWTITFxKyh2XQvluq4Kg7k9C4CbRUTTpVi+kl5tTYIFIrsYG
yV2MERDuintZno8E9hIIodWiz97sbim4IIw15QFb4lUf91bF09G6LNaY+/W4MoMD
33o3pmqcces6NNGz5Z+NDF/BTD+q/ziGHfMRwKJogHWJG7P2LzN0mf3vus1yL/g1
E5M0onqnx83mgdYpY8Tt2gZlAoWxc9GdZnzq1gvGS4LraX9q+AHVBAU2D9GjQWx2
rMcMT/kUY5/i5diF4uRS05BGxHLoCXM52YRQl0v5NfaRtEICwbnB8q1pzRH9pAGV
7jALEPjuBfqDxO+s4QSqxgnFfgQ1QOuMdRKHVJ6fcs//MVLXpvxPgqdAShRqVYb2
di4NDVD3pr4YnUCukzkzQlXZrTXMWt2foZbF3caWoHdaoXLhcbkTPfosWKqu/hcW
RSYUFRYMtz4KP7R9Za6NH8EbVesLM3BOaJ9FfJtWY29zQRVp5fzdu849BHDZOfSW
ftT1U8RHZw/cI7nN/Wyf0Cl8hy0ED3Sr6TZNkrmW+ePueQ0coNHiESPQd+t7ojwt
BTmUTnfwehH7XTajAR7nKooTfzEDUXdJE8E9l27ttM/FkQkso6CK0TTyN5IpCODF
G5fkTKSPa2WxcdPaslDe2u/AweIzuvlf+AQzBYLzX0eX/Qr13QRYxJDTdOALB4hC
BgvyS1biRWvvtqtVFqbXZ2YarlJaabOKJDe+y8M0K0tKK1sfYjC918H+6sEldi+n
nN06pLKVm0dhpGxm1fdLClmcf5HJDv26S6SVIGRVxIhM8+vQFjB32iicWv0gF23j
LTtRR1K+uKZHddeZx6Tyc6r79dgXiOxy1sHOHdi0az5Nhc/QWn/iT5S5JTEDLy4N
GZQSqFDnOJTWY/cvSD9X7836F+useihZDqNfexbSl9OqdhY/MI1aZHnmRxLQ2w76
Xsgiwmw+TaUWRRLKdQqyeG98Yr3V/9ziJg4CviRP7e6bidLZuXUgKI+SilDZ1zz/
vtWJNhmze88/lJTp1l3DqGu+f4ewIOzwdVtC7KRtNTXUuxtBoh+Sp2C8FKPU2anQ
5HpFDDFlYV4kKNElZT6A2Vd6G+Wnpj3l9/vgw0RBgjJTSOkKWQOCd2t+ASDi7Kj+
QaLHtMSf0MrCfd67bBRsiXZD2mv5DLnYW3mZn1bEd8OUgJ8MQtOkIn6TkZ0YQnQE
6XCitZtTBixjT82X4xV9Cw9RgorUGPfszt2CedbZpwyZHON/GUn1jw7NfDz+uR/W
tyd//RdBkT2T8dHU7gBy07unTqA0UgBM889AFP9wn0hQn6p4D1LZKSRzsklkE+8y
CfD3yGiuz69sa342tMdjQmCdrNEv0WsAqmnn2MYbY17Q/ET4OlnrpKkvUDL/7aaM
TasGglOeQSz51HAqFh5UcS4a2JZfibPdYqKOW7jca2VHNEUH7Q58RFcIX9wFnAZ7
fE8JVHFb3Hrs2Y8XrXzpfJsKgfdEiCs36Wm9kP4HEdc2HYFtZlps2OrDIj1KjmwM
JBXSFjVk+Px5rhedFIB19tqy3xJktXLoqB/3SkKIt1P6v8O84DejyoHe11qeNumr
sEhDHEIKTNdWH2bJFOaU6IAhlgDlEyZSL4IfRVhztwM5HPlbE2HsV41n5M2rWkao
JdPeU3FMzEc+rkjO3RivRlt98K+cj4pNgPMqEcRY/81Ks0an/ySKCvLGw9me24Rd
u0jk/++HkslEL55hGiv7MIrl9fUJX432JAqtkwj8H6fC+rlJNgkpfr0SedxzpuiK
tIYL29V8y7kdtSF8HA18zoldmMrKN5At6/X1nJjTFYq8ONWAYM6MaiwcClDegiDO
z4ngAc06rpQZQeix0lBlstR3izOIMyyKZFVHff4ThatWZefERXXXUST6BDMLN60T
oPEL3XpOurgnWEQgDj3M/SoE5eOc6ew/FRv3vOABvfpyyCjhmhDVT2b/hFPVVpH0
o0TJcRnV2wvSFJkYh6nsvvb95Cfn/Vz+JAuryEotW3EmW8RTWWwFTvsCbGmHKKU7
QMqU5h9JwcYwSnalKHWxJA+10JlYcD01sj9lb9F3qDHeDiQ5b1bVMGmsmTGXKLqA
FaojKqAPqTI0S7bo2HprjMFsoCM25J+jLMreoPDR5oVlZFIpMy8t8B+jfrzZgi16
Re60K3LUSlG/TwLRvh6/Q6nVJaYsdvXg/JGQVn7m4UOA8+1g0vFmKzUIYtb1pDyv
w67bmKvdFlnAv8OPePQfU94OmP1Jy3ic1RhMrZtfLXErVgKxgtsrU6AT90GCcRw8
fqFsBMdg204NSAA72yZ/SbSoPXnh76r5vln2D36LOlcDHNrJowsRAGnHfBYiwHVD
QQWTaYWUmUxVTMLzDnQEYCevC5l3xm27035Snk5KfegKiB+q1nu1DT6qrq117p7y
Bj1D/G8mbZnRAi3jRiUoSi8CeGMXvwPVmnoriHExCzWIE/GJEs5s7M+Gb50ntaFY
2slIDHdtFYHn3g2yPYwOZoEiD78egO8sH5CNA2g5BXcyxwNWyEi86YOBx7Hsd4pg
YE/iBSuS4aId6QWREdaI8yo10IJBstOwceBb8AroX1HDmVToUDqSQMI7WqH60Okt
4Wg5fz1h55HdH93ir/1XkeqxxZSd3AqTIy7M78slPs4i9f3/OBiQVDKBbCGYRqs3
A7PVEyApMMx5Pfry9Jo1XAtexOLpKQxL+jChmOwRP42Yo/lSUL9kxMAedy8n/Qdf
HGtO2l7e0bvYix6DHBDipyIupFfbSoz3/HkmhEH9wxEyysPvGMCRwGxYKxWTQQnF
kumkUpug5mnZ26fWKsI1f6ujbq8WKrMrD7Tg4ycnSRstSkIb+7F5HEVXS0VhmzPP
D8uWzWI2CoNI7JEajHS1WGLQA/LbW2xBsyorwwHCxAvAl6KAMByIywXGRvw60Ngd
jie0SifWrECW0pCX9q9mmCFUW/9+lWhi0XgVLRZbEK+fMd+QY+dBcUGFc+W1/5Jb
fPPwEnH1Zy3/oYerYowvZ3+EIGu/75Ssw0RkhoILLzsLInKLLvC4ao6LujK0gkpb
RdLwA8vlu4ufn+5LlTUDEvQZAdIfyRGIyO9OCajWBk0ABK7h0Hqxgs+Pdz7E5HZm
ZL9j8KPoNTEDD9cRhpYCnxTcj54zXQcwmrUVdm8PoJMJeLxTiIiB/sDXZqsJPEWC
DFKcDny4oDfWuxfShRqWd0VosQrhv5eKhTiVFgEz8Wbf8ORnn3SxfE5SOIcbvJyy
EnNRbiaAgZZCZrX5wqKZCqLEbk02SDRA1Og5XF8brooO2x2vN+u7YMzTuJ5erwzy
RST7Xbj2I4U8YBr8APt1rAwbKITacQ+lVs57BN5iMd3yHlC2IyfSXR7zW/GiLZcn
VrNRA8OvArbVNEMW/o1wya8ljFOf7nNuvNDygqNiDz8E68lMvM7mQozkf8c2luvR
JCUK6vKITvcP18k6Sh3N5fMApDcuI/CA9Pg9sVPyXQxFF/+p/b7acfQ/AppHYMtx
+TqZm7ufa0124k8qQHBHr3+MZaV6ZmiuRYm84oCrO7FXlEQg7dzOnojWS7YS77vH
vjlb0GMLhfwREnA8kOOhwzQT4DOLnX0gP7dICPUtXBNFM6URJwP64PWsYFw91I5O
Rkpfx7wm6c1cIH5RxhyuHbSiwaQ7cCKGy5kReND5tEPMUw/Pz/iVrBka+sU7FWqT
JbNlH3WLRXRY93CoCUCponN3vJnG7viBH7xBHwCobNENke9eNKavpt6i0bujGqBv
SNSuP1plBYfYmZFMkCCMYvoa0RQVTUkpn44kEzAuOt1KF51beicUf839R4EH/i/P
2E6Ia4UQ7PxBuLl36kpHHN66Nmfylara++BmcMgBY/FCW/hXeeWzStvunqv6orrG
X5pRQ0pjy8kKacJLU5Thm3wM8WFsiA7E8mHbRv6XIyFUf5DtN6YHkQExk/Kl/uxq
rfmpr/YgazVhbEPUrkoq2DT+6N8A5i5ASotYi9l2r2SQ+m0bUoIClFmCVR6DZHmX
BXNkd3m+IIr0IeaB7MCDJ7+hjSeurrAIZYd/Vswl6fR1d/vzXccZJTKb+PMFvag2
Xvw/PMB79v1lh8E/7yelalPHtZLiTtmlDWFnc9a5qAwTYxADIeclG/bY0KP0uk6L
mucaYoqlDJzE+dsUDBMCPPJ7jiaFiWMQ5dDvXssG/vjQembQVj1EdmaHHHr8iWi8
I1zsOlKu5rxaqcrZMILcFUKL3KQqA/svmViteyZTjY/e3yWEgXgu8TljbBFF8Z16
qpDvSwiWszZqt3ESwKcrqbJxDl88j4FUZrUizDKZ5y+aWrgYkhan3U33gg0TV6+3
9Ub/D3+pY9choafRF4wiEqXoFIKLyk/AKanGQ/eT2ZF8S8alDHRAD/3LBlpaUvKL
dtx3Ia+DciJcwX1up4zCE3986YN2DxEJ/anwhShHyqKWtf5EXvN0TptMQ0qE5GrP
S4HGVMBp7ZKPOI5MpJDv+JWmJIqzcAQ0REUNiQrQ1SeWzY97TiykGtWl5VFCD1Ny
OGh8TWa/nvo6J1oGiJ2wqdWiLOcqJ4RKAbTsqkvrJ8x8k4VhnVjtqfYNNqnveoz8
lb/tGP8djuIYOB+FgK8XkWmvQ4F0wjjXag9SSFX43ze1+bfUYmCyfj//mBZx+aQM
7U3cpmf5A98B6FU11uyiaz9S5RD4LQoLafqdds0FKh8AROOlKXU525vrUJ89YX1d
eqCxVCqKQjFYCwFeeHwOqCw86d26fAp0H6ie2GJ9yVhAaxnBBgRjCtNN41jXW7GW
Zw9QN48s/uEKOEnMyzLIubYmbRImKtxpp+I2fWkbs3KH7/QJKBqKzMrd/EJZpt3E
HYvT1yX67VBVBQibV1mQ3i+uFhMbL8310fkvqy2TSrhXSfE5gsd9mo2TRfHR85FZ
hp03tgfyszw6L3USexKx8q9TKCZm4murXQbaMRWIt8yi8cOUQxE1zPU3WEZ1qVuc
WSuFpKk/YJ1ycHRhrquBu9X3b9WtMzbNTCj19nE4Y93qB5aGBctdYe3ILnKdPANB
gRw5W/sO7ip6n2gTuruAte9L2O+UNL0Eys/coNM7xXOyVGgzRYsmhbxgt1QzWUkV
MSy//cAj22bgi8cPxQofquE9REtwYhV9C1sAnF1N4KSX/HN04WyftL+9FLmTrR1y
BF6YU3fdN2ZSRZUBG+cj6Rr1P/8Lg6TuvkVMczmtd5n/hTjEnmn341iQu/3q/kW7
GvbhksmI8gt0jip0vS6/byJRZ7lWUvzM8ZXqX89MYwHbthmKyiSeG/Mk2u/VYSrW
1S3FDai9JL3dAeZHDeFy861DCVgRZM8/M47cHGh3555aLawzNEV7dULzV3MRs3Ew
6xWuiHIB9nEdGvbLqqETrGYJnwL3lQCbxXlIJvP76Ptw5E5tYEK4W9ZCijZpto0I
hEDA8mXAPlbc8wFiCn//S96blPmXrdIJDslkEDtOvmOXW19J02ZG7ZzLKsEEHqXJ
bay5CPEQqclx86uLu8g4lrPUwXFqbFOUemb6+kqh0vF26aknWiiaz2z3rNCdXjfB
v8o9sfmnufCR6kUk5O/WM9HKSLbyPG++P86ypdDRKpa9/7u2gWM8+VwAfVMDvLUo
kB6j1s2HQhFtdZGeaPm+/TLEPYX6iD0ckl8i38cdobgiAOEslkgl09lSIZ0trkk6
wxXgQzwfN6nDIoSvflHCiUIAB0Kt0Z1JFAEydiHih2jG0reuy0GFX2X799WyZva2
vALjiuNzBNu7Mxll3EpsB5TnViU1kNtvX2h+wqeGhbWMwWYalYirQ8bIr4OP9LJN
y4LPMVEub/3C2Pz/CfXPRtuDHyhlv3Jbkgf/eICtIh9NbABgZVCC2R3LXTwQjjZT
cEypsYMFtFjQP0J+yAq1TwmgLwJeh49Dhn8BsvhmJ7t2SRXaPrJh6lTlNTpsIyWW
YpRpu5T28QYGxo2x7CYTXQXSZeM+q1AOb6qJBWRAyU47Jf+g4waOHg5e6tNFOI1s
BstV1VM11gQj8c8LrSmSk08TwwfvFpOCdZgDWNl5PdpdV/uoBMYj0rZ2Cx84YuMc
4iJPgcTqG83Rwr95RLzzLydQO4oLxCDfs6iIMUxId393+GCMevlc9p4d1JpY6dvV
4OHvMaL7XS2kyoBvwKedqvLjv5qJI1v8FSUHVHbkg22sXm2BqIF18oJMp71Tyhe0
gbaVzSeL/9Yw2DqQqjgh+OIXhD0u5aJfnNZGvikHV1CMJ6u2343XvCGYyhxFPh05
SLMkc0lPwXAV8UUJ4bK9OBqcoIcQ3HTdnU5BRHKmNUnXtMIYMLnFwxBnBNlMNoo2
t4Z1yV1b9mm6QQA2Z7c8PFMCxAqgOK6PRgJgHpgGViQi5+hBGloHqlhmcCUSd+gV
6Je9qJPLE8+Bo3kVIeYC7Ec8eBO5rjmIRbL4d/MOC67vW69Nn067T/rTBfjlCmA5
QrgfjKdloVTf5PAM0xBoqxmkwEI3ZRIWfHSirZk7p92ugTzf7/63O0uz2aPpLw6r
SIJB+K3sgvoiKFnbJF3mLyijnoHgb2y6vZybR88AUWbfDI08rxgf0A5a+ziRtPes
saEQJTh9TgilGP2nKXUJkkWjxTk57kWit2EF8Yk6jter86Na7TdtCs/uq0PlsMd5
d1JbvaXGdtaOycVSRY+VIxSDPGvkuVJMpE4+zpR6Ane9mtR+gFEVTEAC0aZGneFo
zUPnVnHHHe7Q45PHT9LylQPBfnzlWqPIOpX3gtS+E7TVGvCDf140pcnNE1CMYzOz
FvxUhoc1oqZ+sDUsjYlWNOvbNXJI28SX60WjeT/43QUHDnVwsr1298XG/9xMoSBO
QwI9WK+TCo3c/3fZEqIIL52z7wsg9xPvu+6IRhGlRyPqxHll/sYR5MW0kOF4sBwV
MtlDFotmJ1wcrMSSwKAeM5aiWq8z/Bnpn9Ie6ETeWmZqSR3lZOq1PaZIVqI9cMzT
zmR+roO/dXGW7g+OJ+JRcCDm93cUZ56f2jMz9iiCZOuOUCx0RYID/MuOeMCKe4bn
6KtrTlgeGS2q143+uJiHeu1A4Du7Gu1yj6hNfZdmyycp6HM3WkRvYGo3ht4wQhaP
CaSx/yAeEpcAhPpnHVLECT3ijiMjmbFz2N3RFu6vOwS+JCpa+asl9jP3sedXqcbq
bV0q0PXq/Tf+BCH3eVJkATZQQ1Uh3Q4GO1Fzoo5/1mrwpt3zUfktT5neTIp4uLqj
PQivrIhLacVD27k0GuYiuhOisMVHYXUEAwTF4e6i0nvWmxF84XmSdARf23QkIM33
3N7hWVNtyymmHaLn8LJy7iKBAw9Jk22nqNjaBZHQwRQSByfbSmUMg+d1d6PxG2/y
Dw+IQiP5Ne2AXRca6lfeCOXHNhEPQ+FgcQGJEUgJEsqabnSGcnahDP1CLZLp+iw0
W9wE98ZS1r5BR/av4s0sRX+g9CE2K3xnWGZjGaEvy7w1xi96LU7gNZjSQ0cLf+gP
LizI1B3MSKmyVrgKHHVPvByZIlt4CjlHHN85xB3yxXwMO70pvQI9StJYCD3GsP/0
VLDzMZyhkOviY7cfzZD7iPKjLTw/WTPjMjYKFmogn8qwOkvrA+exe6DBCBnrLKTn
XxFG0dTaCDEhoIhnjTq94tggJrDIi9/S74CSC13Cb1PSD06ezHoz6QsC9Yv24qOy
AzTvAnjXn4WhxiqdIEEa9W7SQLX9yeU+/iHjSkkkNALviZAI+zykf/uXuVbx1thg
dr5EVMN+SEZn+E5IvcNficsH8O7JMJXhnMnpmkI0sa77GCa159F9JqJapKTC3FOg
uc6hvrKL2jxrpThZ7bo4YsHJA61p06Q8UmlOVxfv5ajLPU4kB80ChnMugcSXDRk4
bcuF7Rbb5edICrJqAuZ0kC3wYmMgdoie57ZnqLUfUMG7my5TIox/U+c3bz5X32Zz
7JVEZZlWa1E2EyhqQirsiQixshbM2UYFyCufExFL1S/fHWnPBot3SJPOu03WUcT+
QJX1QqrP1hdAP87AEJD3IGyt35GWPxJ5vx0Ew4M/hsUO39jyd4+CLuPHaUiou0OP
6B7LwxXMe1Bu97rkekwPjba8FCj1G2851aS3a+jqfLdd3X/rUIvOZSw2PPIB4PJJ
tQ9sG0hl3JfjQPyxysHcyIu+N7pPisBcshlYnsnBgClkpUoTsYKpsiZ7UzPpMtnV
/Yj5rf0IbOMnvm5VACGhtvJ0G/2yWW3Rseb/naHTUTQxkIZQLVj4HSKyMDieL20/
Qi9A0EWdsnmDnWhNnw1Gln3QZxjmWsWHLXdF8WpbMxnFzLBFMFhqU0+bqvIIApdN
kOn5Flp25ZP4rdxYQB+imhFQeEDD4hecw6pfVIKEvamOFkIY50HjTCsc6HyFJrkx
rjXZ3xqC66/c3RllTsXwLjZ5G9tIM0BTgOeOWMrl3W4gjsRUvDfgX6ryjgKKqG5V
uPkc+IgTh/F42EYuGQdmwEhK7X4Gn0Ya0NNp8zmV3S/n5ceAPNZF8uA4UUHmOxPM
WDSldPqXZmtiyBzk1MqEcM0fpKauTcOUD/V1kRZtlOKrwpPtG9jdhjrs0zODvE5x
3yxczuOQN5ZB5kTO7SRWNDivazHg6TOmOuThyD3faQswTDdP/UDVoEs4yQMWdsfa
LjH8mibJ0G4zpl3yHKSt/0JpBqSN6YzrPskFD8BMtRfi0pvksxlG+AurxaxU+FZl
Z0kktdPP3GX6EoqhU68l4QO/3c5pTB3pk7enP3c7atHDOCPfCTu4Dgm+T8Ld9ChW
0Om1uI0E7aGRLf0Deecc/JvkNjY0Z8Ok5dVOOZx1PQpLJOUbtkoBrBoXDfG0D7iV
EN1ecTP5j2+vqGKbjWYU4P1iaeG7HQq3M+iTsIzzQJz70S46tLzEcNJMRaaGMEKL
3VCRRE6zKafjRW/S4gKZss9LDZ5yUjgyq4ws/vqJR/pSSbPxZMVqB4qt7XSUrf1s
ZrdUx8AiS5lpWxMXR8L3JQPKfbSkPCe6xDKp2sh4K2KAU4XDJnkZKvAcCMpaxKUw
9SE8nJdyB5cBnC05yUkb1FErV1JAWDJxaqjSxIHdFgqt68tbseIJtp9Oj3pO2Awf
KpR5rnZ57A8V7nyYh2AdQAeohamq16NytHDjghe6i/5cknkRaFCBNe6L8GORebhr
qlgSKLPPH77CBUeE7l/xNknqmVLIdXi0x714YhwUqQLkK46Z6ELy8Qwu1mCZDIxY
DeX75pTD1/DSAvz68pjcItV1tiA8sYXz3rTmf4ZkL6YATS9kuDddcgO4Curv/PwL
Pcf72TyOjgqGkc+L8jSJZhucAyppmZ4xz7MPIjxWl+g/vMlvv6daIke5dVvwmQFU
rGFA2KKR7/TIb0hIUoDvos2pXncxIcwy9QdzTqLn05KaZaIUd3tOg+eUvX82BnOy
NKEsP3Vs6r8P6fakGZKpOQcC9ss4FuUuq0sJ0VOHM3RS+R4NR6MxXQ7x/3QJbji9
mqH751oUf6DTLsxuY0opO7mgwLXzY+Dxzw8P9s9+3Z+ojW5qbWP+/IkYsOalymF9
72vvGgNQwk7vn6TSjmGBFaoiSUnoiACH5N9nW0oAtMSm6/PJeFpJACe1rLliEP+A
KUipQGzwVayKUiLD+R0FW9G31sQitIbNRCx+nt7mkFyXrJHqrG8nM73rieAwwAm0
ay36Fjjm8ZDDQhT9zdQ70SC4ddTYPaMrl9GDIf2ZmXAuX8OSkxBrngTcLceK1KzI
WtWdFwUG1AU1DsPcFJw/IRGIuewFF7TyqPSwBokZ4qAdH/ajsfuLJC1jnUupxEYH
arkNA3BPlFH5yGgcngTazulBohhEk1TtpKp7gCgG7U9XXpOosSUpbxPPBGlmR48U
CF6E/APdY+Md3L3cA+rpbbCDMqsU+r2RdUR6zIL/TJdJT8XgVtwMxyY3rV10TlWj
7SUcIIg2AD/nYor2UcVk7n558zB8aWanoWf4IZmlw5juk5PXdeqNXEzccgLGXctk
SFJxqAZuBb9sam2lh9t+5+CfE5UDmpqC3GJzB50ORDslwSvi+Fwzru/v4A5HgcSZ
WUWV5LkxZ4FrToyp0BMwJk6devPd5OYold67oX5vSkR7pYwYfEzA13MjiM9qGLLN
o/DfVxIufpwK2FlUajQBCMoMb05xoDMZZ/6DYOgGoV6MRfYsN30tuKD6zYEmuUkh
ByCn+Oenmb2bHtZEzrcne9fvXqucMdEvv4m73YqXweUrlvkxaR+CMbE8YvsOk175
rut15HkiyTBLapbSkUTSHoMWFbYNZQelCivUJ6fRVuX7Jh5t5qXMQtQyIjbkiCTn
nlM2VHw4z7J7afWyvzNR9/9ARtsn17kJysMxdxv7c9MV9aFsRlZDKC3GOgMyrkbN
z+MMTGtVm8HkC/zW8O4bV+6CcH2Vn59YkyUVvB6cFtm6vP+Es3RPi33ClgsmIReu
GDwIGTvR7+gr4rpOK3rGKfqt5xmMuo1NL311VxN6yG4huj2C67qjuFc5w7BmKZ5L
mBCU+4QJs9RQMUFoBrkubCbuyQw6pwMFnUDjz6lnI6BiGR7cBI5A3mCqxgDZFGcy
Uh20M2lmIddEErD59rqMRPN5L9m6nMQDweHllede+vmZuSbkZKLCE77++QzWNnkh
jY0NIqHa1z51uZ6b2WqwMFPdG0Ic96sxs8XXEwYNtP2A819rISeAuxRqLkyLKFEV
0fRBFja+sENxUWhOECNGH+UCRcjOxiAPupHCOwbVAKvxKV6oSaVG7ghZlpU6VVe1
xLZyL7n1jGo/2TT0c7of+rYopsDJTRHOet3LgyxEje4Q/XXmaRk4C3g6b8DYY4Ba
X2tdIaOiXUkh8NEp16M3JXCvnW/pli5gKbjFJcEJ2mtu9vqornZYoPgSnteAggxI
r9Rd7XpyyHuX39AbqQVBPWJc/E5/xPCLebzYdbWW8F+2H/UKLJkH//Q879UTAPC/
LluKxsIxo4paH4dnpNw7BT8KEQDoZvz4tE6aRhXk1WgE5jnbOC2nxgwmPsMle6Tc
kHzrlC+1iXZ24EcIuV/iBqdxtiv5601hQKfNvsTQJZYKl0V8oFB/E/O0yzSrtqe4
McRwx5hWfzNyRHa0UpMszXWKiBk59jhT+rqgKBu1pW786M4iHsfHlLAXnYSzMsmz
7qIBIQqOMpO7ugLERAWoBiYhZhgpB8IV2qvwWPKEQESY6iDl9wtNBEycd270r6R8
yfvMkfIMvb7RhqIB4i9QCVNsS38n46w4Zg1NAUz4WCDfCPxYvlCplfpvaWXx4m1/
N8iPJtibtFb+D60NbYk8OUuD8XKv7PzZmgdhzMrkE73sMzpBLcygSg1D73Uz8ekC
Ln8iortMLiMjZ++MxEc3Z+1qdP0eGqULs9cIAH2NIhGAVVrVxX/iP7OE4jF/a6sV
AzvUy3bR7wrj5qokO+E5ZqUbOPxWoDDbrW92W51EW2VMfie9aMdB7pT6MmQkmNDD
YZMQ2+y7XoYTMoF+8wPmbaiIKvi0AYxkbFyYXDGNOJGvuPIXzE4adFIm2SxFRGFW
PiY7VvhBSwA4XwwhfDA5LxXQ7k1yQcpAuN1tQEPSrLMKc9qYq6jxFoYxv1LN/zqb
NHUbQHnqYj5l43Eumow8vZT3f1ABf9WET71D03XDQNayjP+eTtlsdbjqbMeWzxSL
nagmNmBzsFi9p/OpmtN6MNKYYUfNHg41tN9thLrTV7KZy6oMC8gRUdLKCKuZa5Lm
H5XsbhDlNOCmcvTher+uIUCQ1kifyYmonpf5jKQwfarKAdu1LtFfgxoea5obHU2i
zh2vorD3vC/1cW2JwxS57knAttPSPlJlHyGC9YU36tiGdOIGpp4tISWJE12VW1vD
DRQez40Uk/fATjmSlsVm++VXZvnLI/eNIZhqyigbPvP/miBm/hKmfF43uRiHRwDK
zbfKTxw8VVCnitfKCieXlLDCMzHhkVVC3FuGIQReEFS9WG6RZ7ZSfrre9QqXZOMr
TtWyF2EUe0Br3SPwG/0grBtoMlTTmSvCk5NORctK1FUHxa0lJSf7RPE4nbQSHYdw
x+B+k1ZYbROU/WIcTw6JesoIxXPDr9bTKis05Cu35WczUCkKFYMzgo05cm84RERz
CkoMpIAsAmmiQ+9xgRxastnRkY3ylmqp5S/yyIfBqftylKnNKyTwNZ27xpAs9AVI
C6YdxljMc4UWBFL2Mpnw1EHCZHA/5a1rSZVf3WloN4/2Y0PXCvfgW2kwNybfLgbD
xcK2jhiksux8R97NhjigCcGWjPeBuhIRXF4xDHR9EcrCpoGvSUgVkhIFnTAkB8oo
VdDVqwRMliiAUZktc6OE5jdYVy4n84jJALodPg8qgrs9poouX/gpEPu2iHkegAQi
1cy7ZYTqSrw1/Cd34HNVnGFog+CsVhxSRIrHNKu2oQj+PfEOMQOv0B8pv1k3NjFd
WM6NXXjmEBkDNAIsCn4mb01Um/25fIEgTJYKogwcDb99VLxqA1ff3BnWnyLeyrIN
r/AFMAkoWn+DRev2jv1DooMNKdKhOaHHPJA3avhwFNLRtxFkBFE9vtHN6lhdhx6U
XqbTb42iu/rQo7QPyPS8y8Z0bhDQIiwcq/NNosfMRW1hk4BsFHKA0hQ1UiN5oIau
If5aUyxnJbHJNX4ZBVpKhfyy3/ATJ9Fs4g8d7l5RRiMknG/Aukbz/q1yzAW9o+aR
BGFKDLp+z/R69nPklc/ziROLCrhzRCWw4WcYLs7sB3XL6sByLEcGUvQp14u7ua/p
vwrRJmTY69A3DappuFRfVJKF2JlBj6/gP590cDZg0a3Nkn91fY8wefuHRiwZ/efR
jbL0Q9aJFPvAj2hsDGaVOIglI1UyY7l/t4ngmwYoQ7QxKDT3h3rVT6dArl9ccSXA
eCvF7/CVj9byixSzX/4SrFhLh/75X+0OhGHU4giPyYCcir7nmE6K2J/nsyv+Xtdu
eef+uWD9+xwIUhf2X1F/ksvyaVDuS6vo1uAboMcxBbnNpTVBiRcWgEf0ocQt2aui
oF7UBUGg32jQd40GhnwfRXsVh0xeq6kLWLu61KaXJEXNMXBj/F9Y4mWsk1KTkoJa
etjJ3IuAcARsJ+wjxGTgeAJXhcYpBxXxO2XEYU6Hjzu/MetncXCtnFepIruRYkgI
4HzmSGWa6/9fgBMcO0JAIe8JblqFSB8mEQRWuXrCjaKuig0XIjI46C4ZIUxJAO0X
FD3O13mRHQyDgaIfv1hJTrySUSRalg1yPVJbKg7Cghwhmjy4pLY6wbQfLwa0Eugf
3MoIjQj/YZPXJN49hCZqSmpgN5TtL74PN5VZ36DHEhSQ5rDwvijYLYUql/qJbgG+
WVDtvGgxAWdVx58vjtbqvRVuv+J3A+EFHdgJhgRSBYmemU0fhzQqev8V2ClFlitm
MVR4AcXWDcST9jpZJsfrkbeLH2mNuvIU0ihm+xZ+olrwxPSj/CI1uDbc3gS/k9rs
pm954zguH0hKsWv05J1ywQYQekiNZ2VT+eaDjVgHlRNgFUHrFL1wthmMoBB7AaEb
wJKLJAh3ZEvDcJDUSaQA51YQ7VoVFME/NWhjL46iCq/vJpwfrtO+v3LuWaD/FTXi
Egmtxz+S/G3swuLbP48gurb89GAPaSonUp/s4l8fEhbVbRh4wdUO7A1P+uyUEZoX
hgSBjizw3Ruw5kPFClZOmHjo2Mv+Yauv0t3SBVGFunu9MDZmCivMa5YYg2fHfS+w
MNyi12jvhbS0mTfqaL4e+V/jXnH54cz4Eh/kpP+apKYwM4/W7DKHjtM5tY0vEOdY
+1RYRIJAAm32x4245khGpVhARGxxufkIg2gRMFr1bvBEnTwru0JtDDuo+urT4wUZ
EpqxaVpiT9JYZS/GY0Asw1gaSxtd/utAg2skXOxLhiUBb72HZANCvfM2ygGBS+tl
p0gNNmLx/WnJLEt/F9cWZM85Y34nNQscKndAr3xfndmqg6HQK6d+hUpIij4AIN9B
0+XzB4uf+etQvbrwMLOku4OLLkVlWoq5UQKeJzHRHACZHVG9vC9T+8+rU/4ubuae
xgqpDrBjWYW/jECzlKvjqJlfr6EthEtXN1aN5sJqsRGo0g8ERB7O8uuR4pK312K5
NO+1JfM1dKejULCh/mfgXXIJiPCwTBF0XHgzUq0M/ZwaClwWzwVn8DIZjohDnLSd
Dvpkcsf4+ka8usDeFl9AmNeoaWxIBs15cDJStd/YIceNorJ7cOZ7qOAln2Gr32GZ
/jkXqvqtJHYL4GOg94z3wVpNVVOc4BatSKcC7LamoRsur26vgZO+FnmlRP4Svl9z
fHnhUnPhbkfAZwVv0BCK/TWk2scUYtmaC4Zt+BFuBXaikHDGpW4W2GNlx2IUlqfe
0PWJF+MXJ8LwgDq38HluXg1OwOKcHFCIyZJwr0er8LKiu9bxZr3hNsjoE0ZbrDIs
zFo+wLZoz6+vUiKgOBkI4VqTnSIY1/BV4i55vuQ7WzeI8Jwk90drZZCQEMgeOgWF
X3FyW0kVbIowcu5/lcvia1rtFLVPpwh9Pu3v0OK0xlfExmxtrvtjrvGqIpN+14ui
CfseE3WlTS+IGZorzGo8fSqBmEF9n9gyS7CQJhatzXJ9x8jAVWsS8yJOXvKO4w1B
UBRU6SOmzxQ4zQaQqAnYcv67wwbEA/ddRhA5oMwkeB7QRxmMT2gBj+jxqLw+vLDr
hoGfmqC/vXm+rEVaykWUoWGlk3LkmazZ7a1DI7oS/ZdtQgNCNocjPUJCVzIXv7Oe
k0566YLbYvIE7QOH8kUzWzIcdmbvmgIS7yYUhhVJT5WQVjcrkl0tqmGmg2YwTEyJ
oKOAsYTHeYp2GuJJoSi3k7hnRoxo6eP0VdgIUiAr19ZVn9KrgObrLbYDvrrjA8l+
5DL9H8wBJVQKcnE8SADbmLrnlnU+Pd/xJ4BrCAw5e4fqjs4pixeDgLBl9mPdHjvk
x01fbZuORTAEhBlhprFZkdUKVzG8KF9Hz1GEfYsAEpnAVpbQ94/DZuKuAK4SUpF2
yx1aZKQwDpAlSMAFxJAg7wI4QWDW4fb9ICy42ulG4kKhKQ2zBZDQeAHmURhw2GkX
n6KPG+fai9lWu6fCyKQb7iSw1f7M6OUVYngDuPCUCffbPrIPvco7i3eN2tcnufbp
5KCQSDqKBUZa1EYKVxPMG1ho7EDcefrtFYPaVlmCAqfaA5DZNnCErsKQzsvwsGzs
16X7FxgESariUb8bNGg+hR++hfT7VkndOE2THKCisyNkoPUY0Px6j+QYtWmWJut9
XLwJ5/UALYvwoLdPoeU2MY7s8bAa0dNgKecCbvdfPEhgl/6bLolhYHL1ONw6sx5b
LXNfe3GS0A/v3CKZSgwdsjsuMiile3skie8WtlcE9M6GOKvIOsrKn3LuH4o4Gx0T
ILMCe3MhxqwFYwI4KcY6rGRpkqh5rMc/LAwQFFXaFGDVjTjwlcw9hpzD1FTrd53H
isQHUK9Mps+Zb1fYIsdwDnI2D3ym0K4FPeuv8Vaf9hgBxD0i5laZSKpmwVqSH9jq
BlOaOIhr9bVJpNre+V1X8yIJ7KX2hhKJRYEsZx151lZLac3YFpW0BNH34uUdzaMy
utu52kAs+abXWOUB1yjnzKWZaA6FgIU4MSsr6hVW4oT+PY1GaxVzzZijpmTm3A11
M2uGN2V+2XwrcL/0oO6w2CgzrDrCO03j6OhqHsr3eH04xLofdpIo2Oiry1KKCX7Z
t6Cw4YWbj//e133L80R+zMTetyLkXxdAMfVMXXbFj2O0TQ0GJoa+m7zjjTQBPVJy
nCGfwZadPBVFL9AlizAq46iA3o8tItEUOdpuHTb3HoLuh87d7EvxLyKkfdsqrFmw
FXNjzrlpfwyk81GKU/oI9RTQTCsdw6va0djavRnKf/tD4n4PY628SdypkZv7sZGx
flBEHw99ob9evIBV5YxgUgP2SKIbLkVZrdBcbcCS3qjo+dfNbLamXkeRrSio5/zJ
LUVTlpkSa8ooKyA7+om86iH+Zek6esqu+VYuYBHJGbUbRBuNaHm6ahjxChTpCC31
BbhdsovEUHGK4gNM9JSrby8H5BfyYTgRaTjZOwKlk+nV0vSGDVJI4BFMw+7lFm6O
8kPs546JQwwC/4fpwxc4gouPKibjuiQMj/cI2BtX52v8kSLEl1+hpvbuf4DdBLIa
atJedml+ktEDBVZ3mmzfZbT3UFoXDRsAPZEVQthDCTJKRLO3IWGzT7z/aebHktwf
8ZwLYuMtFmOWkne7VPjoDgl7Uwv7zukQqevh+/JPQwSPO7M5FxcB7YdeVaQCgrV2
mmP2WJY5iUS2R/5Vi1+9Ozqy+/9u6UmcHzzIIP3CHfJZ1yqYsPH1eClLSw/fOwdw
SayXxDbRWOn99t4JbHn3QbWSdyVQHpLaoscbFV5Hat7L6yvGcwi2jkaNXplmPliq
h4rnZskgZ77NhJdzKVaIYJ84KZlLqpASI1p+iXkFfNuMyzVO+qk6f7l2CUJLTGdB
qkPSzHCcMSN/GcN+xw2aZA9LTOlBvDUg/FNoP54BgQac4c3r9t/8aSYjwdvpslgs
tUfz5ePtshOSCYZbjahiwguAJimtAwTa0+9lP8+tSwMihWMRV7+LJfYTFusbuRQi
hczIoyGzhz/4Qy6oMqFFS1k8ek8yB+zbwUZyV/OomginbWREYBd3NBidRrDqCMjN
MT6EkcN85jAMfw26O7OzxLybYrPdp4xrxmkw+4/LqUn5fGJoKjjP6DtqjMsOoEy8
op6pj+LY7uIKKbDpSVg8SNqIc+LT5nmwwqQlT8gifBco8cKxBbN/ph18lDsM1RgH
gX38hXn49PQBWbKN+emgY+9TPQo9GrhQJSG/h66uiP+/kl3vg003MIPTThXjBxsP
X23CNA9+geQfRTkirpvAk0OHvdyguKg9Nko1nw0qGjVDJ97lu4HrkbRYsiP45b4b
FydcOou1hch3wEYiBIyUAWR1JSW7DzffmIHzdDnYhQdpSRWGWLv9eWrvNTKD4UCN
+BajvLtoKhyp/eFcDNvX0V1NvR70Fv9owx6FdMsaNDt97xpQ0guOGBcgW2HLnloX
441ioaG2my8RoTUr9I52QEcjRokUlnnpTHIv88DF2C3aIYf03hhq7+00Z/kRQZdh
qVV8XMBlXM+5fQYyV4u2PwwqdvicbZ3xTVKashdsL7BelXQzjpIgNnaFPmoi22aW
8A58M6azq9DOZn+KkCfGOp2Xo8uJ7XgOuwuCSdIHU3G2qCVwEFEzcf9V8AfvBfZr
IaeC6IQppfzxyMtNY/FqXtiN5IQk827AWhBv/oulTyT9PxeLeUX71u/Mple5dGha
gKCKrGZphLIHJY1izKj/yl83P8vm1l4UjH7VCfA1CnfD4GiEPUqC9MXb0/S2NsfK
WLnpxuPqSn8x4xpCfmSrgAtik2+HD12Eo/TvoT7ZPFdjG/Zp+nPnfBKtnYGhnnaL
82F1F5eW676I1ulBvlNwtL6AjxQ/H+EZb7Bn/I+UTmiF2v5L3FBH5ABLXEVGMXzt
yZwyIzTd1cSqfW9WWBIPBPWvnJTBc0Wby6OG0vYNLyHwS8cUHlrQJfo2vwjQxOcZ
trs5ehpsB78Tj2dEdkSxFwf5lc5wO63fvBp7z8HdVxrEe4TKpnjupMh6bvPBBK1m
/g+bS9GYtbVp/0n/nqsh9iPf2XnnDem3LNkVjU/aGMsyrJdxK9PLhWATUuEDSLsx
F1eStZYDkTXEMF4YObf8ybjOCArEuI2j1071+iVu88pyoqhM4+SAjSY+uGDwBvKc
75fm+EGbpwG6idjO+VON+YJPUukI7y4vWrkWszHp3Gsf8Ni/jnJVj3m4qYHjkn4s
ry32SRn4V8MRq4rmNPYKUKUHAs9mUY0QxVMNOQwvZ7CCvHbWSpua78GFilbeuEtE
4vg3iydnk0C0hcZQ81SKZRmFCe2NGCYNCdv3j8kBySUsmrlnOBEbxhHAZe7aFYP3
VpDexJRzBYn3n0hmIyLzsFpPHA1tPGiQ95iJqg3o7GuisvCE4HT8ct5hBPtyNcA/
d4MhVjrt6XWKYKWz7gmLVAOEpM/uM3fWmHbCPaRLrLvfuhr6rdKjVCd0VPDIbaLM
cyXTv/03tqIbTDoEDx4c3wsAuCPgzGtimgbhe6hXfys9Qpwp9aIHg8rQJPJieZAj
QqhnRFz0lyIMCe1VumgV0ayK5+jZ158YjpbUPhAUy4WiDmz9j6uaZYhbVUqzi+LI
KZwQ2vzC0bOSn6sm+4J5n7Jr9+DjOdmeEYq3TnBsscFWHdFG7MugDHWUoKy9hCWp
7JYK0/ad9V/FUkH5ECguv2aNBAHzTCL+xJi7y09rqgVVkAuwn1bSYZxBcVDe1UBJ
rhVET2ge/zDsEb4asHtc9HSdmcVaD4fcQZVD+JzwCQ6TSZcVpqHBsRaeClAqNjWf
VycE3Fx5vLCZGIHCjpuiqERIYwxBlZ53J20t/ZPimgFHlKU7TCccHQODsgaV7CZP
g2nH9IgMH2JOoTMzSTNs9DFEULkYh8n1dHH3YCD9M4Fz95s2mbmzwuGDX6b5XnED
ka1U95xWfNXjYz1H3r1IEtC+oc/8j44TxO+2dIQHiuZ2dRN4Ci5pfrrpMWZ+mk4Y
vydpz8D0K965SOJxfKzchTuvOhSgijyteX2z11yEyKo7tRW2KSF0CSAg9KZsv/1n
ppUdBWVGHG4VQYJuZC/QRM9tTi7JXCalltZfxzxxlENsxOu1ugtCjo/3vD4PVB3W
wysUCpZ1/085Qqrz5yMRBCW9l0kIoD6by9DpUuoMjmsrrplMZsNL2BI/Da5yK5AT
QXnQ4S3mVMneJtZRTmsT/by6yw+hb5k3LksZmZ5io2YI/HzB4pbe+trhHb26BrZf
itdONz1qwqyfxyZ6CGg266vJMdRedV398ZqFouf4lNedlE8yP/72g90Qx8dXp6p9
64wAly8Ovv/DchvUVOutxpR8h+GA+43KL992HsiU9tOQoHZBrEOKQBJzCLBtNJEI
2BOjFQ1Urokpo3xNqgWzlj0ayrElODFVFD9EHMyAWoLUG3l7yk5NnJoLBaNQADYn
MQYE1Ko3/PlYc4b5HDggSG81lU1YR6Y8lmTmcJU6b/V7FmAwq/ONeg1gTS/AOddv
3d1y81iq/+1R6qYk4YTzh8zxAgNu7KaeD/6jDOHDb2p79y80NtgY9rQdEAGuLk8X
N7tN0LGhmckeMHdNCqYIOwwZRqKvD15lDADQhGfDzzgNTRgSEl0FYxfhpX9Jym0j
QKgS4dmP0RSKfRenenx/I9OdGM92bUtQdSrz3lL8PuF+GPcXAi16orMwpsOFnCM8
efxhpJU16j40X0W0R69yFQE1EPcbFt9KXA2ZfRLgucFMNTDVR8bMOU5nYwyjo+RE
dHG7winMwcpyTUy9AbRWt+5GCIbbL9r4MHxIIyMipvIBzzWDOuUrlud9lMLxttkw
K/cf2zcXmZRhMwpaAl+nHaIgziVFfGdmJ721Zmrox40jaAPPW9SN6AdYPfThuyGp
682oSDFjVlMkugXr25Fx1g08aQmCdYbmpLO48zuxEisePk0k8bC3coZq9efHafTr
2bKi/X6LTS9s8v2lY8MqoUVVyO4qi8XhvlrNa9pn7nOlSLv7BaSvTMgcp5Pe1HC1
O16ef0U0YS0FS4kvye07ToqN4dfFfDIJplNk2MI1Wfd9gTi1+Ei5bBFrHdzyGu+a
oI/fasf4VOS6qCxEqSAYncD1N7qvq2o4+vupnOl9cdVQWNlOUoRDlnBkidY/E+Gh
DdXnfhFMS4AAlydTzNGYkwguW7G9NTk5oSKQCIRp+26lzlzGlQrf/tP78kwS+9eG
RVBg0ZzpLO1H9Wq/OuvyQHVPaUS6izrQc2zpMJCwLcSjZ6A3Mt2n9CMZKMNe3ijU
zS9l5vkYWttKvEZAMPjePd3EUHPaiY5vheK2Y/IzE4LgTZ1Q/fUa+DoR2ugtbw94
s5f5f8Ss4apC0pnQFyLOrTGuPu8cNgbwvQ4FXXpiDL61kDiBIzJ4ApOwc6yC2F6U
vd2LKjRbh3qmf1JiNdIwZF8FAnk0Tobalh1ihZyChgRdeuYCX0vgOwNPiJ8UxSBK
QqizDoNxsRuh/GuyQ+Lz6klqg0wSttH6wpXLsVUakHvapdWqLHcTsgdiwE39bRRK
P9TCjgVYZ4Y+hj4jElLH0epoi4rCo1FvxxsRSVShUTSy2fS8TS50W3PkLzIA+ga1
XVmoxuiHH0aVh35mnng3V8WXb9jDH9SWD2TMhAWfSjCilLF94jsmhYu6n7KLc+i6
L/NcXVLa+U/3pmrhJl3gZZgVhO12l0R5qUaixL8Bo6EpUr2pS53+PM55n9CJcsLe
nGjRtYMO1poL8a2cvjn0aeoI5mT2QyFNR16B6Go1OYLLU/BNpzAwzIRrsb9Q2hZc
I+Z07SASXQB+CPdc83VdqLNS/0dytad1SLkB9P/UsdN5qZWxlnQfGhu9m5eY0fZ9
b9OL6r8rCqlxJixyghEP8uaZcHuBicUKtcE7/9pgpQyJ402W/VqlXeU6ZT3oVVgZ
3WwUAK5o0JasqgMMjzFblim6u0ZisFSiGTdMtNqRFiDfzkKm8FWgWOOn/elk/LsE
Zc3TKeVSNlLoGplHXjPujeBnFF5fvXvsILA8gyQqdCxHnTc0xLoMrs6GGabnJJT8
eUm249ovNuPTjQjWqmgVPlrImka4aMzpB6xOTGEgFmC017UjFLzBGxQSqbx/xAhQ
sCzlKUaVSXYvGYv82GHN7vo5iW6wj/4oDiWnoSinKhwqPq4lE06fWNxFhNhkA8Wd
nEGRkRs0NJCTILBOJbJIVjlCWQ+kZAcG60fFlHxvj3dfGmep0qJ4syKpr2lOW+WE
XVwEy2j7QRB0AnZGTyPqJn6SRs3sNnei7X56mqUhKIa4Ze6rZnKtDnVfKfBhpDSp
aKutIEcfNevLNiEyVfuSC+GWMY3tMNGvAyq3HMi59MEV8swTcqZqGFlbWByYvG4O
r6tnf6Rvg/dQglzVL4cAXuey0dtgdRbqFBKOf0DyvN4klVCJALbDM1xULqIAf//B
8KkiuP4uu5XvonRdniwIO+lgifkXUE7tLn8DfvuHtJwpcgpwr1Qt6LUluCyX1sdw
gkkU4KfRCG5Lq1ftVKfI1u5P8d6be4qEKe+2BsJ+VjozJh/LgF1LMZj2Pbz0gtxS
CG5wFHIGCmiFvl/TsvwN0bY3rUitetGTAw+BHe+rHrE/abs/TqdG0uMmRCR0B0i+
Jjht0GHEe85BH2o9EzLODt3lngeKFFT8sCJ1GoVpUwv4FEVz8PU4zflEFT/c8jk1
HJx8PpaYSvqhqWAQROES6Y+kAYJwjema/9m7lOC/iEMck7mq3klsvpdtIFVB8CxR
BqatQbtFMLInYkIYBM8Rqy6zXcz3kn9jRshqfDg53crpsXI+RvYJT5K2X3Hd7rzV
Zz9hNzFIHtVyzMNX4o/MxRvnDazlx/utJCxe3S3CkEnMpRuHvWHrVtzKmVY1IOK8
jEWud+itJyeKf8opGP3nzLpjfdz/VnUC4D1522plwOKDO9rvcPDISB1+o6JR38rf
YaGyKTYoi37yWPa0sX+5/zzLeGdvf+fuugi6SBSo6GBn5nooFGj/G06HrPshbfiD
i5MES+aoLP6D37YRT2couzfl/16G77lcPS7sH/EpxI8oGFbBCDr09a+Os6XM/K1R
3+8xTClmAA5OWGbL9nHfCQgTB6iqBZLtT1mGYce+PWWHzgRfuyk0x2nHLuNpLVf3
h6h7PQYAs5manZVycTcJ11ZrHz2O61yuNy5FSZ05MGftkZqOx0s5XkXUwOaXqEn8
TaGpc6lX7lc/kUxSlqvKc1EaNUUneL59WrfIslqZl/0z1q5n1RKrllrGwOSFy8W3
jCudwLTkj9ODtaZTDFGvAJp+TPbUiRZ2hMqXOO5mCGcGZf2HlWqbLm5UIit30U95
di+22Esus+UoWMTDqgcAFzFYSCvNA5aZ9lh+nFFDV6xRycShPtq2aFupnnAcGdM2
ftcPANz8fGWVV5b37oAwnO4Tax1HO0SbJrs6+itJjObe7mw1n9uxMPFdC4h58rt6
hRfudnlgAD67Ac9Bm1eh3Lk4ueRobHuP/qA1iY2H42wHzkg1mLs8igp66Y5iT8qX
GNq9gwlP0OrrAQFnjLnPJxiOV+kwsb2m1AY2foWCQsPnbUO/USYUHZDQv+3jFP0X
yROHqrZNJ/9H7KMW1aFgkUfq3ZNtyDuPjnLyC/MtOFm8GZSh7621zAbe2NgfPann
GzXOalGqB4xH+wILJr3Ug+4IkZ+riKWktUwvNRj0yzhmz9IJPxkCR9BbB4J9y9AV
gdw2uSbt9TKPJEdMa5lWt0A6gTSZRTooGW6mXGG87tOGNLhVSZ3Dgmu2MYtxWC+O
C5oGlpLdjnvmAiJvap28E/G3LRZnwcz+BKOrRsF9cNSJlQG11MLzOyQBXicCBDi/
Jkxq9PutFi2cJ7VX2tj4VP1U7hs8ioLKtGuAQPYyEhpVN8R3wZTrUI6QnREoJzRo
yd1+ATkXYwKljJKlB2OAbsRJN3AnzlyB2MkDIG2G1pES9Mch8q9FGQGsp6UG01+A
cZ2Uu0+xSHn7KnFVPbU3PXoQfqpvEDWMkAPHKPlcJdnjfMU/0bMCcPvoVDL2p7Bv
KkjXMfTpUH6y2oI+XNtIy43Hsqe9DaTEFcbdcyklIt4z8zsuOwyj19ubINHM4vI+
4ZY02WFQbXpw7ugYUIrPSmi2c4YxWroSzul9r+Ew2z6zKPHO899jGf9zd+BP2B3w
CFk57qsS/nzUu3+GEoXo32ug1jZqLRZJzq5u2zcNK7W2WfRHUywwN9B0cafzd5sb
0bEbSIoLASN1SCJ+W+7+gvn+1oMJ/zmzDLnRRi7cbGqlc0UJMZ+qJ5KEqvPUOuZl
3KnfInnCgDU5MjShgyaWlt6vT7ju+SoghwN99BqyUqDHnGp40Oy3+5S5Ss2uaQfd
UigCbwnCw60GY7i3DIKoJSDhozzHwzAXxGgaAwuCi/FGfAC/ZgsKrcX9T5kW1LC4
UEKbGocPwhGukiOKEew+xLmNVFUUPWRvwOvotQJgyl0JUBz/K/JqIz3D2PT31xW3
P7ThGUSvooOgPpuWcv7WXNITmZpi+3M5i9aE171Jfo+XyhkBDMZXGy+QDOnRhkSa
b1f6T79XS86DOBPDWLYqgdL6OPEehem3waqLFH/Elw8sEoL2wCsX6rvUWeK8ijNa
4/2E2wKqc+2zCE9DRuk8eNq1nuIJpSoGESlRX1dRAAjLVqn6YGQmVGrtsNyYes4/
kIoAsTdfSHNWbJogZvoKrVsb7OTDPc6UlLyeYi7BFTeS/s+Z35kN5gdLS95eu0Lo
RcDyLwBjjXPFzeLWLD2fcP1eVnkxv5IEqeYuKoHYy4KA1l2PWBZDqG+n1PRNO97V
rM8bCS4DA0hhhdkveL5pWnSMGVSymHT0KH5jghtldqMsnlCGrSrsuL+6UVDwjMjM
h5COGGMcFQLIjhAzoXSj5hT7qZDzIAaHbzU2zrilg5uL1Ds3cbWWslh7V0ZTWxtK
57LdEZnVoOhQ+YG5wB2jqgUKmgPBD7YmR6LlWHnvfVoQa454O1BrCKrJc4Cp5JBz
GuhqRUkyu7VzYpUCqn3NddXrpYHwwm2zixvrdIpU7CUoa/aAIq5eEvBijvbr868i
+r2tvw34ax4ebiiwTFovqptBkJzIlpzVIIJeos2K36wBqIJtpKuOAS15WVuVbUIt
hD07ox6kTgVOaVrjJ4wfXbERqV3LdBIuMarseT/gpfZ4dZYQ86gtMHlgVj/pVxOm
AoLHuiRq+KyME4VHQy/z58jBOAeT3JdKu48ihK/R4+HenTCcVAXayt5YaF7TI5hb
CDtBCR347H28vtRqt99jpxa/UMen8FaBSEgMXHfVx2mXBzDuCxFBjNsvD18oJ8XI
qX3k0vvIjioe0aoANIX+nc8RDF2gkgLGbJlR5RBF71FjF5OCWEywWERHNetuUvow
rF4SIjA4cEQOPK+Z3CT8ePJbWeErfwpSnn0onGRokyne9ofOaidv+3oeo4V2BPSy
rTVrSX65mWPXEy0Ac4uvUB8eleB5BypxIdW331lZwuBWq4B5pACP8LXn604YPfSc
HsaxkqXN5aeHbkCZOqNm/YRgCQnL9dTaGLfh+W/DatG+oZvb6dynKA/k7r+zMucy
0/xuPTS8Tk+V0WzPCDdHQmJJCmRsWYzStFOtxo8+qh602kZ3rsBI+483oAjt4zKA
bElahIoiOzI9b4xUOj37At9bNQXyKWvjPtC/DYoD895CddFjoG4ol6qP13qpXIwk
2nK1Pt0wvb7wz93uvSM0qiekzhvm+WueD23FgXbIS1kSkCcPjDanFDioeROz1Y5r
k77gaWv1R1Vn8oTPGDmBd18PC+iRYEpBlfSKZ+chfa5K66/w5Z/jex7Dpi5AfVtR
P0nBSDEgcM5FRgRE1ET4enhhoc9GixBKFFTlTX40GRZm7fRaibn/6xQ4FGt20mhN
WbEcPyPt0uOiZg6NW8FZqKaNgGgZLoFmvX3/HVwRPkOC9WGsg3MGrLz1+CbOpQUu
YVVUVmOtGJ1qK4N+IykFZGAHnl8IDIV15IO39dBvqCY8MkIELmzJOgeyT/r32bsw
ehDpM+/+6ZyUluMOjW9r8lBvbCR5xARObtJr+Hk1ldXIJoHTbmniUJfYg3t8p2/W
6A5dxhLkFtNEAH18rMzZdnQSYpvbDn3n01x4OOeS7+F2mLathXy/uXAA4immO5mq
tMDWmtbcIKZ+QELMzH2948sP94IkDK7RYEbP9dwJDxlak9s63Z2TFtplJPp2nO4/
ld8/l9G1t+sU1u3bvBAhEmF3JvLefFOKG3s6IGObtFLmYFP8Vk/IhG0cDT8d7XeI
VPVgSQuVCWdnJr0SBpKKYjiE/Z6LFq2X0bD5xxtZ2e75ETUowL+w/YtJLIJh0X34
AbnApAng7YczHSY5L7xs+7KQaGksoSw7p3j70jtqcixBk0i6J+d/OQ/zGNgxiU3w
UWcg8XjOLbCXO5TYZyHFTyi7Ml2I5N3ODrCeo3ONpHzK7mgwBjZB/q8/paj70amo
SVt5tFqCooLUcB7/np/O0OJNFkLSFBO9VfHXjJuECbiPYiW0AERWPpTTjZAUPMwZ
9m6VaLnARxdntALnsTYNX7UcEU+8aiGbIpLpWQdnkWwSvJUUCN2tuPnVzF8nbuie
guDa2H1YJlG+lunMJnwz2OALVW86nuslsi5NJlZ0ewn3C+LsO3pXQN+Xgsa85AqS
VcwGcwzxXw5lO8/J2FwQvQku7YVokvT2y0V1CZbOM0Ol3elGs3qBnBtpOQvg8rSU
p1AmO2PY+9++lnuOcWjcFxJ92hOBZ4Rlac2MQ/vr2Vg8EKcCm/Pwz7Yziezb9Lxj
aC9VAl68CzwNHP4aIfjOUShfjxr9ZowTxPFWYr78KoPzFa5y0Lx8jKv5owYFTKdp
rPxs2se5BeprcTr28nnPvm7v0lazfb11YsKdGTHlABFFemSHy0VGfJcHB5M0G6/A
mzKQfE8GPy/gkVjj1QqUsi8AJUMSIwaLI8e5D0rp1Qs6Qb6KAk12ZW3ur4B7GY+M
amR6QmDEMu7h6KJoDpJQ0IBxHAvMdKQ1U1iWyN3TQdxu2LJgm7wqNJIGOI7cFQtu
G+QZEdAajLiNhaApx6SMqa8GuAfJncCapCThqA55kA+Y4+8GcOuDEoS40VzuFjA+
PcW73cWXvSNtH19SoQf4SFy/2BEzTT4UXpdoKx+vyH9e6yd5ftVKRi3H1anEfAC4
p5PngVNOlYOakxUGF7zG1g7NjcE2MhoGH8WErp2knF2+5YliF95NyyB0UVGhjvaA
0YXBjRhu/byydLo/BnBMhY13qOQ+UVKcxs+MELDKFrpbkIKPgYbZ/iTvj081i/91
QRNYi+g7TIbNVbtRZcRGccFkRaYHI7AGML9WesiELRfcd2uO4qt7LUKz003BuS1C
0zf+av07p4jw+psEzS77A3ZeMhLwCwX2rw5xjikhacyAFIMg0xTBO5WDhFei5B7Z
uxWmvczxNeRZbOJ0xxLu3HHPk8KXjinH28QvxJr1sI+YyuEjLB4tdgROikcj0VxJ
UsPLa3aHumLLfKr3+mtMX+7+CVzwd31dmBw06hkeCnok+S5cp/eHwT9QfVtOo7ch
NCa1WhZHGSiadp8Vtz5tia1mbZcaxVqbR4+bo0Sy0p4PTweM1niF/AxW1vO1nYOB
0wkuFgcuD5rRzswbphtqcMBXly2+1VlEwTOGkiTwLONJig81cdrXows4nUEIFg2A
+QLpjPXUwWgPDPfefMjPM+oEKLRNXk8Mxi1vuGdNA359FEcWjDQ50b9OxmThOFvy
l/IPnzOQ9+w9sYjy3KI3V8O72xm7ImLwFXpwdc4cw2o16jGQEmCpGXYA3bgTyvWd
6SGP9Red6TaKBGuwrfpQTBz1JtYwjF0SC90H5USZv4bPFClKmPK1Sqt9XsYzVUFS
WIGP/1RBi4MG0pYGKtcKJSwGlxttHt57LBBpA1FVWm/DZq/R/LOEsKeU5fv89BUU
KrGMWiJbxXPnP/nC8qHiVRgsrVEvOzkUuCna5NpPEeTyZXejej3fPDRs7bkCzYV3
7ZE8tM0Rka5BqyJsCmBBUxN81gMQSpY7dOAT2Ke0s8fV2shftqnZGQUXNolvB6Vk
Ss7WHWuOJH/tDuYO7c8sK0OfmKtrgV95TvGFhn71ESfE+31kRKgqCxPpEI6pyRkQ
lrmGA61yqm+BoDSc1KCe3XjEOUB6/bnXZGiHoeaFPPMpng/7wRy3plC7tSR7Gzd3
2tZm+Eyj7A2E98WudLRiaeZzuNrl68wlTBlflhSDuW0E1SOOK7q/9JSq8deLGjA4
VO6OiCQc47iaLsap/jJqrFbTy1mz004x1mJ+ABgZA2O9RppYzwCb5Bn/iPfov4DQ
xCSTXJfzh5zfkUBf4dQn8XIUVB8frPtQHUix/KfT+zqgxy+h27KNeBRpNQAvjPwe
thQd8EZ41fAt+0QEValhVadB1MiXS6A8eDYZHHEtGWlSSiDgnPbstWCVNz4xw0vi
ZHwOqi+6Udtk6iijc2FrAFi+lqLaavJCgmyXQId0+9JA3zU/1oygKDnpD2Fjdf/l
6G/G9Ls6N9BbM6d+xdoYE2Qqeiylh+BCzv/i+s5CL6qPtG9xjf5YVIVBw+2Z+H4t
l28dJtG1PS6lIMl5TXWeXtAbwmEsRdQ5vpixPynIHA0IGfmr76r2zPmITJeyJc11
Us4YLUmX8k9kfXqcb4av8vnxA9C0xRvgKqc2zKP7ld27t3DIjNADJ3hOnfL19nKU
MwT9hrpNUGRrkJLOatz2nUrSQ94R3EGF//+jdWYhpbkVxlGsjhZlEHyI37TF5qn9
1nWv6RYkUH+lqAGn9j/HWDW5fwkJCCzGbhU78YpKPiEtsqF1UDDhvBKZKWvyAqq8
hpc+4h1B0UWvT7KIpfjlZXRJVpQKipaYvD6O80OG04bmJFVUzTnIoRNcs+JCYZAZ
PDvK5KFV9PrHSeNebc38iWVo18gMS4XEVsmz3HEFZUsvuy1fuP5EwAaT6mtMrQTM
ZwTI21Pa4opa6DiHsXoabBgTq5+TfzTyama1Bit7q3jmpRndFfwtF7R6vu4PBCqg
sm9v8OPHaEdQ5+geR/2I/H6RmBlIfYpd5+mpj+PKlJSvBUpyIO2esq///XFzegiE
+SmBj/64TpJhnZRWTeVGwU9ScpgSknRQONuQunVjkOUI7Br/2T+EpiFNKy4N91fK
KaYw0facmf0nOp7hLWhC60GKW5ltjC5sdiFhH7TlUXbP1Wehbgr/Njp6NLNxiMvb
AM1JYiCnFW02fQWWhGSOVOcXjk1G6BC1VIDpygtK1DuPuALViD2Tr/uim/S2RJQj
znHQhDH01tmwbjBsmZBHdDntRWqPxuH/3Z8Em1spCVz42tDtzZDI7Eam2NgBnd7Y
rTkGpCXNaMN61wg5xeNJJxW5qlKdBxNNawCoOYR1ogoJPtILO9sNzd2u2bkQJ9aD
ZVAb4rwTYCTwvrrMBzbPlShvOlVtRxWtldzlvrUdWzmc18WKk5y7R7qx10jOkIyY
FbPrJpi2NqM7BQ/yl5pPUuwzUCUvSMsnmniE5kQC1igVSAh0qFKt4VDSoeVhvLUd
djvnGYKK6ADwswFOEn9HyqYAu+JA24B8aqhhu31XYD6rQCSRHOMcrIfCjwHBRsLW
cYLcQ7rkXj4fTSIbsYO5upjmQEYnLAsGP2lxGc5Tz8pkgLRyOqD/DN0CO+U4YQwO
PzmABbabh9d9aBDEN8ptqLHrwiq6H8vng2uwORm8dJN8PRfz5oSkvt1GHHDCBCpK
1p0yTngyZKVwXOPG4+K+g+3QKeDjcOtNx5xgBlRjJi8u6yG6rmltaSkzUKVq4Jb1
fQ4R1R6T1eRhgMTzayPAX8qtm6m3X0wqbb8JFfnFb7qA6D6QXTUdv/JEyugfNXnV
Gr56qrRiKPc7HfBsMbSmepbNRl5FV8EKHMfTg93xjIWF/J4Qgzkp9dT+WJj35h1x
GwqCAz9OoMttAPRmuTXsiR66kUvVtLVrQPokb+b6heCHQ0uW+BFU6fdRA1p9khpv
bj7KiqKcmAXF10rGBUvWPGyajK1diTw0YsVf77Fy762fcUE/a0FBXWxu1qaFoqU8
keu1D65sDh6lpBdjW3ulbHucLeg7Jd36oZC7ndXtKukewNa/LDayGkiHg1Nt33tK
COyhP0pHxHbXhJPB2w4juiM/lpB8TscyeJUM+WkIYoFylhXlhqmroRxv5ZTqwfJW
IbrC+qSkXP5xJfAKTz2abv/OzqKBDdYS0HwRBwaB5j0QQ3CvxrtsRjTz5f4h1m+V
MOD3nEDU4JD4JrXyv6qF4bV8MrwT0wq0DmNn9jsjOpELoCxFx0VLKRmPcdTTGpt5
xbGfIeNfcEVEt8DC731tybSsPtWQnJWV463YLnBQ6FZ9pFAp8ShOO3OHVzbhome6
djZyA/OPFbe9n2kiHnMe1pZdKk71ZqHDH+FUvLV2P2wifpj5ZzL+Z9LlbxLHYitn
Zjc/3DAZ5b83qz3dAcLq/RGqM6awEerRFz/r/R8uwr1DLEq9GWRo8D6FKfI58pxC
q2C2IWPrvSMnZ8+0IcUut9pnYjSCXl0bRQNAUkv6F5zXktryMUfkm+Ya9ZsZSghj
QAqE7gKquieCBsICqOtkecoEjNHuKTn0TCknhPcMJhkKosWnungz+cudLhohDB2z
WDQeU0R1zUVhFp3+tFKPl9bnDhjSkbKO0ZhzsrI79PTWvStbFhf6a6XFGTsnmBOz
uSLI0KPycg/ndcV9Q2oNpaXcG/DrCai4huH3LndoYDvP1kJTGU7fsGM+loEj/yZg
1bWXt4EAOE5vJpugxxqZPUoKXuEogbttJ/BRUUK1bUer8g2D5mm5jCkI82Rvetln
hjNp5fD9Qar+3N8HRHcCNaTak0nND86pyFTls9QKJdDodh7b5hbpQVsYu9Woi2gp
vUEBnJLZzSO1EgPUJU6KrtbqAbh6dtmV7MpWqSXl6fT+jo9oH9gPgWe+q1HZvWxn
hRoVZP7knacpDlyLdLrfEtyo9KBFbBNkI2wmnDrOm0t8RseY06hn5p2cwNJtFfnR
plOBcIjbhMOHMQGNkUNTYMeHSPeE8OVq56dcS6RYfDGu5vui3fyuomhfWCmPt+P+
yMqFGFzCQA14OB+4j3czbVWn6kOtP/5dlirpvZQabC0rIs5RhFKiXwiqny45J+RS
hIzxGAP3XSNIENkMXD33/ZrRbiPD4OA2ym1B7xAc0zqpSCkEJXkP50b5n8zRKRN4
Xah3o8ApqPhKBa/f3utvP5MjK+8dUdW3RDpt31WpMmttO+HHCOx30pMCh5Kox0FS
dJARdjYdDHF2aqH8XHSkCdv+pTA8GfNuSivFj6Mawgk8d0W9A5tiZXIzlNEcRQfx
Yqt9ypGIBCCOTKh3vR5uqzztl71b8qHSR36RNhOPpsDTSCRy9d6sgaoGY7AibGcG
dp0jnDo2b7t+Yshga3oICt/p27FKjedZ36t1M59TKtgFYxL5ALJCzgKibVzL75is
8IuQCQUCKgCWIu2Jqtjq8I1BNIYHUYrlucUxI/S23yfo10IAfqfDJNuuNzkB3Mu6
89GLsBdNpE+RDk20i/qA3psecnFO7cQRfcgtiuBb5J2tn1X7doczQ9mgzG5f+wJV
faK5xlCZ7eOESxUVSa2ytNc+pehHnwG3FFylgOVvsGXe8eJNjq1BXNX1ctPpJLL7
Nj4BV7G0geDe+Mbd1QU+b2PHJP6GpNnl/D1jv/jxkdbGlTkKoPYmvFPEe0I6nyaJ
OGKWL96uvwPeYMKFkD3uI9dESjstOkKz3yytwBpg2G6cEpQqm6ZiMppWeA80hSvR
MphPRgZPVkzb4u8Krpqu4JH4dNPSeuPKB+XAZPNXGFedsuX7p2AY3O8lDh+55ksc
awTmbJEBPfS6MKrr6j6A7ob2+HZwg6YD6FRnYrOhmtkQkH6ouUQP5K0LRrz1fA/y
poOFCYMb2Iu5nzmF4O/oP04w53Nd59lIOWGf/JKhtWyx8MlC/bZeeyBcu2+8G/e6
GtbtuBEHi3OlVX5hrvl7sWaugEd0HZ4rEKXVwQyO6dWFJIVmlZLMJ4vH9Xp2+vSs
4rUEu/xLHklOijeN6tO+ZdpMTK34pPaz6SGcDDd3QWykg2sPLF5WE92Tojijy6jj
2Kzbva2NEF7jI+JirvrpHYFDhozZ2rB8O5QbdyxFhZon5Mw9ZuH9vg9NvUdyRXv0
YSEC8lZEVFD+Vpt4uOjFRdYzkM7souGyfZREiLHh7qWSZaNcvnzt34srCRzriBFa
NVI35aLPEMNyBRN46jiwGN0t+96cnbVya6e6WzDBIm0tGAoJOEQJXuuJJo9FEUFr
hKpjHsKCykPHVSpPf7Y1PDjgTxUZ0M/ICijqjtFOe1Q9pEe1jOb1GpFjO2NyMfLC
YCIVeibVC4o35U54pYYP1TabcXEVr2cGi8Oere5ZoU7V1yNcODA82ZtbUrvyzPLf
GHEYIPdKkVVJmZQgwsB18GjTUVnyIBpi2+WHjbBunR0/7dffsjrcELrZYiCTsCpC
3myIpvlVNU8e4LiZClSV+WITzLXb6SE8McYeNE8fJJ1IhyhqLR0bPWn0Vn9KxOHH
xXsGzEYk9wUH8FUDhT5rXzGGmocQ3Q6+xQlkDXGv45hjidpExI/R0x5/5LiyPaHg
7XXROK3EnQgyqXkZ4XxOyHvtjHN2499OdEURPSEJv8OTk3LkTSgsg0v6k1uNgoYp
w3B30kCPRn1AVRVQ5B0d6le07F5Mi2c5+P0JOnEvC6IyZaNLJzStNZjr6CJ9CNG0
rf9T/UNOeGFGdQNmfHjz4GFTYWq4/aRchOnufriRle10SGm6CKoNfPRSOGPNt/cg
gnA3HafYTazojPttoCxOubAIW8Pd/hh/4mJIUJ/0LjnS2dkc3eLR2RK/WS0f7OTa
eqyXBjgimULjE7DumGDUJwUrj4kfF9sccN5mWY+bEDSdz0vvGSCTxd1W1vxQ+9hI
iNpcmwKvK5UIYJ9+RrKwHVEF42MoKV0SnGTeYDt2tPMVe7MTls0rrUj8y+IKhVmT
0gvh7p2wnMIZ1diquA8703co7slkGRkCaI38tq8/jLtHp1gfiUHQNouRqOzDUSV3
wmQilf7AfS+/Z9BRqhL8MaUfjhT2H/eIHJdF2EUQ4Q+Js4Lp7689SGiiD40wT91o
Stx+cX64+pmQe5S/EhgBs/NN9jNRxz0Wulcj5Ht2PMz8Q/AB2V6eumIxKPkXrcih
Nx4KPadbGs8VIQCY3u4stJIY6PIGm8wUO86CHghXm8eQ5KYLa6bEHjSEFkPP3d8D
kbM/Dsru088UfbBF6sqsh3g1+GPczeRPAJbHit2fzXS5XBeslkd0eUfWtkxg8HoI
8bI6KHbz6OOevTaizMsnwiSTOo1hWFElH7mLat5aYWP4h1RPsAti8qYkB0EFjE+u
cSUyDNXI2LTbnTKTcW0d4ikZL1cMTbiyzYptpeyPAy/xsXgqn0i3G12cWPHiZl0r
JI6AjBtrZir7ndrIkVvCRqoDfQR3ECYdC/LMM6pCzKMyMLMu8fWGsgiRv59RWrZt
T5iONgz8bQSNgrBVDqjRjLFQNPI9kZtc5HIpPnvIfygkNip7NzeByA2t2qNkK01h
BIj/Gr3CAPt5TyfrQUJpp52n7aqwYDSboq4LMXkSH9+kd9291vFBDohrKdPta94C
ezTwjl8uYUMUxFG8aiEi30nS6/FAslZYuneJjOQ2Y8n9lYe2a8StItkCABrUkd05
HaF3vagNohvMh8wMx8bx8Jc5+Szd/3i1RYyh+SSS4RHBV4DDObRfy4GcGouRTr5X
oeLxy3y9/0t79J1jlvEwpQncAvt6/Z5s35gvyi87uF/HQc3spgEk3aZRmSkqw/XY
v3o2HzkQh8Zb+B9Vt0W79d1eEcxfZiFeic/KCneAYw1fg6rsTAETNVRBfM2iMteB
8brmmVTj9JeIMlqK0V9YuQjs4RPii7nE6izrfUzSG7f/kzrb1vNOFfZe8A8c8LIf
lpNgWilVfeJ4/7Jz/OgOu498dOik4zwcu5RE+ZVmbYJ05SFc+fJbBe4K1HOBp8C0
eOCWT37E1nYWHbpSRRWJdxqsUDo/iRbChSItuF6DMzfPdBE+qDyjCVfPe2UPgvjD
aAlamFwPCkTVW2GxiulXRCUVZHzY3Z6d1ocU2JbxKSL/YYyI8NQLTWVG2ecdtI6G
s1/7coCqDHbHODZwC3f8Ph2hGrJKaVCwqOCndAt0th75tOl1awhKcK3MMdbIxy/w
Bzp1pivZUlQ2RNwAFblqZkepZwnDhzbSynO/c5eTfW54H8b/7cMpr4Plq0j9ZSzn
ma9NX/rYGwaDzwvZqdgSqjto/36QOCL1CwO4umHul/KniulbLi8BY62GOob4a222
ZxRDQD/csX1nrmqHePiLtF7Ul6HU7dpm7IWIQGMFotFb0ghiadEMqBlAuEiMAra5
655V6OzNtpXujWZMQ4P8OQV/SdG/2MNKgtBH//1/ikiQBWH0WYzljw+B4s0+F+We
1Ooet3THhAq7xj0Ss+PWSt/BWbcnxGc9+jOBKpV33y/37IBNn7y9Y/XybAaGi35W
1SkUWOMhLnOE/iiyFaUYxM9m1/6+/S0uDM3k7WiVI8teihnYcBLzYKGq6ZDDRfQu
0eLGZN7NRgFer2KQtfGSfkYlEwPDW7j0EupH227VIhhnjGkomJNcQNW7yNvtjbS7
OzWPMcTSWrMYSCw1Zs84w9zGzpsVJuv0j1jVl0u9iTLVzO6nFMNIMkVCRM1pMV+b
15SmGdWnjyW8WM2Y0gr3PKSoDl4zAslAuHyf2V3+i12/3KHEve7JlRmQfUOlq2d2
6tsCkzI/sohtAt09IMuKLlP3tR7QYdkv+NOyDdRpsetAl/nvhXUvGqeuDHOXxv1r
ZQ68gv+sNaghDjz4aKR+8Kht/d7Jz8MSqByOE78yA0xr33KyYqi/3odADeGzWUSG
IyU09JUywp1Yui2Bh7crB+GKLKFMyGzKwzcTYZSUeaD02kybpTXmbTgeVJSoeueV
faDZAtRfRtP+19wNfWFyOZj50tL8cvcQ5J7UClbUfmatXLAwgG1bcY8kAXOasBC9
VpHNShFUR6pDnJqaWEK/Z4aaU6ukqv0g+Llc1B4REEIpYLDlQhw8Eti8bZHVGRme
kftrVv86WnDhbO8fUMmW4CW4ZuBYKRC8OIIwvjO+L/EV58RBK/ckAeTtzrrsOMlZ
QbdhCLvZk+ZkezF+Wzerx0eIZ3N7cMQep+gQlV/OY4eODyUnVYELvAoZ5r56Klas
b1RDrsBZsvnPwPyTU5uPTG7Fo5tHYIBBz/63ObhXH+iP0XdYk+ArZZH0u5zTOlHP
UJvWoxPZNUX9mAsxojcWdFU5rGFHYHTxTRHVpHY7xwHZZK+7q2cPzoUp1+BM0QvU
xActFyJ6YqwfMgeGYp2NVVbtgPi//mVtiNUWgT9x4ajiaw/kUwd+2CiPHeJV2FUu
vdBIBYPp400UNzoatEFE0ZyUppxaPPP6T5Ylm8tHt8MptQi7ObGGoNFHEz/Fftp6
hi2X84wRok5zkMgvhztMCnlCLC4YZ7KoJEZMfylfKuVeP6gafL3n+3sfCUxIwsn7
RXDl2zfzAVZz5yeRGI9eypVzvqXwCfVbg0f5p94PfKEsi5MLNtwDMiyGWRCpQjDJ
li/NygRBEuyja8Z7vobyCZZvGqsFoUVsvCHZhBWly8rmTtlTenED1G8i4FycriIM
pfZmOehU9+sbB/C8le8GHd6fbImI4yrRRaYzKSDiyeRvcMnn9406hRZQfBzheTPK
MTm9KjCDxrTfzyR+jiAetcQvS/s0J3L9Jg0npTH6duvBTehPaR9P4tdqOAI+aAo4
1JLcLIcdTM827XKpczbEFEZfdOpCsND5hmrXpyimBiR8oXxt5u/BiE+akqHhDTxe
7XxFNpcD/ZfsdRxHzF81AU9dfpkj4W8AMEA+YaM0Nm7CXHBfDAK4cwA4hQ5z7zU4
59ef4N64WmlCiKAwgNUG1/L0Sei7N0rk0A67F7P7jwuM21/JnI280+Uh5aOW3g9S
QvKGl+Mek7emDXNwm0eD5A7XAf5d0om+bwQvrdHmSySmxU7PmlTlPbkzQP2iQL1S
WuqpCpMos4R2BF9vwt5CPUrPDGnTT1SGSt8QP5O0myVrSY3eu/r8dfSiHuVtKUfk
e4MqBzjHeggDbQwoHxGlxl78/czIZ8KVe4LMMIoh2ulfWc9KDTdjQPfrI7VSX9QL
r8F6gSIeWs4HRZ28fox/SuLHTWGg17G3psNASs8y87SMkvc3rsjoXf8vu56j+c20
YjbZUStgS39ehazR9eIvjbmGRkw+08Hc3QvFfna9WB3oVMswFNNHgX+qq0d/KnR4
qisFbRaFaP+ESBZ58MuT2PswG4xP8U9XHxCnpYQgArE0EcnH8U2AavIHG9u+iAPw
GjYaeenQazTPC4M/i0Mq7EUHTagrlxhe/+yQjXlIGBGxKXQdLq0MHtsWHsBtRaJO
ipZUxIaO7S9krlcUq/zcN8iM1AZNAbieavbaYgeJTOJYG1mZGFJsxOJJ5ABlL02l
KMAtMa4CgptinQ/9zrZz6EhQc6f2i0S5xT3DpSk/jutDvOS61u8M6NJI2e7gCIO0
qTYN6X0rMqAjkJ4fq+7RQ956jpCeJ4LYoRDhO6LBtO3cStOrDSQ6jvM+qx/ieI9P
6+ZRtvDwe82WHjs61oZQZP1aN1A9g155A2/H0bQBGEy19o2gRVzWRNxMRRD0NCbB
GrnLkr68f4NE+5zrn7dI7/1LGlPDHm2HgJaTEEG2dO+vEoQw7W5fE8GBCigmaQ3z
zFrUp+N56lCQOpMebBMQ4UI5CqC4cEvgiL8S2D7oyy+gidrDDLwhm8nfxoo4EEVD
GGYumYFVHfHC5/YADZFCHP+OSo9fjAxdSjjUA6EH3UamV8kg9ASYLZwEr+RkgG2a
QLQLTWmkbMqa/1SWwMdVHKwOv0WlG3gxdmBDflh43HPkwaCDAzqu18/NxcuWQcpe
hRUFZ/vUJjGxXvEc/Zpu+kOSRub5aMsowu4rS/BSRru/W/MON0KYT1eGl4WIoA0J
EAg3sJuhjVQ4vHSqyQqChgRh3Rf4nhSzamJqYrB+DS9wVLjGgOHCPGs1VQvPjO7w
bpgJrfbDTD77ii8fauYuilkt3xphFUck0yKk6nJvr+CavsdfPnxiso9omWlZNZBO
wqcf3WxYlbpIKBiaZeMNUFaLhfwxKlc723dWdzTB5dI9j4+2hAIgTYSBiFlYBlvW
EUDkZhE7cfbonBLsMNJ2fSg1k/AVqPfURXZYT1cOMbhdwPRXqMqHmDAawooBoxQp
2jjvCvYKQfayh2O7eHgaksr8Hqlee0WBL9VLoIA1/aG40jXEEdIHmQAK2wTKjAPT
bNzDE6uIcHe4o6qPQwDSb+O/f6kcebQlLmmSG+QYr86q0o4VPnKPgtfzF6JjE0wZ
YQj74szppaSuyFwitvvgUARIl+1Hhn1Upi7dW33pMltGpkypINSwCDULUGPmhkGw
EB1S/qLMKVswEOkD/ia3vjhF2cVzFcaT+7mY8FGb66e5EW6ouVDTrq2c/9Y8Mk+U
FlddgDN60kTCa214rxgNRXvNZzzPIoJP/SFTSALNSLGkygik9UFefp2B3KzZGnOP
kYrmL++TlS+b1TKcgZaKTby8ZzrwyyQJb4yvrASIvr9pz4kFeG41zgIlZ6D2oGnp
7AqrwHDpW2lq8pC3EoseZzlrkqCvhzyFt6sCmar9IC1s99CNc2/4lanHI/0i4M2r
SlzLvzVNw8boExgNRutM3FW09PYNtFQnOcKdOPWcna2kFxfx5SDaUGXUjd3IVntd
Cg+8vSnm5bSYtDGhB4rfXGjZNhrlWkAHO8cCxQkcbdrIZ39XNAutrR1/TtRfFTA4
wYE1o4rnmvlINPFcC0ExCMYkMGNuB1P2N8tYHuRmikW96/8w/I8dlNFJ7U2thSoy
EICD4KUdd25S3Tv50lj1uqbxcrgeiTFSMrGBxD21C5rt0pPD9txdZFJbNcts1WgM
MXd4QNVXN0UQXjL6R5BNb2FUktoDJLhJtirCSjdMCf3LmcFvtik8TwUEK9yviAoK
C0WMv5EjW0heS37UkSlKNzuSltHtzYrqm7kiz6fY1z5cOFbgh3nSvhcSauxNGmPE
2zSkSqoCRBy9PWczqglM6/sJUJAOnwcOirs4I31XKCksYhbvEvO4mhIAYO0INudO
Nb4lLBFwkaLLMbkB/xnO8BJi5R2uYYYbXOvZjQClTt6nU2+m62S2InBaGWhC8f+w
aD1lqmFKZ/edbSLlaUyikk3nsJ4C5GGRpguc1bRKid+Qi1gmVqA8nrxqyYfd7kpn
7u2LLYZUI/YyFjPTlZMHdxZQ9rSr70xbqNv0gd1bwtpS5Lpd2iaq5vbs0m7qinCp
lENNIj5i3kb87BJngKpjoMejqXfYCZzEAmcnd3j7dcnMfVfZaNjcSCUzXHXsxMl9
DVg+McCfo1dXypZ2nGugQ77aq8PlTpqGjYAmJ98mNWOJF7w90HSnUUHUTPexI7Ol
EhO6rgnFZ7FFVNbSIaclLSie81hahgthnmIeI+ducfBF6FjBzB3472Ux1rN+jH5P
6beElqL9etJLWqXrbZPf8RZ5Gn4FeKEYBfPjk7GZDGJCHK7ugdy4Jp/0lEFaUGQN
YpjtSl9TQvDSSFb2U2ycdMd9F3JLhZngw+qViuKnyP2ipcr3wRXVdoCmW4s8Lq2A
FIE3aWdwbp6CLbZml7Sy0weVAdNSM7v/6zt1lHrGz4gqSfw8yRbtTRQQsBcKxbPd
Rx4T7TG6og5GDRl1n4gt1/xquQI9WeQ4h0y8Y9HwK4baVtXko0B126BE65eDHgYi
MadLdlCGvX243SkAde8tn03Wl7NvNUejFfhdc/oQs2PkT7jWN8zu5L3gQd3Yvtrx
Kbej6rEmKwLS/WbliLq04vIy7byTT+W1aM9Wyr1IAw1rzYSHm3p8K/EK25OUjPkw
rC7uMJk85uDHe5Qg4kPGxuZ65vFD6RhH8xYjzam0laPzOYQiyRhdp2Y6ISlDmhQC
kzxcb546B+6nRB1bQoaM3GGuVLF9MopD3JCZbWmDnxrJO6Z0dX1BJN0Fr8IDLCBC
V55+tb004ikF8+DC9qVZWZCe+mI1wKYn3AYWW54gExuqclTLSZN8KFG98RyzXjR1
bm0uq3eg7wvctZ+fu4mtnuJ7OGl636OwDIY63HQQAMtkyMop6RVkRAa/uKeoQ8W6
rK7xTnkHXyfem69YwDcXDLfPQpg7K3IN40Uf747fAq5gDUtIUveFz+vTKU2w4fH7
qTptVXvn8RYJerz6tpoH/rGfC6ZgeSSofad0j8FLKIkGLxc8xRAQk88mOLL+6YvO
jEvet+gdSwuT4HZx553YGG9AjQTz89ZzwlN5c9pc/GODfJO9B1R/Ug+JoL5txz0C
bVAZiwtsk4bPNgsSqXm+T2V9RV8lAKNbQevL0BaQi/yzERurghigwn9vfMafOviJ
TNzSW5P2wLuXi1vNMineCrdVuEXj85pyj1dGWOz6rdgfUVziWHdk6HBYyZOb5VGq
se3LuUHILQoC4ivTYeVB12t8LNwghf6my60EFo72G6bXlqHQe0FpobvUpUyJ9un3
ycgICl1ZqplgINmfI9Bf9Yv6uLu29No2AFQzLZwH1kTV9CpVuxL0/0t5xSuxZu6Q
DkePSbOZvKz1kmc55yKAyEswN06AU/FAbgBrFmhWqrHdOCJPQ8ZJebZc0z0o+Oig
H63AevxjLrzPFb7X5leMKgHO1hoUQxNDCKYAaxRIVrt3Rl2NRGd6x4AWKujaXV4W
voF6xwimRKk5rWkB0a9RcYqPssaq6vEesJPyjAGt5QZzcUbGqQQdo5P7Bt3v3Nns
pJzbvUCkYlfjGAiQ98iDkqshrXfZ3ArSMJOl0j1QtmfAvu2Rh9/1uVTE+91zqcb1
pfPTu4+diqHERdfYte+ATAuOI69MG1qn4JOu75ufdov5Kiuud+FmqIsZ/U/o7MQd
a4sldS7DJzY4U5iDIr4Y+H7FLNyrfciX+DFe2RLrTED7qyIOnK/kAMwUY+A3gEEn
HKBBa15nZ5GqiqzrxWcubhbtolHrY6NzT2GtKn0Rq5KDCL9ccPT5VB+zPDmYMfZL
KQ5dXOmPfmLavR3Y6GLP3IebCmXgspuxOi6kwguaCY8Zkwcb32J7LaCzBkpkUu8L
dlnkqEWwedBBpjB2RpIttvHt8MO4xQNiTI3datRWkSH37qD0QXJLfm+W+LRup4eH
qXlIzJZ+C+E85WWlMFb2RsNc6p40vQoThCQiSrgwr8RouOkv2YdDmAvR/Ee9nPWR
D1A6QQ/vH/lNfDcC6OoS+jPIkjkRkeQez5eu40r2a/KwXz8t09J1Nk6OWqLgQw26
8MXrtbJaXlNueSL4Y7cZINUmxZholdn+GZAtH50eUqTIL2QGA90l7mZrmBbvZTbS
mQeNRNY/Zqgtytfu5KnWa1BpfqTQ4zPJE34w1zf1at86yzI+oD0Rnp0qcX6jzLXm
NuB7YcYrJnkuAgvOhzM10BETmoHlHOxy3/ny9RuyQoKqA+4WpE8ZFYdSIWusimNY
huYtZudViNBTkYkB1p3bvg/E16s0kvNDnSG23Hb9OSkyqpbfwadcg2ZeOPeQDL+Q
ONfvdbmQ8JmpWt5CezbcySc7DVCoLbMOhwcU9XXhXLgXzUKqQ1R2C1wEzH+ryAdL
If3SdcxqaKH8cxaqri79GpL3hOWBHOy/DcrjTQRWpxzjE3k+S1MJ/reioC41ByQ6
kkJlsd0prII1loqf7DZyz7cYKbf/i8Njbqw8n3uVKpgLm9q9RSP/3grt4hPrxA77
Sa99IKJQ5+WuRQolWG2wMrEZDKRcwUre6iR+WJpYUAn3rhHf0QYypqo688/2pTi+
N7opRvnYg35JEIANkHRe1G6JaGBz7a4u8sfNsjK7iZQxK+YekkOx5bnTR4DyH5QZ
87lOmaFBGwqgfOK+aSg/xfupEvgaj8i1B5sFwqUx9bDdQO6D5c+w+QLpbPr63pOa
/Cq402mODKJ2FtnLdBrYrRvYcMzUA/blBq183PygSbOPFQEHwL5cSM9mT3w1V6fI
7AWWvPGdXPNQ5KSytQD/dsdUwWk9NemQzLKJf7GNk2IisBOJ0yd8qFSpXrHVRo/Y
6afP5A0fNBXpDz3UoXlXYMWzatVPHVZ659F5aFP2LXoQPNwM/B0lUeag/XoP2Mn2
WmvXteSHaWcYrsSYEsslMiDwPKzioGiT3H4rorlZYrudbt4HUojSbZTjP0Vnr4QR
lDQrvlXLN84/XqQiYvtEMG1lv1KQzrgWYWvTKlpW7LJVqsZLiZMXxj64PD5y2cwQ
p/lvAPVthIm/uSSBkvavl892OT0rLZEDtyIzkbG6CmqCLLQHbGWK6uv37HObp5j3
KAd1VT7REWOlzZ7dLsQ8A2d1QF83KSo8o3pBcv0MmFrMUmHPcBSBg7D0a18UBS56
4OmpTmL0GklQYJ/0k046PcdCkU/R/Me88r9S3QLS5WD0x4hkhfAsTO1PbhSmwrJb
uqFdzNPoIs0ZkownV8IwlHHcyhh3pA4mociMkC9e3wXhJiu8/q53vssv0xngzQaP
npsQLbHoKlxglmfsUXp/0DehW/Ko/UckiI5be+FBVvgwdOkEz3STjPplGcS4oU41
XquU009IKE6TIPLogggqfddTk8hFh3zuMkQoZSDiRAcdK3XWfGxM7AyrAhe36Ut/
usfDzrA2j3McKL8qSojxJl8we+fIs6fxwJfr2Nzc+Xb8OmoTYJSqrAZLmmimzYpe
lL/I+b26CB/20Husv1WkzQqcXsLY9VL3QWR+T0lXjxTDcGJnB0rIH4pBkuXwUK4g
ov5lZi97rn7/qGGX84oxJqXBI3ABX77Wd+ITaFJ8rBn4mubtTrqPTLSbxAwvCXD4
3EpCBnKTSXG5UugxJUJkuq8hd+Ro/3X9NDWOtuiGMzXEnS0ltlKMpolKyJ/Mbz1S
NjYsMO8LIiV1h/iZKwcwQhHtNZNaE7d748z4+91iOqK/UpcVuLkM9d7I8aeUW54B
caTwnohBn64R8aKqXn+3/T5nVy3pWGJbnZDOKDQYVALLJ5GITj61EaX4rFU+OMO5
ub5lklUvr4MEfgqRfdc4RaxyVImhoBzQjZjDsmxTR20QEHzoW79yRlPLkLK1zYqH
bp8sWHEf09AseeMqj70FYJsOx3X8bPavq5ymDcQ87aLQaxD+D7i/5PHwDA8PK1ei
1Sy9r1YFnDj72uTzk9ofavWqC6M1BmD6tuCZzjZ22Gr7S6TlombfOo+4F12Fk/eT
4VteIZGm82iNs+cTe2Q9dnIWqQizXThDFJ/u90U1ayg2z/dHQbCM6oMMOEL88mG3
9XEXvsx3O6FleXCE2dMTs4VVDd7NvUj4fJFItX5/HdkbMuOa8Lck5kTRSKXCsiNA
5BbSlGDZMC74Sxl/FGsxxurhR0gu0AOujoxavhT8p+Dlo1ld548QT43DtRhKKNr0
/49mz1ejbPViMR5UVnfbVLWC5hRt836qy1eMs2oNW8kwX5W9O59YOpp/70a0CbXV
Yk8D205HK+k0zj0W4F65IxvCfn6O4yJ3v1dR48xMcVLZiWR/jsj9wVDCz0YdcWKJ
xQuWSYXwR0iGP9OwFXZuzJ9oVcPvE8PF0NEiCyQsemENjh88Ggwbeyf3mH+M6rrm
dsJIRnYNkvuhlTJ88Dh//HR1XY+O/tsfgC0Zan2eUJEkxTIrGkMEJEzflDOi3SnU
8yAlgljMn/ND9gagYTRsEzvTO0tCDK9FD3EzJANtfh7D6wyN37Pd7KUxTCiFop3C
x37Vf7dQQ8b8fsJm3kd0jVKadLoVSVKpIhL/fczFA7WLdhIK3yORxQJXWfVFvaev
6qXatvkKZCk5T7R+E6MvjVkkdLQJZ17u1Ugu0zFqBpQJJHBE48tW1TPwvPXERdua
uu1Jd5YxaIEVYbyYdpb6mlmYdBIPDfcpDRXEzPdz7LFqAqvPETE6QkWnqZ++mbyI
ouJTaJScn97fCMsDdi4q36r6UUCXJRpDgYb2uEnE8V5UplX5yP/yzcmqE0fqT+1J
JXrZbURlSMHIOzP2OeJnO7lX8RHqBKzCcFKrrJZBsarl36ImmIfsyVj2pPyDHQuV
NvBPjxYKEuOg7zEznuzCM/gcU0dS2FCasociM5jZeOsoLPFk5DY9nzGTcwWuIK0q
j4jD8V/0js34Y9q841OLpe7+pUnwDL10thr7F71J5WB4LHT+73aGFuHMf5HJ3RVb
Xm+dNt/ysGA9i0DGQQVjYLWSyOaK2BjWSVzh6YXh7aNDqma5pLUwTfmeNh0icrHb
TCT2LOG4VnhEEWF49KSNd8AEtp/rNo6Z+yPaQoFr5EOfcXG6VhIOe46u+VCFFDw6
+XSQMK1xiudiF87G4TOMo/BkP8o0itOLsoLT/sDYjiJr4qDhp0rwDiVhqqumwMLR
irDk7rTkzJI1peEAAQNvd7oSKdUeSEFXOpxpAOh9aAF8xfg73569v1gLi5woizJv
spCdzmogmhRFE3rvhyVzJhyEaFXy1hbDiayDBN2Kb1iU5SwpnM2v/ukhaDZSHnFv
zz0KU9ICvchzAM7+wUUm6OsEeNjF/+MuMVlUvsHtCSAgASvykpR2F/zpcOADKO7D
Gjfb0sLyoc4ZrCgl12qo5PPLtKineM6uRoUHUR0solTt0wDRUZlAAcKgH63MulJu
wdVq6WURnusTHtd+Y07UZ02B86TEdusAQfwAMr/Z4WnQg7tcFhD6KgrnwXq9gDuT
5HPTdqBSFuS87moatKD9Jj6hJX09rJIKM4yehwa4/pavNNJPDLZAZO7a0tfjkxVl
Hs16ETgX/mTRuOxidID5d3Xohd+oiZLx6NtRRhn44O5VGfcWPMfvVBkoWoecke4t
YfOQhZePbQYVoB6YtE4KklQA7I5g53rZnturmb9p6GiG+sYHnIAtuMjAVjnWa9EG
jks0qkF7gH1irqEiDVTRlHll532NAYZhYlhVqv0OnIqte5qIbbJ7iwRfS+Z9q41n
f+01S3MwFxTJbj7jGjZHXbbvt4U+0WptLiq+T60W+YtrdI7p/KDEzEUlEoRiMk4j
lNODtHsNrTbl8UyAu0jUjqtj+EOsDzlc5tUbFilVixT2MVa9xXHdLW8tDPm2niEt
DTcuXMQFu9T9fbjOKqzxAmKzj5huZkcP1xfpvEhursp/Gh8vuNx6iyo4tYyP0S/K
2j4AkmPVHtw0hYFHUciK9NvZsb7sw2HJdIMBvhSMn2MCVbnre6ACtqtQ8KUy9DJn
8EuFRwdA/94mo1TXgHFg804PfO0E2+cW+UuQ5xcNHV0ayUsOI4U6IUDrcqyl8Gx2
2ZYNusBkHdM8yfr96cPkbmviUfC82bpzBpZGOnrXQ86uMU0KInSABlSJkm6DQ+y1
f77yBnsHbov0JzJuhBcJgYY7ZEPSoFEljtJUbM/fHBV12lwXbyp10vYlRyvedFvI
FMWI+u+SVxYr/1J37UyOfx1wwUpeq7zYN73BHseK6AGaIfpzAhRTKQiLchy1Dp/j
LDtQqY4YB1qLtIkQw36vd5cBnA7hsXpByYZoeHn6tsaNYMD+ZYtrGv5wPsgMkCd8
zWDzwVpMAZtt6Se1M9DUoWDARXtf7KiefIHgr393ZPI+6B0MBxLdKg54QHfCZP0Z
rysATMn5+y2T1YX5CS7ruwjnz4Pnym460PGI81LzRvUrU8W2C1YuY4gK8vWgQIfE
4o0s5ZbuVjKirght0dzCj5bBRyeM2R1xMQHiolihK7MNYowYpI4WUV33aUI6/c5j
M58wyECeAuKbq4+2ZDdLGZgX+IXUCqta6NOQqXGc7QTHJG2hB/vXB4QgrAZix5kh
WkF7gL1/LYcEgnRJ2vD4VX9MIVwwPQOCk3KT5cbYLE0rZqAo1XPAJdXMvVHBgEKW
ovfy667z7km0W1cgy/Zrka+CGKOSCxPbU84psjxOfY8cN5IRrzzD3Pa0WosZyJsF
F/3XeZvZA3zNpEJgQxW9Ms1iFS7qOEDP2qjaEF/CbDdGp3GQ4ySrbbMcvRvQ2MbB
MBsCjSbnkw5nb8mHRspLMp+TPpHYdM+/fHw4Oi/96D2d1UMlfqyuHo315kjApDPi
Rcf6OG/ywFA0X34pwp2YeU6jIPizAPiaKU6NXU3ZT3V+obQlN/j0ThJ1kH/jplAg
oPDYaLd9U7HSAR6NwVFRzXNgdhY3gxzaJV10yG3ZdoPS4pC2EIdQbZDWo3JCUSlU
cuGGULS9bGOLyE5dHcDbVwtt5WqwRuayhidx98GhzKSDyctcUwcODqtnv6O1IETc
tKlhYPKvaEPBP7do7yaVL4KFd3LtjORl/GXmaqIkaTwKe9Vo23pVVQAIyX5saLZ4
2xnGGbeLWC9BFwduis9uTPemRNHmQmfC1puX6bVUFZED5sdmitqvHp6Y7lDfmTfk
TR/NR0xo9BolQK0rWv6KbtQ8J6n6b/iW+gHr33DUUcfEDrHVvkeDH/9H5mvFqvS+
jnaMqFBaOrpG4iHhJ1FnPjBjjLgIjFnyAr062gQ656vo1lzyDOEokEuq9DT0fD8y
huH1PUA6nLWmFyR5Gpuc+aC3z3u3Mbu/Lkf+NX22sBAHdcccsC4OoK89LbC7g2eW
M9PvXZXRU23+tWOnjS5T3va7z8LD5eJj2RL7NRYq/fGLBKIzeMKNQiCFtsZmiswj
6fP5PwjdQIZ9oEqdl9FCvLVLHmGAPrkRBiAn2CgPqwpzBUrwzIBXIGP697PVsuiy
qkYCLBKQJLD9sBCI/ZmVTw1DmMZoBkTK9PNV68i/hGvnGF2tPLZXLkjHs9JlJkr0
Zd8xIld6EUxL4Kq3NMDk5GviCikbH6uRt4HpCmeXtc5WtyhrjHcd6cDhVR/HNSiM
CQ4j0mR6beN+nShlPN1od7lRU0uBgUu5zXUxjiZ7HNQs0Ldj/xMFz1iRYRLXbYU1
kE6N4HXX6Fsi8O/y9l3xEEae+5jahTs2s/doswCQ+GOfha6Y0iTduobRlSC488eQ
Gc34J1rs3TxJAHx9+Xm71bzj57UTHlBs8kUhlG+mwLCkNW/rZ34D/3LeyQeVSk+J
HZ/nbfVySHCiYr/ReDumSFhVjJuSYi//TVjYgp2qSKPm5PwPzI4lqCMTL/5tGERu
3CUUuVRcB/jRDUl4VoxjUN13aOrxRUXGGJAGPa3KVRxGIlee0hjKxALIiX28NQCu
tO6tDPZKXHONdlvBUmmysTVqIh0IZF7I6EcwwPd4Klc4cK9XOJV0DYpbmPku9ii6
ZKezn1bVoxiIUBrO01ETIb7QlcRmep/drzF5abchXeDqr2zhUCh149Bn2vzBWj9v
o8119pXSYxfLYBKzwo0xRmWJLDpB5v583jZyORtD5lyrANOx9ayoFDUWLOZLB7Dh
QAQrfpTlZkj2RTwvR70ucLFOt0hE2dq+nSvTetWPDeJeBlij9TbC+DaB8xOFPGzf
Sl8E9QW3DAwsrRLLuUftWlN8bM9yFBY9BKi7qjriYn1toyYY2GC+k/23WvuBHmOL
YWLIS68g72Hl12IFC2C+bDP/8N9w4Zk7FvLIZLmzRAaYV64VBIZKLZhvlh165Rmw
E3x1wlXO7V1+Pgp9BkCTaYHatV17Rr5bQ3a2NB/wU2qxwAGNf1TBrYS03e6/Gmuv
g56f/xSrJhVrZKYnFqMQ/Lyu0dEV0FLTwRS4ASTf45CM/2L7skLqyv7TFlwHg5FT
vutasnRKeZ/fmsQrimHziwbCPrKRw9OmBZHWi5w3+5uWoXWKOCIPeEO5r2d/9yRm
1rsfdpDYc2y7n4nmuPTuwi7PIDhanankbsTqB+AlJfqhIhlcho0mtYRlq6HxNfAm
GzFykKanbs8tyROyyB4PGtSx0m+da0NXNdYNVkV7evp2zcJAyVI0ZN3/AHb14mTZ
xss63UEdDqbx28G6f2z0FJozQKowOAYmx8NimNlfeGeTf20lOvaO0G0OXLnw20PD
1jWnjvKAU8PYa9bG7fZVTwQ3HtgYn5452iiQjxt6pAHF3SmUebfqbe51yG0ZzCIv
s6nWB+7TRDV1iZ1cjwE5ENvMeYXq9a3UOP7gFQLRu40a3ldXVqsLqrIQjrGqrkg/
u8Z51cyLKKfCygBLSYa7yMIOERT+t1eefimpj49asgmOj45sYu0jp5XzPw1gHdL7
4NOmjXZZH4+sY/acMVYjkGGGIlsalgOAj1TYP5R2bnwxttWlYXvkN5RalRr+0ONQ
hyXmjUGXjdX4dv8Z92wryil/f2f4l8lrEXJ4TJ4VUNQNaEgzefW4HsHTa0jbW3v8
nrXDaxL5bH/ptdnsBst6jdPz9BYo9wS1zKxYaubaV4Hrn75Q52qvlJPb1G2vrq3c
PUDT4jJ98lB0ILPPB7K4tWnMc6c1/Fg5nhkPDcx4ceY2div/7IlUCS04iayO4vYh
dL98YGPLfWSgYF3X1n0HB3phfTop+dERkhBLfw/dcssjgcwVpnQCbbkWKwfzG5pc
0W/zUgnfDIZV2d9mnkhMLZod63xOEQ1KpehCs1K/7F8RtVKTFdc8EDxNVxmCAJof
5xS2OOdY7OeP01sQlvPUCC6kFhGlsDKTBsgxwB1ZCOQoPo8ex4bt824H/QoLIxT7
eV8oBpxapiOYgiw0f8X9hK6rX825LyQ6nwJ6LSHv8dCUOyTbOHItcedHeiA28gyH
/88QcJD0zX3FsjPmGMwgSH1ttFjlxHmDT4CY9db86wFYVo/uoSLGsDMTVB6n+RHv
kFIH+lcJYTNJgaYsatbm/w9PSx1gSiZDklP2x05Nk+xxBqWWC+8i3zt06+QaRvmf
61KH5ZHOaiILW7PqWsA/hfZMUhpvYmrorG2YRtjldWhBeOk0P8JCoLcryF6Jxye7
45aakTtEctLxtctAFLlkGCN0xV62w45+892QXFJxX7fWbd3RWg/ECFPhvd3wtIys
mwlE+EWcA+B6UcJ56QpDWTaoTBgG0oGQ4nyHB9sHxl6xJol8VFO2Kkbjz2c+G74Q
r6uOWraGyMMZ/ob+CP4nvYmw3tSeKXYI0XBtbiJBUW9qGOLMzZpnYiYeOkzZ5Qce
XdVAIcqw/w1OlupxkxVDKhAYy2zcwAkPin2gSqSas21/jKiuiJ1jgFqHkPEPntFJ
rSnHOwF22y12UhxHRdpzfF7mihX/GkbOdWUXEFz/iaCgiAmd+VekpkpkR1D6roV0
2FsvhgN1MYFoiyJ6K/rT/mklIPfY5vwBiypYLNFfFNF6w8H6nPZpGCJXvakaj8xR
JhmIWZ0Q4uTdXmSjliTL9LzATYqOm8m+RuCWweM8WHzMOqvsFnixDHrfBh0GNMll
0HKReKoctPzCwzQQH8bSXiMHVbE9jAcnAMVPuw1XdhKYRrN4QHlo5AnZcCXujwoF
6OVFxgIyHVpWISYhs6gDsu9r/F2e2xzffpByDNbuBkYIb1gzwdChT8uSkWGUsdZh
+eD1J/zsbFi7oHQ0gbzcttDsuDpsNH3DC1lTUV9LiilkUKksoE71cnvX4aym2TiD
suJzSH5hTJ58xcLfw2yJXK4ND1U+JipnSSCrsfw76+aKM9A2S5Q3QElbf780a6NJ
peLSjBmbuMuyBpEe30hVdwBUmXhNs/NeB9t+CRIRK7fcBtRsh84KUs71+s1US6u1
SbR99dzMDO6oVkwJEwKG1CT/MRGjJ+1/QD2zjmtCzVjdkm6AM9PbIer+pNNUdTBg
KE0zusjn2KsM+tCIhIVDEMATqcbIoTzRDhPhmk3u4PLoSO/XEIXDEh3m7SHrnVOj
FwPrKw6Apdt/E16YvDBycdItFsAk6fHsZkC4KeaGySTKdT2igf4KJhF/egncVpo5
elO0cbNlIwUfd2jvH/9PHHg+PgHw3phrIQ/jOU4pNCRkZLZ47ebPZU77WgYL93g1
I/1nQperalkncB1H9e4GVi3qCSm/QvOQTQCZfAXwW7RUcQksc6atyLPgpqBSdQmP
zGMx0f+pAJCMbEc1jH1sZ/Exp2Yv5b/+K8CcvSFAmGGcB+hvNbN5YrQ0vOpnb5+U
IqiZ3/2ugHHl/ATMIhlJ6sAm4XT2TAjSomQRHbcHwTMaBpgfM0mQSwP5y0LWM4W9
FdGLqKymUJsCXFcPJMcYZBE6+gnKblMIVte8PaUj5h7SLon8Bz33FdDuCXvgtuCW
f2eD3BXCi0ikrDq8xpS5rm9v77lvwLnAw4/v0Y8WWPxM2ZggD3kPuHkF4D1NDy+k
YTvTT3fzjhmrkJ+RUcmbLP9KxG/E1KrV26Pu6q9ewJTNJptxoGLC2fUzOSQzjDSe
r39XIWK8zKG/jYv0ArIaD4JEON2gtSAd+dVtTejpFCWfuF1MoGYuhsna0hHWJbbt
IjNNUNCMz0e+4VHW6fVwO7kLcNMmDn+CGPQUexgtWdTDaxju+Sky6XzupdKUduFd
Yc+kJXgRjtnJ+r45zB64O9HpnQ7F/ulh0PlIOdQ0rt6ZpO11CR0+THshmSMDxakB
jdgwXK3tyw+itsvB6b/S4FOSqETiwYFXb7aZocHwf1nF+O8cIl4BPyI3/iG6pik5
jzs6tb3+b2BsVSDTqgYM6mAC+BbOufOwBeeTDCUszi1b1CemL7WFyCsvS2shiEcw
OeVfUoA8MfVWJYiO/4eHJoE5qhu+u0NIFjq7BTsB+S8UjDOVEftlYpQ9IMaReTTv
YB3ka0wk4mNfz6HlKj+anjLLMvcy8/n3tpKJGx/ZwfIrdNHsE0MMdZYFfovPkzdE
PL4XPvfo0SKSNrEolz2qeuU95MtnDzNNm5p63MoQdPyII2QyNI8Ri2zFd1V5NNSb
RBZFdxbxTTd1BqUM7h5umTq/CCHBMug1ip7cXn0Y60OZ36JvJqpsyuprhwfGj81m
TfB+ZTIjYpW7er2LFLj5J326BFVhAQ7jxVEmImz+jtqiLRqAoY0Kc9jYEsiBprdJ
Bi3Uigqg804+aeMiUNJ+Ek6fH2UZSAxxlEGpR5rfFgB4Ha9AFrKYJxlCXHybd0g2
6Dy0jP/ywPKowTYMn/GZZ5W/PWwfZECjyvtvARwXhr29CD3errhU4eNd5KglxKLi
nj2qcyPdy62upRHPXGct6XXDDFTlKKOaFBYdic7JAjOxBvyW8+CHxN9RSm9dsN0+
XJVPVHdKWkaH/+u2HFq/5qaXl26ZkNDweCjGi3PEEOgaEX9MzEEi78sG2Iw0/E/a
Xg1Yh7j1fhMcRCZ54o2SiagrYKLhNfI/ccWAXE8yi6OAnqrPDHgi5AoytE0s/Q2J
0ZgTgIdVTHrPxy2lFeZOy3TaDfrklDeFHrvDx3UkFbnq3WvPGdNkHn0j+IuH9rL2
m4eVQcXfgUQZwa3BlVjAJXTEFfpbTULpKI0JcJQ8NLrv5M4vl5d+ra9QPkafllrF
D2p91VqbLa1yYeia1EM1/1kd2FeO+ykN7feyWtDHz3IzO7w90mibtPXd9ij7QNhL
fym7unx2RtdVtfdvwB/162jzDipx+/u4uVRlK04W9Yx3ZaOWqqinNhqn7eRrH1zm
4pKHV14rsRJiwJMa3fPozWumFp3zZoe3EFzoP8zyNVeI4VmWYYfNaRcHHWniqTG8
dTKUBH83E4xddG1rZrysMq1SP2DguqZYkYTLTWC5KNUCnuJQAVUagR+zkeB7ulHU
XAh+nAce2kvEXqGCi3SANe/BdB+29Z2XPHQjPPg58gafkQCVXTjWHz9AE4sWvZJJ
Wgd2lQvuz1YnJFfSfp+6WjqpZtoPMhC/NMRy/nyf5r0pRZ4eWMYhomVWEZodTLcl
t3qAJ3I9xv+SO2ZJRZKeSxhouLF2zWapNLPd+u9spMEC6/8jppIdmwHX8+ZjSNqD
CZz/+KW0ESv39s0E9q2HNzm2DOydFkswNXswmb5Kwqw0lyhsZOUGBux6nsaQhmEh
A8gNHsQwp5gYQgz4gEBqcgOSVnBf1xcbBGkS9omU5SmcsrRTWQOdYcPtrUR+xWtA
zbsnh1wC9cTCk3Y4gjvwTW6EpD6bTZQM8U0Yhstcn0TsDk1OEHWP51nuPWQpkZkx
W0TCD434psoDEIRzIeHyVoUpfqycnxR8ye6Af5EYBbP+YEfqjEKUTbNjgHtIuwBb
Wvdr1mNSf8Tf25+6UaU4+A9YjqJVyxEOHdo0/WfANOVRfe0082vzSzcITh56t4T1
jd28rNEQqqx3i4HKjuDwJVzpvd8k3dm9PxTxPPnhBm+/N1Ouk3aRmrauVtItm8xo
Kv/5FGgtSyu68//NX5F2CO96mUWZs194zMwdhLuroQlkrtZwzm+mKSwXYruKz5jG
SJxBuU9MUgbGNu0fTC9NZKZsEppO1Uq94HI1p3t6M4x0C2JyVhqaSPSShYwTXVhR
KvEDjpa8es+jvRMhHyoAtj2Nr0ers5eM0vtcx/T365wJLQXhBYOtjWnygTW9/GMR
d29OPZphrNmFpxjkpevGeYldF0nIx7q2bzny9UoOz9XzjQXxK/4OETxOxZz1qn9r
ptMxZKYszqH+fQ3S6QfjF4gK57+Wj0cvwXPo+ti+A+PTlRWf6AVhkliqL1mPeqr9
xSR2TRDBlB/oyNhzMdR6hlKZXfQVhzP6pVevRvLiHTDo9DUR1flBru9xEktAjnYC
t5ga0uTON6zOTVwzds6oToaXeRrjNfV4xpzG+PqNV+xuBW5tobd4B41eDLYMFZ87
m+08HF2yERXBo4dCF/NH0s8aei0lZNsxlsLZ1L51KWoSRa7wD7a/TS5nSm+ZA144
Ej/EbmnQ8vfeS3u3Sp781U0cO0ZhTWd2XxK1MGfhVpmM8pIZ45V+4xcKI7MkTuSa
+NLOiQHnqJdp1IgL/TqNsDscoWzELOBY3xg65oymvy9jLs066gDOY9a8iadWDu6X
HCBR4/exK1RZJ5TCEAhuizQiLfAZ2fcwcgtnk9en0qaOHSYxCC+/Sevfa/8lGYWv
1yGAMFdwOSpDtcCgaYUpZkCv+klcEo6KszvZD/gafx+RJY+3LVpDeIZsjsrte/AH
4rz4sUIKKijKiGxCSj9EzmYV5RPY9AzflHpKMib5X9UuQR5JEI+5gsgxwKqcoV5O
F3cwSrP3RDRtCHMU0Tv/074TY0e4GjVY/7nQXQg9g/sz0CTwQU7MZHiLpoH40Uz3
FhZMloAiM2WGmXuL867IUBxkiss2YEXvG5V65MiLwRS5V0hC0cFvYDkrVw4UMLOi
0S/kYYDSOw0ZAIb2h/qFLGe4ptov+Vdk9W4I6xCRu18bZlnoMuKCodwrhlt8tnnR
cSXvlcBPbJj98UPsBw85zs4X+QAeI7urKHFBmuaNXyXbdWBIs7LaQNKPUZHW0Cwb
N/90TZ8TUPsmCd3x3DCZDr8H6m+I+N0uFRG4O3qTfpzPf1Iddwu8Nwyq7a47fwMT
d/NJsr+hBC6yui4ShBuhh7+jiwMER1cTh/vzlimIWbKrIjpSkM7yhh6KdII9W3/R
ysLYStPm/Acd9GYUd6EEu7i3Vuxzt9OyktZlAMFaMpi5mN+9bp5/JH25slhlEbXu
bg9dFamJfTONCnZGV+UNjsrTzJXFu3K2Ut+5tOZsn6ZTf5M9pOAhWBCq2wX+4fMz
cSN8lphYfLGVURqtyNwI+gCzq1wK0qeMA6pyzH3HDAEa+ETalkDfOKaRY/F/CXZJ
LAAzLdILHRb/JQ5cDOEBggYcLW1vhbMEuKwEZjf20PL73Oyt6HswsrH+uzqwvgcB
BrYzacEr/oQNQfcncht7PLxPLQEWeXb33Zzcwy6mdzGS3pMWu5xSBGRxqI18rd6p
vqlI4p3/f13sioa34BDwGjiWQI5PMqm11Ggyc1v/SQC3zfnR7Bw2Umj933ad3JMd
1rsdz4cZo1TZDO8GnEA4l4D8pv0F4FHXPMunP9JdZUq77KhqZrEEm31fmNISA/Oy
jAogym+zQdi5ADbFdPWE9dENuE4Fe+5b1JONerOLXMCGYPQCq/zSlVD4QUWMzDV4
jbsiE7N6AkgT0Qa2cZYkPzsNZFD+GXDUpj4v7az8u/pS63++1xtZL5A6MRqOUVsk
N+9SctGPOKfu72VNOUX/HnV0f8Kk9JP13D6+xzaN7h+VZyE4X8dg2iUHqkdx9pj8
cPHXvtl6VLq9L2f4w3FElljy+gAhAiiY/Kq4Xid0B71YXLe/sZpSfv7gmatMwRq+
FJOd8LONyUywqbHetcVj67lm3eJ0cParR4u9BcIPlI4mmPrglQaWOtUtMCEJoPy5
NjfUNRUCUMKE3ORVTU31Yhb6s+qnsfkhXhhiUJs+pLCQbu4JkGbMout9mA53fiyG
PzUdJ0Q6f+m7HYLlYfX00vxCFT03q6WuUydztMhWmB66eLDWkgdyVIgdSqzXBhAb
g+L7RGBSTeycrjWQx2nMwBPRWrrW7TxOWjW1x1U2IfBXyM7Zgf26NIdBv7nxB43m
OyQS1hnjV/8bh3qSIKAEmd58OUShu5G3Mj5eWcHQh1JlVShkMf6tLDyExl88E7Rt
cG0Z6wA6AUA0SD3qw/23D1uejGrXxbgaXpE7uQGLGlGio1Xlwm5Me+s+T9pA9uvD
KsFwZXrJrjMvdxbfIEFmClzEgmhgHB49ixvqQdlG6QuwzxCTFnaaRHjLDILsnJ76
8XeIuhAMS9dkEj0rfw7N5x7rtdfLw+ItUAPH6JPnjIIndGTwNTHbmdjPWQaWY5NS
kToSQoIUG+R+zI3tnXC4nCjK3B4XDRvn8bAGjj+iq5aLhXVlKtTZVAL6IklqiZIa
Fhxc6OihDA46xS++rpnDTZJS8EZamxfyoo/X8mebWuW1+WG6o4D4Hi1ou7fgjC5B
FOfGasUIY53rZK8+BuAeo926skg1pgDjdOGraiukJtu1O2IeHKdx1qbT1sg/jisI
IWRBaXawVcZPJtkhj4WNjMQQ5EFq04wns4/gxiygH/brlaN9Y2Qbd1beGBZh1zvM
73k5DyuMKBFDhyG8uqnEe7HwJabdm6cxJxiuj9mo0GnizvQf65CBagQbPiP+iYDu
k8gh6QaOFc7DEGRlPtZFmhbPvxmOmrhJAgvUV6F5vrtzjVmFG74v+aXCEy7oH626
hf7LgjzhMloFg8wi0cb7MRWbCWF/0AktUtSIFWCCMbR/Lj4NnOuBMyENDD1pCCV7
b8JD5ZJMu8zMh/VpYFVKFQlQSR9oP9+igYdXsFLTW6Cbtwqo2BSsNsSaduj9NTfO
9rmsWW18FCwPPW/4zkFSJkx2RRxwUtl5bAdtwXdYx/6OIWfHMjB4xlRe+FT//+rV
IqZq1+80Wd01epM/g85hZI0VvO7uiXCJNbNWj27tDCKL5yikf0vdwWN/fZs0Hq12
ekzTc4R2swgJGo7U3ZwUvGQSXHY/bFn44nE0Y1H7zBYGj0d/nUmFiMQhH+QuLrIm
n4ksT6Q+Y+ia53avEqSXpYsskY7vd7yXTWrOK3OR+bdggdmUXuf73tg5TAc5RvSC
MzPcs9YGLQ0v5l/ae5PzTOQv6nC4KY31ZnZzaxzk655HIecYiay/1AkyBxv99enV
2c0/KzifK13FKnSy9LwNpVH/b+wBU42WnqBXJIJmOJr03jX1uRU3cEKrUXrXJlbp
+flAFtxmeIj63vtEwqIl6O5pnlqNRo4hdM2j+WEwBzJeE0zH8wCJYmbRwpXZMGnq
MykIpMdDl9pHELo3DqqHsuAtP31n6yR8iGLoGQmy3my9ecWR/G0P/nYu0raaWXzQ
kEbcBf0vFFBcS+C3PdyJtAn7KENpmfpeFiM44B9jAPNYyg4yGXDxjyyS7YboDzMo
OtnuAzPXaRgwzKxT6gWp1jkI7NsOCgvU25vfPkBPqgJR4qnQjnP7WQszixgXTc+7
kxyBhxhZcJg5PmpomhaLKjzrUdyTOCcQYU8+uUPXV+6pwhpa0y+6kba4PNGjTTXl
VlPESSJyO01BUcMIF+kL9xwoVQrK3etkalidZoerNk2Zt7ZGSN75UxDMGRRs59QK
pAmDHw0C5vPqfbZB+6Nr36pL0h/DVp89y+swcQAV+H5z2kYj7BD5o+zdBs03bjRT
kvcpcoGSBaiydNnESX2/MOSj2FhYNAT3rwTP7uK/hSr9fWbsa2BjZd0cSM7n31sZ
/BIKPb8aUH9ApS5rO7KctD80zIpO1Tuh3s/KUcie3qzLiN6EaVJGLt8XD58WFgb+
EdL9SGynOdu/YG2Iymay8FDUAqBu5bS9JhhNCSERv8SX9XOVq5BmDeSpA6pLV8GX
tnEva+DJOxvL8UaGSlYDo130RVgBaIJSmsBzbFeghi9AdTVUfV99usJO3mJCaMFG
Rrq6qn+WHNIFNDfQUMlqQmzTTCHxF/OU2fq7oIh4batdng5TZ/hpPvoXGGWeogB7
IGX2Z/8h13mQ3EozN7Lj15yNwo2CbI13dIjcj1ArCBfBxWErFVh5W6eFWyuelGA8
0hLT7T6CPUtAzsPa181y6VHLeqIOdWBVoDWjopoteL3aM8LPQLUbzTxnWi06slhK
PgMq2XI8eMD7DkAnosXemIuc3J4XFCGrxGY7OwHjDEHUfAQB+6DPt72bPG2oAUb4
auwmMMrNn52CotCDvRIypxF6pHSxFhozIVp45MKZn0k0ijvW6lelP0v7l5jOXkpn
WwGOjeOyE1MVRPeCbnE06k3wDGBV7Us/jqxXcdniJWZHTP0FMYqB2yWahj/VEP07
aIcjdEFKy2g/RaUpN73I+62Op5IjN0UNF2QC67/HB7ztMOaRC4VRGTONUNRriEMs
rlw4SgIy/s9+/KFmILtN8K9HhC64umDwnUwiinsJiGbYmyLahKz+XB2lIpQu52Z0
ZSgwzvXfBaE+KpVbKKZjwOw50frlVEVP4cIJcjZLWw9jeloX8wCi8mJfr8mPeqRI
01loXtNPqdS/zqEPE9xxoI62mEvf5zY/fJkeeP5W8IWmABxtg4E1z0S59CKn7o5U
ENimwi/bAL1VGuWQTdvXl5tnhhX1lDhOtzmKv0WRevwjPd2+mMvuD3ukWAHK4cXL
ECiCZOJJfK/4sZ+5T7iOJg6iHE2e9Syys+Zkiti5esEoyosF36INGwPP6T34ZX6A
Crx50iHOtNy1Mp3y1rwJjPiAKvluNTBaB6qrKOeFKlJto8lV607eo19AbN0oOYHw
ts47EJ1+nuyTix5wRx+o6D4saS62nwo9zHlVAo7jckfEVJrARBR7o5U3sm69C97U
bvcS6geqNCkTziUqfB2F5QiI2LyZ2fLdB6kMOs8IOvL3y2Lkubc2SwQoxzuyYwNr
W1mn4IUgazHxVRrPCTxyf5fYhZ+S0cAowiJL8bK0nNnhJohPMJy38IaFFXWSzzsG
4BVmcZBclZVE+220xAa8Kr2/HaZsoEZeblNvvD9jnCR1RKhHQ9ALDWkuG7DUnLjv
8RdHZylSbEuP+6mVNC4numqw3UdRMf2TFsdRoDh/jwpLUDxzZwZDEzalTuXbQjlg
HjW6ZxAKsflnww/o7pZFFVlC8hach2VKaR90kdIdgNGYVzYsopHptTDtrAPrLNbx
oundvVIaQIQMjNsEJk0aECiTIlyu4qgz7tSWdv7Q+aprC2iTQgOb84iF3l89581K
zeOfxWBaZh03S2Y3gEbiapjog2wEQ6xNfEzp64ZI+Hpq/8g5VAoWCQA5wqY6v4z9
VsRYdVa08abyQNzmQckuLEg1l5Lq56ol3HT2YURL0bz60XW23W7neMnZfuFgVly0
i+XCJ3ULaQak/N/Pxu3jTMziCzzmNOOQoh+FuHFG7ki9MVJbuPIgV/1R/pBEBRo3
/quE1GkG2rpgi/BWuNjU+2v4HWFN+YiqPQQOhk3wdPr1RWl855spxKmPf4gE7o4D
RWvdwzdfd02IhXO8V2BaALN9YQ30kBo8bTseGa6eX1u0b0c9IxDwCM5hqwVHy+1M
KLaspmXYfwhoaSf3W+HCjXGoQmhnVISrmzgNTDEanrTPftAFBoL/6jhzXEcr7z2M
CVXN+vWICdrSfljnMCBjmQkHKpuqe8M9V/0z1tCK5Mgxr/qK8dt+lxKL2w5XIZpd
3jbYpLGUz8y9gV3S4LAPkVhlvLI/VM/qZln6PqiRAA+NNDzBjnXMPtYlsoQ6QMJi
lilHkgEaGfgqsJWLKHL3taTpHqPi+9JPFpittBSkhqKmRA2FmhxcfLyYmT3/Gh7X
ppEssBiCemnzx7ldL765ZNyG0fe9SdoOB+/SexWtjhJQ6gsYZz9FRLELIvtvarz8
gmYKLUjO6jZm0/jdtmcvKrmJnrt3rqVzRktnJX0v8i0BdD4EGaDFA+Rf6u1eyMYy
wCEq9G99O5VvrlMkoYcaUFuoWxsDH9eyPt9iTNjGBPlUPaXzCwHhvjeo2IIASIU3
curP8VQwlyDoeDuRcbRQA4oaeWEb07I5EPWfDrQwZpRIoBudRQ8s22VP9k/EbtSQ
MoOcPPmrcGs0QhASARerXLQ7r+nocN1tIixFaotINOb9dyBXlADVSlIf/DndyyeA
03IeO3eK+TKizii1Z6sdZq91einIZUfewZuUIVrrz8FzzAWN1EkHJNFW53QhEAju
2/LyDq4Cze+fNJZj/fKw3IVhhFD6oqWlPi6Km/s2RFOqlVRCLGtp56ejKkC5lEZR
fAakt/E4wHt3MMtaC3sTyZF+z0TcSDZrUjtDkFKMZ4VB28/IXX2dPUNnJ0FFFY44
O+vgKEVQO94yV+54f2dIaqOVoyswZ1wmO2Cz1EfJE8vH20texDtJFByPsYAfHecC
g3pLy3X5aRhtQnMfwa/Za2AmAnAMQ6oClJImchaXb7UHqLXNviPjXBpP+UVNQBV1
IngVfag8q2JQpUjT9f3i3wwnbQ96KouKVJ51DpXvSC9LjuJO85zEREOEahERnCfK
ODjJN06XSIlNtapQv+avEG3KHRKdrZ91pK5dGU/7PNU4LtSy5Zfd5bPt1AQ1NM2x
hDSSPdrAJuMuruz1T4fyO38EjlmF4MOLPzE9fO/bFO2SDzorWKbpLxTnZmSoWXYO
SsH5DGvG45bDdnn5XZecq8TTEkzirm+Gf89YMu1sNlWjew8HujB9+SiqWQD07cBj
eP6fpmqypewISafXyavjZywH8knzdxHA++XnPtxR/493yzPNVNcCmn6O/3fTAORP
8FDh2BN4QaFGTJ+wqO4c3xzKhK3vyh9aWzMmEhXsPbdO/DLrwaVu761FKjv5xcmi
4x8W9pG38b70haNlW/Iy/tBbfav22lR14gUupujeFCZRL5yugEsiIX5UmONyrOwS
A/+AO8dUQRpckjWVUXX8ZbGzqm/oDU4qbldObWjCl4Loxtgi3P2StEL/M3IOQVKs
8EhWUumb4exfMbIa1m5YObHoZAbXNRiIBrsFCwkhw8qfeSdj96PVZPGfL38SCv/v
suExpdzXC1PZU9s94RKHsfPM7b2TVVuukihezk2veHjFegNEhtLT90A7AZ/s5Rvd
OFYoLWuozFmrpZkaZUlSYVEpnOm8/4gPQnnzx6zVf2mmpomFfr2rCJTMudq81muW
O6moItwidGTu/pKSZ7Ak1RWS44MboRck5yBIoWvNEgfHueZ2Lb2y6Wk/9voMsval
MMNeorIWQ5lIdyqZJHRquyztELydhLvpoE72g7DbXZU182Lp0rg4hFm802yyPPis
JdKnB087pGaWpyG9SFXuoivDUmpIbNeypOizqksiLSatkc7ruBEEPDvl6DubG2jR
+HXqOJoJ9fC5n92Z5dnIQLWvM6h90V9UuMc62QUA1SXc3NgTVNIRoSG6VV2F5qq7
5ghMlW3ZVi5frwdar/t3rMGOd2scrJjR0aDqVXAsjZhNqcbGOak1r86jSgSLGi4P
5fjYOcOdKAgAPn/sWwYo+40DJr7raxAdatHQkPJO0J+Vo1WkVe0LnfyCGnhAdFa5
CBbXR12mLlw5E7OCs53F4MAblEzNCjR9rNBczlrkz9ZC1PX+Pb6s+Ip6Ksau6R/p
c3c80yy9Azuy21F9BAWJIgUbu3HVqt4L4vywRFOQZ1Czgn0hQT9jq9DjY7SXc4QG
MN2pw7BqdHSOTtjwdDHGilUWQomOOnGLeeA2Bz0yvlAS1DEylq+46xuqt7hKVkrt
ae5pWBHycL61BWGMlPA6C1Cz760OJbgwhzJYjxxYJGZR/TL+Ux99dGIse4LV1xI/
qo0BDrjIH8rS1Pmy1LEHj3MN0btwXOFSv0jL4VBppdMKUKV/vQ/dT9b+471g0gWI
hpZbQj8cPoZgIjCYG1oY4oYZKLUNLx/GT7DLzpgU0izu0BB3TnmDuWYtpbWOdiAS
66EbwkWUo3lnqtD99Wfzaz9UqxoHCOYnZwforiE7Mxmen4DEvH03XoMCD+adIFFd
NOXyqld4x1USrnwmsqq8t8T1e0Yo8IBh/+xhBDXs7LQ632m9o8gQIabpINVV1Po8
N2Sjz/DjEZWbS4JfMO58bOKf5ykLunmdu5NKHSzI8zEAuJZd6O7j2faWBlBrzv/A
wwBG7/g2J9Kh5BcQsyJln3gPRb6O0aVlRPj6sqyruz+nOnhlA0TnVNjKQXJE2/tn
5tMVl7zWGq3m4TrxP3bOpdoPpfkfImn0QsYKZyIVwdwMgHp3XsLoC0I7IMu7AEsr
W++jrTlogJFkGhzl2iTaSLEwkT6/7kEb3yJzYhdzHRBcGAK9XI0fVMoApt/kkEww
gFzuvzLWhst4GHRfyGXb34NGUTSy4TUmy5LCmd9lihW6sB6TmbKQgNGTvCBnuiXj
09HvGv7yvnfxf9C8+HD8NMhx3KlixDackguDC3RzvaVrFQrttRq50qm7IroOq2hg
0fVlwNehmZJaqkoWMYaq11A3VR5LGjMFRgonDkRT0gxgnnncNpUs1ovzqon+Voq/
bQU2teVtrTd+VHm9e4Bvi7rA9s8YMOx6G1sucX3Y8gvbeykT71xQanJNyvmdpMSL
6DVPGrxt2IoRsc4zuK0QGtE4med05PMFZH9t22cwyBnDQWnSkHF5WdfeGaYPN2XU
Gd08k9KMJpGKChj0kimvgLHmyiIrMqRftua6qRXwHpr2hjXlxqwEB0Jolz1KlqkQ
usegDoT6Tlo2U1z8nNTRyEW+X6XPpyRllQNIQ973c4P8DvwXhLs8frSCexrADeLA
6ct5c2SpQqQb5zxIjEod5ipwlr7qfOJp+WS6WDE34LrKzElJzizepqvu1JdVeSGv
4bltiHXFipn2vp79MNg6BTlPxZQWydElP+Yh/RREL4az0hjwNI9QDoa1tNM3yB+r
oZOFeBdpxR/pHAYZAfZkBKepXOcHnzHlv2F/oP86+l46cmJssgNJu9mdj88uheMq
TFfACr7tQ6LC0LlkHHO5/xoLRvjP4wFjLRbGJzLReFJ+OtY9YRkPyg5+nXMOxVPS
hmcfDN6S2g+weKuLM2zUVhlLnAlQ5njysgwR3QT67FzbsP24PxV0+OB25VYBICYG
flfCPLKswa2d3F4CVyJ55can4SMuO3U7l1P1rKjEsJXNoHYWIMcOJCeyygx4e8i9
fxkeYR7NdBJ6AVxGDrnfdBU3w3P6HkXwH+0SE79ol64LvTTX7MakiWfnlzRmF48t
wGsbJrL+L3zwXCZt2spJpojEQMQEUsCFDGTekxmbIf0XJJEkRISCSDwYKXNnTkOn
4med2LPiBZtDd+t9W3kSHIZVKDzFi9BebFoq5lkOM6Mb0S8M/aZIjfVHxdPhjMRk
3sQzTrm/BXmriNVqAOVeeO3QzM+lffL3EMJT4zDR2y1rXDBlyOsMRfC/aODm8E+V
ERB6UwovyESOZzFIJN/2CUMY4KLFJcDwKRZ90qJA67rna5dsCVMppIiPoMOKTpRB
3ZWTqrxCSh5Y1hAqpOghRatF9AiME4keMwYDX5CYBdPyxWQx4vAyXjJlnJGtJcxa
4QnLAH7c4/hVKkF2HX+albs3WI4UUnr8XDj6gU5xUoJumxuPLsRXkzNCo7cTswpK
K/xsExEZk28eIn65y+MUgHRpyv1f/3B9GOmk9KKkRHQlCt1Mmh1yqUDpCH4ugCm2
mDKiqCVO0gaIxxNadSizVFcjMXfevaPrMvnMh9bI3sdrpUvgv8Z2cvB6IRBQcC2v
GXsVFbPtPJWrO4M9gpSBeUx0xa6oek89hAXCVaBO6ajrZKhLFGF1JzqmJCSN9osU
AVw+mbRbSlc0P6zULsWBFSOac5M/PteScBrvFdynZ38uMWEtp7FBzM078sFXiKrz
3Oy5x06tPNtQaDngsy9d55wObfZtEl2yI8n11yhivXFEt9Lb/N6f4BPt/z73Wmro
+yvP0kocqjHDE4tjTTxs3zIHZFXR5hg/rSO0dragdHmjslYsPZLE0o0FS7TxD8WT
Jwgk1PJRuYg9Y9Y1UBRoh85+AC8jlBZrh4Fx28qlgIDF0pyPuWgLoM29YI4EhfrC
8re3JAiX5s9fJwgjp/efUqXHpbz1At206tY/M8B8XumebRhvsZ8XSs6uIT10E/ir
LmnlE9RK0308JNrXbbwEvf5RjTy7Ou9Fu1eUAnUzy30jiCHFL+oXx+KBRGbrhZMg
UEW7A6C2gYMh5Ik3lcWU+LxBref4mkVxdg1AcM3E6kPs+fbcs4BwMLP6vqevv6Yc
h0icV4Ggf0H0MzqRcJ2J13zGFzlEcASvq17f/75IPK0uNpbo/ZyS/7Ge5LpHJ5o+
bJSlmBpWRCr36B33iFdmiYMMNUofxhAghO4g7XQgDrJZKX9a7JIXvm41zJDv//fV
4qUqnsGazUbKrh+WfChXD1HvroQLhF0numY6PvqP5LK00QTwCthqGcZ0aaqQtbJu
BiDYgGvLe7/gpKZLg0ABvEB8mXKWBaPXek2/QcKKiw8bSNbGZaAE7nJRHdZxz6ow
u79MZ9r4ptyYePeXFVGKLxGYxXwWtJdbfuy7HpgBm3acMPCc3PsgIBrqbpeiOimZ
cvk8pdC9IgkQ0hVkx9iWfN1yrUUBVj2xpYAm3yATuCNNcbCeYUnDSaxk8oWOLMa/
Xc7CLcH2yT8fkDGMOatwVp3Hzhkmc1T9Ls/PBcuDWBNCOmYiuOUQsm5K+XnTgl3Y
n2jY4Sz1l/R7HrDXZib12Fc03GQOwwm9yNe4nN+PiL87CJRS4xQI7Div/p/hj/Hs
XADUggj3bDbVdGxTZvVcuCrl4Q+S05d9lj5CxfsgjX9ihjLpB6Cufuc2lZ9zxr7B
cMggtryjAFvgMkPa44RTNX0UvAP0R0yuGSl+xqm4yAcWDUwwD+0LyZ7wTDDKdjcS
zDtYWmvnfNqSQBUBXB+XPWKgaT0N+4I1fBUHOK7DrFXmNWRyfaaAZ+u7DBdWvn5N
JUWx/3OTpZznZE89ol7RH3JIomJxErMmqL0nX1pswTgvZ8IEFSwcTcdQUwHilkvA
nQsOpcUvs7aiJGDnVmUjyCqbgM31ET7g2YuSgXywkfHa1II1xCPHt4o5u++0MwCU
rTvDvQuTq7c9Gc5+u26vExrRpdi3ypq8Dm2/Mkhso4KL1R0d5Jhb9MQ151v1xh82
h6hqSmZNYdWvDqr89/ZepxEpZRIArrWWfLGCPo2FlfLDH11Re8cKN9K3jaav7jeb
Dr6YY8JIsBFoAzGEL/xz1vR6BXh18DCJyO8zXnc6XOu8mdEc8bVm9IxsyMVxFeq/
iJ3o7epenkXrPUz7OqezCywXYs24RQsV9zGWOtvuxRv6JLpAxRD5U3LTTRHK7F3q
vjgM5miFKNWlORaHlzyZzAaQBgZykhE0WixyfBUsgpXw0sK7pp3+29vh5hOhnHgJ
I9KTT4CBrMmmMUvfhFE3PKD9HeDpDBWyEOGL31Qzznwny2XbZEA6JMD0EuO6fXzn
P4RiX8oW5kZCoMQYWzLjNBKhWLOTjtSiOTJ57h1wcEb/1GcojJacJejJZMwaNfRM
RD52tdvb+7R8vYX1LggKco4kEyTQNvtT9Rj9y3Y/Z1H6ifVAWnw5t+69UEGZTh2l
uWfVW+9JCmP/YcUochjEILOHQpbrILfe7vDoaMY5zWflmeSIrGOgxTeVzfEI3jYq
qTFLTQbwQAnIVjIh56UrkeKeNLAe1wpBMklwDDXyGz6+A9ltJpJuzT7dgPdr4isF
WMMetS9UilE34X/WgU5E9//Bng1KFlM+g0RkjCjsGTYCw3rSGurN7OlwEDyyHs+W
fUdFBROwSFbPophsX3mSrmdgMmaZyi5puilZvhSTRIzjmSx98Nnmkse4U7GiMtIS
u0o9SMR0qFq4mfSlUBh9tlx1Tx1/Urwv7o1y2o5/OvfFRy53wWWqy6mxrhr96etQ
sGLOWSx8iPcN0nt1uAJZxotDHBFVoBbk45XVxX4ePqxs+fp42J1pPI+Z+s7HW3Mi
NssunrqBu3vkR98gEGFukM2YdY0T23hvO665TtETZjCHgpcfErhOc5b6xXGakbyQ
IhE2nxerMstqaoVCN3LN1uY2s2hg84khfWAJt8OcNUSbxmtpmBe3LIEhdAGwSdRQ
QqJKjQTP1mjhOlPIV8iX9XXqqX9m52ol/qXMWlC5QbhrZFkFHMGbPvFm8gOuvOEr
5+wh/cmFhS5PjZu7S9pWIOsKwjGIpyTGfUGDj/KdvCBUNjoFo7RX+g8ebmGgS518
KNH2g/3cdxxWHhtsm1ZTOZAqiBTxLd49iab5imbVu8Jw2ZKsLYnj1KvbCfSQIu7t
dNXnnj4J3b4yHPTDVKMvu8HTJiVMDCayVk6WAM8nXZiQK7tPJ+X7u0nT2pz3f1wx
TirjfR67M759ythly2LefkmTZ7R/1eXxqZBwbGxO7ok66emj8AYcKmHc768JJsBy
vmbtVIFk16+ultTkWlNStpcGnS4ugdKkseoGghF/mxWLEQr5actKdlsKwN0N7e9/
Qa9FMrQufCbJca2HtgqL8uOSLVbvSasQzNnNMRT9gO/m3GSWSIU4blJC5Wpi9pGD
OosWAP3cw5WphhMD8eTcQAtq2oarMR52GxUgD+Y3s8/g75vQxB1rrZGsnPO3uLc9
kyG9MeWzoQ0PAmq9GC9Vyzbqr+Mjxladc4ZEy5er1PWtW/eGWZVLB46BasRnnfLv
jXkXn4LFEzPkrZjfCg+V2MYnOOK5ViPpkRx8hzaGikPeJRNbb4YZBpTZPbj5qsuz
rzm80K8Ew/Su4kgcUHmfn9PWTCtTRKU/CM/cp/e5UmSuplqKNMv1CgYehFAZ8JQM
x0Fm6jSC3sgrIZjwtCvlseJbfgi1pAEGWXU1TtolZchCFSCkHUgVlX1TmhlSLI+R
v/jHOZdVpZEo6mT6ZayCNW3OCYCQ9QPWP1/cdj0W3vpJn/jpXOg5DGe4grxQMbfG
mkJkEaCxZgsBFOg58QYqOKi+gYZkGxqeth2HL+wi/D1cM+4d++8FnfHXFfdht3y8
VVpHUjVlreYiMGt/2Jy91S58zUazonHJw3+t7KYpbqjdexGVMQJYKPSyn8syAfEB
WxHJOmZv4vzwFQF8xv85y7dzgr5x8/1JKBSlx6UKVe555QCh+jgSARYAxvOUDhqe
vR250poHQRdhmx0WPfx9peQUUqJTxsPgTURvo3H73wjaTMTtkHVwk6+UIs3C8SOv
xWjK3mrE6gnNrY727fS1hHryDm94/oUxFK44JNncJKSGXm3maXFPeMIjHdydTPfH
KYbJf7bdXDx5FUG27YdBJhf5i66NIQ/acrfaoa/WPgqbDDcBPbuL4ZacJRHZ9rOC
E1iOwKymGLf+raJrIl+6UM0lKd1wYAFipEvcVO82dLwbjEZJCv3FQRwzvrT+uVDp
GSBA3AM0JG5hP3EpRVu9HTWUlxgSh91t1b29nzPAjFfIVQep1LOyO3b5x2xqInLo
LlKsFSkiKOR1H0GrcGYYqr2Vf3JmlWYln/QJnQu+eaXFmtwqpn/oEnJpnB8X1ngS
5qcKktdZB+Z/DelU/qYHtcEgwpz4vwY/jlw1wyRhYSukIlitmdyf8ieQ01YvaIiG
CN+rj51hoGjk3RefA+qAHpuOZcr1G1IbCtcfvjYLtyzl0FEkmXAAhRchFksU1XnK
8X1a2lL8rH3QV0FTQmWDoPP6BLB080KUH2oVwFEtrL78KnJw9DSrAwX3VO6xZdIl
JaegqNozN56150puRs9m/l8TLZ9XfOpuG6HtAvivAs0pjDUsKw/PcTaix4eSpwid
8Ft0qTGFS3Jz2t8G2Qf8lyUUHofvJdrQolIqLgIgf9HSwoE7P4kKOfvBQ2Ayx3C4
Mr3G6vGqJp5pPYNQsE5CEmKme19lGiiiQ7HEOrZ/qQWuprXrYOdC+peAwimXlNjZ
3/J6N7laIHXhbAZuyP8TnA/w/bbiCTIxgLAjrpWFJB8ePWuQ55oEyRHRP4QVgIGP
CYAUElbvHcYlTRJruFsSwFu1XduxUXb/T568+6M5Wos5AjHZoMpVXRqkh2esZAqy
59N2BYBqFr9Bn5+b4b4ijdHRVQjewv4pF0rfwhczv219SFjHRLgr89TIocbNBTCU
gpQ7xeEVWuiKYgAJr8OEfj1ggKe80UB+iajUGJd8NHO7cjg1KG7KuHBN/8Oy6ZH0
RF9iWSKM1wZMItX93SCn8rgts8yXWLVih6GR+6UAbQ3Ayj+uLSHXDCX5Df3FnNXz
rYF6j67YBAMWyVaTp7MsRUpQu/6/CX4GFv4y/bq2aP0agyWS1guMK88XAY4/hnBA
IpDMelc6pPnSEBR/FOtiqc44fhUVC69Kpp3mpFLEeVSdgjgKyw+4EdzPEwKyu7nx
+Hrl4bYCPcb98CbNGrV9Ngj8APgD8YUCiUqwn8EXsoqeTH4UTEJ0znp4l/wwtu8l
Bsjiv+cSyY9I/D86HLoe4bi/tqmakzvGD4TzS7SewR83OviSrcQGPDk++Jmhn1zO
+n7cgoD9lCzwZsuzxn/soGIi5r1vO+XmED1/6J/TwdCzoEwwJBoMeC/4Nxk3RFyK
eTeQClz7OsGA6uZwAHOFyz7BKVc0zz9rMXyy9woXiZchX59NUjgpO7tzjLPjhvmm
RUHvjcTKQWo94LF/LniTO2AcQHnSGqTLr56mSsi9gU6XNyiN0SXWlVNd+d6x0z7A
yXrXKZr817DQSJjwhTdLVBnuvdSFKQldUKiI+E6uBo1b5UDencfr5A8dPGgGLPWY
TEamSqNSLXltHzkmgP1EgRiuj0xEnrGX3c7TUPM4pvEfeQA93ZbKetGVQ6T1lUPF
4f1nDfmX8uDYmszGxFnSRQlYSooV0X6r78sVrWYiY5Y3pH8u7A/GCxk3hx/9k04K
HkA/Dj8UquUj+oMBo2m+SeBrCL8YOnx3RX38hQZDjV6CEPy3OZxLhgsqVgwCngeE
bnBbNQSFWo3AhToSn5KYpUSsHpsiXsUNFOIcF9mIDiKw3Yo4flpj9X3R0YM92hrH
tBo5Fk2BxoIM4zncl5XPOwV7bWqADtjPI9AYkkJq5azuVewkvEJtve1+YagPWR5K
7WXuXDQiTr+n/EYBC3a8mEFkXDWKO3QClalyxluZqgzQ9sxznEJk6ngF8ktHS+ny
TJ6zIrAyC2shn134M3ALQWbU0i2k1Pjov84nYa8i5hQ4T1tJQ1UBhVuK/tXNzzrt
HEhgQnXoCyqUBD78N8St/wOMbHloLtW+lEacrdhMICBS9kA6UftN8Er7e0QaRdHt
UUsZuwulAL2FC0ROkxDyvOBhAe+wpTywBX1wNg9I9xHfSgeRC172soHa6VeQ7wxZ
mh6VlYbmOCiKDt/yYWNojBXrAl0hgOL6kmNTNRkG4R7AWkLp1/lxxgqpWxnW8CQI
X5sYaNAC4zo0jtmtgd5iO870U5D0TvlBIPLEiJUKrNWTntL4UPneeLYrWexAII9n
eg2A8Y7w4AhIP46u9bksBRzg+YpmAR7y8o6dATxlX9OXe4kFWocwqgbjyBwaeQzs
QE6lfKjIdlcwmQaAsrxSDd2gzSSLdFh2taynMt8iykppNAcPzvcnm8FhN8eKWnJH
CdrPi2HGfak5FLTWmBkDMCYYUgMreqADagS7bF7yZqGcVdFZtkJVaxTEHhw/V/9i
MAfCp9oOuAueA5mmFNohxY26IcqnT6vExinBfLo/0ypgCFgsBzqZA1uSGnTioVwq
XYvHglO7ZOToJ09vdX+NZnIEL9xxIpW6h8RzacOWA1HM44S0pumC3mUnkfKgItPq
FEq4o7sxcrkpd8ICyPvw+nNVRnRqWe/qyA/1IPAWB8t2SSfT+8obEu2bWWsKyGos
qoYq2q5mnmwzSdo/ECtyX45AZ6ZVOb2aygWO5TbGAC/1nv9g9QJmYR1orWH2Fnwq
uDLhVBwY6tITTL8YJZYV+bcT3uMx9nW/zS5zougcVHiKHEcbd52SQCvCXcHPiyBy
O4wOqdoge9Aa9IawN33SjsWcqez1gUExIcAgGsO8uOWTLXNIdDigUYG5bTiiucwN
/ojAmPmJJX1ohfRmdxwz2VITOKytadywXAzpv55r1wlg/Vz4G3/0U7c8ovymANwg
vOcAvJ4eF4l8RiNiXdAdJ4cIzAx7cGdcNdpcGw6yeJSTl0uvj7mFpz7gf+DXVQaa
q2RXH/Xh0Cm2KuuzTeTq3n0Q7txAeKnj5GvZCcg25/3h+h1PUFVLGgVWTv/DRDC9
2XZsCiY73J2HkQm9QlhcJNCOrNzSJ+D9f6ueFsVctGxgTznRqJMnjVOQc/zGxMqX
TRjWdo27b1c7nTYsZwAJzNJjqwEMi3BTvEOCAKjbhEvvthd+C8/oWSEbWekLp7rx
VPDNuDcmLNI+j7tgqEu/otZ/1KjmkvDIDNpyOA7KqYU6I1Gar2xqGfwJTMPmF08X
YqMjuOJfKd0k8w1zVw8f1CU+USm7glsBrpFuUrGcyVoLkESpO0AfaK3a01MvlYqu
+rGvy1tczK4GJkBGBm2KYmDGOZERS3ObzSCW41Z8bqL/Uq5aDBXRckXD/oYK34+d
y2HzDSannD6QRobY2RtKytcBG+m1OBUeDyqYAcpO2vm4k6byPX4k0H5BEqxejOmQ
yu30HjYB1sYyPkugGCMr40eu6vNiwo6HTCBan/8zuF+AxJRTm8JNy25ElNO6HBPK
izqACcXXwh+7bsyzN3shA1pxlY3BD+y/lSbBFw19p+YhlrnT4VflBTROorn6ABUO
jfqjFXApBb2Q6Q5OHIrpoTeVwoAl+R/ByjJW+dTV3uiGz00UQ/jU7J1E8pebUf6a
TsJkjjrMFs1vLOxzZbEcbAwx5DUTYFOFJvtze156VZOP8buPTGvtzgvWtRvUTE1I
ENdZsIBRSq7JhIwi9aPYECDrMC1JOBCwlTYo2FvxnVv5M1C8+9X2wElRgNP6NvvJ
R9tu7xG9Wo1l6oXYshXZeFH9nNtCzfRWyod/PaXoU9RR7LA9cxy1T7DvbX/dxsMP
KA7yVT3UiC0YBoyU6vzlTRyz932eJ+kiPshdVbemCAOucYD6rV0XireCAkPXQtyf
/cXUNukqIgyyVqS6C+Pv1+ZToiRiKu4mW4BGFRCbiWHkkRRtrOeJa1TQgLR2N/fX
VxrXNThHsmxNiZO+VA9G7zZrm4e1Bwde3xhx2Gkxnc35HfpzDylXxA8sy17/1sFH
ZS85MIyTO8O+7BSn1QMf01yRgToY8gt5Nr/W8S+kOOC6jo65CoFwiUhY53neHJrh
ZKPtuNCg4H0k8KZNE+EWGRb+dtwnBAC4TWFgPIVh2fDhhppdiHYYxnUDn6UKiZ7B
S6yCHWbO6FXbkSoroERkVY3rbmNuX09JrY3f19dxYolrLZ90J6QpVf7nnXDFfssO
a7qorXxzZRQZ8H7VXzCLNNMp3+s0i0vyFTeDmlIIOF+san0g37mPWlIU7Q64XXTr
3rklZ2dV4mEXf6jYtlO8QpEk8wFefOd70TUgsPCBqLgVDjwl7aBIl6TOcT7M62J4
Q+rr0RZ+goRwfjKT308HV9JHVo5wXP0VbBUqWmLGpuJzouX18Jm8vWntrvbcKsWj
HpKBSgxxa6c+WmLN6iHaAdzm7Evh57Z34HxLMnUJ61S8WS12K21dUxYn0ymbgx5Q
HVMjY0tZeqXzD5DeIGMUeaSyLeKTK/uRFxdY2PSLHjGxBRId99WkBdDxiorgVY29
eFOwQwgQZza7zJNnxI/TiIhaRj9WiR07KBYgyCccJ9KkphuHC4uIU3iEBE6OFway
gSMzcFml2ARvGWvQlN2xzigHmu64tM6rdvfuJfPl8gH6PhzRIYBMb6grCLyTxhf4
jnHMHZFfmbzqrf1eFI08Ics837vZs6EqB1OAI8YspdsHg5fvebyW0pipdSSc4U+r
q6+UT5Ick0fZ9eixKX3kyV+shNWsCyhORtEWZ0oI964y1B3MAnbO7ukKq3ZiXI7C
dpODoomOzY1bY0//NkwdsCf8CsBFS3MRK5lXzrnzOeg6B0z73MqABL3r22QBM0pU
MGnxhofXgXUNmPvoKtWO05CWcbtkmpikVY9oKL/2fXhZ3qHbdRGK9Idw7KWIj2VZ
0rvua7fyLfk7nMvOaa8zevuGN8thUL89EdofVUn7oStlVO8AReRQeXxgjff6fUxP
Cr9FsZmIF4DUZW5EAqtN8mD1un1d1igoNkv9LreWWVaHl/tHSz3eykVDLotqodDC
3+7c+BLPlEmq3betx2PPVlNQEgDTTF+KktZlJZ32eNNmSsHtD0y5GK+N2eiBcQ11
LvbHGfW46hrjcx8z9Dq3ivsvCR0QbX9AQJAkuNRQfe1eDACKFrAN3UryvGU3lnfM
Ny+11oiT1bPB9GbrY2dCk7SRl1QiZISQYR3u58dgUuljAJlVEd49/Bjo0Z0gP4pi
AWBwHkcZyiqFTqCFcEmbPhmDFe6k64GcvmQr5nHAltFX375HaQzQSxu2PceWmXsj
h986RXD9rCEtUis6QFdpnpBxT5I7oAQlS2SNiSXOKKYSjKHo6FNoGMqeWqBzW88U
jtwrjPEwweqamj+3BAsRmCjKVgx7WmosAmFS8cFb1C4uQKADAgBUfkClVlsJ82z6
8VliEcWbxdHLBDyxaEUTT7Hxe5Q2i4Gg5F1PHQKUnWZNnF5x83gL6Dsg7J1bbIms
j3GuzEFWj/K21ParW4D2IOOqP/wsbaZ1Jd+uDolt6W9r5H1FnGyFeyvO6NCuJvfA
n1jUMVnnvdAi1zKGCiQnEy0sSm0PptdynIRJ2KmgvlqRZDq5qVbcLqLFpIxLm3h1
UJvzuaBx61buzMe7tqMvnSEoK/3gNZYwnmiFnUkYiqZXwj59XoCYTAMQZPd7HZbI
XE4g1VqpnJWa2tBhpyze7UWyLYeAZSwZJo4gtLK8MQYAPmzFYy5OVvqI0d50ryS8
7fy2nMU8Pr5iSE5VquKGidkZtKaDPGCG1s/kXeA2jkG/xNYdiFDpGtGW+DwfH3wD
Hp1ZVUjzhOgsniUbiQ69hxXFOHQ/s0TCrU45qx+Y/JV5hOQ9zM3kjsi5wCYZpwrA
9eVS4bvgmPev1Shq+O9//mJu+hdVP1m3wxhIHWJh2coQeyoSMbSss/QkLthoYq6a
SU+ENltGx95CKuuXKIRGk8dlZS2SrEb4dm+8Rjyhc/f0TULhZkJFpaB3Kpt9zBc8
QS+HbrbLTzrS1nuTgKbKOCo8/N1fX+RzVYdJ8xCpRYaT8raofwr+VDAPPLTBcHMl
FQbgKAvclnjlQl+goitT8WOsjCrbllELbd90OsFRxPf6j9+utlGVGq/7K7NgyIJ+
Ww7Eij7WSIJLZDQbHvyElBs1jUXZP6wt8jVDbJc5on0UxHbPOJ2q2/cAMU/RaI6/
HPqMVYpLfB3NVc9BzKJUGdZBaKeM2u7prIQKoTvlrMuHyQHTF8rpd8zxBkISAxX+
IdAr0kUhawyY4H3Hfeq4zhiidGru1vsz4QefLs+Faro28xdAOLH+tAUvlu8Teeix
Uw6lkK9voJJR8xkLMjc6nRY5S5nVJBmVts7Vxn+lK/MvPtJHDsiOuvZFoVB+EhLt
9V6AOmhZsMau7FBK2dfE3+OT2mlcwgX4ibxnQEDsaTTH+UBJc4GEghU/wRCCgjED
3UgMH/eJU+9AWA84YKF4+Q8d8Ra20H4Ry4un6lzX9B6aLCWsIMd2U78aD/EEhBGP
h03MCGMGdSNKBlFJEh8Qf57Kh7SG81wglfOJT+weaVWPhzm35ye1MYsLXuLqh0g1
2l7d9e1OqtLy6UgnghUwmQz0b+24xOjYa/wP9tmSWxeEIDpTPJGXeXYJNgqXNRxl
A6rPh9U9oX8gbkcFOqdcgRKeWZT1y0XqeWUfy/Xq/6k+j1f/IWUOhcfSVnaPQYDL
Q2bm7A8x6JpT+ZENqzFb4i3oImQ4qNPaZNmxxHIyI43Vu982zSSSlfTlwv9Movcv
31vuPvxncU63qOIHYOwYmumSCC/f+8l1/gOFKROvzrTpNmqvPKGxcV0tLrx0Ul0j
i7KcweFQ7l20MSy9Ci/yQwSnAcrChKNJ25BX+RwnzYvS/xYGUWQekM6ctJ3d7WXo
ERno8j67N1QtmFXRInecHCV+AnLLjZdJs9gTm/eFjGkUQgkjww622n+UW9vKCQj/
4WBcjtftyaynY5jGUgdzqtG0T+04Y2gwYCAVtuPo0eBnEjPrTHuH1Gqw/Bf3shQp
Ann0NDLFDF8zmaJKpU/1N8F2aj15pMsW1gBiBsa57LcdJzjPrGPtlwvNEae2Je5P
Yw7WZtE69kNwB3flbvDCwPjYrWVo+jFSzkuRCABik6ceUo7RXSgYOdp60b3by6U9
kOMcCk1YcPa4MawvRs4cG/gepj9eORVAvLsxggoQFFNflUNEKXwcCNjA04JU+bB1
SeZFIoohjwL5G3FBb8k7vKNPpFafC3GDWcCCC5VIXo9IjRNr40nomH9HSra4z5Hm
7Hok6p86Bz5U8DZfmLT7dpkpi5g/Zwl2s2+o1UOIrcbWJnVEAETQj9I4lm43aI+0
215POcbU+GbJYsKtbu5nQ+DpGaLJvLGK1G3JCqQW/aPYMvnX/yWFL4XxP6LIvvgJ
ZDnC7wCLTVsddmvq/1rvo5A7WVnqkUet4325zxUQ0OuSZf1LnGWMonX2ZtRULVf9
aLmtkIe3C5NV5RYy+pG/Omc8yDkZdImGfTjTfTCf3enm39e1cza23ghW8wrwU2NI
6KHeqiSzCu2jjRNQZRrc5AIk+2Dn5qPvGUrQrPaMHsoUcjRnlMHrUeClwc2deyPq
Vv9CKe9Cz02pmyuX565P+xf06Vu5M0WP7DKfpnzjf/HXRkbf5MpPsIo3RPjXtuV/
6zIIHRAbaQSX7vJBGi3ZkOW91IOlbsx6mzYXmA4h6ixX3pl63qIoGSGwpmlsWxnE
2RrrXlKNiqtLL29bLmrp/QxfsIO12vKIeLZLs/SDSU/nqQrDHsImWqBUi5JJGNS1
zF2EDpdOj45J5+bQZtZfax6S/vLWbhr2WBVfw07FBFP6h9N1VELJbwAbRkUpSTUb
imOx/RcfzhOyYgv0pi/IK9yV8M8VexwehKWg74x7N6sQPYiJ8jXNfeITfbd2W1sD
2kI5IUO7/a6Be1m1M7hZyyL7EYMVH1LxK7HO2YQ6hkjYQQIcRpuh6HkK7MQzNKWv
RNkFeWA1yurc5W7B3ib/w3g2I5p2BS/655R2DmtrdTlkfWy1ASExgNNHN9xIhdl4
Q4QhXFlM1Q5IJFOrOttMMHx8PU+9MYgTiscVhkJd5N36VBMPMJ7DJi8AhjDQRAhp
ItnrxJHHkOzd/PSeooUqLdtPaaClp/zF34hGJbrZrNIM4TjEBU3bHtvO9lhw9xg4
sxi73HUpBdUQdAPyR/5CLLFgqECT1nDjUzPpbC1XlY1ayS217McY+nTDZzG/fYFx
zmLw4PGEj2lFl02D/M6keUa70+Tv2uZOioVHl581PlN79Z6fm0D6vedn3MyUI7dt
GGoYTvOI5zkJTwkE3izGR62dW0WKCipeVoRyQgVFO8naPAxHS5JEBqxtJqEGCaEe
GltMGH014mmwJvTxIFxWu92MjuQ3F1xL54eY81X4oLQZgPds3swEAr42zT+YhR44
vFBK51nYZkXmlLiNjjcW63IeyybZQedKL0PqHkACF2ox7L2XCkFSb3XMIeBiljml
+Zd2GFmydUmZNJsdPsfgRSqaUHj1m8wE4yLxcQmjOsIUqJia28AAjUzw9ybB4jPb
5oXxRP3gRxfaw2rFgM/8mI3FSBPRh9eloUYqmtMVLIKsp8Lb+C56+gok30c9diS7
T7jTGaIAyhPT8/fOIXPxqO7CpZGupzvhN7K493eZ4Jb4jLudDEEZYK2t3mmWlG7o
+8YnDBS8b1Zl8d2AahrsJj4j3Y3ra0O7du8xIb6cElJfyazB6P342vNaL3bfi0kj
FMm5RS69/qX0aAaeittuBTl02D7sMk6qiMRe939juMHtqBb7mQVZwWqYVXThSzHQ
2DLWcEZNEwrAv+CIk3e2jI4iYTa0wBDLXncuHcVqOP6Eo+y1noIARsRJo3WCyLn0
nYzON4z2g5+h0l+m56gNjJssftgIwf7UG98s57Utuhq88ZPKQVgskLoA7egF8l3Y
2LRciyvRc6O3TIfvU9H9VOk8dQbS/nmNrVDb282vHYYflJlQZ52haSCWEGFB4X+P
6/hhj1typc8m1R6pB3OSwGN+fHO89+iy8ihLmQNqpZcsyjOD92TdjXhMLZUZBGrw
3GfKRJDJBM5YIRmU3nlRS4vylZpjM19g3XP1+q25MIs81cJjGKSzpqYwOwFvNC/c
UFpGbDlT8uBtKUJK2KN536e2izRTybgM0/DlMIjUkFnUCD8H6Yn1MNr7S9nKkaz2
4PxM73dhGQhJzzMKx4088LFA5UflnFTCxcQW6q6QrNZXKbzmR3h8yvHUUrKs5FO1
N2v+M7qUNLOYDXVFyVA5OgkhFUAFaL++HMBdIgFNHcxVXmXGCJSEPGxMluz9/Zi/
8L4uropKE7ZBq0/3iUYzSPRLKURjuXQ4Jw08Jrsz9Cgbb4nRIjvgQCQbogF2skig
os+N6qTZJvuUvG0RYJgEV2T/UkV2vWOPIDTGOeqtaRyrOlG3dbrE+ssBDOXyDsmJ
+r9gK8QCykE7Cxj3etRGI5zX4dEHx4ANXI9TC1DYyO3KStGP5B4thbsDOMBtUfl1
bYBQUQLejX5HDb3JhH8csA3dgo4CR9jQ/p7qtueiX9D5ucAiXSBA50DWX7rci6Bl
Vdldj7ej6sWHvePACl0ZdSVpHytnjMsEupuEVG4X9+vCRLJFbT29sKB+pLl9j30s
qYCDpEftJGP7Ten5/M/hYuSW/6bQwdFt1rFClO4md4mYSntZ9oAI9KsgTHPc++Za
O9qG9ndZ2zMf3FVoHNZT0S2faItITjT53+vd6CuE1GTsu8mBIMdnje6m5ZprpQ3z
5wyc5mOGRoIFJnDsjBoVXrbEY/0xheOCObxEcn5Xk3LVbFtuVMljoB6L12HhorEq
m3Uc9EB573foDLeUXX2P/zx8vwFjBOUnmqE7WpMqBk//O4D45Vfc8cFlq0eJHvlC
plIjEeHuC6ziHyNQFf7e5WOujMRTuqIwJqDHPfyO6985xBtO3WnYIjqqYPmyOw/9
7/NrIcx2yOz4ESbrcONxv0pJ919n36kC8whD2D/08Y+bmMlZqEvkvB4xFwrT5wt/
kDNTpgI3CzaZbSry2axhjCMh4zvWGJTTFS/gUmdTOidmbExU8pyEIeGpjTQepg8Y
rORuodwugk3rtqmFN49UPDZwf8e5iP7SeH5ZKNctW7NDWq+rLrYjyS3yWPix2DAy
zyYQ+9xt65ZJFd7L7DhuodAXSUe0M/u7zOUdGSxAuyh8TOFnucUAjkKopU8C6Jow
ktBG1NdgXDoulSuTDOe6c70OfMAv6Zo7emMNA5J+1TA3bwfFcdbxrqcOIyG2rxTp
tIDtVhO4LCRf8VPpBzDBPYqSxCh36VynZAmSyJF2SzMQupWUNoJexzkRSm6vx/xg
8QttQu5MFVVHW/1aK88zWkKU0uPpyoTba99arT72e53bWj9pIcI01jynpSz4WR7S
HEJb1XK1BCzHXVbu4IofZJ1RxaCy6q4PDFP80q71s66+Y7wjaFlcDXEgWARCFfZF
cQt5jYp3bjnBLlPyqiPCAGjjjchq5mS5iqqbZeqqZZRSNtAkCTc3wh+jZnJism8Z
kzr51xa7LlPv+WbwJPwCEdsFFFkxnminweiHUv1MLI1yPrlMQ4ZwEjx3eG9w7a+F
geXQtm9qMOsNLiPoLT2PXdR9nbdB9s2ps1/Mh30LQiBRqqy8+Eq9lVu7XnzyprAX
2pG6YYAMvDL1p2v8PABOFSpkoDSA3JhZO6YLDCN6oLUxP4SMp+PAlD7i4JLfIPIw
1WCg8WQnPXDnXC5m38qM6Ura5mHVm0m42tIbfbh+NTCM/YdYC/yGUr3No9EAHMk+
RwxyzpHevlrLE5Ihpn31vyBUy6mqru0PSa9T62Ms9x/BTjR4Fg6nz9eKDpnVpkB/
q+5/wnyGBIHnoGLrXhe2TcvGpyi6dOLIBu0RcjD6zvDS7AOEZI1OG2GWynN8eqRO
LxpUeQqpodKPhKcLXYbenIvzXT0Aj4SlcV2gCaDJqqcwQoA651FZnoFa8ECsTx38
Z4QZ7mvDhijTHqKriNoGIbm87pOfvAzwneoHx6l9D5Kh5ZNSQ/RlD2n9+4HCn34N
eKXfKkILbQrCqNPifv0rR8xsRq7DAwnmSW8Kxk/WL0XqYckPcvNp/I5vjr8zBKoQ
XSc8eYMEQe+zxQhUJCdofgln62+5i8PQydvEak11ro0jWWrV/UiAejJmbmv4sjHk
BPTet7mYXMNu6I0hai59ins2woOYUWeJdMrCs5u0VelIIJu4/K3A3SNS3Y/5d9YU
LfizEd6o5RSvmGF/G2Rj3GqcUMS4+7nPTF4ZrHmjU6nqyJ5oW3jMof54bdZGxTlH
OsG4l5MOZ27UZWAbcd0NQGavLSPrmHJuEkMP7pc4FLhri4FxMoRY/J1D6Jl/IOsF
PmUJEKU0KMxkhMWDc7z797/APTZBNxtKHsl4c2uKkg3xBR1gk0mSKmEHhyxNdNW3
8Pat2xNdneHWjhzbACO5+rporKrPaFVfiSXFTSOSx93R4ean/BwMhlmuIouUfeU9
eFUXDcH7yzkJ1h3e9xIEYECkB8kneHHvXy3j/bgFn5fFT8gJwWbaNcR5GpV6yguM
iifnkVapZRAHXWnywjgP10ZOBZFWOOs4ZGFL9ZlsNBBBb+UmeKePgiV+jxtskUN+
JwS/B0Zwp5Of7noReZeiQjHhMXNwnj0fBFkDTKOgp0kgmxTDyWbeWbPoYHrdk77z
pU4Fm7NWQ2fyg9jDV6NEjUZaO3fSBNcOg6R3OwNdG0xFAbFQG0CzZFdrMCxGuKfh
LrMFl+HFXoyStnPLbXJ+zEsVNgYEDQVaHSURQ1F/mmmzmh/xwfs/p3pV5OMbdg4R
dtR4V9rWdW5+ebsh/+40M0lGM0HBnA4EhsbCWNYCRBwY4utinpqybUm9n8LFYOvW
zIt1P9sir5ehzrgUtdJ4L+IvTnebkbUa865n07Db3OHS7FxpXXrHqp0+feiix+im
DHVKLGhtuGnapUxRb+bvytDtB5yhdr22dEW1s+h52g0I8KiCBHaMPafNywCkl9Ya
RixRtSeajmJXkql9SMycxPzZWUxGRYZWukwbVNfK1JF/QHM6Fyygi0M1GBmowQGO
gyFrz6fWa064xZrL7ASL392RVuNyS5Jr3T9MzaTmp85xEhFxaDo/Sf4WUerzfE9P
Hbx9oeJxIwvFWPyV/2tVN9rGiWrUu8wiE3FTsJ4ha8XGIXD9CofhOAAD6gIFM5qm
OOBmDaXx5sxE9rTUOOL3oKxtGcIxCL+b6Y88nTYCt1uBCasJl5+rzOYue5MMb2D5
yNsMc1VmaMoCYlhX9xOYbKO7cKu24c2T3T/E1zQ/0ysNbbyB8W+njXuZkA6NxxWM
LtS4r3eSY1kbs5MzL+h9CZTtKqae8ZEOE8kuC5KKLmAeZ6g8FZlTZXm8xlU1GKpM
x0J/oWDvxixSwOm9fxaScBaXgaywXXvaJlOEiRxlMHkV0rXxfRev8k7Iy8A4Qa1J
ivLTT6xXfwG1ilSUaVZHLaEP9Gd/pEOwQhQE43QPlOyuJVxCeCtuT8ljM/qKK0ee
8GIpLtGGHmHQCS5WwPCjHSm4sE6BrxDFJKwe9CHPpAZ/5T99HTAsjDbNid8DtcX7
2d44nN2a/cnPtIJECmXDkndgHL1oav2icMQ5NYsOMaLRj8zTUi7NsWu3gaFrLoIt
Wx0g9kxjW8331nsIO0XQmXzsUa0/jGw7NGKQR3wFc16RyD18mHuRW0uYweTzDsv7
60e6p2/6bZz7Kco9gO4FObzn605k8rz4xxnuwWYwMXPZpEUnPz/CvK+PLJm4RvzF
sXAwvPro0jJUdopPHZqUceiy9gSci2+V12XxyRy4/SqX8bRgJ/iIBUzTJcTYfGkR
0ldVFgZTnIlVIInPkpBXsNaBAf7m/r6zcdfldJVwATOmHCkOsSxXgbELgqh8D4qq
w3mGSzU3P7uolqrcB1jSz650SLlCZcR3uwnO3bc83DUNNUCbax1nNBPn1VTrMZ+x
eFUfs0JlV/TPAp0cP5hX8kZjTIkBndSWthFc1eTRR4ugvRYW0ULiWDCwyTGDrja4
Ait8fevfBlNCLH3rrAFjNZ2WDOesLYQwK/7jHbKwGcuLOF2a3SkG6rnx9SYGCh8M
wigrMvSAG7RAd/7BxcwZnVpxgyp4rUYV255IZ01kYmJMtHCles1S83zL+OOYxbMi
apqZ8fcDRxdCdIU1N73nl48lmNRl11shyW1vrAm/2YHiwRPzR9H6G7/+uYXV6kQQ
1AsEpFhjGVzpbyRdbCIBZu1qF07na13C5+g+jbvyNyixg2xaxszt5trg1wT80gLc
t84MwjPG7cxEQ2H2UiamcuWsoCT1B2JA8sqScRD0lPSwknKq16diQhkWxybA279V
7XXwDbaD7oa3D96aPJ3vAzxkasoSJoHRmwgj2vGLMjh/IWH8luqqHILmyvz0qDAw
dyVy2BVipNRfSBcPePPtUA4CSm9/5Bg4dvpDTKyUrZhEfxna/vEcfna9v3zKbOb9
08fV3RaOvnFclby5vKV/QVzBvsWtyJNHnOo3XXPPVnKoCcwGgD+hWchGXOJsh/Fw
C6T59MjjWAofRUaQwJqxrMpbb2QB27bpOEGT6D5BywAc4anBwfhbBp7NFZUAOsT8
3CIhtpEu9ewXb+12XV/I2l7cujW5Po/MJKAXpvPvoQzN6llwZsdyGGElYht1V0A4
xctkPTTzvKUjJeBrAjE5EJ+SwXFAV4IJvwXaZ1rlsEQztjjTy/IxCK9hbU8l4p+6
cBz6IMrg007sH2YNzuujKvVo4kIsyuGJ0pMVC2peVD4A4CDc4iWIg59elqEDhySs
PUaNgv9wusCJucRfFh+Acgx8v+AWQtGbnt17vfCGIlb8wLOxPcwacElTmZqoIiDE
JGKQ25J+X55Cyt8ooRGr6QWdV2cp59PGbuS4XzKmQ8W3cD4VtxklmfvNcw95UNJ+
o3VxDvAmqA5o+msYSHUAV2DNwgo25as/ouor5T2LBPKjT0h+esWDOkSNSdnfvZan
nZkP9eNU7xJ6GcHdGCoNC1YsWYFT3q4rWBm/gvUNY9ttUpOQioBwhKlLlY/af/82
wjEB2ObD0/35No7u8p5evNapcIkNkmG/2dQTnvVOj20Eo5kK65R+j3PbGcsYg69F
sNBSIPVXj4bRHbAD0sh7mVieEcrCvWHyENA4EzhuG+7nXqAKdRq7Bh0jkaTQi0ee
Qo7RFOEypVFb9xagP6SB76iRzidW53fXJcypFV8aBgpthslv0xPFoF3HvKgzJBAe
2DHKdILAKTJmerzMHTVvqzvCjbepMKi+/HVUESh0xwM8n/Owo8MWgzle0aUxoyp/
V1cH7a3BgCtnuF3/gqehY6dM1MHNroQiWfoCaq0GsEvE5VSFVOwVgiri+eTWUdEr
9PsmKOYs4Y9dI8mvEy84TizFtN2CO1Kg2+j5zjs+iLEcbyitwb4OyqG1Uco04zho
lGUTv9d74gLZr2OByKEYXj7YmhpQnfVXIbYmbAredgHjW/cIekzRUvdmkDu8GLxG
gnxuIopD5HfzmqaqigXskZwzzKKyMbppNh/5n3Gl28EQ7FQUX5bO6AyNXor/Xdqi
9XJuo4Ulmf4s8bvpLre3snw8z+BYcg6zaMYIY3SyqNUEwuvTVI6PAhkPQgct/2h8
yBJF7S3i+PWM7CvETQjxoJ5Vyv+kw/nmw8g1RYK+BqFjL5TOoLVURziC0NfRQOhP
eQtM0SFVWHwS1NYnb940kzIGjqLbkCPaeIv8Y8E1uANg0ZELEtmyeo6CukSSyOz5
r+ZHb7m6yen6Kj+o2imKhWPAfsjWLD2kjIzDJaBZtOse3visR4oBySkoHb50KaGZ
3hG65q+VvZ5vDSLFXpKsJrU2ibMYSE1IvV4rUhjzTOkd2inlRyiXxdOi/fUejR3d
PZjCILXJTkISQ9IPt52Bg5GI2DBtZadUZqxGsF3tczf73g8Td4Br2L/GbPuH+pIk
tN6aaETJ/BIuOY0+QE+5QglISZXo70BbdAGFDFc4SKjvu7nk5f+c/YZ/eIgiRO/x
OJAmObhP9TZdwYjz4lFsOw1RoeD7kBUFKcoKLoFEVAMXUOt8EqWiJA7UGuN39/ag
xB+r7ER9+VcTXOTFmgnAyTFUooEExw7SDJK7pJCbCtcEafDLesXcuLWrPvoEh9R4
j1D+kuRTgyNFUouaYD66Mh22rLcYFt8H9s1MvCLDnvk8be0QQoaB+pyUSrt2XQ8T
jo6j/D/9iONuHpzCw9Ag7dE6IfMfUuNgIr+a5jtWGYuxNM8smL1efUte17YP+3MV
IYHlta3lyW0A2YabSgvCWn8DK8zrZ3H8qz6kfKPIU8jCa2ZHuLUGgZbxh3Cd3+B6
8lio71XXFsRohbaI1PEV4LdKnmYdFGRo5bfmnDqeftLS2tGzKKwtPxoFnACQnsIT
VAZkTe+bkVLfDQ6AowD+TANJuxEMUKn1yQ0IvPmHGHP2bz2ee9j4hx4HP7s2NZmJ
TR57Y4zwO4Ws6ceVwp8ywAjgqMhHAquwsYPiJn9lagriUEJs9Zv5oIThdgJqwWjb
2HZdwoHmMkbkJcuZXlAgzbEYAlLWD7x2HEhjeBqe1g/DdKRQ2SOgofVcgKm7rFo9
zQrUevuvaCk+35/RKlLPmnSIX3xsV2/m0/4L9x20yQvlbKrLcrJTIzwGB0h9mONC
fGqjhVCYuCuWEt9gVGt9CNBsRPKUBKFKJKYWsIo+Cz1fZMi5aZIz30Q1IySeuf74
cIQRE6gTGsYN87w7Duwac+FJ9PSGNdyK1jew/xuUhlXWF4OmvO0pxXyxbFYRy9Im
jBmuXCD7efjZx0OXtGJyBKGZXLaN5rYiWwMD347JN/qb9P8FaknTcYU/rNKwDgrq
UL/gzUuD10N2kwb28ADvOWg+3T4BkLS/RA7Jvov5FJZ2RGce4TY8cwz9Wtvr++nQ
T83y0FvOXuBDaR0Aw2hDRYvyq+eMUcPe526/S7gjc2k++tC3g+FmR+h6ZhIUCLaJ
K4RifVzTXPDJngLb/ByLSxQZKoQI3HEb8LLYCTeo+LRT6CBLCDoI05C3grT2oIzk
59hOr6QMA1JYKItbN1Bsdi6+P8iXLHunShZE1dukEt37I2WAj1QQImnBwhEC6P5k
SnOw2TEM/JDPFJe3O/qRBZIM3JqsvjGYYa/XeE1OJQajpkfzPO4UB4Av9hmDI9bw
XzvA+2DIpSIO7axSZGRGoquZqchv4ijq/QzwnWq+F8a2GWWtx1lsf/zM9mdf7yHJ
5IRJiK4rts3WoCoZwN/jw0IL6gzkKwFi4Jrayerlfvg3EFta7MeLfHvSXzBij+Gw
3kRT7kj4vVXau0OflDSmxFGzziB1T5Htm4peMdUj1njy0QE+dN/Eyo9U4cdAlUB9
mcPwUTOSF/onWrjv3boacPU4k3iSWfZCV3/v4FYJd8P0T9R8s6ghZXqAVNUE/xBz
SogkGKv5EzUALbKMz1rtKN4ty85+HAnBaOxjVQ1Deg85rQMt8Em7Yh4dRhqKCUvX
FlYX72VI91kIEox23XsJ2qx1v3riEmkW9IitioV+tcfal5dWrYOW0/s76IdyySTO
IdGZiFuet+gwJgIkt+GC1BB9wEhVOvWR6YklHfuWhZ1A6QrHQV1ReO4rHA8yxvCV
71QgoOmdq1Mk0NRHHKppFujdkhaF0/ptvnwjnH/pIs2Lq2l3UGjUPmaIs5mRq1VW
r89JvkRanmI/LmqIoDua9UJ75bRMEDnUjlT/mlcV2kS8PtywdstrC//ksYoFMEAq
YvskneNHsS5CwHcwN/TNuewAtnl78zqxpvzNaTaCNftZPy8RkdeTH4hNgwiNF2Uo
upmIUinLaZRiT3Qloh+1rBtU7uwKUNIV7b/ZCH3K/5cI9bLA1IvcEUCJttkIiZ2K
47bU6sEudnwZ5SZ0mmvcHPFd4JFPFv5d5IzDAxDFJETYZ3El/iWN/LSQPBhkMIsd
Jq1tLrkO/cvw1ubpMUZIH9pvgELby39swR3MOI2ALP59gm+a4xQMgNWLAIrVo1Gt
uWfIuVkBM75H4HI1MiwkNRDGTn2IDeyTGve6aGg6MnTwrAzqS3nblvwORly4+nM+
GjoYtmwdV22kFxNZwfF2BHDtmNU+p92iGQh3IE53tf1TnfbONuIjls1sRJKTrkTL
p6NLL5BASySsVCnkwU1sX2eglOISk4E8LoU00SLwe0xTLOHaMe8O2dl7kiykgA98
RbamesPeU1gmgLj//ZYd5sh7Ep/Uyo15ktpEHQ5aNYFH1A/AjuEt01oFhHFKlynp
ivwQSc6ZV4crJnJdUSDtKAjL5bYyLI2IUxAwEm3UHFFDHyhtrm3rt7DppIHqYkLv
tJ1QSlHtlX1bcGWDcF2nmbS6KMoVQauH3sWJ9fXS5ACV5yqtEGXM4IS8Ybrsirxb
NX3mULrSIG6p9ixt3Rfw9veyy1FPKU0Q/eeJbNlee6C+AWfcSS3RGv9XkS1AobIn
Ph3cuAfcVHHGCCMTV/AfetrEmVFTPx+9CGNTpw6YAexGi/SUkGts5ofr+dlpGTHH
YIR4KMNXtSp74xAlpZEfbhtGqUFK3j0kGQkvGorjWteqJ43Y9ZFIfrU8xtIXP+2/
5X41g3jWTQXqvFp/3KlN7aKtBI795XNjPbZV8ZxNlxxPf+f6GDOd7NPSLR7Dot2O
6J+/6npyLvzJ8MdaVSw1AJ8z/wjbZiGD39tItX5EFNx0WAe+aZ0cHVfnPSWeJlPE
Ix9phv0H4amxzqW0WYqjwnMtfN9t7GBfD3jMhXM7bHJDkZTFdhNvO0GrjCBpcBB3
AINkTeKSoLK6PBK73Cn1GE1GhS49kejczY+q7U4rbJvWu0HT9lv+pJJE9V+oiio2
q48s91+e6eqI8FhViPEmbMfN/L40n0mFEJHHaubHJvfH5q0Omw4k2rr+Jd1UITJh
a6Lb92VJ0CRfxArn8vPyI9uni199Lp44Zf1FgxWo0jvEYPL9OtZFSnZsfL4o3Wcr
RKOSm5WJ96OPySTz/PVCTgs/x/0Ob7f7PaxDIk5pyY01Sj4FeY74TslApXbdAzdR
5oXjSYty0UkgOI8aUvXIJcZjxOtL+NtihtJEnvVokZjrDq/bAm4hsWAKkCm0gdmW
Bz8ZRdg7v5XJaNjeSldj8PgBzX0p5f+fvLqbJfqU4a9XM1XFXVuVu1VHiYYVxNkx
0vtVE63a+xtWmwAo78RtvX5ABAe1+wzrNdDn3SCanOGebxlf3RJQ8wzFuT2iw5M3
wVOLNkkbWxcm7aVFt8ytAbKJDG8Tx1HYsrzNWJu8xwng6M+d4wej24aKjezAx4U3
8GhvFqnUOFxBm4WvMQSo29rP1PimwmMvu1dYKHXoGsMuDU73iHCxSd9Ed8K4JlOc
RYuwS5gKOGx1u9hfoTHdcYVjSAIeF6ac9JiQl3MRtiZUVVWfoMuA7HVMfqaSeosq
J1hyImnF9UQwZOqCZ5H2sEkZiyqdVRpeBSGsZoa6c9KA5vHZWU0wMJfXBw5HsFSK
i/Q1MXhsfU2Sz88V7FYEjzbPPFMdYvrIOvhQPnU+jmLa8PpcqNMGAVIChZdJWygD
uGQ91/cyExpDFBsrmMPqJiAOyyn9NwSdxqC52XbvhgVMia0Z+Pr/Dp6W36zYUrYx
c2bGmofd0ae0X0tXfEUn0yW6yjifCnMk3G1Aubw4b8N9M3wVYb1pl5d0NiudSCki
JkJRIYjrzv9eCuv99GtAgBgpbzNb/KcguJo+VS4FBuex6cZQoiMiFnKZy/4wIxTl
Zgd5FQF4djkqx0RXqIdEr0n3wGX3wNb4U7ximyZYzwSYisAegIRQ3cborMpSd2Lt
EkCOf8JrWSLPvOzqsj3EIDu6wbW/ai6FU+HrbpFTHRFGR0ye29L0ryBmuN3aX/rA
kh9PXBDEbF5AvBql9IZGi+3Ii30ioWr1sfuZSiOZ7gqSQieQTaZpn+37yFTs+j/g
16gTg0qnsqg0LXHHumi6j4VWJCgP5d/GVPGMUkjokRd5sGJGvbfR13/3OHHpBunw
jMNceTU0KhW50jezkstvlPhFdsx3YZUZZKo5Aqsk8P9EdMKjjno5cd7Mutg2nj5r
PCiYrVNP3lfUAShkTIZq36ENSKs9t1NfLOcfMkBl/AaWT0hJKqT6sdiH2wPtQ5Ur
JrZX1Yz4mvQaEu7brozcN0jbGkgB2Ex4HjGmcMq+Q2Ane2KrREJB1PF6kAahR7DA
2YrdtNhI5K39H0ReWWN5LjhrsP+ItMvGhgI85qMAilNaHIb/Go2TgYcXLLPQMyDx
+PnC8zjBomS9m3v9lWRWSZeLyJt80SJ4bxAxnzsT5F4746j7dtc8JzvuoEa7EuOS
lrU7A8chXCx93uAv5/MX3hD83kAjKMd4jz4523bFExZVUv5eqSn0SLLICHoZofDJ
6pm38i+ORbhnpHnCKeSlyvwlQSbOzOT9GqXk2fVuvmU44FvwnG4S/lGWZa1OZeBb
C/sclpc+EBe6bLdiq6fLTr6itAHh/W1q8SH5PxL6jkQjy7mbCvbjUoUQux9uXTwc
3cNBXcT0kdhQUhh+FpH/h3EBKg0n9QYNxTSdgHlGpM784kMqANQ1+N46rXM50hd0
4wYIbI07W/YGhURHZYr0D2kS3vzpnIAR3PbE+dOWccChFO2bbgzlA3RbRG94fjUA
cPHrMFciKNNgESnM7kPO2O/XjUeQ/kqjUhb6k9R5mDRkLARjAMkrciVyju2ccOWS
IPjMOg76g/5qgA+VdavJjWeo8gOOgk/T3KnkyQtZSkRf/6Es+FxyMjJ6RABoRmKX
gADxzMfMNoP0WuHet7KBvWAyFyT9WJ/7yqN5vOii0x/5Pbo4CxGExiw3e8IiPCxY
QyBjb8MYh5Cfx+7CcWF/91s1JPmQ9vVkQim4JhzD4k2jNrx3H9TBFup1exSDbtF0
Qad4YJqcEMlpbuDyeEm7f4f2s6xbP3yTBB4AI4bcR0+zlg2DMHYGfmsRC7YJZQBh
h8QR5F2UnMwaFnU3QqMQCLiPEIJyhYAI/zGBPJ1nszD+UG83tJ3SmfADlDQvbhV1
S4NZPQIKeeAnk7PtYnBGUpnSWIHvskvT3mVRMc4Ok6/htImTNwsH18NUxpRSfP8u
tdkfVo9gAc+kGsiGa65LRrx/Er3tSU++WsnxYMNqj1hWruwGbTTvDvHrHebXZpt4
2yQxxUX5Ta38aFlT4B5lk/8k1kwU5Z2Q5EBQrKuSJZHs8ijZHvIooKyRWKI1GN/l
qwO2oBJZ0bdPxKvi5gZWUfFisxRTArjclQ6+KDYPkWW/UooWADEj2q0yX29rQVoa
xiuN+CjbGhDa8Y/PfqnF/E3Qn2T62W5I/4LNhmvUHXL7X5xWmvbVqkTszGPc7xMq
D5M8sLwoGCy2nX8+NpUXtwauxO8OPBIylpg5ra3PcA6YVU1xUjdtCzhAOFym2bDw
fYwk4/t0GGMEIINuFQocBw/WBHatuy6Q3EjAMuE1NK//hCHxeWrfVL0AEq9RseLl
3CEJbe9OCt7rU2IHcG6P/S2a0wvsTHqNMLc7bDbWUUUvAy0YJe/eyu3FAxJW/TJL
0hHCgwtJ5+hnJsBuS+MFIKD4041nRlKjhebremDjv3+TiswesWn78ExLsuTMsfsa
8+t+fnq9JaNezRxQzx6ZSwl+vMLdj2k1r1eyF1HsDQT1hGI9wpPUHGDG5Egs/KGd
F2ajPimlM/yvuw9nS/n/6DWLr7JqIK9eaUHW2aiflzOXuzezqkg7n87cuJzGXSnr
FQ+k4kw5LKsy0+tGTemUGmw7I6XvNmkErnKSwqkIIQW8f20Y9cv3GOAoT7yv3fVh
hcfxsFbGfPrCxDTheVaJwrF7zDzRgAq2XDz6d0/0+0rR6L9X04OcXrFDa9eu5DL3
qtndyYDlZ4e+km6V7Fk8Lp7GHLXhfgN84DnRc6umF5pDSDV4jzdxgqs+vOv4RERf
edq6hGphvd6Pf5BKnXaBG7pEF6eUSujkcWoLd1I36nGdVMkN1njXw9c1lRnfadRX
84WMGbTqJqbjMErawvM9O5CmWdZTj0pwzxQWYzvuk9Zqqy0sTcncoFYnjgYyVNWO
HsT6GnXWOu5YN3kC60S08Z1fI06QaFgJo9EbFO2HoyvDZksc0H8hjOsIYv2lvlgP
+t5/u4fior3OoDquQSwNopo/WVSthWqixwEmntnU5d/DnG4iCx89z8wSDr4GrG5A
ugIBZ6lh7wMaDnmdL2OjIqJ2ro+3aEtnS7bG9mb41dWAixTWm/IlQR1BAXB9ftOy
6kzcEX5PmNr4PHesJU0XclLO6V5yxOGsI+b49sH20HDPTiRHYtYCOXZw8dCqXDbd
krUZXkaxbWluwflHJ9WsW13MealAorxeEfu6mA66COzMA93Ej4Ce/JswkOCwHs0J
PI/kdcg8OFRxBdHpoCuhn00jU9sbTsHBRUwngJqLF3w0XsamIlQBlwpuBqOxOYQ1
d6Br4CHFTCDYI6S5IfQ77Ld1k39/cDJ1X6UOX8KYa5auVtSrdNHz6782HczZeoIR
QSTzDuq4+zWhJ7Q4pQU207ujbFheXq8Bs+OjbxwGJS2vddnyUaZB1iaV6MhYXAL3
Fb/4urU0bMoxDWr03vg8n7Otv3mgR9nUZKBPDxRpzPNMJ4+UVJszwONvxA01Se14
lmc81LmxXituJuwW/mJDeEbirMb5u9IFRRj5tJ8ixSQnRsKaYdaemqhWb2VBfuED
geuylXoQTIdWKP2MHyeW5KjPhzldQ76244eYS+OLuSji43TSmRw+g2gbQy7YSeaD
kLa6/YttTH+N8DE84gcdswd39NlG//tsvoBpLLj/OKNtcJFhmzYTlaIm5PeKODJl
rOS/VfFEMht/Qo8Oqit9Sfj3diGzPoBElfvWEyt0TVfQeTfqfqO6ZYD0bdDC+sto
bqAcHMCuMarnmsfKfFTseHASAQaqOviUujbDEdlCPdWSalbE7MrbnTXxCAyOKQRi
2yDPYkrDO4weJ4YqdCyV03OVmFFLw+EV4/DFB+KRY6KvNopv7mbY6cBxOnwwwRln
lcOrAOr5CXT4W2tBUYAtdgwBt9u1XRWbDjj4f4mI0cjdpRl0wVdcM0CxruFfcLIt
lo6hOcKkZwkzKr/VXhpgxuSBCm8K9Gws7lKrEaRgLts7BCTsemgtAfAVd5CEzPty
wR6RBqOLJUchhzu3uVMozEQ5KrM+tIqALahQuFFj2AlqkQoWaIUTO2xFWNSJmHQc
JRPTB2Ce6JJQTT8jdwlWITCWrRcnt2LZLmMyTKAlcD8876OcTK5GMaYfPcVwAXhM
kX7LHRI/TG8NtY9L7aWHr1by1nNpT1Q+lGdyO4BZF9N++LOnajntW6eSJ8dk3c+B
ZP0Oym3fN1/Yu5EZtUdNMmd088//kXAEYvNp8C58wAmyRmSJgBDtZpXMnUKGl88D
rNm12YclY/h3UtUa+19B7fgEfAoRKX8y8IeY7AzbdHBDPzN9Znf7W7TvN2qhihtS
32KtCBcBD8q/lUankLum3prcRVSuMOBkwW579fiPIKihLSnnxgkbEj/dFRvMJD07
GE+kuc9xcslyWlTrTq/U7Ynu9imu8g5bLegkdiDQ9L+/nkJFcxgMcrzD51JiNoiR
zmZbnXsO1Oj7d/5nS2RpXaSKNoC2tSNmGtYX52Gy9WrwS0Wk6wybGZiVM7zGzolj
ysquhjD1hqGfZaXnevedjwUF6DYUEDNRqXzO+TIogs3Fbx7n4EMDzlaw3N26cDxZ
LTlODQT607caDoKWN0N8AIy28D7HNuO27TQY30BGZFPFNTu1ehP8x8OW+3FO4UKB
du37sY6X8MSSRHxAdxaTMP9dXXVjlgV+iIIq3ad1+81Mv2azkPy6Zh4Jrh7W3ZmI
EDW1b6Z4E+Er1eisGBbP0gFq//g+zn2yRLYoza8Y69RVZbtE2UmL2Kd8Bt/BHJbI
1uDSzOn4LccaslbXlddMKUSA7wN5/3ZOdjPRL3T5/7XFg5Or9sIAC4EMcxf2q7Hf
pz99xL+beA6Lx9I3U+oTNh6Pg47w2mAHihoJ6bj5WE4HTQFEp7rqd4PxT2XINU+x
gsL1lz/TA8EGjZ51pmQvqSBvOU9NFK35VQ1hJm9F6INLcXosVZqTCeh6XcAIzlAn
lDUcpQlv0qDx6EFzuiRXhimppPIDPx+2WpxEhDjt7EO77y6TPYuORV0ggqvecbiY
cTFAaq3A6WGmMBX1WqIT2h1T5xlsLziv/N7AAWae0yhi0382QmrnRXLnRnUvZYpi
/xTPYLGgvGtNsteHnz5suJGJVtXX3PT0210ytHSfUr6Ems30nFywe5A4ZeiWT37J
cyQE+krKOWke4FSXmVBzSJOJTL/SY4h0cAc5YDbx8IlOInLXICJNRVWPa68bIzCN
Vst/9WXqzMA+ncQdUjRg9jBj0lExLnafIUrmH+jqK5RPCslP33kzbyM3XSfPYn98
Jj+dBT3SX6Px51sT4zbSAvi57Lk7SbRZntzEItxXEzeVb+fXo6rPVHhgLdoNl1Sm
O2ka1ZwykFpbz4UlB5f7isEjpGTkktq+yUhp21oV30tYLTruXJ0ygFLF/EZgzwUx
lP5COYH8Bh+2jksEl1yhfRssmZ9OSAHJldPeYwYVPgRe7DM4jltM81Q1QW1zDHzt
BDcHVqWbmWqx343OVp0auhnatyyHdapfA56i14CcoDQ/wM5ASQ/qHR5DR5O9Ino9
TngM2Cg5pqdeeNLi6+dTF03sooNCK8PGFPPSp+gq2JnMFLA6ZzpkfDhPcSZqAdaB
SkGEmYFuZ+Uqunutly4ifhudf25EKcizr+J0O+wl2i3BYDTQ2g+ot4Xac5yNAhBV
cisRWeJC1By7/5/mW3WiDAUlLVyNp2KT7kCLLI30kiJbuaZ64N+8Sj2rkoAChw1H
xg99qJlS+WIZuhT5I7rWYfCTjGagl/mMfAnCaXVZ7TnLQSJIcSnHi0zjX2m4Lukp
rvcPl2ulwKVlI5n19IQI+XvLoou2FpUjiN6469vWXDRjfYdwsuSo2Ru+NvdpCOl4
ZUmNef1YZtsSlhjUXBNFQhw7W44gQWXO2f+ZBoEJcxEoSAsFAo6Fulm+xSeF19Mp
dnPovIAlcDo9MP7RAptjVKVxMfbFeQPW4BdjI0AURfLH63WM5NaU4CWd45RPvozu
eBJh40IX8cDkZuJiwA9L+rjH1TQ3qyUCu+xLXk9XI9zyyJ+asiKvALK0OHqIqj9r
z78MiGLp4t6j7ab7VYO+89pNWcokkxx3FVl4Kiw7gfhGKwW8RW3/qUryw4VU37zG
k5UO/zBkO5nZ1/HaO5qmoA7yM1HwYLUcVaGQDCGR6JITMv/9YiZ+6jkXua1hjSkd
RazJGJYNP38PFglGkLq9RyzNalRFv0zIWbpxoHIFISwjKkYokjRDKGyJg+V9XuLa
nfdMwOjsqm5cE8hEMJvZJzFGVYJNqnH0zJt7wx0DO1M8ymcRUOiEcdz5zZUdnJXq
DgKtt5m6/45eDIRq1sMDXzE+Omg7vf9SAqn9oKXJWdW/h7QY1yrjXPNbyZty4k4+
2h+UVMXK+MbWw2tUeCj0sokdejqCT8PIFsUmAgdPRKOVuaCQB+l1PpshsrdwS2d6
sjc1pUrzczl1H/Q6Qnp2zpGc09SQ7/a7BvYOHQeYu1ysfLWDOJ3zAepducrjr1s7
Jx6jB1tqJpzEFjxGEzFQ3Sa1v0YtKvT3yBl7VLFunk/KHgx/wAz19SDvRMU6xN9v
Rys7Y28FwAOBZ4dEd9qBDUe3+1e496fDMD01Cm6kCfm/bRRDaQnZUJNKgixoxA7h
WlV5ikeP3mxCikNFyOCE/BTBgIeNTVwfCN885G/mCLud5t9ndcZ1m+djTrF9Yp/P
eKKXpHMO0ZIx91RKPyhCjOjvJ6ILoAVO9Nkd325D1ykMvhZj9fXnLNvAne2sk2Hh
aMDkg1ZJl+TQsOBhBz2IZHIU7nsOCtSY7w9d8Wci9kkodWR+tZ2nUPHayd8z0l1k
v0xi2xTMWVw3zUdpW4u9Hd9J7gCSZMlGbIgKNcmh0YNm/0DB3+KgEFg5FIlkvCPr
lYteiny6pm3+KaG9YXjbwXsl+2JG5fBNwCeS9GQP8Nr3WNVQ63QnWYvmYDTRNJ0G
cs2DW757eZvOzBNHiJWbLocufkHXaXA1+OnJK8CvDfoaBHgIIH/A5Y0GFiwZWupN
LP0Ff/KMuH/PwVl+C4zxz0HGyZe1C7MWYVeYEYEKylexei1Qpz1Hmp/pFgd5zC07
Z5Upygek4pm9sBpP/mzB05gSZrmMB2gMamDTzxJvOzd4kJXWdEm2MixphzU+GiDy
lFq4QRQ/aeEVILq2Y96FggTHQvVGzuWGlbuJKh8M09vRdVoCCh3BEh8EqB86qB87
nGSBxyvL1mp6xumjpfO+x/++bGzWX13UBo97CccT+D3rNUg4Q4uo9HuNX24xB2Na
o7AR3UQ+b9zYq1YG4wEt6Ei8ZrWJvUU7rKpTRYgTLtYCzgc0PNV49DAZp91M6CJY
tYSr18kdv2tocpMY3u0eI0QJ+t+1/+2OQwKQvDNKCmcMx1WqXc7XkCpZBSs4CdJN
MBAHBs4JUPNmEc3ddO3iTwM6920OBmWxW1mdbVB/xeMrRx2Fqwl2G5OkuYVxbqCT
bvZouH3vON5lvtQxsPTpAzXeWZA5QWla8DxHJRiyjpLMwkbdw0YyToiWRCVn/KnY
9NBwLHfL3nr4sQdIV4jU390btLcfEa9L2sWZh1OcSR76Q8kcXPwBSGNKYpH82wso
qlXXel+O5PAcDJX+ikvb/AE9n/aYjnNFqwfW6SLImyyN0dUO9nyynlzY/7LsyPI+
dZ61Ndb6w9AnITZqNdDr8K/gImkbRO76Im+W7tm1rpboToai4LED8bQaeTpgvde6
0Wd2Ih+kg1cf8OUS1kZ6C7200tpZiAkvpgTNHle5Uyu6DV1bOYQ6ihnIfhXQDlI4
tWzU2FpvEEvW8GwVbngDDyBNf/LQ+oM8NFLNDBIHhlrntR2d0XvDnqHCnOk5tzf7
H5TtL8ZPn0NTAJOOPhTflwpGAt3pJRaNivbrVQC8TNORlTERdFsmWN8qi6R591ZF
xfOhydjtOevgy18AcF6a0o2vzYn5YeDO64Kmc8J35lsElCqqb1BUhT1dmAO1Khid
MpkzQ8cVxOJyMiK2GI80w7lCWzr4+aLWyJZhx5X1KXDo5ahsmvkVted0YnlihJEP
74eIYhcSI8ae59YhjicQCFQwc6TAr30Wv0YCvrQU0u+YkJZhVDcIm5UUZu4gNR+0
qLv2XepGL/7bQ94CDgUL5XqJDuyaa7pqG5Js4wRvblCTi5t5ICuuRkD+fzp5oIVE
6rgrokPRWR64qESWLtWtpzYPyrBET1ZAxA8pQT0yH9NpL4pnAc56VpOg8Wvi89OY
1RvzaMJRVgf/KtoeiWvW/pvkdrJDRAmj52iLHvy8M1FNyGoFZ79a5eE0KAJYlZL4
Qg5W/QWZ71lcRDo+fyf4mOmUStHPwq87cdkjxczCwiNcjet4TBDtzS03bw8DxUL9
t3Mv3cJ12fYhpmV2jXXDXL0uXqzBIFNMfrLNOiz2mKXM9qlk9jUyv3KK3s2Y6mU+
XJjNy48L4V/WluPTMxeiL9gtAcN+qNeZaH5S2/cPzkEbQ/Zu1r5GrIYck7Pd2Q/v
CGQvSlGR0EGulUNS7buiYezPqwHzp/pS6//CgIACeROhH8oJ0iukeobmf/3Y2oT+
1NY6J47mihCjxYdhiBUcU87VvxW58NMKYAXMUFvRiunfyzNVeFBeHnMNgUQmWBUu
s3V929LbCaUr4X8HbviLcf0kHh+R2hPZgGkvZxRBWDvmDWhB/eJJB7MWRUXhYI80
xfCHXydv6t02eddgSN4KJnYnlZSsEXbJOFcF5M1Pf8uCk7WkNLE519VPp3EJZxJE
nBTk1XFZViFWncVWSlAjQ2X1UtG7ww7yvLeT2LLUgaU2FPYTv0SjjNoLwXHjHu6c
yQshsuS9G7Mi1JMzfHjgxbqDEYhdyqdmLvQ8n3Mp+IeoGH4yAycFCkVuWa6wxtze
snyPkitzjQlSs10mCD12HC94th45b2c/psQrkooXPAudkSB6XzzfymWsbAeaSsIS
EgQLmDquFR7zdA5b8jNE9KPzygB6r6enlnq4S0BdCK57yp7O31TUmyMRL9eV7FHO
C4WPPdEw7IEPyP5GE5pJrHM8NJeamT7IvKURMtNccLrYpUxlmbHg6/dz5FEg39jL
YtK0DV/psOlJqfcBdhDu+FQHlGEFCklG9UamxQnFfwjcNh+TZt8RFZktpyCWm0Q0
BVM54iRlCxAGmkHmCBjiqwqVSZjJUBOhiOkEZsFUCsCmdahNZR3kdUrs5bnlp6qf
vJUEIj26eXXiHDA7J2raGN7vw82n259iJyVTYDKLN0/vylJ8AIBJvYjL0NgQ+l6l
5YWNX2osvjZEyReaHaHRX2bNfQ7Oy19oQJkJL6Hku6Kbi5nyndGH6s7F6Vx9hYiG
fuDrmCjO+fGr2fv7aOh/oW+DQHYuFfDXpA1FXEPgPQThDoGGG2kgDS374qhlZLzi
YICOmvuND9VWn9DRggCkYt3sc2lu299TW+WNBO9WHwEIcfRIG3HKCMmIUbQHldM2
K97+3I+C/2m6of4+gVVtwjNOXzSgUZq/1k99OuoTxNbLQDCmTWcaqhm1lFt4GUZV
BdswjzEk75JhqkKCDTha7WwzhsFlCFnpBOFnT5j72IRBgPDjf5dRgpDRx+k/gy6g
LhFmcUBc5ZKUAT0qQLPTyJrxCXL/i0C4r6IcVXHnpgmkdBH28r+4nPm100bTH4Fg
Q5ZeSgjCKDvIUXlJWiZs9gzc6EiCxr+AhmaJyesIL7+BtSTYxF1L3aHlME1nX0f7
+XTD2Kq+3mKGpvLVJ3hAEi09pRTKAPL5eUpIN5JTu97VTMvcmX37H/JYDFr8MZWt
KyGZgNzpBQGD/AsjjYS49MvUJcM2sdIr+al+AA9MYz52lvJruuKwlYLgUNFwDEmh
jdUeZPPCXBVweT8dDjBGXrtE9M7hH0fu+Sno9Mir8+kPL5QYJ3ITCulKkXWTPba/
VXU8nW+qvYpZoBz7AQYLGFnN4YdLrJk9jEGCibmpxUQlOiVlbc3RlZzBj3HCjsdP
rTMbH8brPyWsO0X5PsHDhqcWwWeIsFd1PnCIukf6OS8bPMl+D2OEgf+9mFhrVzMU
3mIk/RfAyK11Ft5BZV8Id5SMZXxz1PPoCY/lHeGgOaTtKDSIduyUH7emS3QarMZw
ximUnR2xfb9R4ulMwu/MjaVIqDeudAapyTaCXPvipV3u1uyuvAdEg/QdM+A2u9wR
5YZGYb1jqG8gXz488FzOmrlsN44AqGENWHzlsaM9dckouEeag6oFZnVj9gEQndbV
N2BpXdKdRIz8IEt3z6BjiBwK4cNvhhKptxNvKZA0jZNyMUo81970VTh10e1CCSsL
G04TPaTnITdbxJYbFSnwSQ4Mm+Rlb1F6qysPw80fJe3lCvjDYda8KxZAUV4IQcIa
LdfLDvcFys4BipwVUMrnHXiM5WMTPtTpzcxm+Vz638YRlh3C1EsM38tAFmhjdwSn
IjQqTSQO1TXjFY8wBm+vxUom6+r7pM21ukAATJiQihs+uBB7FNQ2B764rOhxZAod
PE93D7+wjAo6/h7+anj6AKr1SVtsJwRyqbe82scvQdjyBf1WL6+B46mNNi8PMpxC
Vr6puVd8twL7q3MDfK5wlBufhfLjFQuPmvUNaKwH495yKzi9jnB37jADtiBVqmaS
Lo4Rao+vY3JPe6dfqP2P8xBRz4pQN6sBYEnUAobLSfp9ol9j1BWth+E6/AAz+E96
sdT2iz7EbCfQoBNOc60BHwRSjrwOPTZR9A9oauQwbP70KnQ2W0MDSw0Szk8lzp0H
8Z+4cK5hE49x/OCGVm8KVYyfHgqsouytGOvDQHlbLEJYspWQlPp408GtnxgMQ5fz
U9n4YTQ5flefnRNKHU6nBqOzhZXW/hNNhUjRxIH325gu68AbVPXWqx6r2Ys0hYuX
fa6j8H5whhj9kfvTD1/kKeYta62lCzQpNGldLArmYPGOZugTjbvx81gnEDqmvChZ
8yrrH8eSod3degvxiLK6hKZ06EMAb4J4LLKirl0iP1U/mtGKn2MRXTvH8EiNCK6E
6MsKGW/GQQDegvO0yX2YzCEvWZS+WyX9RJgW45MQX4QeDVZgf0/SIcScPNPTdvmO
5Go6HmAonsFEzR5/rRhHh4vQVbrKQ7+Kt//+lZLp2ZJGYlFH1odWct1qmWIPxbq7
BODsXxJO1D3PAfcFCfNS5QDc29iEkJoQ5sgYCAAzGA3j9J2HyGUTgxrKMmEVp9kT
gh2d7W/pboE77Ly0EBJ7GNeWQGETTUSij//zMnc4c4PpLwE4pGx13HBSfe7N6MOZ
tcBHW41zcN6FwMf07ukLBuCWRStJ4PRNuYnsTTuTmm2AznODGSSogQoGdEsa2rPv
hys2cGRyvw4z7ThCQ3KJ+g5qogjyU8u1dBHI+vLnDtopuEl9pCY7xuvqY/j9AnaA
ywvoRXZikkd2+Jpun/XkwvynNl9j3EMATmuoXs+fFhmPzL/5TzcxtXLHqJNInuUo
wnXK1Ns6xF2YkNZbfLmfsGpWXyzVfjwIWFv/+z1LOBd8JFGY1q9nPxFx7gH9lk+N
eTa4/fX6PEM0qZzEP0zGKKCdZzNNwz5mdXJ85WjuoC/ThZCty7Ta+iSYm5iaDHQB
vpAkrN58PvbkTF4amyH5j22x9cEG7p9d8VbfkxxjTLez76aCWcMzW+kp9dDP708r
AwGn7kJk9jPoRYfpxRRpA+3wikWZJciBfTUWNOG7984HvKHL0gH4ilcjIjBSh3DO
J6VH+Jpdo8wrUr2TE2YJv428j9C4W8XCq7CD8EiOYr9ykEK/gApyh0++dh4YeVQC
DnIDt4K+tzRQEyZ9po6iBAfcOrJa2aod/FJEUZY/T52NDITzNEK4gQ3aK4LlgqXO
p/afjtOzuPSBgt5G7HH0ND25H2SjnzMC7y+PQPPebLb11JDHIt4qnAynIQKEiJzS
CNhZ7tz0g6rRD+mAGLBJqhqQ26bqpUlFCKwof+nTMPNOA5B2t2YjM57kBKm2IPS4
NdEvKMvNjH2dD5k9INFhuE+XWQ7Gf5HAkx72J4ddo04MBZ9lDJE8ZB9lLYSp7Pp0
+2zVMsvT25lotGVfQp/N8FwoZQkn7oCSqqJYg6XI/4dKwkRyALEpImXsuQLUjl/Z
/i9ePfPD2u/ezqRINwwT9S7IiQKMxqLogESMXgQA4PaAsxs+byr5hYLNoiWaCcIy
+YdaQPH2mtxuauTukJROZJ1j4Z5vLeet11SVgxtSICKfEFajUGvfk4lEyIiBVS1N
Z901pbWpJSVA/6iC6A5RA3Xr6wB3Qho7CW1gvfbelt9sWT+NpzuvvEDF/9PoxNcu
cLGhs0QSrzan7jBG4Vv0280pfGILgWTXp/sewOIU+VWMAOwXsRsHG4XacyKKZ9gA
vHjSYVnfYWDcRCtNxUIR1SzpE2qnnREK7Ibv6wtjwHN2cZMKXC4oknJ2GffssW5v
rai/4R0/z65uTby6iag417rVnHaWsOsIPsCq0MKk4SyledA5Q1T9TWbssPvW/xFG
jZLA1cYkrCDATMuCai7Z5ijFrTnvbiOMTHyI3uDrK98XiRuErVfitaRvhklhcrtk
tuzWzBp0PGJ4IMJ1g4/+EAUYPFE0S4i+yCzKA0ITbnPSAZ8W9XOKWfNGaIHSVxvI
GsSV+5i0+ad6RY1bJXYz67L1XFyJP8z8iXU1DQd2HUOWFfRz48JalCDf4lT8Br3o
pansFV97Ih8O6wGHBwTRgzoNyCBdvL6Hiql93BUTFcBqalJl1Fo8AUqVoLElm19K
T9Mpb2LsO9i2qdL/q4XraB/HgNWl25YGVIEWBMoxVss2TMDbxx0cQQsYqTqmu82v
V6Xr8gA/1hCvvPbi3J8parWz2LFu5jKPAUHAIZdbzo+JfI3aJlaXDCPkEe5oLisC
NmbhuCx3FjALeFQnIs0ECo+5gqbRYzS2Xr33vKbh0lJugiYkxRCWD5RmN0B51LG8
KBlR+03mBtP69zE2VfQvbltPDFvP3KFIR7fu1unK5dKJOukP6BHmOmN3XjHs7z+6
hJyMGj13iukkym136ZQ4znQgc7GOGzUHMXuzSYqjCWgqQwYyu8qdGtEIzO2Kuh1+
cXVrgn8YRY7QHAipKDMB/ls1BFiTeqI5ATQMKZ1fmdHjvQg1gIPJIvNViPqtyEHI
iKF7LfkcQ/PzieZD5UuQhRsSensYRuOUbjdiY63Hzc/YWWYFEGvJNICtdi4TXpPy
QEDI7wHYAU8RoxaQPtKTeUfunJHEa+OBYFueEHVtzd2dwJrp2831dEIhiKU/e8i6
xnCb6DM9ikk/APR3Vn96AoaNiVpkl1H2HuFivlJ00/s9iXdwSBNlNgEVz7mLBAsa
pgBVgr/85o5c+FTDCrWuZ3WVdGe/w054X/9cJfnDTN5bSVinFM11TKeLVTmYOb03
RTRnCrO/F4SgeMMgFKzs5A+GsrWWpT883AUsN9OskObDrAoVoUZOCTUJIA8iH5xQ
pj29xJ+OZEtHJBcY+h6IgI+Ny/zkSSH0tTBEZSYiR7+T+fcGR216s5qxqX3bN41Q
VngxwuN82v4gm8eCPIHAgG4KyhIu97c3xDet2JxZw6ReG1taEmjwHk5OAkOLNZCg
0B+s7N0ZyZVdYJCfVBFYOay5wvohQ1xWlRdEOxhNs2mAJs+5tTjytALKIQ9K/Vq7
jClklzf35CevCymsZdZw8tpVD/Numhq/rK+nlH3FEA9y7IUzQlkY6sJAiAeM6s4o
8Lws5gS7D9cki/ov7Ok66/hALOxPtmSX26b3r5GUOjAbBJssUBHRcOGTgFDEYEIk
aoMxSg2V9CzcMbMz+dWJq9Q2YQbtdWjKqCRii+pq7WyN1Btw5TntVQzVX0OrThBi
dkYoQuR1aced88RPfK8XUYGl6twBx6D8HrbliPdZKgwZ6swhFV8+dYtSp/++irBo
q8RtSnVKbSWLlv++VKBpkZ2RAUP8Gcx+wCATfU6tkyUix5U+AmkWDp+8sIDjc8Ie
XoRhOr5JTRpr4FOYY8BuP+vzQmDazRxW9MDLDIe9bZPRHN/9qbxGG7x76JpanuFP
l6350teI88nbTlSOMZrCUoi5s4GCxePnWmOtmrWpA2b54y6QXBambjcijjLB1uBk
mw/Rabmhga3lPySAkaFZ+E5JYRqsuNebwTBPyDqji2CnYmgvya3qSg7i2UdU0Mga
bly3XSLRbYc/n49Pfa+7fNElnX+dXU47BD6jmSbKsWJE6HYmW+r+/q735R66fgRO
R/3RY4E0VeElbwyvg2z2RrBrgSCnZd/A0MnOhTZ0HrWH1eAdqaxepHgAsZINcDVA
o3Ri7ahFAu2U8TOyaBJ5LfXqFrpxrsHyid7GMygDqIOvOz79AWSWWaWK/HXdi5gU
aIeernDGetnXREWzOqeGg7Cf8GfLWgY57opnCkTVAL1IkbayUHIzMzQfojTXC/3k
vDCP2bhN5605oGe5w+7fzr8DMKZnEdCFtjzraHFRvY/fOzkR346k63yv3Y4sMYRA
VMElMvxyrddZJF1KxObxlyRNdp6t30u4+wvtYS7olpUD+sSUUCCMBV6gxITo+myv
3aTRZe+LH4NpJhCrLoCN9o+1xwbstb1uRe18DjPkLinGHpw4vQMx5NW9zKI0NYGD
dCCWe46xaCngeW/IygTdRizcmaIouOqZ2WQNTJW/Blij9GZvBujZD2WmULMD+LQ0
vVvuwsYFOQEI8zisGAz0L61oBvOygcqG9y1ne29bm6cjzXDUbF8Q3u3arpie5U74
MLNmDJ8MJqNQHzqm3PgYtdbB3u7PcanzIU1XF55IFlKJH/xr1R48w+XZx3fF877c
0Djn3phKpPWHLIgLRWnn67SxBeP2Nlw+8L/tvVjSuH/Z8v7nDO2OWhlUEVmcHke+
UJwSPPirhjErkUUIm9kSJxwfoy3c85oX+xR3bVL+jCG/bJpFLLmpTqK6yHB0lyLy
Rg/53j2AHTzDXqPZi3gVD60MabtgHZSxAsOeoBuXpnZO+GGnUJOMIKqmSwIIhFgd
A6uQqu0rCuAP/edK1tLKxL7sL+RTq4lEZdmD3s0mOGTrLCmuD8MdHC5T/D+UbBeD
6mN8u2R671wWreZdQINLELuXhePWmVHRuDGyyC9i40Ioirh+86A2TYJrxguZCooo
HXjlXWhS7OJ0WGrCqsVu38KrEtOsEbSJXqh8Q7DJS/uFAeoZrR32Ygz+xSLuneQW
ok5wdVcCfcl2gPC3O1MMrKxST4EhYKb5vHpBhwklwyrHFRPigxFXCHaM8+yHGjlc
6I4I0paiFgT2MVd9LS08WpMSJ63SDGotzPe4lHG9E4I7A0t4b2c1MTpYo6HPJQJi
vf+RcufGL/AJbX/TwxrZlic9s+k5RIfUpw1OzN7686ChnFnPveogbJhOJGQVkS/m
+olacCjxmv7V95X7CaHZmS02MnGmG4SdZTcaZHNFfI8YZCNU3HulDdRtQX0Gg6Xn
Gbr1l90FR6a6NDkwuaCiCWrbwEwFvnPwF03ohC+xu+kvp7Y4cXMeiPL5mBrBzh/J
3eT5f1Zi4qDBze/qn9Eu4o2Pcz3GDWuL1hyPo+46WWU9l3/3CAkaRrwSzfQMOzDM
U1vwF9rCnwyrX3qB5GU/5t7MNWRC6Fzr+RvKETe7bKxWekT0dSl0umFJRlSc+FOE
xnoQD/pUZtgl44OKHO4NoydMVO+BqQ6PxQ5Mdxgbd9aE4O3fqRrMVRuKtZgrfG7b
nGXQUrz8M3rMUGml3WMNp6xR37J+JXO3zPhxlVG1+y/UN9FT4TVlq9SkQEJMBkgL
3FeKAI9TY2A65cwTBL2xUX3LEVlm36C1Db8uTfStcPJLpngsCX8/r+WHKV+eVjtc
l6Eix0JLQORAvbXb3G5fKiVPHcuGY5Y+2pBxuKWlloZi5sQaergUdhTAqzsvKgiF
JSvbXOq8v/BdBAzNOI7nj4vhRTUt1YZDh5S0nOKQXwSpl7tGYrCt4027pQxmoQHl
VEJqoKjKRKFZ6+NcTn4lhmqgcN8fm5M9AoBIa6KdrtYrg78MqxFnKZ7P0jML/HTG
4JEao+wY9WRv/zAQvIKjcx/ewGbtVDtiXTYpl2OvTn5pTnsoxu+CSj4i9SFr8mGT
oR3jjxrv5cBSSdI8irLHi0oyuA+yvVrXIh9U2RhNNnqwHbfglSudAEC84WXrJxGi
QHXFV0w8DLQvtn76S4YUIi2uGDrHbDctZ04HmWmosTAD/z9FFMlQUDcRSq/R4T4W
CfoWrwHxgRMMA6GhppNmL/S5dS6snCqXtozlf5rEZ9WPa2lbOMQbYHF3c5fkkywT
TxNkVyAPuJPSB96kFpL6AkMRgJpjzGKnhloAUVcpGmu/EurEpo+Kl0CpzqsxVCM9
qi1JRJuzwBBgNHsjurX3tOpYNYk+4y2mr1c2QHIeh9fZyCytaXuCZsgiLH9raPGM
UIKncEEF1471KoDDkjvAyEU2afCmShg2xcq+7Nn2mbKXbA1vnPWFgBnc8LI+r3su
qVPDpdcsRIZnbhUHCDh8vtMwemBe7fQUgXspxU4Pl1MAZu3SEuXfoVsfjAAHnqVS
nId+1iuvMknUtySz4/8ficBuL5P/+B5SzBWr4PNZLcKjsaPmZ/9K1QiLVRLS4enA
Q5QdaRMBcywBnImm9xfdFqtLi9mHUMWlmV7OQUjOLXRqoWidgYFAxi0oFIGmIqQ6
HOetMDlx/SW8w39xiF6MAzf++GoCdOTvb+ogxpeLc4oRTaRAo3shheKnay6B717v
uzDuIvUFNk3FM9knd58FgJYkFKzU1js1TsJTptc/UyFRujz4i4wzAGOEaz5uIPtF
KCTzUFdrTTaMWQkNweo/wAP7eX+/ko/3sYgEB7rl1kEmpDslkn7h9TU9dV0JATRN
IQbGNrUCF2mEmhnEvxsDJlko1NZ2hi5jN758iTFL3adkKwfSl7ARY8RaL7ZvUJVW
/jCWV9jFF9DoP+Mtiu/SxnZz86zwVKCLuiFzeceDim0R2EQZhwqZ+9FIXL4UyjHA
jQIgUO7feAe+aNFWi4MM0xj2Isn6IBqBRFRMlcqS9AhtXTRhWOXnxyf8mw5ofmlR
3bW6HiaxOep8XSCH2/TFOiu79pD6BBWL90NJbdVQlX7RvbvoCYg1D38WC8c2OKQK
74F5KUXBi19zLjZTDfZTH9X3cLj3gD5llRqQCXgrAhcL5M3VB1UQy7+RYnizo9IL
siIminL+y5MbD0u8NV6ztbKHE7mSz0lIEo5uVGg+nme7dLwlgOPKbMIZFYNA1mW4
10bXi63O7GIb8dRppKEz8hNqgMuYr0iKLKuz8eFkNWsfMRppFlo2vEMeKFhhLPgm
2AbLuVY8maEUQdkH0/URya2Xr+1Nv6C1GIKrnryQ4wHMpN3MnNipcoTH0dXwDtfr
8XBvMuWQfxsna+9Bo6svGCdzW7AUUVFiIldNIwskLcZVHdHmbaGA2KkbIQVA+AjP
QSjlIK9wid6nzhUa0QltYengO+durOaf7GGEZ5a0EZCO4/YDw6fD0XFUdiQ7Mpd/
pny5SDHv1DcE32NvEGSJW5yk436jfp8Qsd1HWQlkuDT0OYAixlGiPuNA13SBI/mL
n5z63LAunb5qy7arSGJRKOgYGQAz9+Hcl3UeHMLdrUsevDvg4IjndzNZf7nZjgCT
8SA/1LM0/9tX2y6nZYtrx99zfsK9gnyS1HWcE40ZU0rUUdWBcCPwUvZ8JUd1bn5J
UgK1uUnbKaJ2oKI0LG3Lf7d03uultBUQn5AJF/V/n52m0he52WgFw3n6eRECcn67
DVyyc8ZPzgIW4+4ew105U42LtsSols1Kg+5i0RRUtyBNOX1tYPFmAiZj02HAfBX0
J95W3idPXrX+d0Bglq7KFFC2CMP7TqhyiRykLGNQKYhGksLNRpgD0QKzN5jvufDe
yreb39Ad/v96JbIeFpAmxvmmIh9RjyMcLruXoyxDUkZ6AcGNo1SP9/2Xk0ffdvu7
+g9zP4KwArA/E/3TIajJG4uB4h54vcidoPJo0miCwnQU+UkK5BpMugneRBZC9pEF
lNLdtcNkYMJaXPILMm07YGWBp/6+ZGbBO/1r7zaEOT/H3JSenRgqhlV5aD41tarC
YCyiCcGjMTLf/smAkagBsacbvCmScD0eiII5rguGwtKJr5c7doUrhPKu8yeWTeLl
ZfgCaqjzLhsflbupo100gNZZWktk9OKKNQkV1s4AfdlZ3fGpz84cxo1xs5HNaTsl
xdQjEE+Jo5zm8tmTfvOrysn0qtoA7D+9XqTdxL+lZoc54fsezlhzPZqsDSSuNHN5
PoQRq7GF+cj8m+51smkDfhVZyS2QTVa/MqIdg2Fx9MdIsOJZ7NwFho4L5q37Tkd/
pJ6Jt0jinOaKWdt9dp/wMSv/IjkhDt6M9i3cgA9oeRpFkcymGm9RXObtolIlMwQW
qE+Cc0Nyk9v+Z8SJAcSxfi9RStrKGwC/C0OrGWGzu07Dl7PeZhSP58W96yNahq9V
G5uBcnMdeZG05F0DGogWaguMjG5hA2KN9piJxiSZ8mVr7PKzN8Rxy+3uamz8dCGY
v+ruefWv11VyhwZB+C6IJwiEfsOnuamu1zYYyQ+ZZmZ5aErrj8m6YDlJowmFGFc3
K5pbUB+Y5Kz2y6FS+ab4aojH3RsBOg/8JgVCnowINj36LisRgXdfcX+1GB01vY/Z
UDfBN8FcD5NBgwdbLZV7mt3eh0P8vLXpOsiXUB3k36N8MQ0DSphOtUF+IX4j8HNS
hqV86osCBAym2rCijiGPAB/Kx6Ga9ZjjSrrpwbnUD/5hHs5jT/uMlEiZs+1a0xeg
96/2K8DVicSh4KKh3bHSiIdzSdYCuWCC9Bd7112DGi7+AWLh4hndGkQkTCV4/s+S
21/u8z1VgHmzRTCH96+2FbEuIbI4hwJEYfd38AHFSGNHj2NwsAjneGoxDzVblw/2
+/sFWjsi6SRAQ8ejFom92KIAQB3XZhPT3yHsb/aJ4bQxHKntatdi9BHl+iijf2xF
IBoLftONbvY0XWEhDOqjfoGskmrDerC0noiqA9JW6laicYxHatXP8TMbqmJVvIll
xhVzQ4K68GHg3rH0fi0sY43j3JIWjouW6zCDDVXJrH+AE5WNUyMXvtOxs5ltoiiK
skwuHsFJDd2tUsm/ajat1RRGU19RGAlo8lN/q+7LOizYc4gWomY2ph19NqSOHros
zd/Pqj/7RxDgKpKlMAovUWgOx1bFkgtRfArWqkkA8+Vw0g5nR9NI2nq+kim99V8v
CvRkVgvLAa2nHfeAuZVp5FQFkQ3oAiLlMVZKB/qA11y6zqFCu7dpodUkKIoQO9Iq
1Sjp388W3XJg8Nn9UlovJZYjfZFyjghiZuF6oyStYMQ92HApF5g+foysGhKQMLAL
MDXIEZXrca8nQunx+Xr0hVkfflDtNNSeEbLoiyssEnfqRW6vMVsVW16pp8P++wve
vqO06i7H6+iLxadWKk9DApt7CI9V4ODWAK6clR3eNAQkq8edJoT4I9EP84mR9NFn
dCP3B7Q8U0o1/CtYsW8qWMxDIkCsDBNk6tXE1eSVoGj3+acI6mqYyGbohOT+cDdM
iJpsokxLPFuGExNPZeC1kFYj0YfCvPQ2uBKrDA6sm68xMdBLcGYSoV872z1nNyv7
ONTwsxZm9bMMWcuyDVnpAn8qerI5pXKULp5vAlVUWRPATlal98004O7cXBlxm2dt
SYoABn9KyAh6IvsuLgc+VANNv5Yz3wGG1SK0wz2YSD8nldNAqTwgfupODfOud6Vc
B3INAoeV99AAvwbNzTsMUhu5OwvjG1a8LEF0IinfW0LGcXeXdgf7WC3jxKzJ7XuS
eTqev1tUz9THk47n//KTi6N0qJyatI+HWoD4HEVvHpaU1Y5YcVEMcSM/WmnvvRaW
DhEKjLmhZ09izGVNQyJOkHVGvo/S/Z2DmevyZo+aWT5BNQoQP2+rKrtXn8ks9W5Q
Hb7RYc5jKVPWMnaau5JOmYntP8ST++zxwVwN9nq0Wgal1hYARi3yQS0wDQxw2MTw
d8wRNlG6XW/57+fx2h5rosYIbjyNDttOEWlsuP4Ft0KtvuzTGIt8/Fw5f6OqExsN
7yix85+TsoaUpykwWPxeQJwVlLMDHnE9FzR5HCN/xoPRTM5cJP9RHNNpRAHs/zT1
Tmx1i4okfV0J0HFP3dSSKzDqeUnOnVkG0apx/uh9Kmd1xJNKGnEN2XgJhZsQ8A/k
ZlYd0wZ5JS3zC7U6mr6rDHB0GZIV7bwd+qrPZB+vS2qfR5C9wCXypaN+8ALSxXES
nI5YSmSLr73uHLWJ9Sf9dl1xvYB1SmtzY5TpiIpakUAqxgU0+W3CawQlE16lQa4e
6hUrC+3FIh+70UFpK1nKyF3RPbQ6aZ+xuctRi+s2ko+8+XARjVfxjT/syM5zFU31
/WzgBmnSni9BNZ4hrUnHaiQVCcar8Ia0dNpfYbL1Lunv3oMWkEyiU59PZan3IlBd
QHM8CF4m/6lJzsE4cEEx37VZuV8ev8nukMHoR8QDQuQ0Ofnv7SSc5090HuA+Kzi2
nVPfQLdPk0aKoFu59IXjYKeAIzwc+KubnDgne06mRgggUmOz73d0KxjC7zHLxOC7
oWs01nQU3ambiWLDa4XbHcssrzWuXYX53ruUVEEC5QMuRfZcftt2GKUp/0TATRIV
MNxgOu+FLrWUHXujCultEXce/kSLKpsEtKxJmm7SK4fabVy3jf+ZPC2bTN257LCz
mb0XDMD3jyZpoD0MgllC1qkfgHNKmSrz9CuXM++VobiLx7a12tOt+rtcej3tGbx4
qKsa1Iwt74reEXrv21tTA6Cy2PeNSL60ueewJ5SFTJGxwDNZ+/RIGrN5yn/6bMRt
G7Mzn7vx4iOoeJ6VOR1qP/93jkicdRnX8N8MqcYO6WTbRyKI9n2dp6IQAZ4KK+ku
Wtl7d1Lj01rQJMwiHI7lK9pa71UnDhif7PX14zn2CK7zGbNdWrAV/h4g7NXXlBZc
4GEt8/zNcAoETeU7jX9PaCpIXwMw4Z1yvHGfCbx6846yVy2O4m43vG51/BJTHylk
Xbz1pzYk8wgcPtrYhkXqsql+4eS7JzS/XGmp+IAmIBwSCDEICkBfOV8DChV5iKwM
6q4Kf/1J0HX3TcXnJUMrVPWAJKMTr//koPpmqaV4g2l/3A4EelciXFcpMCKphPIc
Nll1mP8slHXblEO91t6RVld9VCztbljQlgPSGu8vCmb5B8lKmE2WSKdWt9L3qoFR
SozAYyfrQBFqwyKhQRfmstj6FcE7StpEogKJhnod6Quz52enFZFVwicJUvH7x4x8
y4YQU5xkynoTEGNBcxWmi0Vs0yv5XDMg+dlWpPz28jTBDL5+lAcRlRcU4EoiF/JJ
3ZLJ6qKPOQfYrswwl3U0DceUqzdN/930EayjmgNELgHbc3N97mS+0fLjZBMUYQsA
t6WlJcanHVS/+vTBOqO1CylYFoCAyy7bCSHwebUly16GndO+tHN4/4Xq2lSjJhCH
Vjxq3ZpXTmyoN6/zjvUO8hIl06FDyAfP206YqKdQUPPdW2XrR/+L02YzV9Ax2BDd
EoVloAzErQZZD3WJBCEkGxkW4ek57U15rVgEC88eqpe29b1WzShoetrlZb2thNNo
bHH0sKseTacIcTs/E6JoTaqJRsqz+v8TNdhvu8HpTCwcp4wqH+nSvboKekpU9ePL
zxlKncaQN5O6TJl/63rX/gBc6wwTb/ofOhxqxKD3RD+27kBGM45HubUeL+qxUoZI
J9rkGfnzgUZeadp2jptjx/JOistaY1St2W4CtU5kE4P11NJLt5g/atD2k84QQPdr
r4PDqzr3YhDf08g7Y01NFw2jR40cA2Nuos+hQ/bxiZKLCRnufqmUGId4FfAtbm0K
wwcV5EZHZS5GiEcpPlvxIWmfpZb8tZNBPw7OKdDcZ4Hsc3l/iaIq0XI6T+5AZ0lW
OR+4hBVb1ONtz78fntTb3ZGFcyI24iUgdqNKbuSmNwq8vIvHiZY0GCgHe3jdduRS
zlv08pJY/ZnexYipS1VVsd5bsO40Xsb69tTBY3+BB+lLbZQeK42NYueBTZpex/BB
h4nGNahGJp6f3P19hEC0b26Dx6JviuAafmYDJiRSyAJuUaVNDlnFXQO3NciemrPR
BtiQ245u5JfQjtnRO6a9nPXSbq59KH8yGq8B/y59SRcAowSYk/GEfihZm9a9w1m4
MxeXf12gj+hqqvl0MHv+CCzBrTJw2wlwFydMgfz8HNOiFLNXINEJQjQdS4lz650s
dAGTTozNMw8aFpDbXN1SbZMhh0jCbzdoM33lmQeWzaf1+uL/vzDcSJeut3ZFZ5kh
0qNBzB6t2v92w8I8tVx+qsOvZ3pmYZ4sp5drtdE6gKMbL2THgvEb5B666SY8H1rn
ya/jtTzv4+2IuGVLbn7cMtrco3nXl01XqBTFPkPmM4DQ2onlOlO8/TZH6Ph7mktW
TTELJzhRaZdDcKRtWPUsCAoWicKtlYAhSnukgTSkO9T8KJUS9PfCdrLSqqNOIYna
9BTLf1u4IqWgIpX8+IMxWGDNfhYg59hGTaSkw22DTgebSW2TJkNihBWy6dXvNF/b
a/7d1lllMAWuBKUlrSF3UYVLihjnnhemzGz0fCEXuh/aTxuntQfqawDAVRwUjbsX
GIOPBKD4ncJxp+v8uFSY5q9s9zGLRI5BUnOtjfX7nL8K+Yj/PqfgZE+2Xcj0iouO
wYIDT8IqdPsDKFc2QpNxKN1ctUm2NRXCEDHvE6z623wU6jcGWr5BlYysZRLp+NYC
zgdzUPRr1jmy9r164f4y8+9M4gnACobjbZz5E6WXKEPQxHoa1zxDHa3Yb1I013Td
V6nNu9j0ywZwv9yiDabJH8Ex8K6xBtZKBr/nugfAn4XustMfrqHAUMtZQPfz/Gx+
MoAHglDlkWr67MHZzlfEuUMfXYDqZdWdrxdJxTberuz3uK7FdXveZNeq+5h6SK0J
mjF8nDgMIc0wq9CgKkdvu8r+xwRUfuytNTv0WkDfO9f9wsYKMcl8q7RPk/ipnK9a
XrlQ3aNjO03Q0uB/xKdUjWwIxxiT53V8u6VYWR9PSf7c4f/CuSfXxkNh34h4OyfM
ykjj+Vq2+lrRZplEb0FlTBrSr2jdNOw4QHsKp+y6Lai8ZjGvGwlqogLCAi2tlRF9
a0EwuDyquK7AFqw3UU0dCxkGIs4rn5wBUaGfxLMFrX+0lt35Ktm7i8l/wdxOQGIt
JHo2qMOWpZAp0nRqCOWKlcBtMiFWTIKKqOfZBjeid+NDVhXwV59bgDmMXMrIticI
5srCkSkwPll+Dw3ukBuyuonnf2HRtB92LlDw0+FH0Z+7ntNway6TZ9nBNKE0gXfy
xJpbN/Q/Jl6Uyg/y685TtI0YVl18d1Kf46FxxQ/+Qc6+ppE5OwuFgFqv40hWCEES
JpogZCMEN5RUVQWSapz8zAf3sAueupdQslGodD+vvOsdvKJKb2C3grL+Ncxdah1k
9+U4oXlRCogkDDR2Cjmez/N8DU+cinSco/yUCFOpo+uuE5CVlcXsWnnFW6dmi/B+
+EfmbTSPtzhPNSuyyPXiYLT4H0xZAstNJC2FCVO6Krb1C4brZmxEUCQG90MBn99M
TrnroQM7gE6aYUqf0gOwu1qmhQGlWJ8GRPHeIj6Gg57SVq2QHSnFMcmrzI6HmbH0
9Pt+YBbF39wOoDgwBElwQ69Tzf4Z0L4L71Qy/TBck1qvjUBwpR+KhnJa73wOVDnU
+wwD0irA6ApFqhwbrxdEqgBPqmJCl0MpsEZEsKheunRwfDNEXd7y3rVCOeR8Zgga
LLcFssjI9JaASNQXbByy+z4rO0je5JJJnKJAleYiLVOPFo4Bi32vE0ev6kefgBiR
gWGEy3kr7T7x/N0rFyg+Xvt0rm5/jQvoqoUM2hQK6POhHThxLb27gLkeoz6avHT0
OI5adgjHVOYnTxw2iJM3Vnvo59dJPznHVs2kSN+hFj19pvIWeW4Ms5hqS0UKTcO8
SAc12aUw1jazzUAe+bZ4akzBE8ySat5MNu9FxsfB9gtIBw1UpmcdaARhYr1L/JCJ
w75bF6GmFtWHNIEjsCU2nR98Zlm17EJZZgwhu/z4VRqI/zZo1nhQNSNc2nLA4wZf
EvpwJrEY4wq27yql05oG+7qesnKq5pNOTYkg9oDFWRpuu41rVrSRMFGMT0VWV1iu
UFn2BKmdLO/mlUpRC01rocKW75EyeAI1EUQL0v+sRGzYU1cXXKhEONxNRFQ/ulVy
g/T/rXgUP5qKqRN5zrVjj3lkHxfYyqU2JSC997vgbV+FEKsaIZpTujPXiNlktsx3
oOb788WfzoEWeJI7OCdVUuBTtWbzdHqjgneRPgibMJbg0c7szymnObNWoVwE4y1T
0nqPB3IKURLWRrKTTXwuWcuW6jlbBGwTQeBW7XEqzV1sySriUcU71mY8Mf8ORXXm
bkdK9vU6+f16Io44js37JOtYPK2tYzQF29cqKMXL0kEWp2PPykNkjA2rlUwWccEF
lITtmwN5X68OzKAwnlFfPMwXdnki2eILX2y4hCRp8DOzRV4QuRRDfaQ8yIMDe5Nh
U6zHTYnZN8wlUJEDmBPo8xxp5m+f6qsxluFngXYJO0fZNBa5rYYKs6UdreZJwKF6
CCp4rlV54yP+b7bTwzOuak0X8nT2PQwSmdwAQB8S9n9SXHmekW47PGxEFWNZhb9L
DFZmjzj/1zwtRqjt4/7pyFsW35A2iAlUZ/PbifCwa5Y76JdYgBrMPMvzowCDgYyk
rXtOYhclOOLH/a8DcNxo99NdBlXS9ne5S4aKIYR425BkqW0LO3Sa0FZ9vMMOgqzu
OdyyNKe4IyrWwBO3SxuB4IA2WHDVa3elZKd39JcG4R10P4STiYmj/JzdUwg6HhdU
7WjyrwynPGAlceMu2v0bMK3HpTbOkQNVnibRb7OIG93Jy+r4UjJLa58/sLREjptu
y1usTQfeYxEAxrDfTBcnSrZXZ8h34vybpERGh8w0X8pc1Y3lEg/1OAa4Qsv4ebsx
4P8XSR/m8zWRvKmwBtgMbOie6wqriEI79yqHOLc+W/lqG94RFNCD2W2fIRtP/8l/
/UbYzeAObQgf2q4+MmAMsnD2c3OfmlMRkHu2jtUUK4AHuUMUw1ttxzyRSvcawF9w
qOI3SXGQf86P0KAR0NBz+Sijd55CQ4CwguCQfPz2rl3xIDldr3UOwdfZhQqmAgSD
cRj3Z0MhOXfuJFKZrefuh9bQbjpvbKTWBV8Gm6Yv192rAfvPx8Unp9X4tDafyABb
R8qURXeqmOBsOgM8waZfYabAskaEp/5ayJbGho8WiZllgClprfSkKKzQhGrj9s2Y
7u0B+EZ0c4tB4ZjLMsX01QyZUfhqHerv3jHvYQvzncrzRuLkU/rhLf5/RbLwE561
FI5u2V3gqrrosjJ7DSzENmHdBU50EiaJXlfF7t6xFDX73CwYrAjP36r+aOaBHQmf
RV1bYAaG24SzoUAncuWsxoDPnQa8M6v4zZ9PXpw0HKTJbH/Bz5re24dbfXu9+gYp
pVzr7rCqVeh/LpmpABV5CNAGqbrOiHfsETnep041mvwZYV849hOTBjN2m+2wRxR3
1vN3+mIXwjXGvscS/vdSVg0ntELi+bdhqDSjRAKsIqsBlWZdrCcr7RinG1Gp/W+0
nvKC6nkTbiEUJpyvOtC4E+V9guXDyzsV4Qd2yFtO7eOuQDuSIM/8JEyx+KkbXUO0
76E/wgo4kXbIFDx8eIqbToaEpuw7uoo3Zc1F+Q2+uyGQ6ctaxGKENeGuPmxl7o/k
Cqy0K3yJ5TcwrPnDc8WfQo6xQT7jg9DrjQ3k2OCT7f+lIPJe/7eqm+m9XMVFK3Qv
YZrtr+Evw8zMZ5itI7CT4Pjb48fiGPaHRrRMQcmbhR8AQ6c6K7zwSany+wmwpqKq
R+/FFbfi/ZC0NJhEvhw37ibjvqtueRML9Fz2s5TTJLUlR6ahF/3833qbut3bJ0YM
v5nYeDbXcHtfsusftYtlPNmJdUIzxJ2HyNakrYQjfjKg9ufbyp9njVsewi1pJr7y
xJjb7WQBXOrIsGLuQTpH3OwTXjaiyjCtJs5ITw4TRaFW/kxW3m2vUB950Vr1uegG
Q+BGy9jfiewwPNeSydBT6iJWc1YY15hY6l31r2JWtVDKKudKP+V3m9Rv6WmEpiwC
z6awIyYOU29mDFnmgxdDUc9nJ/PQRHuy70YMaFUZIYR+Z3Mrd4VCtwLrzsAnlFZC
dXEBh6ICpuuvRn+rSc2xaCRXUiV5zNrKHg5XAfi0j69NEv1ugP+Wswep5LUWYBbi
g3aa/SWTvpqj9z4GwBk7LK3aZfBmuB4UE45ZvlMTOueQjP01PzqU96uaI5WIs5GK
09J8riFZNd2zrkRtvq7KYhdmCrvnQXX4AnFTwdGHF6+V//7PNGjLA3WMa+Si8xt9
oPybcmi0lrhBp+VCudS0hQ6V2QBHLm4YGC0XWmqIhNSPt48W7trgX6e1mqUgsxIU
LwZQfSizqIhGPsdvH4RYAXPirVBe9T3sbbkxCC9FhobFTdeQp8YaHj2fU9++GjKt
m8T2ASjRumABrOWIoSMinGk9vmbdBysAAgWP5SZR+cPzksEaSkHf5TeX73fDi9Il
LAXGupnfAsIaHOVzQAGXqqu0cAcB5ljw0RPAkQObJOzD0zN88yDZLe011GL1DaOC
WvE5sVNefx1gOQxmbeHRZJT2z9ITwhBCMGN5L5RgiMtlyJB034t0PSBdvhZC5LsW
r2m/PV5YVXQ7ozaH1WOclOhdiXFhOpY7Hw+Sg9rCDRxuQKunkfUeEfM9vGY0wGgz
gvFcYnYEclSg1yOEQVUMGFRoan3UF2Yu9kAG5A2zS0KXwhc5YnjiMsKAfMkT00M9
I+DM5X9EwDqz0hJjGlXXLZFuw4DMl5oZuvrdUVkKf4D2kNnORmg2l7WMjikC0MA8
mMK4UfYX8ed7sIiHPb82su7ZiNfV5wApqU7GGU6JLwOPgKqSOqCFnlry2rGmEJAN
BiGxHu6jgSnZmZ8FXz0Lucx3BNXjYDFfZkJdlPZ2YnV3SEIvAG8BLUZrZFv+c/W6
aUtnvzrRC6YA8ouhkmtyLQio1C+Cl9iV5wqZzDeAwHmdpjFbwn9TBubau577rHT0
eNvfd9ajU387uvHZzekH1rTurGm3OKJQALrwoZiuGhkyb8Fl48Wr7DdfnLoTHSfc
1Bgcrnyx9mPbJNMftLAGzWKw6nhjpCKc0V9hUF0F2iDkmLtxsv/8rC/Ycf4DSHfO
/NPLv3JbOkqmS72gySfFg2+jmdpYXXsK7mb203GvuPSUBv5d9vQRIP5gGv9rWli/
K1vmxKiVvOpnNVtFPw4ek9rw9rEDznTKfmB91U2z/TfiaOWAJKMqTeMbN8GlARW3
SAdlevwx+H69mu74M6++YqpiAN2mmYfVYkr25tpSwZZvxikxjyOYEhdA9Zio+Psv
RLYNioNqkg8V0Ing20TTKS5H/WJDukDZjIuDZ4cnmQ/jf8FE/YGe5xaNvw/EO3tr
rPR0EzhvHDFTDUhZbcOOeum0C7HIiEOy9xeR/eFz4b0wG2TbG93nCNaGVPvEwaeG
zfatYKV6eh/2s2n7XtmztdcVWN4lPlrYHUkjmapCmVQvwucJ1BTfcCe39Jt2Csa2
05MzTTeDMYicjKXRNjnuiTGR512O9cQHjF/wn51hJSOXnTgPpoKvN3wEbvlFyHHt
Je4ZN/WhUAmKtxaZPkhOwQok2aFgFuZfV+iz+FTXxODYy8VAksc6A6M/pmQYz3Cf
f7BJUsxJI+rLTMpB64M4+whRbiErGu+luJzPcA13jPkBXBSYk3M2zOZT58XkcgmX
Pj9Zig6n78KkGnthNu4KDQN3qZiqMUK0EQz0rj51Twouso1RJXcpJe99GAiGUzHS
lM0y5XB9BBamPPAU614H0Bbm8YkA0KimZmTMEX9/5BvSdVlsApEpuyVaQFLGCNJQ
haedjTVQXEMxgrQUzLmrIFQ7qW4T8xtFIQmaiyqw/i3VXbviYhtApGuF7qwC7yLt
axSIu6IKE2finJEFw7NHZh0DAkgTdaNStUG3NLCwjdI4GxsJMax+E+/AkHALGliF
ZEAAIg4eflujtOPsvKwe+GmHsifcss9tbeN1Zcvg6huBTYxiT1LU1vdfmhw1vnQD
Zg5uHTLvYnIGz5VAFRK2vsMaVK12bnYYHAIKilb0MCYGZ66GxZdYJ+5/wUkxtW47
6U8LUUvpZwrGuQEsN4HSxtoqD0aKAf4q4hsVa/cxBO2SIEZm3acdH3Lqyy1lnlG4
z3teXIL/QUp++/r8KARye7fNMZmAXis5i/yG4fE9npYeX0VI9w7mI96o/g0Zg29f
VIx7mvV05/hJTLRVrayrQYnG6s7R3w+Fc0zTtt1R7LSAqYlSO11I3aFlvf3mFSgM
2DWAxG61kTKUIYuqKfuTPf4WmTHNNyQC24wvBy7NujiUS5iEMjcVXjTkycULI2Ar
iXBa6PdNhxQETt7CzmgBSMMj1O+o/+Bej89aTftvYz0rSmwZHujvmOEglZ3djSz3
ehPK6e5L3KKtV7S5O5OfHAm7oBx1GAsPKwjLz+JPTn0r95Dgmzm+ky9NH/WJ3uCh
fibYSggG1fHztjsYDlmAutqazKtLAkMwJfEemP8E3eSxtRzzVWOKpJwZWzsF5m9b
GlV4bRy0HCd2HllbZxwrjYN31xsQkdtVqAbSgFJCyyAoKZWEagU52V/9zDXoN15U
ZWNT0gI3+lFxB10X39bVZDJW6DLAnS7h/BAWXU1uXlvpoqD0h3MTbyNqghtiVhxP
6rVrfOrTzWkv9hXA3r1qX7EOMUzdNLzm+iFwlLhfm3LHAjOmGFSei+Ao2z69sbz7
SnJzcOL9C2qYrVFeQTzEBiM2fRmfk2U7cBvvqPt/a8BUUnzuPMBhMorJyIt9PaLy
BAmDw2C2MHQj025xTBks44xg2EOtalX3OWJ36qFc7mXohBSl+VlVgK/EkFHjwMee
Ax3x6lQVaEWelqjsOXkMdJsMc+EZEgwBrUPxQA6sCrqeh+ISndR7W9ZrYYyoCpQV
p+7FhFRm97k4x60BfIAdl4BPXYgGqVafUpyL/lw3/tOwfkOsxxcPnRIdBlyK7Gc2
KqBjAUDuDP5KhGZaXN1XQ0qVUbqHdxfJ3HuNGAQSZyUPjc0kSnZdbg5wKwkR/Rb/
7JRxMchmCY+9ct5ayBbT8c0MxNmImJ+kftV5IMceskYT7IGCKZ123Zo1Wh5nDx4G
2MYHiGaw8VI84PgZYWl6tbZNSpnN7Dib8OqFdxhnWd9jlcKh4s0gKzTpR2lfuwVW
Vca1X74mWIrTgBgU6ICMkHKInImvDDPPgeNUg1pMZ/zs+5oBjw8lYtOD02yJ9V1s
yyx3ljMy5Lps5zbNZ+RlQ6RYx1zUmE41+ak0M3lrDei00Kc+7SZJQ+GgsCKfv//8
vksE5T1apilsaGyJk/XOsCbr7LSghktroaJtx7KwMAOzelJ7xARpVc8jJApGui1N
m9YnEm3xK/we5/Sdhb6HOrs1jZnJwTQT5CL+H3uzRQm/7QFTfxO3mk2hLutrMQRe
unQQLKHYs3PCmFHMG0COrr2cCl0SUhOx7klJ2uP2zI3pkrDM+RjCnUUzQHbasPxT
yHs5iUzVI3yptAW0jqvMs0M7tHZi1HvDluYTKNtKkHMTVh9anacgs922L21lNKeZ
Ws0paWgZLr+yDZ0Tzxw7O55GKty9oj3rYURmj1J/WxQc6pLjoB+HVM3zo5DRs7+N
PuUiXPO9PO3bdloRVAESGz6QbsiPXw5Q3ibtcw8qEShy+T+UtzpkXH2CAkBMr1nx
ig3a0UA8hCb7BO5R5Fap2IpWh/7XCdfhAd7BKAOHiSrb6pajMCMr6yUk+8WCFXv8
N3/75U0+dTToYF7clNdHmlf7LDar09rh/rrBX1Cpml0ZcEb//snif42mryHiKTgp
/PpIxhYLxJ576H4hag20Y6OSNKTsNKvLmxeXSzQU+ZtjWidBpEqKdhtaIEYwywRe
JvVA6PYy2v3PI7NXLCA6ZjFyqQ8o2yH7LahdYoQE9VyFqmkrP8m1d1hu8dX5APxt
MYS9im0XIzpUtQI+CxOZBInKJQ3bjnR2ICuI7/htfiokrc/ue1MbHGdS3NtxQc7K
mavw3O6gyilcqEEXAJ5dg7fqRLK8rnu9z3YNU9aFEmuQuNlQJkbGJrrH8n5CXhBg
mH+19IRiyzveOTdMoH9Hs35IabG2KHcS6uPZEjUfrGC5kWs/4g6Iaqv38PAdXdw0
m6jvRJtbOZ+8653vPtiMS54qams6mhmj2+KcH7v53oxt+yDsHH2/v2/qDHLZ8Ncv
TVFMRCLX9zh2aODfM7quROvNOhs9DmnHuakqg+U8Y4j/EtLLw06FbfyYWYUQs1bH
zueiE5QwNJd6jjCo5ldVwj7BBir73Y5bVdovn2IjNbjMfxR49JV6QHBKnec5ku/1
/ncSwhzRbYnTH1N+KItwxDGjS1g8zQ8zfxHukJczAy2Qzsnbi5rlmMrj2BXGmwl3
lNjkLrcl+c86kPlDsXlzQoWJk/O+dRZtz0SVa++/5cUUZe/haxAnPaIOBvfMY1Z4
70ktN42gyeAPt7LzLM/oILHoslI2TLzNYv8BamEoQdggMRr+ms2oDcVVD1VR8ffV
CHD/seVsmQb41cgHMkwUbzTfzsQj6LCYJrbCMgPdMo+U/EpAD7QyZZCppMBm+jRw
AKSDnp+weOzd0H9xd+yaYSQZWW1df6BNogTOL6D44vX+zeF9XT9PQjUrIEf8TlcS
fRZqFBskkmvNE3Tq5zM1vNGTqnnIsISdSjwu0OuB2AKf/P3SJVuP/aNa6ndSJ06z
clckcbO7/BUvrEFJu7uktitGBZccLNlz7nBkvBoquuI2C0GsLUi04i3N3LzFtTQZ
7t2cmPoPlfWW7ShO0Dca4316wkduW5yuDJfRvvb/qUbpGnF5jpS/xKEb7Uz831Nc
GNgc3tez9K4udkoJUHk4VvaQoGMPjMIu3urYb5gc9OAKe30/J5K9+Y0dir+aUfzd
uimO3EFj9hoXz0+00MYBTtSrQy2ZLtDlfAINJb9YxFdAbBP9mvB4puAclM0KAE9X
msIzeb4gVKXhTm6/F+eYPNqX/hdKkve6R1P8KXIMS53vg3sm55t3cZVmb5rdw9sp
X2e88TxdDjq8IThieWWEoTF+XRXq21XJv+9mY66QuSd4cfsfudRPPEuKAGq/xJd9
13yAYPFm3tR6gmPMbp6pIqrRrW5ef+EGhrQfbN3U6d65lOYC7ioOHQxUv/HmAGY0
1iyuAikvnCOfEBGx6XKMWPR3p2vSVlEQJoSBH5Q8djYImGyEW5/XiZFDPsEVn3Jj
Vi2yTFORVfMheM/Dv1RYw/z+vjnoYXClAyKgspGlHa4/hVUatobKVV4l5QJo4SsP
xZdAGle21jFr7Iq1HyLHhTLmGk4s8vOpmaDfh0kv/vRqtLk/Kn/CJmnFTtmX+zou
vWnBn8Tn84OrHbB4VE+t1HUywGsljrE0bRC3DIyOUmFCLV7/Y+7ulGX7nllpR/Xw
dlmNX2NxApqO9M9cqGHcgy3N2YmbjI8sZjC78BSLThxm/7+U6Aut6rYdSn9tq+j0
Ly1Twp7r2p/Nj2ECH3Uozk9jCsQBdoyuVD7Ep3/DnOzD4n8KsDhIgsExPsDhf6PQ
SwJWQpuiSaVx5Y0uhmjK+SNaX9JoCkUVx6qxQM4nkOdPPULs9Dp6bbUmq8ldCtio
1Cys2gdY0RArr64PrEXebscC3lbcgd0rMz55vZE/KJNffRPM6NZ2lxvDvUGgdPls
lUpRO3/QutnYfa4czp+N+qIMJzbCSm5biidzOIxs3wjFRBLP84pyDzJTTzjWVQ2+
Hgd4+tr1yBJpfeDAiWC3jsHPM5Khr+Lwi+EApRI+GvkpxLxkndBpNT1oL1MmKiOa
b4XcdAK4iw0mtR/K1i2g/1RuLI5VuimlqBmt7FNxz/62/amJvnwzSQn0CF0x2U58
Ou7v/LGBJ/2RHcduGsx5S2P5r4KIlf/A3U3Ioa5b0pZFmqWgMsC1NafO2GbByyft
McZH2HfkR0GM0kRWIfJh+vYozNt0zZiUvfdaIbTjg7vKk1W1bFLLYMoSK1uyetQw
KeIbNtK3tJLGpMaLruKluRw+nozGpVbJjz/7C3N1thLM1pF7q+5eha5PDQgjZy4V
JbeWLsU9nY+I7LZ7vtM6YrDdpL+XUceG0EN177bfDi9yrIwot+6SRCJwOUxdm+SU
rvAM/9BBmujkidr6/83vOot5W6KJxiXRDtWto48xjYprrHcmIhYFoKL97FzcH8/i
wnH7OcTr7wwDNAYlZl9A8AI3b+G2hX8YjQZ6Yscf/kBfSvpu5gBQqakj3YyjC1Tu
jNP9sFoa0Zrw2XtUZIZuw3n8yVhgmzFLQ065Gc+hQYnHpYeqH7ueWufHe9HtYe4L
A8J4EYEezDsB1aPuoADTpBhyvz66X9WxcSzi8P/LNeT5+FmwHhjztuBmgK1G8Dms
o2PqvMsTeWFDNkpUIa02W+YAg90jL5J7I8/RtgPaeRsyqRpgqXYlpS5LTViPfT4s
xlFF5GP+8qXINyqcjl9QWtJ++xiY6Nn3SdOOExzgkNyJZuvBdlD/Dl5DiT5VT5cx
j4hrEkcuSNNiXKl0dhlUj7vuZsDyqQR2hSZbfA1RZkytfz2KqjUY4XpxLveStqNM
rkY3DdzNivzWbxtCPR55PR0OcPTKzmdZPreycjwJIdlTOq7IZfViQwpCwp9PCG04
7yqxH+ZPft/nr41J+mVBiLWlgF9ybL3hDzX8MkX7jA2DWUXxLEyr89kuFToWyVfu
bK8dPBGN3/7w90593CSarJVL2nFAFEhlhxdwx5IxR4TGkjPcJr8lptb2+afqdwOp
4hqYAFlhBrdsA4DaMML0vrZAYpZJ7HL7VyWhLmnpJ840B/vaP961vPlM6pG7h7fk
pV9lR213a7rue/nZ/u4ek0jksBsHxeU8T5xN3isxm8+JLxQtmPBCQC77mPooHL7a
fDaYsAIDTyGUfcXxA2zdDq9CpzX2jipkhamzXnsUzUDg/kLdKIujJte6fBh4FKKe
BhAORx3TRHzIA8wqQ2t21Vn3C24y0HfTIOQnMW5kqIImruGHSL3dRU9OI99DEB5n
theBboMrU9IKTn5fR9GhwJjuhweczaD7yti0j4Y/eGFnnDZUQJTUbypaL35UTL3g
U3AByWESuaeur9bTUrzOaopLts3YB7gCJAtFOVdi8p3vmVgf1QZ9sRTDfLFMesKb
FJaihI8qY2rm0anb+06zpUIArJpq3Y5doSGNDXGMa9QK6FeD+BfCH08JBlWvSJzI
kbFxbKE1S+qOjEVItN4i+V1+ZhemHf721u2H2cpn0qZt5Mcc7Z7i9grsNznywFKP
57wTcqXtG3DWspn3PfJwsNzxRhsrOIoRYYYXQ6UbBi+9D19k8YGDgltU5xdD/u+G
RfaStnGoCtALugZ4ev6LHpFBrpSU5pyFHtvn18Z94chjpxXO/w1JMZXedx60AjP5
nLMvcE9wQPH9126F0AtktKOSElg93l1ucB+1647VgEfEiWhI+eFpQDhqjjlGYwN1
/MoHL1kQpFby92reCRM2CEVMpDRxZkrVwhyLAO8XrLZUaJ5ANs08nvZmYugKFaQM
xUWZdlecSIZd2LKQ01ZdABbB1x/cd1CmFRQFD7U2yloIn/DIH87+9TN+zjceCw6i
kIvVnvDh/T8HjApE2kY9RpjHijP1Re1AvbMuWa1lIG5oCBo5NaJ5gFWNgArSlnNF
H8rgvZAPny/h0Z8AmltGREc4iRIG/s4uT+i2T1ht4ZDIB7XemOfRE5MqqTxLj+fU
dtmvGnG19K1IWKZHh3Z3qXTVNNYkgi0fGKAIJWUViv6/u5aK4my/tDlTnfdd0SXW
bS+3cxt2cZ1dMM8Yy2C8ZQTkBiH9HrnbN854o9Umx4Ea0QmCbF2RGtvA/Bwj96Je
dNB8jnkj4BN0y3lXvR0BgnYbnjzx6ntHtI8g1bbHz/WWCNqtC8bwleW1wsG5Mjw7
j0X5K3VVFvqMD49JLHYnDTNmtyCuj1einFd2d+bB8vPCZ/7Kg7bKNMN88AFbVKoP
HUNS+KoY9kxQN0cBa/aVhTvsAaATiTC0P5cOHPlzTIcFp3M6/k4kQRUHY/5UeaxF
fe7yvFn2vQbIthcK9nD0xH0iNwHkPRfguzmOAygSnbPjEKP/XeYF6qnMVTVuwls9
USo4k1nzRAsVFMY4zjQEIwOW3ZdncbulmAZcfS/588Ojbfe/dQHIjERuemPtugzZ
mMWrX72W3VfMFCf5H37EacTs5hKxTdHRin8A/ZK6mW8zhQodBBHOZoiHfh7e4+77
hTh47z45SJ5bpz0bshjz6nOh8kvGGqqUOwbhfxZuTjWMaHG+T3PPY73nN8hlmH8t
lKUaAnwPlgKUlzjxwdeOU9JOw9AQnEoSwb+rmrNZb4EcB1pYSuKD9DtrARqTJ3EO
RiOYqCTUFnr2rjkhn9j9jg3OuUwOP0KWrzsu0XrLatCFysvgXWGUHumN1n/k6iKd
q8hppuRksAPzdBXxlkyyzXsi98A2kzRlVZ1/9M09WDPu402gxBDyfPCG++6qEcvH
4IzvtnNN7S+u8TDPw2uIwfEfx/+/sYUdBgIwEsX5MZzmtrfZZiICobXs699CtbEr
bk5FHBq1t2yJOlJo+lkHJOXVq0d3WTrwUU8q18ZyeRLRgSY2rqtiTPrfloTLOdZa
AE9QzAZ8RI6mrroapGAkSoZUtxlJOX2oNl1Ivmbvf9FXhMgUxGBsy1Tng8vpY7Dj
7uBSuN5NFGTCjpqbuIraY8Pgj+Tosu2TC/GhjIWARNWChRJhFK7eF1wG8Sm6k/sy
PgyuQxj7heUxBFXH+fpgoj2B5Lo4N82pT+mIEmchbzhPzjr2MOcVXA6QFskKtefs
g+y4RV+4JdRzmkCjrZPlJfvu6Z3kpr0oZ2Ixr/gFb9hNOFjmTVenjPIKz9s1qbYH
C57d/5fD97+fFlLBVtjdiN1xMZWP7Vhc53B9Ta5IIyU+AYqYpGqfLSThJ0W+Z2T7
1gztdmGXnPLRM9nb08yL/9hyoQlwySJZU17CmOnknhVVo7nnMOQTqePlEYdoLer+
Qpca7RGrl82n6HLNfgEjA41BWeJcLxuf57Awepfa3c/vHCjF9eXbQjTeMjQV8Yaj
aW7l4ZhKPxalLr2bjabXzKQJQXLFvxmumyESBGhWAurKTZc0aPfUUXgqpgauqd46
wpqGOl/8WDpXFMk0MBTiA39CXbMGa/mJPtU6bQB4pIDPoYp8rMRHdpZy6iKh8el2
G7siloE32zt0quVnKEW4/v9oXm9R9XD5ELvdNn9aHtdXe9wNXVWN+2tOP0Rl/aGJ
vWZbGt/DjNOnvgaizO9PWafiWWnX6KvGvAQvB/IOe0m1jrvm9pM+z/3TumTKpTvj
i+4iQI3fdj84n2xEY+hu0mY5bGFyIh8EfA/dS2FupS02fWMeMnngFCSIwQMJ9cmy
WX/PBq7da6581Le3J0wUMxVkdV49tA3Ej9C/XiP9PimuQkYtwcK+RCXWnQ7YwYOX
iI55zwNzVO39r/uh+KBEh0TQof6Cw2YwHnvuKgAnH9CRjx0cR2YLOwo0tlADetK3
oYiXb1z2aG8zMhpAP5uCaQyyE5WLRwhAXsqiEnH2PPWAHy5PxgkXHrgJ09UOmMhb
Te3fAl4puRBaE8WYBMsUHs10jfsb8wwp4mxv2jSFPh70vJ/bXdBH1kmJCEmVXAKN
/vdBfO2aeWzBlO94NuRev1j3iY8p7qXe6vxy17xIuGDt+3oKsZP4QF91HvoDralN
2BGTS2gD9/NVue8MqVaWoXCPnJcXpr8dyZJJBPX1AXaIuXj3oao45gvH1oAQDpNh
g7GKG6OQaCjGAHOsT5V74bUSREXBMO9uMS8tFV8Sy0D5YcLgHHKWtU2oHPbgX4UF
83EsTpUX2LEj/gB4QgvCAWtYrVIPxp6FTIxbJLTs3gKvHRvWILShlLhYqF0jYAOo
DrJN94MlafNjliQKTE8HKfH4Z3aFYuZ/aENiyCtUvgluS5fZnLjd1A+bTmA+rWOG
mvHlog4OgNrKnuRePvNANIuoZ4nbqQc+JCM1mW35ccsNNLlRIA2VnLkRdmU0onCi
eBOTmvbl7Ld9A4tAFoPfIk0kKH5HuhB1x8Vjcet3Dx94M+TBMGcA3fDYB/jgjvEQ
mjUkHo53zwwbajaibyrxzfykY9eg3U5jM/lkVDeCer3T3zhUeky8liymIuIuwMML
Dsja8KNhjYHdh52Se8gb6geSynDjwhHTDIBeDdH/viAdWz5JcLK8RoY5HQeK/gBl
xYTxACgyZkdtqKNN+ttjMd+of84Ycg9nghbJ7VNTsjM6Eu9Ik2hOigkyRIwjtn2N
dPMsEXEeIN0vFjOOAX4Vj06caGR84JzRrh5j5l31a13C90LvIHnEKS+JgmwOH+jE
a1Ac5qJyq9uVAT8KZUQH3XguNFtYgv7Il8CJ68/DIVfc8JrDx1N3tSsZq340EAY9
bI4HBR5eVsEzGyr2fyo1aJCHVglJ0MYI3SS9GWicNL6eK6IEG3viS9TgRu0gbot3
HLH+c99F6eHSTPf1OrjPBhHdZlIN5tKHZXvONqse3/sbBX86b6DXsYq9i63js2wU
4Ok0DAMT9IwRRDYENlBLRWPQl+6ISq96o7isynGResl9iBq7qVWMatp2KNOINTjV
wzM4wlEgE7jGdwtuYkGSPmIiZWO24JAB7iLj0QORWrbGJzyWzixshFG9XmBfWMLq
nw606gQKcBKpdrMRzbNVUZnLiFTbQgOdgBAkAkZTxCiCJc7sN+WwY9fVWqsYNmAM
AT0gmz5ok+4K8EIO8f6fdDsJ0//Hx994iydBFmdgjBQxJtbM/8hqChJcl313aCWy
hwQqyBGwBY7D+1nLwvwVzh8jsZEwRAlZmhEHnGajk1bAwosQG2BErT+hCMvuUY0i
GW4PGNnoIkN7MbvBbgV/qRwJ3W/Kg0A2DehuH0GQL/IxgII1eNFSUDFFS9EIE0L4
msndaiVgN9K+AO9FLTKpwvAd5a0C6wdaQe/ENrs4xJIPUW01Xs4wEyfplAGDAYmj
0wGfYXsvpgsJ5rhmkeKJZTKwdfgmGv/9RGmGzuWefTzPN7WRqOBLDNVKFxrTOPkS
Zsp/TpgLUwNa+/Ex2VgqW22X3FUbDG07USTRvvUzIurZbwAW4UB+46vhIpuWe9Wa
VMyASQDnr58lItTAERKQI21UJ2szcU8MAzy9ub5pXG12/y6Jh0l/Hj2LzLNnZawP
1cbGQ+5GFW4JrSnvBT0+XgE1OAiA3C/Wrb6MxmTICXx7rwmlkHDq8bogm5/gnPly
3eSA/eYOmYPcWYBQtmYrrqLlKsa1w1Qkj4TWLxFzMtIVnGM9A5jR18E3/YDgx2MI
w8W2b0QjV2HlpHCwVsaDslhUbIU1ZUB8KWt2X+V0FsqdpEu5PkFcPWX3v/JgA0kZ
ariXqJC/YSZiX7PPWJVBG2iCEWopTP9VDKGbokMmY/Jihl8U1AcTpFI3zb604cY+
Lpli5ozQnRfgyNh8A/WCf8W3es5a54vqlFrCMFytguAgS1KPt95JLMDLp6ybKJ/l
lnhSNz78N44SpnbwWyl/hKiF2Ln4p2ci3rjS3+Srb0s6F4R2gvUHrNaP8GOHA8ex
pOYKzuf9JO93sTuXhGg97ldT2OeXetEYmOANNB2BGUya837slIkOYN9voj16hAIX
ESWgD3zDE5zU0LNgR5dUv9geB0nQN3DdmU71X9fs2AcPNixbo2MiBmTNBgGPgldU
8M0mZ9UCY93y0rdZp1cDU2MS4utkcKm/6xgRLav8H7V3xjzk49zZzd+eThj/Beub
UMnb+n/2dVDta6EVyOdqfG7+GipDRv0G2JK/MqU9sEzlxw/NvGLLl3WL0SRlbIGP
AC89WKKU0Vy2j58PsvioeiGsY/HDfOFB9LqoIDeH0fOg/4kh7q68wbssuF3gSuMi
1rz2kFCImUPI/hwhFP92YwFZqe4iI9mx4XBiDTV9+lsufzPxtu+wd18KJ7nVYzAN
bsXb+B8qrBw0Hmjr3TvMoEv5rh0Vx/p9jOYu3m1eg/dhN2Fe6RPwkHpi18Cg4S1l
0pEGrUiEVK+c7THhUPam9pOrBkvhzPGXZIxkywSNCRCjuWCcm8cjL3vHeG+WneCM
5xomeN8hPHKHY++OJWZ/+QjVd3sOvAR2/4/cUx3dBrISFXZ1BJBx6zeaP/aM0KL/
Xg/aUha4S0GiWuLyvc1yIu7gkovGtHwXO9zjuee/by39ib+vUlvq8FlagytZaWkk
tckBdog68y5nTn7K7BSKJwVaSl2mJepeox+f8kx8j7eUQticMApv/L4fbf/PHRqw
ioN3JvtbtSatO16+pjqis0KnB1Hsed30Heu/jFT/aBzThkErzErPpwAG/htP1l8J
CD4BZyIq+uMkpNwTUrQC5ZzKiHLKYo7v1LdkEhroXfLUSYWycjg0qx4t61OTWpkZ
BWhEum/Fa0gN5GzOg7su+7uj94bQ8LqJz6mN5xkVmJ4hznQBo0nWPFKn2YAh+4dQ
KB9Thj3YQqlJVtIeOui1ktEQzBJBPZkV/xhg5QuczOOcBX4OqN4rc9K94GERxxHC
Xq7oWcJj8AJxfunEsOPjGjvsMVVxRKWc3OmX5et6/WlXnghmhn2e5Df0LSQOFY0e
RonmLyLSVhvQnVMeGNQkqh6Y9zxgQCw7Fiedkp3cwbZfjK4KujmqJB+iZP9UwwgB
CJQgUozQFnYxaejKGL2USS/IB5/JciCViHUyG+3xYA8NB1uMhXElT3bTol4uGcJX
WkpjqqlV4Fco8flWV2oy/RNCZy2P3nj9yNbVpWVxT/cvfkuRewNQ6pEpxcn3Z8LR
zkUMJaxUexEiXW1WJSRmVgtWSswDi537+iPr6wYHvdF3a2ZIedDdgWgL9SeztZF+
bIqaVKSibp3EbDniMAy9c/wSUuzSYREEIUbGgUOEwelRJhiXlsoxZaxRCn1VzyAd
mZjzJKIfqlUyK2bsVXsMe2S469ZtMr7NwaOM0/BDog2QcAyNdsKw/fIAaJa8VYys
2VSOg5TqW/d8v1F2hyhRbDpDoTVDz/fFjBiopZKqZXvfrViAf9E2lO26KdLL7PgH
AH3xJ8ArzhzVn/usCH1d1EKh5sfdmwR+uxNQK2Pxqo3Wp/P3l4z5j7wjNn7E3Sru
AvpyLfH9wL+is9axamt81FB8fxHotQletsohHNNUquOhO4c2kgzHtElKOM0UTZHf
ROvxrq4L2E+h0ZIG9BpCRznoVkY0Cl4bLHBqz/LettJYbPw+WAEQAgf6V+XVFNlH
h8TvEm7HpvGFfyLEtVUDqfEFfzgGKZUC8a7nRB9jfbLURlN3bssVR0frqSWjroos
fmF7PEpDYqlv/p+wy5/vOTYr4UfGdYcjz9FNswcjbqn9uNfonqKxl16NQHuMG9Dw
GZ/VzJYvbDgg+/Fb5haGpFfVttL5rRsz2+g5/UFTtdg+WcdGVKoEhc2b469EodM9
ZdpnHEvVhrFQN0rs8dSGBAWF4UH+/Z3gSdUnGCins/vw2Pt/E+Nxp7DaaNXqpt/G
dvB5dqrCHCzFlOG/QeuSEalpnVK3KqZvNxjw/S/F6RbDYF70rzqKKm1lVNA2h45k
FswvVCP36pEL6OmNR8S6V7GeaerHJ2j6a7K8zk3gGGz+mUj2qw3yc/ZYk5WSKz2z
CK97lwP+6IgYpYU5RFORR672IdBWN90kXxNI3Pb+KBlq1VcyfEZUJZpXYCIoIWY1
sgv/4gHnK44TLR/1e8jqbyrVcUWs2QuJ0vDAKSPrRZsvdv8GSHWCxCAwpjQV52GM
BfdN6hlbqUzVZcnrzaa4OdgIYto7eZ7i7lgYmXse/0euMpuLNvxzo9CBANgiYsvJ
R0JmUVmusYtFIsNU8rUuhugl9+KC8r+0clTlMgr0Ua2EGsA3YtSEKeMuTkXXY06O
B1uWBknWPNrO9yalNSxNXUJhU+FMa0Ph1pYn/xiT/c/DtcMkc2fRZPo1adUqEKoM
f2yr+M5i3qjrkMyiC3/fdbuvUbqAnfWmA62UN95HXW+fSO9J8atveHG+ME+Kyiwa
pNCxS1AZ8PNsDH2bdi+6tQZnxZAXmJ/hDUAQIrlpZT/peNroGF8rtmZJ2Q3qmKF3
a8bgcDuYpu2VVcnFnX0Pxqe4MbQ5IJGNFQbRLJ7kqvr1vQY+yLQGGqj9xOMgME9A
+hi0coXpgPs9AMGA1tnKGPcBl28ItkpxFuSM7HMgBK55B7/SzhQg8Jbibi8WomFd
t88stDG3g4fuukr9jxv8senbTtxNxpTlhrCRrjreYN0+Nmyqzhigw/osdRTw6m/l
FOJBwJTt72reJavmYDgaErSTrBRrtJBOv+35XscA99ioANyTgzTplM1Fa8gC8da6
MYCiRSTS9mZgYc4ZIfAlpdunkMkmK9OM0u13zaRUz+61dwyKJrN1pqbdIfKyyJTY
ZtnSJjzcre6BW4IajfjSyQhIUDF6GOTzLyssbciDjv+kVAgCAo6cg7UMGhXZJTYn
hNAMQpMNBfkAzY8kHwh/NkIBMD4tD3fKodHQXhl64VsIVlOp9I8jaGTdz2ef2w8m
TsrQwpsIyqHvhuKMIp+4PL1cgxFGdtxq6WGy066rBBHE9GJUFvAYxeeNG2R7sAG0
RssmYZ6ML94YMGpOsfH9n9vQvcSQec74zcBDeV7B2gRWhHhpZcnJrobI96uJ0YNL
tzeKSzZ50UCAk1talnEIwIwUvV7aD/g5Pye4sVsOP2xBDdh/sXls273au4sYN+Xh
3OQc1utwcCy+fwkljdVRmGJ/jljSTBAFH2kOqQTlBe7rTTpt/j6ogLollVsRP84N
07LFcVe1t/AA0ta1f6CODhUdSlR7Xjb3fvxHqr2jgJcclsDEovD+L9oIxk7W+wwy
hZ+S27YsGyPikjJRw21L7wBzdMhMMwgvAYUv/l/iMoH1G/KJQYOSY9avWpTvkIVO
Yq3YfbHTdNDZTEnegmEQ4LAu94V39PmkuLGRl90l7jPd/hu5uth/4G1qkcCLICUM
4VZTaGbyupS/Du78w/T1vjG6/99wBCB/FZDkV6j6k05PffrJYunILAKyAFxMg3JH
Yu9bE/Wdf25JpOCvdV+4OA3iq/jtJ/DiS3WLVczVmYn7O4SQgdVYfElq/m2J2FMb
XayFfY/Q092hrJukhtgtxpU6i1n23Bn+AMcsbj87qzJ8MVa4YIIumUt1C4pE6Tf+
qpQunUD/VnFC8uQRhXd/DcuVNAGG0odovizsyjfumtNVoNjDWqfvyXI33bGGYgKi
ydb4r49Cjnt8l93RTpZlUnO6cSkPjNcHKt94YXuPACtmeH3g3bB03mSFK+IKJjkB
mAy0a+OD53qrZgZ/CISdruRHT2tYasx+smUbSpR8mskCPHCkAtk+t3weHkojfxmc
aHCfjBC5qKldKswJLpjr2mGxNpSf4cZQhl5/ZSRXMNJF3I8KvpTuJHfrEVydhUln
6BNuqbKDvLz8Wdf/dW19sF3k/vjq+cB+Eoc97lZlnamBKJnXRNbYrvtIWJqpxqo/
3v6kW8paaZgnUBX7VYEqNOW1NQHIS66mqhLJuP94BKgI6p/wnCyJvpJf15+9ydrZ
xLa/Ngkrg0Z+OtjNYC1GjggoP8WjxjZNQZyojYygtENRFPEcVXcCG6rDaQAnTYlj
/Snp3q+Cx8QNm1MbuFROrE/P02p0RE/jIdSVE5BkA2wZOFRQRuHrSOnR462vpYig
vRjKuF/iBL4zTRoIdyzE00WedFFklR16zGXQxyxcXS8il93WNtWdfkwuv22dSc4v
mym5k4WiJ/TZCmgBrBRhWSOrw6QKi35xDctNyE5APq2SioUFa9ryDax5as6MpQ80
QD1GdCC4N9zNIe6EICtLArOaqIyarcYmicRL9ZMYnIEbDNc8natxbUTsvxJlepd0
MPqB3EBbiATAh62A2lNSi8aZtY10vIfe/K3OhbLqIeaHgaf/lRSeqRLMX5IqyOQM
ZEcexQgEG74PxOZ9HQwKSsfCvur94YvBzmDb5kz9jcxAPgxz0NIL8k+ISs1VDQ0v
9pSYzspzz8BIi43GqTu8Po28ouzM+TbTfUV9VKrtAOOmmUmciojhgIiZ4hnqClKX
/K89AUFN+4aTN4HfVHJ5GtoWSYs46gj3Kr0YDZfbxNGmW8pxGbk50F3DQMa2SZOk
Xo67JsR+HHTzLTBbNT1L+JFVnsTWvUEKLfNUTpE3f16VsOsskLeKE6qLjUc/ZO1i
oU1gYn0J222YRXQ035gpG6hwGnitZsN7fPyjo16Ct8h/rFogK2fLq5EhGrs9iy3V
GbpXYzsAk9takAuFtm+Ls+EOoXTmzilTudAffc6pVPwpWbxDiHHd73CcIOlzPGvs
PQQYmnQMc1FpI2xpHg1aleITbezdz7nY7AmrHrmRUfKf/j/xwPIkgf6QQfhF0iEF
akR3SbW2gwMjySDPgXmUkNb4doMJsYUlETPitOUWZQqpGsBikLZ9DqwBsu182XGE
b+hn1RQfdyk7mItlC++Jemkz6uhKYgbhO6abvMFov9lGjFNndaJrM+quCFnRotq9
M6CS4wNk92q63t9lFGbiG3Rr/kY0EywSXuDBJktpqSLWIIEYiFIRJY4XtfcG9NEs
XzZfpOtKY4l/LFNkt8ZG/DXo7OfyHfIzqUnar7OKzJUE/uro6BZglN4dwdom1psI
9ATd01rurkQuw7/qTRqFUyf/wikvX+ulO4v+chi/k+1uYiKDvIgInoqoEr/+2eNl
uOf0C1k880AO4kl3Ei1VQAS/I3VkiH8vs7FX6rijp8pLIkRfO1TBtpVksX+VxGBF
8PHp3EI/h50Jszd+u5qWpOmUdAK42tlivPwLmpv9t6a6sKv0eylP9wlURTpTQGrS
i9sX5783ZWzCTBbeJGAqScYpGD+dAW+/bZmBdtVNp309Q+63DnW7XLQt27cLMIYT
ZrsGBbmm3K+0PKBycJmNQ4kJiYHHpmn5JdDeNr8nc+spv6wDIMleylrMcEISKZL7
OU9mzBXD8myOTzLpiTwyF/x9bPyX0uWGPjn7DtIjlLzR7VzH+CymLyQHjLA5MBbe
ZqEI2vxB4M1c26hU7xa29JHB07Trd+2Ku6EFvsdma9XU2U/Tfk0YsYheNWA3VPPy
TnfNJWbRmx8ENe7l/QjWMNq3pl+BwaSxifKem0/IOuItusyaAg07BEF+Ft52hx8u
4sJ5XoJiD8MXUQL+6RNGc5IkrBkXiVvM84kzdKODSPxTUtHC4Q6CIKUR515Ah0ZE
yFpBw7A/JcgnN2jMAFgf5DI4cjYXGu8ukXsEn6fcJ9AKklU/zELLRnA8KSrc8cXT
011CAnVz7P4ZamS0duL5ZHgy/fkXMghRn8kdkhmL1Yhf3IE83oZYJls2QkencOeo
OsyUS/KMzS9JmAVOGH6boXLFa75yrp3RWR31TbQYa4/8DVDprGHNVgY4YRc2e72z
lHZ1I4omnspLJr5rvDV1Wkz6SpLjSkuacquA+vQ5Q48vvWOraeR/zD0k3Ie9x3MH
G7jzXyyy7HfKjStN1T8B2BPXUH9TIXBhMhUbhyLWSDLtD8Fq4QFvVsiH625KpUTg
SWuRtmEmeY4bdc4dSlSLTJhOe7vfIFRxYeoRWt3aE+A5WByw91riH6utuWbGS6Hg
JAFUdmZt5LOoFDv7OlSdmKh+k1NNJV2JrFDb6RMltRs53IqHtNTIMMR7WNd37z/0
cDwTVnjxwsjDK7XRn7KEh+5hZ3C/QAmOWBAH0RcEFOtbgDwyrXgbhjDn6i0RadLy
T4PDfeC116wF3yNQxEIJrgi8NKIpY9512rY63djDfiAHSu4STIMSkm0KaYhlQG2r
xz4xGhoydK0Bn+HVdW3Z6wX7Bs9mYt/5ZSg+W2wiGoc+4LMPggpMZQLll2JpsOC0
XcX8rAtGgUFOb/OHC1MmmkOBRvt0x3/1Jdq2NAEFVULGjX+JhqKY/WUJM0NPzUxC
JfJIZnsAWmJR0YP26u7eAi95K2eGHQ6xVbb92+dMXdWIgA6OpDHqxU8Ny6qTGFXV
Et6BTcqqGDZog5ysjNaSoYVxcShto3ZGEhQYHfBr6BbK8usVCUdJ9HcRYV6i/bvA
0wQog6y5UcVetU6SR47qgAIb2TXjer/qDM2rt8rYy0qOxjOBAz3KpDtsXr4H1Md6
cdiOMN/h+nQYUrZDEJv4kjDS0R1Kpi7Y6DBTM5eWpW+bWqyjOyCnHx3ofYV+MPhN
K96roJN4G8a8s3Os942Dc0Aw05xlXZBdcOWzpB9I+vOKEj8rHAlOAWlcI12GV78w
9dADkn1rVeJUkPoVKjojM6HR8wjkbFNwpsVq+aPMQPGkYypws4FeB/dHl5upQi+T
NOkYppE7mh/5/UYdbXNklIdEHlLDDnCSDFJCO7w2HERuuVvpgCbL8p96zsF0/ABM
t42UueMYueAxAFceyuHkXcpmHNPhPxlMsaoDSctTt5cOSFvwk9ykOoG0w2b/bwcB
BRMogYR3eZIl2MV/4C8lislH7hNW1AJUFacmWfNwga+7S4+ItPZ4hm7/ozDc3Y/s
LWbDuKXV3+4pYAPOL/QalVfWOh4OxL5oY6WN5buIDpwag/9M0EW/MI07HbIGUK9A
36aj/qqxU2qCsBwkln9Yq32TkNmZy0cFB5kPzVtzOEEGQHsmvhEDM7J1MBdZnGdV
GDYQgmvYKqtL+BuswNg+TgT3bqQHbJrcDgBmZPPjBwo2mBDF6wIuT+w+WMht/aRq
zF4F2CRlXAt+wq9lZ5SpSdKGk/xlRnklA9Vd+PFbGI3gheprhFO/KMuE/NagxZkh
Zq366TQU3rcW3d6oI27+eUW+2SVcFJ8eGZWz30eJ9Tynvq7sE6+48Y85LBQRDIxJ
HbkRHDPxMcWvwU8pFfjUd1PFhQ4mgy/cpiVXwyl0fKkRE2jG0nF4esXxvQSEmALj
3Nh6x3DhcAdTPm233HuoZ+ZRk5gXGzeF2ikrTRVYpeyHa/6HeqYGYjhhKeqvbGg/
KCWRL05jHPpgHQ0roFUupCRTlFuqzmCVXzaep8v7WIPi5jT/Pfp+JgUoD6Co9Vw1
5on3xSdZ0jQ92GWrTmNhpcu+AUWX+bEEWVb0CPowYAS+vP9wNC8G+eFCHXVrEjHD
V09OH3u81dq4cZ7F727/3wNrlBdye9NfULJGYqf29gWaVu6rMmZ5VxullETiTBzN
DfZEbxQ4LSigGFvLr7t+ntrKPP2ICHmZKusfI90z9eWlmIdNyVMmtpafWzCoY5pW
v1BlRRuAbhDWze3vhZGvu4trVMh58gEi+15LQmkGOSCmXRyi6PDZVkSnU8sXuLK5
ug3lxGvvNpLfRoWVo+Xb7QYtBk0J8mH7ONgSRGslRPR079O64EMx3QyHyT9FVdWX
y5X9T89/L/mCv6I/CmYBmIgMzcz08HkdT+eUl01052ZrkYKPERwnWW0jkOmMBzgW
9QI5ZLcnOsJLeGpri5tEyLs3cVjKR3WtloIz80Yzy2e2exXBEmR71G7Ewj74Y55p
9zu5m8NE8iKSVGaK1+KSTMG8zSH98S/j1dOurNUMML+MuGpnqRa1OyYp2R9ZGBDg
vtiJ7qrcNp2lvCqmPwgZr/r4l8NLvqnj/nJEkDGRJhtqvo/iL+ePnY7ec+9k9++E
J/nphi9WtDXyiVnndzeiAIn3AA85PQuNbh3dPOljT/4mJW952LdnuFt53YJfOq36
6bU0AIM38YGHC0He4gz66xErbl30N4G3IBHQ++86e6rLMt29XHL04yKap2FkV/W4
rzQptIjc8Nd5Cb96srfj2cKDZJlyHU3O2GkmJLH5128hEQfaPTuVT+V1nLnWjzdn
0XHghgmWpTP4Rr4cxhPGmtThLqcRmCdZ08WQ+CrKMquIt7frCQwAsHGgUjDkCY9G
NvPOSezPWhg1HS00akiiis28+31SdoEeLTl9ytKrp6gwLaN0BE02k5zkJu5tirOw
LIEkyn4lUwm6d/Xy6BBmrtfYcWX1UQUqfmGGp32gS579XtX7Upon8G1lJBXbjU8w
WARAU88iWx09WvbGzF+OEjq/AguMTSpaZx0Z8HApldJdPI4CVhB7iyN83HP3CFD/
EBdAc86mzAZME0sQYA/DFT6Z8EYFdf17EXwA8lyB/7U2XiC0YtOoAqm6JvkixFcp
+7ZYXHgWJxbhMx5D4azMOqg3itI2v7k0PvVdx8b8TU89XEBlr0LHIdfpL6OMl8YJ
2UcEkhJPbUy5KSuvX2WuPuIowdPl/+1Q1IFmKWim4Idc4whU/6yrVIRfRZONM3Rs
fNfpIcDLjJ9YcTFieWM/oZjX0IA1tYlB8JabFqj8JzgYogy9Ya4bh8/EJoj44NDk
XGvzGGGHenjLqdtOEFzAGfLQ6cZs58NP29GgHWC2MmZj3x4Yqub9lEZjdZFF9mr5
GNJOydPfq0nUEX6ercF9yzElIsK9xBjPVsAUitsEIOubbVaihpuHlIdpxfACI+qc
tUZZRM9Ozhyw2lPP7h9mzMnuOzqnzYJ22CjFxGUWojsv/t/R7xBP2LxFLSlOug1Z
91wAqu2rmSgFhwvziR1d5DAiqXBZ6fgfHHDHRpNG/P9WjY4a6xJwPW4sdy4a1QT3
s5wBphVhm4ejBNf4b0uO7qgqy37XQu3JIa38t6st33mK0Vw6COesDctGQl1T7htJ
D4wNZ4ih7DUO9rgiPDEIHB5X7veHoDYOWxsScSKj3XyM65KgjIea7QlMAIZ8jmfn
oVA+FzSRSQQIR2x3dhldVfbMzdaX1x9gPBvF5bJSfdVVjXcuLoDzelhTrbbqxCY2
vACkx+9+PGlq8HSp6ZaIvvhyv+OI2gYX+ZfRabY5lNPnKbS1Nr6WP+PKEABRLyUO
64TfJamNXyQBxDnqPLQyqDaK35ag7KejivPbaXYjC2RwoH/pj9Gq4USAN9ChspjN
Rm5NO1XWvYA3HyHqK0CDbw3lkTTFQ6QqBo9hYpcQMoEgeej/mRdzAmAo1xINpxZV
Jhubr8sHnlO7atDdOZ/pUwrYJzcQGZEwY6HDbT/1cB7Eno5nzGuZQZFWuVYk+DbH
C/RLvRBDEfCxCRTfas6lvfN9jhKRxmMNGxPhoBWE+sHpdlxVoT1RLamd2sfQ92m8
pPND4mBhgcCUUuTCjTnwZNHapi6tHKAtwfJZaGjRliMzFh+Y7VzqxXWtTqkoA1OJ
TDVgGUSe4HAUyUVQL2CvwogPGgPR67u5xSDhPkqz45wes5sG3b3KgwTcEKe5/he2
ufkP1oOLWl+WIlVKslbC9wEeieDPzCabOS/fpEedhS6nJHm8cN4b4QYHcG6z4983
ewlhk4rA8EYRtUWX0H5pNeob6GkfJGpa22wJU/Uirn7JGNarBmzn+yCjKqF29Aj8
tauW8pdNIRECzGcGCwzvizg76vehqXNhNHHJquMB/czGlxQVSuZ5FMmYAqr7NDBt
FxU9VOXeq+/IKKUYDII4Wn/gY8rAXwAJEMF3HLJR1mEsjAGvUhwu9rcMt6HWobxr
yyULiMnjUpauSkk+pH20nfXMIvkrxjFUlgLCE3cKbhJzixUfNtr10aqOMcPFs4dg
Ey1pw0E5S21/afZ4VYWfu59eakorIjo4KXIB4bd2G99jX0kd9wWBbGZyeRR54z4q
tXQSZ6FJuCjGBTTb5+dkJ44DjOwkOHktADxzTEPq3pWVRnLF2Y7G4Wtw1s/LPtBM
XEImq7TmeQV5OoMPjq7+A1qFW5GwEpBvfpm29YG0y6t6Cspehafrd7mB8nPFv1d2
4dwEpDELF5raeILbwxXM9PzsNUJk5Vbu5rqbsSWVvmbh67sSWsugXP122SXf1S2r
TbNv2+F2j89vbGlCKUlWi8+Xhf4FQHc6OPNXgUD1sxMnRoX5WV+TlQMUu+PfjbxN
3D5LFrxMIwSE1kLV/KCWUMrEpxgH3DIqeoD8BlIIGdk7QJvifOL70dAnfkHAY2M0
c9yikZl9VuG0aC9VmSMSTs+N3FHtnj7AVncqXKzwOO2n065iojmPsXl1If/6uAVQ
Y8k3NR9nOh17aiBfLak0dfvb+mgQEKgcbFzKjCSds+83tdjSRIRIZUyRDPTiHw2M
5UDfWhLZ2jh2U7kN9vJ8DJQPleutAs8WdTixBQK92eRnPF1AqNGPcvYjcgCk2o7+
kLc3tWCm6ZQYZZ7tzNwH1kvo4vg426+ZvERjg8CoMXIAAtvZfgRQwgrswkM+Ygpr
Geiglu2rWmunX8hf2EWDTiDJu6A9goW/QK77R0VTWH4vInGEiuQ01dqTV5hoJ6+j
ZWZdvlFLtEv0lMR82hpWY17e/7qF81OzwsTVvT0yEHt6O+JNKZpbvjXKi9FGHiXl
ta1YiKpOiJm0y0H6bwrW6iKZAiS3QiWt4Mb8P7axIW77Pljm3yhSTpgPsgC/C193
Phegf0CbTRJ3LhZwvhwgT5RMSNX4iCjSRwUe1ZXFOKi2KSy1q9qbtA1WczNkJMyP
J4QPvKdD0P1MHxKptiWrxf5RiGAnIDThNfBE4WBoaoZV9V9rhJug2OC67ar6qWC/
1GXJkLW5RgKuFyngvjBil0osR//mKKX3afxGxYaaQibO1Y6gXrxZN+EoIRSFB5B0
cBeu0IR96YbYOwlva1/uTAxl2OZhYKemeoOaLxDv5whrKVWGbju6S5BaW0zrN4Yh
VOHxfh/Pda4LVajOjINoT3DyPonDI4Vh54V+u0gewOYuKlseX1wQPKwawGe6BJLe
BEH2LB1mGz8HaiDZahAy1u6VYG9lkn8xjJEknKKiSVOrRo1L338dphtf0Luh77SD
QVHP/Xclsibm+qh0abMgBrAJEuHK9rfjydY7Sa2UB22+p1OwcDuA3+CJG217BDzg
vj5plQ27ts+ODxSB3dIXxCy/VCn4RFA/dxr+Eg1RMmoY5B71HBrbSoD/aaan8lDI
rM7CmoEiktyxDpBd/Nkd7JAM1Fa9SmksB3fD9IvL6zytyvVogDIi0XWTT9S3XaJi
T1AV790YZSpgUclAe3o4Y0SuBzOGps0gOlfojUWfNApmhDmtMc4LZkpqdJRt/fbr
bUPPpqUN0sXQPonSI9achGDw2tOk/fXzfZvyiBGha/cYEqPTRfsEky5aUDOG5VbK
swiV7m5+s6wpkaJaWJ7y2QvQywCg3igZSpuBuNlN/xbhTuasiGP3b6kCU5hqxkP3
NxWi3qJwYEj0uOwjz6pzCQ19e8fBI7sCbhiH4Y3nupwmdN3axc9KQ6xGLrkn5787
Bs+oHjJ3EzImzhYpUxwosWODtSvGHLOz1I4oDSX54ym/gsCTh6yjWwt/eVWC74AQ
H0GwAGQj7SnzWhyxyQ1X/eC7wVaW+z1E7xUzGvpc7RGzAry5MKxHlTOnGYVkDWG7
84T2tbIC8DxlMsRu3N98xEaGr8RSPwHd4hOIQsI0QdSpowME88KyiDlF0RTiry8t
YYM+t6rdPp6SRnYHmYHfcRBWJWheulZoEHj2lRS4Rnb2rpzyFHK6yTMvC9kxY9e5
6C//B3iKlTCsJPpcT84UYgFguH7yhyP1MCIhX5H00s8o1h6DsedsHWpRgyOJ3pwA
GQ2BJYIChdbJ8HvYZVvpTzG+SJt6wX9ZDT0yVsQQYyzZmklOPILE6nFq8I2kXTEj
4TDXWueXj2JHQyGuAEWG2PIdg08rG5SYyi3Mst9S8BAKuUYkk/asbxfO4zGPCUhT
bMleAi4Ja1TjebOYugWjLs9zEsZVEPJ72F/4CgN1E8yUH4OpCpVV65sFNR3N2jTW
iidmPpfhdlnbMdGCyE1xDoCTO8Eu+BQQo1KEMmZyuoCT0OufDM6ctvY5Smg7jq5H
idqKXkn6gIUbO1BP4oT2B1tGqso7FQj6/PDEwhi7kaKGBiDnA1HTn6Sx5ETRDfNj
MxeW19izrTyaii4EVK82TthTkU1jzwJtEpbre4Ly/TjLfLNaPcgcPD7XkuIUK9db
3yWeepc12YSIFtQWiDktvYIocYAcCDD9MeRzouanrEiFVYMXgtFNeG6vnq08+miz
hYaoTmfLdXYg/zPO6CcgJW+rHkq1ij2+DE4cm6nxsWdUczvvXF7hJ7twGuI9cF/o
rHH0kcgwXPK4G5Q71DblsOixDt7TUN3BC9ttxSEi9NJk1OBRaMTvTbIbpbqFd/Zy
MBkQcgfdKCgLu8ZUkTtcyGOJmB1qyHGOl1TC4vH5RTIdWt4qqvyOBelAig50b6xO
hqcioplZgRMtCk/sJOP+UABJZJ11SgXOPRTdG87iKDyyO6rVCy3OiSFtiFR+gAKa
afZTwKPR3VN29ooXzdhfL+UHOgBMsTGU50yI2c4YIH1EtAf/oad52b97GHv2xVXp
SN73g/ZP134ZNABfBcwEd3JlklNJRfBFSUaGVENX2RaokD0zSn1tPGgtFVcgYD6g
AMr0tPoUsVfbkjIWidK4Q/t2iYTXjDcv2j7IWp92qTHMXdZkbgUg6kWycWLz7joj
nuM3kn25nUztktP7ZwTtm7nC2+Zkto01qKbceyF2lUx79C8Qgh1WiUtnCdpZR/8l
PNFsrxoRRo4SQnYaFA8WR7pBPx+Y81RLE86/5ytqYKJZA1zVa+xzJvwN0dvBDp84
djEDVGt3PjmJRye/Q1SD0u6UkbCaNo5+x6IG3lpBhrOxdGrr2Tv8TfNRmF1useWD
jPBcdQ4myI3W1J4tOsOhFkugFwh3cOlF7m3BDfJjhHDxeYuFMAsjJsxUx4HHaZG+
uaLhCG55ppM3/xzHkiVzNAsRdsoa4az/d0cjFlhsphB96ihEXj5GOtVc6kBMsFSM
rn6AhKgB6oorxVbd1EkNY7qdPf1oEpHlhsc4988rY1M95UneepNM4A8rCx6wM3Yg
rasUbqpniqXB7+ttIu/mGxRVxFdP8n2KP4jL7+9+Xkzygj3+TAOwErrDzByKwkPW
as4cKmWCL6Sp7x/FnT+32yT9+ZJx7kbCG4GY1lw5YDGfW0AQszwAhz0gje38jNfu
B/9Y6IkgvIINIiszsDtNY/ucdXaMKFKUAmop/Zey4qv0ftHtVAVV5ZyFwXP2Tf7z
2KqQWEy6FcgcR7I033WzW1b2I3Nms9BUKblr5ReY07ZovcI9NRTIdmiCwc0dK4a8
45mPUxvvrLqhKOp22B3XUIcKK6Ldz9ho99+0kWURIHK/dF69Mo02SXcIGAiIzZo/
iF9Z4Vjm0ETCHm2oIA2j2a9lMqCpUoDFIKyl51YJavFzMavqMsZXX5pfa/UwoJ+1
uHpf8Ye+llyJ20pusWQMqh0VGSIbM4gfEX1lziheoZeLyPa6Ji8/lt6rAaNDtoaA
WoAgeMKCq/Au+bg4mRDio2Bok6nlkw/VDQEw7gMRGAseb+fuEwSbNpswy5lv8/Zy
CtQUDjnaBbmee78RH9x8GvS3davHFlPZoafbJ110JiylAY+LGGephYDZ5r1jQoIe
4HR8SFCV43Az8YEMtfjVTHlsXkgBZxgplY7mqw+MyRNU0U4EXn12vj9bxwoVUx5t
yLe949t6oEZ4Y8pV/hbBBKNit3UlNYHSMSPGpm7q38gdWdJ4C7EelMnp8IvqG8aw
CpJCjMi5Mrfz6X4sj/fb7pp9J8uXlaQAkCIOIS9Kx8ttSpwfJ8Jk5xYZMV77I1c/
OlvB6U7VL4LfFQ5CBUtVDKG6+wM9Lwbg91EcHGmWPcHcQWSXClNZLeqe/wu/pYEJ
Ogx1SAtJrgss+b9YcnlE2SjJ+C1u4iol0aH8KGtXo234oR4AxY4r4I42ffvCktrH
pB6bO90iO0J1GEUjQHdkjuCRMdAd2UNzH+E45DyAPLJoGo9sPebYu8t5ez5gpaGJ
mfih4hh/MIGTpFSqZISNJa8vyp2dsRPxc51Dk4/mK3iMf5xzbYF/1lh1GHjAAXvN
wX9dSgX0DTNxrAJp3fSTakUo0YNdT5R7iKQaiMyN7PBnNTjwwS8NXhw2Ubq4KGZe
Z+kyFGcgzodpKjLfXcxktiw1u70MPzS/63Fpdg7+w6yRZveyyizp7prVUxZQd9Hh
oW8LGSLHZLFNRY4XMScKLBOvGVD/nmtFH70DZw+Q6hytAwir/f5U+BBnKJQhHGbO
40eZ6fafKHO9N4/xFNYR2ONm/LazQSX18VB8ABpZxpYoLmrdVYtlf7at6NGtaQEY
oQ7xFJSeAcZR7nXn92eQC2zDaB216ieBsBSQb1PmMJImHyqAhPBTIChJZJidw7Cu
YaJqAAUHNIRk17b8j00/7AiWZPStTqCNB92taWSZtJRQL+qCh5jpO3rjQaO/I5Sq
PBtUvkL+GflIrqMvJApc2e4235dafrq6/vFIX11uTna8XHgYOoVCKXKCQHYW1TMZ
LdvsoBR6QzOmp0EllLIbMATpATCt5QeCW6Om0NbocF7I9REWYQpNhKs0mNQgRUM2
IPf58O2ek8iqeDXo4Xlub4zjfFgbyPQuta+UOYdiSqY9+Xf++/rTIbv0lP7hgsXb
orAQ0M/Nefyle1GbhFAE7WdC4J+GlAvhyKyjMTnnZAJICeh3QsNqjJDX54NsecVu
V+laO46aNBSJukhnwwS2XF4StFmkmlRzkuZJKkhVpabOcWteiOxinZeaRUOgd3gF
8495bE4YN4E9kv95CbgjR8a88Wwvfqv4SvZVkfYmYtgTX+BXiIneph3fIgWChYaY
12ZGbbt3CeqmkFn+k0SxAvSJGcDzhwRWxbAttXdYgDjXz1+LrtvGe+8twNyiUgUe
MNj/YU7TeF8D9ZXz/RMnH5kAoSmsjfVnc8wSVWmGtORLkNdnfu0FqywgCiWkfpJe
wSeEUdCPFQSGg238zRZGkvr/yrXpBv1MBiOgNJsyGhmbdu3TPxQgMLbxoq5ixctJ
KbM2F/WaSjkza8FYKn2Ea9GYcEMQh3UfaOVBsZpsu8occNA++aoOxGAxscR0yKzq
DVg5icb/VgfgtbfTCUsivxs1IzPIyoJ37u1BFiNf3N+08xVLvBc63dtisnNhIHGk
OcPT0Qpaiv8K0Z8R16VnhSb30um5SUyr+FIrIMBkLXmGRKHN2SdZOunETXlpSPIg
JVzk2znVzLD9jlaqsfBKgtOqLN16H0Ttc+e7wFIlIRuXJeVFOzHF7kAQFEEprRlU
WkdWmuMkaUE4QWD8AMhyT5YZdxalpWeH9XLW54U9yc8hye33za6oIanBkPyplzpI
LFU6xhBRlyAB8mBI/81of75eo/6HWm9pvktvL7JRSg3k6vnvKnvkeAdNizOH/Swl
Km7UWPQpNALYwhXUW+4wqM1HHhyRRK/MG7u7kCHkW6I5XUk2PtNpgz8aCCQZ8RL6
Uhn3TqYnqiXQ+jNP1S27/uqnF8FxQHJbZt5c5nRzl4gjVDmmkxvAsQ4JDFsJ7Pin
HOUAO9omeT5ULoCo3HQcntXEcueLz/BUTNTj/1xiq6TQXWN1gmjM1dJsRJhtXdEu
OO0OkuwkAc1de6MoIjcTJhxmt2pL5RQfLCjUJeFJJJmL6nHwDJZ+PzKDV74zDOK8
mS6VrXP8Ymm/LRC+nnpB5IcnQCiJU/3UJ6zXtFVg3sYGPLZJWr5MjF3OnGvYynKh
5dZ8w5/8Ao7VnXzkiY52zHicRj3/F8jJ0alYfEYfPKvDWPdjcGhhT2QJOsIB6dRW
0nuTGsi2gG0cvjU/4aFno3C9S2/HqQGBiq8oyqc4T0OUYyydJWa2aMs67fFhyblN
HJJjOX8nfdTzv79UGv/xwqo/giS1T0iNrKW3jU1zXXoXRgFHkAm3lR9TVkL/ajRv
3zMkXas4+m/JxfFUgw1eb9PMVwxTsNDanxlS4YIrNmMCcJJRE23roMu4sd4k41NL
NrH3771XoC6cYcN1F65qaT3/J3BuxI/RmZJSgOrDTnDNjSp3RkmxXa27f1qPt/OG
yN6K7nIbaBWjCrXlHtmEaZ4fhvbiP34QZBKDYTRkwN5ARaXVUWPA/Ox0dFSJNKwu
LQWPRGJ9kQL/BpSbIEG3ydOu46nhrrkISmrHq9ixevGGzghpd8cAD0j6fLA3QauV
dGgjTZktl0l+8s5rQ3uih+3bg8FGm2PNvxNEGOo4pCQKq+hxgQ3ClTcaa56T+W3f
2D+XIvLI89Jt93LP3uBXRliwc4/oMMTbH+I1PiS8uGX4kgLowisFAoLrRVIziC/7
l3AhffHOet6Kq8jz/zA5HrZY7qI64P/2dcs5KbkNpX6SBc1owDSVyezWdt+b0hji
bj3Pj3fJNkGjelGN0Qx9gLAmVEKP054RHHQi+QlQAgOsOhF/fw0EdL0Ubb5V5BG0
/rMHuOHrmCMV2PudDo81I+KyGgsbC/hy8754BAbSUZeAcEy2otHag3Eii8aUOXRY
ZoRJgOA/2/JMPaTVMuS4qK1qFdHArcJiI1Slr+ultAk1w8xGwhzim5fGvbXPKkHS
n6fG7uBRlsZAmjq1VwDdF/18EC4RHUaR/W7Do2dBFPjXkpEorO9peey42auSUpRJ
c5HplLA9vOVh5JLu0s9rqBwfuYMyQNfbrcH8bhFCHIKSJZ7sC1xIUTnUCmA1ObCb
b14qbGEh1IAHmUusDcGwlzCWJVo9Zs7fWJovjET3r4ty4y8RvNpgwk/ArquHydK0
gNIFZ+Nq9CozNNkNUF908JpEnvkIv+UIFMrs6mHrsvI8T+o2MW52wqcFWSlsaYB0
i5YJLVZPg4GDSxTxWot2J6xRyHd0EAFaQPOw0dm+Yp3bkdSUhI3rQr5bkDzkg/sx
Sj8J0MmbHkowS48o12M1WCvno8cAN+r231gZL85n7maBJdlN0ykY056ibjUSMWOY
EJe5h/GifOMmgQOLa0b30oPwMD+i/hbrOikmemMJxH0iK0hF2+0d46WODsFjE/EL
/1vSyxNqwTYH6inKCjBaxdXN5P9wJu3iRPZ/o9k3ZqUyw69g9dR+XlHv4XaqymdQ
pN7onJkeRF9PkwPGW9lhiyTz72fqyCOB+O6SLVj4CzpBiBL3xCMDtk4p7tBzH2xd
vZx03mu0wzbrS1AaavRZgc1LeOntXjibjbDFRvLg0GWA7X7PYuU5OvdzCAEhQrft
/BH9Z1GjJMwHN4OOfKKXZGlSLEPeAkJ3opCojJZNR3RBfpWwcYUY7Xgb6I5PUsta
cfGz7pDUrVTkGQ4QA8g6P1EfAExqP6YxZRNKP1NQtpuv5dNtLzbVU43f90T6v8x9
OA3X+2eGKicC2ix+hyZMZAANxlXOSd0QzxjlV5rpdYnDdgSlV0oNMEJIat6kR+If
l3/n2IWdzXHHQwYbNdTdf9BIo5XsKI6vR5a84TemNu4YbErY9HRNyhX9cnc3d+9r
h1VqzQOzjGKbNDlfqXL2Yjal1bdLmsh2Hcz+L4DwcBbCHTB0aGpSeZVjeu7e9xt5
jAAoMM9TqHWMZcclXcgdf4nx/fxlAz072MlqtWHu3xMGqwWUUx3SJhZpsQ+W8X96
Sjq0m9AJVLJg5uA+aRE976N/CxlJSjS1bxBSnU0Ppdt5CEL5Y47buOHpgkxzw2CD
Qt3ztWKYYipRV8Gyp1hbCLjtdlUKJCtq/RJH8N4nVQQeJ29g3QFu1I2ZjpymJ5s/
wLpjRG6vp74gGM2wDvyVEJKZeO76vD++te3uR5cGUbDxOkZQoJt0UrEnzmv0/wd1
LIZQdtc/nbcahg6mgsKReG+VplKeWWjCnpK/at3ien8jN/YKFBuLCdfDbEMHJlyA
Uu4Btv+KD5P4oW0keYB8AAocP9bcuYBlQymTNQmD9lGE97gBpQTB2CKzqJ2ZDkFc
uuVoee4ymtcWZxCFh8vEyW+DJDFAS0M735CXOpxqYmnyxi1w+hpKxMCgeVtI30AS
OuMcmgZoswogcDGKoZyIa9oQA1bklDAuHrJR6b6uTMiX85p2uYaTtLsV0oXM55zm
ms5U91rn662QKVgzM7Mt8tyvLZEKU214ton1qx9RAMu6exXvg/BKOv1Fu9ITLv4H
RE63qvdcPoZvSP9Ww4f2lMoKFcgFPlaDt99/TKewXCmOgmRU6KnATVJuNm61RBiL
AfrwRQfB9U5da1qUGCK58GR60WOxo03NyV+g/Zzlv/WRwtznB7r4iP7fx+6g9S4C
6+cFRWzM0OimVaIhPPgMZ1UBl7M2O6Dv6I5Y9sNTSW5jdCCnJ+KaDo0KrBruivD6
0EsbAibBCwxv6z5YDmgV7bVVAbwe4PN7SRssgUeS1chz2A3SVwXuxP6JvjNgPMpb
tezKV9QPQL1VeRtTRYPsNPEMMEGs1bZa2ztlvl58Lp02Sn/TSUgduBcJ5Owx90Pi
fSQ0tuM7dJO0eeYv+n7D2dDGDHrkzJFEZctuGWAlb2haxT1QmaTrpZKRwuJYsnhA
4EPJ5XNgyTi1OCb82J4U057puoCkvZ1I7nPr+56KrfEPMhgfrrKerzA25PezRZd8
7dAinR8GyIGmvtllUGZOjAR5dKXok8E7YRbrDwDL62BWJ4xtSMjXI8apnDdeeip0
sewH0qboBU/i7PwaBRQzUw+XDJU8ufkJX8gXRm21/PaabxyAGgvMeB2UPaA7rUqF
XLP8qzgO7crGSAjZpwPYA64Vo4/v93pYkAxXEtdwutp6MboD6AjN/acE9OEz0p61
ACNnygAYMi4Z8SlL4LAhT4/t3XtqzaMsoCNCL5kU7NWLksOyjHj9SqSZDlgrBOGG
FxSNa4rOdBLVO18Ukx71AQxxyiWQuOjUg4sQGj3TUmqZgehQqRhnN2gFK9OqjE+e
l22243xG6ATRuCSla2Sh60+ktodAeG0P8xeR968qbXio+5ETJwIFqeeJaqRWpopU
pC8Dviqfx03xkU638i270/qTMWtGFcfAnWJFmq2t+4jt9NToD+ui86o0fAm2C/7h
Hx1AFE141+hg/rEyMCq/o+rjq3j+oxFlW7/vpQlDcHRINT5T4qTsUZMf6C6CrAjG
6PLnauvxoNtFbPjk8gE4jXUafDU1FOfKMsdZ85zGGeEOdWiOjfqC79q5jH6S5kpK
6qMr6sYFclXWOQsK3Kub6LUMtz0SrpMbctmsB/xF0zOMSKn5uqgKmnnKqi0LBEe1
uVwcZLHM4LFj61XCPxAYjuSoXwQAAa8GwhO7wtj0nsNYTbK1sOH55q+DvjNw2Odi
OzhnU1iPOZmtuwoZKLwFyaxUk2RMeCQ5tnq6ieC+E8+tog0A/pC8cgFmzgiNF+68
E/kCHuNtJ2cERHW5kEJGabgDIZzHENprZDY4Mw8zkJAV8ZlgrJDC9YER1IjZeXa4
c9EHZsF47p/rS2gKNtwReoqzn4oqctGNDXqBxKmKIHtWygyPvgyqkSVY65PWMfon
ESDgffqL+tNUzsgCUjJsXaUfVaxcva5GW+QpUSFds6K3zzK2ZF0hV8gkUjq8YggL
xc9/cJiMuDHuQtWSWcUTBfE2myuDDdrUJWzn5Ula4GtWB4LIOTFCBviPbOtUQC+k
xUO+upS4cFnQk+htPMjUVaRA95msdQ9nC1R2hAuy8wylRy9ADVibXA4qndkHtf8g
Ko5O0tafhx4Uxh/wgc5YfPKTVGZyTIRJAUiP1auGRaQTfLDH5s3+Wo7Gw1+SLPNU
ZPJZP5QZSJ4WGBoHVYjiTvHDVTsMA08xEfZSGPTcsL9fYVvkGPyc15nFxo/XaBkt
HEan9oZ1ju2DAxMqwV1XILXxLN7syLJiYa4WuApC+EKzvXoWZ2Ci0UCDKM7ytpvE
W/TYqoHWwvCRZeLz0Q6BE9lqeugOx1daa5oBSQM7oZIZvNVFTq73+y1sKFwq6/D6
tdmzpeMHr4blYyNGjoyh24GePqtTEI1zmVwBojIsdI9xXM3dAo3UKT7qgHE5X6JW
WO8iIdZHrqMoI8Z6O9kuwebCEH3Hyx7EeOPB0Ji4JHt/fcwDYaUF4YBXLzrJqQZa
tKkYwtwqsHrXc3XAlBBpRnHPJPCIkY4PJNLTebI0Hyc9rkDQcOUHbz6RH54Nhb9E
1lVVMLh716zZ1BXLHmPDc3VOkbmSPvEclU2+gQk9WCeGTyeZgzl4WOAl+5jbj7Ws
jnY9adCpBDsfhnamMgnfrtrH64jLx0aqnwK81L0UpT377w6wDEh+lP+4yIUC2jSO
a790INqtD2ubA0uaBwKVh1ULsM9CQ6DNg8YsO67OKqalOKmOV307IjrcTJFR9zno
zcJCMGGV2DgqAa3fios//vF4SRGOxlv2fK4UQynDontioNka5HJJpcwwh8fGrKVh
+jwkxrWtyp6zICh/q9bqHbKK+iCIBRxbRHqUDQVAMn5nUAgUfUUPtAwty3sSMvCE
C7iJDgFvNcKb8VGJlZBh72C6N2+a+7xx6gKrh5Bz9KlPQHMOWgh/02z7QZpY3B+Q
HZWu0aZgFGB08XPRDZDQaHyo94JAETG8JhRNrg0jj3KNItXnWBEnXQLdbAHRXObJ
5gBi/DdqcV4E9R4WUzOCv31JsfTtQMtP/A5y/Bk40o4I4BXSkeZqX0QYm6588K0s
8SK3KHyqC6K1PWe4ptlOP+oLUpNU1zZUQ6TUEjJ8UvRQNXz/tkfs2huY2iXZySLL
0wBQabKNGXcZjkEb/veeMptGjhF0WQKK2Erwfgyu4jEW/e0foSXcSPQBNzrhIceR
RUWMKbKMJnn8ty/+S+kM71ddc0ro+aROsw7moOM4sUdOvJlRl5eS0lVhGw87Atjg
ffwDkKlM5uXVCFDlBW4UToxZzjnHvPqBX3Us9IvEToPwGVmbBOgMXINhLmOV2c/i
mkB7KXZz9cjN9bnh09TOIhafxCO6Or07YL6WBdNrZS1FqaJqIKfVI9T/40zQ3yhK
QGihQO+UD53QUPlT5oVmglQCQPbHj+g2JALp/CcvimIlalhVe2vGijUgWWVyiKDl
2s0ht1ntdvcGS0Z6nCx89pma6jk6WdE0QYaaL/z/l3CmiO5ecvhiyoBXdLirDTOa
Ng5r9Zus0hDN5ARb7ij5sUyLQWKF5dj3KJacBPlwX3mUYkRAstLURCW4L++1V9N2
A/smaed5dmBwLByp8BHzLF/A8kfQy3eiKt+a6z7RVhk36CGTthiVoToOxj7rl4w9
ZMKhieQdv7MQXNnC6HAhHwSL7YpEEkpMH9uA0PU3r8WO//P/HOjnFeWl5+07lpUR
SwpaY6QdntK+bmh4DWMLxBmEQqnrmooAAZ+O70ZTpVLOMt4h4FKGl1YFzh9NjXXq
XtQVWSb1MJIx+tQUJ4cVB9Nggthf5NwTT056MOk05kxlv1oMJYTDbL9kLVCpXiqA
omC7acLXlBA8G2CCmiygRBIwsi3e9DHAtKkeIGuI7Vo9Ow36NSmrGwPpBtDQ3hmJ
xIU69Xakvc/QsFbGQn0PHIKQqwFXL8CFKW4/WQUfE8fDv8Rh6TN5BUCWi3KSzrdC
/VpR9H/2eyAV61TgTvROWmTgcEN8VAVfpDQrhm8aCbN/A6LOFw4+mid9gzHLwq5E
I0b5NnP1Kp0sEznI0xXNyMFpKZMyN76vt0QxtZqFUfPKymWu3krb/MA7kiQcpPu0
GkUGy7sUSSYftlZ1ptBn7+x2xW797Y6xE++ypbayuYKzcBAXzyEjAL5PS86yWmhC
VI/6Lthvpg74mZayKbXOXzZfhqU8SbWs6uhOzv+gOk8YICKr4UWF77BZl74y5pAQ
QrIRWZs7wfHlYdukhaU3gE1LpPkpXJ7UKofuOvxRRW92NpVifgEdtuGAVrpVGhnt
L1+DeQclIue5b6+NslAGH+ohD+orpyE4N1o02GRPcCpHgoFiMUGbbUHOEMabBtYG
9WhkMCfK3dRdf9oxCmSeYF629tb/RzNRPwqAZCOqxvJNAycJJZ4UmJAiSOb1WUtF
U7Vk8IHgWFhQfi/sMFMcj5DhNH9Owk65AjrXKvIHlr/4igVNkkHsz9Jx80MlMDuo
5S50O1hFuihaELu27fB3D2TNakOyHD9AdOuDf6iG3Kk3shcZ1T9+onEuoq1/Mvk8
BNXcmq37UOkm7f8J9M54B2Th0FcV2RH7UlznZx01XGwBlCKUPVJOz1iX9rqRM6pE
4IuxXk+2fh+8lhD9NnXh7wuK0UiCOnnGO+N5JKpUqQlbsHqvz51/OJr4SnS2LTKm
y8W9k5SGNeU7yeovud0CLrCvhA++ZZz2YqCQuskhAClk1RaG5sPoJXWf/zWbQlbX
smsgDnw/Vac4wv8pp4tfKGY/dRuJyUpQf1fI62KPbSZPagASj/T0qkmKjze3vS1d
ffi6WaO4pnhDuEH7rAEbgvnFyFXfAcbf3jilpCdj2Aw3Ilok4L3Wi+NObcP678/z
eS0WHY3nQZII69zfDrJjheOrKPJlcthowRxOrmnGgV3MRSt87/UtxW5/P4eCL4f4
7lLPAju5fHBMrarFUydyIU2iiG7TIwSsF2WibRdzpS+xOYAqUp35M/iKZJy7Hswq
YyikYM3M38zsr6d5lnSSV0iLbu8wZs3VxJDlvqcfogHnjH0WB4wivS+VExpN5/nc
Xw184omxzj9zK35P/MxGyxE/7O8lwTYLi2IurkmZrc2Sk3/cN7hLCgaqn4sKl3Gp
JWbYK7JBPbApfHmGqtDoaQHoti8iF1gjKklW0CpTe2mNBTQkf4ML4ZCUHUYcUz1F
Vj9IFR43yi2DU2GtuUTPcx1cq0p9+3G+5LRNmWHIlxrcMLbvjsgN2K9tUkeSi6eG
G+OuJqqnXV8wUMfYxrtYIMWcQoB65ztyZcSxF/qJAiHH8wtOZ+cLJfGu5OcxlIUE
ugUb61delrC1DaXTSPQ/71KQZCXqcZjlFFvdnQyMmwXUqMChQzlgjnI87RLURM5o
J9kPpbonLAHK+MV98HU36u7x3Z3J8ZPKV4x1dY/ngWeBVvPDm6iepZg8n/mA4GyG
BcF93EAyhDxXjflCBIau17Y1DvmFfRUf1fRjN1GT2WfoW+uHAB/nMX76rJ9jBsKQ
U6mVzMydfViPM76Icct6CBwd0Mr+jnrywVKu1ORjG6pRxNK3wGztKmafxlx8KLW4
aLk3TAf5a/Hofvo859N9wFgAq7LtgFdGY8F+BdgrJms9QY500fEFLlyIbZCKlM9D
S5hsDW5ssv78znDq/sLnG431S+PwQp5HCwXzbqUAFBeCLwqduGnqMq7petNetAlD
T5GO4PHvp+W7CpvQtWLYLvNi6p5D0ukQeJ1HzKADTbhrT0wVZUtnm6Iudl6n7CRt
PzYFuadiL8VlsPo3urOR/oPk39xQujb88as2pTqjc+OJZawPJuje8S8cf4k4Fv2u
1GOlEug4J4fXr79MYZ4td2UkX20LVlAD07I0s6q31mZaX5DnP+398DLmP0Y+ZFMb
ilDiP+gnNPurNe8ZrC5SI/gBo9Tv2s9QuKBl0rpGfFPl0eFopWNerbWDtTx/SgBf
TkL2XDJC6VL7Et+VArBYwGim0FO0rZ3gKU2zE+3G/HMFWjismFDA7pMSKDLWo4L6
eiILjRQD26MR9s+mwGxPcduDJwfIsFO+fZnKy2AkpP6a44F0mv34KpyakY2rbQKZ
nIyRzptXc8YUbr4EFw+KQFeSraQJgPFShbXDvU0N4GFBBiVs0dF8Z+h5nl//2jSY
rYf+veOFvDtNvBTPaTg/fo+rE31XcltZ84dFCe8zcax46j0KviGFhHpHzpT015dH
FBinJeGDU/bFgmvFjnx8bY77gg/qmk0jYi7k/mZVgBsELemPLhCSoVWuQqm8cZet
gQo5oPydmGFCkhO98paR7y9Hnzr/x4K+cEeL3CrxkEGsXfEK6+G29R/JFF0D+eVa
uB5Qhbqqd/3h6PqQZ90EZHvDv9aE5qjzeN6wt1oEbFhK5mHz6Gh8+F14WHss6/jk
DTG9dCERgFt6tbPLyHQFuQgb+zE3N5jSq/6Nb/mahd3izPXCK2bqKeVhD07updV8
NEPy/RpG453rlkT38MlP+U11Q9efuM+0kwDCAsHQNeqtQ4JCNUh6ohMw0+lUKV4q
6qhGz66diKw3pqJIvGmUNJi1QWdL6xWdGZyXDrH5Iq+HHrvVPIGO41GDcb4RDUPf
PhAzseKruIh7+nii/ZMeVEYj3qTi4x3p5un3PCAeILXkKkY7on0fXe9RrEOLEDlW
ddyfpgzzzUoNk28UY6nCRHljLkI0T+juzku2GNV0SrbtvJn6xCXUbYaODc2hoYSl
0u3SoXqxRMMt2yzfm+iFpu+Q0YApxwRntbXnL8aEaCiXDUgus7ILiBsLbmXR0wU2
d+BYfbqAMmkGKX1QXPkat2uA+Dwq3MrY0N1VSYy5OzyyMCHng0/nmt0X4NntbbTh
DGDVpA1ZSdC6XswO80ws/aWzeJey3Mh3c5KcToNJrLyDptZ4O/MK6melCteRwjfi
PS4qocbGddm5XuDwJCcKnWrD+aHAn4NddRDxRLigO7tBDEPPPz1GnDxaEeiTgFSV
wG7O3kIXIWvIXOgNWAfnY2a/Npwi7f3CWlsR2oSnZ7gOeRKZB2RSHK44LfYb8jvV
981dORUftZNdLP8w+0AzbrEWzmnyfPrR3U8zkk92J5rC+ve2anDW65v9uiit4V1N
/skQ4hNS4HmPguyYZXgwN6swB9jVRYXfjbfHQi51f4AoGYJ0Q7Uzoknv+0o4YgDr
QMt9AjghGc20w1EUoK9jVo6UOQltMb1RxKcjL6ciGNL+2ltTIGVo4UZT2dPp5uA5
l04mBgz8ExIpnW7rvhwJ8CB2unfucKZ8rHmt9IDI4nHIFUhGltgrfYv15vQtgaQ2
rjfQDJe63LdT90O164YqtRUwtr7tgK8MmHPGCwIHxmklW/BGbITJU2kGs5DLdDsz
V9GmtDm09GChunLkEU6zbcbBsQMggMapDnzkNAbzL9LjZuG9BbkBR3jzEUBUDNJc
hUPSplEC3PwyKfOc2nqquXjtZ4iknB3FhNUkIHCb0f27ohT5EaN7CuXAEfCjKOnf
JFjkIceTi8vl5ybEuwedQqXa9GVjam8G9gyam01E7vohoLG/i4NuHVYVEmfk/Fku
+QP2iqfnoshFAwvZO/oFdmTL/yXorLenKPntUFpth5fnak565roBKm1g3dlShwD1
qmVvgrxsxEzVs2s1/qKpwwQbEPrhpHc24TcWTEMPjVU5L0rgygaAQrPGjJP7qCjQ
w9w+z5Eyx3J+4qIfFqHtijR5DaqEfPelu679UDohdIGKpKMS7efMK2ajF2BKPYYF
fTQjTPfnaliNkKIJnV9Qk3ORk1XJxVvmrDbleU3EuG5ao2CBhq3GpffHQxsm7OW3
tqKrEC8GQ9cqGfeTuy4/dxXPo2ZUzgU5eNQP/ebHjfuJZNkxqtSDpcJU3wS99YSq
nJSlSJzVOi3FU3Z60JcrPfwelOWk0IzQnI5cYPyILAdKQpPgUf/XDk5o1DS7rMN3
JAs4Nwev5ZJYOMk3qA+15XBjZxB/uDaZuYRNVxWbubDo6umlNdLeBvsuutOr8530
4/WUQthZgO05gMfR8PWnKbnECzXdZDf/1yeui424VFaP6SVQ85e7ItaOxWncQtcw
3WQa6oKjviwD3AZxLiT/ABsxBJLtljOi+uRuJYYObPIh+nUC+jCd0S78zpk9Dr2s
7qysv7PxCPU0O4uJkbK06937XZ8WbEaRV5DLTvOiN44QJvbfwXIZlPU5bweq1WKu
dhwYZ3+fcqPUa6rEd6pj9mXZ04fbl5iOpXCgTwPfK4VU7lq25xEkdHO/C9BiQpnW
yUU4uxsxTN+SqyTuvYDm7sqekt7vAWSe3ivb0u/oEblvuL/nSQFokrogJepke9Eb
1ngNu6BhhcC4n3u2xi/a6KmE0FBYUOTuIAk+b8wpNorTVLAFmG/ME+wdeNldlWJg
auTjvJzMuNQdmA0CXuKGCja9sk/njBm+IG4a7FbDNzbAFYPQZcocqVZr9JSJ95YW
/dzoN+c0P3mkt7seioSXJZgHDwgdkunErFfsXfJv+5uxzvQWycnckzv/knauvCXn
ymXmtiINIuvQgMzk9IV4eZWJNtIB5/SRf3H2gRZAyfq+oaRfmQLPfYWrDkcymgkz
aJopNDDmQrdDczA1wQSAwhu0Z//4Q6SOUEBJN/EAMjB325Z1eWAwt9+AhGdX0c4Y
aXIJ+oFnoiEdcLMERQ1uyUur+2a3G339vnxqV1EDHPxYMaE3LLlXy7el7Ar6hxLN
C2gkl2uDJXYdA+JGIrGc+6WdYEK16plBP0YFbGtUR1VG9a+i1osDGVbzQbOzka+k
oyo2rPWO9F6mdt+EQx0+cZn/3WbAiFtFoDAuWqvQHOqTkVig9qmgGcriZsLyXJKM
YQsFttc3nIDHAjzcaVCdDFWTomg0JJ5AsDDucRlu8e5tuyw9ZuaCC/YspOHaFx6Z
kYwAMAGU33CvaFg9d1t873qrJJaeX7uZoR2KvPtF78U7iOmWBorCIRrrsCNIeEOv
x+9TDalXZmvkMxsZc//dBMqWLGIWFnCiixlbrJICRUGY+VsiKskfxVWux3c65yEe
SiXH4HPu4YESdRV3KoxGd3dvgX1jnGUuWJkJyBhP55zZPDxQGCH+UkydWVNjZCA/
X3g81LoocmSVwRqqFlG8GszHQCvpEGgI06WoRBpwFvOV3wL3p7RwW0VpLZarbDZ4
MEyCc8Ud/BxvlkU/p3nTtANfSU7IIUeqQPeRhzoCnkUOx6Zprd3q78ZztF4IRlkM
4bkq+4zc1AG6YXLZzpZ9hBRnsP0Qf94va3EIrZ3ZpKtwNZ3uD/DOke2NSnY6r+/g
cmyfh3XwWMawS/qXi9JZz0G6nSWWwekvNb4tQLq5VL5zIwmZ6Io0jQbNm8x3VuPZ
sgDLv9jR1SdbAVP6GHgh/R16YH99XkMMbI9dugREIm8Yew1p57dI657VDRHbhstv
WHnjYtq2tvnFzlvSub6ELhOpPgwqWyZBFYdJUcQXDyTgzAIjGfs0dVHfXLNKkgvI
koVGDkWcWdZnzfDbHvy305qOL/vl5bA1fxGihQ+YJorEdPODydCK0dncdOGNHk4u
PMgxa9sqlVWsuoQwin68WgYTVYrQpJfjQY3gyMmCt/f5XY8yBwNjQji7n8MZ0gLZ
uWlg4V3VEUvss206kLWbugh7e1NPvZUvw/HrLM/WdICwfAcd8eROx/zuN/r7JsZi
Qy8CYCZisIpWQR7BHIS8XAkWNhqgmXIR0Kc5umGkqrmgWlI6ZirB8bPfO3BIisjm
3yCBLahdQKjbxJigFDcSF/c9JyYAt/jASN8oAWHuSA4yaRevJtcuJIBon/Cxr6ZW
vfGI6pDakEM/zh9tzx6Wce9Cx8kHS9h+vWsysVZujYor0h6dsfMlZ1ROuP0lTUAK
1EPNz/UlCIpJbDRsIneDGgdiwIhbXXOGyRXAYMkm2CJGD6Doq63j8IbTnwCthtHi
/32VLJP5gUbr+ESjdBM908Wi+fodPmZAdW2TbnX/XQYolmOrx27GrSA1pAXpNtAs
GE3DSDR+mu68Nu66LU+CgbJs946F7P7pMa0FWuDjuPFcr/95UsjuqxB7QEhxf15o
AT30duVxkc6AiLZv/M6SzdK5MzwmSK/kWlRrjJJG77hwIlQFki2lPHFZxKPXxeCg
2NcZztivn4dFczgtvksbiUJEp9cfJYzenZJRCx6mIyDg/+4S7NBg6EjMpU2EH+UB
YVWvLatsJYRfyiIGrFtmeplQOdUgeNCyRRBbhSzb8CEFr+MQttdYU8tW9dLrW8NF
mAv9ll0YRSpjp7Ji6iPwMXCLPYtBTizNsQxcCshqwGxO1o4XEOPuPpv0hlcCN0A1
elTe2hLE+blL308tIuNJyk5mgzFS4Yqn9hNuq1hSDVFprrw58CLiZUVHgj5lIhYw
n0sPpz6Mh1vL7pHYPa9E/p1ujQ9fn1zglzKbCo7Ta4S4+YcVaKYYFd7B2jhXEi9C
iLQcr4JIX3/AHjx/yI2WP5VV7Wb4hZLdQbwbpnjbazgV6sPZONjetdULkIyh0y7Z
z+2IOXMoTpsurW48v8LeYyoqTGf6FcsABBzDpcDPGH2fbxtXZST7TzaQXeIsHVnk
vESMF6ZBiJLq5XZ4uN4borseYI9CsANtyeFzibxUJuNxz36t9yNObE/vVfLzUqA1
/Bz9oSDHgGfI8gcHDlM+RtKTtRMUrzO/Cg3iNyHW/bNsxLnN9BHNwGaAsE1z38RE
X7r2MbCINA4+ZQEDvbMNUd/L9GioVgRTOVYH3mvDALd+4zvb07JMJJnLHD+RWIXH
cfzcwZTjpBC4s6f9ayuYkIAtZW/bS47HL4o2f4S1YjYubny+REZOnEGsfKWXSDM2
p4hEZnwD+a9pfcZ/cQGPhk/1ZYPChJ9rfCOiCLvjz10ZoVr92Eypir6DRt11pjWS
rbYbkeesApzrLPdYYEVcGTxLCmY7ieQYVClxMirAKhMsX5KaWzgJRpdZTwGWAcNN
nEqaq0hC+SfWZG/B+MQe1quhiKcuN84s8YIoOqHh+P9i8fAQVuIyEsmp87rMvRu4
GuvIFoV4w5A92M9PFqilS6KziU270uEi7hT03XGe89OfsA7ZpQDmFhkV/giXrXx5
KD/ycVQBec7yVZoS3EXAFj23G7wMi4Mp8g4WkEKBjlp/NE82e6M+3hKdHMWv6w1I
f4zbkjq1ePlhhzdWOU1IEY3GFF33SNKoS3qmb3QMocpcgHpQrC4rnDkk0V2AoBjp
HxIn3ZGqSQ7Opnt2f3D1YldcNmxH9Lr6jX9fJ6qzvtC7Pee4a7TsBTxMmBWpfWww
6PYBbSOr7S8KGyIfXAaG1svvCknOdbf18e0mPhMys9c03DGdLbM4PkiP+G0JSo6V
zlI66aZXn8PB1QQ6EyUZX1Fkz3ZnkQymgeW9rMBTaJzshoaQStLHXYLFTitCWMh7
wB0kM9Grz5Mggc6TiIPSW1zTMALfUGBpoQWPtiHNHHlfnqjrZrGV37/dWzpxwqEg
Yfw9YDDN6rDn3/BIoZcJbfwVA+gFcD+9oRhr40j2ljy4ulUB1NltfZ9MqCykDYB4
u6BdgrBxwow5i0devQXz5s7kA/JJY1pcR9StPEAO9lj74Zumf4OrE5QasEOYgXar
ffRM1swuZ1IOwqZXw0BPEGoI9VzQsiCElwEsw8AxoWa+SGy61SkcMGeMoXzi7UTL
NnDXkK1tYFrIWQsUrPIPhsRHsqPskoq3uwm/c7vGcHzOPHj6m9AO7ktjJWFNrfAV
e0dHatZUxbpAc3PkM2msDpGlQC/sD06TgfJUR62juQH/ESsUHFm5OQueBuZYSnJ2
OgI6GysqwnBgqwSMhjbMkeRL7e0pyieibsabnnEBUeWI31YDBHxuXj9WMwavh0mB
1yg8dwtLC9/kBNUCLr2ISIKD4oy+nTPeZPJwGR2BITbkDm10VWB7G7lgLXSWW993
KIV/qGGUkuSADWU16IeZcbXepygo2z9X15MsxPdg+FgT9WfapziFRNNNcRRGoONZ
wUFHQL8vx68e0H9Y9DzTyVnCjuiEthRpj0XGm7lopkuLS1KXmkRgKTT0PRdOF96m
1+RtPo2p1TqFVoGVbw40ln60dQBZe9mnOJCfrjhvFkPz0mRMqwyctbKME8jviwnB
og2dn3G/9SVQEXUZDSd25mISoj3QD8vLMoccguwRk1N0HsnUxAa8XaGDVgOqp9xL
kq1n/GixZ1D1EcS/Gy8QGAsdDt+E4GEn7xtwXk2Xj3jDYqdph2b7xSIl5O6kG2kz
mIhY/umdpmsTUf1ZNam+U2BCVv12d+YPG9/ZNwJZir056VhFywmetqyjjx51KdaG
Vdfqde5R6Kt41OlPKWo7nArN5ofJ3rysUtnNyotIZli8XFJgZ+eamnGAZaJv57il
EBHsWu/jVwvCyZv3veGrXRivWiB42ab3BZOgA2nLgQt4iORK+MfKGChGVHoJX1eR
J29yz00iimK2Ft2jVWIdCHiO4XQEUNwrSmcHw1h2P8eOMA3sb2A7l+KM5bntqAE9
PwkRtnJ8ucAyMXVtpls/mEJ/H/m5HIJnO6FPNLDpv4Wvp6hVocjeIZLkR+OzmuFr
HwZRCzE2TngIVrZx9ZIDrki0ZQPRDzeL3YpDmg08W1S5AJVm4Vi2a20X25QnyLau
T7v2/Afrq6683hOSK/y2R25kMyLcFN+g8eTdrAg/Yt042WKWO8xiDwMRB9fi3qdi
2CFC+fXszni8j63wAkQAGka3Ug6pEB1UzZhYrHyA4oOggQ++iLTarzRMoWAMbVd3
jzLj/OynnTAf7/2aGXW9yz3frVN2Ap8FJOwG6Pq/9CsnDhrDtZNxc08RuSfK6hLT
GNjNsgRXO4tl7pcG5iNvM95tMvFaDtbBOmd4J9UnUEFSn4h0y5tuRsOdlNCs5+K5
TMPTIiv0cUl223JV/6qwIk3MOEBk6OvXO2DHSVeTDbN45bpvnEqCNgeNmv209Z6q
C3DKN1R5RRg0LMLvQor6fRpTklXBeAmIEu1xzBVW2omEFSSNwLZxcpFlUtNazBNZ
tyyryja/6TACEMR2JH6nfsAtzXXPbi3rwpFqVAZSvA41O++QDzoLQddFDZ+tIgg/
KI9qMENU4CpHSpcsiTFcc38+mNLaOMha4BA2hKI2NATuOmsek4xFgJVEGhI6UKld
5Y89p7OH7SZs3a+A1zGeAEOV3uY9TUHWjR7B43QNpue0HJ1+z+1I5rPKi26b4mmh
FB9bVpOMtSgdMEkZrJVWHHvZqTGjHiQedAQdy44/xG6irPiojKqAVe7Ug6SxkEGH
mu8Gpi5AxuBUR06JPwwZoJabO9dVxBv42E0QnQQKtFJLOwyd4WBw/JYFhJ9N75V0
Pa8h9MPXirxUoedI/hcPwxuCoTDlY5pBHhRpdUiCdz35q7h+8CO1K/WQnrI2mhtE
4D1gzTnv6Lsa2aJ7VAs0JU8J/bzlu+zcaKz8iNbiWxp+4fSuxBjPo8O5zE8NIVca
TjRSxtKt9hA6sDFwgwQqEu9Y1qLIOHhxU8J+YBruazkzCv+aOD45bM2yAtBHHIoU
ooRPkVqcxHeDJeikMaBg+ANpflEj2FnRhw7alcEpoXnznbSqMcFiiFo7eFtho1WQ
Xz36gkDTEwMd3G55WaWGYBRoPJB9z8IBOxoZJregGKJYtBX5i/79hl/6bFInSsuz
iaQ87pz6me1fEZmZ9SoDN+nWbCyHjUEo5XyniLFzVLQ1fcgXHZjCyjB4uHN8Q1bU
2n5vWOWVc8LuQUK6g0ify4mhhEottbV8I6yewh2p8zeSWsrqqgOMaAUtiohVHpTp
iJW3pTH6AgLPZxeJSS+2aoUbuVSkBElRrfa+pMQ9l/kpviFQGJ/lxcOx0hg51OFH
MCgAVRW11+3IpFX3olRW8POltw3IxXfYqW+K4QVinKBcHciedd+14AqieuZLOgV0
orzqU7NuE7mxSQpRhbK0n3rbkOZkvVpywWOVadAwB1h52nGLNIn74VszcqvEBmQn
fduBURt1WtCOUYjZ+HYFzskVbQecQUte6kFFg+ovV7m49OTQ5Q69TgWM9c4HCIe0
Bx5sZScQYH9IQdLT8z60wGR+lo+h90bz83rFUshNNXUgFgDeM4tfvFWSMQnWpYJG
vyIDcTvzb+KY8vC8RGTo8pDg/X49Ip5fRz6CwK84M0GkHag4QXDXiZWmRXkCpnoy
0+N1IcumCDae9m8n6e87fNf4OIzWsrJPUcqEolMgKpDHijJPPGpemzC0nGwIbYG7
kQfoXwrB0zjBVjunAlhmuwwnvljlJR2VSgNspfIAtgyTiEOp5pNuXeFFUEzBLY8o
yruNCGH+dQesZfhNcxYK88e8ke8bsbkeVa2V4ZOpXLrmFUzY0o9U8kZQxvN9xdDW
EnAvSudUzTIaIIZYmhvzMvf2lFdxGopN2tIORefpfoBfp9mdYu7HwI0nqk5tIaU4
fC2pGwnFKegXj5lhgeK9rcSuhHg/+yxW1wV5n5eWSTqBaSxT3J3oYYx1R/QaDn02
lePNFVOd6T3VG0B4uqHopNxW+LobL/2kGoTX1haa1V9GCQ8tBjenZz0bmV376svj
ONdO1eFCl0n3X+ZY9lWDP648kpz0qUYzQZ1PZVTJEPsc/URy8zrg/16jNoqoxdBT
YRPQGisLLH9iq1Lw0tBKKNwIYwIw7kFfEuIfa4RkY5J+urpD70aqDmhYsgAk132j
EWr4YooRXC48XqywxvNgIiPxKb3fG1KzZXBugsZbRnzEnyxT43kbIenGjIvsX4JO
Qa4P37pVz6/H8E691uN6SKLoPoqAriAt6PJY+CoPvj5tEhUtQfnwqPsdg/rfbYVO
Nd0tmR8W4+XnMTdIpJURlkBPqXHwIZ8kQqQ23umIihKBoHiDpdHv9EI6RhLPyf6a
IH2xgYenpoQlqLJE0LuA0ZA38sPVs3ZAUpE4PXZgKBihz75yLJe5BRNZpq5gzD8q
Xes/asfTJmpUDYntFlpSLWsRvkQlsAx4DTcIrc0cD6wnHItuIWoW37/oQHJVloiB
KY/FU4cxiJQ5wsqqB0g3pwG2Iv8yGFrQmhDuqXdmtakSdHfwT/9BYAfcHKIOjuMY
kcAAbnGlo2xVWYCk68LB7L007gupR3YivUSw30HSbQULvmln78jV5LAtoHMpVPAI
tgx13tPQ2m4w+cDlQs8Ktts91T9s6pSuwXW28RZAfBb4WdDZYl5hn1VoIugk8/ZO
OQ6P/PKO4HwFS9CKbHlYYXYayUpmeQuQC1vORJoIzDxg0uvIob+c1vPiM14OLpqY
skOd4PCV/iUGpu15vQPlzm4Z/ApYfqLUokvVa3Nm6oeI8C63rCViTKx3Z/oOHwO1
R/Ixx8HpXoiOz6Of3SlruQRCotBANH1GpaIdOBXauVG04x7vNPuqm/HFXkGrcmMY
Lu+qFaiy3/4DGkB2R23hdAlY7vC/oViwfdQ2nG3w0JcKIBgowk8hfhBbI3x9wGxN
lWbBEj458U7VoyWX4xJVhScRXfqqA4EAAGXKR+mW1aMpGHeFC+cxYULhzI0oc1kR
NQhD3m76DeS+sa9XANcpPXAA9m3kxBZXP5UcEPZKGaXTHbFbUc9PAPx6K/5OqWzo
FWsbJuxYISj16ivjzuOg/q+eMpo03WNJ+1rc+i/OXseZo6QVo8XrZr8ZCm3EJM5n
ixKBNPpQ+Rx4CxJgw4WVxOapxT/IKvMTCJHL6zJ5u/+DqeWlxse/1h6jtxOr8lvt
epTm5a9HAjUf36GFCRYqpnGnrBHq6uRbFtxeS4gjcZRoxe1bTrWPWguJ17xzegNu
qzIlLIK7CUzSBHwBc3xvgH/epAEWj/oauBFLApLqH3x1YWEueo0rlw2ItJFhSD+F
Tyw5yxz20fsdXxoAB/n9JK5lIv2JaIss7oUJWuZ3Rkr60Ror3JhRm+6OWBxPgM7O
wGsuBC2uGzwsf1lE7hsADA44oUnqAm2rnh0Tl/TSTEHtobZm8tQEeXyN591bO9NO
Cj8e8yrYTBte4xsBi4Qhv0MoInP3UDbAdit99ILoXSHTpIGwBUs9E6Jbw905fHwe
PKCruLg8AmvncydHGFYPejzJu8CU6cPY0F9HZzDa6z0Ubvg9j08hqgjJwqwgLryl
fNCdCQA0HqzzFs6YBtvvLvjsQaB3yqlLQfwVMvnFmFcLPlfkPirkDoCiYErsquRh
oYjIwqWvmi96uts4b25P+aK/87iqq60SiL3ZeY0KG9gncVB5yCIQAPGgy6bdfA6G
7ynmWSY9e+fVrRtmJ3xTRAduWsmuXwlNLvOrAjTFgIlBUbU2r2z7LFjjsajycS8h
x3ueeMC9rvWmK7ytsAkhpjVrPqwQZzKIuvSAAfdyuvb4v3lQdYl+BY+TU+vXUGFS
DafpsUVtjfRpUmAxAkd4NOP25S0Q+KXE08AIzPyza7gnOrgeBmR+PZ0yvRdI4tEX
eKl5zFIjD6PrvdP6pnL4mQcD4GdBL61bNc/f2j7wOeRlapQkr4zve7CZcQ63SJ4/
lPxxrFyoGX3BwzsTPfq+jUjsCQcjVJFzuhMkqmboj+pKxbvSEhWPFX/x7tezAvx0
es+FSRU2wBSqD9J+wtERcQaPQmTwhLVQW4vJkitXxdLzV6Ai5WansINyLrmnLRXz
l+T9O8BkmEptt4hOlxc2Az66XEu+5ijqHn6HwGRjhDt/iMebq72t2MiN1Kh/MAS9
MYnVsg+Z+bmNwQXkSXXYTn6BSn6qm0MCUtuvNTUTnQhwAwQxM/ym/5+BurVYbRsu
zXvx/n+AzOS//rTbYQnORx9bEnI/D4N6fuo+ipLqaYTKIutT4MLSaMUUGT1V0aPC
6GqhflOS5GOzsTYhzEh2LgNl9l6FigcPvNZOyNYP+jwJzlvul9wqH/gpCIPftXxT
buWpmu8t4aQmivRGmac8LfWQWhqkU4FCY9UFQJ3ax3R3DINjYJSuL49YPYosDSyi
H5uU8gy1dsNkW9VnwkKrJAz+PCmQIy+PbOlmn6dgNYm2MeYEFWIdMraDNB/R+D1G
I/ZyYUJj/05tCS/wCz6nLQG7hfu6sJYJSi5TeU6eNPPuI4QUrZ/Xmh45fAROKvTZ
m0e0tvNkrJ09E/sPMxck9nlqxN8DPf4b7gsZ8j17vhH6ydRx5uICik78P10sTed7
2EdqdTfs8KuBp9UXr7nYR6WWvge3SN3KlVMsI4D1NB+HNl/wDHGicV7bCMNwfDrk
bu0Zr16+rkchbTgxI/o5xS9Xiky8+QnBBzvZ2Mi7HaiA8fycxbVEO8Od3PC8UJyd
zHe0yVFaqsEJv1i5L/arXnUJh4CyJhvZS3mhDl2Szoy/fO08dfq9mjyx4wZnwLnZ
tWmqpTDRSXFldDwv2pIm4J81HCO/JPHdJ2IEOD7IWN7H5v3iXXekPMKS1LdAkggg
lgOGvwrmlEPNSNDZHHQ2tiTf+yaXYBGdiUok8/tuRCVzLWlTkrA/JWfKQOhHym3j
SnysJMBZ33EspeVic1uCets5jFPh2qTHzeITOInrmYEXjpTOg2KKfYmMPPyenYy2
4Mj0FzkVM+1uvvc/GvUeXfZLF+mkrwXWLJUY5s2xBO/u+BJscbsyU5VPQpP9A+QZ
8Z0UaltPS2x6t9QNAWjtEQ9eZ0kV6SKY2aOewtO7+AFLvKCROvgR90bjBKVCWa/X
CUL6+KA9NzcnuJAX8Gzx4oDb3gtGWOxAuoQIiUVELUM2FgqyyFaD7ChLFRi97QIR
oFFCPJoufgBvAxiM2GwZEvy/0613SBGzwBTaOcrfOAJMeh/L734D66tGGCHITo5F
+2MPvSf9E7S+IhJdsi78JyFey9/VYsBTGuJxynAgeqtGUpF81yzjmXfiFrx1y1oU
/lm9DFxePOo+vrzltqH4JiQvjcOfMdM4s9rOtjjwANhR5qBRZs1zQsp6DuAu91vz
L1+fQT3Yb7f4o8B1wVXs3ao9vowPIproQ1UlHNVclkZ4ZGa8hjNFCjfkYEV1GMvO
VdIhZM1Nsud93+H5vhlO8L9wp386yarqKXuZmkDx76zRBAHmeuVvwB2Tl+4pCIuF
54FezkRacCaRT2bRtR0Mf+DeDiz1fQwDUP7bdl1ZOY4mGKwQtE/SPrk5npuldw/d
Ti5K1jIiOFEi2KBKYMz2lNubg0QiElsiqutokWQtRH9C4a+ORUV17t2pZICCkwYR
Fh1CMnzegOKr9tZRsgzE0gy0Alihhjh5X/JxrTX9MVt46w/6pJs+L8R5sjeDsKmf
P+kNEl2Ft18atRwUBaMLzZIuZWu1qiMalh5mB9YGnqMGDQ93GSrA9A8073ijg+GL
TCOkxLRY2FrjdvRroVlc0QNNiC4OU0agA5msEkm021nYlTmMm6jlIsycPCK6kzjh
eQ7ZFU6XOTgaoebaSeAvX5QjiVIIhl/HPCcGacbp1x21TQGCnaWCSPcON9MxJrLx
qNkTx3PPW91lgtaOo2Q74wLsK/VZH6+CwXERHnFqx/iE3kUeC+Yatw28L7G/RwzI
XE9BoqROA16FGNVgw+BvLNQYticPd+wmpnYGky2IpUGIuClGN66A8Y2VeLwXQ3Bm
JUYu34Fskv65BSndCMfx/1xKPD4ZG8xhAoZX26Xx9hkC0nUqGnoDSiqvenVyAaRm
4pyXPxL5yJ/tTb9uyv57AO/OXAHQu4JFTVXUwqgRx21cm6WrQh1U+4Oa2tiPaYBt
g7+sG8sGDbkgahsefSFne5grxpsCv8IXbyQslHzC67+cIAjmJpVuZV+2pvtVocCG
2XXzu0iP7rs0kGLKtThuGepbm9VEgMtX4pqfTGbrDw7gfNUUZq3pjw6HEwdhGP0e
3MHcxTjIqO3fEdORNYXYuW6eCO4aMPWdwbMUBaAsrOrFca5D1XJjFDfJnnz+QJuv
E1W6T5EL4FK7RWgdGXJTgCsvFIo7BvXe5AviavO/W+6EPEylkemeq3W4SxXszluw
3SbTy/rebsNygkA+57tQNTzXVdLa99Z1g/rEHdz5vNX+gwwVb9wfZSDijW7gXRbl
rJNDD6YlsId5ft6bGbsNAwL565BPbaFYq06/9J5QK3caBxRCRUcwLN9UfqIZvtth
TenErxbaRtu5/sBH4Qvj7Atz7vyYLL+uns6U8ZrlKv8qfi+8inb0wfIWUUu14DA2
SBOXkbEFxWU4ZVHc3+m2Ti9bYWXZF5G0tcU4D6v++OqD6m1/aNEl+TOeJkweh6rg
AQ8DbbM3tFKSoUlcvpzhy0TBfB2djwQdAPyKs442Cv/J9H2StrEL4q04LBvwh81l
4wa/r99hb2xAUBZ0rXP1rRaD5vMyVfOhOHJ2Jrj8JIP0WUIkB00xIchdOG9pG3Ez
6k1r7rHdMt9CrAEFVP712PxJoN+5cBhHStDb32ZXkWrewHJa+zhKZVm3MRRiaj3V
F0vcA4wWmDd9xLCDLxWYuOXfV4/BupeZTq9CUA91q1jtyheJ5zvrThre/nuqseF8
H9cFAJxi2dm3P17ear4Ic6BdhHpxmE8YXrF4CmRJPY/dEBcYVARAYKRzKYqq8hSN
ql6INqaLr0W173I0gjbpzb3+S9DU1R0kJPXsxEfH7UZr+9bPTULvf2hCp0vM19Kl
XAIfC7fqlDSY2N0IS9FzUiJC0k9u3E4IiWBeeQMMkRIHMt5r0siqTNcoKFGU/MOs
LdoB6X/SYlFc8ev/Ab6n0O/z/MhX58LTlfm6BEdMZ/upZz0ZxnGBwe5C8U696H1j
lGXjoeExgGQyEE4MbTDfSvLL9mBY4bQ1eDuUSsN99Mugy1nwtAnMlK+yn2/FzpGV
6EvYrKvzn1wPXSK+mvoyivTbGV60xDxiu/SjzDzg8ZZhoDM0MRscz7COFiro7zbz
eIz2owcp0ii4rz94fGFgSiQ1IbhrO5cbPlPbOB3U0qccnoOC92gRl9MBsqAlurI9
wxok/ZZ3HSMADBmR2hJjY6rXLBv5Crkx2aus/PVHCif0nImdtOpRoC1k+8Yzrt+E
yM+XiLLjdf6JtnQkO0VbYznbmENZOrEYdtb6qXSfxxlYQBYkJfBG5vvke64n3ttT
+LsI0VFqbaiKRPm0ciXcgL/nNnoEcLB/sr3WxeYKSKa7rKNswmLHnpA6ojgWK/Ej
JmMdKaq71FltaHhvf0uKZndulcRKDYF0ypCQOvUQuG4zv+SS/4gbY83kbYdinj8F
Kx6ydDFrSSoz0BRS1Mx0a/MCa8xkA7zWlcWvcnX7JvcGzP8//iuuywSqH5YqMyy5
vawXwvdau9/2/waCWTrfybX3tyZgLZ/dkj3xCzedef6MRuefP4HOsFxWJxoz0SqD
0TSpxLVndqzX8I5oqTdfZiPHdUtwI10TNFtZBE/wCPm6VuxNb/6BwV4WJedGUSsS
Ctmn/gN6t+dwEJry+pu8l6reTNG2toNF3jF89DJAf0oUZvQtUp8IU2T9wZBalKuH
bBgWfABk9KArlGxzcqzbQtyiwvKz0nD7uWsoZyuDu/7Ns4PMz3oD87ygaggboqtu
jtiwCtZP8rxxTPIOMOkCf1cW9BFuh1imVFo5vX+Cnj12Jc4iohRN/96vc331FE2s
/KmmVja1geRa+/R0Cq2iLm0u7JQqEeYoj7mtzrcKsz/KeveI62zeFAGwmfY/Ch7w
q4xzZjMPPlvbjjUPZdkB+J/YOqLt6EOjBowi7Xe1BlQyIPVeefojvC2oTFKEz/r2
2nKecVTclPaGrDY6ZckVLLKZJBhJ21ltiA9A4bvG7RXt69+8/+czxxCUeomhVvNR
HhiNaW/eO1he6uPC1T/1hCu/iwGmZ6OtHFIhQhyIZlA1kdYoB5lWdY0Q94f5oWrF
ijTzkj2WJ/Pq1ZKYbMsj+YAxcbpxVGdCvQ0gdawWmvFF/Fbi1aUQAOLBpM6COzlh
K0NAXCRpUyDWjHtxISaHXA6OXChRW9PW0tBsT1b9w8EHmALLkiW7AYP85PiKQtIk
j/6tS/9tt3lbI2kLv/p3cHSiUIsEUG052dHGjQAreZlNeNwsOoV5lWbGu4fxQypD
LWOrCJXmZDO+hK2VFO4Yd096wMWT2v5TdBPyqmG3x3aQCm7zEg1y18mFbnzebexr
hkcgWy4qQZuXvb5TsvcG1Y0AnLXUivYmoh+twFEms/ONpmXyh8q+7d+ZZkFHYSFN
sS6NsbJTzRCHCRBWrYE7l+IMWtmX9yYQAWIhho1AuHqAcWlEuw0LWA+o90dcQ/F2
p1Zx/Xb6CRjDl+MEe5Y5sVYmFay7UieuYN45rTW00KzRCtGsIuv9Lc/Am61J8ZUT
SPuRyI5JsfMwWDstvKblTez4YGdm1p+H+NsAik1Fa72d2sxJ8ezP3CaTAYG908i2
QDUZ0/r/Zjwk6PqtoiVcDxSKor60ssr9kbs1iw0RjmPWWf4IrxzLHuiYeli0UC9n
x0ZUdF6E17uFg5rDg8ELhUE5vHr8cXSd6pWuB2G64h+OxDHFu5Vsl/WZZSPJGSgO
B7GqPkzAumRchQ8Dz0WyqgNutydQ5JuG+aVDxOr/pXEwTKjBp2o/qlnDb3Q62iB1
h8g3KyWPh0hubSV/beH5g0xNyqWJfgzsVchAT1SxwRJl/b3ZND1I8kjJ9NbP5cFh
4yUaL0+oYv/anZxept+t95CtjVdxfQmWq6GXbuBjNBo67hrybilTofELorrVFUjb
7Qj2+ocQ/ade8UygRcdWe6cC7SVzVfFlCAteH1XrfO1GXkaNEXTp4Zn4Ykpvwlvj
Dhg2w3SdBn98Y77UPMjyRUYzIgjuxAQ8I7i9IzdQs+IS+RSipj+Gb7Z25sPaFVfc
fAV0IBgL7sHfhqK5MBRtSTrMzziJ9ToQRmrcoOYXNNINNnDdT5Dyfsmo9PqzvctC
iS9Ku5AoZrOnzF6XlUlz7X5ktmhX2gcpMXkE+F/5RPHS7NIB3Qfjh49MAVsuiLyO
XYEEJyh61DLejb+rG0tr20oJUi2kNTHbJ/i7ACtJVXYjbimK2dRnXou8cV1TBq4a
AJ0FJvpi5AwRz1v737nc60M2KldEG90NQYRZqfwRdrz8Eooifx97V6LTo5mA3PBD
HEENo+5lnH+rbu3gkJnUJaWIBFWHs/C0WD/Q7UbvpKsURuB5fB1xTfE+4CAXCota
AJOGcH79e4WX7Jq0nYauuoDiQnCrvHVVz8rWuTmqGvOLi99qZCZ2GlPvpft5Etyo
OocNdcVuzL5/IzpmXwlehYRSpAHr7OxlgRbQWbX8XT3d/adLahU+IKWBwTxElELj
sY21GpiCZdJF7CsOy0oiNHVN0+EPi/+8PQuSka4muLww7d8gkeVEwCNH/nCjlRl7
u9d64eXeAaCAnDRb8dDkEIHVhFmc0OO7HXafmkqCx0XJlRpox/6toMCHxPjWlWPi
id6wiU2XyPYcZZsAup4VgpiNW5YY7cJ0g031xUhXXwvAqQG+8msLF67oNaQUGKk+
mqD9lajnNlfLnMzO7vlp6Y73fokLBFTort4aFx4A0WFasIPfgku3t1moNAmLN38I
E+uRbbS/Fni1yw2gpxwGyJi9raWUeF1c4BBpeS4uFGAfjCwS+aYKA2vMrx6UAsk6
Q2WlllQEEfrYJxm/Xu3ASxa1B4znqq13lxAUZqBaJALVTQT2q9Y+fbyDcz1d+7az
muDIKhTC4eWs+Wm7J9tQOaqZwldugnbnTnljfoYb1Czo+K+acnij6IB1kJJ7yuFq
hyNCyAec2nIuBKeUnRT6DYa55A9qcdi+q4fe/EXg5r8jbu6fA6nQtg+iAPGh4OYB
hCAN9iNcAK4FxdwSwAYiMmg/AG2GxqOevUvX72gf4q4ngPkUAvIhc+4B2vSLaZSY
VwlalyjrfatH3DG9vKdKZqbf/Nu9MR/ON20DNuddTz2tp+We03Me8HBfLJrwumyM
1yZRzu7zuHI5DMPjObN7YwTSxyvkMD35CNDhyjihjjH6wCBBgqcwrNZ2T6XUMehj
NNl3THtPczaInYS4VNb1sWQRrGyGGb1DfATNl0pXsRmnuQUaQj/JNxpbdfcMoAkx
c+yJNeyi5WIE/aBYhqamzHlorPOTXdXn+xve1chT0VZAWYrrdlQ9BNVfwAPIBYzR
VDhbWLno3fQl4kM8g9cdWwcTGMYijKC00mDTQojHRBGMOiYiJIzvc1y98BUKDRdD
skw/zWGH25CU5mnWuk/zOr+NvpWK6CN/AweO60f9shTQhjBBPpWWAHlo11agkenH
q2dt9f+IRs2cNLlfvJ8MoLbEw7Z3E66gtphz/p0c1Dk1sfDfEyJYAcHt8olydd0L
hQJwBxzaeB+DSXwr6jHAeb6hbpDilMZ6rWSRRoWAp5pim/ipcbf/6xw0ONXrrKXC
3tP2/zaDarqI5pL+BWyiOe1fwKgkL2ZyJFWCWnef/r2TfhsOrIEA9m9D5wfYjfxg
I+KQ0y+8fqwqax4jrH7F1mpmudjAByuC/9/VFGlMuBlROLTMlT1O8mpBjrOZLscC
/j+d7FwFolaSwYioFNOqfbCVqpFSvtjc1UXxmUDBDYLJv1LHFfm78dA+VbbnxyND
P8kjfHmvC6YHuEybTRDelH/rHnP7nXwjZMYLWl6XJE7p4VHHzwf3ov7TXlUplOpt
tARw6iyMqpIdqMmL3HafJYdc26wGBMGlSniwaEUiNis5ygg49gakmf3nT4UxREuF
GcRVPX4OvmOEuUC+Eenl2QUr3qccTWl8P1e0z4AQkANSv5RMa4dbYmT/0URu9N8G
II8L+o91X2fcD2JRIfYmQ3mPo2ifl6cmimwnyxCEQzys/WpzJ/h8/VODYlPBs/Xx
/T+2so7zncc91bQhxZZ6B1jM0PetFUtlnoWgWutJBdyiTy8HroU9Sp69mfw60uie
ZAh9KN8iJBF59GhLyhff9hZoAJhNIT1OvHdt+SP16H4MyCa+hqKZtdeO/dPPujW2
yJxOl4Bzn0w+FcmEzIa2HtEVyoE9GBa5vAwClAuRGqNY7kow6VriEpxK2KUrcRkb
SBSk9D4cLHEOGV6XC2tYfdPKEqjmn5ewVpkcHPM4xLoRLU6qhGJaXdgiO5nr79fE
wg8APGTU2iqDpqdkYRnksQ6Za6VgDSxIZu0R0dsenQmA3MFz8ijx1YMeihKoHEj2
kzlaeiawqdrri3PBCi5d2+erIswj/7C6oX7joRxaS3xpcC2qaA6IjEUBr+n1kp+n
xMjHMuf78XA2aPYLd9e6IFan/ClEv7C7yvltyXzsi8ShylXTsXYODdSsneIEA+8L
jygjqMTKvslVhqlbJIp6FvfWp/VNVvRBWqITj/mCpvkUe2cGuU+0dlSqoxQu2DGj
ZANypCxcv+duo/wpcMC5xwtzDx9Pak2yeKAYVtdnpnMlZ5VCqVubSs4Y5I4O3ax1
ej5drC/jdjTPeihzy+cUNLuPZV3o+4bXnpwKj1hCnvkkdVniH/EWo6On1mCTbkR2
k5qZcuSni/GVa+E+kMLM5qy+OR9+OcYNc4D+Oj4ZGQCaFRAkbThFL6G0/x3OQbtN
9NXGEOusmx/nSFG/CdsaVXNbYltLKnOuUoBM9rDlpTVKS6SOVqqWdZagtEOAc6a+
k5y7VdgzjTxBD9EHP8CsOlnOxhNJ6ToqGT5D+YoEQf4St6YXbJ7rnQcuY8QtkHHR
9+hIBZt+Zje7XQLEaQpoqqgiJwqYtUidPuUsQgY/JD6iDGJcNCgnWF5xm1OMcHAW
n61HapeV3g/8m2Z/B3y1p9xGOlSS9jfHJLe6bFM8Xiar59MSGu/HI1pjzCx6xAIY
cT4YkEO+VMJ4P7OX8dJAMCiXxeZs0IVOkx29PHcEBKuCmtswoRkqnS7JZbrEZi8R
bO7fcLTNt5wMpLw90r+atR+gGoGladrXtVisPdF14E4AapJfZeyUer6aR3tbczKH
JAD5R5Tk9Tw7k/opvY1Heh6hPcBYLagi4ZJ+k2W27Dc2zA1dM9Uk3S228DHvlFzY
iJj8nf4beMyBfaL473UUHi/qWD/+AMeMy07a1+dHAYGaFR5EvNf64n3mioO3U6+j
4op7SCcA3NJtZ96u6ZJ5Y+bY3hO8KG/mvLkVIGsyDusU1GtFUdpaf7RdP4y0j1UH
uzRGYySjaQY1CAK911NNhpYF5qEyKp9UdcxrowXGnb7vZBYl37E0bU+6r05BosUE
u/m80PeLNmwPP0lfC2Yqiig5gtLFIB0kY3NkUwaU4DcZdTrg0nQ9BRIQUUzlgg7J
z+dn5S1Ue09zrrevLyiaeX/oSkrlGXVmj+/aYixJiD8JK9gTl1OAcCeWm52II2ws
h8z9WjvWuBUCKMdKisLZn+tnErzbbqfnsYDHvog3C8t9YVYTqPUHhPrAwRTlzBVF
GyLh/AQVQSyUkaSC8yAfdcbID+9q1rfyY6HkEqsiVVAooWZtIJgJmgJ3CdmM/Pwp
bgyzHhuyIZnX5vevKr6+ZKzWNDwELPySw3RL9ZBx47xsNgO2xObT/wZm4L9SHfBU
aLWqsB8FFxneShdfulc0GG+yEwT4JqYjJQoZDYN4L1Ac24UKIi+JsVhb9M/io5Qa
6/J0O7Nv3+BfTOAcEWBJUVjanCbgqkc38y+V26/Utjvb9/zp46IQ086whbsKxecD
DvQmiBjtT2b98uoMwtgp25HkHu9uvoI0DhiWCEEYxfqa7oIV81lDtDNcg/PzU/r6
gsIOty1Grmxs46KONakWFfidlMcGRBcCkhJNgp5IhN4hDjYbP8vo1OMubV+FM8YV
uGkzn7RbuQru6M9olOfL2Lu3bDvX+0WC8js+NtqcFv8C0aFlzTckLYdyaxPnpgF3
JACoRcWYhYuGbixbkhrTLZHcQk1rD5qYBWxA3oekxjODSaEN93sw9cimJntJ4fNa
ltBd9Y5FCVGJhCeE1xw56R+j54lLdYjYy0rlqYMUxmoYdlSOUgbjrIT0IJcItCxt
Pwr0YMMVKhMgdD9VUjQumyVpNd5Z1NWbz5LmxVhwJO+EAhMZeol6bYYkE9eGViiB
ZUthbAFuSzxUgjJ9PzGlIuvxleDleKOcdyJa+nzkCDNoNjMwNyK3uBjsEuql2oYx
6j2ZHoiwebjV4lRljr1W/yj+afa5fvSEuiyIyYE2ScUaQJ8ApIFv29ozGkHW6PBV
ZaPnAZyGKviIZ6f/AyVDdE0LlzYrgNrvhDBvxPfOcQaZexgaNGNW2m3KgJEuKyum
4zI/MT7z8W03mzibZaLrsmH7p6f9HMO1vqbelf3IF2uz5u7aT/6LGZSTS1KiGdYl
OLvozpJzbvsOM8ynrjQPgZkznVQBRJZxtthXIZgwUvY86/U5WFV9ByuXfYUgM5KJ
miJI32hFEd+3EoWL4ss69dVV6PLllt44THLBd3rJHbd8EHibsdbtNV+beNtJgof2
a39gsPeQb+p9dZ7vmEo37FXwbgIP87qWSNAyLHE2FdlmkblTDidjVh+wu2MAPGeV
UrS7w4DgRGX1TYwueClMLlXGTzpY3ZK79xSQ/DRtuFcZa1PbUn+gbVwm0A8+j6p8
l/WuwOcDTbOk/+JKnXPyS27PEdTDCv+sIaWbrV6grPRdWCd/H6jbIrmAMxVAnl0A
b9hJpIu4fmr3cqxE44Y0NRwRypY2zQ7VyTQ59VCLYZ0dBlxDQmm4tIy8aardphQM
6ZSm3Ud1dnt9C44D5I7EKCb3CYGIDt7wXG05lhQYAyvtv/bQJl/62cWeHC4I7V4e
KSCJkoa8AqgHAK3JarcsmnYES8+OY4JHOz+i3O19yYgO+dD2YdQfDsQjtiqy2qhL
uG2/PNghveTA9zPvCHl1KpzxglwTGvTNgCAA5rJl1n8Wv9OwPeVrQ0s/K1McnNUM
YGd2huJLGI4GcQAAG6r+tbHgTvTfLUozlqmkBSSa3xjiBUDqGlNvCgna8XzFI6MY
asWk6bFCI4KnVwfF7UJ38ZnCp0VGKi33YswqGyExlRrP+CSbEJFErt4LcYtmkMs0
Qg0HT/+vegADMtNIgIjU1xil5jU2PvOUm/YNmnpx5Zh+ur3HocE8Lmc4aClNdrbz
y55QMBs/h+H0fPkSpYlS0t6v8qQx+7FTwuC7mMY4fpeqFe/2JjB4wUL4W4EsNiU1
IK1jjV9x0K/3tzTUbAdeZ5sakIcgUeIAupw6+WuNi1ouOhjM722XsJ/sPViMu4fj
zArQHgWTVUPoVynQ/fQ4r54tdBF4CylQnIIHThgcX3in4Bm9+BIWnZ8yudhvagPF
QZuqDg4KMJXui7tQrCrX9XUNHI0sGrkpSGCv28pktcJIkO7jM8Is8h9XV9opnuNo
4Vg3qw35Zm+TtOuDW/twrS/M6zCZG30FOj/afxq2uTQrtc+d8McHD48YrqSn5nt0
WLg9PR1KTyUQGzbkaMBVj7SgGqp20OFaQPOFMyUYYW/QHL9mDgMbNMYEyXgYhEHD
PodG430hqjzCEZ48VZ5XwK8m7oTot3uaVEnpQ2o7fAz9vJY0aqBY4w3YxPtr1ErZ
7KW+x3fO7W/V8qxg1BY5SyNkShevFqudmPfwnwqVCQym7vusDUgSswXGz4pPKB73
LQeGMeJfQ+33q6DorgcqtgDrIEfT+zZFb84cS4cWKdNZjveta3wdXIGtKO5fweei
M9Zu3ly7bGcXaugrxWISHeBXlCrToz4Ao26f3Wa3xg/0wJM4nTfgX9F81lANsJ+S
1zsqIv82atjmfMOTly4yz5Q0gRaE0+Hr5eDjRa2ejECh/DGN75Axs2u5T4twkKlA
ObMaBhSxnitsQCUnnLfJAZtsl68TKrna3cCbW0tI7dUs68Fq5hHuSyM2XNUBIcfw
mNq6hSUQpT58Mh1cdIx14HdmerbTyVqcQ+IeROByTNPiGIX/v8QvjBVSqX6GQDvq
o3Rym1Kn2qdmmwml2Z8mI5gM+PNoOBs4nJ+iSKK4rxYvSPRqKjeESj0ep3wzJJVj
XO3MosQX8OMvxkvtwmSfKr3Yvjwi4vdHbiAJZ6qTogARGXk0sQuOHWT3hrOC5Kx1
9VadWpW2ghXynKipoMRiU5+Qst43F0HxL4xhih3XIYVyQqOqdMjVdV3+qPTnjIZX
dGnpLlgFTAldrUX+dkCpcw88bfxd2+oZcKzlNuRzHN68fgGohM1p5xGPbyGUAtQ4
qcxZoCejXGF9GW0qXVimoayq6Dgf+1vr/LndteNayGJ3t2dM2klDk5Bq5zPrhYnD
hAcgPmHZf4+hNAKnRSvhe3THsqOyh3yhSGeuY8q5ovBKTDDwWQViCbgRPRle7ZrW
qsA95ToI2HvECNQGzGPHHX3kwyQoP5/eIgzSuzDJRdFRUpveIBrg+/lRdQhIIcxQ
/NcZ1IpdV0LxIuGJSgZjj6Br3wo1i0UhabXpzCGFONTEgCN//TWATPjc3yM5N+9k
/skKtEh6JSp/d2wsX5CZsxlAWMElOj4twtWQAwF0CWBLRKK02otijx+qc7HAPiuL
Pn1SgecC++QA7fJmwGoQp+26PChxnOpRQfU+xBe0r7kJO3PwFUWODYaATjlcePvQ
3Ca4jrFanuHhVWTuz5O/UF3FWN3bXaX+CqWQIX8UUZzys/a89+uhmjPIlic1AR6B
gARnMV++dGMU4VHFMsmGH8NjiLteaEgRuptDrxZMxWPPFx6MEPkul904dWWn4FoI
0e6yBtEkGkFZh0HWK6nnAuOdfsBquBrQp5QfaoHbGV4KVmNMX51AyUq4M9F5Mt2U
Uw8KLWr5EiCLyb0rA0IOoKI+VkTIXiAapAJT3G5VFYGcO9b8ttvFkbyU9Gi5Sjoe
e1ctsMGVNA7Fn9gNDY5TQDZmLf37ffzoAUvvddmm41BNeeAEk3PpMXbz2PClM1qG
YCvc5y3h8o0RU+KBLQjQhR0VwWT8/KCRC3tFMc1BN/6G16QQybjcwP8e0JjqJyH3
ht+0Jw+TeaU/RUxKjyOD+lK8Q7fSiGlmygHFixqKOvxO2jy41hztWVrxPmZGfL4V
EWkHtPK79vVd2xI8qAAjM69R2Zfla9vBWKHy70D2n2lkvhcbe7W5VX4ksyYF4f3t
T5BQ223pD9TmvNqLlP5N3bOqr8YUL9jwvHxGnEisX51zxA/I7D7S14GBe1b7yHRy
Ku6gPGZlw3+QCbmJkAEbBjh04pYLv7a9j5y9nZQxCouRTKtzR4UMj45eRSf41IUw
4zkzIJrnjcWtKHODMC+x/HpDVbh0rXs73oZKvQbGYhc/bJ9/7yaXQ2oI0/fFhi++
NpgoFwKNH+9upVreMCJ2Fv440v58hRVlI3/lvUoyCCFVSESaSCUzCNWWDwXFnTJt
24guEalXQ2NAjManob+RVieRwD3E3PO8LNYfXM85FttZCu8+0IzWpwmOXID6lMzW
4sd3t2W6Xzmnijz8VSYfpB2nya+HMCQ1xZ+N5T6EKLjqhHQgEw+eSytGi5IKx/zT
ivSBm5w2sQcjjr1A3CoI5sgtrvR1053jxT9WHQ+klmAMHW0UJ84p8lyZme+WGDfE
Y85JgnF9G3EeSQ4V5TU9UUQblH+IVv1aF/c9JjQY4+wBH+vF2/qNF2HN8+0e2R7W
rYIAg4h5QHwYhzlbTKHQg+WkkDKtzSqN7FtiMERZXxARPlGVt6E6lkfhpPjLTtDM
n2cncIFlMkxXjUrMgBmEtWlAaK1CCexkOgbzwtlSt+CT4B902vGgdPXGFn+SocAN
mFChlf0udyt9J57iSPB23qXY3GLXFF/eLaAQu4C4i11JlbLaZhQfzrF4vd0NC9Ox
KXdXWWDulE0FlaDX5UoTTBCxhRKicst7gMo6KlSKz0IAu56tzKymTNMh/WTrLzPb
4kArizOZtWK8MZm2NxIpSKthtLB5w30ap/vUCkoxGHmJKa3DQpXL/a1BALmThU8X
99nwzVkh9px0n5pGXUhY7M56W0GpfMrfM71p7NNArWyyFbL01R+ESs/kzX/oMzzm
2jo4g8T0uCixxFfZj4M50aEI21AeIfLdn3BSqMQwFQAe1ZYTfXKOlBN4/hezeiOr
AZYV7nCeKjjPiso284x09g0884rwTa0mSkSSFvncANekhvV51ZoQoG03bXecCWzb
h+uD4PzawfxIl/vAmt4mWylzelQh92Bw4tiuoM7pOUdWVidObdvrDPU4XHHTM16D
5P5Ce8suS8Kzl6k4S0vQ7SCknMSw7HLXXh8NivZ4t6RMQzE9LsuaXoyORWsL7Sfp
Ang+4Atfyf9Lq7y0r1FEelcM0WVMjxNvjD1KXwnkvTO1otu6EHJB82plgl3qTHAq
WThVr++m9F3WjVhpApMEVr0qd2kvpGIy6ivYNBESUxnI5tYCfOvoVKfxNia2WDjN
Jnsh6qXq+RtAZJmQGX0Img4pRoE/FQpOvsdSMH4rbPZK8hT3LVO51CW72t6icAMU
gByao0Q0m3CLw0RP4+FAbc9Qz1Dq4lSdrZBQPpP8J4+85AEgaFE19ZutYNA0ATlF
7RLKNKP1q5XAwtOyMprstXHR4OO1tYLvjSv727onlHNi0aVLTUfeLPWigP6wVruQ
KaClN7vKdprmF96YNfzd5v77khiHufSm978OC0Lwhwla4s+qNlh4384CfK6v4dYB
m22ivVgq6sAfa6VIOz7DDJu8pi4VsFCMLdt0RV/H0WLS7XdeKye4KiZjpg/Nu/6a
mTNPeHDxYRUd9psLI8epPCKTeTItiHJpo/A5HgHnXfKbzPP9fXxFz7yhLWigpQ+0
cxu7Z/VKdOi+njCWK1dWVgRLuuqB0TSovN/sNu5fE/jXxXZkhyRlopJ93K9ktktl
aBXfJsgbm4XnvlCVxmLnp+dhIdGLESyb9cldUIOmUpz6m8CKRhxJgGd6bw4Rjdlp
T/ikK6XRN9TiKPhoQf6AO+1eona4oTyLh1hw1uBZ16V4sxF8ql/Df4RiDogDm0Qn
Nf+NcRmsJBcho9BZYMghvfNFCkdjxnqoDb/IiGaM7a9Hh6/eV7aKpwDe+dAbBqcy
Gdb5KJVhZkft2Ok8kKUI7IPlWNEJ67rLaPgOjJ6CceKyby5HbqQVHXsYKOU/ZlbK
CT2kZ1AdGk/rI6kBl9TsrT2+d0JdhHkPNHs0VB7Rsv/rTrHu5YK3pyiL6jf6aH2b
uNx8REZm20uyR6nOrPwMLWpZ7gb3PN5NNBqcPUMvaR0A0aE0y2RznldKGjS10jFd
Py9XF1trv5gg8O+MMqSu77DgT56uWfsdPDEKVG8YhCUTTL24DxiEWYzp5is6Y89V
qEqoIPcMlyS4XMJHKsDsnpjeJFa4on2oy0v+fqpvKb/zBlO/sICbLkPBYuiZCeRk
c5nNBArai/Reyd3DhNoXqdSC541oWFEbVT51bioqps9eNjAA6vCju+LMGmZNoWR1
YnrzRFZjdtizW3krDS1rfNvIk+7hqyCz+H1trEd/O17GqchFhxq/a2F7n6CAPxDZ
7OoCle8wGXx65NRsLe0huoVvFHb16D8XBrgUXxn8+vO6022PlPFZla60KY7J3VVg
vnH+K5Mna0wrGoY4KcrpCI5V3TcZtUo4s8ZLgEVZVvDh6db//PeMRSkq+Xk6iu6f
2h06Ma4XikCRmweResK0beJBI9k2t1JukswJtmNl5HUndFQy1OVIqaZBwkyl0ReA
pamyrTmmZVlozspVP9py++SyMmSh7f7xOjnF2H9JJqmn3AnySv1JNIMoIBt7CBDd
mw2TFW4ojmcZPn7s5JXsxLZRH5eACUI7DZCfWt7OAU1hkAy43xj3M7RPXLCLYY8/
cAZr5TopGfXAL5Choz3MCkITRo72g8yvL5ENmf/9yOOKPVFhaN1vzGpKz4pk4CNT
spwmKxAt5XS9Iw+PUhAolsWFD8ZDefb369mfnbhrYGJnSFXoXv6w7HHio9c85fv9
Zs8htYgirNNcTVr+vWqbzMFJFow8L41YU+nGSqYUA8yalhT/yqfV7DJ3rJv8mj8C
ZtCL3TUEDzOkhU3zXRUkHSFnOPikMkSIRyq8JpM+TDQr57nXBNb/XTt2hjne5EN5
epc0T9OD4tUjnasC7bit14xajHPwUDLrBpLHgyUbbIyOU8EX46VFPV8zUL7GmNPc
nOwW+KtxiWlL2ic4SgSFvMdhpUqJYE7PMtNQvj8vp+HL4sxzysHO8hBVsU2Nre3t
Tv+J/a2qSBm962LqqQ1bLIwRe594EjgWCWxurm/hCXMLptg3oRvjyZVLjlbPu9cd
mJ/ysrfrhRB5qDWVIq7vQrf2BxtFawWpu78+REJzk4UZ82gx4qzl2Y5huK+EjVHo
+DECixlRUp286C1sI5L2c3e6rTSoQ199k0iqLWUIO5W7mdDKRY4HIPstbWQ4mScI
M4QsGyRKTo7XEbd7lbSFCw2ei6qAVfw8KJY7YQhnPkhFl50lZW7rk64MBMQsCx5u
d00TXWGwjUbYeOpfIzMpZObRndIK0kPZbc/lyAfW220GOYYF1tcVIYDeHostR3/y
/9bbfdTXjF6hGtnI/DU3VtrnSAZDP0/s7kza2guPXCzHtortWrsekqbDWIJn7l2/
HbChQ+KchRfLaSFnyBydImu9kk0EwVvWUJn4ksDnLh5Bnyf3z7I1odmIDfwPiRBV
sY3s0RtUrx8lUG+vEphPvp58lfGwsxquyCRuxyXianB61kF54QFrx1lzR6UE5n8I
4NYEO4qHaUTn0EJPc2Ok8zHipGZKAYxw1kFGI5Djh1hG6Ji90QTjpBReu2gPPJic
SV97iu51juuwB4j2Hsr+w+OdUqILuWmApnANGbzIT/EMvGjzKfDId8c43sed4ppQ
gg2wsKQzzIkJ1+fHauCVRUmM8MgEXQcoZ5gEITnMyQAs/TH1T50jaERo17KVoep4
Fk3mBmR787PZqXFUfz0vn8KCJbTd/gPUom6rP9hZM8xSkeGFMjUF3MQG+BlMGCY0
FeAVwFe6C+H7ZkSbv71k6UqFJhVGUYrfEJsi96wngBEGmRVrfjL+zvze2ayT5xxS
7LQ3aV2g/RuBYYynyi+N6ZVhqXC8xaj2J5C92T+wGqideEdw/LnfrnLSlO2aiBbJ
boiLojxSdVLhOBcRS825jJhgLlW4xRcwYw1jTRO+HPxjEsP4nkZ/fk5l10S+6hrL
hA8iHYnOy4ZAA8W+N+VjPvqwfYoX/5local63YsQZmfOspZbC+32ypVXWwAR9bNv
0uZ/9LoHJrMkQPJ6u2OUcwkFU+c/wke5/QTezjg2QV2IVVQ1j0juTZg8pvwJKM4j
NjeUr4h8UczW/7o4Xx0Ry7WhlwK60Uh5GGaVAbyRY9prBSFgi2jR8zdiV9iRkRoC
G/N6LD5s39WPv2TpUXhZZNPHxsrHTxLkCYZdY0qJFYm7N4r8Tr0JOs7bO8zTS6PM
gsRbyYTfa7u6oMAGb7caZRA7FUDBFgnIAvZcnATsaYgu3BO90y/w0EFio7gp1rUc
58bqLLGa+ysSBot24ynMnMGqk7jPortTStF7VqxPhiLlIL8GAt/L+lo6fVf15rXH
yXxkTrpg6TrUgZmGBuawNXC7ow9XIwIu4l/Rzvv7zi0EsfBi5/Jd4LZvjn4rP2jU
OKiJyMX9HlhycH1JnxjmY19gNvvsGehPnB6xske7NJVjVVBc8hKBcfmM0ujmX4R/
cWIAiqD1XnAVJUWeKMU+Uc23V10ncrvmbr6XUXpxPlUc1UEFiLCpNmfLNmIWOD05
1qLjgo5UY2kXcGmYQS8WYbqvdUb90ipuMNTv62vlU+OzPfuwzte+Ls5q9lHLfxMb
KBnWCC8ZI+uNbh7IQ3a8vSNytIHtEMnwnwej5po9MnjnCqCvz3E/aI98WKSuYyav
mR2/iabAIfMLetYniKF+XgI7e12GIZc57I1YxtrMK4raoROWMVdoo3Ch9LbMqn07
Jhb92kz7RbMemzYuyu3qLRvui36kfYOFeOisGgsK7dkYSxkQlaqsOu2ag7lUi/s+
hxkQxfwWrOVl9Vp/TIPgKvltDW02hhf2cssRAdBq6Xpjtzp3A/kkY5KmLwuXy0RC
yJwuvmrEc96UdgfLy/9vf/sO5dIWRsj1yToRRjjqwuM2GXzbWOx8DMrnfH/fcTa7
7kDLXM67WFDJbrRQxq+oDzMW9Bhu0t7sZOrU/HBbatxiiIGAeXIJtzAFfv4DNvRc
FyqIBxY+gx0HgBzIJ8Fzs9ogko/WjLzxia4fdxozfMuX4V/CCntK/L046KnIqnRH
1GSWRbO3okyTxDPA60nELHX+yikI7L2Z75qLuSBxh5FKbE32X0c/15ntjUFt42vZ
56YaPWWr8SerVmk/jL884YE3SHVVlBEv8j35ZmWgPhF9sZj+XjAOAf1JJl2qqWat
GjyE8JiXKo+2xbXyNitQ5+PrNAykuX+yBiP3C2+cIj0UAlwc0EwmElAeXUPv8+pp
1LR0snjNzgw6lCzErA+i/THYpQLPjVr0fzczHphf23cNayZQshZK+Yns+EZQasxo
QwzEl/VEh6kzGNTjPVJqKChPwnfQdZg9oJc805/WGBjy3eW9KUXbvyL/eEp4DLW0
yR7Vm6DgnklGoE1IC9qTjT+8RmdvV7phaJMl3hF1QnGlwOFymAG91J5ix/r4yLxN
h4CClUKL/5+J/OEOdgv1A4lmaSyOCJSIKtHf4npTcG0Eut4eXCCfCtL/ksvd1bCZ
b69YaoHK8YTSpmeMLTvScVUdAwjDScosTRzUjihHBXsSZw8iMzLb4QojPYrSg8px
tzTWdWAY7zNtPq33m2lcNSXGP/ZPOs2JGKrwhoqS0ls0M8PWODcI2W6N4e2W0FbK
PiFadJ4GYSYYenMl1QR9P5uIIYPnaqriUIfQaxSDR4KG/hzRjh4JZE6cm0Jr547N
eN0cXn8S283Xdf3I+N2zAS+gS1sbNkGzXfacHY1AfinsXq6CEhnXytTO8rOY1DBA
z+1PjTBjYfUNPcceFmDE3qYFbaphi9uJOEehKNc6PuvxsWal0pO1b+gtPL7tPPWZ
wRY6ZBUXdjDez8DtU6ZUzUGs3Qq3kyrq+tZUJ/iktIEVoaonfPIsoFdWqOX/QyQx
J9J4hiXcKZcfl5r/X0La6/4cdZbycph5J5IWjWT64lG8Zos38Spk3gos7MWXwGcB
p7SmPuB9zCd/oKttrCo9g4G1DYePstCLDULgfUvH6hDKYiy/i732/RRl8ghKxRW5
dK3IN/BdbL2GM7B2rGiDI6A0uAIVvTbEB5Df/SFW3Vtf55HQxQ7mZ9uu4SdsunYo
guQcHXuQwdSW/4UKFj9xPWdSeWD622A27ZuB59BpY0GzWZZk4ZpcytSn9nVpRKGV
qWo1fMq6NyPBCXBTRDnRupPXZoVSNTfDy7YjOxNqQQXq4A+0u4W6w7U5Six8Yz6S
vQU88oe0u7ukW8IshpI7HPzkLsng5Mnz3rrx61nE2gglJ0otvNe9Pmv3CooBSmKe
bkl92NqMZSpARUKjLMQBsKCjtKkoI+KnwqcDRoNjYRJIrrF1yLOwQ1OKN3lqTucK
HjHmAR6tdARAtn0P+QEh/4jDL9KYkoB59bfXOcmcuWQ2UWOsTLJm3IE6BKrj92rp
ynZwBC34GGSWD7JLU8QBAApN+QY99fPAUmvlWT5+Ekr+NFe3QmhTriHkfdtcAdcf
ielJqIguLAFW47dkoiJpdpD91eOO0/ju06e4rjgWUwo9DCN2PedVv45OsYD83eug
08yl8Y3hJ8WVXS6JFgmBZ0f9dv/rGulnzExYrlzG+PRtB6YphRoz07ERgNMiMRFC
J3cF3zpWlAmEax/UkgkaEnUB+byQ8GeuZSKTKs7LfdVTTRHWhkJx/calU3Z986qR
Md3rGLhaO5KA51R7phdjm3Mm31B2J3yviAGkID0eKl0BGnC9JepDGh5VW21vOOFM
gkTqdj26s+u+2MwDYS6RX6p67nFns84/jxffTSxLEraSTX7iT2eZ/V+ms7L83XKx
OpqZk6YyeDpDo9YKMMGz9jTSDI80fxWOdl5VZXv7uTfHEujfKvyz7WGy8tz3ALnC
Tp+T2rI5mMJpPqYyhg2qRk+rNp7MY50fZCvlEPrdKJM+Qh0xSX9cbE8Mf+YjSzww
LAbIVul/o3EdTNQje1owFlLAE39Iqjk4QQ3MAGgKtfKczw9IE9haRyJB+6oLkatb
Vup7eN5OROA6L1Yd59erSqUvJS9v0Swzq9AhfuSptyodQAqJpHHPRMOeLmil7m5l
JW6bgEMZq+/1dAc/u0Voheo/VwDeiCtBabBsCdAtscSWEEDGzqw7oae4lbr72s/c
IMohpGcvqujGs2dRigHCbRRKTtWAu1BoHWSche0LHx3VKTe3xJSq3WOJWZFnbfFy
Yf3kpj8og3YZq4P0gFqoEIsodWeMOYKo9xLdFEuRGfo/y0Y2rUkzkbg3pMF2RLUC
R0Ewn1Y1ZPF8Y7DiEish6QRSUVvrKQIl7+9bhbiV5Kz7pTeXUTaCxJYrByDlmBCg
6zKm1zgpV+zp8yX0JBbT1sujbPjZ6hHcE7yGLXYefY9bfcmdCI6pway3nFNgWme4
ejIk3n8akMWrmZCk/70u7zbPz8fdRiCYRFW1LtZCk5+G4Vh4aPlnVpGO+1TWCvMb
6133wllUhFWPkZj0wiO6SuulDNzX4nCBQHNJus2+O1BImWbvJ+kAKF7pYRCHMGlg
dEdbtG6CCf/2ma0CQkGZX+S/YfIlEsGkrwu6R9XlOidHg9ZyHjlhZK9bXjfAcy/3
tYqXs/XAjn46coddjzkAfgZ1uSMXAWTaOofLadh9x0UhvEiTHYa4RVQ7SyyXEeIw
0+JdCur/eplpfSgpmXA2VXKTX25YIwIa6yvDTArJXluJjPwwRMz5uzwkPRllrG+7
YXLcpmPd/bgmQyalp8IDKfdUi6zaBjDTdhFZM0/wZ8g+fDCqZnIERxlZqwbDDnnS
Co3ZE1pgZhr1XhwYjCx7AUVMXK+6hiP8lqkaRZHFr9k3xBaPpp53Ozor2f5LFW1S
UfoMSoYX/bzgp87inBij7P4IT22GhhOyAazoJHVSN2Ok3kr3nw8tahJyiurhSXJj
/c3cdO2tRqbm/aq88Ga9tlZgc2yrj5IjpscEAOrDfh0wbXRXeFuCfzmq1V4Yntu8
zrxA6W3iAwEJDfUL2CwI/2qfOoadytWOd6xM8FygUMvFH0KUdMcPGgF/wZek68Bu
5p4LyFgEN9o+ourhoyAE/eo46ZCNdCCWFJNvrb4TQI8wPv3wOJIRURsfsP8TW0TB
hegb31VYATkGVb4dWfld4cMkMqLVqMxm9gdQu49HgbgrdmZnDx+w9YtQZbCFVEt/
AqWXbcbVtbS0uTL3vK8vwutcnPDr2LkIs3+aNottERAl64IYojwMh74JWH9gGBrp
yt8fwleh0n0lW6DED8UescWFROOsvpLFpj6M68d2EGW/Of8P+GqtxVeuwF2M2tW9
TQbM3PIZ7KaQYUqENgKyh526yQYc+FsToO4E9PPAVrbQ/w5swH09KojGusVSHnWd
06gfL9fX7jhCJxbQaP6XgRsLLOIVkI2dpGiAfvMFaGUXhibtMUMU2KXonHbRd62i
XR2MF9/2BXUJEILHeTN8/TeRetUM3YEfBa4KzVIr171ByFw28BodfI0ZPral/tFQ
ch1NGZnMc2Hyqf9k/1VYduq1vUhu3xYTGP7Qt04+bRt4i4XUU+YT09aM6Whh8OKQ
cvNIUi5j21muuB/cUfVz3DqIbfdNigEMK36RQt3I++4tC9gdJuvYT9KHaCdvbZtC
35PaLguZp/ijs1mpyQxEo271LEtSE/bleK+fw/3SBePjxdU1evEU14OED5u16ix0
0F/+JKChjiIPRg5RsGlGUBWSfgrOZL2lpYuSru73DIEMHMiJGrBmYfoQZwH/Ra2y
/hz9eX8Ki+//1r7XYoGmiw4jaYia4TT5zvc6Fh8KyyDGAnLbaswO4mDaEDgkcHA2
0vnimEh/6alY26B9elo/9kAHDLavA/wH2493bQMtgm79Ag0xfuU1LwcUa1J7aV47
/la2mbYel/7dwtFRW9Fv6pJqYgtyyI8fBG/H3xwDMxFLLi1hpyhePZHdPJuMQr/7
qN+Sfi5FfpUV43f2/yVFmzpE0ha2DO5mdE07U7vdTCAlePcigJ3s4YG3xJ8kZksh
xGOZ+YaIvz06dzFoXoqFf63Q80w2SVeSnkB7k4ZeVQ8MyEFNPQMZZLm6h8xrhUJ5
OHRjqFIvzaqHyW7RsoJp1scIiB6TscHwwhaOHDWhig3jgj9hm4IvMG9DLq6EMjWG
GT6eoOlJKmxZTVLegpePOdCrKXCytW8sDZ968cuCedfP3JSrvgIrqFswzosSQa3n
rHYqYdOKjS8gYKZAxnp36wLMeKWACBKK816JiGmIVVTkvrFPaaJ4OcjNd9J3vxLA
cEP80Y9RDE+OkocYGJy/Boa0GpZsOTWq71rAWJuk26ANry04DcF7HV6H8CmnYDJF
o3cR+943RuwGYlUb0s0zIKVfT01mNzXfkXH5QKika74LMk4POFYJQ6qMbgGjPTzE
rhswkh9/L3J0ApbdS5hH8Lv1Wy7na2feJkS7fmtDLOjPDonQ2nQnudaG87h21lSO
OCqpFJ34cycEp6WVKoryHOJb8hbXPtpmYUqtB/qLbxkku5qDfEIf3DUaAWnm1Cwq
ZW/LICGY5dstr7Kb7plse5TN44oJlpNSwd4sHmpw7U2HCNaLBkqO9bsIW7Pirrhw
vo9FkPDtgCjgUvpYQVz++kr6al1aYeBCAmcXzxtSFSyvS7uKnOPtyukTvJNBHwH/
x+4fpGa2+Zso3n5/9p1DqqgZy3/0YeTMcMW/T4JLImfjD6S8WkzYPGnMmOIfYXZQ
IMTA9wKUg61JShM7DE64MDxolRd2hzqsLB+LZ+LHu2vXjBkDs6CvcfMsG1nzRYYw
UW+bHctDlzUnN68sIVIZlpYtfLyhN3pubkcSLZ3TShocnNdXrSbD4Ky6XLtxPSnY
Uc75yirdUVQrQAvASR1rHbn2Vqb20LyGG9Bu4LQjZ0DwURXzacX6IGiEwSRuGhos
tz4B+Fgi55hVq8WbfLi0wRKCtjDdSOZU5P7u17IxmVlcrJyEe9coPlrR69xGYuoO
zF8tUREXnAip+nn1cptdp7BEruGeFEmyy5lI8PHnzXLWVD5dOuQPRBR6SpYOS/Qs
jDzEfb/pgcdD0OOyrkd8QwgIZzmTdS7c/RV/nPuEIYHPYvqeouhqiqu8SeWrFtb3
0ayYDJ874j6NUgJKLR72LaGc/4K9g48flS4rwpKLUhLAeIhYX3736RtCn0Pp4tyY
GS5JSY8f50wA4osvc7bhnksSwvjgdXTjBexdDAe7XYX3qAzhbirh1EFduGxMtrPV
ZXePUmKH0RR9sgyXzK4XjtEYyBYy9bJXyN529svIQWcfYovN8gfRx+kmwJ0xIYI1
/7ikMN6fJrSZmaaphIK1+Nj6hRKy/gaOYdWZGdXNCoE//19lzbdh4eF5WQ2WHk7w
/7716PiBcywJwpdXOiVLUZ6/7V1Ad6nJIztO7dfGAizESOY8y2gUZqaaAT/YfboI
nCPdE9EGIDAhJbXigyY5j5uF09Obc/rZScPqF7pfSYZQPec0rnaXPY5T1L+PqoWm
Ed0MudQzdB0BKQrp4n4L44BLOjcWI4L9eXz99iN2YwrEmxgiVLUL0T929sOBhEzG
KVySVavnodIYYMH6fHguz0KDg0noaqt/6BNqlfRQ2tr+Zy9ZWaqf1bcn0sH1+pRX
YPsYp6uzySRHG+10phu23Xl8qtKa1hmPe/NYFlZWuuCXjwdcshSa+YGdEQ5H0aC6
Sr9oYs9qAaKIHU1PXfJ2agQ8ey5JEiSypBq3PICHqagpSlNkyh0eR2Zm8w6ARJoO
e7C7DwYYTox6BNg9QFDlk2Az0XRDSuTjfUadi/KwcE/Yf/cCyE4tDy6soAtEa68i
+w8Ea4x4jkjX8lLg9cjNWGbSuPE289LXl7tqu/W3ngJ55jndOeriNQwZivysIbq8
nzJteZVNKD5CHjlxhvN5vEAibvWl4VkmKWoyLZhs+3a5sR8sjHoi5eYJLrdD/4J3
Ndhy0xEEYea7pKyjRbah65di41DCv+l3iSESDSVaB0NRut0SeNOA+DgmeY0Yu+PO
ntKlwomQ3Qv+dtu2I0OtAjGZQ68OFvF0ClaP3L//8S3I3VcTt1HFgpEMz/sB8aXm
2YEMK6zrDJfLISGQggn9E5P8TYVpEADlQzJBWNLc890doe/nCeriEjxtHtiML7qR
/u+4pnko9CCfR5EVujKylah5a8mtOv4SpNaTxvTtwp5wHuNoVMQ2WZySnmXfoyyb
mXKr0FW25Kzer+QBBzaEf4Sr5UOg4hcBkr63qveeWmxyrCjM1h+yoOcf9S4NFB1H
s3ZViOrVlL9zwzimVfl1As92+e9y5tqPe6tLsNpAqj+YVi8QSlkJZgk23iiYDz5u
WUnMpfet6llufYHs08BAQUV8JcEswNnPCazMvOYnD0NNFvml/IxDmNICApj1XESu
ZJ2iALxtArA32+oOK1HPOwPvJ0PgUG+Tr6wSlr1IVa2DZKcemjHZbPyK/wQlTNDB
+fWHEbCAaXWXT23famv5ZI9biV+ul+oqXwjD06+0KZWOfZxEBLLb8UikKRtwt2J1
1mfpRiRkU5z36wY1eYDf05ZOIldik2KPPqFmDbLWxQwSXmYXX7WQ+0NmY9jyHCXm
cQ3iO7gi1dWBUn/hBUy7pZCmlDrF85goFf3DrYAn4uV+XB3O+5p2WQUzvg12IJln
IH98PKtgg6NT81zUiBSUu082m0NhXIkHHUQhM+MRsZ7t22huMDNbp42TBiBO/e79
uPnM7XM3IigLjOncDtl5aNSZsIEThRE8Q/7boViiu0hXL5emRciReqToU3dt+uUx
nZGLtdhj2ESYUByGft6hh3gBKy6fzwxkTOYamLMFZyMeuDfKcdatORD/ty9MaToP
qdDJ7dQgN9KAVNit+yJHfD1IoFPTOvc3eUjmHYn3vGV0XcRiFoBsPFBl/lYaruN0
HWOfjr6yXoUVqcN8/iuy0P2lyqRJXeG4vEZinFDSKlANuP6WD6FgfL3HtIXbLUgX
0h2I4kc4694f7EcNfHf9UEhMLu2LFTntMrgIl4LtODM9rCwK6QmV96MmggFZd4W3
EDMXe0zxSct/JoHedUJNIaqvhTts9AnTJn2DRKYpL19GzvGJjSdUcNhKHiUSncGR
fwLdpsqp0jrsDjD0jYs3oTbO52BTPJW2gwUBlKszfL0fv3QSPOAcW1EDuf7O76/r
lc98Jw0C+iAUoR0zhg0N8AG2N1HldkrCtC6wchdJZSqdWh/3Nrxge+Zy8hD7fcOJ
k6bRCmP32vaHI9L/aMjyN131O6utuCJz+QLkKTmeCI7YJZr1S9bPMWGuZe/LesDw
giMxUVSlncoztP7exK8/yYSWIjVungnNQG4uoocGa09hdhaDqyqNZqkf+LGT6C+j
nHRx6uN4N/QmuWlhU866w8h1nsCbUcicq0h/KJL42LlRsLWE40nGoWSo0oyppzJ6
Hjs+aTDvQPjIJc8Bs82HNz5ncQ9ntaAF7wYIz8xHgV/BzasPZVzRRjG8BtQz3cRL
O/WKPjG3bDDi0uzyT9++AX2+ArLk7JLaDtS6RmKDV3kTy5Czs0C9jtkY82Uc6VEy
4bO/fhlYG4zfdeamA8Gkmzf3rajBRmI8Z6NVCePZNn5Mpd8KEhNj5LdhUig2PPU1
rGSW8aGSFoFGfr+Jq2RQWJjm8t2owfY60ALbsllOCqAIhkg9HkzA4wR+zEnnZtKc
oTwYR+dGdUbL8UppSR7wBYLV4jrUh5527MsOOj0aNrlBBMUefmtYWirGIAAjhOWn
6gP85H1893YnVNlCCPKZGCxkYKISL0uU0qaVWESNFfEvvKxU0L+HAp1ct9uGWhni
DHgXbKatETFERDDCwERRfWfLJyfC6Xcvnjauzah4Oq/fF6yWSpe963GFPbx/zQLQ
5GIHr0dlopK0APHsdBAQdRw3K57eRYzIcZHlMt21HNuG7Gr4LO5Uc/4D72RDKBJ7
z4sKn2oYciT0vJpt8HovPZx46/5hy0jOg6fx/JYq93FSyyMbdUOy8HiY8IGhIXrX
C5iQMPJmQsxKhiLlfmsJyNwsysq4UBMR2ddzgZoEVPXzXhsBMDW4A/uYDV8UoKTY
CT5GbdCyeypMfNOeArfgXqyW6Mg22fn0tJER/zv7d7I1YgweSIYbJeZHjPOq2sr9
DHjStAOlwWzmYdZCt68i4gQJ5crTuoUWMj70pXsa7gUUBA0ulFWIccV4WlTK2Wjw
Gp2nDE7gretZ/i3htKeaFovH7BMcwt+QjOhkplrLi3lN+UkYkfq+8Fe7IX1CbPI0
5FKQBKvzGjU+nZZlQOCSH/vb2hnjqQv7Ukms9QmpMYc7Q1EX4rS8EJxtWYCJ/dN+
F777HwFaFYPz3joCb456lVXsCvyyBYzn7xCOEiPCCP8y67IXoITF092XGoHXkOjZ
o/hX5m6fAUE+fTYaEaED6m+Apz4Z6WtqQM4zhJIQn0jiySh+p3qgWp1Gd03442+9
bVmMORDNunT4cC7Gigq9k5823VhM3SUDst8tGeQSGkbHo/MM9VLihhUjcyxqhbOr
XCLicDaW3Ep93hUZ26RRqw1DZfC7B8C2i4FBpGrG7/UfoAluKJ7EZLvixsSPsyNP
QadaqYOe1PNrYKONCBihzoDFyPund18zGcHRAPDH8GE43fTm1W9rd2LZH3a62qNG
V6ztOv9h8So6zbiTeBnQ+8WxOUY7mWS0g7qgV0NYbzjapwGXbPb6c/1lMKkjnGET
N8E7hDkH6pjUU2PQNBByx/nJhxSRsjStYCkcwR2sedk5ZEqPjIiYwcfMiEE8KdVp
bCv0Tgek8X9rmcIrPlfWa6J+t4ZRTO752/N6oXy/dnNbBdi7rDVw9WcWIR0Mq6hk
XydLgkMk9nWpTGGjbqFSxsU4KQf1nD9nOV3sSdSZ/189W++bhAF1jGfmrJBlmfO0
VwteH8gxaHrgEaB+8/ye76tgJep8ryQGvKKtWNQo2DdlWoz6nJirzAiFNLYendBB
6kkAxWiQQSEDeflCaJPYT55WqqHBF7cN3lwxjcP95nbN2fOMb5gtkdbzpv7guGk/
pb4ozThPWKxKs9x9jCCFuCgqMhF0jqgL7entdzPI3Ou6lckAllZhZW6RPzXBc5rB
4TVGq2M7wTfaddHaZXV3tRaB/+I7X4Gw/SPUB/2Y3YNmcoyklHxxoBfLqa40zAhN
Jo9OqVpgZoZPz+F62bDDxMtIKGCon7mAfLLvRrjooOxMoXcWRGvWiGHsxQvzpcLx
8CaIrRhWv/hxee8C7LDjqRfZLb/MURq8v5+hD0I0pX/TdX+JIbYc3vlQvM89RCTs
nvf1LBK711xiBR/J9Q1vJL9LRzsB0X5tYeJnJU3RBcPGeiiPG9qVw6X0iKwlZN8y
tRwnbi2oEayyvv4lImqHT3hrPhWzWZDYU5HaHg90B1CXHedgdsKp+BRKE3cAAw2j
VFWv7nLHc5HBOLZIiTqA7iytvw4XOMjC7G21+VEhipUIE4G6mfGDA9sFZfPGo1hT
9ktpBLeEowb6gD2MJdU4XWfxXBAx1/fOd/80mH2OntRY3F5dx7h3ca5JtZDE45fy
fS+j+cagPXQatav5cC9Bad2UMjnfXOWuqjme7m0eBYe97zuFAr83YLbRe9lmt4rF
MTSgokntKfsnqUKe96aSjgIM2A1nC0qj8SWRRlQT1rkz72mVls/Mwkr8EjYrUvmT
/WmGwtxsZG2fCh34Ex5RjRetHLENlLzMJe9B2c3RV7usz00cug+bvGWvsYKB0tCC
h7CuU0EUPi7BF/6qhqV4x9EaLJCA9kwIbo57p/bRWKlehyXsc9lqh/Q+5OyJmUro
rBT3pJgMbu2cl5i5mYni0lEBZtgO7e5jJutrl50OZbQv13zcqKOPTTv/Z7iPErSn
DEicMfL28OPg8k2kea46dvCJ1ixsKF+F9LT477EzbG7TJZeGZ5HPhQvHUvwBpMUG
JKzBmnpE6ak1i5ODF9Tblc1MAB04eRFhIZjfRRxz+yPV8map45NxRONLDi2kx0+w
u9nUH8UiF9QsAbHdR4LpnA1PNS8yumHK5aS+9gVUc6GQnH5TGTejYn+YBFzbrUMZ
wxSkTjlHhzsU2tDW6y9jEdChdv8uc0nolfGoaKwlxInh2mfDHihRssmhxgzPC+bQ
WwLBNUdSKnuKRlsnspntphoBf5yyoy+xJgEmkbQpW1D4ioTvtW1KNQdZmgPnsYSb
Syh/5DIMXa8DBeuWepdVeTP8vZQcfCGlUJNxfm1eDAMKQt4LQupv50gNS0SwfgCH
ezhPL8b6NHIfrz/ejs2ypU9SzIsLQLeu+MosIKb+4zUUy8Cwz1NHRu898+JPEXOm
hJLS7UVH9LB9Qt/dFuslI+wUIjmEdFDBjvDCiqGYUynmrcSU5n5TdAFuVh9MjVfB
6Ut27qBFuNuqXiAxrOJZhD9GMXLd0+cwuuAnXpwrI/YUO99VtwlWH25gzKcTYAWN
Tyn4/qGHl+0nvC2esDPUh/Ogmv7Kv58JQCSLPxcAPKh3RI+E+wxcjVRfJ7ovSEvq
PaKVejF43xmgwM9bYW2MV40IjfabAIGW9+aChOYwLkV2C4oqCJ+wF8YPJe8omuEb
3GlZUEgs55OKL9PX2l6Twpby6wz7bQCcfXtlAKxYIBkwHFmsWmw8Pi87XyqP5EAx
IfXdmjqz4CPt/aHBiheK/0MhXAI8zayxOizcDvKAw6vzeG+AxOFWUYA6ANt+bC46
2YdjAfRk4GEblS0DYxLQAz96EfgpR4tAU20PxzeA3ZPlpsYXcHCFKwy5HxMU/+DK
9AnWZIsD2uL3UfkGZz3Rvmexk1XMCEl/XDtVkQDKrQ3i79a1ReivR/VOYeQ6SSdK
kG6JPpfbdvcHNoP5hk4FlkZyLZVx0qG3mdCVDJ34PYC7Y033TtlvVBu6woBVTaYa
FyD/oyPpsbLa4jONYyfOYSOa8Xg+aVLzKBUXyJcoiY8Dt/6iboSiOANvX0Ki9E0s
V7JrV14/yhxpFBScftTdZDZh7rvzQF22iiHpR1QsStwLkb8tKX+0uszai8p2dRtt
yLdqGs5+BFyz9R/4yoXi8c+hayxofASYavSHXFuNs36t060IhhHqqq/TJGPv1BF0
c68xYBSkeT6ik3gvcmnvqD5VIyv2nXIe2ddaeR6fSQCMVCPzk2RQzSvsUqfOzjIw
FF7e9CzzD0KfFnrzzJPdvFbzuuuL3K4rjH1Y859TEBwceutdChG1tpb+wAQIrAL4
5ARklfixOvs4gaqWHRO4lRXpelRvkN4k6guj5tb0ewm+j01B9egVT7zPWIgTh0ap
DNVFfczmngGXvsbRjCmsQoGNREzixpqm1Xqlmc457YGDCGfumD9FhejWUNBbuPsB
ZZCsdwTpA3aVsUDFy4wQ33Lz4rOFXv5T8WNTzQjFjc9mvftN2BwWCB7KWoegQeXq
e8OnrYXXl/CwLJdh4RKdFtnLx/4mdsC8LJ+N6DcJEzboqiQ38md7g9wY4q5noBDT
ndVyh9ebruVMSbyeycP4WWTsOKdQsg66uoHnPctg+1YtUgyswU4cinBzBnnAslG3
+BHvnBa4vO3T+jfnlZPF+Nwd5t+WmsTY6yTJVwz7wbm8iYKjthlV1dlXRtVxh5K3
mgGszbcA5/AqOCpwzKSxPOXWyhFGieNQIQw2WGSs/zCVnGtvmUofW7mSPCnGk7Wa
6UCPuGKZtHSv/7jvzgzOIUfuWpIdA3Pfu8alzop8l8d/2BaT+6HKsYEybHVMSK7n
yZGYpSozatU5FX65lytP1Mbu1MITQWs6vln1GjJ3KvSXDx0m7uYzc80vzBos9GuR
115nWYEKAj2ABXiMhrqMchnGvfar7VM5E5lynPJdEaptpkAFJBf4bgdf8unkPS47
UDZBIDXR8wTIZJD29kteU8Qpa4hwEqlODmFJnrHLH6fsC2KuRd6mpC223v0pECG1
Ph7I6IWCyb1w9UZNUrSdNb2jPGFe6IpaA/vPD8EyY3th08BcsiZjf1EDdh4gGnIa
dVFUgXLpRbKbfPaF+lw0wO/+KQXIy2FRUVzjwwSsIpZ0uLtGWLTdDcbtc7L4wEwL
duST021eIMedltwUFBVxhRXPTWQ2hjczA4OLP80jNqXKF3M0G622SwgQ0IJQl31G
Y6BfNYA4VSU12t9kH0Y2lLDdRrZXmxxNXms4sNB8mDkgbx1j6bJj6En7Bv/FqqI0
Hx0iHtlf4V88S3i60A5DL3goVH2ZFedgADFRMhefG0GtgIkjO2B/ZKc1WPAF8WUt
5r/E7waJRTWe+dKIBXmNqE5EHQupVU0s9XyZ4cWvzDmWSDjR54PFdYoEVSD8OyA/
ZNLUqXCgyU/A7Yj+SqOAQ7akykJZER8ygnZUQ36xeE5JQukbo7ckhpemzNIc343Y
odEGGMNOGLDdqiOIjU2PNCivkKC1hfWHEjNtZ5ZCzaeLXRbXGQQUqggy8UKvbhc/
ANDE5ITYUIRjV8XmRO8fNFxg5gGMCgvCXq/lxS3lypyLgb5idvW9cubl17HqwPgR
53NQo7Ab/P5IsmRPe+S0p2f1UhpK7ZdBH5iIKI3HlvD3b0yVz+RyMLADxhCpLu71
4FPNIUUvaaNhYWecgYzoeQ00E5UbFE6ypHAr76DZyzEG29Q34cILONBsjXb0iIco
pCDhURFbtVKIg/3+kCaDaVHN92z1r3flKMU1rBfZdl+eY51U/WQ0RAWwIvP1b/Gr
LBK4jE5SK8RWT+rRkjVHLtkA11sO1g3tjC5NFlfGl4ci2cM8La+ZMMXHhoYrwdMi
QyJnS1i+217khdh7ZQCfb7P9NH9FxwfNX4QLJUnvID40Fxm50+ye16p70ORHPwAD
7jQRt0Rq3YCROZvvfy4CHC1rI4osNuNI4XPSqcaiTR3Wd1dNlUhze5fYRxi6UQjn
e+FzS+TtSSBnIRtnseXhjI1+turAo9D0V+8vtb74Bgkcth9oloXV0k+oQZDVmwXP
x+qM7tb2i9u24cHXGjdKzeIZdQw+LzWjKox8p8miAlgWihFhs7y9F18U90ihdvmQ
SiWf82QwzJrePnZUMvyJ9/XZPJ6tLd6eDaIXblVlNhusmisRLHk+t125c+IkVVu/
P/JxprUtvrO2Pc919LTxEhW4xcG9yvfGQjIyZhYUXGJYGTtSa9puuCiSPu3mFlPK
gg20k2QWyZuaUUxuUh4xgzZ1Excli2zOcgE5EkMKJ+oiZdJlpHkfc+lj16t8IwyF
obyUQBunWDpEAHy40HvJG23cAikyBaQTh8q9JVc/IlhYmpweS+P3mA8R/oprwYNU
S4WzNgSdeClY9FHpq0dXfew0akkEwsOO0RP1+RQ+B7LN6xriRpynKCy/hHV56Ef1
Ia00AN94kayHhWjfaqUB+H+jEOzYGDzUSENCYGGH4RTbhST1BmrvPcgL/CyGK5+I
c+cMAxlOv+jR11rvou+73XAUJn2OqCawugestWvJHdF+vHzwS/11bn8YTu0+GETL
tIKyTKLr5zUdHeb+iRqA86dmBhXUJ09moskh6hEZCk3ggYZiyfOSYbbZhTr1Oz80
vbui6k3TG/5zVBa8CPTIyrcCIlRTo0g5p9X5vbcjieifiGyxI4VawIbh/GXW1/h6
NOCTMMy92Mlv95Ei7OhWBBUN3AjANlCU86IAngv75mMjg+3qwpOeOW/lbVgJW49n
p0kJiVy/wLMdIxGrf/CP5rXVLxlmev0djkmNRJzvPKtSM5J8tb7n2vvDbSTj0xMp
WBIsqMvMb+LSPQ5gnHXqyrYUBp3Yuep+NLJTTNQzdX5Nwdhp5EJwjD048IGEgTjU
enMJJKDyPJ+FCC+JVTjHd9NEsqr2dIazLkz1cVVRfZ5h0t2KbRAXpZYctnsQwVN4
k0RiLu3vUPfWD8vXYS/kPNMP/nU4D7Uf/I/pBZuHJ1qwZK7COSUjHq3PtmBbtNY2
771hCaOt7en6xwA5YgWWy1Xx+JyXCfOUui6wbqW3xVObdfVeBc6WrXLrZJ2uL17s
dnxN9NpOAD6FkQrOrvuY2gTbR4s71YHWDXWBMQqUzRvG+7Wz/VdsBkya6CWi/bf4
hP5rxkoJ+2wWQ1bKB3SYvbp5R+PQJcAo4gAaO66seOcUFyMyFMVOPP6pBFCJt7u+
FxYasO5Zwb3OGzTUhme3TX3rVHtbZkh9el5xqPtUNK1dyvld1uMfo3hpyqesgpRc
c2JZ66wGE1xbgqkxr98VpikwaqB5cud6RY6Re8X08V2Sv+UHYG/B8FEMcTO9FG6J
FJPX7lHw9mCLgHNqYt+/rytBVOot8sRkjUz+dY9Kx8JlXGVhjBtrNJi90cxWQKN8
LTjyql8xb2ynifnw8Fis/XKL73IP+DEdANLP1FGT1iMZWkRQAXqJmOTz98mC3Ixa
a8a2snR0GNjntJgqqoIwvIR9uuKhpByi/wRvPNm2qUguZHXsW3ZLhtz6+Vle83Wf
u2lQvs3fF6jXjO1BC1pfcR5EovdzgUAP03/9bMRh5lN/Nhy3hkouE7cOZlCYd6Zn
6GrYUpYEYBAeuw1CFjnguTCkukwYNJq1BV6NJV/Pavx0zhn/WCtm0EC58QXhNUvU
qIjtPtK8B2Rw7s7w9OOvgByYBJs2QHvGzRMedPBzoP57GL8yHP7pLYphBCc0obBG
PZOIABhAccPGMB4XHQVag1WbYrFyYM5P6lJcajT7CC5kS5d+dwjfE10reZZmap6B
rDLKFYaM4/XMys2Sd7JT7BNxMhoc0/rjj5Dc4X6Dpr9Achp27TgHu9Kr8mYnTAh2
plvGBJxbmD9oUTsyN5L0KP3J1AcRCopcyDJapqXiWw5fe/a4n8leNtqNcIYdwXc+
2DFfD8Y3WAH+kCvUDMb55cH/ETmenxxj4az04TLDK14KGne4n0jjI74UI49D7xSw
rD1DqvGo8GYnbExALyeeO7HTykumm8zDJEqwnj1Faum5W9YS4tyX0Y3N43LvJrb9
CN44h2/N56/NlCtmUM3DX6svb8CeN9aAzwUDTIkumUPKSJTuRpcYtSsaqkoMS3TP
8s85dR7s+ju8MyDPuMtFnHljYNOog7u3LJu67PDfomGzHiQ9HQuZNXSdaXgo0mCo
+Tq5T0JSG4KqdoZp9dqG3KEL7LuGgO0ydPpyOifo5ePpwpu8vznqrkmq1afmTxU0
sCaJJkLDoF3DB0TWNulZsRiPPl6YCX9kUnNMbGKEvw5ZT8zfI8elM5NEnbNLiz1r
3pqmRIJx+5pogSebX9SdIG/9+eiNaJYJMxGaBTljFrnQ10PEp4LZccSN94/wuQf5
zaxP+0zwcZG/kx0QFdyNcFciqVDBdnur6nid1c8/MfF3850NOLHJM1Oi6CFpuX/z
zPJAQ6i/1Q8PF4ZiY+Z6cjt2gvXO8gk2m/PGyoPBP82RKil5xjt2lo2Rp3r0vCIp
493AAngwWYS7o6YMTmdRp3ebscZqaQcL8qBFWePA6AlFrqn50I2WP3CSsdT/GoCt
ubAjS2+WWsddutC06StLd7gll36ewECpurEkL+GEAQrlXXUMS2d4ljDogbIVGWTo
3ff19hzM61CifcdfIp/jJTp3vBHyZX0TR5iqdIQhCrw9LZZyXovgj4Q+4xC9z4tx
HV2WZnOz/0SjGNQCduUrTB8ksK5D7ay89ZeR0Suxds0qWcQLHXxBOgWPRJUU1HV4
7gxeBP/UjJhpBTsbOSwbqIwKx7xyN1CcaNtvae2pg2K2bh9qobGUfC+rV0WOm0/s
CNb7oA5b6qXkmUOWctOPbak5VY2v+5z5SoP7oOG0F51xmmxbhG42EQ/R0xTL1ms7
ONikJB71llMoqNQtLcLv9CJqOYvPds37QOeY5B2Cg0xfpssZJ5dxsvlA/U0MiBT0
wSLdgOebs67NnRh5xCAprHYChZT3j96QhYjGsC1ZfKSzwg8+2EG+chzd2Z8ge8tf
gUHbcyD+ydOCf7QtcUPEUHUABUKOOYlvmIOt8eFgQQRAfjUuN0vlys8hXlc9fSLg
DULNZybhZ6LU117G+udtKmt8gCz22A3CXebOCypkDI/cXJRjZk+5/d1IpX2H/Ps2
Eu4M6wiNc3Fpuyb5GdM3zi85xWXbKSzJ5uJWBNo0faiu1N/W2u10rhy5QLMmts8b
tmB0EyV7qtKS/EaA4wTBMyrIWNLRB9MxTAEbP5rtSwv2nUU5SL9k84nACyJ3qR/P
5crxoVryBx9HFEFnbYmaaQEIzNqH0V0US+m2sNA9yWmn2rPxn2taWjVhnAhE7eR7
1qLBiAWej51XxXuTdd4Nm7aU1HC6+ND7eebUbTGUY8SKbR/G9sKidJiLfERM2G7s
tyGuvq6FU3fOLKImQ6b1+QyTP/2ywMM90mrVR9yYl+sZOknBryq64mXEF9NJxgbw
9MwfjoTHiIC4CDmD2ibXq8DaVkLTHjCSA0f8/L2NfzT8UfLEK59AYjsJjbIu+b/P
q1pK47Hm4Ag3C86cCZDoRrN/W5Ed9/2L/+XT1c6592RMf8rtbuCN9XTgQKD3r8s1
gvVzgoRlt4LLVVl5L6TlRzdzqbruLN7k9JSP2SUKJPlRLzZJ8F7Xo8MXUtzNi8N0
QsWzN50e0cN0wi9M5TnAiYTJKfJ3lA4vWrXJ/vT2svP3MUgEHHAHPoVM8Kif2vTw
wIkS+uQuYGja8EWhqsjyvKLKYN4TrP1LPQDCEm0mvQdTULShJCKBYEePoGi4kNRv
QRxYcp4Huio6sL+Z0YKbZGPPZKDW3I7iyTvL5AXgNG7BGX67IQoRyAaz2p0fk9eV
XAz0dVHFHb3JQ1IYzHqetgAa7cMyx1b8ThBEpi7OLiTgGttCbfqTofv4rAORWkrA
9KSDXCM9yp7m+sJC59vEVCE5Nb7Yh+sttA2CkoHc91S2Ii+jHMKNqmPrcf1KS/nh
8PNqUh2dwglYvC37ICuxQltybt47c7MiDcEA+itRsX1go827AcjayYPgE9afLAez
czVly8+LttY0A3ZNx7kfxf+v6HGjAKoPUNvFdhVuqwLUQHEapk2yjjS0/ppM0hCf
KEmfZkGOE2NXK1maSkUVxFBMler97MIHpyxtHildEK97sDhrNmuTntsNDNtN53hx
azNSloviDZqYKU6V18//2GRa9cOcby7s6TNaNQbQWedkwA9aG1XbvBdysI3E22D5
vM+MdK6PJtwcdkv1AXeY6GD+qbDUlu9cNQ9qZTkE2VH5whwZ5SNkHoSZyPHxAUZZ
ZbFfPmJj34k+9sv9vxzN3FtTbnZTZwdTuojnx5iAzkRWq8m/V9SuspuEfKj9rYPf
jpitwIuQA66NG1lssX6cUGOx6KScO/xPZRgihkmXwZsIyRuLvAmnQsbzFMKdQ+zQ
UOBi10o9fQp4qWgDpkwFeUinI0WZE6mMpJvXYFhtLmd6P/qQbD6k/d6T4azRCDjI
TZo7Ozcv9MGmWlRvzi4mAWD1r1FyhDXOsSTEYSa+Iywj5NL7VDVzYomhXKUJ9AzU
9mTtDydDGi0xgjvtl0JBlN6SUgn3hWJwfzavV0qaybet9yudKdH+/ehjnxz6I2wB
6teOZQfbCmhSrjtkq4pytCBdO6IL+r6ABvroSEeLY9N8j4qyQom7k6n2i6eHwxx9
NlalNVRCrJX/fo1IoZ2cKhHwX8wWWjvji/H5IEX2WCSDTCQ2kyBsFK8sYENIRC4H
NmjvilMzFIbCSGTMRwYWqnA9EM+Tz3zL3MxJSLWfrs3rDjy0IC6gYiThO77vpuKb
x/kfPhPKi6brBq5C7y5c2MeUoHDnEHXcag+zyCsqlQH78Jstt9Apr37fOwe2mGQe
HHbPJUEBcguWoo59gjtNqIYyG9glUR+0VkA1NKaMmQiSnmQ7DezZ3vyqWgZKWRVs
bqph0+DWV7IXqhqGYbkTVJvg415z5ls6BzVJc3fUvpQwLG2veob5jDHI/PvM/8xS
FXJRIhL1KnduPV8nLRDGU1ZJQggSeLNp0grAOo36j7XaXGX4jTtq+E7pTlvWrK5A
oIhat/QLqxp+XYGq4rjIG06V2ujzEOpYKuOdspuSzjADawtL8+VGX5RfJYRGuCti
iMzaQNk80bkqeYJPr+Gp+5ufLlP1SPpIGmLvWmVy9GCsp+fYQYcumGtWOAVPHrY1
Ot2KfdSqnul2u2YxW7J52JEEIPfzaH4mvf77ZReFgSs4jm3GD7hDLm5dClsHpQzM
cE2csck/QAVtwuJK/z+pREAqLWmfWLBTMBVjMyxrNq7acx9BZvIMhXQzb3MNTR5j
AG4kn3X0ZgkgpJd4uL0as+4SnUijEVJ5thi9PE9rVVyX6Y6EMIJPblJBPoujZX0L
b0ILbUT8Xo4HAxHkjTgf8tNBYslvoSgi2F2CugMX5F7B7I0Q9fNyBqcUuKWfMjhs
6eANr0v9F089hcsaJrm6JBZrloEes+SWAnmUr2KoVyXbZE/nBRbzW5fWU5ijpV+W
b1VYJE5ZFcyWP4jaASlkhi1WjJJBfRZeL0uSCfNeQJHa3qUm2NcQh4OLqSWrgeYn
nUqtFbfRZir2wnf+FmnXYWSfzc6vKs2N5FHKeX6EsM+FKGZrTdXrwkNAQ1V+j/Ha
Pg8jkB7PQe1CdixihKTn78gCFuFp6pz1nhHQzNGKo6KrG84ZOEwme8j23qABmluk
dW5fLWtdlvWnoaqBgKHaVBPk/8dkyWvA+jPu7eZ30YyLO5msG3TvJVVuEUacNcMn
c/rzuVA4edwtwGEDNSjJdfNzmos1Ya5h5qM5FfS7ccSKxiDS5A1YhygnLNxILpw7
eaNRB/Qv1NvPOB0RGnJg5hjJc86DzfVI3JXzhoBRajkO0rwPhwG1HTc4ZhNIkJMQ
rDQ5pSxTCLeGDiNO5kQ7LoAu0iiCoO7dC/Copjn8Iw+xet3yD2kWH/zwEuNm8wl5
veb8HFEaRSsCZ/Ixd8JVvNyMQBy7u4B64sb8DFyMFMbSs8bgKxqcqP05Vc/gyXtV
lhAIfV2wycY6XstV+z/k826AKYv1bRuw8kYoL8tDM/4FViTGmrlrPQ5/+Ra64jCm
KapszV4PJy81fGX+eqjq1hJMAuTNSyXcUyxjqgNAdJmtlRaiXO0iu4COsx8sl2Kw
dCZUMN94eeuk5mVtlTCyXNB/HFJds7BzNIoXaWB6Loez7CrSBsNuJWfHnLs3T0ic
aC3K+jLS/oZB8IxTkO+fWBZxFVtPUc0XYPrZcbuNYpZ/DhdTNmC1O9cGayxlLQuh
R08ee6N8Cp88q4OLrFp1R91kA++axo81pEoLBVaiJ5Aufd1f3shY+Dfi96W4uYfp
BzXG0zaBsGa4Rd5yWZ1h58w2EgVt9QESQVMspAiiES6FEs5yq0x/WV6+alwSD+ZK
TVIOAobcQmYV8poFBvD7vzZf40D1Los2SrKFLBinJmrQc8GhiicORoI34o84mEge
WljoFb7YtZZoOvrKGTkD5H9n58u8cCNBe6ySR+HsjLUrsxdMC3XllNliLEnMZROb
h2iXGWjagrYRjxBe0+9cpYKWjqK0g5zza6sH80thTVYqYHMk2XT92Y5vkwy4VbYe
VRbslgvXq50HiOQTG7qI2TjOm0WGhUqoinkExtvd0FVAGEhZ3OUl+cSKofu25oK+
bhFz9J+zg2guz9wRuMvPncypcMU6gqdSfCF61vLlvJV36bulLMMgk4fgaiZn7AQ1
jEMC6Drxq+l3T24Cq/aH7Twt+7547WdvBO6oT2X527jvRTh6Qw2g7e6CLFgda6dd
1VSlRpNFIJ5zsY6gQFtVy8CKXkZu8uRfqm2BdICT947z2NrH+P1SyaWHlMGCKLfQ
Wei976SwPUonutgE+USWhvqFuRcoOE5OSHcO+pdVnNCguIwnUE9ompL3np8HobvZ
4ABXzAUDWHX31IZv/ZWNoG7IxmR06ymYqAyVJ0Ry41Hn2G5Tbsqi2ENDEPZAW4Yl
xuuVgzHuzTFDe/POgeVnV6LbogfM2ew6JJNWV0NAmH/1so7Q/jOuYZTiH4kTRlyP
CdtRjw6zvmLzWAvSfo0FiC8blrq/NL0mlKMxTcWhh9hOMh8DrzQoip0nuvq5UjvT
u/CM5xhugzQruA2AXUmmn2HP90NhrDP0iJArYcnFd7e87hwZIAfkduhzyZXvIAnv
UDDgwLS7qG5S+jqhiBgBgreZx27NkZqnK0tUgEdPaGPMkm/BQIhkfupqEI3cEKll
5m7S82lDu5P46nup7svhbQ11E1euS6/GhHHjZKzBCn7zdN3JMYFuRghmJGT7Psei
qnYM4cWUL4bFiZZN2FXtRAJCz4MfmcFn5Pn+1xGLdxrD9jHzhPCUZksPwlB4zXGk
4s/afrNhZwcvhVQtlP1/OY0cFB4v5b2RcCj8h5U+FMQCTorODzKiZhf6m70YW7hf
1yHglmuyx+99/N1KL1NzVffTvcEwVDHCkQO+q3zDDoHWc8Ia0eCMH7vmq/bJLauV
wlYoiZ0d0E0hP3HBORB3DNld7/tF70rlQ21/yv+cpl2mGTAM9IiBsVSopCJNXzVC
wElWiqOm7O4MnsYP9C396DaTqdlrAfdOBftONiUlKwQ86wiuEOf+31us+XgMq9jZ
qOGt1XxFu/iDMhkDotHl7eu1K6S84c/4gGywIaT4h9StKN1Lkt+3OFOVrLHvLZxJ
7Tk9Hft1CxxapcdluO1c2xIcQHJdPjWwE6mdabD/1OKe5qeZlQWBbtw6xmuSL3TC
4akRSuBX7WlWs5Wgp2xe7bFX5ZzvNucBELEIazfpZVMLhlGk5dZYW1lkLTlvW0aj
hd71xiQmovA2nK228YwGYwa3YYL5z9+fsgQ55pZMjJQhCuotgcc67m/Trzlya17V
pcaDLrfEaXRuyHbMfLSXB0C7pFkA4ZBFf2DWD0Amzj1wc8GHclRkNpBsY2f9aog4
N79vBGpAckcSNvPqu0wU0DbjclAl5UdenH2Otw/SiPK1yIibs0IAm0GjBWHSWHgp
tUBZ2/4MlAgwdtJsoUaOpYJnSaTkxd2WZn2Xl2tqyQejxkMJAmKTriS2gC4zeXp9
OF8YtFapVrWcGF7YALav8IQivJoN25DObViGS4vf5haynoWgFkHXW4/mBjLul5hH
IlA7w22whrVGMd+UJyohJdnWwFUXdzjj0oKK0uNEaotW64xPrjwOfUBM6NZcrkaa
pBMCdIUjCXZjfSxjbbqaQCeyex3DthdE7rYXFwmQ2Fh/5SWJ59ujhnytWTxbVNOD
7QWar+K/gbzmHKViVKYgV+4vPpidKaNI1/FWHDLNn6OjBETLsysepx+T+48kSDVU
sEyIlN1sybD2mC7JW618k8ShNH9UVWYVdcCjTsSTWJTTFQU8thdK2cjZWvaAF7ca
eIa6jwtFQTHLOh0JTM+3BU9/vdcurK5fYGArBC3ccpFHZkcUv0xMNDN/Ff1qTqcA
AlWRoBhA6vU1+ixSJlDi+Mvhb3pyt4PMek9u8/9GWZEEzUkiyYk3MprO4dZfom9v
hNiB1G27gOzO01dtKdkPUeqXMetVqx0uwXt2PPBIoxYdCbcufFoEObkij1vFxdKc
YSxe6mbB10m0H8hYlyQZc9tZ5jxPpbyn6nVcCqwIqGx65MGb5kXxLT1WhTHyraek
Vr8Jt3JYIvjKy3ae2GVZlgtnv2nho4ON5StHntr1pwMKO7F8RjoYYcZENf3e5d1N
34xIl7pwN7yd0JGMbgqhzKhVUGeaiWs9EMo+CQ2f8JysXgYotC+JlshOgau2A/IB
Ad7vrtirnO/hXAwUowX0pSLCHymWau0RX7JuI0BR/dx5YNbfj2ZO1TMuRMsHfa/8
2uBhNnYS4j6/KSNBu+fxmRYqEf+XgRBx2wNYZlKt+oLgP2p7ifRoh1uBMiZU+f2J
c46/90GWM8HyOWECAFlDE0ihGkH29KKIaw8Ce/j8xg2gCVBEc1yd9ULbxWQ5PrNn
DgcX7SC/S9jn0/Ix6wrlRWDZk+BdXT0CabMigDNARGN4HanUoTPB3H9q/154LpgF
vgafQBwWMFjyqb8fgqMo+5WBUQHCpHL4GZ81kArcSUau46mkZTCprjQvQsZNNYH5
W2jmM+4+Mr8J6vwgstxPWDkfzofUdqxzhdIK+/sCvsMZ80hlfYrEPYnpyoRWLhTc
BRTojAVwHMmNuLvjNPvpttGB71X6i6EyXlPNUCtWmPEv/N604bua+axkjx20fAhc
Pqx0i0hBzT37PPwdL9ZTOdC6fahZYR7w/CA7uAbq7/dkoj2TG4SBAbUZTFh1QXwE
uUx+w1fGVTUygWSl3Cf0D960vfeEnC0tNr6CfJAOMwXuvA4j+e55q2P8I/7fNWyN
1OKIEqv7CmcmaP6558wEhb1XnFjFuhHyUUF/HYjqy14L15w3UaT5rdo0kaoL1979
omxtai1SVTaE3iWwwEcU1FuUyHrClCJpKScgZP26HCV8zroXDYA4EuQ+7QMdO8cV
F0sLlp2hGDWY/BmTaIs7BbiSWSI77qDJ+ABx9qcFPNS/gxF/Al84R+mNu0skWwn3
Val7SFjTuYjU5BlKZng46GykpjLMUQ45QXAdoCwV+gPBPCgaz3+2OL6wILmQvzDx
A4ZkuFSXF0oxA/7xElsgnLTvsgUHc7BLjW00cbC0aD4WAtyne9bt3oAtODaw8fmp
X6X43qpyReauq3a2SFQYzgWak3eYRIGULe6jF+R6RlkIdMwE1mIRE1v335FSlWRc
5k+ck8ursYbXJEm3SrQ0K+x6th/EdRF9PoS6Y8eBCWu76BvSA5nktxkcfHr5omBL
3PDobGO2ywWFEZHJwQZsi/m8sXVG+cWc+zNGCY3qDEz+oHbN5Jbu1mLYRgxwiG29
i6FjpN8H+XjMEFD5RmWoWHiP8HcW1jRrCQ5/+Yh//MXdz9INc8y7feoLPprNWYKv
fIiSfI5ASNw+caZUUqOyKmXhwCwAZLkdiuBFxx21MKfNRSdpMzDqLB9ShYicRLjl
LdrGZHDEdCeSn9cZ8ZxA0TxBnjIT53cDFj3Jd48xlRLfTngiP8Kq1+5mMm0AqIDN
WjFN+wcpXTxwNvF6TmhCWHfOYQXwoMpz1zEKH7P/FaRMeInFdxCiZOuXuvUNFPVH
vXHJviAWWY7Z+TDb5Rb031IBDZYX/GPmlFuCZ/dn9FZJv4DaEcKVIaA5W/tejHR/
E+E682SuZadALabEd1RnO5XZkjWtNRu619Kla3xHpLM2XN8npKolLmcoAG8zpuJq
4U7vscB1W4ohFE1xiSAadZWWI2VzkSqMYP/UrPD081n+wFbDhtRRUSMMPPH+jkeK
KRyomm6nuqxEiXLXrR/KASJzeJscPSwWoEJa+/3jbnvJZiAh0L7TfMKUsASwE/80
f7hYNhTgQxuNSwf3K8Yh0ie0qGqX2cciMpCJ9kCUEo4d2wsYTy5Wlk0SibAko1Xg
FCvLV3AntuPEHd1asdGBtrQX5aIrRimTl6y1NkpqJruzfK7vjeUUE8SD8ajuhGat
76KFvbc3ydMwmKk4OQEsYKtF+1gx5/2PMQBVxyyoUUhbRIseVvKjFMCLgCsgTj5/
wyD4HCDgFp2asSWxKjfE7DoPBKa/weeCUheq4TS9u17QypRLGcTPByXYUDx5U6if
WIJ6dFw+k84Kqi1EOyTHRvs8REElrvOjJ40zW3xCZHqaCdrezxjR7bgdfL3vJ/84
0rNPEkiHDFLk8ZEtEtN6iZpbFeqOxpM3w8RT7OaqQ4hT+2XVE3sc5TiVkpvvFQeJ
jueHXATqqJuKra5Q80WLNJQ7RFv+gutF2UffhZ2YWanPhB9TE1ergoH6h64MRGxm
oJZv+rUQs6h6pEJSliWgGLdcrLzwdAPvvSo5dvcPlNZKwLmEWxJOTBEDaczhpF9k
brfHxQrT5e83b8qmf09Lg7wAAcFgeQB5oJqqIgibvf6D20CFR5Gn4zeckZkrLb0N
PB1ccjIadFWahs8LPCD8OK+x/zKweFCe7loToxggwlXQUE0QICgHxNjN0Z/W9I5u
ljC9FWeKmA03TrROQ9kIror8GA5SbvdPu/nz3rFtI3J1tWRmU02C3KMap/f6Has6
LjL17biWj7PSaHMxmpv7tGa7cM5tQoRMZqQp2zFUILPBDj+DHg2DdWQmKnf4kyXq
+uoyr13CPhnW+khLvTT0l7Q8qIgIgMe0LVphDJt+Pg76R+cBXs8fecYQiufgStYx
xBCyXllYVIDjLdftVRPGtsuBAAGuSAdtBkltxoGjJnyAJWbLvlqIH9RKvDHRsNE6
O780MBanNfOVVBXYx/NhGOlKioJWpqnEMfmEcSUCgEaSqoHzF5IF6EgOcXuz8cNo
g6az3z9P5OLN7MY4XRRlx0IU9OCdaZGHL1Z1b35FyBt8nndreAmhP8mLdVIrMOR5
BscdlAFHWyyolE2OaHTIJ7XzA50vlEu2QEvl+LJ/IAkEogz3vl6DgkmEiqrRSZeY
xNXDCBbJevH+w4mNxh3BW8SMngljKN46KTt0z4xXQgdDA1ZkJTMsQULDyyJVOsKW
GjyK9sYU5O+AMP9AQ1EZfuBa72j6kVydpDJKDJzer3LRn1QZSWu40Yy4oRBtQ38P
lB/d0Rt0IlJ/q1qvwrp+XytN0lOuqS/aGJ2vgP0gagzWzAcTFMI8R6AWNVrwa5Oc
H8GPJhgQ0OL3m2/8tlAYtw0N9ozMXSM7hqVP265DOnnI6Xr1z419qoOqEUf0EgJl
V2uhz1UPyxO18kv1/A1TfH+YL3Aq1a8ti/u6lqsmuLj65Ei9Dl9v1QBqAMN18aXC
9Q1Zw+mH/lRwx2HDXAt6w+tE85NaoAJklALz+CKnD5b4n1dhbnbsFfjQHQ0Muv6M
e4GU/psWLzgfGY03I4flVSUUG/kvPcRCrGa6cyzPlfuw6YhvztdlCTbWo4opK8YE
LkQmm9vpPNHWNCdK8dPugW4MBthMuG77W1EEnz3INrunzQgf+F6dr4RMcFu0FTbM
Gs8VyS4kWKVSZEqQOca2FSZhKz5p4wGYqr9+bI4vtQGajRV6z144m9dGEEBVLvr4
S7t/Pj8zExooZki1RRdicdFPVaWBsT/wP1vbN1E3s/78IL/1oo3kO1Md/BpAlIGN
VMo31FoOgkJ8WY75d92OK5ytGQL5XoT30y9CV+1a9yc9sOj6CNigcG+BlxqnDyw+
rNpZclTp5Lhop1Pw5GXzsVekU5nzzMn59pmcpz5Y7auN7Yx43RgJMcyhrKP3L5Gf
z6Y4LM8cPv07fAsZ1/nyC7Cozjv1XrC4E3djTE4Pv21CoUKBBRwXUUncpdISe91k
7egcFPGOJ0Fa8nAbEHZerUiXQ2EK54EOjyLIqRZWv4YC6/RZjxgswQ3y19v6Z8K1
zu2delRSBMBtlTSpQpFs7P26gJlf1+MGonT7V0eag0MAE2JaEYkLEEuZb1GnT+rl
l++w//R6kvSJjYHiE7T5DtS0hYzLJSYmjE7E/vcFxGg29TzqY1YeajEcVZ1ftKXU
jM+Vyq9agMubtaa21qj8rpCUQ/w65bS+anpBy3d9CIAGHje6OI0vWjyWurUkT/wz
F7AgBfel5d0gOG3Dm10tTpa7lbbPtYCmoxvOvOiUOYyy37kv47vsAhxA2hX0DrAJ
htstJnqwN2O7Az+OyZfLg3IMKr7CprLBRa/uoEDQoQ7LWF/7ZRP/fXDg7Orqq/Bc
riItD95za0yFFP7att9a4yNoo2o5eos3iuiel+H7BpF1tG8S1PSsli1OPDKN0Qu0
3GfOoVn5YmriBFJ32gr0tZ3Ac6HBOA/AzWiSuu4tE766AdXtp8VY/CklZI3zGlSb
2PSBmVST9qdIsCk1cd5fIQdEMxmLujZkQ+OPlv4OQAN3BWE+Q1mBeZVoSoOtQ42z
+94i0CkKnqIbvskAh82bMczoBH87H4gZ2MOAVZAt2noUpJQ7/AulWxHuEQy66/Ou
zlVwTp+0QmE+ueqepDCDOtLgrxAxYiWpcMChHTxJy3oS61caxVgghrBfs72GVNS7
2I/s0J/5xYZWrcGxzBSk/nCgo+eQXPRPEF/qm87LvWoYrhAIyzWMRmY2KFRQrQr8
hMD5iIHlrLlrvxtXof5P2AGDYNSCJ1gNRIz1oDUwbZb0Fqrg0b95pgSnKInshQpU
XL2YOzJQiK5yXM6CRc4uByH2siZ2W9OhPfSw+QPJqb5/fEoZe0Mh47yXVCpAn6Nq
WspERXdjBAV4l7lh0HVRrW3yWUqgjj/TPzeHcCSSZJ7NZB7z7WFEf1W/6Z5KT5G8
nNMWY8MlZm4crb7/ya5SoQWo45SnpO9vTy+titzNTur7ARq8G3t4ibYyw0mQBJar
ZxIrbTXxdpRWBtyTmpsEEAYsWjRG580wTaw+xtWYqdoz/6ZL8V5z3hqnnOwiJpXR
Aw+CtrJ8vm85oELFpHR0/rxfl/2uEkg8e/WCU2xs5qqKuaDTLxmBcfhLcSLSqVv6
qxox2H4bNTZLZlmvZByytwReaZWxyulDhGfNpCXTX6HBrYpjEacP+WYwkbvgLlhP
6H2ymGgsJ8mbIwO19/Rfuu/7N27cbwiWL1K4tsrYzUqgcOj//r7d1B0mmjN1uYfy
1VQdLWUE+h/iT//uvLzd0vhUHU5I/W3GFxIVvJQsjMf9MSytYvPCp5qYNbCVS6mQ
D16xeeJUh1JX6ORe/3NkKrzYsfVz4v6IVA+pSgQaBrd+V+sGX4zbUz1aNioohxwE
H8XmlH3FFcdyU782b9TFq7zNESWN4m+vUhrPwedPSHbv+oUHlDxoHDwTTyjk+WfD
ktYQv7TF4/LDMlvHqbbQRmQjOkoRipsWxOZKNs2sNWzllWiADM7UjiztIFO5bOBl
GBL3RcQ5jU3zwiUD75z7os8azlE3pPrDSnAiK9KHFjv3dvUpjqM8BYJEIDt6TPp7
5hhm/fhmbL07GJENhqUideEfjMyM4wPHGKL8fAz04Fg1jur4vd4TItdNY8FItoSk
tvLXR4x1FaQ+VfWWmZmRaME7pLv1tif/ypTabaGQn1tFLe2Ag2qHwZJWPyOwipI1
wOO43B+czpUXfJGNJ+exLwM5CTjEUEim3JbvnZZGyRLPHhY+uFYBbgoOMXRDNMza
xHy5sdJh14H0Rmm6Y2Lk64M5WeBXQfO5h/A6sBeFVeAP5r3wPjMJHMTTAvMV+i+X
dJtbQwubWuq7n7/q/Hu4LkaDc9LY2s9a8j7AFxn6cK/xKMNpLISo14a+sl6bPj2w
b7wnHQN5pxetOfkGRnGLhIgLFCw64vHu20NJuGEIhISpxVbWsIzn31qMt2WrvwLh
MRfsnJn0FvxI6T4GG9kdJXUJKIL3r/x9i60VRDHFbFxdF4lIJMM159D/SAh9PRk3
CubogaEPU1RxBz/1u8yiniZl5OiWZAg+IAB/nvfp1smypoa0kzh9DUYonLmE9GRP
LtdTMFufB9iDabJr3gm5fhiiPcb1eQEZ74Lu1QRBaDXGOcwAyMRfmsgZyW1L5aHl
/YFT+7ivezoyB0doKmE3k1XTYvyxyxFgdT63Tkz2yL221Sb0IrJ9eZSUW/QUqwe8
AQpBwucsMqrvZrKgto1cdiuzbUnbEV80SkhjpzKgZ7AO0bJ4rpmp4dwa08TC/lO6
hBhlBVx/HmD02o27Lm7WHxnpdEm+e4N1FizHpPcZ7FTXsrunvaSzx+Nnnl2IjVWb
9nmbKlFmZFSRbSjdnKj39Jh/7P4z8wc+RZC+SuOSkHmJ8Y3K2qJukl76Zic2bYN8
q9HncdWpUO+dDGdudwyqoEnWefL+r//imqY5JB/NuI2OVmQmzWqGvqizJraR8Iif
P54/yLzXgiuRekH+8WaDQhpOydcjJfmmhwpto/VPd3TJjzqBf5AM27465E9OT2lG
j6Uxl2IzlkRlUnIE1JimwPo2s3Y/BsOAa2VQSezLbwge2zkioBHUNvGztGsw16Bp
u3bMBPmpZt0JJjDqQ605CggjicYC8uEOHXBT1jH5dWWyHAVS5YRpBfZLEz9lMfa/
AEFR2qXO+yAnQh68uKeQmI+kT7C9F98zJZIxsTrb7kohTeUV65lad48cLVstf8MR
0K2SxvcG0KpxI35/cycc6jKSV0kGX6ztKrumZW1Ci6jO5R5aL//EcX+YWenPLQq3
xFpOCMbQUB1k1B4Z36yJn5MzgpMNwiAiHwZgwHTCo2L3SuUFl+qtiZEWnzdKffgb
XaJPCki1obuFSxmZmk96RLzM9Ild/F7Uy2hEHZAFW/IglCoWAJetofeL/0/GQTXG
ZprZVQskkYKeQuW6rUG0mA8qxNcfKOd0s4HP62I+SDezfMqaylICJWGmPvaFrYjw
qp9Tt7uvZRqVRj2j1vyBk21m/O4+jUQKjnc8izoB5c/H8TiKyBPbeTY56+LucFjN
INSNmiX/xf9miciEDJ2yCFT96QZk4XuHmlPIO9O8ue4Z8nDAyqQTo+4U4WOsXQOe
V0fBy3CpS1oojU2QtzbbZhGfOEzI7DX3gms9eXnvprkafASU4dljnX7zWqBqxyJw
+ytA+O6nxaLfiH9DHWcexFDwdFezurapVi4MSd3iTxFYoC6r0N5Ja+50Bna00VB/
h5mZ6aNng6ymFkn2edPE72NwzfV7CDMknf8Iu6hzBTOxRZv5yeFmlQ+bkWYPpoqS
s/RKlo5QzHUf74ijVS3eIUv1aRxXZqcHl5iQkwcwChn8a1Cz9QMKU99/x0OzaVR6
TwEC/xP46sM3UlYlepBsARF/LnYKPGTcyxjcH+cKoBmxUsRkyg4QIRZTxOcAQLtd
GViOQ4HgkSu9E8dBLGyoFkJROJQ/hTa53RadjWYupEOLh6BgzziHtPSPdp4xKF60
BkY07oiWOG1vfX+R5+Uze0Skd0+Eowc2SGxDykdrUQJk89FG/ajP/1F9A5WFFffU
9qbYbec17GPFeeKcgqzvz93SrOkDalYM8gy5W0xdwYsTK+V2rDCfoEq5Khw2k5nr
WL2HnsQsIgrCd8ZImcbE/DVQZx763xGBI8nHBLypy3mJENV7uWmFJogeTqXdPt3S
BYUuDuHyQxwcqA3V4AXvBky+Hn56bKKC2c0cwjbnIYMluuxzrnjCd8i8PS2bkoxC
nQeLYRJKzEg+Oeuws+EcRDViN4IkQo+scymmh2GIRuxjqgXWhyW+8W7ZNV0fJhAI
+H8yl+gCs0d9wVkRCfgxFtIdX3gaZ3j6wVN7RByW1pKVSwAs1PDUPhqOTuEy0DFS
WQ+O8OGz+ZkuxAGlTNY9e4o04+fJFo3R5YVMWWsXDh2VGTGUZt2vi91fpPDHI1k5
n0Dtyc9Z7H3caIN9Zz016Jli1xeCuzSdaDsrAhutzvbXaVhu4hwkRyCEwMGUSuCt
ZUmWNXyt9zduLukhRIVhMb04YhLA786TAUxtP2z0w+Zil2CW/WL/NQIyeFh57dvj
0VaUoOMhvfniy8u2WqYE3l0KW3jKDvxBXsfPjHTXs53C2Fug1Q6cv2UA74zizRRI
+JQIvUghVvZkUSOmbcN18lMM3m1ajUzMKTgW7MGIWGficuyFHxFRwxvMtT3dIuag
o8GWcssUBSNZS9jA9z0H1UqeXccCjGVGRisFxW5ndUA3nYervVPbsP+rzE9CN95v
sOENxr+olgVIpjv9BFJcaPor48y+kJ3W1naj9qyfOOk3Clpwlg22cx1rj4XUUc4L
F3InqD/edHXmTDWY8jnzzCHjRxYC/NyACEJ14CHkJBZsE6eR/uETBEdIjcwYulid
aabY1ZObHeSlQ/fIGRmsX8aGl0fqejWulHzkBSt/zNgA6UYegNoPk7vj+USla+fs
bW/B2qW61tJ1QM2E3N/WgOTL83D2HVllQFyA4xoBObseCcCeXrvfTWuiEDSasaeZ
nKhdIq3Ayl0xBdK0QVcfabiw8NzUeLKOwjFQOksi2A/+s1Sta6JrMZ8hm2oF02c7
nW8nmh4BVh4OLBeGL31opYlog0oqQvALMBEo5YB9xku3XelhMlDryUwmW3okuP4A
TtBL3+KLWLS/XvqnhdG0J5mhqZe3i3a2oIn7lMchs+0cppq30vNCS4S8Igry82Cf
tiWnwPnzxkx0mURzQGSklp2H7XbSGExGHK+KWIumosvAqbF0JpjV8OWgyd0ofETr
e3civmrihdr5AWcKiuRoXYoKEE6Iey0QpGdzaZAACX255jywEG42fVTj51aWBuL4
wcJe865QyDDzpSTAnTZXWpMg0UIrPBYy//G9m1uL3P0Y2FGyd/GyraXoCm/HNYrx
RWeJLge+8E+bMNfL9/Xbb5henFlHCxtOpAo1V4/L5/GuD5BeFxA0hbPaj+vCDLzf
A0loC3rKanz9VxqyQXleaTLowlYrCT9paDgcxZf9x/IoaW1UmiCosL+kCyhcXC4l
If65VHCGXfKY5hewKGa8cxpBNgkzaGtxRC+b7wg7kuGzuYoxGRFT2T1t3Hkpyi6A
QA5qeXa2CzWXE33eivFtV7Ovo4Ne1IhEK+LJUADRJGXMj6uzkCMZNWlCJtQHGsux
9WFEEsgk4OwF1O7dkc1JEnRERCGtU0M1h4Zc2xlhUl1u8cO/gJFCHB+8jD17cyBh
Fyu3VKEJMK9q8WNANm25GEz44ZY7QsZkCgqorlj+87ghwy0dKv7yafiRBaE1OfVa
cohWfRcJPO2L6a/48wxcNHWB67yIOWNwd5w+9BIaMqp21YrqYDNiNWiMELi+B6Ix
Aps3Z7DLWWZcXPYygUX0BiVEFIZ77tA2HfkxZpP0wDg5qc3mYEn5fJfPH3vRukiY
RFsnYRbFQBGL77GBXkRuQh5KLgRP/BkU/AuHnJ+DQdQ7QxriP8SknO7Ze6F+ImNg
VHMZ68EgH+c5zVujkd7fsIGUck0IQKwSe1u01fQxmCI35qbZKjUFQqmuT6nrFWx5
V9+tK3enIeua8HZtczqnY5SNRS2D5dLQEPtFUQJ5GzKDdpKal8RuBt1gEUruPShK
ZHeLjFAxQF6B+sUnjxps/9vyEWimtTjcPDfTnZAGYFoiHlDQph7mWrQ2mMv3i5T0
a4+qbuOI92qE4V8s/GF/22f0mCGvjUF6B67qVBbf8yX85gIZwDEjDyvp3uHkC7f1
qXW97EDsEjfMZAShIs1JFmeqPfWu9sOaVKxJMnmaPMAb8ELKh8ji0oGGQ7rW7VCn
uApcqtCkF0cTSeseDDxob/VfvfRgT5/03tKcHmDCB5s6+9Z+Y3Z7vavJmA095M3p
lXqxV2VLwWOYs5ce94a4wqJYNSBPLNChn+tC8VJtRGnZTYlQ3xkbU0QmeGGm19Cr
QBhGv5v1qcrfYoxNjfinR1Bq1kpcmkj4J7TaHC8oIBJ487BTAkIxLm6LXVAzX3aR
Us4XvSRLC8WTap5cvstpSjs6QfaS7OQyrnZTz7sqWK+BlYZwtv+ZyBPJzq+LLOEh
gjlIeTY0ao28cZiBDkpsKf1HykGrKUuuIUaD6qt/UjnOTh9oNrwM9cZ/J84bv67Y
nIOCAS6uuPegb7C9wE3c2qn+4SELka80/Bj2EqgNa9ZZKVqutoQY8EdPpaiLpXtx
ipzNhQENDleHIMGegM4HMT9KHJ2hMkCMUBStkwPBVB1NmoY2nnR0fJ+NsJ5SLYva
Eq11yj3WCugpcHVGBQ0KPqNksO09w56GU2KPSVMMUZqRuMqaNWbHYUlCFIN3jIPb
QOSgdANB2eDaVcwHqI9I2w2kzOckB8xP9nGzVhEIk5EEgI06yJ0BgGo/qe0np2lC
tHXND/0LigFrEgxrY0K+7zMDfU1pdPuYbZc0muKQ5f/pWjt8fHsgXC0bvP+m1c2g
RUQOST5TGMfbI/Oo3/TKCNKaOdKyczgLka6TJ84W7O7g3Pra0akxMJG9AUUnA8yX
8Ic/F3oBc1J7iQjNnrAuSEL04FHPftivj+CSDh0KzIZHjWMs9NVufpyQ5BCSdARR
N9Xam/v8+wd9EhgaduOPntxiGGpEw5ihIAmGPtHdAFzcf0K52v/DPj+o534Ru53z
9VqnjrR4MHozl3Pfpw3AyHDcYY8Yr2O1f1KKhYQcLTzzkiRMPIPb8bMReMXdxuOG
0WLOgGSVp3DcRDoHSivtfhwK0q0hOfrWrHxsIQlhnlA8MiDH8SnrbMjTck6oYYkN
Tn2pSLxRazLpXwRijlsqNwQ8aK0XgoF7THz6H3jWmwEt4pmn/yT6safrESwFgih8
DOUzYaMM1jAfKVhTpshIuJXROaQfhqf/TDQLYTs+EHceIVmElpQ6h+v9SOXeQzrY
MXju1fSNOm3LCjfS7DKbVaVoKeVW9chCSP+IAoTifhwVZVnOmUwfANo4FChN9ytD
mSIJfnGI5mgIC/Hdv99T/KaDUoOGvw4j0pDUO/g4PyClnUMSXHQuwTKI9noJzW14
8jmj8Cm5ZIj0UHwi7DKVuMxGtGkHiG22faBOUcIgZKAXo7I6597mqavDhOH8hgq2
hHmK7pyYE68ih277qnRYGe9G56sxuSJ06TfN1Cc2/ZLWM1deZDzbW0mwJnriDwG8
PdAB14yQ+nD/par0/obU3TFg3BG/WX055MPqp9c/+gipZ9Fhht0rjG3tRojDl+gm
IDY0h3fEQXycbUeL7GQqvQ/dmTZZdy9/QaDV8IxUvW1HkgTiJxOnblicCvCSudmm
CV0IN7aKBem/JmDpcnCTv49JuQtxM1/LSPcev7YI1NOQd3dApY7ysoeUMOUZ5flF
Okl+iqWBdUIk/vmTMtvabYgs3MfZIRvpG3lQd+ir5qA+NgATC4eppHsOOOs/dO4L
7bJkofn0hd97zAAVjZaJijieAEcvS7nX7HcQGMY7Gh1DMEx4nVslHC2L7uMDNnaB
pQvqEL5EJs2Rr81noG94dNhZgdAT3UDnxan+9Njw1+4Io9d/ExqUrkg+n1vFXHq9
u0+f8mLl1aw8QiFZ8UQgKTWCSc73uKd5HWgO+QkilXogUoG2VkoWPza9kF72m31g
BBT7k0Yu1jDlcwMMAHa4rGCNJGVy4k8LAbz098e84mw+yXjM3Dh3+NDUsMqDL3Hu
hYAJZmCZwA5ge98SyOyeRM/oYb6N4aAA5y5hORA9LpZlRvDU7V08/PjWcqNBaL4J
TH+yMiA/MtBsb2V6Bkw2J9f+tkOLDN9KpY2q4xK2d62AO+o5kj+0iP7X8gaiOwfG
RpiJuooQ27FXH2FD45ro5rzity0V5u3gOGYdCxgzj1xJzBVjLxf12+6N3NgcxMzA
emMMIqdnnVuXaItjc3ACz/Md6vu5xYGWOi+mAN8AvHAZKOux8eOpx9xqqM5jQclO
NuNfz0QbR6MeQmnPNoGEX250l39yTt3DhqJJvuXVM+5kXLR5UzoATLdf86xkM09M
Cbc9pDbkyKozf3S4YTCcsHdquxhIJoi4EwNi1V5EsOeymoO7c4OEVDmJsCBPppO4
0sJ3QTNniknTG7fy1jDFXfgGdLZF93pwfxnTrhrE0hhVjjS+PZs07IChHF4Dg0pJ
eU2CzWENFt8em7mJDwlJR5HD3QoWdhBJaYElvhvoXc57YWEGIWRVnajjN3Vb/+hz
o1LI/WczURup/mfDtF07YqBehP3MdjsKUaarocMf1LjgYUMOvWD0Ky5/HH8FyMub
1RiypheQ16VEOt3O05HgbbMscWVToUEU7LQJASYgv39pz09FUOb6zaUvawJT48iv
DWTtQ1SBIx/kLe0Z0RfhX67y48YVNw1W7jBuRwDqk7tDHiQmNOd6f8oeX5Es9DT7
35TTUZ9PU+OJYoddi4ArEdtAZTfwCjObob5rnG9xl2OiHX7ZBQKByygqIBQ1nCIB
TUlJdMV/Fj3YepwaZaETVXiKHMDMrWc4YBCw9k/Ynpy3YiukX4DhvPHW8KyphaOT
Go4wtNMsW8c6H36iq9d6goJV2+qF6QYY/xQ+0hnpUoEQ7rdkoSKcrF7snfX9sVv3
cr+PRau2wGJ+eNK63HPDnHBRu4dS89GUp7lpgOqa9vQFOmJy3hzIidSIhhoT6ZPz
FDETUKeE1JcSE9xTMEzJGMHZZ50+zaTr4j39yGefsD2oP8M5k+vXc6A4qb3ckCMb
+/7QD3Vw+qTS7CzlAS5IO5Fl1Q9VYQz8UPO0AVjfo0qUVWOBJhLChgmreAx+90yZ
lYabHFLPQOIgPiwAQ7HC2FAtA7wMGdbAle1GghiOZLh54ddEwAiwaiQR/3ekJI/T
hY8ddgcf7A3pO9Vnr2/BHsevF5cyithkt1yDmSMI6WS6eOV7Rsy+O3Z356s4Rv41
49k3SJ3EIJgQYUq1pbbd7UsVfgrMUcQugHyr+Ogl7Z5uZBzPlsTkfY0SBXTdwYWm
5JB0EAkMOuaO6lSsoZeM39J96/Q0NhLCLbgEwOsVZjEVCYJrQUNJwv3Qhvtg6mKA
6W7jb7gHXfeI+KWxSHOtrg0pL6JpSA6TQdczVKaHhA+0R/HtCtG3tEmjGJsm22yu
CgvBupPvCFtdPXhQp8BZFvTh+VfuxDRMZ9W1eGUUtYu7FBmY336Gg0VFlBO4m1Uv
wYcKepyABPRGq9DclWLn3MaBz7wEXLzZBA6LWXMSZjEkSNrLwHfAMskkHflR4Bu8
OLX3MJWiUaI5padZUJYa2W78QydVQSNYyshB/9fG/GMbTuXmc9p+OinC5cN0cbO8
sEVE1WCN8lqIJxYZUTQX0KJPV/PXIFDkyJ3zX5KCL+ewt7zM+9LFlrGI7yoQPvR1
/SinyxPVzseK11zNChcG6Ot1+46Bm2/BO/SS008H1HTgtbhqKV9BD4jW61/O0NqW
F4J+LmgSja7BaCsnd8Vedixnsaj5sv2ZzLKiSsC0gdUIK9I8yIP96WTi9gyezSMZ
HP5DD8CwRqsybWtPRX4gFNsqyIbfdmZunKeONXUfl75WU+/2eV+CxFaCdtQbgM2E
4rkf7heAzFOKmkjse+25iOiyfvyVWjuL71UfdBvvlHcV4jZauo8wVQNRbiKUJHNf
ISv81168CNyvdJZD7hNMEEIwV4Xl1n+dUjkXievw2QjxBJG4nwc3GfHyTe9hIrrA
cpHhsSCcvI7leF8IlboInDwqAPktT20E+XYosFu2XYpHOUjems6xQDuzMVWw7RYw
LgKCYFwIIOhEXzkBN6p1L2p8xcyxE/6AGVPrx3DwHbD8nJrOJILsHrsreOtbiCqj
XFByBdmJjwRRB6BZ23Fru49aXwnKvu3BalF1LVTsBBrUQMcO1dBBLvLxDvDOcGQQ
oP337Qa+M44Q2cYEiz+A2c9nZPKI9EJxdvZxG4ZdICvfMZtmCMQ5a6JZl10Geb6K
J3bhPiqrciEcoUxPc5zDgFyUbdDa0n9P9/+CwDLDwf+HtSNyOmIJ9qH6hctu2uSn
ghuUr3pSRz4Y3oOAKoMwZsRxHH2VPxpXja4nTgJJwRTx4hHbPYAc+D2tnpgEncpn
WfGOfFP0oVKkpyjcNWrFi7PlNl8bsWKXamWblh1Tm6JJ/q+ofwvgTmQstcxcdSM/
NFFjifE//oVCU4UaY5dhTwFiBH74yvAFG9CE2cnthTCF6HobPZYNtq5/fk5iYb7C
7hvLL6hwVuGIB6qE265y1taH5ylmWtpAQscNk47PDLpiTMm15umUxoeDBmoGbgiC
n0l1oX+uZ4izQiI/QCjVrGMEbLM0gw5zIRpAMCvYX52/Mem9tl/mE3OQItvMfHR+
QA7Po90j7bOQ2lzaHDDpCZYUejp6LrFhAXrSG7FzuTm4pY7pu4yQjrYgtXHbB9Gu
me9OwKzk+uXlznVbyQ9ZQOZLcGIdQn/CEOihuiKp3iyNNqkmEi3p1tQx/l/Uql13
j7D1uRdaaUAr/Pw3x3ybdhMPsORmum7k1nxZ3+AxSqwzZgxbKPm/yAWL8eewjEkG
kktXUoRd0mF2sbEc/G7PnPCV4pvELwjI8Nv8YY+NP++E5gH9jky79P2D+DTeA95p
BXwN+xCpEqsJ0jj+M3ZlCKyGL6H9l/N5BGiLmhXaFfhFxpzZnqpCts/Niz5xi9/2
13WCMefuYKhH8/mlslF5sGwglcz2iT2c+u7neIRGpV0r+jLa/cWi3U8YLesvrVV4
AL/uStLWIC5Bqd75Hmjl/MuGIWjwj7OgycpXwNeMrXZHGOQCOK18hDkdHAkV5o9r
RPCInT7pO931lQWrL8eT7IEwdFhuX+JZ4tW54jTsH4PlS50Q4NfUywjP9zPJmIZ7
dowNrzjfKYJQygOkbuuzoYgmyrVWkQDOqCVlnohHAaouI8hecWzTEHrD5XWFzlDJ
YyTZVvDtY4SJI+nLpIL+hVVlW2bOlt99mZKlSFjzjL7ngoSP611MTlzRejz8m3M2
MWpShzx/jg7OYSfD9dd7JQ10mmwzQ8jyy28YzCTjA1izG5hMw2f+K6c66tuHy0+c
Co2veEKdZflz4hRMOTagyAqNNTqRmfgLFcyP3gMzsJTy4fckyAgSCqV8y9AYYXqD
Vf0XqklgUbgbdrHCiJWGeWfaXPV6KsJb9OWBRMRxX/zN49Uwisn5wtb27cqdXj66
jhybQPzzu1+YUrZYWFyNvIqxniyvXIp8LweTfbbIL62/oFrYC0eTEuQIO/o0ov0g
oAMcWj+emx7bG/nYYtmPMn85oqTkypTA0Fb/VN1XcjE0eWc6Qu2tue4u3rJEU/Qi
vaJqnZWtuAzfvjTX+GHa9/pkF4jVMDHgcwQZFPrzqaQu2BvyRmibknVc6sXk8JAO
YJCNBNLL/5+h1zYoPrUZtD/z9xcW7cQ0GuiytYN5BL14Z/4vZq9//jSGk3WL9cvy
XiYfB4Zcm5rjaZXD8ljN1IbwI3/fYwkhRhdMju0sScHEPmWYHTCWW4vF1FqKau6B
bqwbouOFGVwP2+vQQ4erfWHjEjWK8tLiWBYSWZeu1ev54Di8UVvfNbsDulc2YQXL
Pdcpc5I72UCZ1/GeWfy6FIMh1JsD54mrjLQGh2kdPhCYLIEHAoqUwICQMZ6xtYa7
ss8RCNb6LMNJBLas6CD0Slk7oMdHbrGz8b/JQdxo1C6+I6+kSjzyMmtVUxU7mq8e
2vSwqMPsnaE285TtH3TmFBcusiMuvtoPN93iCc/5I1BKnykP06SsZ2XgdyblSgG2
Th/WTlYjspDsIpp04XGodedECbSI/ghfmvpi4h0gk0K6q264Gz4qJtSEM/3Gd4+l
1tIUIVUAP2DVYQySjbWU0vRflCcjNn1Ncljp5xuzy6f8jRAuXucYnE9URSJopb2f
EIExcGA47cXug3CCEkgymxPxbcAojH+ckaboalEDve4UFZEK17tvH58eLdwTYlCv
l4PvXgVRFOBWDKI1egQTmgnJpdlJ5CW7vvGWg2RRrwLMf4VPoKTPqxBQl7Tc2vdn
RZT1DPx3Ex9HEQe5GMHANdoC88L46HDktw/zeK94pHqCCd269O4TnHNFsyV3jzwS
7Uf8M0NzLAJmBhHX1peKKSF6561Cza9yo1fDEgvpDnyLIO5VqP960IiNIacmeIGZ
kbuPMwcdYoXBU7kWszaXuA6OAfwHRhzn4DzBFgKNEW1I21kxib16Zv4dy2Qbvwya
qSPkDpYpQj8tm/OlpSjdvgqPyIu3eqHRbSPyNd0irCW595sMJ53QCLYLYYapYEzJ
oNRdDGENdqg6xjlgLytZKqT3PVgcu5vpNm0FMT96OzfB7bZzmkuIi1n74iob22FW
1Ln+jq3X5irIXP1OoHO674bH+Lc9Ec30pwTwhXP2tKe///U0WhI512ipS7oKEQUT
MXERTyfpnTJFNQpPI2Zedd1ycrSzl7gpQjE0Kx1QtJkim68C1fjCGvrICsYoxE6b
fExbUe4BBVvCIXFR7opkufGXBkcEMd+1pG+DS63Iq7wS+R9HyiU496/6aa0LTF3c
CCF2by3sfgcFO0E1xXLv4GOx1OH63k3AdPDqAR8B05u1LZEiy5eHVTlg9nqAUOIr
dDdkSuFnO1qM8At9SwV+07HuZcFyBuY/LESwjwH/NGkoV/1oNEbGT3VRoGtcP2Rj
IkeLO5n61//ruTn+7jYihbCcdDcSxrFnMIEJhhhEJk8YgpY9+kS3ZogtqgDEM8OP
ONXFNQqsmaD7t95+DcoqAnHElQx8s5KwUZb0wkm+xM2hbFbG1vakbzFt2Dm9er1+
/y0DUijvN1zgSqJmB2GS0gtH6ZgMMCvpByi1JhUWjZdLhRHc2qqnzQMVCyplhpX0
sflaWFOE0rXRoRDgIQZWQaZMYvKcMp5u4YX3hPxbt0cfqA0KGkL1RweM/6ozgqTQ
EjWiMXIzmL/8AhaCAk77ZLFMWRzfYzVK3wAoMHO5tmPBIuMY+kLZ3ecei0OqlqDe
DVeyEWXwyAniqVoaRq5qo+/a+PAsaTRAg/GxxtLS7wzbl0CXssdAm0XxU+FV3wzJ
wkrqtiJrZy63TmpfBlMEcB3Uf7+sxeEdL015DYjKliOVvFGTM/18hVhGcb81uIfY
nMdx7K2UW2sClkS7Ba3c97nypywzPWwO6KkHE5y2W6WX4+rWhFpRodt/CuvCAYFb
gFwOfomdThJ3SB7B5ZvK+ICh3Hv8iyFvilskFIOWPkTqwPtVcdK359yFL52wTzUL
espm5HTAQXG15i9coL+v1VDa0xGi6o3gt2eXuIiyaKLy1SXG6ZMgsP38U6JS1VAf
QnSZEE8Iq0w4f77pzZff4369e3bZ3MyLaK3BJzmOnVmiZxSzpZ1K6mavAeEWjeQ4
xxEL3t/3r/vUz6Udn8Vp78G1Z+G1s22H0JM6wiq6DXLEdi7es8vMwXPDq1bG+p54
oFGEaT/c3VeASeHAPpCkNAiHjCE5RfObCuzu0bHTkuK/f4n+IaoKydG0dpjNbPOg
HSGH6Oi9+iKNn3v7Fhg7MAxW8OvyLFgI5wK6mYfiRXIUPhDb8sPC2ZuCU30h+5JR
r0nowtFgGHTWNz1b3mumxieR2OAFPqJw/YvYDaN7q9YjRTpKjpb1+fq+y5kakIuP
TQW7WESJL2HPJqUOaQfetVM7uVBqyFQ525bNwanRgV2DMqClJN1niMq7QUJbX2/I
0+Nl16Cphpp3MvYXkuNkcl4ZWzfjJF2xd2llKcCE7zlYEhLe1Oe+kQrmIhDQVsB9
7gWzfVce5K7CUFy1tQ04ACPFRZH1YWYudeidmvTxqhkHpd6T8SlSPY8k+PCtyISq
bG+WBsaF4xivOaW84y5StVM7oiXR5+zuEUWehA0+r5H87KFKGVcPIX3yj41yXSPt
Feo6WbETP5It29n21QMh9wq24UaLCaT+J8kb1fD9Jea2yt0qhvOEtkKd1lo53sdC
wtNgRbDUcNs7HW24jSs9CUaYEthVAlqljEQhgyKQBGLTghNjqVbxTVdvu/CvGhSF
N02yswkIDQXja/rua+xWaKyW71amCN09ak/TaqMZjxAMcv8RiPwJh1Z3XiavhLs3
WNWdYDyWwdnZC77LrqOXi/72ilrunmv9YCgjpomGo7hJ6aeinxpksAzscjxp8Jay
n1lFIFZoRulwMFZWUSfZNtN6BxA75iKX2F+iK2sEVM/fToVA+qKBtarKb92drla1
IXnK6xt79KhmFFB1LXJCy1TUJW9AlD9BI2HUgubQrt6eeaDe/CTDnJLaOS2ti65F
1eabiAYhNmUFRefbKd8D5wEKCBlMZGh52ibIHrQFKEgXT9DCCy7IIUVVxHTcN9aH
MitRAZOOIPr7TF33f2PAGkVKtAwJP97T3Wzb0XcrKjOS6egu+WXpG3Aik8cf19M/
5/FHosfgNCHVXbzzyaDvkv4sr0cmmAv1sJm3EvQZnss6KQuooNco+pjCLehB+bBh
iTNY3Z+1D+NY5QUTBn1obdYwnr17T9GqdX4gRv5XrOtrhMU9CFqmtT2B2tO+w42q
nd9Eh5gA6lWGhCe/13DAlYFKZrSUDAqTYitssZCN3oq2TiGNXsZhi+NPPjuHrMJ8
U91f+qmw1rlYY03/EVvmRx9Bf2G76N+y90oyGHmpv8RQ6LAKUE+pP5xPftLDGOe6
5IJIJZzCxsEbmgeMSZN4U7ul/IFXq56zB1V/PkGFfDvOq8to4HvspbTBXgQBIIt4
XJzAr7ldN0T7CjiWAFh3/OCVx3SHgScA8F/vxvPWwy1Z6sCT/UxAfIgQWdFzCACO
0uk3uULDy+vqnzawwsK9WIdXxQukICMWaTaV5jdkLOqI6H+aY9YLTZ/JmUO2kjdQ
/bUea5zQBJTo8uMBBUy9EekVRi5X9wK00zwpD7+QkgksoPD0zHbtrwGgOQx3qCHG
88UlrXJFfeoPfwG94gBwutgrvely+Xb2RS1gDJEXB+SYxvDYWRw8WvFUGW2LwK3v
vP/U8W4MeX6pLdbGIuv4j4HAGCaJsXuMBnekKdIWA6X7OGKtDkIohCIpCZUQkfsj
QxrprqLTeoHf15aadgestzEm0zzlAF7sTOJrN/q8lxcLidY903P05IA0DTI/MY3W
F+Ry0RC9a81crewlxmnXqwk3lb+9dJ89/yQaklCdg/L8SfTXN2lnC51FWnDr3Xf5
EJD0C0KVlDl1ZfeSLojIowjMqsPlsJ61tpx71vbx3JWWvleDcsr6rm2Z2mM2R6Lp
sslYJxOxC6IX+RAJj0IQMTyc0DWQqjW1t/UV5nn7XBJhWr9MioNVLABHnTS7d7Rk
9p2BUIfviLmGE90Mhp5G805I9eJySpYW/HB/zhCbMXUbdvSseEC3ZZw6qDK0h4hm
QeCHwU3E5Lz+1kDp3Ptru4Ga3UIrPJmAEwuZ6zpoxrfPDP/qGUVmisrBX+zHvPzC
s7qWiDjwBPv0eOH8toAE3lQanR3G2Ms0fBIJTvc0/TIXmgPGaHnqx9YDlHleSJxh
TndSyWS6UaSPKGL3Z1pv7rs3aqR1Y42yPFtF68TbtaXdj8HqQ4BzndVuBgOYOl/l
2S7mczL7kluWVncS7ipYtuZpS2GYUFK/l0Q/e3Ej9YsVhZa8ZxotI/KJ4d+/2A1R
8dksPrtp1iBW7AXo4DVZfnsxAaPRpIOSiFpcWhUFN2ck+yBW1IbVLOIA0MrGSVOw
nFbGSvb/PBD31bjO4W/4NW0YEPLTQ27SJmJiHN87Vm4d704ioHFZYokjKD60ZlPx
rK9y3lU2XfVS0ltJddbzq8lzYWsW7p4d+taf6CrgoXHjjLXif9BXRzZYzIiaYLHI
MCpo4koKK1Z/JOO21/G98yxY2fez7G9B4IvcDoSn0nmgAg1sZCpUkPWWWuulnlgp
azyFk5eB8VOCmdtamefUL3NRywAuo6VAuKte+/SGJoJikyGlb8brtwnSi6wlpCE0
yIsfVE9AJqn+VTBi9MJ7o08o2J4LajkkLupIj2jHga+d89a64LyAPGSVtHPf3J9B
prpAju4D+S6QLHVSijHtQEtnauxfeKiMtmDe5D/IpisSJzqItM6cpTDxoCvx/lOY
f1gRJKIHiIS6Gz8eLXgZoSc3afPEx4oqksxk378dKQjiuavfaaAWTvPaqiBRB5Ut
01gfnSQC2IqPEAuT4FrVTfeYFKJWDA1eoNURdzIBp2OSOhkDhdPs4zvQuSlABDdU
YqrbvGOywqcpk1Zf0yxMu9NAFSNuHVtvO40YUiZ/wKOKrDG1UWFL6jcRqW6L7g14
gcFojPSJ3a/PrThz3ptGyp7v2e8B/4xlnIV4fDNt/HxN/4OjJtPbDFgEI8IhTlz0
RwTAlXKAc9QJctTSrNwRufrzwjbtfTg2Cf4LK9m2nF/b5lD1dotQmtbvuZXvQsK9
YeXdNSVx5tShVgDzl0/tmPe6ovqa3RBG88e/OVlQ2HdkKuroeJhhnraud0RR8gIU
6yrmAIWEhy8mvqkfjZ48lhBL5mmF36RCY1ojJQmfYrNwAY6KItbXUIzY8JtOnSQa
qqy2HyjSt8tjwqYDyzL4D7DMeFAjAHogV7GJnYlgwTLqlOqUep0ThgvqWpDTbftl
5VGMEzv/PQyKCApfx89RL2y+56I1nMKk3UCKtzn0bc3mZTbR1TJ/W6J8+aTVL+Qp
7VIT/VRhiSM8wVrujKYozHCOEmJoKJgPpexjjdVfyZs5nKSjYS2Q1LQnqxQyHq70
X3fwzcIk/7+mnxYFN+oxiw3rCrAToszsWFc0rLhWYTI74/QaNljlSFVaxK89NUZn
QZC3BIzeS8QN/SHAFoumU8gyiKoz8K1D1NGTN54NLu4se7NukT2LWhVZGr2QK96D
ehaO9fr1VBE1m2UyQ5VBBgwpN1rxsvbsAGgJFBZQbp3MPy/DA9FEx9+HtoNbLMfa
hiBO3JlX/+x/avSCZz+Hw0tCqGni8WTMp+GDlUXo8Xll4WzcwodfpKgibybrP10Q
kHvNU/BUxFe57EMu+dK4jXk57U/xAb+FGHcliBxHmChQnyxIzBS4b6HayVCCeYn8
mTy8rAkT3qMjp4+yyU/iRoJMCT5pv1xaTbsxyrOGs15wRY205CmgQFU1fKP8nNq4
RzaW+H9XunRus1gWCUaPMclHLs5+FGrdu5Jr6xR/vBuA+R9AeC6cFMfpqxnItmq0
GA013UiLrpxeNsG4VeZ1PAJKpkLe7ryl65y3SvRxIbvx6dIrkjVEZqO7pZnRSWoV
vkRuweI1mrvQygCh+HdYVur0rFHBmz3oPJCPudxSrTkGQrltfQZNd2+b16in0afB
uGF27buT+uFxoV/7ccPLWMZWLLYIBMBdhGgejkcvo96qMjlIMIL/ZIw34dMXKOOT
mHXjofhJ84VUOSQC4h9dKeMArm8woiOeKiPTfd+OEV6SroHJZHCADyPWMGh/6GRq
AXPT7mXFRzxyLj0Wjq75sQimTAd3Ost/Kp0FEouh7ktha6lyqo2tXF/PVEJI4WFe
JDEc8x6pLr/mdqTRFJNBZ9I6weTpSPyiSQ0POAsPZMsKoSBbHqitcHDlLzO9EpmM
pKFKZbq34a3hB1IvO4Il7W45GwMfgSgXFV8/jg1vjWCd5hKZ3fAwwziot+wawFUL
3Qp1pyQ8QQn9nJ5iT+89KQwOXhCDoHK06ukDKrdUCdvQvAKsXPB3ZTNFmDK+oVh5
9SHkNRwzlyx3NSo7g9byX6mfPMN9in0Yruw4njaxzjWkpyeNVTnYxirY/w21euGc
MMxRm24NCg/rMo9Nu5vyfrP2OMFhqQWJ/9FiE6AySvS6txGJyP0+Fv+zFxVC+zc2
fZct8KaiRkBfMNVqqsMj4lw4DIE9+KnYi906mF9RWvVHH6vjbRcAXR5lloiyaZAg
ykLPKmtDNV/W4X3BDI7UX87T3UgHQnG/OkxPrCbteihgT2g8MZE1K9CMd2rZkaX2
FlN/LYuQawGNCrF1+BXcLDhO2XzA1P/4ffSmnKFZCilAr/5RpEXEjX2E5uH8G1fX
MyhnfIXb2FJY+9I61aXOSpJTCV/PBrMYaphYIQG9qj+Gi5keAALqNa4tVQTtUOAM
KXa5/qt1E/H/N++WIS1oJW+VQHi6bHN30wXl77I4msS+8oC+WfXOFcQ4syBKK2s9
ZzW+zQ3IhM3Ve207sBI9QwO1TcZ3MMg7Nda4MPllmjmawKRRF64t8ExlotdmMB+z
GQc+8nWIrJxM+l4gSSLgRwarahLqBDrfEzpDuZm6e6AyU1QG8jRtO/B56Q7rzadF
8huyT2Ao3AlpPA6wUtfYTjjFrHsB4Jgxww68PfoQT4DyLPWywbmeExbju/YxLsw+
6rhTXb8LpaqfPBj4bt83JlRTkWdq8Oj/Lt7DGDtQFrFQ9nCoW4uqOCU2pQOUy7dd
W1kbYPKLG9dqcqS/OdvK107GJTC+tcN3AcFeP7PJnGW5pDKCpX7rJdYC+9s1jykw
rphqMsnf4ZfmINhzYPVB7M7FyNBYBvhJsTqIqEfNEFGvbrIeTvMIu5sMky+qLE3o
bC1dCFoKjL4+G3uSdjCraht9SvBLkQIy3Csh6v64iGQB891Wsy51Ys5xEqNQR/BA
5QatdNchpqUXI+Nw7Ttq2JQudEFa5sv58y5qJfOFgKV9Emq6RguNt4j1p3vP4CxY
LurubOyxuttVMgtSUxaeRa9I1A4wcj1AYVpC2mXz4zHajrWRbcto/45uIITAwmI7
lpmGWe9dBv3FvMIMJSzuzPWsxOsQVUjia8qE+hpilAn2/HKtsiiIMnxK59vAmuTn
DHyhoYcEAxxAJB7iq5ER3na8jA2aqH4uatHJN6C1bHz7JL/jCwB/xa1owVHY7bAf
L5IYy6IiXzrfoh7kahiKEKNZ1XMuuzh9FRl2szJeifEK9wJKKWoCD0WPi6LyLQgU
6Jsp/xYxGBNq5St0NbJDw62zl+3fXVE2zGNBWHeGozjh+UV3cwtZeCkvYLWrfp0V
Pt2Yrz5vK0ZHllkElGKT3RlYuDoFVG7ehPqqtEcWqGB0P6BuB6EoBa8kFVB6zgW0
+b18U+y52R+xxDi8TvPI7GQ/6siaFtEDHIu0gC7Zd/0tr8MxPFt83xijjDWobqZs
diY2ML4F7dOVhX/klWBsgWLV3AqxcWUyhP6Sn12UotoizTZEVN/CAXKSTaNg8qpH
UkOMcakhpfMZUIaAoYHpuA9k3Dot0x1g/b2Rdy55bKiI4NzGlSuPDd9yB8yto44L
hgaSQ4rHrlNgCWO+5pmcvVAXhQTddIFLhQp+M/bw5QkcUM2N4mA6QQDpCjBfUaD7
YFgMTYvg/CbDJpeVDSXsZIBSehqTtGuTJrSC8vFV3FNLnBPoObRiJusW/uycRbtD
wyxWkQtUSPCUY7JQ2B2RwyryA3n8uls++qilH06xNVCkGGSez/iyQoOIVDt/IlnJ
pRHWK5SImm1ofbLohQFjX6KSGwf+MbHF5idA7ZCgiHP9rtHChEQdAHUe2Odi+pki
y2kYZQZ7M+aogVlgGsI/7U9Tt4UanFV9GBvIZDfzGUhYNMVVBmDUiFENtRWyNeBV
GHCeFOICareSNlkWwNjQeBiXeHneKvDg0VV26yuKg7FdLbzrHzf6YaWmQvrGS7Vr
QmDk0ZiThFh6caBigYZAm6w82oFebsrlVNdpHyM2PtFGNHfvN+Kn4xrbxKhwjbQI
DVmWqlGGGVvP+zNvkteLDTu2zIbYgiYbCLURX26TzRFDqiuh/DV28e7DPzH9ad/9
KQRk4Uc0Qbjv5DM6dZ+5Fr2NGhZ+zqZZSnnSl4yWzCh0ZMlZ23ST/W96n0tjGUdz
DwYSHOj7Fd7tT7KwgnLEVtUNeO1LK5701dcGzvnKgC8OTYQ0B9MybtlHIn/evFIJ
DqJ7b7DvgwUXktkCVapDjmXwxlh7cd1UgV8Xk9iP/cmil7EFSKZ8GOfVFKix3U8Q
w66ujRCRTjDFDWfKGtem2LwDqtNIH2u1MbhprC04GjlsT+dTOlAv3Yo3QHRQ2G0A
nbLYC3IVo72LvkQwJdbcTrFHE9NaJsUisTPKNuDtLZF3JgrxI2nkQrGBqKWZrAwP
bLPSCNiWUsboKIm/AgfZVeaY7j705uFG1zY6+8bZlSzlvQ7vfm14HE7fbDOrfshZ
JFwfCCqc7pen9nH8Z4afpWHVNAv2as5HtZrMlB3ERSLh5GWKJewqN1BAbdLe3LE+
ge9X3d0XBDNY1idHc+6NPnPcY0mhXOceplNTT0QANKIJ7KGg0s4R3XtqPaQUu2Jd
OZQn/O+EfqGx+RIoE7biotoAzIo4NHL6sPRfuZhPQZKYEtSmsbKjaBfQ7Xap26H3
0XwGYUyLX/fYUV/z0QMCd6qGeexc2j9vqgJ8Eo5/LVL15LmlSw9yYlVhe3CsvvJV
mBnMGZrLLWZXgAdwkHaG6xd69l0g8MT7/t4d2zECoxMXSr+F0TyDJy7PapTuG6V0
mvCUqux7MowPcqPCKhNdsGN5q/bwbYb1JnGLdmQpqrHIGA/UyOIBn2OVYBLLXURp
b7wFqXXUx/nstWqXbkeVcK7OAz48P4aLdEqitIGrq9oYpKYviORHY5xokxDgo5pz
QPGt/8lQimwgEB715z519pK0Wlq4SMblbzowOif9sL1UC7GSE3J76Tk65zomMOJu
3OtX3gosTdPNb5vnsOIF7I0N7TBSjRdAxNG0kha/PNtwDf8iENxgSmT0bDy/aZiv
ABG++tLFu1i5VWALPpXDIY4Y1R8KANHubyK1UIwGOh/F++em0pWX4DB/YLF3qIMl
PXCG9OCxAeDpb9DHnfTcuSgzyNHlJVKVTwsBWPSJ6ZTDqjfeRUNBJeXCto9Aaw63
EjGETLoIWxdRRcxX11sja2fnqzNYphshmeCpKQwCdPu0a1W50abNwoo1Iw88xpoQ
6Rwfy+e3nKnlHSdCTKN/ti6E5AAk3nEHlpVBOugoDE02OLDo9vtApMHSsSSLHW2n
Pi8sA6G38ma2yav6kHEZIX7ABpKAxPG1zYooo3VG4IjB/mLinCBvIFVitEkzwpTl
v1y2QFK0x9aoW5NoRdDrQwr4TENqGnvujitYEizrv0TJ6u6X2yGqs4Xq778yoP8N
OGe8jRNytuMtgr92VQ04ICAghsM3WumePeVlF84ImN/24Rsnt7GTc/KeSAEsUS+1
Vwf4ribBTjM95MphR3qjUSZoDWrqXETy6G3W8cTGWiSIHxmTTyj7MWy6CpfaKcse
kL9SYJYpI0On8i95EhAjmNQZwVgmp1SyuXWkjgRLwwfqPfI7frM+lnRb8I0j8e/7
iU6klob4sBDl33mo6aWnD08MIuE+WqPztDgSoyXJSvCFaXS104CgSCuKE4MFuPZM
tpVgxpX6Z14ahM3dTjDtwKTqrjHfX//pkHHJzJPdFYmSeLn798BBc8VpNI6GJZ4p
0nSrjxY7B1j/1R4OXnEPxrjpcqz+7R3W4vSuu+poe6yIIUkHE9Pr/wXnxsmLGiGW
nA9zBvpstGnPpzD95kT+3ggJ4M2FZTMZgcwDK6B4tal1nqj6HkLPjnYBYLGnfKHY
lTxoaDoalM5M0BcphpFX0otydCG0rCvYjbJ8Exs5tQq0i418sojr2/3bRKJSnjoS
/xTfSUCXt2JKxME2/M1wXNE5vSH5jVcZA6BAIol+MWKx22FAoyiTn6HNywsOHkf7
2czM5ClttznSONPhfJPpoYLqnnsjuKK2zzkdSG2aF6r9oJesjDFRiOb3txyfytXN
HBickmTXg1MceDLrfXDCFZ7U8Sa6C9wWQiuyBMyum+R6Leq1uiNCLChu+NIMuR6A
j1ji5o0NwRF62ECRCZSNy+Tz4i69jCnFR0dvXsmHvFeYhD7g9eecIFFXmrDwSwE0
x5k04ywBUwdn5y/+oQrzakqOa7gS4h7ZQkS/KwotkXNjdPj80DHK0q9SJLQOBYvC
wEmjg9zRomo7aDrCYiIwQH2ycVv6fSJRjOvcmPF7He92PvX7gwlPpmdGivuY0Abf
VPw7h2HQN4l8fCZ/edZGc5yrVegW2DFhApJXq8BczopfxnkR9hvJmWGylWHywqxI
91ExZUhbg61GTay4Ktg6UzC1QKmH+fB+CxI7Q0uqBeqeh5D/4odPPSXy5UzPiph6
nQddxMtjW9EuXdTsTVreOI1eRehVxwbXeKDV+u1TgcZBb8AA9vvwsrhHnTlExcZ/
4F4pXkstUxSUww+I+HY4cILAWamjQrOySb2P3aNU+6N7BqYCzgg7GEFI8UrdE46z
okIRAPJ2I0OhL02HJcOc2jtCVCUgb8HV0LmES/Fynb3M/gwiDGSMUE//pNTB0weo
6210VWHfAlk75YFKUPLI4JTzwf1TTKyNq9isvnLZ9Kgq4Cn0bYLB3SvmkuDkQZ/5
BHojmDHOIimBM9+wCrpvQ7XAJaFy/QGA7diOqwePNUO1x702UZznGRDaPDU1eiiw
vL6vFSom3HM6zNz8yzt5Ey3O9veaA+UN/KO+2UmsMmzA9nqCI8dwCg/Rc2En92ju
QxeReJP5ra7knNLimLVmbYVjWqpyd3Wr/K4DU8jZ1TH1jLlRuqsqIo5c3c85yaz3
YnJAQrd1vg29rEGITIyjUD9/NYsiAAHIYTuKOkkPuxzFj0pGebyNsLg5RK5ek4ox
cGMHj6gw7bAP+sssWP4YfLOCLC1L8jf7KM5fEAvRzqmMMGCefaTuGpN5ZqGgDZIe
WoRwKPYVS+5BdJaYElvSzqxnt0wcy3VBk0fKqO07u4epAkUd7/J5LBH7j0EXQ+tc
hSsy8qLA916EGZScOhZfZG1XgXYtf5gSaYqFBolEnS2Cswiay/fjzjrKwEr4E+e2
GXS83hkv31UO1oz7AuMhSKFSJF8Q8h1vSgZD9GIa3XSk1HT0ZroVajttvnZRkTlu
d4TfYAsEg0a8uqNMXoe/fjjpINOHinB+jwjXo9spFf5nWiXJ38BUz/Wq0l66lXvI
dKDyAQwrO+NlLAD/kSnoFH6w/JXtjF5wbp7St39kmnfAckFHwmDKXVAB+2R68HEx
EveclESH26ZHcq5/pSHB6EAaEVPEOJ/m82sE/b1Kf8rlfzpBqKuN5zS4szFcDJWp
zKhCd8eXRgNddcxWhR4FAqvao/70h1l2pL0oSYBOLIX8+sQIsThwIHL49k15/6Gn
PziquPTbtLy1g8mWU/aahCvJkQbWHFFqbcDTUP0KWtk+8OyRGpgIs8ftMKVU9Y38
86+S0OS7tcFIpFeLq5ely307zOJuAxUazHLHPXILjFX+E70HNDpJcuoGcXt97tS/
b2pRyH8IkokTQMQ0y5Qo18bVY6F2+lRmc844a9iVbe6BeRuyGBtxj+Ain+MsR1mN
DtjiF7SyWSQ6mqe15cgY9gxdLcYemaMNsJukKyUo3lQh1snvLVUqxkFIR2IrgPQX
Aj88ceHvU8JYXyXOcT+NtdC5+v3iBkiWNEplCAJpcIQjqpCvD0YPTr36S3pd6Dgy
coXpeJZn0vZaoQmvLuoahrcgQVkoBlCtXdzStH7HC7txpSxo1G5QQDwR/sR55VUr
mlx6yPl1wx2iG9va6ILdaTIc5C1ve1vSaeCCvNLJt7JobkF9nHZr521WPRQk1fUJ
VMtK5poX02J/2/H/m4ouL7NOBiUpTqKI6zmx+2hTBxwEAnLC1z9E9Ylb7Pe6mjp0
X90U5DYN6J/CEQuF6pOe9g+AGHTgu6BxLwd+KXkHCq5KZpcKd2NfxwyRWRNhcJu8
gMh4/AfPrUFJxIDgOiqFiivB5Srs5sX+Flh5JRUOkKe3wVBo8d1kscaeKs4wh9tJ
cIJsAZbUOdLfmbtwGutMAZZZMcd3MoeB5BaUE/00131jVCiP1tjWY22+kg/2f2GH
mlRZJLis31Sikho50bWIY8nDoMPZUEpOSdqYpSTX58U909n9Os9MT9WQ7e+T6Qk1
cMgg21cR+ADDvmQ+IDWeZZ9WS/UzVc72kH9tlGUitraPT8f8kyre2PesYVqVh+p1
7uaLdin3fJZWLP9eEetASNPovHyZp1yIf1O2l/U/DE6pC2F2lcCX0e5jg32xYQtb
Xn030iuqY9wfRpmC0wckWLgGsaVbatubirAC1qJ5ioq4H+UHXdWh+tYCoNVAHgsb
uCE+Gd5/SpJoTk1o9EtWwVeb0V0fVEA7tZbo0I+xzATKlwapZ86bXwxMVWZ0aMZD
fOhqUx3Njudh+SCrjThb7tbx4QODUOx8G5nNzK/mGNLbq1T2TJHVOZsqSsqba5wt
JzDRxC19IrAHqdI6FiEKfOG12kqv8FCx2UkNI0iiUWIe8x0T0QMfGVObbc893vgY
ufo61WTZExpGd+las3ymfsr409WH8CZKnKS6Jq/tecK3TCA/ImbvL4lZgFvCHnxW
PUwx273prwGCcpiOUy2hcBQQ71MKusukuYFnTwTndl6Qi+H1TnJbaYCDXe5o1lJK
pPFezvAvBnT29SB+Y+L/dUyVASndPw+uovgIoUA+9IagGODHohg3Xz8x7wm1NdIz
FI4m1l4JcGP2gRZpmSqNDpHQaWhK/hoky8ckvzqi/bdjHf2HcnDE8Fy5yWTGIFSo
J7Y8kFHsgfApN5LntlcGzYgiCZkpyFZKhFCKAjz0cXp0kLtFlZ6ktn/MU90AeFXz
Trpg/dxWnrH13Y5l05n9MDhqlP+PC/k1e/tL07u05ptbengWbnQDTGW21KisqeYh
MzfxMhS7aDkisSkfER4WrlOOQIdGrkoaC7009mzEazcS0oAEcDMFv5Qmww1c0deq
fioHNwUzeyIeGUtBJToWDZKEchUnUWIM7g5KssJZJJtKyitm/uQ9ulRnbdtOF+s2
5DmiBDkK7+dW7LQi7qJH4Im2UddXgRQL8kBKykA70vtG+oTLHx9IEtwBFm1OMtcm
j/1e2n7t2sG+pycCX6484LZNE08txxcGlo867ggQhs++shxAnxtazT3m+hQjVzzr
HBlRO3bEq5Z7UaH41XsN7UiGpObnI9kr4LoFH4fjWkol6ebXzn7Xfr/5sc46lW5j
fL1ZNWV0Yn9BgyQyxLXrMrUq33bpiz81aVfBzLA6eqjXGzeXqgOP1GnDd7i2zfx4
3PfnPzwye+05OwUFkGJ/XXk0h3WIuMLoiWfJl7RjdGuxlQrz2qkOmyoZWszkCV8B
acOQqGLyQovytCbwVZsKZUznkehjuMhXcUsbPjVYn9wmLFQkwhIklkO6AcrOrVJ6
M/ydhvar3oy5mBW3llnAMzsIMoSmuWa3ap23NBf0Djkk217egiS+ubltWggqQqrF
0o146TPPHQgfagxdPRF8i1tlASZpZeQf4HqqzZw4A2B+ylUajyTjV19I3GNKd0Eg
UeYc8yniaj5x5NzMnlvBH2nXGoHkrXc6A4vu3V1fz+2iLhxun49xJ8DvOVdVNHxX
/NT26PNBt/NO85e6dsev7gjp8e7wb//EWkWMNCrcbMSG9LJ9Uji+OLvfLs/kTLpr
7EytLU3JPXN5lk0YMbvpURtKGr2XP+UdON+yYZLbZg+89moEHjd1M7wkW1+JYYCF
Zyja6xSSTEyNcNejnOvpcvv1vxUpcLJACK98nd/2J8YYPSq4PwD4nKz+0iiko0cg
VKs23aYaB70a48o7ZGQsqAX54cInAv+krR6xtoqOrfFVYuUdQxoDRuohlW+zjbaR
/l5nbD8FC2ZVCZs+6mGME+L6LYqPtSQBtqSXxFuyXV8tuORg7Ee1RstyDb1tuyD/
W8cFSl+BPq9hmxiCOXzeVUw0fnIhvA0Arl0sP0SA6K2syItruQ7/Ja3867GrPI8T
zPAP6mFg4g2scT0rqxRocvj8oHKagiBYG21LB1OOiA320NNqtaUQqLNMF/OEHzs4
lcYx/9IFfIW8QzAKBqsi6nwBrSlAtS8RVzJ2nsTcFDQcZAUw0X+mfX9yxX4phpns
waB4Jzac4a452ov8Va6kSg08jCt6gH2qVt1w3d5OJr3GR/Wubl2JIRymYgx/L2MT
I2dwcF7WMArZSMTmYzOV9+A4aI2YAVwYE6ZS5VTymFUTUHU9HI0enxrjc1A4ZhX+
iA27SxTCRJQW7kdPlWZKdRPgOSeCMuWTl0dgtrkP6qfoRL6HxYWtihfP5AK1iHWm
SfIseILz3N9xc/A+sIPjLn1zFKRBA/fIj7OAnXSAZGD6fIqOElW5Q+kZfVBe1+cz
E2+BFLL5D/UVYiFS8ydEtWtWvzGBQR9fYxygYvP7mT/G4rRn/JzpmfXrSSZDr1C6
Ad2kjCaGxH2vlPQ30SqV/2zpg9LmxPcFh1Xno2tX1YUVp4b46dKRZ9L5fZPT+WAK
QVGNyCeJXCk+K9E9dNvpq9XoR20uYN54F2MPjR496wTpvp9Y1uBbBNgUeLId0Dbs
VCfgNBjZzxSJZ+5x+AI6cA06Ho9jlaec+Ehh2KE3q0NrjWGEQfOkqxMTKeklf1IY
7PryHeVT6WZSJuhPEkp2uaIwEqlrueYjMLHR2G4ZQ5feW+LAAr1J4QnKbn+XLLj1
HHmmby8+u+m1O9ni/3S6gjyPJ7vYqDpFh7CNp6b1AYk+9VanvutWWzZ6MkGHEyUZ
uuYTjqXtBbY8ZmyoTug1XoSJ4ZEL7d2DGXQPkh1Amxqcd//7DEz0VbYNK3MsxxFX
xtNx9vqV8jB6q+gaRQGHDkt0eOw7f2FB03rx6jd3m/cW8/v/SKHzd9Hqf60krXTC
HK3FSvxVNTUdRYtlErw8jD117yCGbLbZw4ns8xd7k1JO5D66GL1OipqQmZ0oNwBz
QqZWqZbQaP08OHVcidPy1ne2TKvYTa6wvrVf4O/ufy2zJwCiKP9YTnZcCoXR7a3k
XTXGJrn659h6TnzE0SDno7eO4pifQGWBSGO456iC4HX6T+BpoFl1FWmnU20aKKHU
mzfa8cbaPHUDBEvRf7allfdosiS+vTT5UAVXJH3fHW5czw2/ESRKBCB0CzWD9CzL
SVRuQM+ERnk/zDPqpspEQuTruPAlN4hG3PnodlKk86UWI/UgeDrR1c1Qjs0TpPm/
UejxIDQMORYvdHLhd5Q29KQD57IQcZrp8pxnHhegGBoEjTVfFaV3o1CH5Ys3WE0N
1rbkAxdtMO2FC6+LgA6tIINBJS92sc0X5b6psKjXqF+et3EpW6152pBKcCtZb+Ip
JTlSo7nOebvjpNlHot1TOby/mFSvAeeXfdAGyqRFFu/towg1MQ/aiAJNFfYhYExY
rmmJGDRCV0VaweW3Y525aQrh4iWiMaAkM+I5m5+yAKYv+rSFxh9lWgZXSaf6VJeZ
5xA0C9gkyA0OfFHMqSO1U4d0lZuW1DxBIkX930Z8iQs1CWayQJvHxD3ia15KnvHW
sgXVdRmIh77d3ntKW44+cxbFNcMhOKHEhkS76fnmyCT1/1hPeBnegmFthNmBNMFQ
2FqwZI2PgMlCP/2XV/rC7fXfnVDzU19nULxItH0iD993rPWqVsqj24OGrn6Ps41q
mnRTgeIcyKMpQXAwKoxdWaI1ZmxtNBo47fBlgTSnKIGcA5PAHmcprg354uxjgVH4
iKZfmZHTkWACpALV1r9At5FJ5GFd+P2UjCgRo5h8nw1HJh7XfHMSlxBfe4+bI0Bg
fQO2iK9MTIBi9z/talGQN6KfRlxPLQa/MV4z8OteEsTYn2inHTme6RB4pqSZ4Qq8
13Rn3cNxdYyEjQOdW/xIze3n1hXjRc54RJQs24O0k6vU4hxz0cl0K1QpDUPe1Bn9
8DGoDv3Al14dtPoufNZJ3dJdw3h+KCxDwH7swkxA1eFC2UhaSTR6fHidyLE2aMJS
BfE+jFGJIEQUvWbe8KKRmGMEf+wkKHyctKJFdUjYOixcOXJOF94kg8YjUcwXFmrS
iuJNYcQpGbSwM546qWYTAJJwKgSpAmds38J6ucgA3Tb8Thzs9dorlxJ47q7YnYtN
jBOzFMW2qGQYc+O10QyClvh+dnDwnlslmGJQtdmigCa/a4/7YJpRz/JucUtXZQqC
6j4BAuVUhKA1Isce0kJu9Js5zEf7WYwg73fqdSdGKEpJ5w69JyfyYT7PW89CPH2f
XGAs99lNl4xIAvFlXVyNslF5hmmJt6mPXT53uUxEonZcFXYwooawqooEW9Gu2N1P
7YSYYpU3gKi6ZlPKjwSL8jW7CBIhm7HuBxy/NQFGk5k0mh/b44kcv/WQRKdWoiYf
byYS/8R31hNTAc9rULsz6yLlNzExPou24ckqwa5Xz2FW4kR6ikpPgkdDUsee5R24
eOT+GHryJYTYAt8lCyLqWtBNv6eAoznbQwO2gxvzZcm/NAiFCiOnE5Nxfj2NQeMP
pztWWfcyQBuvpOsCJFioIo5n1b1jymWaMtME6B2e2X5ngEOrJgLictwJa5j2gRXH
Vs7QzY3GMVZRf1ZPLK7QCCSnf34MpMD7BZOhRQWTImxxTHMlwH1O1V+qijACwWeM
D6fZ2+VQtrsleT9787VBsnA9xoT2mCR7zVhLlw80XenTdObtZK227mapchhfF95+
/KTj9RgOoJFcw/HqGCOjuW8ZqbUeKx0GB2uD5JpdFDp7GAPkaYI7kXKS3h2hkZME
/0VFWN1LMK6qGX/PR85ZeoQVMfdLxPFX0JTLxEHAagqtoGNlzJTB2HtYJRax4ouo
o/Z7AZuzIshmcQxRinICh2uqo2juNfZ+eAIL3xJvwJOXQ8e08fmF9tyb+AvlYKwo
oqO0F3wz68IGbSyodOX0VEFf7Y4MOC2c/qvDZZmN3/Xp0xKVqaM/pvxGP1au1HO0
vnIo1Mo6E/+6wucZUoUwN1SjcLmFVJ1xpeh5Gq48me6l/tOV7w+gfUxPel69d8oj
wXOUgiUAKRja6iIx98WMfg+xIP1Z4Mmh81tRVvwXEt4mGqShBrhDQR3jXdpJ9QEs
u8Jmi3CaKL9NhVbU/Ac5Qjr0BlZYU1kCBypy+qI8/ZHyC9o+i3ixfLVXeOn4szCZ
aQmMoKHs6i+cXm2NcqlrHustuZ1xozeHt9QYpAugUTyTBmzxzSMJU0eheudTmJga
VfV7/vW8UkN4qHnr9FXPTyt/Cb90YWna49q3wYS24x2q56OzmJj3BeCkF77Fq4U+
23lZQ2OVEHmy6nR99Omrb0f8lgMqrwvWcEW5o1Zuc59XJ5WY5PpORXm+a861QhBq
gwOllrDAbYE8IDXgzegdf5MZuf+OAIwMqna4sRq7fbtYjNtejKT9ZBKcVQdLRs38
5aDMo6OsZd1r6p2AaC7bYSYb/Xoh8XOU6pW6XnXiWFiqNRgKDwqFtYf7MK0QxxKW
vzTjpXzJMtQN0M/I9B0clU6A07dQheundw4Qs+2aZ5bRo6YKE7hLuNsYbHN53EgK
3EKT4s/xS6a5OR+5tdNazMzKP/tKF3YTUp38ohTsiTu7BR0uGtVPOHZVeh2E/ljR
EVyG4Ns9ObvDa3Wi0uo3lbEpK7xit5KyT9FLR6tEd23xEfzdQKxP/5nYaz3NPmMc
FUy2SwqMlJTFZAv/pH3d3hSvcvgRzgURXk6XDeSaFDZI8CmpNZq0M6KBK+RDGlJB
QGivbwbJvIaX/5X58I7rG3GnRHzJv+SRCKzN7PwmBMtGjrcF07qcJOxxEGZaajsE
KrKXTSf5CpSZI2KqX5QDQ1oObwIqiEWUesVK8U7RZL9hiU4pxbr6sey8lKi6rc9B
1Ex9PwenyMQIRwj1M0cT3oQJX8ocQUKuGm5M+9CBQCtVjb9J03Ft1tR1m1/Jb0Ju
OQpgwpSrx1wNwsGmpz+Ik82OCzZG5NJyINgunZgUWj+0G+uJwddsYMYRV8YpqOK8
84hTXdbODnIu3YZuMzfJSbZVeEJojJSCtc1wyn2UuXOvGyRSCPwcOVoy41QU/8uV
5AyHKw1LiVj0K6Nk2JFu3oqVpk6MPPcCucv1jz13UGdqTON+Z6zk/3pH9FlP1VxT
CDrhgqF55zazWmsw0AIrsAZyDUNtg2BGjODZr0OU+/qryjHeV/CHa956x6rhinMv
AB3vqKLGP4VB3Bn5444nP7Lml3NqZqT2MdmWNwJoOaHHlPSbCvCNPXiDsbIsPRWq
Ik3fNCjFniAnR9t7Vf8rg8HMda+84/TMTZnlPa9lj8bqLrQr6vwBgZ/oKHnZN0nU
Mzn5cb2GC1QlRZgx4pR2kN2X1RWlye7s06xxUO8UNARRYM6kUTVpG4lOaOiWVhJ+
t/Y1pr5GHHlixcSxFaGuNKby9RVyIA4Xqqmjg3ZS+0VaIO2x9d5nTGb4E/Aqj708
/0qNDuCAV+7NgSdz2SFvJlAUTYVUSQWTnIyusMXrTZDTaKekDB5I470gPPzUusfW
6DcOSOKkTNYyLTLimdl/e0Oqh3aZ3diuHKpBbb9QT9bNzEzLazeclgtTmVsFZuMb
1tgmFyeOzeDNaoslOE3CmlZKRDVvd0XQeBWvTMrHsqIqpVxmVneUxxibsTkrQxtS
wUw5MAdoRRDEgIV9HJGbDHkiw3P3+6zpDOvkF3q45dVr5Ng9VFa0nEVj9G+Dl01H
iunKtF//GB2fXgJ+vxt+O1/Yl6KOsFIHxyeXjE+wUsvC5ic+gQEZ1mwJfysy98DN
FyVZPhsKHAUfRqyd/O68wfTyZijUcE1ZL7AFxSFVWNr4xicfNk5UpYdIu6yKxAci
7+0GymVtLPDyUNiRkLYDdNUKFk+NKVRP6Fq4Xy5gFO9Fwy2uW08o68DS4yve2Slc
VVePcIUHO4kEuxaTSKfGmC+qGg7T2NdOmiPZc3PfOd7E/eqi01imIcWSmHN08ZBd
e3UzSBn7jOZa7M/lOLQZ9gd4PFgzXP3q/5GLduv7Z2wgiU/yQF9GCAHAmjzcjHTF
xitRsnztal2Q2g6r9HAzMH9fV1CKxZhgszqDQ62epcKW7MTVepon9uyKG8Tnu0ED
mwj8ZgpadQ476AtZd+G0qQnExKPguOhU/jLVbmre2x06MJUkE4gadGDHWML1B6nz
sXxCMC1cl5vfTCT4F/7TRHV/IpyXdxnVbD2vul+Yq3rQCPWIYpihNo5H4MEoIjOW
mGQgGbjWJnYZ1a8bLVgwJ90hE25AIefyoRP+BBaCjpd5FdapX1kGm4Z1Z1tuQoAv
ODh0F1uPBEgHUvpNDvYEW3ZGykdveKhXWmC/nuT7CDdHHRXFF7j7Re5qAAzK0iAJ
KMFPRhVkAVS/Lnz56DdYB5RPEG/+M8dcJt95sRIw4O56o/wZIuAFAs0wcnkrgyeh
ASyve6SYN/q8zoeFS6mZr9A3XUs23FGj9ppqRw1jo69mpOdPP40Q6jIQgaBv1r41
5XpnbHn3CsOAX2208rCIqSTXBtqxQ1QTzELCu5Ky/TqejeSbVYX3WZfmjJttGCBv
eXn/+otzNVNN5qwEn9PSzirWhZFa9UgY3VAG4z1rj5mXxEqnblisu4GlYEe3a3p3
rYIl+wRAQd98s5v8Dbv5Ku2oAo9rlwPw4v8IGFUbRFUWQxF/YqKBSxmCMlMXQ7m0
BcARpt05lwhFyDyq1F49Qk1C0StvhgdMpVecsWEOwfCtCuK0vxbKzyXA2hnqkHS1
NX/iDwvDOeE79fYKMc7HUpvosoROlAPxOsl+6MEsbtsR8tk2DHg2xg5xJbku31zV
ONFgYhFAeLI0rzATFeipDadSNbT5hmXBmmBO9QAxavzmAUhd7m6RYVo8KPfwyBaV
BrgVSnLuLVdfC9a84LF0hXLCJrgaepVt+0eXGkyXlT3EGzbX695yJ/m+kvLMtYHT
RBPnkHg0YxMwNgDF9ysxh8r2r+fTmEPyUnr8/nijaHNE0DQ0K1zQA8PMDmMqpcVp
s0MZOB5e4jtSLOpmEph/0d9Gmyj2366Wi2t1UMJkEqVzNiA1ZPbITsX6vguQLLON
/jKY31nSHUnU3YFKkXhf7CBFbhWKm1VxBuKg39l0UBrez+hPiXVfkqVocomQ9P9k
0AycH3qLmGZ/oJcLuQzTIx4rrWS6t2m69KY8a4n6M1bOUpE82XpZLEQ9ICevZtuj
k4d32XbuMp7N644qQpfbvgLq/s7oN0e6J3JTBF5XxPiXMLnwuS5OWBvjpSye9bte
RmyaIjkLyrmzZMdLZr9VhkGl+Usm3RAEzuodMBiecnBQhTt41ZZJOC3peyG9SaAg
gt/mL6N6ZsiNxDd46oopB4PJ8YQ+vZoH3CfVbYjZOLq0h2rh8vTAhfYXwGbCnPNM
KqX9sQm5N9uP3UdcMyJ9xq1uxIaZ7VBDA+mbvH4+xW9gV+fyYJ8udG3VndhOuIt7
mZ36UjzNH8OyfheIuz7Jk3Cuj/R5d5xsB3Dw808pTyW2ZAW80IaGT0uKi08CgEiv
h7zZvxbSvOEEC+TCv6arj7EyccMy0R7z5YnxP+zj2cWQYYCx86R/1GqxOU0mfvQH
Ymlf3zmHCoCHgJEYBYIzoLrcZyfsXq5VFKvS8iViuOFmNaWgUAZY2J+wI4yycx2l
lGeafcHz/umdDr7hia42FnPbSd4xkoVg+OKT+gYA7I3qfDaYv/nLRszGPGGea8s6
udHqPlCtfUiYlrN/8Sf9XVuXNmPN6JfvQDVE4guseg7EZ6R1xswrimYfdNeEI05n
nMk6p4+JsehEOzMlgnBIzkaDftEy9zbFMurIFytC8YvRzBAq9GDt80CUCGTf+W4Y
FlViIQbHqfcW1QQjl5238bzldYdAqpwBlzA9IcpsV4d9vzYW7GbbKuCwohYm4zLw
0M4d8QxnIiy78qxE21XapE0ESTSwOytqz11/z6iAWmp/GyaVP+YfMU7N3MTi7DV9
ETkefBeupa+/3BSPs13kjKlZRHWh5zL8EwWhHLVtd0S+UbCHEsQqdVylu7uEjCGT
GF0sAsR5uqT+Cf9+V0VQi9/nMEwDgYDDrYJY0rMw7hn6zmEo4Wty61c/GEskcAO+
AblwAso3rnzLcB+s5V8/OhdldEMD/ZsirAJUAhwPkrCpCm/J9yU89J+Hy01zvmA3
ePvzH0nyJn/4AcZ+3cmUtGC9qx0cN183BG0e5wVQM5XBAsicHibeH4FqPuypm5Hc
ABTW56TSigWArpUTshdHrBQPluUQd9MrqRnvO0aUQ01wQsugMtCWWf5HVtWZYOUQ
uRS66j4cPVLNOOkeJLFY/EhqhF45IEKVNXWBi9bPVOKq5nsEMQNf7Ga7/1cEIjh/
IONlZNFgLscrthrZqo9/aDRFWDuL9ebjtzmpN91/hGZ1VqWvliltEvNktzkqj7b7
4O24viB/d9S1xnkIjElgmRuX/fO9Rvf4dKTgC9iz1gjGVX2BVJFCN97z1Y375ZbK
d4vwKnoTc+3O9F0owh+u70iB+4rh/4FwSXPW6VCsyOQUsQiFil0ziKKEf5niMt+Y
qvLQ/pXXfqshmKDkcoeoD/E8IEmwqE9o0BywZsEsteziEIGXTPkcBN3Iytxmr/wM
3sX9dWo9ExUU0MkNrdxECAR/p9Wm8IfULeU0yNfO4WrbWVkn49vTKIon12nh+/cu
BFE7uWFaOPm3wzsP4/4secicD+cSPsIXLJJIHec/zzKgohKttv1aOVjL4GF3T7G3
g4HDTeW+Hzc/ATT1E8zdfJ1hvJgUnUZn08NlIv9bdzoLe/L3sUFvGri82k5Ib4K2
YVWmRThIA/rPmGx3sTdBEmslExiIoVThF4bNM+S3Tgq2vo1DBDN2OLTk2QJbOk0J
FedsZSfKOFlFtlpWHvtgVuLl+r4Nov/aib8XOBCn9M+L9bGjgSg4UBmsdfttb9V2
wdBN5S0ZUqoiI7chZhIfqIQm0h9O4czEP8hEpKqQykDXHl15K1dXKYCNme1T3v0a
ZKK+KPdy6or+KLGTlXJ/fJgjt66bPxyh3QwuZKyjs0l2GQ49fqP/MlOPvqKBzDOm
x6yV48Q6JUJDoDpIsd0NkCwBQCaR/odw2rOwpNddtYsX0WUdlMf8K7C35c8vLOj3
H2wip40T3Jm4Ba4mOCod/30PcyTWB1/snWVJBpWJVyTdI0q9EMeK7q9RjBsFFgzX
+W7c2VxS41OLz0Sxy615/KeEUp89Y2pVQTlhCoLkAxpi8er4QFh/eBAL1p9timx0
aOWkkUpy5+TWx1HO3p+XF81w4QACkCCJtyynJc9E8LdL2Vn/cPEXKqep5P2/aHqT
Q8nppCwFdyMS1288NqaUF80IZO6H5bvPDNX/zpJXsIH7VqCDDLtV44A+57EY6xwk
JEIkfL7J16nvnjCW4seekTKxeelx1KKR9NMxIV+y5msRsNAAVWqdyhrbhSZoGwhk
E7Ku0qOvrkv5RbW8lwuvKcMuTHV4TYKOnv8uY0MzVWnNz+DKxIVukfAMJKeY8aEF
c+e/MufqvCJr2aIDdnQ0zHL3i8rg0VOrtFFZecYXck5oz2T9hpk8S+ivNko5mnpR
3OYvI0YA9OMUtNT9l7T+7+ua88gSIxt3720EDD0dJkAHwcPtxsJMArjCrhSEmSOG
rd5nGA8Vn7TgBM0GRuxgVrXJSIFQBo2nTs6Z007PoUC/2ymHcbTXasmlPZi2vtfx
QltfaHctDLfZj+uY7bK1CYpwNN9ZTrkwJfnFacsluA6BOK1Do3+Nof8cOz52lPHc
5yBOhkW0KY530FSJdzkkRyKk347tEQWXs8eS4z+MXsaBhZGOpjxzMPRPRrlMY1v3
tB9JTzfJ2ExlK0MHLhLMKym6lVzl/3SfWve2VWxUDjhIvR6qAwrduTMRJU2qN9OH
ASvoYkc4jsk4T4AZruTQj8VIQbd50aqFf3RXKz+JS1KO7Adu5RUPkRz6yt3zGY+H
zgPofI8THkHyOUt+jkBKdOj1gAkgi6igmp6AvtHNgaTbR80+AjIpoSOu8iY5GUOE
FUc3uyQtjUhKaW2BYBamA8SanJxQRTBpt/4/+JX/owvKhV9j/U+hSpMwGG8WQIKn
8xHv6Vz2Iu7k9bHec/GXY4lXtZxGebZ2eC0APQYTp7yyEaPdHHv0AlnFxjl4Yb+k
AX6EYiWVTneYSBPLIooqgMgI7za+lX/kCqZun7000+/NRhwW8iQaqpU1jKPcXm7i
v+py3i3V45cxSxN53hna4N9nNUjZYx4T34eOooImUxBegBSIf2Hg2nmzhaNg73VB
oaDkhVIV2Xd+BgCzSUUgcpHJyvM0jJAzQm3tT5JVZutOZI/2YA6GUe++KKaaNC5Z
szeBH7Lb/uN+XQXksoJc9++XX11kc3/DA6Ji/wWTQ6B7ZjTQaJh3p1Dtrcws77iu
hw9Dwok6fKwW/n1in3vSu2HFAPLr9ymT5twFrOYz6/e8Sp+ZzsxQp1sOhicsGtr/
cR6XGo1HidzE/nrvt2P4DUq0tVr7vN01vb96blaL8XsaFkcwOd6vuZti/amniRxE
Qc+QvbNncMdgdTloR/DVRkZSa/e04VNVYCvTtk+6e/2GVNc1IhWBWU2tKG9maiJa
Bkqy3VQhQVYemAON1v6s3u0tYtvzzxmkbxUBeLeX5/ppLFlFNOI/aUQUHNt06n+q
mBjG8rP/zzp9VzepNV2hfA/IR4ihDXzZR0Dm9lKFqVFzELfxdQhM/emAjfXB1p6N
MDFlabjIMbqWMERpwAkC15bR1AuJSMoliZ6TZkDFaNzjThtqz4gTYDR95V8VBdJ7
KX4oruA/XcVeZitwqMANkU3K/gcaBbyjTeFfLnHOqgxpCzyNC5LvCTlSD39N+p3D
kJmDoeSa/7YXnENVZVoaB7Eqvr5xcLxmPHJ3ql5UIKcsCEr0NJ46vMEpm69fzSAO
9uNMj0qWByE2uquU1JeTPvRryrcG8Aap8a5aNAo7D+e5G5giOZZ5zUD49Y/MQpoY
n3k0t80OhLKly60lMzdy57fREZvMTfzkr4gJLIMW6Kk6UigxA9RSNQqY9mXpol9o
bGC8fsAaSxZ0A4hTkFtnWHXEEZeIkc1nQpLSLgVyF/NHFimX6m/ofed/DW+4VrRN
lL+aN7lT85WZfJnKEybh5QV24+n7NrtwHgj7M/FfGtfEXujIptORD6BTuyHG8cr/
n2oErLCX3cvvBPqPUyV23tuN6bdM9BOdhOXoYMI+K0kItoBEfadUodSqV0WLgvaL
OZ6LKt/fTP7rHkeE18X/tKKyz7Xb9WF59znoG2hJakaI/KFRBl7HiYNbBPN3Lqv3
3QBCvSsOUmW3kNUkRVSBi1XljVIdMf6x/X4emiwaht/t2wEzkJX0/Bc161VMh4am
vsH3TtlvlxH6V+5MOEAZs/wt4l9IasOywoYn+P/yxWUIf5/Tpc+FHzgbeIGNkbVt
who9jS7zb8VgAKy+fM32D0xbF4r0HTczvZQViXp9PqX9X++v5jMQikGjQij0+RE9
D7hyfRsvd5OcQXwdcyg4t0/L8g9yveQDiyIKs5Qa3Zh3NN258HzV3Qj+dLJy6dVL
LHNYt+6EsBJgIb5mls1qO6db5v4bqZ+SOhIl1qkr9KtPFi1r04A1OvdcvRB0i6PC
QkxBfBt7JkZwpClcgHZ90FIr0hBnRsYN0l4+Bt9PDGzinpkN8KcBkOWrROUF2m6e
+D13ri/MQbacS+njV2c5REUYG+rCkPdAz4GmIEh7ZY75uCCPehol8kqX60MkPtvQ
TdeqQB6PPzyCuYOjg0esTHU62wSUMMbVI7JD6hAfto1ymGVoaLIB78r4gGoOaM9o
HSNxTJtSzHN4nBBvscDz/LpcLqkTOA8CekX0agEO+X9mGXBl7h7k5j0EM7e6XZXt
FPoVp2wj62xd+Yai3OtfS+w9/BaiRjWzLcRaOeMoFLxONYweFaiv/KD/FCCOc69I
qzOw9hFn9/PVQhsZdH/kdDpDWPlBdWPuYWBhVcw3Q7v1XkUU3oLGZWzdaIbeZpMN
B27R6G+TzgzXNdkkSsPu0BFdb4jg/KYYowBKK4q03mjhF83gG2NYJNiTMAg405Dt
S9ThDERxP4x4ojMNYErybYJzsCOssYNhto/rFnsgvkYZJkl9DhG3XxfkldQUilgm
FL6PlyCnP9HH6AeJNLFOxEaA/fAmnN2UwBKBLFK/e8ZWA4ZpGVo0uG3cqyplr+6D
wTcKbwmhw5tXf/1sLFVDSg0CCsnukDeAATfYoP6vI8BpPAUycahwfhvjselHlPKL
8jJU87VE8mwyLdoq+pJ5iof8r5ACJQNFfwiZsOQAiHeJP1m86MFKF7ar1hz66haa
U2gTTffHw3oWq7uAn7Ej9yDTpiqQ0+aYEsfY5PuewuTbu962JwJXeA8xYrTxkOis
LBM0pB525GI8+M22LWQ4S9XrbiGFLcI5Tx/0TBSk/LGCAjhXny2qf8FTBlyV7Slb
no0ECVBnsOc9ZyvXdQIEGb9A5KpxfVJq09BfUSDtfu0XO8PRMMoQ9kh6EMAvVy0N
9+ZXBTJaFqw3UieZgeCXEbu/FmV2CMeFu1JQghoD+t7JGOpm9yZYW+45m/SLNfBF
VRpU0op/lNz3m9xTEIzXakykPELFWWyy7uJiW7AHtXAtpphKQiyVd0PMuQWnb60Z
MMsquZP8phH7bstDf3q7qc2akndlijn/DHawTiOcmXhJhJlRbfTgJsnq/WFfqb5x
B/oOPgZRJwHYHNf5Ku1QvdXFNo0Enf7bZlrxyGIqpA8vopAOIid4/aOrycqD9ODN
p1l2+8kffBex9XXA48wwXVpZ7R4oIkyC1qJherTjRJw80GA0apZeSlLb3CskDR9x
yjC439D5p9Dk62KoUZN6Z4lCj2jbvvAOQUHCpc7sZT54aNjRlJKGQd4abRKuVXEl
vWddDkFgUFbv7C3qr94b7MGA1X7jFCCEjj25riWyzPNePR1Ycbo2bck/qsmRZnQM
QUxuaZIe/25B8AgedWWdXgHyf+cmuELtx1Srx9l5ezmoWxz9UXz0yixYDkFwFrJ3
6xJwjRYOaI1J91Ok6ETB/RyFzUWQonkZJYukIClpqWr4sb3Wmcppx4DVHKC0ZR3N
2odXrADz6ZH33GMtG6XBYwE5Lm4ap6SLe7ZzdVzwz5y/p2x1alhfk7Fxb5ghroPY
aLzp4EqE4noUxHmC8e/oZbEcGUE8q42HwIHyCzUMxLxMQhWO+olCSwe2WR6gBaQe
7MTfSzLrR5tKNXeWmi5YIbhc8wplEEmEOpiP+EWdypMUga3lfACNlNQWMB9GlbGn
VI8iQs1MCU9sQsSXNT1v3fUz8cwioyJ2ArYOib2EiJtMbTsq8Q3mpMwea1hxS3Lb
l71gyjplIV2AIye68CQ+wlB9wSDa1fr2/b5Gipo4axaK0P2n5LDLDlebN3+erHrk
T9naCtMMiDWPQVu7zLxFFdPgtk1EwKry6JGsoBCGGDIzVnJlF1lFQsPdSfxObYrr
FN/6+3O/19txUm2l6A7KstHiXC7s5rV9Lsjg0UFez2g2Qbzb6I4iiALKvmcZOI8G
vX+BxfHm+7I7AR+3vn/47NO8+Q2GeBg7YDrFBc23dSRN6Dt9WHwS9IX2uKeV/f4u
e0pKlQN9Z6NHEeIzI7k7wH88+KSpIs21EUZJZuxWIZImaJW7QnfCoUkFDNK8h5cL
toENK4LFZOGO4kjm/pPmoGtuTUpEUDcXo42uoQL6OuWJrbbc9PEQTBPHnDxSlDl/
3Pq1BEWSWna5cZ/1ElZVgC5TS7M6RQOVATMmYSV7WFBq3drqyoNvke6txBTAyTRF
cUZGDYn3aee7nbi+6gj/Ryvpk5+85p1UmMlOF7yHm1NYMLX0iP1+u/0353lfROgk
ktQn4+vflNs7lt3clk5oO+OX4Q8layA30FB44O1A+WKKY97Zwf+Z0zVhZ98Qp23S
jNYjKSEhxcq+dwDKJaQgwVnoqhQ5OFjN/bpXqpuBLXXHPnMmP+AxzrIZVPKo5B/k
4mEm/axXXOfJpoXUMSWX2GzvE0tcDpX0hjwueyHe0sjuB+wHXnG4wUBYu53R3xNO
IyYqLjUoH7ETslrzdiZGk0XRYbxSwKmobfQu+FgejF28xoCuN8Z9+nzFXNzUS7Lp
M8MZppEwt3a7R+4/QpnaQYOrTM7qp+7SJJCvB4qk9T5UOhqxOO/0595z+L4MC6FE
rYeRyczwNI5CLX1YPOFAPeVvOPfyi1WO+xe+EC76XwuTz4qSSSIUErtIfeu2j2wV
Wd0aDAu46hDmqgWv5ySzbMKJSIQOriZ1gUL+StSwDj5VVc+gEzJL+qU6FHwNKfSn
rvbaeT1P2GIUi0IHjvYOTDSAANsOIvdtlpuzDMicpp9b11jLTWU/0snSZANvyV+y
d+6kQE6+yI6le6pCEj1sPE7Xhr07c0ilK8qLYzIzZSa+8QHiZjk4iN74RsDebMwj
hyfjn2Wr23df2iTHFpzovzyj8/LGX00t6+besO8bJBrtMR77FwvaKsrWAn5zL8KI
BCCC2MH4Bo/5erMBkvOR5oX5NHyGy/h7+z+RmuvC084qmQAw9fIsZ71U2IY1eGe4
I880/7VbkRfCfjZFnzT4PGAuxbi4Zka7+FzBFaYbaY8Viz+p+rtRsDX3QG7XcXjO
n03XGVs5+HMw2s5pGx7D1o14EPvD+trUbNyYDKjJ+0K7L/EPX6byYgCq2o62a4qb
zNyfVnhRRZIVBBbsDbXZlusPpvqVYObSipqBx6VSx61jAZKr1N0E/vnTtEh+Zac0
QukBjCtQFA4ovH1oi19FBAuwtumpJQFwkTHkWMl09QEFdPv9kCXU+d6LVwfXSqef
ZVYgEXBMM5L45F3nlN47HEPv4qSt87ge2Ga/QM7A1hiDtf7E56F6gP8vzBVCp3i0
7LS/wCMxF6IrBsW70iD2Y0URkHhE+bzWHRGeW8GqdDMR5ACohOu06eiKkl3ZwZBA
fWkqN6jXZcIURe2+2ncuGtI3ZHI66sVMFSkCOcteS2KCjfN5RF4wYwoiwzxPfhUC
5ySAizrWp6agf5KMITHdFNLcCvgxLK1SRRx+GpLisYuZ9jWUT3RM3sboM2MXQD3T
aJRRr9moKRw8BHk4usFKQ68WKrKmcMGcaZj4uTef6NmbBTzjYx2ULdLQPCqIUL1F
Q1VeQ4GRqGaka4ilAGT5WzAb4LZdJOYKAsc4AKnFl2P3iosBu+yaDr/sD4DFUxd5
EVyNWBAjVs0icYn4/KKsGMrH87t6HHMTU+c8GSgPQZD8skYNpc/PPpEq7ZbLc8w8
PcYSSLZa/AlmST+EknTc4vBaf3skeoVdoa+dqG0Wbkfp6jacI/jhHFdOnO2eD3ln
IjC+wnoDCsp1zL2KS82yz0TwATOJEawCiKxYM4IVjtZLXdCY+dInSSj9Jc6c+vOi
O6H+8Pi3rbFlTcs8QdDnq9lH0PQrm2FdaMKhSTohH63AfB1pn9QYFA/Wla+bMK/7
r6odG6R3gGnV1y/nI7p/hq19AtV+grg6N/Xx0ddZBlg3ZjcntQE0aqD9JoB903cB
e/DyPJs4UMIfJ/g59zmWdF46JT2mQQ9fwbb4t23LHUGvS9XSYVLlB3Eu9elpsDnc
LcGvrB7WkFHcvcawsrho2i/h5NNxPEzh32QNSYzlvlPUJ4kKRArLfEpJpGpowdSy
Ropic0FB7hhiO+f3RBKi6LnaYe0G+A1lwFnYwSNna0SfhqUoGTtCldY2Se9qoUzl
+yVRpyGtRz8UHITzPskqNV6EY+soYjyKV01cNiUQ/8KWoaqpiw2Q55QGNxtv3eUj
mHcnxlHfPCW53PHaUkrT5HNG54VSTgwAlu6hTRmOBVdt7nW1FMKYfBqg6u00wAoF
L8+3VLudhcP/l87MI3i4d20DB8b0xWdeedzXUqdXM00koyHRLCn//84E87Ya1Ygj
KVfnZd/oE7+uXck8tMDF52SXl6o1wDt+xSh+XQhYd3LDGEqk4CayucDP6mpo9QCi
S9p6Gv8McMlRWzJSjO4hPpb/s9cBf7HOddbaAUFDRMDnbiz9t8qJArZur3LOPGZf
oXDAYmsA5PW6iVlWMOeeOGyvZ9mjP3/rBbstHngUFwEz77aXme7qAHhFUQGApibW
HKYDNIyuT66IzgBTHi3RYz+r+5ro9d6mR7U6QGjhjCb8yddz/2X7VLWaS+bNB9s4
/eLNp5D9V1V2jqT/JuBODJJZvoMAigBNpeYlKIo9IIQ9PeiImrFYhrbOTxG+Gkp8
Q80ixAOnQVjbJGN5LjofJyb4H1NqDkZp4urBGVoWjLby/OoJdKgvS3C73ntdZ7xy
k5L7VZSw6Z8cUE8OGUb2dv7k1bFpyJa+c8bQ63OlmRfgBJbcEWJMij+jHc9JNssP
CZeiFQUkDPBa1B3tC2pVeL7IA7ZwSw/cmE/C+wbFX2jA/3cKfISvU9GEd0yq9rUG
9pnxN26thyQt9d+5Hp/DoH6OHaFymiRB2i8sIQbgkZLm8zGvFj62oIh+Z3U/x+3X
LyD5Fw/dWrvl+/SBPetzP1tJgpicKz3e2ret2cG2LW7gNABCOgbV6mebDWdwwGtE
xoDWasvya6SkyrvZB30VGkpg7vFI6bPc7kBk62em+RrN11M9d10rXFWwQpXVK7jC
WtTcc7UuPXUgoCwBRYLaQSzeWNPdVWUldooIy7/dVl863IZKt6t9HPDYX/IHLsqi
zcNgNopWQTrRtHZ6INzPXR3JlEU3MH77iOnEVLqX6aez4R/M3YSnU7OiJvKVKIum
jWWud6wUHyfzEV+OB3mi890s2WX+XCfprpNkoI2NX487jDTrR29fDVBMsPRcfN/a
FOQLTNAP/mueVh4xZh8RNjKlOQIWjxyVLbXdavdhtEA5CivdMyrWul9jIv2kxgsG
tOEuxdPzgRQShQXT/5dIRX43D01kvSZXQZ9poM7jbEI4l8vTfDeU1MP2Ea2CUltH
vKeKV/xRvypb2XYmbK09xjZgKQLsSeD7o2jf6nQ2oJcoZ61x57NrawIoCcj5ovTb
j62sl/YDqlmVWIhUebMKf4YLhHOO4y4XR4nch+K2w0EqsyRDdnqP+YJOI5+7lHgZ
5zUbEOjYsFYUmA3Gu6hr2RpQptUsKVmtWZlVxLWA1kOrZ6QEaxc7n+3PgbdnXC/U
hssGfz/3prgKJ4AFkuwBmsOVtZPypVMXnlCsD4C9MI4KWMCBo9G5xCGAiTBaTRBl
JL9Asa67PQaOfvqDzfApL9pIRMGZyKxhgHTJS0c5nom0iURm+D1l0faWMojcV+c8
Zjra72FaIfAKPUH3O4FocyZqIsexbkH+egJv93/ZZQtsS8diUQsfoXYOdwRq6abb
iOEpHQRS//dd3AX51x9soVcyM5IhGnm6Uwd9DM+n46u0wQw12bKpYtfk+/Om15Hv
UPk4uRPvNBAm2MinWGStlSZNdsmH/ITi0FI/dv98rTXFE8t6BjLrNehSGI9LBnbt
HdCqPQNqJlH6WwfvnvIbT7HCbVoFG7eS7K5PoeaYJGnvrwOezVtEMz5sgLhVqR1o
/IL7Ds01N0f+BVrdBRPkU/P6oUPpO8arHxri220X3MrU2y321KKgw7TGVNj2QYg/
PyQHfCmuV07KXGMP78KoiQiJRSj6quiaUgLeIq2nU+NtmFyx7DU8PpfIBdyILQKX
08Qj5h+e9/SCUWTnmwl2Km34u/gLplWeugzL24PXcOU0fhUx74C0JVPRDD8ziZOl
6SWZEV00ouAAtDrP352qpJafHy5kirl+fJCvh2IaoqXQDlOR959N6VSIKDEOdqy8
un91UTqElxK2o8GaAT7Z697xdYgI6lTeaVhsSSRbNVBi4RawvFlnj9DS4UrfGp/7
PoxIM3EYu+kUiiKbhxfAK0hhnXrWLNvuO8xVkiPGthYDJkTuetHNC50PFvdhkdKo
GoTdHYwb29zaXVzqK8ITQWVjxvIC8DrD5kWLYQ+P4oN/f8L5ay72ddzXMtakTxCR
CtwZFG5qgr4hAPxoS7bVfEPl75bQHluhOgvCORx3pHaP+r6Z3Yygs73Uiy2TVeYI
V/hF7OBNtOI8JRAo8IsiKr9dB1tzB9szauN3p4fFN1sB1PRjxCj7fVf/UOfpBesI
LmBChB05TWiHDmS6eXrG/KXTXcHQ96QKQ5ZdeS72UPmB5lR4ju0rttciisKprp/Y
PxJZoEChFJClxU+yrFjq4LObJsNGjiaUQZsXiOa09lap4V6jWigvoE3VeoPUkdo0
hD5Q1WI/8j9juKQL9ayrKQL0JQsrU+3jCR6zjhE7MxS1uyChwmrAexWITGG2yF9h
a1OTNxV08iwfXJn/AhUrtgf/Yaz1JQ92Xn0fQKY+fYH0fxg6GMl/1i8XNJ5OwjRW
F+RoEIOEwo8M7Uyy/iJSf6ifXbtvaGS//jU3j2JzOFcXfwZOzykUwxPSrTLHoPkL
ei+cwHMCm6FSWvKvhRS3gApkdowc0DOvJBIGxuf1bgb65TtWwZPsCcoWZz7GV/CF
HGjwb/XiCN2MZ4W92HPwijxDdCiydYruMYUKpjp+YC6+08xDxUQFB9YXe9tQ7yRu
lL5/LaS/lr1WNKBHPlnlP3LQ8q+tpoa5kYqh0SOq42KxHZBYppSXoMMr4+Ce5bUb
XjTC8cP9KfNmH1CXLObQB3elgHomyAEkFHgMhefUlNY1sIUYwhWa1HZh6kzNwzX4
m3nUwJjKVXMWTogNV3ZBtAIqs910D3IZRClOF0BVEzPtBpFybThi43KOLexswr9G
/7B57bM2X3Izl5MzfalXSHuq9+o3mWYAg/uMH2Qtq1jkROdyrUKnYhOf/GeJmHV0
qeYgfeXUrAXfk7OHFeOCopdCuqW84gccyB4A/6BI2fr1wTQQY73brbVbl+Nk8zBI
2Cs0zNnGjxlONeH0Go+xwLKOGpFQOdU7QDozRMqnrJts+IVg+K/TQy5eSnEk+DyR
CO5VNRTkgVR1tlUON4SKGgH37oStMSoVnu06mY5TFL0LrJRkUCRIo0k/Poq5Q6+x
hg5MR1lF96e/l0wCIzgT0dFQmxDkRBBAadn/S19sYZbfRCd+ARyOWs92NummZyqN
ZsspIyt4ZlJCGV+q+3dIvqgA1NlKT2kUhXEXMZsvK7S73VgGNzv6waezpVnC76AG
9uMmyb1DSFBLl6OlRFbF000A3IiR5lySYSJ7DL1QkFidjEKzPM8UdNDCN9PtwzIG
y+VsJ0U3FxvYDbtBZ6BUPLgOnoeDBGMNidvaPOkUDBsRNZmmLsQevXu2ykkXk9Zs
IK0FlD+eVbRJKEe6G+zaMY5CUJY2FEbmnXclcXa+O6ir7dSpfE8gjZijGuGNQwvi
XNUQaBqO5oPDz9iSdWpG0M9o9OL6VY4wFkksF5DWf9+p1QL5IU1ETXwY2XC3LBvl
G0zpj/BSfKf6eoc6T1I3zm4KCs2sVkycRVTmJyNmgJVePEghv5iuproQc+AqajvU
ahpsqbgRbwHUFhq1dkYEAb2OxI7C8/OSEbFneqWiM/BmCM2H7VY9TmliywwS17sT
KJB8op916ve54zEJjwWq2ZLFQJ2RKjdZvdRmz7/rCZ55CEQNrQGgEKKNUK3UsJj+
azD7HjMm9w8777RIsO9Z4iekf+OXLPvVz/pttgXhJVVHBBjEqJHZR07BVqvMhOfc
Y/zVsAMX6puZw0Bh/00OXQDjsoSkqVRmgp+yO8yiVDP/ftsqJ1nM4WcZ7KrxO+5V
4tgf2CJWej0blAN60hs3uzcB/IqMe3GBXNtYXW/WpI4IvuYSO794W6DQp1uCvIrc
fMz9nkDLYZgSTIENYObt8HIPcxZNhLOpc91yqk74Xfv0XbNdt21OogJPkOuTQ/3P
O1CdHrOwwNgghfdnI6rcv+1emFbfEE4uNN/LEh2IksPPP01nhc7b+ynZ7DtgI0ge
v/5b+UiSmmZ0FEK6mk6nNPltCGP8d3+qYRQzQlVT9qibQNUivof2dvby+uorZqkm
2e5BqHQ7DbYp3akzoKUkkK1+qa8DST7z9FNErSmibahAXw2s8JV/3XmtHXYUzC7w
kfj3PEWMdlWAu3neZ6BHKRMX4+MTXaiCnmnBa6FU/AwkjVNXi2ytzBI2ocr8e3yF
a9XcxoPirGebsGnlBmLpSo/GGO8dhqZ81hxIKb9GwmIMFNNtreGbL2I52MqyxBss
p4gIFMngjo46G6IgSXBa8bylB4YTxjOgtGVIDs5qIIlJdk8hZed1wzWQCUj6xQY9
c3e2N0fg0nuNtHDm5mFxK8d9lO9ZRjsaZHEcphP0/Bi/Ca+UiKCN/+IH+jkOwgbH
uEgwgGvtitIuTy38rUDRPqdgpkqCu4dOiWWc2OsyLyK2s93ZFAMYnz41zTtFa9eT
k1pD0drnDLt7XGbxFyiMzEybmkF9P55Tu11KXf7jWpfNAdxRcqaqdTIt57G74YTT
pPn14AIBGszyzfHl1mMqQ4aVeRZgDFdwmNfHOIm/2JERpf5GFZGqgF6vyrwzvpVt
e09AsD9DG8sU3bp4MHuMJDti5kb/z33qxdGAphKYcOfSNPgGmGM5rpytpsq6sVw8
qDtsHi8HeqKwHXJewiu5/aLCPKHhHt2PJgN2RIEUU9TJr1jjUsHqiAHn6R25Bvhd
iKJ0AM/NoKoGt5UCRnMQN1WHGGKvls+RIx411us5v+HmFBld84UJkfZvgsuGNts0
Ren8I1hzIOlNxfqmmOgRuunZ0v3iOZWM2Un/XWwQXblwUCGcviBbpoRvrihkwLro
8ZUzPUF26oNePegTMnr/Np72aVRiBTEX9zjaz0+6Vr/dXKT3Vm2Qz5wdmspPvsPF
I+laoebbbCiHWGxmH9xcgdNa/pjZeTpATQbWZpvFaSQHM/D5rtQleGMQz1coJ9vN
PEP4e/2bL02QGQCCTED+fF5uuZJJ7hTJBT2KtmucB7FAbwNXO9/ZaztdZN5kt5wt
pMLNVvHflllr+ghHdXoyDcekFe0uWwPjavFvyuotnHYiGSIa6uhhak1q4K7IsfJo
u+d1qZ1wttWFnc9YIkcyB3BOHOYDILreO7pmycqDMke6LeopNXq6KcdRag5OeJJI
/cnIVqiHzlXAs53C9g34kxMeC4UsP/amz333tIb8rvv89vqBSoF9VPLGry/6COm7
rSusLvx3bY2/ZyKYevflFRXaMrGLLMaTdoxX2Gfeisageg+wRwAGsG4KMgAvLMg0
B6Sqs3umfWL/5PjkxYezferXTouqJj1ID2dLiCf/J6OgLHbrWCnVhMpnkOfWgcJ5
OfBmIMHmMHQHVHubhmDuQv327OqXXir1/sFQ+hlXMXQ73xMVdiLOLQ52vNdjqrtz
DZmLotum8P8pvIB3N7ug2uxr9yhGWvGftxyqVcfK/5M8NKR1EpoHb3Fkds6MJDrG
bSGMJvccw1g2EatEp/ZruAOjt1rZF2xZB4hygpVXXES4LGA+c0DBKvOME5KlhXMr
cB45MBFP/duHtWMtfDXiAVa2lxk+f5QLXFgAcN44drw8LHBIBCwbTyerAC94wKMq
R77i3q+qtahXmkD3rtLfo50lG1jj11usk79UVGGyP3/AIwrczfECsYO3DVFuXjMp
FF45mvYHUDOj/6uEGW3Q9JVPwm2dHpJCdtn9f1Rs4IJaS2zpuVSWktf1UTHOMzU7
iszmgvoqL4TEtFm30DAHxKz2GMC3Dmvk06SY4ICxzCyFfy4Huh5OBoh2SBAXbfxF
3BJ3PGUXpBlArfUUxaA0RM9cdqNEHuXvS0SwzoVgSbg+OLZeYpfMcmHRA+TGH6JN
rZ0U2MgKuCaFV+rzA9TeQZiUrTJeNzYjB26Sj3IlHsNYskvI3WBEr71iq8K84369
bCOUbkT/grXaZDoVukjJ1vids6emPfK0KDUpuQFZdn383ihUlxgoGbRqvLtx1rkX
hpZJ+LrzuPwpL1ZB7CpTHBFODMgEh3MQiTj4Zrhql4xpqitzmFZQxOG19X/kOc/2
lJ249w2ZA4lswXqpMJ9X0K5vq1tc/Dbsm7+QDzHbvEvb0UT/yCvW8+4F1x2ZTJXx
C9CaEMgGx1csmLF8NhBa5ecTqoeD22dWoz+f+SUVD4cVEA6cZP3TF3H5gM/H9IA2
gCfc4pFIlgqnRPHspS2HpOjDevvNfcZbqpzkmo2YeMAwupA7WjN6I0/qFWB7yhgb
cJ/eUUZSvKFy29szwLqXfxe2fRDfUIWfLgbwpDsAwHyVWvY8reVw/CpjvsmQDgd1
64wULOJSjOaZwA71OeBxH6qI8Wi71EdYcu1bTRyxQ9PWQBM9GHsKbwhFpGjgdrgR
XDwXhABM0l0BzKn2Rgv+1jEFNO6VzLMD1aXhHzmGHf/LCSSWn9y5iSDtipDb6hdt
nfFhoqfQXyCgcf/Bq7Fzko0MH1ToYyyTnZaqtCQar/qk3gm98rtRAP96X0FEcPIS
FkDkhzy4hVL/d9VYKwMT841H3jLmgsv60fAOC6O3o8EfXu9b2K78DE3FI0SgYwo5
U1IDNXzNRrcEiTTtwnJEw/0XyAgDyJAmfr+jBlohdUoIOePum1BYG1NRpSZKZbVQ
z5dlfek6eqqhdlgCj43kS8W9adFCmUKjZ4X5O9Hckx06Pm5lgOQPINGNNcjfTlXr
lMAEzAn9pLUz49njpB0anF+dP84JstbAgzaA4COa0Zfvjg9bEcnvgJezmAYOTWj+
h2BZTq2OqCiwwCVECqf4juqtOap/O8aUWFQqZK+6AovpPBxbxiIW9JMfmlHH2G4D
Ny00n3OYxdnCBnNp9+nIt/fUabk+n9oaTvSR44rg5Yk8rOH6bjKAYdKEN0rkxVzw
xel1IMybbni0N9L/n4GwwlgmxvhELqc1OtgbHLGp4ArapGBNvtlad71gba2c4C6r
JwFnCdTZa4TuAVW/1W8pyNFLdADgqoDVghNvKukVOQgYZXPRe3H/rUwiZANge/uY
ZZsKySylgP+G8Ulp9fMWARxMludET0RKWMpGOnNJ0J03bVxxB341Kmnymo2XpSzl
4DscL3ecMfrA4s/yY1UQDfAPsvtpjBuTRyBkE4p2dtKFLuIkrTrC+c06apQPCEKu
+HTCZ6NDL2I1/G1ldifn6uIGniqLW/JkI3JhPj84DiNg8qBOm4381XhSPPV7nwRe
/c8l63pLLuMCrMkSfGQsbEQfMshbV6BEQwzkEUx+ndXT+1pRUz4haqF5ibR0t+wU
CqO6gQzJGQ9U8OQ0Z8iWLZYfp84bNNO4nZ9wxLL6vQKwk421fB9ikquHUFpqjOzs
BwqbkA1cJpJCHqSbdgxzr9rpQRN6tLLxVKZQlvkJ0lpkJQybBFZQJZYP7LcIY4HJ
+a+tkJ8oOCVKkX/lC4LVXe6KTRCOoDl4Rx0H5cGTE6bO9wbfQQvs11XKuS/fvWwR
2EVJXMTFxqDHUwlhdO8JFjfHrBENNOpkD0SsNlu/p0ay8qZ1OQYDktWMRG03MUAA
F0ZezkfHDI+XrAtHUJeFNQjAn8ci4CISZyxdvzvULqYCXIn8Y4Y0QRYy+OkpDu9C
6PhL+SqGmTbTnmfrzBfRZ3cR3OnLK2Jwi7v01yp/RQp9lfBQIC9H8D1+eU2p+K2t
QHCvUrVKY2hBJlEGdfeXu8OmLBs8QvJnAnf5J32boONGYlf68DZUHhiDYdnTX8hV
ttKuWBKGF0eaYkaGTcGT0wnNJUic7rjMUhGEtIqHWlvXpZeGQBto6sPnCKYQQazY
e0ZLqODLIu//Dj8I8zvcPOpuCn/LDTCPSfnE4F9C4hrf5pEAybFSbuuZhBDzQJTe
ujt3gkBfzimUw4Y9pzhdP93sUYZo+TBICzJ0o1pBmHZkyC+Ajo2PI7MfzbZFnqNw
ldYX8LmMcBALXXX89GnKgxkDVI+UTqE3Xpd2NdFiAM9XvUdsfafkB+Xq9Mc8Slmj
AVnO2tv68SiEOf0wt2vmBiJu1Ny1kaqwMMRucsDK0S4hHyl23QZARXOWqmf1QlnB
aYjj5roD1bS9aSizWxngM8COBiZ2o42OTBfQFCf0vtoHcuroraxpoOQuM75bGPsm
Emj8BzuRzvzIyY4cyW1zXVaDMjf43oL+aadfe67dHCGueE5eOeejSqB6cSTVbnCS
awnGFuHx/piBiQrLmKpHOiSvA7GDSUBXO+MYSWjXEwIGFsfwKRjX7FAIUtQ1DLrE
JqysVyNuRLBS81EZGXJCHjLXscreKAq5Xgad74Slh6sgJgvBu+wheAbU3upgRuot
NylTsclln9Fpk6ZZTFvrO2D80hjcH6IYr66PkMgVPhTgxBaRG3STuHWZkTlqeiLz
OPSfFdI3gWy9mD4Weol1BJ8Tvk7KTQHTZkvGUvIF8HVh9t/i0zHPcr0ovQFdy4YR
pyrqfn3DKM7XXph1L6iflnsRoq/FidAeG4GBOqVNELs/3f8HddNzZzhD7aXKxSGq
8+GHS6aI7gfYVaC7yllQujjLjKP+zw0jXGNF/JnDaLcSAF0E3Pjdl1s1jRugYizz
GuudIlN0pX+Zovi9qOTvRMnvW2k1s/oWcHw4Kvj7rCmbvuEYKIRim7oM3vGp/b59
VMChlNW5T1DevlFTsyjAkzZFsPfL5Zmu3txAlI+jTDNbhc4zpv4SRv0Xhem1EYs5
5YE3mr61naZg1IuDd7M0+Lfwjy9dgNlTkJpxlooma+oZ0ZHbufcwte82cUQA6217
vSza3D3Y9u1K+ytbsF5fswltn3sbbW8PaaOLSycW5xM3WpMLw5FBWWORMPWJy90+
Eaov5dEnEhmDFj1TwYQ4sw4csLRnywfpULu+vjiujz7w1Z+58Q5sapTBcw6nlqZW
uDf+5MwUsJ/Y0D0Vab6IhRQ2yEt47crPMpJ9uE3KtL37D01BCfFvyCr5B/P1pxWr
O/R6uuCxmjnolRmEitP5/8cn3aw+0VZU3jm0cNm5mGTzRn34bW7+OsYTeidsKlCZ
fMvCrN0d5KNmOdzKeZj3XykuVuxp5NvflggQJ/tqclIttf4mOrTvnxvZ+X8uxaDU
TdjfPnU5Uys4lZS/X+c/CuGJjRJmMgEDdF99XrrPg1+L2X7I/dia25zmdIYDCjls
2DlTb920tFtBaK/egPz0QC+lR5fNK+lUEhYZbZ0yvcX+TaU19sjbF+3s5b8K7P5L
nsavsDgR3BEUNXn6jeOilf4rlAcaUQpiN70sI4ePnUYKHNse4O9uUhLoGfmVt5ui
Vu6GUDrv2qayjt8At4wvJDCIesgj/IZ41LX3LTsszGYTwZN7Y9t0vMasgBz40etZ
E5uhmnNKLojomv0jgqnwyulYw7JHXeeRFK53ocLeiz1RCUZsGIUyf5pwtSRMdUW6
0tqDbz3ifp/ai0xXbrTV5IyvsKHpDYD04Bf0zcs7N8c1+N69cUfif+JhPivQQENv
GPCVAKvGrkZiN22bc1ycpQBZFAHj2Kcep9XC5WVN3eR0srvozPsk6YLv2Agl44XU
1+8EKY2ICsKGG18A5lZ91DVIvgistleyetuEcCvaTiyd/bgWlo42oyji9qL68M2M
TqwwAD2zg/A4yqyx4/rNmXsCbIOYqtyCDxhEVpE/64lsNmo+ZNfpgy/Y1USMXobi
BqWW6+evdYhceIXQAwjeOzcCrL2+sngD87XHcWYZ0McubswrZIXo6IPdLmy2uCV5
ldvDrT3zselSkmG9q8K+GSlq9mYy46PblXBHNGv6b3MNrBZhh0m7Th3am84/zpeS
N8OqBvNu+T3KHZtxxPEFpjuRpmWbMSM8twpKQkkekDUxagqAO1goPi6d3yRtR17H
B6Ta7wF6LDa65KyjGDtPAR9H17dm0mcUEt+cWv5OxAEur8w9H+ZkycLRJlZKaC99
IuUrZZ6jnYFgXQKgSxyBfiTeWV2qI7hZXXQSJwmw1J/WBgp20Jt1OLgrBmwK2es4
T2ztBHCInIFdtQKMieEY2rjs0lYF59CGRiS7g6aPFhI/GaUYpEZtzK60TrevN26v
AjWdRZV3msvBDEDYl2YBDLnozacXOTubbE53BK3mKuGVXHox2EMyNDP2cqwbWhyp
opQmSGD2S+yOihb/HuE//OIPhEClxr8/hTKaiw9LE9GSMvwkugfT6NNpPuW58wuy
0IxZ4OZsMsFLy572V0wWPSlHKj1hu3/LkToxf/PJ+MKmj9R6MyWFdDRSiSs4Z4r3
hgVAIB8Cub81g8wxoK3dwi48ixSydQAnnKfHVsskVgZk2YFcY1H0fnsqw0yvp8vI
Tjb5DeruSOLp/EoFVYaanMyTJf1TGWsQtRS3YANydOnky6/gLI1DaAMYrk1KSZS2
m6bGO7mOu6oIy0MyEY+G0PnLU7QHCBqpX3mWjNJZHYlUun2rtQnEDhTxDeHyGt1a
PgdhwHtsMP2gl9C2orHoz+TD09tksqeKPsa16ZrjYnmwPKdP060/oABKOFcZI0L2
94ChIPxPVm6ApZ2WxyvHRidzETFk2X5uxC9xuhvDy4DKn4tICZkSPCjCBm1kb+u0
rG2OqW3iY3UyplQBDYcVzC9pD4kfztLzGcQHSYpKUO9JYnprYyNNj23wdP6jPPq/
Nzyf/JxDkE7pG5Li1HMhAe/xTFctvEbGqsique0qFLrh2TXnw6eUvCqWXHOn1KuL
Q+OiFLzr1DUucTP7kA0PZaOmIbouAET0a9wCkhOgrai0aKCkJqhSgFuar0/O2sPT
NEQJSfMkwGQ/nSa1TBvth53xIMR8oxXI3RrpmX3ccMIlKUWP/o//XBhhwWj4qIRE
QvGvLrq9NsG+x+WYa0M5gv6l6gRgzylDNBsP8kxOdcj2Tb4Nn0i7MagKiu1e6+1I
zlIoNPSXrDQGcDOo7wh3BFva9/3aV/SMc6DwZZQB19jwb6sBiKplCUl+S/jiabBZ
S/8mgfCPwMutB7Ogxdn0SbZL/IPY/5csFf+M3Qf1VvMs9FGz6JA269vEPZC80I5s
roY+lf2qBb/MdzXaAQbh19bwCz0ygmH5tWmaK76hNCLQmTs3MlA6vN4xgFSk5RVC
Wy7UFcyM6PWSBop1KUF8C85MT+l8C1rd7oINq9tp3kYqAeIWQ8GiwJMHLjIDlfFE
JCLIbeThheA3zbGg8AKrHWFynz/0SI8r+UmSGcK4MozVt6vIyJ2eGxNAzr0HSbph
sznsOFJr0yY2n2c5oLZ8xP2lj1QGnTxhxtx+RyuOllWIiV4a7VATca/ampniTO0o
nWbr7TszadtxkkSL7sfXpAd3RhHXMNhG6MMigclfKDVD6p8V3+eEsvsdMgwohh1Y
Min/eSZfqi382VN6an98KJyKCR9lKctfHaDN+ptn2nbMbxniurM3+UshYbkDPcmY
4g44McsXlv3rZyDXZo3RZ6nHIY6doi/EBfmJMThwZhM4J0ny21Nu/80Eou3MwiEr
Hve1825LgoGRhCwSHCX/wqaocWzIRBTDqb9HSI/yGbBqsktZ6GTuFpXvMf8S0xxU
Zi9MjxhDAkr8KcDvUSavPcsSFQRJVBOTHH/P3QwtiZXbwXZf4AC+V1/29GJhnPkI
At1eDTcrCdk1xkPfDnIJFdJXLCTG0+uh9rEsCEj8jtKV17UtyFBWLUBwucfR7bGR
DAwEGltnzz2c+75JDna0E2rHtGrZ+TgK2f6VaPcgZtFTwgbV7albi4ZUS7jcJMN3
7J0wRS76sur7hO+yCSDca+W05IOkVt/hxzPPFxdodsfhd7VnEgeesBpUA4sZSQVL
5j/i5HNycyizr8HQRBP9PLC4RITg0/o1VEd2Um93A407kiGA7Vbn+G3ZJhHiY+RT
H1I9ALK556YzS68ujurSmTGJrGsFf87LOGM5bt7IiDsuN1hUk5eZvj1dauXr7ki5
oyHkRagaQyPGUxzQxOQfH3xIMqtpbS4nFy5uUltf148Cm/5Uzv2Z3A1aCKl5ADbF
OCcvyEhp89CgSWM2gXQQGwUtwyX9ZABcmuPVNQ+QjdxZFQVEJafpI8yi3WO3k65f
jVPEmd8yYKuDLgPpZf+1h7g+9aTuzBybEg0Hj8TzkdOMC6oI2duBWuHuDcmY+6nJ
re5KOgtA/V1g060iXFlWQCu8ig4MoofYWbTXleJksplAu58GCIPBQCILhOH0c7Yc
3ETeYs/rCDXzRMiqNaknf2mWOwKhe4gQkLRkts/QmkzHo3erWAIrk5maspWA+Nt8
2hKLuuTEpBZePDTrEgjmV/IE8+yy+i/bpZNFm4zkAU2cTD55ZEovH6hWJ4iqEurn
F3TRM5a03M//VL//gU3szzT1sMPOpvBE/y6G6+56iRA9RmWv0xk6ikAABe9S6Fx3
q9lZ1Zf6tbNoWVI5DTEA611moITkcmuX0yGniDiHmC9jsnIAK5/PVWD8YmW9ffRf
LmWSgupGMzCFFFvADbrSiuZIkzNLnSvKRMEWCC/fvsjQM5z2vkx3jElCACKjI0Qv
g8uv9kJKDCf29R0VWKkHH3bGtURV59PMWjJw5JovHxcIUoUXwGcJVeLnt5L1K12g
0ygnMJm+i5kUzS0/kR0G3apbtMKAJ7h1qcV/k5qW8+1/yD6srXUeRBM/B4MHYofK
SoG26KStgIyBQDEORI0NHlaGQMoB/lfRaXhnVYPyq2IPZ9BBhe/S9XVWsO4TXo3q
k+DpfTIVX1mxEJMl9vT7znrxyj184ggeHSkq6nhc5FYZlWz/dI0pyW9XdHAeGAuZ
jS7WTAMCh6AHtS7m1/wh8996BulondcmSv+ZNnzAITY/Ao+ueuCV6FM+Hs8n691S
NBVX22rQx/43NylITvmvYlcTXmA56i9CNPinduv3MKBxWl/o1nD76VDEKhIfG+CW
55g1svzHdLeMVC/nbhqFVizXqTGfBaZ9I7X4bmCZqN7IozPvdup55hwmxWr+Cqzl
NNgjCLbllD0qPLwz2ZQypwIe8nJmMWJUldbQAusWhi0ykTomnW/cTjHdsU169fCD
bxp2R7h/pSppqg0xjrXe/GCbXEwfkyx/wOWDfaNbtZyI8kFnMBJnSuESulwD7C2/
q/fpRZ+Wy+59pKty3PwHxZnXrIqjZz+oNa9Svrs6Ap91SbEfLvhVe5P1BiR7Sb0y
xHAErWwAKEiGq1zi7UYPL48yw6ja7L07VwY4I73iv+nX5sMVDk4mYt7PBnVinWL2
4Gw3o2sZG/QK+xEZBYpDrKxqrOzf9+StC32SXhouW+yWoUoUS++9PW8zguCeTmZ/
V9tXS39XtDLGbiPvPAYgAdsrhPupqf86ZRHQELV/xuXJ2IkvsiHxlXuMEj03tGqL
Vdz+UfctAE4mK+bGBWcmrPlpxCApPrkIiUThXvl+1psN2UYBj8n88MJtlSpR6p76
5ttCdnePLnOM2DgwHcGBcHAFkcOM3p3S5aYTFpeW1MCIA3S3LQY75TPHOxhImdJ7
RWOK1HTnC6XKyU7zOVIYbROt0Jnb+3TY/yWFbh8zVBxy9VIf9idfBqNcxFI6Vx4s
/NP0jLQmV01/AiEoZwMLqcLmZnlNV9MmaFPmMA0Q0ppWBohvGlKBoBEj9Yio3s2g
o4nG9/TRXljM7aM+N+tMkGivlO02BhB65qacKSairTDYOwBWodePK6zu+ZdD+VER
KXJUfe5XTsujz8NqUfSI4FtgmdniyStgLyuSn344wX0O7+vY4vqhXFKHQvoo6z87
JLU5wXbR/HC04Zy2CLKkCbGZJm1mU8QLPC2jaOay5U6MFIfMwBIePyZsWBHurf0o
ag4Ydj1q/zyxxQVUNmqATWBHSwHzwZj2dKJRrLeJXl2tdfJUkDVIepyz0VSqkPQz
k9v1nqGGm8EsT17lfvjDtO2v3zFCABeLdl0O2ioSYLbQsPJUYWDzCHu+7M7g1rUm
RKgI7GDaLoav74meod0cGy1cwPhA/1KpXoQWEkCFJsBZAYbKJ3orJHra17lx1CGL
9iSdfrqu+uq5YIvncX9+xcH4Ex9t8b70+LUGQ6b1O1injFgezwCoQ9vi1sqYaryW
f5McRtjPkjE5Gt7OFB71gP58jUbizpQYfLFHzvCLyFn5awmlexvtFYPwVTN7Xaq6
KhIE2/Z4SkQyzdVR4Ks+FCF/ecammva496Kw/2/TvgpL/VpADs+9+pqmUODIu2aD
Mycl5SuTFzhH/jDP9UE6Xw53/d4LMbVHTv1mksimNDlsQ6ElIRfpv9slnSqPEBug
m9nCX2yyzTr2qri1ODxuZcBH1YV/2swNH+V4vPppCwoaE/2o82MZV2P6Rf6Setam
f8fux1fGPtLs6vejq+xFUU6O3ssJuYIleLpw5ZWiiXHUPJn+aYqCeTZb0a3eduR2
VBtc9NpDHRUvmLgQOkrqN6wyMDiMk7isfo+R1OMMGeWMBlGkojUz7W6H+OFdKzz0
ivhgNciOgknyTOFcXbucuc5j1ZF+5e83Ut/uoup0/70wpEM19LXbSy8ARHS6MHM4
WNwxMsMX+76rNdZp7y/+HIxqp0GgPoGCn6Z7W1MKKVg/jpYXSyhp+8vBWE8VwGhj
mjlfA9TzRciiElU/P36mhbKRL91Yq673j3ysHEpAHLXMmGtSrWI7/GIwKjZ1dnIU
MS0CKyOAsNFeNcJLjbyDlW416eMrI4ZQJsYQGcOuU6jpyrysq9/xtfe7TDjykQWV
K61tlUUpHmxPqscmRuMG2wCBJYRx/9TJ6Jx+OB7FwiajBHtbU5VDVNRVSqO6VLGs
1XxIFb9TLgHxSB7BA+eZTpkkVLukiH97+IhWDIkiB2m9AEDPc72sSOHdD/HpQyRg
ZzDYHucZ2iITL3C27WmxjmAEiocbOQFrlzjLsM7kOjrDb33ELNr9Alm8Hq0wdMBr
UcJkIQxxqfZ/lf7Tl3pdVfATP7mIX/3foguvFquNeUBguWaC1VHhuFeagAhUXCpj
L7focZQEeq1QFu8ZqLl2l6ZMANCK5lXVnoJk1JAjBmMBQTY4QFlnW1zVbrLKM9/W
lrMJU0IfsKe7p8k42EWlKul8qziCdusxL1AQ2JqLd4a6GVI1kVSKRZ0OGaC8K/rW
Jf9yyQFSky4JEMqZM5pk4kupravSricJo+EqPx2hpejvxA43s29A6XHr0K+g/xRV
j0G9+a6ktN/Lio0m5MNXxGxI8E3g0gtrr+Veiru3zDKiSmUiuqzcL7iVBnxiMyUi
okG0bq2+lyySPXJz3JvfARWK2EVMWdQqSDeif4K3w+dsbNMWnF/TdM6HhpfS0zqZ
YGPyZvYhmXBVBrRKqynSr2C0Ug4IkUrmn4y5377Ver5pX+TIRY29ia/2UjIADRJW
rJV96Tu1zm/OYFLAwwAL8Y/DBIkiWlMm4pPVwe13badkVYUZvOzp1t1zz16GZaia
uylASeEsJqhLFJIZJD2S/EwIGsdcMPombn7lcU5YnaoZVdpp9naDNPbWszZMfIVF
nbNyJbDJhN2wJK2RUfrRCwVkimu/0vCPDl51AUDnX1pn0bNWionGbXe2fu6J8myb
OBq7mqGoz2Gf6ROm+lENvG5TBDMEmRR31a21P1eTpIrI/q7g6trOuEX53u9Q4MNd
jxzjxx2m2hI33L3aTk1nzmB/prUrFGB47+FHtYybrqcUsC47bNxZzVxblkXNrVI6
NvVBbJuDSMsLXchR95X3ICfAEaQ/m2ssWMI1JPk0fCL2qEphz/fOQl05JCPyynmC
+rIclFTSCXhlcmfizzBOODRsdUxaTGskdyDAFtVlHu6Doyn836XuBXWyG8gh0kUp
Yv+uFv68Hx3YarQhwVTG8bBllD0dfmTSt9JfJXaD/1UqI4GPa5c8cWPm+M4EeQ5y
eLS1w9wmbn5irDQVtqf04r3l/QNruVCB7TllimbG/aeyXW4sUqKqiR+cS+NBtKDw
TscZjcZpm4ambPT0zxxBUHNmQpJBgavWpEZ/QmeWn9Q7hZudwGOk/2qCiCLCciGf
MLJa0pgZrSWZtTc87xlWoUkr+0i6FLM3FOfEzXM3re7wafAKeDYN2rEY816Ffi8h
1KKGqkOlWYdvPQ5ETSjmUjX4b0Js6e1/mCLAX/PsnQXh/6taBS2YAppjn3RAXCZa
uaAWzMW9h3sbGgeaq3bW+huClkT3VMBQHPIurYIiSqArOQJeatYfll/IEwEtq1tL
V2u0v0TBbzrkUPSoKOluGZ8FcDmxGHaF7NKh/V8VoLvbZTwM+z4EudBrj2R+HC62
SE4L8R1zt/lWQ+zF9lv2S6WO2q64VQdYq0o3dZoUHF/RINBPhTllnfq1v/eHED3p
ToSy/sQsWbjJH+/nA1mWWaou3fsvq0ok7YJ2QtXrUYljo7gcT4vvVBm4v3ZOKyKP
VEIIjq8UP/YES7cGpLY1DY9mCOnYdLxKF1slBsWl5lrReEuXxjt5dcDBt4Z/dL1k
sdzaY/VaySo+/DiIOBJ0Rvq939hRkyimZ9/YsjqzFKNVDwstBFsUp7hkUNyry5AB
CVUhdNaHT3q75uPps2lww2kWIcvAMwMNxa5YlI6UJL/BQ7zLlX3+ESZp0/L5ce3K
ymmWte0jCiHtjnpmYMGq7rwPBVpzN3PPia88a01OE4cDK7L940FdOREgagqD07qb
gz7F95zEDaLONqQ/EAVQ5uYiPjOrv42nUSX3WQw5X4bDkH9z5PJ7AscR8e84NvbY
aKUCL+t9f9evhgB/RBwiP7vendqJdbhWxyZDKm0Y5ktxrGTJmJPqpGQNLyEhRWLR
ubzusnsp0jrRxp1HkPum+w0C+YTwwJoW6ubN+12CYRL4bw/4sg31n+1+RCRQrBBA
fBwPHpz86g9pHo5zK0c6Y5Kl2tVKqCEsaUQysEoE8OEenhQ23buRtu7Gg0zJpqgU
0Ckshu1j49TcB4CmZz2fCfgfgaTwEySLgq+pGwBvFbCQz8/ia6BBh0J/0XXh1kDG
SzUOF1nr2SnGFT8A7TINMMzvySY4KDKdPu9QI3riZb2rXFOI4Lsks61eGiacamWK
T/IJWO8qhHSGznVJ3FDgTbbNC80TLgvI1iik2wBa3bCzob8Eg3viF5JEYgt0lHme
9OV5SWx/eJyWiYngBhrveMevOYxNghy0464tpGllJcEfIwM466SHUm7WLrt39HYO
b+I5KntxDXQZWX4MDu6zkFKPp1MzxwbJ7zM1iFGD8zeYydzLtxlhLH22rDhsk59i
83cVKyvc7gtarpwFsbDhf+0R7nUCIubb96N8d6UjAAbpfHgPaOtlpkp8cLlSJXkN
5LbFt3338f3y5nklf984i7fh70dNAjutpAaKBkIRXzwF1wfhwqoH1LsF0RRQsERk
zPENRWdBtRAOXEZqTzCklmUQwzFiDrxmeUWcd0LxfNQLF9KGoS5Lr8rNHotlim5i
Uo3UWrigTjJDrT9GLIH/HnlVFnQ9Na0ZHwp0eKIXw+qs19CGszUx0u/NkmfAq7jm
bGXoh32q6cx14ljxyKRU2OGH40R1f8FdbfQHzPZIbEZtNj43HsdvZkt6VCECETPM
tdWm4Ax0Ealol9j4s7vuTeiUiUgUDsKsMDgmJh4pJdrQWQaD5zqlrtw8nsEPt+51
PzF/9Z0A0FIBPJ0gQ/HUIT+6mR00GY//bsHYHxqJLz65UxhN7/FdHhd7RxmEPnT3
G1GxxwJwT674cTOrKdwxxeHURmZATCbwJWxi2duyE4AGIGhvyyObWwPucjyussYW
2+UAr5RNW7bIseOShw+bH+IiMhpqrUwy2HHpDyhS1LeHGN/+zc1TDlkrUQ9eOgly
lM8EDQ+ayIbvH5qR/rnQ7WTZl8N4k/hJQH5v7ZwcwTbvzySG8lrzVS30Od+EkCBF
qV6rn2eiKcCJHNKAqW6rwRTAgoDjzN9+74/UyiX/Enxv2kIrJy8AUwQVc1crAC/6
YM8Zf7Pdg8/BOQOB7cTLsZrh+WXiR683jwGmm9FxDdSru+FegujRsQ1iPJEJzeNr
bhoGy8KdusDtByM2f5YZFIcO/QDOehJRVbhc4p5vB9Rg4yIBDrABCfy84uWkTVE5
i+LnwAucUFEQW2UN2q5B0cg0NmaDxFQ0OmlJUoGCPOW+HW0fVWuZV4umppvQ9u7W
9o1A64yGmhPhqoyoCN1YLQPfSJlhoC16Y1l2GVjNxt52wAEerUJ71c8/8HFMRkmw
nIFadaNnqJn2YdtCzvFbX+HqKaJsVKm1hhx3ZNHDA9dCfQTWRC5GJFOwaL9Zq/5q
WTWjU7pYTpBq/gcJyvENYWn7HO0NP8dV16CynKveOo9Rke124sqtvxZwG19RXH61
pwomX9pkvu7MMIeAot5p4SkojF3z0Rv4kaluFnG6la23PVF9H38MSmou/4Ht+Zgx
NaMKWjRFxF91rawfN1pW0ndXHJZjnwn97yP9gkRlqYKFkcAL4tZfA6YBq3VAZdOh
E0aV8b38TtxUIYRYVyv9KTOruY0mP+HzG5pvLzf68Xn6AF6eLe9o/FYRdXiUpXXj
vOcOUmGaaDowyneX4dF6cKvVanWzrAoe9Rms7RX05GTbMi5PLkzCnX5P0wjWRng/
QiXlUmDXhic+4EayWMrVGiGNYu6OjEjfhMyhMpgkxSRvVIde6R3jJq8WGie7PUQg
c3XS82lBo+S9ToEv2of+FbT6hIzcKbehmVM4tnzveTYgNIm4dD1AvOZ0B80En8PY
ZHDA+U8wPVtgzc1exsJV9X9QHV39i+MJoE5NSY4KIp+0jjugzdfsfdAn7e+0X16W
wiA/4AjRusHkYIzuCq82hYmt6r+7z4Ra+Xvze5eJS0b8SpdFC8nn+42NBTNFGura
zmgoDqS31b1C8UDi+tU4wwY8Q8e9mGDAV9rzasvEEt8Fy0f6i0amMaKEwTSLXdRV
KKisYiJay1rpSlGLx8U5m8RK4UNCLpUKL8rDYF+dW6I7DzbjHuW8eUZ6mPRg3+sF
fE3Nr5Xb2Jl1n2VA4jewb+d52Ct9yiHr+qg39xeM2oL4Cn5q2dHAArf7yXurDD/h
xp+ZtSF15xEJb6jXupBv9oZusnURT24GeuFBdDwMcS3Kw225kurBp9YTF/yOPUyy
8M/sHu6VysK38ZypcG/LabCsjf4pzrtyVqQvfzNKGuQkdR6PsKqZSg8qde0Rf1lG
t7TTKeXFxpQMSt9sBmTf5PP19VaD6G3u3m++MdYDgN6tvaVteEFYHrENR6RR3TKR
gP487iWaJY7VeXXOGIlCZvA9iTiHCvL212+WgH9A9JfNqYSCoPY0HEqJJ9ZqxJ4S
7rPC+yucho3e6hoi0fgnafWvbIm4qLgKtM3TeY3N8d5Xx3CWFbkPRPDoKnp3v6M7
GYM1QuLMShwp3jggiKqXPmunzyhb4cH4M3Y1/Nvw/9B7q+IA+mQiE1ZDPTCNINdl
2CcwG1C2+nvHqZrjBqoKkoMVkgLOBwSdS7EtJFj34SY7kXaVB58IUahA34E74d7F
NLVOiz1KI2umoKHGqkgDKPlqwtnen3RB2qojpoIIaFx4S3VeZVkwyP9WkoppvH1S
PS31dDbYruNIJzoPkrRgNwtBedI27Gqi4f+pKRqbWjhruvPZUkEFPGuBv4LR7kpp
5CoxPSKG+5+rJcWVogrt71f4RH1V3Nck6BRJCQ02G6DDKHqDpFqDjA2tsRbqnkYe
BikY2A79RuEfT/GgEZAnl5sXkhcstWtIbbMOUAcjff+iLYpyu49bUKltaV61tMe+
v9ZnLBxnLxsnFEsgdKq9kDFVc/7RdEuR3z73K3Pf8XvUuqUVwVHBEQzC/0s4wgXz
C2rJzG/72ijht9dEKxQxRiCyPpuYJUDnpwY+87JMM/LKctv114SjabfYrQN7vTva
HxukqrrLB6h/qBgFFv/3ahMTkHr3xexB4u60PviRKUplZGK3ZCzcga1ec3iYKOFC
jYCLCpXvF4YwEkoymH+LJtBL14TmVDqcBgMe6ta4bTbrUjnXBQnU+jsk2KnGbvJw
I62amVttHaXmq8w1RDT+4oOd9XFqj/YQETAjv06u7HN2wXDTIIIKtK6id45Kwbpy
141HnKi2pZ8PIhdEgp8XBvy5dchVZyETp2Z7laRDSH8N5J17LG+/suty7iWVarUC
g0bK2M41jZlrTPyhk8r6VcCg0cIz+FIQ0haciM+WExx7EL+DTnqOtQ0T2hRZ17Dg
7/Hdk/wZt1yvOdttVsDNgelRPnOsmhOlVmHadNj0ZdftlaOxtW+0R+NFaCJNxJOw
NbnQ3i2es6xBsJRmpZG12wEjFY95LaoOUXwIh5sBARAglsCmF0jsBZHQ5XgFdgwc
ktdtvt0u45ffDiSUdrwaCU+UwXm6WuF6P/S3T+/vu4Adco8xtmIcPH0loOv9CGC1
ub7Ss3sNlRRY/f0OZiF1oa9cgVTOYzt2COr35I+Ok5tFp82fPgGyfTsYj8oMy0dt
KbDvpvYubOewhi+kK1KzruavaN93TfdEIMWDT14SVhZOIc81dqv61g92DMS7VGM+
tqOlqyoHVY1/kEb6lphoNepHuxScCKwEoVKWeSKtFg1MPxlegNb057fxr0r9om8t
KgDIaZpMSMLuodJhpXgHk9jSe4XDDfihxhPN1gTzC6XJTc4adTTb7AGtdEOLl3kU
/5ZjGUmsb1EBe8Plh5nxjVoC3CqJ8vJK9l8Ai6EcHSoj9JzH3QA3AMSsIEVgbZTq
WvZBrOCa52AV1IDg+daA9FwOFI74nFje6FaRxPBVgLRmCU3TD1ahZHGDcMRH67Ke
hMn2O+DKL8yQW7/WnRIOzq8dPkeNajFKjIQOTEPGUJAnAeF4KMJFRNBT5uqTxp66
M5WxLXe8TXD67WpvqT9qRA7ncUF+ay+GgiJgJ7cKThp1wfqoE83a/KXMOC1pt+nz
aK524IUDr4Qh5SSI8D7IWfQdjncsAZp130h8X7kPAkKfHY3vJC0XGnHiC7+7SS8i
e+FBVesp0SxSSM9q6nzUfZlf9ICMG0dNSk9h0w5LgGlW0LeDt8JPMA7eROAnrK/G
kKt8/ZdWPkF2cqqL2GTpDn4hOXb9fy4z6bPEfiXzEgeoXtvYl6LfljQwIU8An1YJ
Gytqw04oseB//rKxouKjcxHEdvVrM0TtbR3MPiU8h8MvMy1347NbZKeWCZhxb4B1
1TVadliD8QRcZmbGzpc6XdYf1vOsiowTg0U3CfaQozaBZZXq2nLPr1whJA0yOnQs
dIb/V4F5E2qkuj74/wahnqvLDWAsH4QplucTKN9U3cHwZXzXYtCIcgb8Muv0PpIr
22YrjUCJ7VIjkK113ZpZSCGhOJBfjF4pk7AkNtDrer8bCEy2JHz6ZQd+XzmO7SbJ
QIO4N5VxI8MFFOo1L/UthgqHjMO/WlGcED2u0MSulMQOSiys+l2D6YnB7AftcqSl
tEMeBmSQDG4ni0FJECJ4T6ifpDShFQ96MjqdsApgytZRL5u3xSkfmMsLxTMC19b0
D6ubzLqa0eDtjOMKo32t5f5behDV8/kmJAL+58cXOCSJqqQbNpV/if0IhHk04lT+
lZ3/CsmsWpQ48o3NYiEuLJPx0gvR23yiJWmNLe3VJUQ9SMhk1ONK9TiFOBUTDh6R
WWLkMGsuLlsVySt48/9jpD8hVenr+3i/O5YLWrIsMmt/8Sop0OkObM+08CyEVHrO
1uF4m1UyWFQWN9j0ojlwxJKdVhSKTmjmtUuu+arNyWyLEg5oPdQBM1GKdNx6RWUZ
ZMAnYgMnDM6a7XeSPCsiWTFtpORr3E2uElwBXG8vR3jCHFaZG1TrDgYEZQWsX4fg
j4y7gO1Mq9MXwOuByopEzDPDiXMcEW+zyEma8gM7vQwJQkA+EFFyFxYDBlItQjpI
RFoAJ8OpsiDaBhUEefcOI/OymINmXdLF0CM6CCqy4YC4oEyqKpHcdHk8TmoY/Zcw
kMw9Zf9Lrnqtp7RyCk5wvFD+p+ENpdyKCo5qPEU0+QFQpNwDn6JLSh3CXp92wc85
giXnrIKbsEbvDlD3A7OOunEaOtBskGCkjC1cVlr7/KBHgvmDunVk/On0TBV7xqS4
+kHJf5CWTxvPIp2Nj4IWWYQOAQ1Epy7C5XkRNpoxLx6Q2yn3Ufy44gtAIDecBhVr
7ZX+v+vkz9iAX5pUV73qBRnSRwAJh0o0o8T5GiqpUm1QxV2xOr3lrzWBLT41MFdE
F4YHTvmzl+cxGMHTnv6mMMxB3LSyITn0V/5yF3WnhZe07GrSLhISIsfnLW9gr0l4
QV+CToJBim2DMKW2Xf0A2tmHy1DCNFuGRnwNXzxZ5Uvp0gJaTlipDmNS0T5t37YG
9L5iecQalV8Nsn0iaMW5xHRxkwVCJQDYzJ2GCJJ5FiANBtewQLv2V82npZ6+qF6V
ZxVCe8fV/bml+evxVk7UvqxXA+fnEWdrYbAafIr2o2OOC+pvTjYC5AkKMU0/H5+z
RN23xLzklB/SYzdYRFcuenlrIvi7wEAPhK/sgt1Y4iKacUOr8/Y65uCpHkY9Bzvc
7JIwJuGHXXIfPqMEYGtyvq61GAStP68tsR6x3rKgqT/7kaD8299lwISuoQWlE3Ef
yGN+qV9uc9thbVsn/hEdxeVMzDMFaNXfmZ3GdKOvChJ/NaYLbAFjd9JyeLRvCHlI
K6+JQia5APCFhqsmSWe15R4XCbGdrNpqjAPR/BaIJxio7I5vHo2h+0cipSqEHbNg
KsTPHYGc3tjNzItEY00tsG95YeT8WEYvs42Qw9GIKv9EEwpWnVU9wzmTY+VE/27y
LItU90JFQZRhPFO+aekXQc8tTisY2D8rEuKuTwgvvESKpvj48lE0WZP6Ki0aDzYE
ADNy9SK6kumso7oCuyb+bZcTEztvNu7n+5XE7KaqX/ro/voen6lzOJlAAJ4Ny9G/
2GUvYC6JlROkG8Ews0EeaUr8zYw9pkQrj/kGcUWT/AuBnSQbnIXX9TPALqXK2tuD
mtjdC2KsTFhMjB2xlCYz8vMDBTOc3+bNZmKpk+guWBcI98KnVkT+QK96B1KzbEZR
NQV/pB151zB+DKhsOaaAv+PXWLS/GR2iIC7CnaFohzuGkZFvAQ7p/nziOBtGoU0U
ove9cFroPlp1ZFxmjFtIjGTcQnzZS3CJxfA3p6GeoKkEimK9alBJ+sOaPcDGHhfW
u3nA/MdjBJDzoPHiUi5alB6McBwffQdISkiR8bS5eslOCTfO76oinY8GLQ28WhyN
pcRgVJaZMWVo7h4m7izxhziUtZqHYo/ntjtBeXXsCLzKTO49XcqS91zz5ShqkQZD
896BCTIhKF/ZepUVEf4hbCS5SnDdH3lLPmdxbkIQg6uBB0T2Mmo8UHxtJUSOmHme
qxSPalfDY6zPg4ZFaXLWuG5WzYLQzgBdEhsQh9vGC0xZ8iEw5V/b5Akg+WhBJ6Cr
vVnWU7LpME8qAcbQZRA4kgr2JRO7NNJTf7jOro2GIeDkmY8tBrhziR4guNQ/QF11
vqzr8kRF2edM73Wy4gIpkKEipMCLllm0qArZEVCkZGWjaZj2tI/AVlubk8FN0bbh
kPu4Qq69hHBFevjhXLc1J/OzWEbEzpZSulf6hhchcZ7HYJsCW7CegT3culaJv9Zw
QaJ6s6c/ZnJzPtnSy2cCYTtMymLLuMJDN2GMuYL6MwNDm0OZxseoAnZwWfaDhMzX
f/29Dubmy5LuJuBDn3QxoSmRAHq8R6HCbPI4rBfVNU8Gl++GD+2VCEMjia0DYgE9
d4YXbD9zN2V9QN3mWPjG2STA8QKULOJasu7c8ML/YJ6NJ2lzTdb9JCZJA5JRTxc6
GlW48Kr0twoPzWhsb9csuui+EYetmwac1Tx6Jy7jlMK7s2BjgPUQc5tlTJ5CDElR
cmzIipofTdWY3HWJRv+/TAdI6IqRv6p+lY0OvuOaM72bQKbczh/Iz42zp5sXtbv2
ejYD0Q2rbaqQWQhdrloEWvti5tsIGJSSn9dAKZmceJxurQgnR5h9ubt17DPJ8S+N
1vmd+wcnpZKORa4Ff2UMLHl1bbl/CA3WsuVGb5NAKXN67rGWWD0bOVMICVhhVLkW
W0s45Q/qhWpRsXeYwWWJkWL5NcieK28Pt2nXRe8Ek/3kHOeoBJnkk5VgZuWU0AF5
71eZOZLvIQMw/yg7u+ZSWqq6t0zhZnxOdx1+2pxev/Cru908leCnrn554hCWiRUG
XpK11hmWHw7T2i1d/6FpK4uAz2HbPCJrUDqzeYOhl5tCp2sh0UK4NWCjw49ljSpA
AI5iYiOAI8MhQSI+s21wKa8HsfNkIZLRmuSck6aSizUYujEdfDxnPblJMCed7ln6
LcZGg1YTpR3yiuIEQtZGAC9psKMpGGF00BJDBtZclvWj1MgZRkxSiF7AHFe5Zk6a
DwKRxdy17XtfLsNdqcDEWVBpz/NLbTyl/sadSuyBNRvaRLMG3sGitNSOky9BM1bN
9pvycka1eaaTigcvKVvc6vkj1i7DXaqj8Ez8X847lzM12jemAV4eP3ZokKYrX9M0
yoXQ1lUI8g19JeP6N2my8veHgIoWvB8wrCIXNpgNFMeSGO9m6KY5EmQLSmw6rwKE
/0qajksjSZSAGnLPPPU7hi/Ec+XTSpBzC0CirqcoG//x0F/WSj48S+deI1gWMgL2
gRsiLGV6nNgib1x/0l8xkaoL3jLcDekSqGK9tYrrW4FTAK9mMviH7X87bRv9feEh
8Ti5aDXw5MumIrP7L8Z6vF2US2IE1RXHrkNw/3klkpBJKx0PDU+LWXGernixvChn
tORxWlE3/QG/g6FLu5DE1NGxYUaQQCcjwWErloLma24VOJHJ63WS8VdjuFnE43Fb
9Jqw7KzlNMcc8hPcykmf12GtffQsGzeh9c8Xh/1mPbVD7UIzTW9yWoYWcM9aeX2Y
LQ8J3YnEmBYvTz4FEJGL5RgHlyACKlg/wMtXH7tbg2yRLFpnnHwgMccGmGsN+aC/
GlmoMbLWde6p03otVU9+m8Y9lRx8Nd5lpgzvzO62OOI9fG47CwJrP2guNphSqJmH
1L37masUJnHNp/1/5i9CccPxXesm0xFpqPCs5hkObpNkahm5Iht1DeQnDj4Q3Uhw
BhStNtUr8nknrqHU31/bk3XoxdosSDnB8Ah3qpPSyJyqAFEi0MAM8a9f7mHIBR59
0JWT0oq16gHFYLrN45CZmcrLjA/bUye1JkYIfWXIa12KtMuixUel6AvchjBvCF6/
r5Thd07G0mM0kaZsVUgyBd72ObqLkb4U7f6ioIQdP/afvnT4PjKImaYANYURulBR
U1y9qAlGLQt72aAiaECVaMdN5D9kEWPZXXT60ypBLjfyT8b9R6+7dN8rL0+gItZ6
XXVxXCYlGc0NsoMuYiYgiA/+xtiM/HEyGrCfyvthHnE5eri6BcFm75CgammEGP25
YxIAE4Jy/kyuqdZBpMrylVXzwZln9blz7jSSH1U8syYlpnfztPwU4iCwaRHIYPia
h+hp50QsvuaqccCTgZFehKjjJr0Q9LjR5fmL2TY3RoRMnjs8EDI+DMGlrcl8aZov
/UtLjE6veNXxsjjyov51+V41desrIK6SXiydfGBELWpAJtZPc0P8xBvS3MX766W5
KSAEd3fUOOWF0jVpXzJrzjjtkyTX41Uh8iET4SF99+W3nzj4zq05TKdjBA+vTfAz
LQueLhWggnJ/HyLo302xELKkPDv+XLAdeZXK5PRdHtlcIw7HrVkc8Ss15gGWx0oX
UycptkKYtkd/yOACbqk/YlrBHBYjUwlSUyXZ6SHveSvBAznKMAVabt0N+dvArz/E
sXqdECYTKJ2zkCb9M0nHSSU6EryGXBrUr76vLuXuW5/VI/h2NvmcLdG6yb3rxjlH
7lVwiOms954RsPygexoIfJDJPONHjMvd+XSWTe7wY4mC/1eVwR48DrYfHUjY0fWe
mZtykS8O7d581EuFLs8rhPMKV679+XJEkGeklDlbSfJOhL+r25dv+9+A0xLKil3B
WVji7lg/eYRdvKh2Os80AxbkkLfEShnOFS5wIic/Lz+uUkSx6DUijt6wdfs7Cklh
96I67sMjdVoBYf7NRP915P/13XFFhAIHeGc4puHfVMejwM6jfOC8CWHce0F0TJWz
TuR7z4LGegTIXtDRn5yCyv5m/2K3Slq5X4L+XdN4PjHrzme98L/UErUIG6jWza+t
G1Nf7K5U3omhfcAz+HmJ7/y9OOHwUA2AR3+AvEJO9PPb42/d+wX13DewFNqB7DhK
VCQdJ3Z3DndtWwCuKY73Cx763jLDJwj6Ru+u/w1PZQ9fzUXztvB5sm32wJ7DlutF
Mxma/i4kkacC0jrwcq7Q+yW2HjAxQn8F06QMNZj8jcOHkuseZExCZALk+dq8YLUh
R7/HFnX+cd86RXwBclR1J+3X17CsESg/vgaWzV8DoJJ8rx2w6bJ73AZlhiQTEhC/
Ve7NB18M3TKM+IL0RIvYyHgflkudEbhxXHWt3EQO5P9yGcgvk2mofpg6U9FiDH4l
f4c4o4UDM0wKPB0H/5BXpoTBzBL4vGbjzZim1eTyKQzHDmQvVDqbwhgsViolYXVz
XC3ZaaP6+3KgVX39cUzZ6DCPaitYU+Ktm6bf1AtVqC4zcYi8AMELhkS7xHlFLgXd
TtwZMFQ+wwzEmfVck5/VC6OtzQeQpwFt6qq4hs1jHDZ2IWCVasvj7NAe/9Asiy+X
4TN2gG9ifCgstlXBTJCUZv/7VTszMDYLeXoEMjK6km9DO31EcbToh/y17w4GFa0E
wxcq2ECdNkrOzBoOYdhCqHfV+pzcgROL5N9j8hyh+bm8lm8d5iKqDFF6X3VzNtj/
TSMgcXNU48bnr0x+GZXDYJpE3wAxo7vqrcLxRL057C9lXW0VqzTVjSehgVYLYopp
a/B+XteSXmXgG3xVA8rQ264BM+MmTFMY8n7yDvHvTNKAXpsUTCv/5dbmtqnyBpJC
v4Q23kvXlr1QeNd4Zu9lfUtHHYTaDu0rHBrnqhpqzNat5o0zP7I13qAs/ME5oSlF
cVYbD0GbGSspQacGqeafFsJQU92txMxkRsTA6ee7SHYxappUO0xQid7w+e2QQeny
MKdyPnGzxcMMDwbYWuEMi2OSr1CdQ/CN8rlvNzyaJgHlA8JoW279HEVIeW8Wu0RP
ipaflO0bDIZz0RIkX6c26EPTmVODIIs4SDt6AmU6DaGZaulLlKbY1fIp48xK7nYr
tn/vnpKjqR3DwdUsq4It7ZmkqaAAhejCjNRlh37BzhTEuI8+1VyHKdus2ch57h4B
jw7DIb6fu5Su4v2IjNXoi3PYl84ivQs2zoqsbCHP/WQT6RsHdS2YJsQX3RJHw5qs
tW08ZVNufY+FjGWZsKrnOnW2CyKqv7VqaUWVck5zZawQ707kmBRrjCOtahS8x85Q
AEd/7ohqzGosQfmNt13ZzysxNmMP6c1w1aJnPjVWB0Kw87RuYo1qKJT7D3O2alxo
vXsaQrnpN1WofAcH1BQFaaixwgB3Edva3PACQB3qoN32VGMCh9C3WLqXewNLeR1T
ffy5nOkfvqllva6XLkRnLBrbn2kUms0XViAQ8dSVtkxc/BXcu15hGAtYY/p5PH8c
IsMgFGxe4CeuVQZGbLx4eZQwVdUZjiuPNAVaeiCE3ifJiZ7hgvpxjc8+pcIYTo9B
xryn40U1MfaVRyJGZUd12hYHihsKZOsY1SAjcUnxZPYzAH+CryKg8Nf3GOrBCAjv
Pm63fQccLMkzn01YnmVdibXMoGP1DqND2/VQJLFFpxB3KpVu+Ivz8FKXrTtw7isN
fPeL3xxYU/oBY363DKhmgeuW2aP6FAW+f1YCuR8R17Cr87NOdmaT3gHPR+BFgJmC
9l3SQ232zCP3XkhXyEy1/Bvr1KaY26veK4z6Vtu3EbLMgrnr70lFRBT2Uh4AodQu
MlrMWt/DEkOiorss1R5tJVXiXZEVPwuSjkIKqyaVn00I0YE/Xp7WsgYBpafXvOUX
vw4hWxLMgEYZXoMPEKa+syYKxTdwychTAKCiFYqJbqP7uqnsnyb1LEXSwR3Y3kkv
gQuKooFnW8K0jTblGnRWQWA0pdVm0CQfxkb5kWl/VFGqs0TxBLph3b+Muu825NyJ
zkcDKt/91T2x+ydOD1OwL0HVZJijnytCMdU5Gh5Qok+T27TwsEE/kYl9BMJE7ddG
SEIh36x9yDfBBHf4XAAnY1c2Erehs2mKvuzTLJKb/vHNC0ri1I9XL0Pu9LwcAzsT
fka+3dAkwa/jJpOu2TnkNpD+OqP7LisI18zd54JRUWTRKCBlZG/FWBZg/RlbZt0w
QhYOYP5dXCCPtpkwAeucagjabNnXoLKuxFHiiHgTQoSZuHRQs195k2iyp3IrV0+b
u1qfyVM4DexC0R0HVJULy5fmjy+lAfRkTii8kQ2NmLi+SqQzW8nB5ZhhNygM2qIp
ChkLCcHW/Wk4NeB6iVP0Bfwar3fMnwVFNvgOtJ5M9F4q/iAjx4sqX69/bkZXLDAp
a1kLA20fot9IllMahhI8/TYHMZOfFE+oZOcVc7BOBTHezlK8kTc0H0yvy7wHrtlq
YJRwriAiWG8wGF3zDRIHgKfwrLYWCOA2lhjB39WUpgdymY/5dn5eT1eQoTQv2lWI
JfSfGAoIoz/r6pA6fEtZwPMoOD7lKKuVimugsbnLU/m5JyCo9tzFXYjMbO/pbPl/
S8+rZpf9dMreEJodpOtQDyuHmuHViYV0QOoTaCMiPl43fRZSsr41noaiS/co9bbV
rtwSQ1ieUmJWz8Cz2PKS5ct2DTVjsfMMKE7kfEbK1oox3NLcVZPbovdKqOgAFsjW
DQnG6fev7l22lfbGqn7fkJviVtaDJ0pUA8iZTbgivUdwhPG8ioIJY4u5GiOXRB6S
XTvBsbDmglmw5gZI3bd0LQ/COoQdBCXQbzT9HStSOg7DXZlFx00NB4TNrVYiKhmT
qquzqsg1ybEwFH9Cs45bdMf2MHwSVEzVBC6YYcMjUCSUGfgLjZi5OKRM0zW9GYFK
R2agb+s8rL6XxhXasGKPlAkBLzAel5zymXs7bfvR8+VeN1XXEkWBn4kd1wuinG9n
BQyeL2Y/EvNw8yli/w1wFJfgFsLP80uLOEDRcOkW75FnahM9FD3RgDydHbMgF9Om
+xCgM0dGGvfeoAJlXr0cMd3Y77hwVQniGKnBZ3jhvYFuAfRLIyiIVuCPrxnO13Gt
eOVLqzwZwX0H4GtTvEHP4Ry+Zz6ILPHNTKyYJ9Yur0Vx6fHhsAnY9K830l2jljis
1KKexGWRBLzHFQ2hLII+8SLx7lZKKT0KaD5L429AGGYYvdI/YcXOs0vXHKK/AnKG
weR2l9lP8RKbU17IGvi+XPjXki8Xt9etviVgYI32W2KUgammncghyQGvcVbuM6Ez
gv59VbrUkZ3SWIs0P/pTaJkhhPUCmA+dfzfOBzJ8/UsHlJb2hHN5X3kckQyFQ3R5
ZCY1rZI+bBKZuowrfx6NHyNyvObMBxt2rel8+sIfiyJjhn3kIzhTzuAKyJR+edqe
4KPKIFxP+ORTjR0up6Gvc9cBk+h9kR1WnaoKFQJ0D0UOHyHbSJUSeaLitek2KfYr
FY0+xIn6QaGEaBIkIzBXGNAXCuHAwlKAfJ4JaTaTsCLtecrBwtxIIIaGTr/oFahV
6f6er78juoVQp6cB3X79hVPhNEKaXfZ2jWxc0IRDqAXtf7c1zTF3drha89ZUlG3t
ZUfx+KGCulyIjwv+JgZ5giCnY3nDJh9FamnCPlbGKsq5xqbxhYGyrhAvAbtGCzDs
pvX3M2FdLEyKe8T6KnDndrhwqI5XiVyQFM2MYw3uBwrva7WNgq87fujPeAOcysKQ
Y3Ju7Vysoge8o/IT2RiwdM23R7k+y7Ib0gGXCksy8rXQ3in97PiA0pxbIRl2a80q
78XB+oJ84F4vQKMVbV1fPXPTLdD5gzekwdNGOcUa3GAkO6vsEu6OqKAQ1pKkc9IA
Wul2xLdTQ6lb45QT7rDFkbcVJWHhHBPopMTN6vd/xCOuYrbmvW2XCbIwVoUomDOw
exU6P0uGXTeyYO1TAx3SzUWAfD8HbhA6LXnR2Lny9Bp0o9gmNsFEZD36x0OYD9Ns
Xf927Fss/pzLM3Lo1Kt6Vl3oQ/jo3v/IqMkD1L+0NRTBOECy+5C5OLQxwm2nDPp/
9rjKoNh6PRkC6tVD1WdBg6v+08GEAuCXOHpG4g1mGQrqdRI6T/ptzNESp2Vf8t9K
j0li/bs2aDog3BTLVNNp3egVNPoZ71Gcrd3Wbdfs3QUogrLKWbBqn15d+l4ARWJQ
VcckiIPGYCeEuEHVJScF3ZlRV7ZBNVIHkBGRvSQtPPbc2pro55coVGPtcrsIpU3n
bwDBZUxK5vXWXA1X+qt00X6VCTfttfpHIHSBnGhZ9APDCi3n6/VYwPAcrI1Hos/8
h8OU7gro3c57YtGAQWlHwUpYFVQvVj+0Q4pVwZexYp2L8WZT5tlR1cz6vWXIlAdK
BHm6+xznpFNt4taPKNZfz08XxTLDJO+pxxBDmAm+8RN8L5s9xPsp9fcpuIXrEN33
TnzZIjZbIAQvMIJTHfcQoeWFAy3lIckYjUHNfJmzce9ZGFkT8PQ5slepczfsH8+/
neCgKem/mPYLFUQfZYEPCdK6R0lbt/YO5Lr7Wn/YtFtU2XgZKXfUhSk6dp/12tIh
tOe+Hc6y0MRtnlldOllcbcB+0AMqeScMDZ9+dulKYfU1raqyOx544Knw7bWK/EXU
JQ4ymsNzymmPWfhP524k548YzKwX3L2G/w3J1x4BpTFzHbM4pgHo8eBBpLd82viM
9u2e+z7mjc4CENAcCyt66Ec+SMZWJj1+WbAIY+enlRkgjJ/2A4skJwaaXT86LQod
KAyiXpVnfxEcs9kA6edolbbN6OHMZa1ZCcm04OH53cK3d+ekGyv5qXMOQp7arepT
T96cX443yWZ5jtvaKXMHtPpFq29WnYZpuTyrHPneZ6VCp4QK3SSIcF5u4vJtHGrX
d+QKQqPA5Ax9hnRXzwEjarAnnwq7rpxbFY70B8i50s2TrV3f8kfzxOQqqGGsOduC
IgnixkBMmzFSfXEriSZ6pw340SHw7urisNISjoR6rQDM8LGs+CFOB4JxQWdFcX3G
GgooG9EIHxr9EiX3XcLfHvo8C/32kl/lusWK9st/gCSEEdg0L9/GARRJgvCS5IOY
r7n+eA1hzoT63hCIqUkToXpMBHSSocag+Kb3VfdLclSjIg1HUPZcbfED1mNmwZSz
BezWzS+8zesYq4InLP5yP7FYzKB4fE33QgrRxbgu606LNlJOSgdbp3BnVxC/iDZX
exRJkkcVSVfoIf/0B7rlmv190/aLuWeyFrOKcezr8/lfZdBZE0ply+Rntnpr7Ji8
wOJ1+npAnWTppS8n1vZ6uTHEkhVGlrA5G0Uxj4ia7El4sI8QzBzbMtL2UTuOjsoR
f4H0nyGAaVCHw1AkEsQGzWgKJzL3HFCN2jKr9fWgVKeAZJvoyYA9IBFkvXgkUxLO
ZEz4uIOUjXiR8YQuKrVWr87mGIOatB5ydyzOMjsr0zPc08aW/OIXs3Xm5zY5NNwL
ebM+FxQZkAbI81StaYV6p92s/t9zqhHRP9mwrrARzU8uWe18AL/Ar1Xe4z07Ux/R
LI0u/MN7OvJKllSsw0bMraCjzxjtCTQ2D5nYjJRZ9Or+ZwVzdgXFU8GUPSoQgj8E
pYz8P3SU9du7k1izNdPhRCCK9G31SBFVDDiBBlJ9tSBRD3VzgBKQwHxAcHf/oWrS
9xQ/dZDolX6x+q1SKNOeA99H2cvDKcLjEPwV9bp+XHseqiAZ0gz4rzigbsD7gFVS
CHHOIGdyPQJ4SPkNZhOYCkLdpN10fN9shRowbKPMJuRqWXI6VJZWT8ZXwFEobykX
aythH6+32p5o4FyUAt6WX3xr+yBm45KsYoSVY98hTrFIJB49ydfbotDygGIkzXS7
oMAjPYxSH1RTZmPi6ePOnrZ+mPSe27hJnKPekeHojqDMOJN53E9oNOFk6bEGVAz1
v/ZjO8QJ/sulBmSC3ei5ixF1ZIxzsPUrFSOSeJ2cpM65bW4xYbFgW/JsQWxbkNuo
9Alvv9cMXlZFuwSheVwd44Urur5a6w3benc4nlfsLDhTFsrpQurRtbDkrogzSGLF
xjtCDTUtWQVSUkyec72x91IGYg7japJaPN3fYmu/IzBLQYKR63M/UWd6DLJhSNUJ
KHUz/hM5XixuJdOi63MOLn8HFnISFoaRysp1YuTFdlnF3vc7THdddON5duyqIsJB
hDXO68UOeLZ4jdVM727VUOpgl4sZbGO17l12e+hmVG/XY+tdFsagl18WGKydFxkR
7jOtlULyo5+q5lO+LxAJbY/SqoKHoROlxfg99GWk1f9Ao1KQLR1tYicQFz3uIqDW
EydT5IqMOgI7ENhtd4nIzlsV6LBeEc81nNxO6PIhg2atSC606OFYMCkukr0sipKB
L3GSkC8KFedPLqmETfZHkAKCmjxBXtYDQxoGk/DYUg4njVbo98tXbbQ9vGRCqWst
JCY1vBCjRos6rAeRGJBn2wHYY9w2S2urbRxCVHnFXQNgAwxB97w2YpZverZbomms
/WG4GPAELbpUfYX5q33ThmNCte5qATOuAZJuEI3c7Rv9+Om4aI8eElzyv9U1vUB2
sOfA4aj4UGuNOZypVuL3k3ajfGqph93BJNbRxhcDNTr7sLjwEME61Hi7CIMn7MMz
rgbmt7swi4JC7VfMOZP+a/cUrC0S8oDYdx9rawsoi8e0EHWKxzgjOR0Pl7eF5ecy
wiIEOWCXUv0cCFbE6YQ0HUD11UsnAcKr7Q7P1ZrHrtR46/A/blhfhvl/fKtydKG4
xeNXr4lCK96fZqwxVKMWoeKparK+vCF4jsgzBmEuc42BOEcCcpDtjT8KuCBiHLqp
h9SDEQ+tSDNI8wsJPV+nwR/y9EGj494l9lm9AyC4CH6F9XDmvMpftn7/tmivNp4U
Cd/jmmISu0DNzxcQ/gelz2CAcr3fdtdjrS8PkY9NXzUjp5hbf/jfTgei+Z3FJG8y
EeM9dButdBqsxLzq3cGGSRlknLBb0RNf50BOAWxcvfW/3LWFkZlC1EMo5A2MbctK
vaAaFEiH2LLc/FsYDbhsEu427p9KfDPe+gfNXaJTjtS3ncM5xfY4jM78igT1JZhS
uKic8gr7WHMMuARIrQ5Gg6+HvaRaJWh0It2UlonWkVBOjlVgNfEilW8ey/v3mHLZ
w3dD7R3MU5pZNTTi6bklHZHn4yJeo0nJmlj0ZH1EUyveczhbzGQTtVXechn9pKsq
Dh9N+LRCxzV6Fe+s/3gDKuk6YgKOd6u+XS18cEWR1A40c0SmH84PxA3vjTh7j896
mCuN5Cc/eZ1WdzImVxZidnXasWDnlDE+87KqoQD7CjmkJKHMMPxMw6tDYNnHG7/Q
tTDXQxBPs9wn4R+AuX4r1tFN3m/Kc1ugyiBAffSAcQQUF/OSPPTE3e+AWqd8L+KC
xbiSFVhRib/lloyBoE3x8MGtSojPHk7v3AF69h8rk2NkFIb1NlSu4h5yFc968oq5
Abx3eUSpj1dG0fgrxDIlhBAR1nRD/dhLpeXp4DbkjzxjjIyEaJnQY+UIm/ilG2cy
utcOKhoIGBQh1gvPP9l9H0Bdxn61yCsOwE4ApLE/CaQeFtbO3tbBK1pfDHo63OZs
6AlDalUxdS0RKIozJomTLlK7+CIihu1KtQcMCvQIzXFTsBW0hayLa5QoO9q7bsR3
XK7jgddwkmztnMyGOTE58PlXuQIKCCGDK+v5U5nwEa5ssuefUCeUyc349MG/OIoY
/s9F+lSlcjWp5zqCaDQJaMQ/KSdB/OAeCaq92HCXg9IGYeKSFYREvsryZdQRYWxO
xk90P29rGJaglm6kGigDDnORcN6ibc7TRxv5F3ztg3SPbZ7lq7BYiBf5ZowNwNLx
HU9e2243/2dL/6Ls3ErxFh4Ik1ZffPvVuPmqRqWp+SiaNdHOJ3u0mhDBPyZ7hYRv
IfXjhYJ3n4ktv1ZxGDWlORgiEerGDawyoCmnUYdmiZp15xY8VnCJfTsuRJZaDZEx
57ESX041CciqcvL6GKe4bbohxtUGjDhDBaoA2JL4XgD3/bwfQw63lt7GXVFuzHAy
YyuehiSw+2klgCuUIBbmqGi15W+bwui0ZFCHCyfmjdbP26uGwmuPbKPGO28yxNWW
8PHGSHZIFkuxGNXv1ie6sQNNVMHBd8VgeLKF+ebFbqT2m1sFNgWJRQsdDyC5uqlH
CdLoPcNnVv6Lc+iugsFWTwvBcWCNZLpnGUlZdD9xI+fVOuKllr1YaseP1bg93oC8
C4eiqIB2KTf2U6hv2eIkolRj2Q6LdMre1UQURfKoIroUryS0/hFw9R1aSi70o0BV
uyh1DDp51Z8BoSB0NpQeONTwIfuhlaTlvF4orqeR06kCNiblyodJCPSspRl5y8ff
y9cYQ5H+reKZrCxVZciMWc8HJyav49akBw2MTb0EpdQcSxBylQtDvhf2OYP9O/ab
0jo67eXV+4asa4EdmGL7Isopu3Ck1voCfaGoUBQqr3sm/JwKGud3JJXvX8uARVcX
bkBHrsjTOo1lWx8YkDPLFqBf+ysH70LvRWNSuD12nE7iH0W5Y5MVulVcl1G3n+7c
3Ing6SwW0WrV5VaXN78j2HKfJ27w86GhcD2q0NsvHnRyp+7X3bgcHpphDLJeqy9l
6jFQPRDj7En3KMxh/kG8c2zJ/3X53GGDnKP0egnqSxWinVs9yTZN658G7i4NmSzr
3SAVmqVEoWjLJBKabJpsnXlRklqWPsPM3zPgqww3aJqPstfBh4zR96Cmf9OzU+11
dGb/JFi93NcDpWJ5RAor8T/KpP5acUUtRGJAe+zH6Uaw0Fj4GBzwdvzNo9HI/4tt
pDVbDyFOKsytOOO4ngDKR17yFS8LeFY3DF2mQhirD+9jUKFUnse9fwXIxsSkcW6n
TIxHGSiMNJlT+T0gGcifhFHrE+OrKU1W5KRbIq4A8bDRHpBKJODuuyVCGa1JLIeu
xIoh3Ng96YB2/XDQMQPWfT54Bs77iuXp9xl7+9ioQDlXjPz+bczjhaC++iYf2UKW
b3tMQsL/WFhl5/Lhpn9d/F/N8N31GdzTxQ9Og/ALjNt4TcoJUf2YCFNTuqm0RNPz
QP+EFa1KZfiyvdPQj2/X15t5U9MWxAHIp4Gmo/Ekf5TFinRLqXI1ShNEnG5YuAnF
dH8hh70Mtz7Q2+ZpQC4wPfFZ9FmaIPJPca+wbsEHocLjx1MAGOwMvBv7VyntUip1
7DBq8zo5WMWduvsEZdM9ndv1T/am5q1DeS/x+wge03+6kQuHkbYe6cALzQfYCWm4
bWSUkHoKLjbAVm/UzBCISjE30GEk0vOCBi5uETvOwhRZpL800bgvouvMv8lkLTh2
xaSLqp2otA4Sn7CG55OF0lvUKk9TlIPIPAKNwSCyLX3aEgTCnmKLX3u3cTQH5xP2
PWJxCkug0GgweT1Fe66P302baJBEa4x5D/AT4B5lrEGa4BRkG/WbkbyAxlStOBQl
Upm1fogvD7qNh7Ld2CEAlfKjZshF+WX++xEWnLYh2w6fJWmW9daTBOsvWEDMjn22
JnYpgHthnRS99viYuiybrJqLdsQE7SdKLjiVzCJjMAGIlOsuqgYs1MgotlZWoRq2
DGJC4y2kcUCJDQ4LNKpF2hF572n6AUCepYyj2tRpo4SJv5X8cXD+rdH2abtEMXEj
pFCol2UdhFoRGBqzgLWz5s87CvyRf7HsvgtwIQ0cqiW3wwnlgYXyOGssJbYxxeCl
RuTm5G3TJaNkAzQHSotpSRuk8gUcHncKEjKQiNpY3PkB65kEnGeRKCvySZJry76i
tnbVB0kYTsXRgo7XA+41nDc0a59tRyuoe+2Qzp9xzN1tRYk1pOnwt5PXr1j5vQa7
AvkdGmr44aqpFUrWDyGosYHfvVY5Fzn5hhIdSLPMMKSVidd7GyfNWQhkaDCj6cwJ
Yxz18FxHn4Ekksp62y1iI7L7F42yYQ3dXLDER+rMFKDZt7SjNQJRptMF0/PJBYG/
SQ6F+hqTTn9PJHUCzWWDo4h3Tg9PBBjl++tx6fHPafeCHy5llNlQenoS6uYTHxSa
+U364HE3jvKkjEiGgpOtaWb8SITzoSm0d6K74gpZwNPsPTqWhyrepirZzOL+IQas
i4Ud82KRNgcbNWyeMj5YKCVVbc28z+cfaRc5xHRkh62g5g3NKQo7K4hrNnuFe8Si
jzfZWCsUPRffqcO9a/5I7aMGs7F3FRtICCrvaNvocir+GztEDIh2vVcztb0+TUu6
TNOk7SiVAXr3D48FJff2eoKhAVOpkqU65jlWq1NmmTxZBC7l73iWPhd1/7WGaidg
/+C7jO1f0q4ihcVz1AG5C9J81Fml1ZF8n+9vE6DcI4cDEGgAWWu8/cYQ66cpCa9L
0BhnkPvaueBvLIOQ+cFGS5DCaYZRAbPvFSjO4BAniTYrbulm194YO7eWRRzSr7lf
j1xhCIVs/l2CJ8fyVV4uhUOXJfsiiHdFxaCaOPUpKHOQFmDNlQnoKXDHCHHD7HGj
jjU4TP6fhlPaIGEUswPBG1G2qb7V+DM1ss5IBop3wv2K9sZT1z+DbDBPQdANeiwq
2olra30qGjLBJsSsxLGi4/zP0zmWODythTqRgpNLVOjdAucs2dRn2inwI9KOIpFu
ajd2nQdFqVtF0hlTIG+VjJkdkfzhJ+D3IKsFk+JsP9hQHqVMShAH2wfBAJdxL6fP
aAt443g3nhf28Aw0wmw1HbgUEKgsm1IsW+NFJENcqo/+D05W/TZFpYw3Gl+nJbjd
KXoyBMdtvka9b976Dc8K+EYyX28U9KjkRalohDupPg3K3fEidr+WEV9aNq8qiy2+
QcW0RIsfDP4rKczqCCVhtU84XvSxwMaU1IjOzeoY0vDFYaqCsJXFt3kpnqSs5wMv
uMxm8WvXqPzazu4TMKqhhejHAEUctJ6h+Qe2jxNAPQ90hF5IjrqCDhTYlE828WWT
hV7KJhA3FYGFiM3aOpyG8ErqNvLfEqeqtj4RiqWz3apOlzBcS+si7lE/du/N8bvT
85rAuHQZnHIFiVvdqwPMl+fyYYnawblrGcFfvIZDSQdkV/Ft9nFonX1I1uAKzKg1
PFlt6z4S1KrTopWAYWRiXOGwoc8Q7lENw5l4wfTxF5yRDJkcZkTbLxce9Y8TytVO
gcR3FDY295NIl7wqL9D+FPKZzE+rWJnpCqYjJP6kfxYkzP0vl9ewlkn6gmalKzcP
4xfxYaGWiaPsdzsZHg8xSaNW89Qthb3pHdjKSTf5DCu9SPwUavIvNS9IkQbVtzNu
8Wd+/AplUi40vsK+ttXBfe4dlQ6JFK5PX0wcZG0M+9yjud+5evvCOhemoJ2meKAi
ytqALjcUsUqtTD8otSYowebzIcIOh557Llt6QFMnClnIGp6z7boux0mT4VBIGBwg
l/VOa+cHvKEss5VeMWDnDjdasgAxszdzo/cGTlRDw6aVr6lgtBZyDVCIKOw/ayeH
Dk448oT4jVmEoiEk81t1HvbvTosA1gKePkDCwdVPUudefJF52PQT+dTWZw0I/x7A
6SqZMragL7qRai4zqQv5nkhMBrsDOOOo/WD8iW8LZjhayCcGnYuehvnUjs/GCLy2
hrz/Vr/8xWwULhBJgWAWdaYsQ+v3J6PqUiokX3ep1jUGT+itxjPU1vXwq0hF0OS+
50nkRJ903YL8koHP0/RQMLFZAeqy2420ukCgnkh6kFdcFwVO1oRA3lZGbA7z9Vc7
O7nJkxzqFprPWT/P5Mbu7U9B/LCf++Ugp613WoQvEu73mD3l0WqN8jxgg3ORHfGZ
EzbBjtz1hBYcBFlNtCP+CXEml1JKbp53iCaQS+Agv06vB5TWTVKonS8MCqaLYT1B
0e6fkquzAbLvGghh8KsL2Qn5eD0uz/wL+3xKwMpH6vrh0C6qkPfRZcsJUYWT/Jb2
TXu7hrewzto4+yjDySAQaIRfAO1GDOpraeWqyXxmdAvDZLOsDSJag4K9UgCpt812
PJyLONYcZMOrjEmGfiegEfZ11tpw1n3XifJqyIFw3VuLrurk38BzO2zFh8BVhhGh
oWhxRu2fj3ucrVhMVctRxEqNjw/gR+itTwc9xwJhJvD9gv5bTKamqR92+0B8BKB7
7Rhhoa2l+4mg3lYWcLHJNm40Z25iBhiHJaBZ5xDJRRXPzF/EDvSd4jAEmeySjPik
siSQPhqAm4THGyZTst/UDUfOcCPF5/ivstJ3zXeKTINYZWTNzrAOucJwUbO8GprE
YUsyFBHkLHu//MRZI74EALadqfaaDu+m73mgJtAkIp5OUv6fqhk/YOiGHWAAVPJb
bJnZT6lFOYaPTad5CVTTDqB8DQ3Kyf/Rf/G1iH2onPOAWHmphkR6SFPNjnCGJ1Ej
7oD07uk4oeWNAERRTBL5QKhF5TOeebc/Ftw4LP30N/QPfKqfqlU/9V+njzkm+vK/
rlTUaiuny+xP8FHM1FY2QbdQ+VP0kqYwejOAhAkVbyvhUmK1ozloxRSzPJ/CL768
/kCg65/AreJm+gKz7VKQoWDh+3LHOb1HsjZRElTgU7IuQpH/rkYGURpWQ0d8OdpP
2JPIdx/2GKEfNeJoDfZaKfgMHhprgAPqwG8zYum1rqyDkAl6rdS3PRp2NfcPDOTj
9tEXzP5a3E/ODRkbizEfvybHF+FjFvCZRGZeBs0u3S2hcVNb//IZvGP0hykVyu8r
OJ7IocX2jg3AF48mIQNCB4NIx5O/rXofKQIisRp1feXuG2aD8+CI8jL8XLjHesML
jEdA6UwPIabL87RH01QUvfWGjWr7tBTD59fX8SD2YoCxHIVECfuDRZ5/1eV8RuHl
iMGlZXa/onvQ2zl4DXTTAt0TrdDHY3QpQtjvUWRCFYoVSmO9/QJeuw0x6eteYUWh
hB8XTuKLdJZoK0z6bTaXHyFurQAvKpV+D+3fQXJfHJvAqPPJ8i3lUrzH7QCk/udt
Vjwt9WAfUpylsIuDx7/6n8vOp+ThTBPiOXd7hMuoTtm/u1AECXSVwiMbEOU4L3AZ
Wnx6K+/fAS92XCR/bHy9kH4ItAbn62v5oojaVKmDSYBaoPDR4EySwjxqFM9PvQd9
hQ9NBTGKdYxMlwCXvM8Uv2PjqzdKSErIm6YGOMcqx6KPlANlrIAuFknWbZgojV0G
oD6excHgpXZkMTyV1hBNmG4wFP3HWKN+9gGPiu1nTpw3ZmopZ0ADNfyy7cc4f6ma
6i4U3VIwBQxAFxAgFNsyE88aC6d8SCO61cudp/nNyTbzjMvWh9gZ6vZC+XNUpdMt
4lud9eAPFcvbjvOahLr6BzPAwjssJVwRltxj1WlImvoCwRODWvJpxWgk+GszUX7i
WCWzCpj4W8P53251OTfcraFC4mV5p96bQWhyr0yPdpiwLGvLEZY9GvJTiuSEVQRb
QuMvzvbs3fUp6g/tpEGzE3QQ1VvtbhMhXGvVh9+F/fo2VmQy+th4rpyfyHa7Rdeg
uTD1CbBr677EK2Rg2q0S/S1Eu0sz5/d49R9hf2bQkSpDQT+MZP+in27YPKlLBSEr
Ndq8rDuqFj0Juq6BZpcz/bcO7JKR54QmqJ2YfzNS12vyl2U5pIc1lfJExIwweaL9
z4HQqJ8/yynV4Me9kb7WbTgZvhdpHEP0kJ0DnPUbfGiO8VopgobiPZ5+AcMW3Tb9
WBirX2jaBf6uujh28QS3C01LzhKpwBCC22gUN0tOL9jsi4qE6doubJ8y7M0LSO8L
/z5r8M1b5MTITFS9I6indCajixLkXuWwnTZLqk80d2loRA6piA/dKYP2dBlQ7fgI
vX8sGapSjErUDSo4z8S1w6EJlrNpaPYym6HZxOH3t6VyjtVHlIm7+EQ6DrOv3qja
/2JgHnuIyLhS6ktA1PJ9H8OmKRbFMN1TexdwA06+vgTrhXPxPai2dLB+dMmk8xcb
FVJcVFjchkZiI2S0EUNtqrf6lKrLOThPHqGPiLpkyOVoSVSm/G6tjTZC4GwkCpql
ECTM+jMBzNsJayzXt2Gd9bYUH2mkHxoCvZzccFuKEbAI4QwLLU92aaTdi9Qi1nLu
SIpzGIRSY83wO1HzEYaMnmGIjO0IIyxP8Aci5rflxmlFAqf4/Butj5x/vNBpfmxj
BtlisBWDR5+Bm/xqzK/NWcsNxy7ZVXRxZ+v4BMKN9SRtBcLxy03WpK/kcjXHd/bE
ZEumPtuI6taSeJQOjwumRWj5Rw/mBvGs8Yvdw9oVoZtRWqz5uuzEw2PPObEWr75a
IDdWz+lXojvBO9vqaF/vcFjZZsQE0aCWO48rypErasWcOVFWh07nxo/Ea7ctswfZ
zuF7BzBatW0LPf1SMzLGok7nW+0u1cw7MfLHmNDOxCm9E6FJn1iu2Y7KH0KkMksY
GfUCd01+3tbbEpQNVZYAllgU3EO9RuKKFxZ9js0GY3hKi1Wf2Uq0RkeSawZ2bVJT
OsWargZZwpnVkB4lmMrFaqufb+czcE1cNhB8MWGKbq1im3lFGemProvBOMP6jziK
5yvUhfb9D+WgTSEQS4wMcKIXioV6GVDDnXOHLvkf6PZXkwBsN4Lcftxx6va4QrEs
sk77k0LqT4TkF+sWeAMGNpqWcs//Q/RcuFilShz49JAWpOyxgZGDeXbBxwZ0ngOj
u8rl26FZ8Ffy+k8cqBvorRdvYWM8br96zbl2OoYMjwVUwP2vzvq7cMFbfenSacP+
JJ1kt8mJ1E5p93VtjGP26IsYxYQeyE3SuZmKCsYI1sAwP60r3ft2Qb24uo/gqK94
oZbPJ7UjMNV7CzuMtAldciCkUdSS5cZ88dqNo4eHpNLH+cSLviXUzyRTVg8PQRik
33PBAyua/lDpMI2Fygeo2qSERGF1ybbH1b9KAG+y5QKUuEXySr2sD+HzL/uss8A1
ftePVo7cQF0WDdGo6QfodDi9LxoCLGWDu9tE5sfNuzpozI2Mgh4QlKNotOzreNA7
Y7dAWTDT+P5pp9qIJ720a4r6SJeO4lCqJk0iV+c4u4NiYJ19AQGSjsstS3JkQIVi
I6FwbfbhP/WjWgUHkX6J0mbP1c5lUgnGk6C0ZY4WXbTxeP5TD7R28q86RfYQSH6m
W3SZH9v40NkQiCuulB1xE5KJSnKlOJutyKiz46RplMcu7cu9HgNr1YrHlag6HYZe
crWMMLFLmaUy/W9HJJYpoO9u+nBDlQVjsmP5lPgQZl/bWQHiJyL/b4X0yz2WwiAU
hUzwgENXLSVHBw7GSHahceWcLhDnPstI1x5FVJ6qEGJqetUoPCIzGVXBRxeAHtpl
R3VPzvQPXkt9ZE3FzKveUCJ7z2gTVftS1V8Vr6qbbTZpqhFW7juMW6PpBaGieFpq
Zvow7qQJXDHKt4UBcyfYTK0JqdoEMkON5ZGFL+flPfYAJ7LevIKmwQuiRpYjf173
A39NFu927Pk0orjegPJ57hNvih5ocFHf8jwx33TrItLW19CsMLq4WswB0ztqTs1y
Vz/HnNPGyEmRWqc4aurqJizmZhsvFWhl9YIhmQla9tv5LG5oGL3eBBCFCG0urkMq
AjlQOuErIJxrNVwMwHadDrTPEvhl3J1p6mKvxs2bKVEAtdAVFPkWJC8I5R3ICGGy
TBMaGTqCYcKvnRxUgoMscjHX5wEvbS/gLElifg6t4Jp5vL1bW8XmJMgpDL26XNjU
bAedo43b6T3BN8zXyLsPoGoLfN1om4c4O4qE+EtjS30r9XmVW4rFOSc0AvZOkIWR
pWRk0k44lih4vMvFrZeIwCjdi5fiMNyIvFSKPKRyRgCysmQlobZZhORx+V5ARUOU
IERnylCV4KCLvJR6OFP5Sn7nXNxRboSo99chmyUmsvUQkj8n7uktkrMquOxnql1l
hSl+vZntuIcCzSVztsJaW6KWghmJOf3f8Cd2XDeu819A49StKbYnKKYd0Sxr2s81
VwcpXlUmild11L0l1ww1htPugIWdiTf3jA5eFfykLZuvgL3MzPlFDlwBkOrfjpqF
iODMDmjDcpjYlZhuJP7m/pk8Stsd7e40hqKYEVijZ2l9VRM/Z8wvJUZ3Uhs8Vy/d
qfdkmalW7I7RahjbB3/NZpBa3RFcWjuK5iSz4mWBnt5zfuvegNP2wW49w1+tKLwF
YKA3jsxIqqirJsTNAFd0bYdl44FSfyH9cSZzkBUAcxJNQqUllYVWYiKvkK+jNEgj
nbKZT7BocCr/4SPPcVRT290e7LtvzZxg9LRRonpQkIAjxXqL9ai+OJ+leRJz0NoQ
EftmeTHUevpOJuWZH5ICqj7pE/w6lEJSAlbRV9vz7blasAAkBsYIa5I6ddDILcMc
hbQ3LTZryHOf0LnzQY0t17fiwoBEnQe9oituefwoWfC4FWNgHB6IV8rFRFef3Kft
aH4GOxa8ow7xBDwXX04YrZKg4eQiS3pxZSxhcx6Jbejw1vGW6sf7bz40kCShcKP/
VMto5wbdbohrtTOeYe3BRsYU6qa/XY8+ciHNJqnnqRPjy9GfyBcoJGUgoi89mbuu
df+mm+OQNoNnItvpLCJdNQjg0XOFiPh4+EhLmc9YVno7HBh6x572GR71sCCAxXHC
DV0vAq/lMjZnm9PVlN1BFXkAiTq3POBr6uFeyKDyBYMvo0PCzKS7HWv2nVzuYHZx
RZDB8RmNQ+KQLPksI4qaJ2R8vrKi/uasT1Ys8v7jz48ZvFFUtv2q4TengmoX7p7b
hJiAyN7ZpJnoOA72BqeHccBfWwARVCsDMcvf7X4zCTYKEc6PkQqXBCGr0VTEymqq
VhKSnKlKBAF0FWj/EPVoHQuUj6ZhlfZVnT/ER5nG0YRHSJE2kiA5IScBNDUYaTYH
+w0zqZqnkXzNl3ZweWZgPo4HiV4+FDdRrZ5gQcdDddbU5KcGKiyKfjJiDND1q3Z8
gZDfmrkoGPfSL1rLV2v3PYYgJq0DkG/3k0FFaKv0VzwAJW1IHttSIGYRvTqlr7YP
9+zUXrlYesy/DNiQvcRY0fXd+gVSYDYsjOXBU9WSY2EpfTr3x/cixmOyaBVjoLr1
SWzugUO3jAMxoeguAyHoRRXkIpU8gRnb2bVBxN3r5WAeYsbUrOLMWnEKS7Od9VdT
eOU02zJajuDyFV2F4Ea+nOhBmbwX3/gcnsP4HqUR5xk4xC0RKdR/dj/sKvqRm1nZ
DbsBRAlymj6NO43TINSxKcODF7bG5kzuqt+RWmPq3QcmA/BVrNqm5YlF4ieFQBSb
OCfsjj+zWehQPDUMRIbmzGl2FTwcfhjRe2gq2fPdfFrP2k3f733c7kKMjyk6jEF6
XTJHq4TszI4bDrnPpNZ/X4g30dPrHZetqcvBLapxp+SXgOKPMq7v3N3J1xkmeC8r
vi3EAmoST1xIqPrqGOL2fZGzruZ5c67FmI3a+mnIIR6fv+hpYZNoA5dFK1IDDSdn
0NsJzAIiUWkUpYM7f4cPN9zagBEhf62BKYoyKgtx0E8puIOc4h9mcRIh/7HzexYL
+jw4kBC3bPlsV23ASBlfFCH5Tli6/Jm0BJsxs832G2fBQHaVacN/yRs5XpOye2KD
2r8CRYbqpEC1T4cWxxE+ORqH5+LC/EQmieWOCfhslo2JK6mh5WS9wyhC481f4X0w
FkHk8TmDW91k96X1n993pZyrNgWXbhy1tM1OpINDr5K2KcXRjpvksz6zLhgzpGUR
M3eeeozQZlS9QpdbHz8QZaUBjRWPOqr3Tbd4N33gnfAEG1f8vV2q7IKRrffOhe91
OCsVcnMx/6WOeY8np2ypRcNY7Z7/TkeAKsM+wKWHL5v7RKyBGjE8vpuZ6bgCJIaw
aI0nLjzMBpM7zY4xDnZZ/pPPbOM5XA/I0BHvvS4Xy4RGTx8rfLpgqZcAnS4HZVCA
3wDlXuWFX2yHeLNZM5T9vmcW9zC2A/YWmmA20CQcyz2lSCT8aZ9U0JBZ0rh9MRzt
fT1V12UBJ7yRrFAHLT/Lg09FPjp41WPwOgCnpwE8iCaAZn+CFTActlfjH5lFrCck
eRUN2nZ5XK3PLjJDCU+V81Iickl9bEF2GA/TyqwEfflFQ9KgOZLn09Nz8+5zds2u
ja02YUkGpnm3yK7S8LUfwvSmcJHg3kPDAisuuLMYY3n1kB5Ty6FAOsKzd3DHwtIC
GQJAYyc66RtxD4qAekltxkyhFO7L6MjNbL9gE0ZozlSqIjnAvPWwVX5cbVdSIjbw
TsNMws7n1vOcuczm8POb1by6MGqRnCxpuAR1to5qMsvpiIDUj0lH8N7zaUCvZju2
Z5qXLZgDsOn547ueB257ImAvtEXjC3b+sWHibBL5wYfMUpg4w+OByJzNk2t2OFnJ
BGMhN8PXK4e6+1E05w/vi52wG7H91cq9nyCRJw9Jxeg+mYiUt9nvOnh46xfPoM6g
hr243Do//R2JB8MS5Gt34DNoWUv8dSGsT7g55AT17BAgILJL4hmqMTsAMk+5IsOb
xkLNT5MhPSGgfSN6QZh5vAQ4R8KucSirJCgsSbvD9UV6Se1Rm74QTOammyYvDXIp
bqyDHUKUx9PaQW6cXetmcH1/Jr5Ef02MBzjfrV5WmXqF+y5NOP0WQFPkaNcMJG1M
C8/uoonOqGxw8YEHqpwnXL+LKf48Ge7yUbjxisQLsk7iqvdyuBPTmI2dEkmp20Us
uZjen87c3AiQapxLVaXo/PGtGM6dih0NidcrtB8ZD6qZiH7Vd5I9lTYNCqmDPQo3
/Xf6S26TmI9RHZBw8EmOFb90DJX20xL5lj7u7ualA7h2YroOXeh50NA5QsPlqYhx
VmF5fwjeNXxS4BTZ7uu3fLN1I2zNBsT3i/9yyfClAL7KiDHtw0FPxoXYdhP7U6lZ
BNr0dbN0154vl3/26JHMBge/uKNAjmhDi71smGWErQt3YS8I92jUNfCJETc59nSy
U0gJ1eYProEUwOgY/ekFYlbWPjx1Ww4Mo8S1wfnNDuBm7KidCUAkdgSIGSln24Uj
GVbLGe4C+AIb35w8EmT+ej0VqP3tCaXyRMxsYogysnoC/V2XgsWoPw7NQGIu2sPI
uGAXbVG2FuCZDjsp6xGcSLmf39AIXsRZRkDxYDrHoFzcrMWZ68lp/NtBLPQOmM3J
2k25Q5MNNRgN4+YRQbuCv90OxcrJwss+EY9jOqky2x5lWWt995dDLHNHteO7QtGL
qhRBgdDUBSgASx0b69SkF+v/9LfVzT5G6IXaXPlZf4Xqep9P6tHkmT9J4B4989MN
4Pj1UFdAIgdZ5C0yb9ISFh0slMf2Nex5cz0YSiLz8YTXV75G6ejegWBAf+DXg4GP
E4uT2OT8QzgYObmAZTTeadSJwHmnQt8YAA925IAsrKy0jZ5Ckzk2BmTH/rrWdyFJ
4n+quLXkCKaczaynVltHGqlukCrE0NN4HIlpQsPh4p3Cm+0TzlyM0ktVyvSbMxne
J0y6lokVMSfTHOoJxXjaRCS5WUOIZ2aaix4GpxV6cq9mLvDc3Q6IZds9v8PeoGNP
7lDU6FgZoVsj+N2pFsvTOfgQbpp1JbrKKABPWTsJIRQsCN5jUK4Aentzev8Wdh1I
YEaIIMqALaVjEWKRpQGzi9T9q9VVu+qgYNhh/vOW5LDE1yr/CqsMTKWhega7H8Ws
cVBjqomwBi55rIDNGnqh4Vp/uYloDAZArTZhE49wPTgVlOY4xE0rzwz05LT7oUMH
4bWi0N06D0lbVmnwz/RrUCHSxE+g9ZZ1g6KaNpiWu/+IsyapdjRDZN5fqFSRT8S4
Du/ILHb/figtOB6nctprRTMKAFIve8KNNjuyzh4D79sJZZ2KhtQzzCEho2eDTZpx
IkK2e4GP4VC4Z842MQ9zgaC+cIBSm4+++P6K9+LwF7bqZDQRsTDgSOeRrNXNr62N
/HkCc0+AAzgC71aPY8pkOOww8tj9fU44wsKffBq448KOs5Xe1cAyzg4Z9m9gxlct
jQdyYMjb9PRhuogCCkTfa87/mxnKKdzbxgLg5mQgxaly1P1vBeywMxglQVbSJ3fL
ipb7xixYs+y3/ZMO5xAa53jLAu978I82citoD5f8ssWSgXlHhpMc/7wWTvHexdMm
KxaSthl+BhR6rQwIpW6BE27GxG4x0IvMB7rfXha8qGVACLeq/o1ObfR3L+uB7HUs
dB/4l6nouyHRTUfK9Cish+VLjf3NagmQlnccgov+3YJQteITHyv7wQ7vfQaGwzma
X2Qt89Y25e7V+tcqiv13yWsNn2t8exw65beS75R5HxR/TN8QHrS2ZzJBkVFpN/iK
heJEt/ec4AaVZurwf8GwjkaJHRhKWRKvHG9yEuY7SvwImHXf7wxIhMgyKC7z1MPF
53EpW+v7N4H48aLpKQ/LQs0lDfn/2UqMWvaic1dojGIScLFsDeC2TyqT6Xv4ITii
rT7H0RkXIW4WSiTr5Oqh3SfPkh5oQWD6rNwcFKwdQxYyvnWFY0H+9wA2WxbMqkLP
qO/90ABZS+h9q7fH3Jw8xkyiAK/gyJBYtfpR1maccT1nVtVs68cyRj+lpeCCoRWO
4kDWVrI/IkSEpL3yY6f6roC17/dwN0ZVT2teJYOi1m6XnYTNOrmFLJHO5zwRQdNw
OlxRioMUYaTU/hF6q3WvNxfblUpm0cLg27Kulop6QPUllKK8E0N83T0diGJR3wIy
GdtJsaeuAahLgwK9ytd2QCe0ohjSZDQUhZ3ArCR0Giv1zHaBzYn70Y3apP+5biZi
xRmXEOPbksrD6oWQ6GNYBI2x4oOc1JdIzu9+QLMVHwEerr7/XqeMxGNZT9VFdoVJ
Mcu5vfF6RcfhuU0aNmxelqf4C3GK7fxHm1F2rFXQ7sbOhM/dN1hADxgnLWs/oFGF
Zr6Sdplug0sD8d7GDXRIk/q3vAh71RspxDCpgzcOPJUs0ON3j06Fj1N1no0GRadY
NIxxjDPM8Ij0VaBqgAB9ycE2VujPUp5XG5dVmH1ytcd2KRr6BU+0YL17Is0lA2Dv
1h41lOo0PEjfEgJv+0AyCm9pymlJpIWJGsQCAXcJ1Toryx624Q/aqCE9ns5GKJYg
P/IebdUiE38oXlUYVXrjosfK0VziN3/MO3kl0THmyLWycLyvLhij7AefSe23iYNR
3u5ki+YEnRuy4USAz0NeH9da+lkcVG6c5ny+SOQtVXN0kraJA89OoiaBs+/QvcBJ
BVsLIyY4miLXi3/x2uOlz942sISxG5cUEzDVpbupNAOduSs1IZz3KzYsf8zIO0Ce
OJuPUtrZvNhL1OJPv1H1OnnWgJpIbWDLofHOlQZ5ZHMNm2bGhLx2xT514IEanDVf
DtbNZHcy9x/+tpjUh3p5fuqOgIlq5Z50k/wpMPNmLPtOJ9P6DCtaj2SRDj7v1+Mz
Bzqp8y5O2gwHcB2IN27HXya8OFH3nVftJVAUOBQbZioVwYUEXC5N4MmFekuwvPF1
fRH2uT4WaA7kgI2WCf979h7ARFVI4Wq7qBPSjtb+jICxGhN0yjEp9S6Va2UtwYLz
d4hwRbQ0/RZW7IkPxobxw/BKqAWeJv/5cAZFxvp3bp9po2CGFkTvr3jjvCCZ4MyR
QBL6+9yqfebb5EzlkqHiV34CUt7wjWswg4lillnsKZWt7ATrVUWjGaZtxgSm8ffC
0qknqQ7IETGx58HvSsBNSAPiU7goUxhiyQ+H6K2fEFAUHAuVW0jfXbuMKUiHf4+B
yYCY8mMbAhzD4PClXkp/TuOsRmHz+lyzKbMMxcnEUG2/L9Alpk9Bqm1DKhfOG0xA
472BhwDQHkipPKAyAk/znJL+VJy+WrcIZv5gECrLVBdYfbHJaEpiibrKKd6UCLbi
5Qm8a8IwXYUSUi/4+fSm5vTLglsjtzzdpRs22zQzlKN9gGeQ+njyB2UnS4tv4q2r
q3EV1jE5jDN47UaxL2ZXqH5D8spPePYDOULximvBsOWbW+xYXXhSUspNAkW6mT1B
02uDiVZfKAmmM50HyN5r12zeWEjYP/w4YDleoeipWCrsADGGLP7cGRBWHkPz9hfH
Af3HbJaX9T2qaLTDmmANkdcNxB9Fm71INg2i2FroXEtMFVr+UXJ8YotD91Zg0aDF
fsXYbkT41n3ZyVSEmTpD6YxYXJNMVhiDinf9t8jx91LXRFc/Pc+x1619F1WgXK8Q
8VT7w6h6qYpjO13ZkEOw5nTXHXZQdrGYULCLvtikIZgC/Ze6KuXEVGtBC7ROIcwS
hS4XmyB7s1M05Wr5VXU158rSvnFdRRFGVgNs+/bIVRfKzcy3MlA4TOvBwOfBrcAi
5SwhYPYxotEhMWKm9jVnRNAj/P31z1R/16jSB57hruXm3wXYRB8oBQBjfl2yROAA
/OQ6rrIWoAD/Atv7ISQ8lhZkdWYTdQjK9ePxLGw4JQ/bKF5EcQU1//hMRBfc0+8R
G8PK50yizHhZodHGZG6FPBfIU2bsnxQQ1WMUMoB9NrHd5FKzWUodgpsIJnvvA5uw
3eMx+D90wU1tpH5/uONUBQZdsAgOdtUvJQt1mLJMWCBMD+4QXFPgOYNbnhiA06gl
+7Sm7+PHUVxBr6byZL/0+C+Y4gSGI/TjPrX9FDJ5HtfaRGng6YQor3zoQhl+hxS9
C9dePm7QVGN141g6vg/+keLSBwea+VXtsOy9RbT1wtJpyh/sDUYle3J7p/G/BhNN
noFvU7tJl0iGvMLoHuebh5ZHbwWs95lE2VVJ1YswU9eYtflEQ/fAtkDErpwAnhkf
kJI5fw/Mwbjf8cE1zQS7oZ9qT80ER/gSNuLkhTH4L/69t3X+mKBSYEJte1z39as1
j1lA6CIYacU8J4Nlzo+YdtYeEDRNifUw5OTMU9/+iKzq/PR3bJaXWCwdg+4jBE6J
aCGdExwOfMzgXOvZmdhv9r9p6Jex3fy3/fU0GXGSdnQu2a6bj6IE4mRlVOTk3HWw
u6M+mM2yh1AzC4IJ1dovmyV2i06LsYscoju3P1nogjTVfvbk/oq8t6ZmHqvOlObT
f3pAwyH3WWR1AJdiDsPRPGp9W8mSNVKMh1RotkdCchyrCT8grZ4hkk7o3RH021xd
xuDbfR9QvrUHjDMcbow2nlVGTc/7XxpyTNI+sl8RSQNtDjdJkNTjuA7Y9KzZ91bg
APbu4v5swK5WvT0eowWyX23uObAc+LPqCbIIE6UC1hP4lTzrFh1pZ1Sby3L94v7o
etuX6Owq3rBsl42JkQCnUQKhDYxuYSNK6d3c9ZhNuVEYCHrQMijGKE1XigIcXhY3
joK+7a16be8Czcthwg/1iStPORoFDenpiVN+ucA95TJhkibebABJSWfDwlMx5HDz
5n9SAaN7/s4sLZUmLq0k/vqEp9FvH/6YU7nFVdgC+EzS3LloCRVbGdrGPzLm3EPU
y2gYwzVnObN4MVA+3CTlwGIjKw1TunAL6hksbn63xKtj+8EqvqE54ptHpJzWWu15
i4i4qtbnQ1l80J9/Iv5B1FXMNmXVzmIl7ZM3xNSdoYWB1bUor2QjqzjXxZEgJ+ih
KDfKRqis2pXiw4YkZvSqD4VqCH7vBHQkvKuhBJFb+nYDBd39IfxRVzGdpu0zOTtO
KIYyhg97I1QyAFHxnm1nJPJbWdFWQrbUqbbU0b1HBkCCC8ihUh01vbUnWW21I6NC
SZEgdZiDIeACGJ0MCcqarA66rj95xv3MT46Kqr9OFPfgI8DdAvumyca+B2jV2Jgy
kPOR7B/NZm8JTStpbcOoMD9nHY3Gof3D+O5CXmruzBWAIvmQnE4TshvkhcDDs6yr
pxThA3wv3TAd8Ie/8HbYYPn0zKoEkna+HOjUfMhNX5Ff3RCVAg05N0XrgxcDmdBe
UTrB8mCbSK7CJ3pseax6jwr8S4tYCWmjH3vpG0kdBD4lsHMafgDFPvy3JVJEgljH
sVBEm33nrsbvNQf7+0PilpzoRpjuzgcHwRWkJLMoFYqZYiuaKQKlIkIoCBvmeL7H
UrOBIb95cRI0B0ySzX2wWiTr+BP2n8MsVA5kO6bRkvlVEB7nqSRM54wArpI+uNVz
NJXAnxsrMzl2L4csMsMqRQfyMQR/7nzTRLf7mtXmmxVkH70TmxKM5Y6flcXQNNir
9q1u39yc9JyyC2OXbxu1zDNgSpgw8Nq8MMBgkRmGXaG76mTiyfLKaFLMivycpZds
s/El+snuC/UQmIkjBTkIX/bHSoacQfRgEFr3kVK+IkRbc+dCtJdCRjC/ghpEmQOP
IxGwExAwFHWBPZMatmR5Hy+XRkTwjGk1f37U9RZVNug4n1ZNFfXwnGoG+FEQn7rP
VrZhZDvRaj1CeqeIxkI1Hk3+LHsbphvGEge07MOyV3sbr21E8GiRvIuZ9HjSxxqh
sBwrF4tEkcs0izGvYZhn8FJ85UPreGvsCDEf0L3IZMdhEJjo+k8TV7GQEDg9MD10
6rOc1YFqWXlZMjVUyGpZqbFZ3vXcYqUkuA1M/YPshEqHWFrGrBH8RWePRzTQoP0k
v3E5nMZw3YhDl5nURBLoMqPF/Mn1fLRDS+NJ0hHu5ADx2G4vq36yCNGwDkGI/tB0
9+uDkKWGyGo/FZMgLn5htTC62zih/UPalru5ZZRAwHBhQLHcJ1c8Yz000sfTbJ4Y
gUMq7Jlej+vreIDhn1Ri2vmbdszFldZKdeu4tcyVLdxCMm/OLTWYPnGimMM1lxzk
v/mTegTvyfF1TAwoFJt6rNYaGgX971Kaf1EuytA98B2mgB9okwKnmatQtUPxk4iM
whXDoPpRWemdgA0Am7Inv0N3ufnhQGyXiaWprbxPUWOJi/H+N7OmTczcbmkNhV4H
dWYAFHZaHK9JjoOIKoBkP2mcHGowCdMOpmJV1+DaWcQ7BfIJul+CooUqrLOY6MIS
nQ0JAhrkBtodsH8FRbC2FuHxmXrpTny4JRTjvF3R9mrLKlPmigJLmVrgsj153w/X
liXWfeptdKjpl8YGMTRj1KPduMazwJ0ApRqnte03JQcrAEGqL79Fe4Y0oRlR6QZk
vWbGRcFv0UduLoLTDnoRPky+ozRv1xKoevuNNfO08AhC6nJIcJAk+kJTHzTGtf82
jszQ4E8+S/uT+DM8e9DkPs1EnA2/i46OyWMXYIh8lMqDP7Z0Gp6aw7e54AXKhwbL
UegaX3lGO3Vd69rtd57FDqx3pjXPPog+cHlEVIwFFjL1msCOlHep6RVcvZP8NS9x
7XKKoyRzRuruMy9qJU1WLY7JNo3sn5fqw038gZs5cBIB9Ias0ASokKsG7AE3KVhN
qXBbv7V+ffanwsQpzwLc7aqYky96lLgTWTgb3LiZ5C+LAdc4fGJFxbfo1+msujzn
6T2iflLxh3ayYwg8e8lybl6552jYrAcuRNk9i3UFDykm6E+F9y4HK7zRBnabMekf
PXzJLAob++VbT0oFNppQ9EXNud7RlkA2x0baj4NYkB2hynojNkzOWPec6h3BYAC0
C8qUPt+HAV4Or1JFGSNBIYYAvapGmvbEv2jQkeEqhLWs0WQnqyzcLM6Rfnqhb4Ro
8PvC7dLaa7l3hGsVsagfPjd4kb+cXZ9zqfGQyaiig0hcdD5bE4/C4H7W/WcJGY5j
tZVah5UqjU96P7JJTnNdjqnAjIvDpUQC+wSQvesvJL/Rm7E0uCV1FlE5uujNpr/v
uXPwe+b4g/YKAEeDTredTNZj4R11J+mezlETEJic39KKrZfI/GStXClFXm2LS9N/
gHSpAVXcdtab48SBO4z2c2R26rRPKUzUClK/nd1/dPtKjjzm3Mo+usq4Q7QsHsjJ
uwNZ+eZIbeEv5vvyUzy4hY4bM7CKOaFhiKF2Ga1PDWIhLI0dFmcpXQH0F5qptPNn
TU6xoo5/+AybFtSJRPPkQjDM9bAP1R/PGcuiupmG3irZJYlHwZjDZUDOBQ0ntaKy
nElVOl0MxVNojqsNtcKL/bkA9G4Xmh5H13Eq4n1bTt6DE7Hf7FZ9lJyLtx/mXOoA
4blHispSXTeEHfcTCjwHaFIWphKQ/zNgC4TcQ9WxWIOrNH8/LgLrcLGuG4kelKFq
oqlep+En71AsVboj4y/bMWkvzufD7XYkROFOV1qE/t4pTqN2nZba265q2bWhqxD5
xxZcTovVMS3TRrSGjb1ZXVOiqt4XUHyWFWGGREBL3Bcyl8nqkk4P4alaQ/ETXYg8
8//gEKSGfJFe8RSewkl3asKbB5BnhQ2nUdqI6Pfov+6PvJX0OLyAuFmHb+40LHFm
0zhqLsmDUau64JUeNu9Ip2Ex1d5EF5myDTjwbw3Qgjmu7MsidfJ+Pyh7R/gW7k01
xOwwbzJOp6nNQsCx6tvWkzzkZXMg11MLZ8YH01OuHvbKjtRpsMgIE/3UiTyD/tbr
tax+Oc6AXWvq3A5q2q+krDxKIhEORj88ikfCmTaBecS0JFFOm9guUbIDhxKr3ytE
0bg7Cmep1/uXwtDWUR3XFE4N+b9M9Jcz+ymBb0Es2z6jAcwDcMoCtpZ6F9nm+tMR
PSDIt4W4qM8GZJ3pff5NwVIVgN2Xfxjgx0fxzgyeG0mmRoNr6xPWfI/hDXtXO3tH
NhbJoyDW9pRQDCubQbcJRQ3G0mFSRz2CB7AEnjMfBoQrnYtytwl1XmSIIIcemSp7
Y8zib9yh+jVzVEpRHRuQUWrByVUGAMq2TL/IE7KwqeCkFBTFmfB6+NBm7AF/3vAa
q1nK+uEFbtUa+oRxOwm4DcHTAYMn1QnsM9tOgCJ/jv92yJgvgDmRp7Va4zkJYEAf
9lg0oMQ5KNEwVZSfKlErHez2NwcE8Qw0NXBlw5rx/TUJ8bbVIp1lvBDFQ9JKkL6T
3BRlp/++w8vUSoNh6c1bAhhzaahlS362kubeXQgx7O4ghgoP4C5P1EJQ5I6Cpzyd
3DXxj9+bz/aTVx4JTyG6mdoPzUBLsnFbuson8gOMpX6LzQXWV9CQFXAr1W04Ioha
5YCk/0dekxiADhlElPRhS1gVzoN2RwGuZ9pPo7IIJ15ENBM9+ZsQb5S72UzgeQ84
arEhxeUxv1/hSBi4Joq2pfon1Wz5xVH9aOw7whyhQ0A0Cs/9PXnem2+EYM7Abzon
d3Tl5hqq6k7ISsUdcg2rg871OmJZM9WcNlkjibpS5/QoUxV9qTK5FoQyeebgAHnZ
OyQHfrWB9R7nFN49WOirKb7wQ5YfG1HYLnBysTdZnyEEKAZW23vLwufh6mLV+DFt
psq07eyqVlVEv7DAAGVDaQZYftvF297yMEIVXO1BwQi3Uzr18MKPIcFW0AEP+PeI
GJFLD9LQW1Kb65nkxmby5//yXhKXwlkLEDJKoZmC6G8EYUErn10EUQt3UWx8rEsX
ESqdBYc/6ZIfBJ6C3R1b9utinG8PnUl9G4vNpmzG3uCdRh9WFaoa38KAai/tH16I
oS9tYTX2BBUpP+G9cQL+gOgZBXajMjOqoGNncL3yFYQfUpFhmNk93BWOl4lq1xgr
bEcgcRRyCk/qDPstkNOXLs2miz8ptu8M2Sg0HFgp3WoqYzkvOJoo9yyUPuxcsN3b
AtLybFQLhhkgwWZnV84+3jrihiCMPuGxzaN/N1iPEyAahwJi/ITELHsmWyimKh3u
GPTqCPQgha8sUQjPkvU55hy5yVH2h/YVI+4loCBtZ5FXchS4jJa6b5oZj6t6ufck
ryapxbZ9BH8AZQKNG3KBSPDLNyuoj43OukPWl5fdn+CTfmYyiKYeW/dzXuDSO+GE
lQLPIxvZcSZyLNwMG1oINNv9zJ/dShVppiBwB72qeIvSBjMNVb+OyHuvhlINmXNK
4eUE3CoMkmU+feToi7FwjYEjjb3v0rp2VPF7P6cf0bTatDvxfNK8OkEUP53PR5wd
kn/ghBautnclK7ZuG/yUo99knUfzQlT4oCwvRDVLX5VPzZh1/Jm4fd++eNnRUf7l
habkuTt0GamfK3NjF0fSXSS+bj9Qstmo5+onbCkTZZJ91RyI9xsZS6/OEwrGKFfb
NYO/AfYU5Pyefi1ex4FFHlJ6/0PwyJPObR7suOEpQeVzVrfWf0GMIjGwft6SZBDr
rw+GpptAdzVbi01eah8XvKNCiR6gSsO32iuspRvEfam1YCXV7krrT4ca8RTNYLi7
KD9niC7cfxUl4Z1hlCh6s4IpZQRaq2P75MvUWrYbS6X8Z28ZA9dkMUhUw1UAlN0l
7s2LU1khLwlnuDK7t/XAo9Yh5hvki522bfjiunAW6/BP+LVUIibmx/Rt6TdmPfIf
h/OMPUFC1dAGMU/vV/OLVcPUxnRymq2ZX7ZaQC8nF81JyS2OFz6J9C4Thyhx7fG3
2NWzWAlCvDeXv7JDG1AnFH9NZ5i6uQTHKzSuozyI9HxOgyPX/GJV20+cw94jawYR
L+Cc+ghSmsTJM4gr5y84ZAdPncUhhdFkM9F5hc1H5G7X6ZRnXwtW283Ee9bcV5zc
CIgo1/YtULZxx4x/svEmhgfG3NghS7JyPVZlWTcnHxkhlg4OCAEPlYbMOAYSN5Kq
jQPIwq5+8qu5VZP08ltUNpcYCQDN0RBAbmPyIq3sm6QPTmETW7j/19dI157/AOop
VoTYm8nrU4PgZaJfhwY+az5w+ffvW6zq1mEiQAr/6FoBV6bvHZuicCY7aVa+wdF0
UpHgb6EvCBxNkaQkDwwqtsJfeDD1IJtMjq6Ds626KCYqIq9lcSW4Yntws4dW6yBY
ObMAd6ycn7Tm3WkpuNXPxRwoUq/j0iLUujCTTuFZbHKD4Gq/NM1Yds4frV7ZY/Ze
bsskcYQF07iqxQoJAdlj3pC5/XN0PMi3CD9kLJg2fWjo9qPuzJklDlBQ0X+dqWSZ
vWWUWQ1g9vcmBM9bYueBi8CvAsu0Va74EmbHnNcocTd0oVvfBP+mcjBxjkV4h6+3
FHyxfOZc/tnEk2GcaRluj+YKdXt1EW/kcRvyu0yWuKDe05EBBNaGOolYyHHSP2JG
g4RvDJiVX0lFcl+wauwtIs0ADO9CGw3bVqOlXAmixE5fOqcQiKb0PFwYNWPB3vmr
8lOu/tU2+1ssq2Dl7gHEpWi+ZhFfmFavHFrfNX6hSMU3Q/WwLykvfhqroTtfhuYT
9Rusi3fRXK6zGo5SNopMESBHL9Luvv/8Cm+w0y6wSJWBTHeQX1UXWX3jAiMrSo15
1+8UeairBp3j1Ol4R7a6Q8Ded1megu7Oz/7J36qFd3J2dNy5oOSBIDSWeI5Q77WI
atgWPnzYoRNtqw9C1yjGbpV+PPvxwuuC+7E6RyULgXxcjcV757UkXGisSR/DfmUc
Vs0eicE27ycUr6vofu0IytWgp7boinFmZ4o0IEe0FMWK+o2YLhZpArMiNVDs5sVq
hbP2zydi7W3XaYXeEdcNO66m+bX7ghD1RKpa/Q+0VisKEj1hhL3q6Gbqv6Q7bv+C
4U4qa8DWS2zg2Zel3fzipuPHkMljx6SNbFQ0z/wFJaLoaiT6Bay1iATXoqX5oX/P
bwA7Mkif0YJSRLvmswE06ugO+ux+pnRzOtPqVGDGs5ofFzCLGobux4KsLUheM8Ij
swytlHuQx5PNxD0kGAFz3YnEccybW2e5ypsTluereJv3Cmupd2l0law8FJ0RlidH
Om3NqvjxQ7eUv17ymj4ZqCrZ0yXWLqh9BVCkk6WN5AJZBcXgwLPTFivI3gVOLnpE
j5j/xNkpw72n22gfli6GhnTACQI4xR4wTflVt/eYSYKtpm39KwmcIpelu962FO9u
Nhjj6ODGGa1ZYaaSqB1DjdHxTNdCNkYoTX80JzpQWYiWzyninxWWsbldWFcPOhz2
8U85Bf6G+/l2lREaDzUqx77Ee85ykynmbuuWJlfLv0bzpiR+d9gE0QQ2/NoT1vrj
rdcBC4UukqaKbhI9Hl5zQih2SMhO8mcN9W4077Hc9/N5IUH5ZqGYyXOTjDEE5WuP
WPd4msLeFD54sS6Q9FTTOZzt5nuBvo8NlLfugwu02JuHzswPEs0aDLy/9RkXdWqD
y118zaK2ISO2HQh4hVVRg8qnqjg2OuauRS+QmlIl/6FTDezAh9a5cntq8ldAimBO
F6KTymUWRHa/YHNVgz3jc7EIri/Rpw8cQjCKt1Td9xrPfdUgagkUe51c967UuCkA
uEEw7dQimLIp6NIRU/Uf7jyi4tfUWv6j9NEk/XGkuMFednyKnnrfWQqpHQiGnNSb
AGDB0igYHE+JI5w0Abx2uIsEREB94b1x6RV1YdvOlCRC/HH6gtVarN8NR3es9TZP
L0MT463GtDryJLEeWxS8p5oPskZOoe8IIuI+pJEgWUL/bNUIgrpHjbYuLNzyZxWK
1i6vIScw9Iz3Q/ssdUSwctMzFtdJTmSD4UvkrsYVyN/8vvqiJPm92NevhyoC8EGG
wAx+QkyRnmN8xHUWnn/KHRsDiX/rYAjEJ/ILJ3pguDJqzN3V2jUDYugK/SHzGogn
2zR7GlzexFMnE1QubS18/fDZTTaNP0T7PCg4uM/zTHXz+6yFcn6hze8S9Q+J9TnI
6DNwjlypxIS9Jso0BlKXaH7dRxPqkRcNayjiuYEWDnN7zEkrkb29XMW2heSNAE2l
wXIwZsrORDLXemLaHHUJi0GZa/lKZckEXX8PCxUrdSF1UPPH9ezdMr4FH9Wp1wkD
kCwDTlQNY/TbYpu/P30Z5mThC0leWPBRdmkEXW5GfNCUia9FHXKG5tslaXSVzGVn
JFymuQDXAQEaAYyqJoqWptyeXOSTuy8yqGYJ8lznC9gtVDLIaoZE+CwnhIqAAsiG
AGCMc3hycl8pr1NRTwId4N6bBldr5xjLsxCNs3JiKrOK8lF/GIM00caNCZd1Csy1
Y50lD2H1mETotJX2cCYEsGCsaGKJxqN2kPxW0cJytCNra0DB3GHzDD2nqBIdkSCV
+NkMXI1Ai8sRMtvkgTE7ED/lCftgBFY0L+VMYUA6V6QDhHwE8L30QNRww/Efri1z
CBgExsP6rUzLvqfyp91KPKpWggOx8gej66qm9CIkQMgppvJvm58W6pQsjOAiwFAR
+p7lzlei4ISufo7bmE+6os1QBuDjMLrliYVpGVNg/wgV51PfG80D9YzKUct95qB2
P92UKPmkX0EsLfnqw8mBzQ52XyxPxiLVrETZjYlOGXpIVoJxaup8fud2TDzu7QO2
Po2QWRVVJYo0IzmHFSm32iZXDw07KL3fS7MNR6pAGx3onPE7ZEcEbBMXGWmqF2Le
axgt2Q4Dq7Mtwjbp8mD3eweRkBp0j0erHq+w9uDZBis0QgixrS+55hTCiyGygb2I
TLVk0a3mdCsucaZ2D3fbHG1XMF+20oYDHd+l6moUKm7gpoh1Bf809f1Ry0T3Z6/0
rPeJSEj5teBJJBDCP7Oe2T+5edrUNxidCjH5GuaGKTdKJ97GhY/mYB+IKYJ+cjx3
gV9mknOhx2xHjryplDNMWrlzxrEhgUZ0E+J82CxpkNcca/KtZkEYl5xfnxaPPXKJ
ULmswRZCHGfkW/oIkvtKL4jq9UsxA/WkdowScb2JHkE3EsAsplz1CTrgN34MuJ4m
uonU0a0XWOv5LEeHeh1/L4zW65QVvbyGlzMsmXadBGjTfHMLEgpmjLLidrO9X4/4
cYPr/BGzg2FkPkiTx3sy9qUGV1paK2nltUUKHIfwe7tryjmy9mKQJ8LuJcrxIprW
4gTXpc2O8EUlY9fpbT1NfC/OMXuHnL5Q9htbjFSdFlmMvybAJqB9Y+CN+v9qtXb7
Z7nYsLce4x01SyIM9C2tEsGHaGFB5wjmipp+i42FN2DOMCTFnOhFsjXaP0IlmcRQ
1q3jPj774bkY1PsVqBGStvIwf8Lbz/8UxWOZA2POWaruRudRPORCk4+16qMv4SsO
H+HILeIIXgzhdbx7bXwV6KbMjZPD2hsh8mlok2jQiGtvBafrJtMwqVJslbP3rpOg
1G9dWWROMczoIE2W+rLpm7pFDKj0Rvbb4Cb19FEYnFhbMVIHmJBWkokgGOfveqEJ
df5HH3J1+iIo32DHn61MBfuyFbo1NdIYYB3cj22v0gWIPWyS8l6UWzotrsZ979My
rfg7zs1XcoMo8n/+g0v7LkfGsLqH4nxlK0pC2jNOWwO5lNhkLRYSKT6h0MaBTaI1
cXgnm22w7Q4lb3/G+tTf6C9GPgOmDvqjtjnJvwVqOyitMHFf/VZ83+D3dJ4/i2H0
dPjAccSHn/lN1FHzJS2LOru+MV6rqxyEsEo8yVstZruXxX5uIgZvQfvoQMTcgiPH
nLZO/xTOO+APNMq/Zu/LrNXMkf/Q+SFbVLP55qPbtZ5Z3/lkgeKYDE4fr4ikefli
gNDNnbMP+1VfVticYdGNoImfjvHW0RWONRKiPgWJWK+v8rW637O7Suh1kKVcRq9G
izSlnF3wUPew6P0wExUoPDUTOJJbnqCT4Wqqpcij6qoWbmWY+K1nIfOexduCyN3M
LyCh/TARE7X89wDZX9aF2KiidDV43PsRXUyRsNAiAiUPjNpE9a/WNPsMY/ocIGeI
atXiLgQVTf9E8jd+I9OYzBfIu0DZ4iePwkWDdk7GN9g2PTTTCT+VKfaOQEIs8x0F
SOac4c56VQjKXJe2YFKgy7xKMpZolvdl5C0NCXcc5ZUOgYNlPqo29I6eUxTJ4Sr6
PCPp7EMWUBJHaZ/CmIJYVEstuGiXQvTfHC2A3HCagIyJphaOWGm83fTRQUnX9ugk
KRZedMwgnfzslRUFYN6v0uQpRby2RE3XfFgLinyMzuSHDjCDWGd2rzNCNcJ050wU
kAOJ6GqZKDHMeq/qFIycHKLaXRt7fEiBHbDwGcciMP5R91a9LWu0JFap2DYQs4B8
DZ2lPc8qowxpEDBwTiWCJzxe8UjR6VsPpah+ByRzBc5tuGdFSManvBOXt0iGhNi5
9J4CVUbImTrS+w6Fo2SlTPPVCHMHERQLXuULGUGfM/dWFLsGKklFScKSEacIoF7O
fJ2Sj7G1b6ZairYwbcHcJEBlxVu1v5lbYthr3eTHy1pVfHIWcmbkJVhKs7a+zalC
We/PQdMly/rE9zscMjctEqlw9J0+eNNFAlgqFHmZJPiV8pHhVk/R8Ubma9lhYkFQ
WYYQBa9954uJmtWOvAiDXv20xgYGgSqHRmPTtv40ldZzfuPGuw740MNBSBfCXMj4
N+IUYrj/pvEmzuOXWayOFZ8bYY8dskHRvtx15GV0w2h7FtHze9nGAE1fsg103nUg
mMU0h09erQy2UPeu+sRQ/LrKmhBYhoWvLsAF93IwrBzW+t8P1RBxJbcx2azL6wEd
SbsDiEsI/5NH39B51yFHRXQWPVBFpeJQhhZWgiT30DT7gr/5O+a16yigfRNq1abN
TetuoMjX3eFqRd9wZg/nGvHNbz+LeycFj+qtYSpFXDT0QAuvBhuXZNjCBmwvR9Qk
fPEfimh4KvmSz1VkUpKul9o9qdKBnTSEh47bUswMqNTP0JrRmOIf2Vf+8trSnx0G
6OQVcZLozLfggfNEtBZTl4ktrDV63OPcJEKOwECV+MPyI3EV6zjJTaGVJoi/Wwr9
I/xsid/YD1HuN0wVbYg9KMJw9mrg56Yc1KLlnM+CdzXQG/8wVxzwRnAXV2uwigHL
PY4S6nCQ4KmK7HMGTtoTzd9C4wPQTL78VJXuCuS2I1STchGMsDuaNtUwklhL1xR+
abyMj5XHRHz9vvtOhqblyC9tyVi7MWHwCS3UFWZ5WYU6RJjnw9A5QlCwCZdiVEAJ
l7ZLB4OOHEtmtxVmsu41p/YfDbzTk1cyu/oXQTCFcs5ZTix5lQSMAGtcXroQNoKn
hiPqxaqPijNQDAjuZ2MRydVRBVOz3RM5a+e/eqt356FFSpBStvpU8/G5kyAPYVYr
4exB+/A7nEWTGGUAx1g4sv2egubzgahepWl+vFs/inMzHis6zfsnkG93UT+9NrhL
m8XmKPai8ATRCng7Bezo/DSt6ioXmGX5BaSyUy2thglf0U+i0wdzlMg5qlW5FmsZ
NfssvkWEVyu2//56mVlyPpSJmGqZZAm/nZBemeeWIhI6paXLIf53awx4QHSCG7fp
rKZ//6qwFgqjNzzATt7wmjYh0izOz4vW+dfHOYotkvaq8Lr1OqjOVmZF4j5wpPao
SkHGGW7VT7jocN+oCDUo2JhMI0U8TkhL0y+JcR70nokJi/cZidG192v1alE9mzDU
4UzjCe3uoyiazqgz4E0z0Oc++5TAtsPLXxpS+I0XM1DA14NOBQ7gP+/k6XzR1zdf
1x6x21MNNhUMxAu3M2bIjFpznHLf9byAZXuMPT7RV6uMSsNpC9fJq5cgalVHjuFG
sCZvEof/EmOn9pHWOwstmtXQlBV90i8uM/WAGjZPGqcBmso/DzvrpKMa5s2o34k6
sTN8T1M2ijdkWUTFgcy5Qbx2S9ZxiPmZ5Z5927HwIvdytQspjHcV6bHnVtrzPBK0
VS3GJZZ/CRseJzUcqKK4k/sV+IGsWGe60CkZSGljHbS1uHFeQ8Pl6adgPStj0PhG
/XqefhorUsr9/wp3u3w2Co+o3oVzC70LqBg8So2XtL6WSyFG0NmjCt5oejTd2yN4
NqJBjxxxrgwn1bx9HEiLg6X69TLmznmBYYAblxsEgshHRZ31YFGLUJuhi4riHucK
7ZOyIHtpM3s5MYj/15lzrqgUTkVzUe1sGVbz3HlxpNUfJPq9/M4U69JKtLfyWUKp
w8eTw2YuOjyqpAg1tLNhyFYMM0tH3xCbsZ88ZeFbBEJdDHjdoTZXy9DdWoYyW9rA
DddSZmnoUPTWe+lQXVA/b30N0hnpXo3zAeDSkzy68OPTQ2bXZ4Vy6g0EqPzwETTn
kLFii+i2e7TSV/Zr9LX1Mv8YDvePriOv824HQmZbm0zbV86+0N3J+EOYF+keroqc
/jTk3Zl67EWZceoHYE9gncD9tybldsgQxI5GzaBfT9dMtPCKqZKTB68X5ScOkg4O
vTxdlD+RkJ6wzxcQ4OGSa+7v/f4iSL0POEQUdQG2fOv6+oHnZuI/UEVA2AJo/qDU
5eyzwW5dnAPZmfFKDBJ85ArC/z9G+z1E9CWsg/tj6ChscSndB2Hd5TeO/N0yyy4P
E3CJSz6IY3nJzB2J6imbyrhOujtS0mycLB2OCVmNevmCyAhAinCNrpNG+n40eIdy
Rcyd44tZc7z8zLKmiBMIJWglhcZBuHoVxIKXGbI2eMyoeXncbUIMExoHUgrHEtCC
IWbgLc9obeQHG7upsHv/OYemqLS1LjNdaLrmdQLf78YdhVb/YFI3FtNOoBd26Zfi
ztaHnZu3ryBGAkmGyXnzJ76EgL9RCf2jVcmV8bIwoZYbmbiHleTd836bTQ25x/IN
rP0h4HEZxDQ7dZQD/CUOKgmwZj3F5bIGxGgtuup42Sl+3KzNvxH8hqVmnRWYCkIj
8rYZlEwxXwcz5TCa1XIQneukmGbYPRdZsS1+Cumi+XxYTUrFhmw4eQJIu5TMPhps
GH+V7LJnwNAjzGzA32GXgFML19xKS2R6dBJEq0gGlYBZzPb8RjMPRFBlXcVHyvYN
rg+X4m9aP8g0ZtaeuijlB7dZtilCNSwnUWvPGEtAkSAEmp5j2EAIgDBWIPRm4H1c
Ja2dVvgSkEd+u8B4blF/pibBLsQc4yhUnbcxaP5K0jl3i1tjAyYyYYGTE+Vg+DN9
X5y4/fx93daIHheil8al9lxMBcG9Umu7rR8xrbCmJAtHy43W8dU3mHRwU1OzZaxu
Hy17yKlXRHC/j1QuKRPgDevbzfPkZ0r8bQDefR9m78VLamz/HiXmoqPc284mYTw4
5QdrEmOOYowmqlN7acNalEOhxZ8DeoJofaLx8kB7RPzpMX+sFE29eKZ5OmP1VfZx
Go+GmMJmT8wyjtjgEsYrLDLD/SJisw0Ad5HDPtr6t9t2v0gz48OYLv7YwumzM00d
FIHWlcvYA8PV91A+4fecay0t8cnymPJ972ZxvwlABiMGnKIvP54tJWQssIo7nVdg
PlxWwxGJXOnQtEYodJOJEXzMKuI6SgQgzx764f8TcPD/UOlm89H7Fm1tXNPiCga0
uQOaIrnWWVi+8wuwY1OEHy/3e1oHHKAlgYskazWHV7Js/zxA7EWlvxfbZKwarCgM
mMv43gjjdRR6MRYFUPIq26pRkZ/lmCS4/CQL7hlk7EDIDKLsAFSjOP0aNFUl9wPA
FG1RkCH+lnmvdwe1H1tKMbdcE58n4KREYp6+kyWYDbwS/7RcdFmhdpKdWMiS9EVZ
70cTaMYSiw9tHYFiW+ptckJASQQNyLc7lSSHF3eQoFd4n55mIAewXBlLghQB32UO
Nb7NgrMLMCRDzjEMKwtVaAEqlW9MD5M3LJVuleJiczQdCD4j59ioNh+zdk7J8M10
TJ7XjRbBBYjvmbRqrEfZfDZHQEBBCUNabc5oLfUFkSO21rCTdAXgXGfTXiYn9AcG
Kq9YBBPspTGxIk8H9RobrP98im9rulqHoEMgK5ei+Yyuk5JMLQK2UBECn2WxFf0U
crdusYQqhgsVN39yj9ERMTQvT3LtXaiM4b9EMzCXJUO7b8XGvzm2er0Cy31c/Kcv
p5rDpyOcfrLfm+FAEwlkajg4GC5cJ+UzHhvjozuTqbUMyA+epcFtHCwRlNgrpJvv
Gb+Brn490iZauaK6DNPgbYqMv7Jfob6iYuQW3PhWnuVf8Yo6zRPvkCX5CAy2RO0W
I+UBEGXLn37en7jFHTwf6u3bj6zeriy7wIEncsT6JmF2f+hPyPxMM/y0Pd2GIUAp
0iL2MkSas67/ydBFH/TyQTlpesGGSFRWbdWQbGzEO1DNA0oOuOqNQUOgNoToWq1z
1nO+zl8Nmc1WL9tnwXBxE7JTNMHG38iEvQpvKsNA6vLGmx9pQDJyjD9sxPdBf2q7
Gw01XXEZds/BGITZns+hd3oCJ/IzY9vkV1H0PgF4v6UbXNNsGU3eaewmHr5VDZIc
9UqFDJeqh9y6WIGwWJZuk3kda+mkXTb+yf59HKcGT8Ufsc+C8hOYlnWLvdB3f9LU
hN5wXuYGruHrsAQAbe8XonvTsYZ15XfkF+lNoWyikXcnzsFXlJX4mRh+yMbL1dVK
yIdAtztjVWuCTFlSuFwcn29/vkr4hWlGHAXc53wzqUpKOefwgGpAkaR4bIfdVazc
MTvmoFy0q3QneY92SHFN9UuOJR2GcfMde59SEl8aAikgOLmToBvevS5q0lHAkmRJ
OsQc6CRCl5nvg8ASM/DD/O2r11S7S3NLzRISS2+T7l/MAnwByVVR4RRR4RUZnF+c
KSXPLX9hrQFRB4orsV7Zh33amDwbJhplB3On7HW6a+J8Oo/4hDhP4TaiLa4hxQJi
qIlW9L63iEo/X9VzzgKKVJEzuGBZ+CU26Szadkzar39Cqto10gwY8HCKWiAX/wTp
FN59qRvFJZwB1ASJ4Ho0uEqjEKkqQ/A8qjuAQ8Ovx6t+gSJ4hWO3tcpGoWhgMahr
R1G3/7yn8GC9/7h8rV8ySiLj+G8XlzQfXGLx5Ut07EbChL1+ybSt8be0K3He0/LF
oYUfx0KasNcJlRKB+dXj6piW3YxBLaeFxjJ9EwHg0hhSEzLQ2pNlkzTJNgrf6h/z
L+GYBRb+K+TNIU6yQ2L+JrC6f9A1bYe+lX4fvS5uxTqg8+BQe3bZ71bjd4q9pM9S
SI3+63z+Qe85IN70SzEMM9vJrpM3FAmQNdbstDUX/Ypko+GfyrgeJ4ZJsiBSEpnI
qhBa3R8Qq7riZEu0ycCu29mbZTRvwlYZKFIkyF69c9Jhl/fIDCqKm8/kcb2bKdNg
MXr2r8tYr+1gJ4j6rj1HoR5Tppv0zRL42URmuVt0KYIRtYepg4w7+Nv6OFH8GLN4
zziMX8LRJfJ/fGSJNRlkTUM+lnIKr8BsB/rwz3bK4TAtCll/OxB0OT9724bm8c2m
uUp7+1zfQ8ubNrOap9BjYyctcLGZYFD7N/xWyvGMaXbV2SSrOHrfbVD9zQiintaj
ExzSlm/uxeJZWGGtAR7j5ONi/OHzRkhW3TxgnIGicjWPqZWhNQ99qTFOmpaA3WCI
obs9djfRJ98L18As+rR2nXx4etFaqGK8IqkkOKY+Cfi76EhniWEgrfY6Fm9Rd5Hf
F8qZhgLvsimux62pc3RRifXpQDHCso8qWL8/RbT3t9kLdwqBLOyFEj3Kcdj5xjTW
tEK/2nr9roewliGFFEI0KxvPn3ZwtZkJdp1AZYbl2ZE8iW4gVt6ZPumqlV1rTvbQ
6Dy4YUoRqHa3NBXnJBy6QWHm1ydEcqnmwr1D2/AEfG8HUOZNvD4Ckxb4HB6ByBth
dAhvRLtCaUgj+KQZ2nsLix9rxUgz9vuQ0YBaEGkY5ei3HJr0eBKfBEHHU7IIIwWJ
V/Dm3WO6u2eKjAKnSPMuIBWq8ymp7QiKhire98zh9I/CDTnOHFmvu/S+eSUE3GkZ
hxOoI5m0WLxb4AYJm1Ykf0lbuRbAjLItaW66vSgT9XaeA/lxqffd2JgxGdirm4he
fI1/08Cnv9V6O5XGmPeocfdfjXjSp4vgJ4R8yOE5j5LuFQXY25PQrIrh+qXUPDMU
FHcqQD15ENdV1qZUgTPIlIkUa1aYJo7nltuTmgo1n9MQSy73C5/dE/pp3pzDBqgm
UeY08TALxw4zY4SOJmJeBliJY+557Mnla1ApcHh3OzvJhlhL+MUrUC8Y2/sdjrvw
OFMXtX+f68A7o03NkkZ0z95Sy4DzyMmXmPg42J1A9+yorWwTOFmkXWaN7uLrERbn
OsU4jfDxtmnDyE/OKU4g1qLwCJhRYjPpQquIQcvDDh9J36L178WjbBowA9OocGNJ
4SznsyYR73x0IQwzWSnxZXV4raxlPRRwnwBieORlv552DQQQMnlwpJ50mSgOttMv
qPrbP0Pgx7/7AcENaUHGsqCOz48fkD1J6pb8Z2cw1AeBGgGsGMHaEK5M5dZZYWbw
QTbhDZ9Mle4ntL3AK3stz3K/pb04R34VVxb1bSQ1cdBkADaZo6uM5ah7oTbLIL1i
0LUrCVBwP+QAo5iwcrHC6hVW+IkxEqX92JTXiTkEymX/6u2p7GwPOvGTKdMDmuAG
WFOfLsQusq3KudgpJ4Yh7NEq7Agl0EqEIycdm/3E3BMTbdzHz60PxxdvFG1RgnMT
ammZIFJ1WlPHZ3jwBaib/av5lGU63LueR/BjCgXEYaKqQSxDDnd0EeB2xfEO/a3W
v8zK1PwODrf4/PlClLIhLswjpoRhZsETcyZWy5e54r4t5kkka/lOP7hvvzFqiQzR
Y7K0YW1QVp4gDQ08Rx1AIhwXb2fLScOxy50Xf8fJh4gZw83ExgBZ5JXArHI+RhF5
EEuvzVbgwo98Gg/U7aJK51yfJrbKVYUle9BNbk4R3aXWE4cc1NXP8TFw1QVJXOgA
wJP440WeROUzqkGyY/8nm3PPCyJ6BrGfriFcXg6/WDH2EStgeqtbifNJEXgQzozt
7ecDN8/ZojcaLkrieuerH1R14ExPBf1vS+RUPwbVEs4bBRTEm0uV4/qwOiz2ee9h
mGSNZn+VTxzP2SeyMVrDJh2BuZCdk+PxZrz2J1QJoUxFN8lNpLxoHXUCae0LqGGM
vUIy85x7p5zMIkzCS5pyDetllOSOkm9T9EhsPV23xsPO4TdW9/Gk8GpcF6FrQyeF
eNlSwArmDk7sWkzCC1cuYIzwDg36E6bl4nxN8/uK65FY7Mk0HlekiCSQ+sd76ImG
M0cHG2hWRHpwKft5KoA0+CRY6WINw1IfflXqLuy4A1VXY3IIxqgMAbGBLBDE0WUD
21Hw4QDZLW7XqEopOeEzkvOakbJT7pLd7+vOQPkPoDjx9Z1aVDiXhD2F7gdGcYQX
MoTxVADZumKFqWOoGMyyp75jFtkAuE5Sn4mJoMJGjXRLiYAjqvaw9wJXgqX0d92q
5ZI08Zzp3SA7R6T1Z/sqX6BUs2TRZTL9uetX4Sb7f/YYlXpC1PF/daUUnT5ALrpd
5dwjIA6RFZfqpFaXgDFU+SwwuDN+79GQExodpsJC4U1E+b51yrVqgkt7g7qgtepw
axJ9zQ5IQTBm7uOstXQ80rBaOj3UbZcdsa9VZzLh5WPypwzZt3kP3Wh6jci4cVfU
y6FEyblWQCfLiJNLKdmxqDGQhgddmbwJ4iJBZ5Az/myIf1N/sOk7oWyiIf7fUdLr
TG9gziTZAgDoLS4mtY595S6Uihhr4LEWie09318jUcHOPl5/yreKGQ19YglZSf0+
zZNOfUhhN3xY3Gfmq3bfOFCVXR+Ed9wq1HXyRVsmg1bER4PEjBBY3fQe5nyLywpT
NSoewTsKLHF21z0Pe61b8OHoeWbiKCdyyZYKaMxmeLXlP0JFlUunW0HPIOMOKH7a
7HQA9e8hztvi2jnYbJuJkrmp+c2jzd4s1dIWjE5U3wvuP+4y3J/0y9qROpG6ax86
fZ8xQV9ORdxz5cXPR18rXpfM/37yBZFazNnmII2o/z2fxJx8TT3qFqoJTwu2TXqc
TYe0wfMLRGsNLQu4y9vUKhPY5xf8dvk0PVtN/VL7oNxeJyzBZ9HsoWG00DF91bub
jDaTYoYnhYdkpXtisghmnYOEKwCWSVH6k12YAQI4HGVa6xpb2Z9s+x9OdUPseGv9
4OE2dkb5Q2XcDzRaM7PecHEBM4uKSkKffsNJojoFcwgDFzoIeVSUL5x9nHz5PzbB
eYucCesmPqTB3goo91TWdpwUjwUzs7cWlT/Pax+NLnFmM4CEOcR78iHgHnmAqNLL
nmVTR72+a/ScXbRn9asXtEwK25J3abpOarNPXYdecQxE48+oAwXw15bV1PsQ4rP8
Z71oXZQnQszg6DXVYjzsFPIoJQsWzge413YYb3uluZ1Iqvrcd9e+gi2WDE1OkXhn
6ha5t7k+meL4zmWZamGV0L80gtVP9Qt4CyvGt+dUQD+2MI5lvxupxLYHZ9EZzAbi
JxHUm+5v/edeORWIn+QgtUTr23msuVuaZHDSFwrpWmu1bdhJlaxVJ5mrMT2qVoPs
J+aO1ppCwohXuAEdi3xHKbaPT6r21LMPdR0TI8aYHVAV4K8pdvmlg9P3yFo5UmPR
PA3ICUjJt6Wao9tlUPDym6McmX/RO+85VcuE5/OEmOCF8rOQP08MIsYrf2mVkUxJ
XP/3PwfnYkc5J28mVJgK3deMyC/XbHoWgoLfGX4ExUUM0xVmRBqIoHb44QoX3QcC
aiMe2ZxN0ocQ3OnCs2xjKw9z8IzfAxSC8o3IbzI5RJmnAyeoV33RhkAf4YeAYzxa
mMIF+37VTb1rvOUsiR7WsIsRbcQEIndB20ezXKl0CSFibYkO8nBfd8CLV9jYB2P9
nkIgezLdamo1i9PA1ipA8mGprVfORqNoeH07znIqnq4/+Lo6uEeEmLOzfalZ04Dt
rFwAQlEI42vdBolDGtwhWEM4V4T4fm1cM2KxXAfzAEUcTAuJwocxGBOdFV2yUp5r
0/N/BifXuceWzxdHeHFtI9zIOxio0kuaWRhda8SvVHK1uNzd5Fh6AZWQLdIERnfS
7gwBCZLIwaREdPRA73VcEMuc3ExIMC41FjRQ91/bDCd+dmx71WNSmlcWc1SYm40I
1ap5yyHDFD8ZFJCWwi4g6rHP8QsrvWFEXi6WSqFyKDG4RVEiOsTPeBEJ5eqovIoC
eePRP0RlTFlrjIg9qm0ClGa2ef6e+/SgcEx0oQefHJFTjHB5z0L2Dr5gMTRSiX7S
w3latJ9PTGpCQj9sUOclLPtH1QqyV7SBk+pK9Eap2Uu6aFKYJRCVn1lqiPudDhlB
SpgwOGTk9ApiaWgvgFMZtvhPX55yqRQCNx3PTN/y1yHH6KKw2UUU9v2vEfYaVH2D
mB7wR3coul98+W455Ounl+XI+aw7DTDVNBHeSTviEpuRXjtfwT5cNh7NOhT1iC5R
1cEuSSgtYM+d1iBfbBuMinCG16uDrcvHXMiH8zaChzkwGYmpMdIgw7cE4+tqX6L8
bDAjX3FYX+WY+RQi0Ic1eXK+N7Hbu1JeI+vam/zJ9RXqBedm6QFqlkc5UzPBn/c6
DPwt1+Gu04gncB+nHQisvFHFOkzWSrT8JCNPuS6vOWxVtC8o1wcLwwe7buG2itxG
S2O0enHlD1a/DUx+We3PHQ6JmBv5SgdZkUR/mox/jPRiqlIfcQL5l4WiD9Ci5/ok
1854cXWJowWPlDozELsIBQFnNLbKSP5zoc3GGelxo2QhdgP9brXQ/o15+Vu/M7Nt
zdAXd3aGRYNf9jgr9Nvl5SM7ka7LX6zg1zrG6Ch+RUe7FIOjjxpRUMPMujQmqWdl
Kd7EcYWU7qm4hYD+0lr/F32SpeRwIHttHkBAqSEAlFqEu1T2VE4SEn57PzllWl8Q
bFmFxVVMNNwcSWFrpIZ3ovu51dSGyBendP5V7Tw8aAIpYYPNPyhkX0Q12xG74G2p
Cz6hp/J5TKbMvdllirw5epAEQhf9bIXgRIn5+JNqbCOvKIJv1RwdPoYEJFLliW1o
brJhRcWrzOSpqJ+9/K+PPPfFdycpiLw4ywQkw4UeM3b9i5LbTT12wdKBQCzRc3sd
yK0oDG53zayXIlTkafgXMf7XbVFjg4lVfkzJ8lxkQqZ4hABU5wNPXfGGCZLC7Eal
oOAfWA3Uh+N3X7jQn8XToFUk99zbLLQKIF1n8d5Vq0QrwkdAV00w9ap0iq33TB4P
i/Ul0eMuwjwLyY8d+LvAhwEXFZYnmRlx9MrcaqZCpOg1Oji8t/xJ796bIH4K1AaT
NZmS7LKwqtY+Bn9GAe0rPhTXkjVvzehLbHKiVJpgrsJ+raE2P+3h9An1KWtgJpfy
tCVOgFdF+Ptf4u+twjFE0qiKBBN6KJBrCjecgtU+xKUxWZrDaQvxtgpF8QLvZ7F5
D0V078U58QNnuPS2I5AOLDdDRQA0Ln9Be3oc97vGjjMCHuDjxalQdVIlxUGVVRN7
RWYNLG+VmU2oIwb8vqRaLF2cS40su6pXNObv7xLuLqzuBRF6gcOh0ObjL5Or/CGR
DduJXrV7cPWJFM8zIO5YqOt9ftvW48h+2iXGzERb/hrl8spTbUnOV5nayvobVhmb
73K02rPUfuxoEJjibNIHTGwLnlMcx7kvfREBqjzpjaYz7g9J4ju/SlXr+l2oLpgR
D9Ilc+jEuo5qhB9lbe7bXlPX6CVwnsj7s46jSITzrs+UhuXfX6pQbobH8y9TqUcJ
GrC1XFBXOcUdxgtbPIW4ZoujFJDXns3PN+MQ8Qe0CZVc0PV94VulA0x3Gl4YKy1K
G15QyiaNstwjkaYM/qohQMAwn0kQHgO4Gif0h4rdr6m/dbwwIaDazAkWZLnvl/R/
5lw2AD+zm58LbIvzc7qQ0tTgiuJtw/H+oTyfi88SNfHPCMl06KjzsmpAnpwNUXV3
pyeCHJG1XkhDoau/cpuMzF/Q6zWZy5jMXrfQyfY/DWqxgNjorU/kB7tzQ4oMN7gG
wizlXQN+Y/yrSwkhG5X6UKqrODkdOz7bOLB0Kst7Lc1eSV8FwvI9qffDXcvq2Ykt
nfglDkkh7WYRYuuiE35PG0Y2Fv+SGaMlt8Tx7+vPPs1j8JYmyJK4f+5ew50TKFMy
iWneMf0HLGPCXJhBvETX0/xfZg/5vbzM5C7SS/seYAg5FS+cS0nbB8BG0EgNhmud
u9ALW22VMlGGu8feQgn1meXu3A+MvJK1F3i11Dan+hBgpEWVcDnlFw0WY2i9JKbE
dSaC+R8lwApvGBfRlBrbP+VELvvoy+UCIJcP/YeI1NCzVmkwDpg2RUNwUG6j+/qO
JDKFQQHbPhG5J6oAuvIHLvckfyIiJ0bWO49XBvoKe31nd0+sJ/9ur3GaFAkIlky/
0x7dloRUSSbIJuUQbp080LNAmsdPKTfxE0U6kK6OXGQ1DRdgW+UCVCk0QNuxOYLg
d/dJQf+npJkRFHjMYn95U170+NEUAP5gdXURHUgOroNhZM0wHQPVDBWd2WoSkn/m
rLqTprFW3utelPo7tiBMLXQwOnF0mT+T/Fie1Y7He587yt4jtBYWtdw0EYYJO9tM
ccdAzXVGVMYtM0W7ZDeiW2N1GcUfj/L17o5PXvDL0D1ExRnGt5c6Jo4Ntg41S3rB
/IPrr0qtoNDmxXYO0c2HQZ8nFFgvB7C3arQiJ2YXs//zs2w8DKDx1z7D/u2/lY0W
aCTS51oB1XCyNWhFy1jj/8B2UA3+HQYSNqlIcaQZd8wKML61k1vW9BHXt6xEILXn
FYDRKKRGAtHKtZtiUd/57Y2SWpumhTgRvmqykOIUn+KIA0rMnlw4VROMtUQ5/C3a
ehOsdweRxFx8CRGwnV1Z43h1+IW1U+8K3+itvZ9qvSP3dv0NypMmRuExO3oZqzxy
6qXZo+gSKykk+LY2jPr23cnEURfO9MrxUCL9kj8ZbjmvDPh9tU4d4hLSm5PZEnP2
9/EBkbjURhJpAw4JChGpQkh7zY7JFYN8P2bnDBGKeroBNwhKyYji1WvPenB4irgd
Lsyigny/V0U51JOOkv9W2CA7WTRO0YpAsXtmwjU3FDpnDmiza6ZBLceWCblWMcux
JuKPyjCPaKNuE/UjXlx4x4bjeTjuiy5LToh1+ZX9iI22QG1FwnstQik5J+jpgfhb
j15vvALsbOs+G+yFrxWk/AKXz16fLUQeJdjbg6PxsY0dAoG+unENuCb1dF/Si5kF
BXGrF1srU77cPMTmTQvG9hC3Lfxh5D2MkNKpncb4YlfuFHqVrckny9grKwmr3wED
arGXAr+2CgBD8cPMXBKHqETIwh+m+lnuG7VzKr9OQ2ohwXx5iw7Wx/2jISqob8HR
2vtANNLc+pMIb/oF//koQDHCu5lSdEgqMBlxcALLE91j1t6CeXpT40PsywimyjwS
fs2DtqXsPjniCTX6KKj77uOE7K3nS4cjNB1yLpYnLUR0cCfozznsHNfRXEwWM0Zl
9fAqqdqU6pY4COB4ycx0qjewKrtt9gucAxLSaVxRbw2TgEj514DkpsiN0qVgoqI1
hiIMw3W8kdVdqmzxi4oJwXcHlVmZWDecgiUpfTPXiuezpLvBk54j3DYMFLwzAHmI
gX88h1oGcbfkRuEnzQ54n2WzW5e/sAnC+QyuaA7UgVu7enNUm2PXf4CT3A+YgByE
EtKDgrZas18iaikkaJfXlk2Ll6vDm/th0oG7bJr9ew6uqSxEiVFW6Jel5hJ3Ry5M
GbE0z6MWFc3VN/6NG+bQCx3WPqqdOfxXNnqQ7+nPt/bUvdwuPqgRjUoKVv3P4umd
NnEjd9R0HZEK8Th+++Viv8pCEgVnDG6FEGsMivnwwP9+XVv+SyORmS7OM6xg0nz+
w6S1UVfO+T682Z12PkrbAlGLSD4hT+pskyWcf2uSaeN6JlEhX0nmYBT1+moAYzo0
xWl93e/EaX3zXwnICeMUvYoBacu2svxElzTNhqzpmSGQ/hl1WOxK2BQoawwc4d++
6kEy/7CcPgdB2FNKFK2iEInOkRExjHAS0pKQnV+3aOgiM7QlGk3XCrUoOO/2npQW
5ZoMV2+jIDeAFlV9aMeOEdXi1CUmtjRK6fwBacCMid8obV16uHf5TfLABuHIJWzX
u+v5CBRzmQg3T69umQe3pBzHbaiPOH1aPDHeQx9xtPSlW04z+AOQ8LtS8mZUhdJT
UQpaoUdkHWPV4UqtJAgma8IV3b+jqx78gZ1v4HSpO1xJxnA2iPY5YP+0beWVOJeE
6RLKkLRrcEHQQDuQP0KNL5QmjLklhbmxRYO/FvKFNK1thtp0b6UabL5JJFyxpjbM
R/GtmXGoYZhNXZaAh4ZL9GH01d5QB6oykyGE2Muy5lSmr4wyNsXnU8wN/iFwd/Wg
JBZaw2eUfaaCYjfscYySMX2fXnogUYsi2QkHKmyMs+k4XUIRkg9MTWBBtHKmrD1W
+ZIkHp2esCrcIudAJMvTtcgtd4y53pRY0hwJUTZApjTGyqyo84SrgGvTzIHv7xAh
UZ2MvRqWWjAqpgZ1As8YOV82AmkWcUKfQ635W7qpghMT2jODuZgdyhZlhkxiPmRo
2bD5X+3R8o+TdobOw1VEwcR7vyPnWGprZT2zqmW7HSsZzuMq3frsRKsiJoXXunq6
4IZhWn6U21ej2gTi2uquMGs8YX14O6ksV1VcWBmhI0pSdn/jLb0Oq5kBLOekvtrA
tUtlGx1oYkO5DCGeLFawjvWPzcqVpAG/FhFmbFYBaRjyCd6RlryAq+VamQ/ZRiuY
AuFT0f+ht/IU7gS2J0KtHdC6WbXpUs7h5elcqdXLlKq+HJ/xT2mhpAvLwahAmQUv
fiuhDP6Frj2h3Zsv/cTnrOOED1yx80WWAs1V9ElFwwpR4HspPP+6CisDlR+IpGa/
nbkrsGmeVeDPllsST8cD3+ImFRrhonypYZr7QBXZLV4Qza3p+d0q1vgTD8Ooxwc+
rWZ11IDFwKx1zYl2fSMF7HnPEpoZrcieHNHyAieNBWxx8rg5laezNtBA9BzVA1Fl
R5+XozQp1/ZV6rSx4zNV3/Bk2If4Pw09LPhMOafdKygARm6xFCW7O7rBYjBt4z7n
TmKlR3drk8V59gIKq8Fn0mySAzWodQoK3Qp/SdtH068xYS5U4ty3edYmF4ACHFLV
G20lwHlQeUaXu2QU5O4mieHkosyLuCZRVccAUXqqG5qCYPZ05+4mpZtytfYJP48O
USDUa7KeCAOcmKnQGJ47RijokKi34NT44MAsqYkdLflY2oLHHuAsu3ret537XgB6
TZXY0rQSzFW+dTmqanx8UqotDS9KZW9JMM/pCfEFzxLntM7Ghx9qGCDBjhvEqSXR
qeOADamUK8Xwi9qUxKgU6GfroU4wohGXq+K/bhPm+4aLrddBV3n0qhvixEzE9pZJ
ohpOlVtMiwLB7FvMLxY1w/pzzO+/wj65AR2G9k5/V3MLlD0w8OmggMjWA8+zyYIu
Lebv6tKI67kHOGpibuQt7ev/8QaGPSFfESd6z9u0F4wE9LJgZ1UEInUMAIPTTeVr
ADKNCE5Cacdl6YFG+yU74Q7haJxOFCLRFa4bJ/9w3ITcG8vH2NvyCXdi34WWMiDZ
Df8q6gUsOnngr7NqMUvpzgYvPSiItbW+y3tDx5DnmLWCEIklx02KMZoWCEj1AvJG
U0lcBuEsX/pgVbcMqN2LmGvSo8T3yRmcv3IthRi/4BoIMwkTAH/scXyi1yZAgllw
FheytErHow471IqiaV6NWCaf68j8ExMW5kH2tdTKfkOvQhD0MxGtWFWrUMaD9l6v
vL9VJOwOc1J5wGc1LeCgCtyUsQ1tY2Ht8Y9KK9Uw8UCq3B0HqgTxyDGsbVSeIP+E
GohBuDO1jbWlyJiEAsKjN7CYnTnzVlynPK5EFYiuF2FXj86zOk8A6NG8CBsTBDcs
QcdnveURu9XHRD/QwgMk5VmnO8qs8qbWviXQIzwy2fnJv5AcRW1Z2XfiX882ktf7
XSzCtLe1oodYuAfoWzOMiTl9PxpdaOUFBEjeozQBgDqVoVqP62RtYdsCEto4AOWm
4TzhnhI/t2w4QuPZFR6klg0o3pUMr/kdrQhUUZgWYgnZAyb1BHqalCge2ei9bcuc
Z6nuuplrA3B+C03Jnn+77A4lwidUBumyyfPPR62DLMGWX25UfptrvUzhFfM1Lkub
oISpY5ULMR6IOaVqUQfjesNlv6JggmTPL/XZWhK0ruxPDEn5tY0lO0USEOl49kKQ
86MgaPpARx3wbiNgFuEP5JECzLcUCO3tW9vXFtqw44fPzlym7M6iMCLB6/UnHbwr
ZhXQHPgo6Gl0BPlyXZXNd7kAOTBalRDUfH/OTonsK4PUuiNjaCf3pdZaOW8gUPEZ
/S9IrBBqjCSJBpoZyDdHoX1iXXUJsuHV2dgJoLj7U/3c29bsjtf/XTvIVnAMqrE/
/XRVrmT87ccOhm0GJiCHNnTfKuwYDJWJeM1uI7MOjLI+MJn4VU54l8DaARavMNhK
QeYQC5CtRQGK1ClEsXYpjKjMon69dZGuEeBW/Z9yBVZ8oqkhr5uHHOWX+WcI9/gF
/b7SU1VSCmRqIo7IXeWTd6SFTvh5iEJoWJI2gl5Wct4d624kVoL6fz5iMwJf1kr0
pHnSiOTxXex10UNc+0GRF1Pd37T9nzLYx3WYFvVlAiuztg9dzbNs2ALizl7sP2Zw
6OJqxT1gaPTTwwnJj5OyFEvMHjyHKPxNcuO5+FYml2ks6/AEQw0I2BChvDSbwW1I
PNXYcnvRHYOh1k2WlxtuxVQCO0VmVOZcZLX+V6A51KsULEXATPU9PoIMLmd7pon/
YtUnLb2emNna3pbEpoBFzuvfMUUAJeRkgWYq1J/Ej70g9lv2vOV13V9g3mxXtOtk
qCbNIhBjembGDY+eg8KlX0zaqul++6NdupsMqjuvki+ybr+sllE0saZznW9/UIMv
IQ85Hz1oLnlweGOSoNuIIdKVulaFX30dkOcj9MFC0A2xwb9EDqNk/qIbu99LhpIL
uWnj6jMJQj63PE4Cc/CnQ5//k5tWF7QkwT4Ax7vU4ibvQqgJnGFFFUZt4lJzpEZi
fgztke7akPHrjzu46zRUulqayaynYb/9s972Goz+n1YoFvjoBPdzlb8kYP4ucRw7
gQf6/85uEjQqBK4gX77ATZjCDprYedYpk9wGXhnwuVrl2QuhxYxi3FtGDzFivsVS
6IqHJAAYEGaUv7xKucsmWObNMX1oZedHpU70ioszNAfY3DHTXP2ocTpuU46zzVm0
qMrIZyeDHmYT5v36qQ7S4Zj8PK59nLFZ4MJGoPlhqL1Qz+m5X9xUl7tayiF8mu7e
9QIp5oLATNAdjgUzcpbt9etuOk5Fkm7eVl4BBCMTS02nV+lwvvE+SHBuZLDL8BFp
UMeQXd+iOWnnOJvUUFHMBPEBHAeG6rpLg5jE8IoPygSYG/QN7WlInDHMABP0hsgB
VloGDWs1zUyVdBELZer5NnrvoowceBxLbFmrg2ton1hIRu8TgAm96gJ3O0Rhnn6/
063Yu4p3DGo9LuVGzVqDUkmlTuWjx7ojJuBVjgGUQJj98/w3fLTcbidm+Gq/VeUH
CUxPMIKPFSBDz6zN8RRV/B0TseVB2LUYW/0DHT5pNiCt1tKsZCTyvN6VZDoOkz1X
WNmtk+sroq0dSX7+koS8rsCJKcuKcUCyl0FitUImQbL+38qVZ7humJaSYtwCLVs3
XZev+uB/A45UyMZD9AkrIioRyPQN/fzqhfMEPFJd8ljfweYS6cpzG/CFhhf7AQ0D
kQA0PBJJb/snPaimtpx+yNcQYskVF3Rwc5/OLYPlAVOCkfntZn5HSJYHt8Jj7gMm
Qt3yzPRh+aD9dROd6WbKXV7+I0shhr33aT1AJGVt8/k5nZ/UxbeHdLmuCGfKBi/P
iasZVCCYovkOorEViPLH96CrnjJB8zwccGlbxUZzNfnvll3/uOA4YCPjDw+GmIHM
nU6J8qbtYMygPpnRanB7By0mZadlKAx+mKyIZ+TQokQ0ZRLkgxCkvjZvJfKAzULZ
HQ9XVikJHHaRgWKRuYCdirPUNXGKtRyIQBRbjDUBvGIV9EbEwshOUlMzxYidESUb
7XfHFQBxQKyBSE0mD3HcK0gVcIm/zt22IM0iCkKIerdYBV55WALpA5/3vDvamuc8
1aBCfvG2cmHZ+hZbaZeaFIwLWO9FLafF3rO4CVwu0BtBauUzN7Ypn+go6+kQpsJf
VNpUWen2PkDgDVLnQmFVel4YP7H7i1RjbP+S8r31/K5h7ZZgNC+ngp8woqMGzO9y
0NXCVOdkykvHwKJvdhWNrwA1lFZerpW78FeO/6R810+4PqReSO6Q63cV6cHbA5Hb
ix983p26K/njC32JzWcVb7tQ9nfMoJP3chWj3nv3R4Dvb81bDlNafYjut1OqMaa+
Pkhb8F/VEGSVbLbBLNzPaigRXtp6ulxhceWXs6SOAbSsuQDfX8OYqC4p/yzuHxDp
hi0uZPXxJGKvu4XyY1ANzjr3YWy6FpAxwTMu3eolC7CTwsidZvUKLuH73gwR/O/T
lFZGPMozBxxG1It+chXYDUuSxdVb3CVnk3cifGbBR+aNbC0jgfkuNiNm1YJOJI7m
e97Nqe9N2fR8RZAaEgl3X1a9dpy7OKA9PRxftgzSeIPyaNTFLPQgItb9C4XF4SUG
GgKFAucxkPR10ER5GZi/zm8MiqrfjsMihLuChNSCtEwZHr7w02i+nxoGay2MXgnD
oVcnUWVVwy7zUrhwuvhcNZ8mVoOnzI6vanCs8o0fHNgzkQ7IOvzCQUyvRZeZfDhc
Otz1s/LyTGEX7847xNc3u+TSs+afmLgru0CiRIaVo+/bbaWAScLgUtrZcB9Hff6Q
lJ4YYoHeDypr2PpN4GGZ9FCCU0gdJYwFdLRw/Uq+GJL9X9a/sztBr74ZScqqDDCw
XGC4f+jsnSHK5MEDFqYvVdcIeGyM+CmKfQPvnpv1oc285P1lKV3SnwAOaW5Df8Or
UqnJOQnV5yHCv2QWlolKr2KRQxmalXzkV2ytwlM1gGtT//KsMO9jeEO1Vk2kEiTQ
gk/dF8pM9y2/1M5lnHw+nTlxZjHljMlh75j36iJqAwNoWtCWHBcB93Q9J7ea5dSE
5sn7VKXyDVS70mUl+nxTlqLYOtob06poGp23sPhOXatlb2RfvFOA1X35Ze401USP
fxFKfrs3KT9oI5Y3gK6IoYF/DR8Jry+wlTo4ByIYmxEaKKs2Bt436/eOMgjqkEJS
vJRV5IUcWvMi/S/tOZGrxhvNM/o8sMYuhLWHje7aSfcWvA3L8I8YO7eQ4upABhf7
zF9m2OamkFsHOGbO8icOVazTWQiKQuZT9Rd9p2J+9/Vbyu5J8aHjiSmZL2idWlKl
8lFSRbzSHlsV8ge4CdsiLM4mx7FqHM9PdDKGVNw1Y34ndPuYHlv5NM5vKx0NUIv2
CCLgb+hfhJMIleMBaS59sX5OhYneathw3o48dMhTQ+KOf9jsuOfqsHkdMSkSQFYY
i4gBwwk3xil58rH7K6wvb8N4vZ2ALi/lCjUV97tazR1y+m9MHAiV92Tyxreq4djL
wHgHLlxP5pT2mSy/ajpCZfm9HoQkO8wDyfaDrnAOaXdqC27/lhRDg5BzzPLOLSKA
95OJZBoA37hoSQPjvu1DB26kXI69FJCHFBTmLBdJWDZOl19yHPa64I7uU0o6G4Vk
L9QUC4hYVKiDQa/4//PcLcn8Oclcba+XeB5+3a3HOu45oSaMDxf/T4J0DCrz0ifZ
CDlEmT/qoBm6Y74azLcxWu5IvbWBgY2PuFrp37E/FTDJBAnuPY2ZKKEKtWj6oBPu
/bs5svp4XsTUEhYDaKjRGIATHrZ+tTPHmM5RTYQOG6GQpX3l7+A3Iq8TvIGnRo5P
e2xcrdnkUqcM6hyCrpxxxtwcgCf8q19ITMTAprQIEefxh8VTvfTHiP/MivbhPY74
UQWw7aCFeWnlR5tLo5laucr0gAoJkbZ9skMK9Pao/Jnx6FUOH7qhPjxsnJIV1rMk
5odA+dvKoU2ngH8oDy0dHg/1zADApCO73Y1qpvKP9w6ZIfCpz8Kwkszpgf36KUgO
VKvq4b9Mra+g77y4Zxcg9kM8KjKS1YzIhTYJau6AZgZdClSIusATxnOSEgwrqvqm
g91bEb3uRV2cLpXrNa0x13UHuKgC/AoMdi4Bc5OIO/bEHVt8Bm6Nc/kY9L322YeW
LRo3DHtVcCEmRg2KMVBIl2npmKjNlpqLWv4T3xLGKL9jBixvX69LSq8Fb9xfnGWy
EmvCP+6blyxKyNSTSED8Jq+uong09gTu8TcUnMIJDCbtCaQZdqW1xkFZxbjork89
KHODR/cw44NBJemN/zMLuPixqp2eouyvogZBeFvFqNLn0uq7/264O9uDX6Ehm5HH
KN9SFWQePn5efAqT8XTQN6s5va4BW+VUEfWykCs2903jMk1k+RC9gKOuwlBTJEP5
ZYkLY0rpCgWrBDjvv7D3gStbwUwzoSVCa4SoR0Jd68G0JFJGI5K01Rn3BwO3HyZN
aersZMbV+CdbLmh0WIHEjsVpe+hHnvwmfIOz2+MpUu68BjPJnL852cRZGzrZ5fAq
+7YrEWeyfl1kVgjj9mwRhWOeOUMtCAFYSboRB7oCaVIrhfrwmTxwSGC1YC99yxLa
ugm7JYXOvucNzBlztXBvD37SleyAj88Pn+uSIsV3Gpaomn/8G8kfcCGh4f+v1jL6
e9hTTSMe8cB41Nz6cNSQ4O1yFTB+ePgzE9GPSgapQuzY2PceaKReiFJMIEBGG07g
qJGpl59b/jft1ceRLjk06/UEPCYNn1Xs2zLW1+TYzycWKKY8hEojHQmiz8o12xcw
JssjIsKtHuC2Xvk9GKtFex32mlxKMIM0z6wAF5YDh2bkx7B0bIjG9wymrjpyg9Du
tt77agGowR92PQXiUBpRRAmqdU4MzwAP3z025PQJvyvOP9epo7sh7Ln3fIlmCOjd
vWdOrpHP9wk+JiR5gsNIUEVhmw4JUKWC03/VQOOOpft/wrmq665oiVoyj5BpEkIo
tNPbPmh/luuQZe62CvuWsEeD7lU9sWlFFFoFBkbirE5RFIETzAfSyCm/vOziVGtV
IUQ5IBvFRcvs+Me4oRg/S5QDnxZbYgDAKkNv2yQzwC98Ze/HfrQB/6tFM0GCNseS
JbIja2wgubVjVGbR2/kwhY4ioXptUy3iPtYqL7KIXfQ38ffnfg3K4GvIP3/UuHO6
kXCwSj9x6Huwa9Gl3TnX2rCLBbqVD53TNwXZvkh+WAUbPfoyMq4tadPxenU9vvwK
gvZds/EN5olUPv7Gsoe2ObbOE/kBphwIxw+hrAZpiS4ERNrG/Y7LrEswJ0IxcdF0
YiuQyc1CxsXLdsalvsEzZg7fAOj/jNdRDPnqX5bWeb1eSkzz/oDNNWc/x9WnmVGz
/ZYgxsdWxsRbLaB+q5DB5feo8HIt4LVXMEPARsK8UZkmP4RboYJQWvmM4FCkSA6+
nX7YqLdde+VOXbijD9TAtDMW+zuWFDp5EojtbqLNj0g0WyStEkUzPkH2yQ8qfAgb
eYX2Be4foSlxloXD/xoIt8F0/3OEhTvAnwZUvxjTVynCd63qUgXsU5sXR3b8UojA
OTM/HOCXc5GfaBwtdfjGyOb8xHOVkg738jkEYLlzFAHJ9F3SiKqZxsKrkl67fZ4U
fm8aNJP6oNsne1jHWZBIl5GbDaPIZB2cDFm+llel5z2Sf6iLqf2gqnrOhzQjvDSY
AFCanwtzpR2ai5JS3cbPSbxi/ONYybD8qzXEYyQISQMnSVYNz94211MVVfu3+lw3
VM4g+Phl5L9B7Hnx/GsMTU9Np9yHoG+vkGdqY8nB7KSD0v58Ws/udyR5VGHJgank
8NZ8sSHyYGKu440YpesDjZ4wJefaTDEB7yl7hVWQtJ7E6oVXNcQO1mRM7j1Qq9Ic
OFoWT0iek3rM95Kq/QfBV/bkamfkEEp0uq6nCUqI/WoJenBfNdvPGxB2p7V4iTBh
U4HrffrN304x3S2VFMCtRSxiyBxbDQrKrQP9EySLlSXc5YwivHx6T8wvrEf/wwIQ
b3eXJe2TC6/OU9ufnnt7IUqSdIi8kpacOfL9Ro6SY1wooWpzP40zmVpwSEM9WXFu
Fz/WI35sEPzKCYU1Cyu7v1b5x+joLOIh63lZOiIML3HzRvXgbOhEGo83CoC8H7t3
l3o6Pblcs1LMeKJObBYEbX0U0F9WuiPAgjpeedhU8lYoUE36cemwYAGIkJqExxbS
q+22IN3SAKgM5flZ/N1E1JX8AHw3pi9qTlUAceKSdfeFpwiT626hDuzsd+p6v1FS
qgQVm9Gwgnmr5M+7dYyiPAz1Rthh4t9oUVIVu74EiLUABjatbxLfaWH3uy8CGTeK
mE6alRpbGOMhdrBLRtKGRsz9cICl+aVBBClwxu6/tEz3tpDU/0S+RO6OLfGBdaxv
W2N2lBUhAWzofqui6kL4ZvVMIrApNUqNargKOVI/+GEcbstkSTIhXif/9W6GkFAE
PSu8SCjhOyTBiwg2+Nro31aLAuB27QeJ/Y0nB8rQR6JxH8DLvg91KFkZOS+bZdc1
I4qM9iP1TQliWPv6yxbSJpDCdBnP5Q7qNyAWIN2zD+6ntQW1Fu30AMPaU7R24Hs0
SVp8SZbjnmAeTDvS9kL/4f4jzgx/vXnhUzqfcs4ne9ex1Wj0XOL4eBk0lddEkacR
RMgOsxT8qgxni385kzRlve7PIeXYR0/BvjWxfGOedilyQ+YqCXOFLF9if6yvoyRS
4ypPy165ic5eXPzL8SMkY7XMsTeWRutFPeAikYr0RKlv3/m8CbMfpKso6W8MfsI8
tJRfDU8RCW7nPI59DFBxLA8O6a4eKHiph7SXUKeKFZ11Rfoov03tNubaAjIsrsGw
gJi81R/VGHKwXhtlK5wD3Qb+unUVJ3F4tFoW+fgs1O5uKsNVYYZDiaFB9Eo8JW2K
LL5xF6cXqojAa3mMYmarfnaPI9nmb9v4pp2Hh3Wok5Kz40Snx7s2sWGpFglrpFAX
hgexe42983mdzD2TzkoOvJdn5zllgoIEtjFI7mkDtocbvGCvt7RdF+1FKxjgmnNd
sliVDRFeRh3O7zastdVJ7p+d1gkUd8as5Ro4PJA+KvwRYuKpmb1fM1Pd9wd1PleY
l0nuP9l2PZc/9NfKyM9CiTM6qK7ulJM7nclhjz7gqmcrM8T+6gg/LGTEO37AhVSY
WL3a9FcMZGnK9ErLsEDWC5DR4Rt/eDr2tSxJRQp0GvUsHK1ye9Z+LQofRrM8EuWM
iJMWHQsQvAlh8MzCbTIV1OeEpilFX4jK4kHOFT2vSy5tBFVlyGVDyHrVLttkTju8
xyMcT2d2rkOR/lexSF1uGKBuKwoGqCH8RTtd2Sr6s0+49Y9bsPgwlA2GF3002BWH
kUtZNXMLkuqmJMSL1q/ORHIYX/o8JA8+0ojzerboyUlfPUUJVcz259um7Ya6Ifck
kyLijuPeu5orRuaADnuRce7GSSBzlMCLEbUGX/+V/AuaynxhheVgd0nAEf4ZYBzr
dCi57yKpL4v6D5pDv3lyueFNpxCeExf345AGDlS/qHOhKp0lm2t87fSvdoRVX2OO
Jx8TlTnWvMTkpVyoUhrJXMDV+vEwRbPpkCTbFTH9dtSEGrxX/KUJ4eX4Gr7VkJWW
mmi5o7VceO4nHlOgmSoKcLhY3jg6jEtWTGhBzCnGMksMnrU9ZZ2OCN1LAooq2EWM
dFm5PqVyzvwfdvHvASFpO672o37aE3AAhGRih4PlqeR0SUAfTbPremfk9nEgWEvm
VJ/3VpXL75jMcdi9mlET5fSZmO7V8lp6HHgQczUpUTFnafstbkY77bXNQcNWedMM
Cbrh9+ofYvgEAJw5m+EGpOvkh2jaWXeMtDlvAZye6Dzm17+rGqZgBeKEH9a5LW/1
FHTu2fio7slGN1ZIkKRYcEWf64PBCtVKljU/4EzbMhw71cHazgK8zNviDTZa5t8g
WMUJwQdt9kowjfw8OQYI5hci3ynvxARGLqlAWW+a5MspfTVsbTYT4fID04ycZVdL
U/6xua9Ibrauq0dq57Xj8jDrFtqIFdzzoD60yNhIp0WeWM9SqZcLTl2McB+Z+XE9
D+IHTVAuIOJ7cl02xlcDgIAQ3LNwCzM6XwYUicLwcg9BoSatPjH/2h9tCTSeN81J
e3uliEVIntHzGRmgL7UZYudXrkF9aggCVbdic3XDR85q4yjxGu3CKvXs1RE7V2Nu
KdjqWaZ1tp3fDJzTUwQaSDHALM418wKcIH/h7wG74GXEgvOTZXi2uTJvW+sb3RfL
Fviqwv+erZnSbvX84qiiaIHlf6DG/NBs6pVHmOe1D3BFl7IAfWlf9muKqWqEfz8r
U+4iOB3XGsnwjv0jTLKnpeinRQAU6SEnHh0qNdcqcCDHG1TLQJ9RJR6NkNlvKlFN
pMzaiHMb3aAbBmWr2TtiyAUDfi7N66o68g9vQQBbzq+N2lD/NrxZbFZ+i4200HVT
A5Ha3jyKSo2viIMwFIQv6iBuy3SwuNZGpGWO3EgZHp4ycCDZ30Xp/i+w/982gY/8
H2+6YnCpozYcsA4Ku8yzG8TbXxnINkMXSv5mxbyUh0kgqItc1YFEWH8gXS1NBSbt
yExKmbiYLMGJ3oimZMrnEel1umyuD5+XROugf2Bf0I+AlXfo5Xv9QoZS4jI9PaLv
STz1w0tDUcpaZufAiAhNXepAkqgIk8m2mlze6++Q7jjLJUhO7jlrGlYoGrI6HP3P
I3qRIxxwKbQDZyFNobQKw+mAUtZBixDVnP5PAouOI5Wy6pfoLdDcHfaDBuu025xi
C+yuLUGuzvm0ZdrkJhFbEiDwNujKnaz6rS2DPF0R0ckjYOTkCAy9S9rNvb9CUxvN
wSlAq7q/qEaTIb5fFuVKcMsJrbRW0EqfL5HSj6noRYT1J1BAg934jnvJg4RHEVNm
eNNmf9vHn+Tevrcj/iSntU2lxx4ztUlEYpMcz5HyOelG/31D4pOpfu1wOeMMza0l
bWjO7VSZjEATktvIcVGWxvMavSDk2XmNuApgVkXzAXUtSBxQdLV3neERPCgsovQP
cHcqSZzB+C0+H36iHMcHaSWLhWjAPo3vyfb/mFzVGXrX1FUPZAsNyNqyVrPGZ9cE
XbBVAmzGoS5qzB29IHHA3EBLqsCDdu9hWUUoKOimHqXwAc1UU50o2QPJ7gdYOaCl
lhzGUFKI+t9OT31eYv1rIoFlZc6HxgCeMCZv0lGN3MbQs2i2QnG+QITjEhXTg3U4
3xXi8gutKapX7nDrxj+kBm4ARCtldRNYkBWcqeMTkDjOsRUL81P1b1ubsId84JPQ
hNu45K2OIeeibgGbiIr+txzEh5kGQBXyHWqWGmgvlorZOUNZCbWk/cuIvf0ZCPzU
4BmJM8IjtxD0UVCCrmTm8Xpfe9czRuxTPkEIDLh/bwUoMEkqhSAiM+a4rKEohht9
iuDIqAo7K+ZhFDN453LyumSSJe/NrDAGDy8spQMNkBC8LI8RxjYmAkNv2oWVB241
2rlLDDANGZmvB2L1dk7W60xJyAw9f3pEhU2dbkFGSR5yAj+ZXOfb8KH7w3zNDXgI
kTzxhDeeWRInZVMRj6HlQIWbpRSHcPr56L/Qt4z27LwGb9BTYwcbZ+NeLBU0C61K
b7NxDb3KqWPgMXacbWsrXW6yirfa9Qp5Z0t8ETZUcE1IRK3ETDrP0Y04eVixJjY8
n/CGI9Gf6u5vYutq8M0MAkoCFifjHhWggNghwnqDS5lkISOF5HVIm2DdDzOvQZPA
20zu8gI2xzMokaAkzrtJTDt6zj4SdTF0UIkA/eXmQG3QsN5VnOal1Yi/LmHeCaAk
a5OvPzEebEBoSqWtPZU7nWyOQr2685riFwXas9iJgAFCI9pRx0kVmQeIZezkp8Vs
uWLDJHVvxDyyBfCHKhBdW81eD72Y3rR+iEV88zgAbXKDpUg8eJxfuz8vnmRCYqlB
wjvt9J6wYfjTQH9KsQPeCSjGhqt7EsIES0QxUdNF2VfvDEN9TOndFxUEgGDRH3UJ
IarO7q09wx6TbDsZyr8fOACD659EFnlejx3wgmBfC0leT+5qkB78Nv8YID7Mzqbz
YdTjsi2zNImWSYTg1lVJke7Itn3m6kRHLM1Ck08qJHFhNy9wUP91IqhgBJVUB5Ok
3x0zJWQCZbBvkXV27i9/B7c44iyVkXn0T9i+HEz4718+g5khzfEYLFdeWSegOEVu
E7L4D80/WQ8qjyt3JaJ7cZddrFvk8hVjNMJXmO7Tc3PP/dh/7nl430icXw06VohG
xFymgpuc5O0zrg0GXE5Mps1GYLzIQt38qjKF1zMh+HeSFqCFis+We+K4Ib3aiZNM
5JdJsL/b2JzUE3a8wxUyQAi5hdEsaoERooGD+v7yqd85YZ5G/dNpvyYvQJFDwufa
PJLolvEBc1LAbMk133SvExcDjfxSICEu7MBmrwk1KIH6mhv0jeJ+R/QonoCAJxCJ
TMsnK78jfNx9QnNuvnM+v/qPaGd/cjApRY8DwffrxVJtwWzF6hELRlsxH5/m+36w
J82spZmf7td9jBSnlus1YdLN3sAkE7k4nNxtd6sS2+uhO4yPOqVTJAEwpn6l2CXS
bUQweAmPgeTagyqxwK1oQ4gnqOw33hzNVLOSSyH7NZxBb6FQxd6PzyWYlYaAsI1/
smKIKP3ILGMEUknK1xcSBKbtX3gqYZSEuKZSwDJn490eL1ja9ghbAffrFjlosy9e
B9Rx+CMzSClLp8ee1heKTcoJOhRzvWH3z1iGH1SA4TFF23zNnBK5M4GR5ixTACTW
arlU97gj7C1YS0U3ahA8hqzgn8VY4cKp3qOv9kgvhA2S/eG5GUYgebavnxL8Si/w
BaPXt9ztaW4ePqFhfdB//pgPzOszrXWRGxQ6aQweZVjUiOdeuhimse7oHB+47JRv
bvTJ7ozQBK/65uofOyWiRSzFud+uOGbMdQJGt2wKAcbQV3tAZLU8AQlXZx+nbD5e
uil+4YAZShDrDNx6/e/IR7lOEqSY2D7fbFvxtud4/++Po3QcR2vK3wqOcBypSHZL
U8IIn/v92JxyweT1MNm4RDtwiOe23pKpr6YpPNZXkxLPvvT+Cq3s1WfhqqO6HWrl
Zvnb1A+H2kKnXARGhPyEDW8AK9n02qscUMw/g+H2/bv9nzse61wd4AwSlBBAZ+M2
7JD72CuYyOZQzuhryd/m2faa/E2s4U8gQp8ylS/hqZim5YgWHgtjJc2GyCaETgVA
coW+53LZ4fNWV7etMO7e1Fy/524eAsBPvXX+I0+GETsaDjoiUtv+g7vYrcqla0Ua
2NOhW8fffkXJ0o6i3wagbOBUyryeY7s1ulBjIGmXvhHQZhmtHiuoPEQHkOeXKIQM
vL/oMdzGH3+hOsH6jylTn2k9muLMh2TT16YUZrg0VB2jKYe0V+AfVJkCmfbHi9VP
UAkMxvl+Pvu7mlfPljit5CzDX1sGS5iMoGqRUhZcSresojeekK2mTVyir5CAZsMZ
hv6oPa+xsGZ2exWglUGyRlOxV+41FbQj8AGeLDzGrn/HKUXSxGHwm5M52CJcGsBN
DZuDT1oz8XAFDAMHatxYQFWb3eWPigXiwj1Yldk5XmZNcoPmmqsXYWEvYaGoMZox
gFKZn+khzVTdcpS0Zg00V4jpD4vxet9JtFBMcFMaMWZCQdz+Bwb4bOlcAnxlO39b
/Vq5J4drPTF+S1bOmIi84LR0VihtheG6jeNK2R8s8PM7HSqmUec5Id7Aq6786oE3
jt4zLIGgi7J44ox3emnclSAmL1EkKofWkF7ASOM/rnkuYjfx4T70HyRcqWMPEM30
yL4Hqm2cNoi+Fc/iZLLz0BcLv8Y6PZtXIP+zc1aZbQZpoBfaIDCouQrZAkUBHOLq
OKowcl/Krm+OoDgzQUhhCR1cINeYp94tjgvoLJjojo3kDTro850zksAyPgbYpCAA
cLWECOCXnFpjLhmIJw7GNg0D5HJUI63mYgW8FEN9TT+Dnm1OimYLkpRPD0BtTNWu
673APzIddhQsFli8m48pkyzggTDW4G1x0UfHXkvEJGVwSaQJDdDAPtJ/JvWemyrJ
sLeYA1cKOuVRcUQbZNFAYT5CGSNPIxBcAaej5qiwpOpSRam8tRTZBknoTjS43VPm
8VPmdz6EOJREuZ8kS1MDn4xWuL6uWANwJTseal+YA0tp/pO9Ba/5IBL3DCEkZRFe
EKKlL540O9UZR6wbAOgHxAXXnWNua6jEWhwnOngwVr/cBOA/xo3fh5JrPriEv6MB
zOyElIluZ9yxQW1rt1HAX/IcJxnFzCvU3T4KzkJoVEwlPNZeA9KaB6QQsiZF6yjX
3tcbw98dmD8cr6fpTCZyC836TqxUyc6OgxKjt/HexlqviMXRitKncI0uLYWBKGH7
GyvTRNhJyw0TZtu7bDVF7OYQ+I1fggRT8xkR5cs8IIrPRF4HV5M2dkXAgPHfWda5
zq5KOhfvJMfUJOPR90puWFdFiWsMdaUWv8MrtGVGPSKrDclbRdzYDkx0yTj16pMF
knibzGQolwX+gYTrFSGJRx68AS/xsMdqIb44h0t02k//deiyM8AZFg1fMBMGal6f
+CaQbw0sdy/NEzXoMpsRniGXSBqpzUBPoxdp99xVDN34eWtKsBFNv3ZpJdKcHR66
zFZ1/YsvR1V0ZuIEzDxBNbVHr2+4OkiCmaos+4uS5VzzqYHmhZNQZ9t/mHbKu6Da
IZFnglvUWu+OigxFga+7ktkW+AIO8OmgAUnsghpXZqe8CvLReiSAUhv8c1AxUGOb
vHRpz2oPIUeG490qIXCw24VsJPW6sTwufvk6HQrBj7zTpB7mo2Kz3D4f7uqIV6On
y12KCNTLWmlZSAaf/39DJarjBquyE3RJJzaoJgVP6lyNDyctEnvdmY260qHAF4Ya
ffynTQI8adC13xGOtnknfG8jV1TW8n7dSZWXbxSwhds1+Z/PGu7jTDMNhP0Um2cR
T7lmajL5pbX0Gag7Md+zG829Juw83swQed6mKeirjSKtUzFCHap6VrLfPbXZ9yhJ
bvQL40ZulrahWVI5xsuyp5obgg88JMG9EDJbWgsfLYV78oIRsiizeA4tcdB2STQ1
S6jD5f+JyBD/R34+DEuR58DvIZBxt6c8HnvlNrvRF5ddqsI+NTgh18fb2D788UUE
T0NxXvd4yQLI+I5pZpMnil5W+4Q6BPiecQd5kER0fXMdXxOeZGHm/Z2tGo6BN/qd
jXbdkcJNXtlkT7tbvwUq/zPSpUcgcYQcsgm8aJOY2NrL350V15m8VGL3nw9fEZJD
/ltgkKPehK+yFl200eCFVB2nGQKortOWcCV37QyWIVRspfHe+EK1pdJQg2hPi6Re
i9V7qA7ai9vMch9gmEr3zk2HQ5jtbinQHMsSOOv+TKGEhgiPQNvQ4SyuWYNRyHSy
+TkVyinDFsfVcq+6Cxk4JB9A8Q+s/ItAXMWM3yr/6YrVj+tPNxsLXW6/61lHKBIZ
kLGlTGKjtAoodjQotAmoa3mw+4fTU6f9rA0qydu9GcQT75Y9hCHCURevwcMGtcAc
hmgxpz0UU7jxPw8ZW7+3H7Edzaj1ycqPtre6TB/KHMKTUkzL33LQ0B61DFo3JUyv
Nt4Sys/Mi7SMZHLntuh+5Q9bTC5YnKaR2IJHs0miXv4Gd10g9LkCNiKoJRdVTg2J
WniLzZG42nxpo0aK2/Tf3gYQt5xHr4Lk398U1k3O2RWHa4UoJmog4L4BEB+XU0TT
de3kVrTBQuyejoJ22NZgnnKYOp0StVi8nlKugWH1q4ea4BoRwJczqr6L/jVbAfOx
fh7reiWEMmI4Zhlcwfyt7kgvvKZ26diMIPA2mh5nICk8v5Hd8GMz1a9v2+ZT80fN
V1j4JLqoXskpEm1+Vp1VHsBxSl8iCC+ZsMNCCH05BI/S1+r+POO2IfdCYeaNV+yP
odgtFHv1zVg9q3zuQJhAyQEjSg9q+hoA9HyUgeevgCej14laZdGe+o7O0MJcakVb
BPg/fdpp3pH6jookN43uKPhs+4R5KvAl4geWlLGw2p0mwdazvJZepsZtvl4fao/g
ToICM6ZybIh8YRl+hs+3LZtMUVq1qvyA7X8qGgYrvVEneBebzi/5NsFeWs05qsCS
WIbvOTExQ5c3KAImadMaQCQfqhe68qt9cwlJU8VKNU57pCbSH51dETpdvvaFY40d
rwKcaVND7rEu/+JwheAbguTWzST9ik4pO5a6zvlhrm07jD3jO7QrD//8vyA7ZQah
FV0ypp2QyMX3xQOPXUKSvYV9ZiC9/lZfjpzOlWoCNS7q4WtAitb358s5QYvn1ZaF
setI1vny7bMPM1nVD5ELL0tornc3NO1BEQy2aqoIKAnTzaxzP1xPSH2qsRDRmpRr
ReXXfjv/TcNiohIgcvyYNk4dPEWewtreJsztyDpeTtk5Ad7iIRiwqiR3SZhp2JWK
ruvTRfVUdE72QcRcrIh2zxXZ6/TIkKWeyuRVHGfCX3mXN8sSUx3ZoqUpxEtpJCb4
GfIF1ZG4vk2Qu3OrA3TTa3IvDfdi6dc1YsdQ0MfzieY3UAMJlmDyk2bf9zuhN1qf
pydtPesJYar4xw5ZT6XKlWCGikni8lsHlEZQ2SoJuw/vVF3gDPCqIaRLbC1CZvEA
AcxXK69C0tUFIhZX60d2ML/yAkpKKLybwdIQaw0nCHQFm5OVd5FPRzKEY/T4nis+
BHLXDIF90UR0gslamZbBaEPF6T+tx3oyuowz3/qtOnVSk51y1oCoi+Y4/8l+NE/z
KTem5ZH2rjfr3JwqQjxczzGmxL61L1TOSHZrn6i8txn/C+ahTNWUwDkAYtDlbrKK
+SXl5KpZu6OjeIWxUaMj2w+Y6TQ1jsr2jB7rehMCK8wWcBFtq0T7GqYc3FFbhyEL
qIicHFnsQxGghk0aTW7xTmWCV7Yc3BiB3lkvdnNq/Y2YkIclaHvzJgwQCZ4JxRt8
edYT0y5JEvuIKD8g6KgavzQfj7gpwaF7feIAlE3T0no3TxEX7Oa2UGtoLtweJ4Wa
3I2WfPuNpBNjQ71I3g2RiUoQLHllBXwminQS5ZzlePXT+CGFWSE35Oy+Uhe4gSQ7
ZjV51Oa50WZhBJz1BWI5T8pN7AhkrbzAmWMf5ZJ4EpIK2kHplVnOXJe6SI/1901c
T10m73auT5ZtDjx/C9d7UQs9xPnx3aA9w7rP7CpK9I12lRyV1e9+h2Rt9e798FIq
A1BFc5ilrR0Nq5ZHfFuwGFlVDZWenUZZpe7pAX/9zWk4uT1ovugUSaVdwiWroQlj
+/lk1jh7h/sCVPm901xc4DrgivnzdJdzIaoWpawJlgX9rQuVA/w1G16j6HAlhAiN
nDjQlB/tlT6/AO0gr/1f6W8p8lz/7pZb7GwJWpBdRR+agN0o6ECRm3dafSXQweAh
O3J3KjmH6dI1teVQtRpHpHlHnH60R5B3ShD4bP3SWVOCF4Kld40jty3+RNxTDW/2
t/fwamwlJmdDDeni4fC7jigdFE9L4878NVh64jfBIu6I6Ryg/lI2xI2vFmpVmqnI
AlC5uEunQVpB9TGKVID2tz6jn16YOMSQ7mbB4sbPzKT51RejG0tQ+QGZC2PEACXK
i8yR+3mMNtOLpHtU1hAF1hkNDpXPe/Rv83y4Fjgrsz2CvJIKB6FE1X6hwtA7VPSV
T7RQiMDr/HuAQPy1I/qJAO7RhjmA704mAzjgMaZy8tPkdBsulN7XoRZtVYYR6zYS
EcJfKSajlNGZ7VHKKcRlHxvKOKmS5+4WbfEQSldADoYxJ9GLgOnrBLJ+Ly8UECx5
aVxdn08RuiKpzvBdTwwE2ytyVuJJ7S7yn9sDnKNRvTZ1VCSrmk3cul7ASnaM/qia
F8rQLpL3w384f84F9J8kSpSYG+i7iOG5IEZTJqzaQsKOcuA3S32HUC2jEYfj4Dbc
If7/bKW4HCIWeyTOIGRZNM0CFo+s8bUZJ3rKvLU2oOgJmfT+h/oDFS0x3w5v9bJ5
pLEeHAzclb9vKB3iZxUXJLd37KWsckk/mKVzpJuvJ0BSeoY+BQFIwWj72uSY+3cc
3zPLEc4u3GF2+c/LsYxDPQe1Nq6FzWUhD+6kh0JNN7bCoPgT8hRCa8mphg0e1mJb
901VpKChBpoC+IsKSeREp9ElBkXvrB5+mruMonLvmUyn8nbvise6p6atR8ewGI9i
UJn5dVai7MftZ+YW+wHVpUgNfGtD9WEEhFmfIGkJMmhCIHiFqVLxoRO2epGLGSIN
SQSlmymSHWXNpOp/FNXzwyx9v25k6YUR80d/PHplgQtKwFkHf27RbSOJLq+51DOf
EY6RxadBVIJkFXK1/0IvEJXSaA2Vp6TxgOdJte2yjRmokBeydyqY9qBUkJwY1MRy
eJuxiVkO3a4qUxPq1P2AtEUstly/M04OTq4XhqXbcAyjzjS1oNE2SQXwA/NtGRrW
dUI1GRjyyy8dUL2Z6XJkw2lB8LQWRPhY8J6PQTulYE9yIgPGlJZaRVrc4vCLJuaY
Hdexph/5e2c7ZA3OzY+KNPCQcsH7kdGc1FLJ7H6VZmUcZRGwqEEv9EjQ2UaSWXO7
i13CmJpLenYydg/rsv6RjbMA6hLjw+2HCropObfzv40JMXcRgbCUpp219Bs2koBf
4PZKGXN/8MOOe18yOOE8wlUnXODwqVLOlZmSJe1JYULpYcSqVBTb7TGt0WPvtqlf
x2wZqPT29jF4faJOx3FFMKM4PYyWXH8/PkcxnZ7OVSwh1Tho0SxElVwWGJgbSL4U
8Fa5hRcnM3mA0sS3oeNUMZ/ib2aWh4tObaZT2YALb+acFOAzftmYf9MExKU2r8+8
IaGwm7aqyvI1TcTIBAO0J/yx/ZUcLFvAHKrt6TpPC3vlLGYNgm2ssOLqVVpkJi22
IRm5y9kYpvHhgeukBhhM+65EVxWMo94pBiX0Y3l4VfffZ1iFcHp9opzlrLH58E3X
ChtDNQ+h30jeGQq+XPihvT7obWOdjVsIHNccif9S31KPRWGUwKjDzeFzs8R7oMDo
RtkxOJksAKyLUp8NZlAnIHxF7+Qpe0MQD5miWrvfUAPK6Vx/+T80ngw6gk3fKNNv
73rjAv4S6EaYu2EdrLiXHKTV6f4V76ocf6Tnd3jw5vwYDHXr64cuwdZ0PZI4kI0l
3XBoH4b4xa16Ab1UWyELWeq9+4C0xFUAgBe7LeItY2VF0H7kYzcxnYcSJgLU/lF8
lMC43XOAgaljxEZYYz+28jQsxV+xv4toBppSjmvcn/4wZMhm6LaTuKmR3STH/9z6
ibosilWabiyI96DM/XgipH0uXYsVZcGtXQiu90xbtRGYNAyfUoUwTfrX1DfAqi+W
QuazFT412hTgeHmN8LRP4L7KxScLmWB0IPSt2MFPIHilg/Xr4DCrH6K8NtISPuZV
1Cz8S83Fy+L18W09k9THhVdpY9lXplZB76/LRrN3tU0yy++iOR3s1hksghGI4dyG
Cp5LUDn3ftnnYbqYxXTCHOj66axKS7sxa1cn5WTJUB2lrYaxU+Qj28lpNODr1VZ5
rqOEefU07JdFuwenFexV4zC9wT8VtAysD8vWWbvIqrQVmLAgTU6XEN+4NonBpQNn
Qnly4Q/3IwnOoWv89JHQpJCfaE0yTc7WCqnB9mUsStuN96OsmogVmq8cnrENp0ly
FFVbf1/ebxMLU+qRbrVR3Ea00FuK83xIKuzTro8iC8ueugASJPyPrhj38qI8CWRn
4uYchfCGX4Qj+rAj8JbWKcVDLqF7MQWa3+9lJrKz3JptD7NdLz2BhER+8rIY1/oN
8AeFU2uIbVY2vkJnkl7zJDyG7uhuGCf1FfAINOtMS39FcuUqop7OfsrRsjNeSU7w
jNbNQLx9bWJ7pnRBiDEXbz1lPFfcP7m+uU/njLopvUxuSqO4qi2dNrRLj7i6tJaN
2lDOWOJiRmfQd3BpkVG7BCfRDo7okC7titPao9jCDvmydYM7VlG2WlVoBJyAqRj9
AcC4qL9PR4jQsK3a5Rwt0oOVeqicMpN/zryMwy1pNeUYf3P5UIFK5MXrJ/wYH/5x
yk1Ljn/XWYDWPOOBYWWgwo7vfPCfjG1IyJTVhIVF/TlcFW3V3cuArdO5AKHEP9te
i2RFzZFcdCEAi6Q1RbKJwC+GhtdJVpj/8Vw55q0Zlgso78DPF0zaWVUQnwqdOQTe
FTj0K/F0/lenOBR5Hgyt4iPjuimiuHpe116yOCgA0FLyW4F6ibC2Vv1KAMmV1Tel
1Pu0BRjWhiPEE9w6PwRd3w6FR5ke+vYvufLasiqLh/UH84kODVWjHwjTXepEPv3A
UimY2Lfzt6hWrjhYyTJ96Vs1nzPtBs4mWqTPXQNszi/Ft4bxVQuxWAHUZgIzWRjO
+qrmVrDd00Fwlh5JPobGih/E3FCpoe6scAq4BCykLt3VB4qeszHomKN/nfqNf6bS
BuK6B+0IwprG8iSF+mNqrAXV5F+VoTpryPnzM4cv8mxCyDumh6xGTX99+AXsMMjM
kSsKmhgR1KIhm4rjFA67Qw0foCkizuMrmIP746qI89gbAKuYrGXklHau0q+HymVW
R4cV9mRlWu9gy5W623Lyn7jLb6mZ/eRi4kcp4Xun4xVFTrhJpvwpIxjtlIVp8E2e
1Q7ItkYLy5BHpn52SLkVnYTdPMl1yhTPXjOGRi1QkZcuAWFMDENB7wuL4y0Ix17J
+sF5YMhpIXQNIXP90nnH9ApzOLbRZ6yqqJl087lIP2RucKvP3PODYHNrc96io3NH
Qoq74TgvMZutFpjkX4QFxQk8a4jYE0M0GJ6595bluY9BNWJuYDVbojhJ9+7UIGwa
ryAV3S0zfCMiufCHppPBI8ZEgJyQj3+PGPHTsPTG/33tTdNdROmsFZTV3VS5xQrL
GTfpBrltDUz+wk2Q1s077UGdACokOb6U0kbDUrwU1hVfOZX1sLqvPvOSndkgixEy
HWm2+5BrHx2bGOSxGKif6yP5ehfSpPnRVO9zdMPX+BcFK6gSSvU0xoXwk2Xe9ZTS
PBOvB8AQM3slIhQR12kDQsPbYeZSxBVju6W0Z36d0Mb2Ja3VwKKson2X1+BsruXF
igXLQD5tpAGdOj3eEGGtJ1AqNllsyRL2GY4hTuTM0azYZ4KTCtAoDI0nkef1BVeq
BgcONyV0mD/wW3AG88CVS+ifQCIVNvzLpyusd1mqg7gdZgJp78d2rl0TMZyFUMCb
mn00xKHvTJarUgSFRVt30vxshGnTNsyRUO9gSecWf9Ad/dhJ7D1xnkpUQdWyMDwj
PihmjO1Y6L+q4rCgq/xTB5rb80PAGwrcdHz4SHl0tSXMEdGYrtN5j65bYUzHkFJ1
ZS/imcvZY1flR5IGIDMfrE+VATgYFagwdhiBS8LFNyOU4QXWbQEL+kxTKW6uDSwi
Xsi9OXPWrO3agrWHKrPu6GQC3V3ggYKknPaKibcZy+snptrMQN6C9yKa1b0eepis
dgmt2hTXKKmqY39wXSCKAPP78lYcdsc3hw5Ec88skKI6/zLlvFFqEY7AH+tiG+d7
HQrHTkWhgukaXOH/sqdV/7eOQWgBGYkqqRgVLOTiWpFYlzhguTuJnWDQTapudPYN
jqo9O+0uysjAvBJ/FNRkEq3o1/CuoTC+NYMmbI+83fCAOhnU98DV1ytVLR16HXbX
8/7RORZF5yQPE0Gowguqx0MSrGtsNctbh67Rs8lXR6P6/xrEnaTZeQjh0kke0ktj
WX/au6X82Qu7c5D6c1ds8xvXgRQ4o/8oivdQ2wInx4XltRVhe1G2rPEHZCzKaeCa
DyNG5wp4+4CAut6tnxDbX1KCvdZ5Q21QCSw33umV9nadMdXJV+KCZj0NSqtrWtpc
SM75WmM/YsRA8luOZpYlV3D92CNNzhMgRVz0v6Si8d2lxXM1SFHfFvyqp5f5doAz
hGY8tu8qzu1ld6yZrzIYx+Dv5NCyB2dDfomgdaNBoxz1HbF7yYI9gId6OaJwy4os
kgITYQkWT4PPdtdUmg25QOPViGvq0aP1kwd4OxNF/+iAS/2KJmuATq6xgBSFPUYu
8DsB0NZZsXQWgm6tg5LlxAllqZlYfZo+Usj7yWeCVTFfCv53GrwQ8re3sx/ALP8x
sh0zxJuJfGZbY/By9Bu92lZaEiC3UR3V8LRu4EKgyaKKhO78TBQ0vdtX/+8B1xBr
GL0+rsauxsJONmNlOQRw/WV+e3+UVNQMx/YS77gYOl9Q/CC/XvV5zSSuc0AdV0bB
d52Wtos68oMDEohSktnnJ5FgzMB1CxjPTQvk4TnUfssxpPZLpogXbrVM6hcIkcDe
YVGaYjjC50IxRHnJYqaWUrOsncZmu/8CzAByE31BlSyK0kfd4VO3Wtfp/5LM3URu
aRBVDkkBa4p6lrl6n/HtgcaO/4G/aAstaN/qZO93NGI3vwJbcw9f/l/fzj2U3Lyq
/OYCXFrDVn2JQe2cUErWgU5LemHSUgJPYfLG/CCnozJViTLiX9lc9MUrlj8cDMpJ
ZxdtXtOGu3soFoz9oqw+aaCyGvZX/uanX8/P3Ow05fPeYJCaVoR53gFkG4YmWfIO
UUxTogBbDvQXFlcvm9uo8oq8UJs+CXw3bPfU7QeaUjaEyRJsYIUe/MrcWszZ9bH8
fio6HmTkmkRMm8MXpGik5rEE0T4GXw9tkZ2Z2dwkGfvgmmF22d0qCpFWYFLquZGn
mvt/CKo4de8Kx3QH/BeIi5xWeFA7voR1K4jFpZK5DJZym4hpdEOx0A335iPqAFaw
mSbnb08UR0JXT6TtE/gT9uw1Lv01jQqOcPFZ7rmQIghAR/ZVQAdzcmKkEl2mVcr9
QfJ6V6XfEZXUOjs+klhReVGatkr1yFgRhnEt6Yh8+WFOmq/bgprnjYhzY1WNf630
fYzbgf/8gyuGTppOVSS7XIcZSYdKLnu7JjL4fEa7fXbeqXDYtOatmQLrA8CVa9Am
0p2CpKErFJSozY1K5T+M4ZVl3INi4v5XRosO2fOssFiADtwFNr6uG5a/TH1SGQSI
4e46Lgw7gAfUf2HEv2/tzjfWZ+AcSs/+7Fm8mFvhaPcz3C10ccFbLjVe3TppF399
NNuBG/NRTD/90lyn6bphyqDP3zbjTAUZtgL9FlmnCQB7YrB5hQaGa+RcRYqdkTYe
omWAaNKyrF4r2T7AwNun1cfwj9gfo6tSeiqsXD6rT3+GB7BTg382NmNgnT2Jr8JC
O3LUhS7UIO3N1XYx7Q/9hkYkhwvxsD2UC0IbTKyte3saGIfRy5CcsWzF8IdGl/a4
u9xVdquHePyN8OWSyba4or5nRTJ5MlxPi6gHTaFEZjYwkROvqn7LhxLGWjWcJi+K
9jLVEYw1ztq4ATDyIRYhrN7adyGeLQ2wKMWXxATOZ66RRTdayJx/SwA4nPhJsrxJ
nOcSR/6gVm++9P4a6dieLdrKfV/JVf2m22vDos7ESNihS7F6KFHtPCqcXyUCsp+k
aNDj7/rSuST6b0DWOjjetYCRHrpnIq23FzTyA3XsikQRUCC+3TzRXHqlAa/nIZKb
cX7cExuAFO9Myixpo4umtBDySnT2yoEaOxnwckKoCpDk5RmaSj0/vODt1EG5Oxaj
agnpn/P7sQVYkoAM4npAveqj5tJEpb5kwndFn/I+YbNzYsoQtULIME/Npl2sOUJw
pU1fUtVhn6w+WT2oqhH7lrqh0+bxdzlkgKDN16MWsVJnVP+qDL/m4GvSdnzsZx3Q
XcyiZytUCOawXEDnNd5wbVo/RXzAjlemOreKigwWdP88JUKTdULzHWhFjG7csH1B
s2Kr115DOYATKaX90pWDF5rdOh8dZ1FHNEK595TNmkTNlS2Z5ahI86bosIY523MB
JeYRjuydbXP1J9TPnpqeSCJgRBcK87oYTV0vFbjfRLijTv8UK7IF86ApPRjqixV5
JRWazXt5NgH92Nr3D3pCLzI6MV+nYBJc+nuWxCs0oUWFY1DWbjAyopy1UKWhxQwf
DxcLz0MZpcDaSPQcB+cpcHz3Zw2wy32jEYMJzhimI+bz0im1CTQgqiSaqPghqiML
GlI2lprv5gZwJJ0oRjZZACjoEORx8cMeKhkLRfWCoOFQhWG8g2AyV6hU5WB6UgiS
LVa6Reze7MFMSv8U4aJNdSuMO/Mq3L+9KfoAoV4EacjsDrin9v4mFKU7IWYIxKPV
PGzWPwGJtP0Q7x8B6/91dtjwKQJzO56IfDkvwiKJ+SzeNPL/Uzwv9bS2ZE0KdkaB
eqnwCTrstvk5HxpcunJLbffnyXl0Zi/biyjeKwLKJAuZ8bCGjnhcR8avMyGWXgLV
6iROLS6yQHgAERiO0Vkc+vPPSjpnbDa1pw4XKmHoFJEmEiqneyhdI6ENgyYYmYNC
22wO7uVOjAHPXceNlagQzqSycw9EIwoJZjAjGN4djgO4OdMQEf4DtqLtNd+5iSRx
Lk5bVqWV7iWhp2vPN9Y1GtN7yOn5jh8EccHNpcHTti3RdX9GSHd1v7Th/mVJTqyJ
aIPltHXxr4l8WJEZelPyOox7SnNOxoMWmF4bwGtikke5gbcrFsF48tHxsymbalKz
E6BcqGRFyztDKu2DG697aHAl8GwMqBxm2/FzXg11kuyHpI4HccErfO+h2oAEYqKL
66hc0/HPHKLDIPDsEf78mi4Y/SildZ6hXnZ8I79d8Duwj7Tf6SgCP4yVGDLpx80K
swlTDmkEIFLHEnGmTqOSvWYeSA1Zz9GC1au/KnOpOfbbQ8X2w/JJhFsM75JP78Dh
ZCIj/YWr4CbEMsjyMDsWW44BztRXwZLUF0+pnGaW88OxXk5kAQzbJJnT+b/5ntJ1
q2tVePHookjYuOINOm5aMif4HO3IadV7tZTTcCi1moBzBi7PDadF56viQDIlYUqv
UfLHAfdEovhaiYKIw3p02BgzisZSn9xbgRlNQ3KBCA6t76JFpU3/l/hK7asFlAUj
5pK0043y75eZIYe3bdSNQUe7sWbsee04YE2lRguaxk3fa46D4HQa8EpsitI7l61Z
1ettPAz+MRj7E2H8101OvKD4IESoY75TEZmBhAtKMn1e8jukf/34J+OuTJBn9t5w
kG6RrN5l5PIYXDAIiKP/gq8r2wmKkkxb7u6CTx39mtzk/6N7DJ4VSEfeenh3iCoP
ighY+B5rggfIlHXiGVU6uvtJVwCsXvMVzCmcZ500UX1wjUbUjupLtdWJNspZ7ca2
Ls3IDb/lPGxf66T1drHnPOkGLhxtqojG5T85pZhyO9MK2hz18p8fggdGWdZfr8cV
TDNg0jqHFoeALl89rZqZiGnJMjxC6J1G3Ke/RfzUp98nzGBuQVupnEcNa5Hujl5A
Q6+O0RpJp0lhoXtqbrLBjFGLxLwi7QNrQqCIcnd5swGr16ASpykeA3I6SZAMJ5ew
8gjWxbOTTY9amOBfxBFoBodfeVbIOi1PikyH/75YLcsg0Wp4QK63SKYyMtRtomNp
Ef1WUNQIGrvqrxxE19nLTlxCkAm8nSOSq0105iOD7bOwbehTAqFqYPFHYfk5qahH
qgSZJd59tu0wIg+/VATyqbtFKEWxwuI3f+qEwSLaQw3ncme8JYGXz11U+5atYlcX
15ViVgKO1/YYvcdyw9oAyrQQXGiHvNveoqhNGaBOa5oI+B6gzvh78Md2h8dV15QP
PrNMOH3gh9P8Sh2LOunUwE3IB8aYlClJzipqF93cOHKxef3UZ1IQxFmHX0oFPAro
098+2Sd4fJPjgIOsyhEWet5/N5KXb9z0l0/b0tkHPgqy0HF5JdyKECd9+XaZTsj+
Btpt7BVl2dAZkB1TEihe/Mjhjm09pyDJPgH6MKRmSL7lPZUqQjC12m7l2mDUmQVD
MEh/cuTArtgtm2JM35XYljpELZtBEgNZpdAcHFDIzuXEFX/WYPDeAqSnUuiWfuOd
CO3e50d5j16BffekUbKOGLBsC5dMZrDjNRTBfrKwOBCHCr8Ps1sUNNp6rCA6uoE1
V01v+qicbZUk2BZEvpKezXM0QQIiXAdOMZs0iwt+Ka9uQC/nh4qKXyJXbI9Qzavg
EieRj64tG0FmrQxd5WMC0MUHa/vUkMigmaKvLdzDt9w0ubzRzM/0dT+nF8/x0Q61
P8ksFf3shYw2BnyCwQGDd+WCB1FnAlwAr3eS7h+ntkx0mxF2tENrj+jK4Ly9O5NR
Ffs9RBz4DWDOpRlORzK6w81NyZrhxRjC9rEm5Yqpq2gk4nbvgxJQeAWHYoj5CuTx
UAjE7GcQ0ws0KkuQMVY6/nL0F5WwmmfygoSIYHNqazOj2liSNGZjeceUDjjw0/MG
Nfb1WRc/wSpSFY9PQDtxgNu5viIX03YHzG7udYxSkmlUlqObXSkoDNq9E1JCIAxD
/YEaNnWU0Wl45s6O4sXcEDMrEk29K3IOiaaQExK/XbDAwkKVIf5H91miX0KoagEF
BldjajRuwDjxEv9QXKjKzyTOrtSeQDO4vTX6AalsBXywf6ednDoEYd46XFV3eHJg
Kx+rnkTVCZVvClQmn3VStTpanQxGF47iCQmxClegPWVuQemuBqnyB7t8WLYUQEh0
xKJeak+c+95+xlxlXvg0HryUazNn2nmdR2jWVbjoatW/J8kDBDJtiLcOjKE61xKO
HGadNewnZZcppZAEIcwhLdYeBrlp4lKBs/Uk/7iahiLglM16O9X/hy6Jrts60f0l
CkVT1NpPzNkZ5pRpPWiQei9VqCoel6Q/eN9Q8v7tTab9pDZzWgb+i9PQJaMSAdBp
ufHlMYRXLk1gGB4GGBtHwbGSJ1PJr9pKzpTvEcfbMxMDlQf4rUb8pUOA7pW98wRy
pgzkNAzPh5RgBr+aT0iIphL/xQ0luFoiiNGJmjLXx0UPJzPmzMrq05eW71aCNHfI
jrwU1QbOi8N/wP5AWi+t/WkEDyVTZSaMwk7wfybuXW/2/sQlxiLeL80f6y8vuRbG
L9Kvq3QlQBVpXevUCSaKJcL1+qgKT71WmXmnFhpNjnbWo61saYP3sqr8rsXCVpjd
gUX66TZtPy8i5UozJzcpqp4p791ZIOta2i5GiPtG7j1KovsWoh79u5cTrYD/c/A2
AhNIyNkuLdFVxDY3rYQqlO3B99uHTF2n02J4+Ir/EGvxXgwbS+yI9Y2qqaDgvHWg
a/OIF8JTp6sCcJ+PCynK35xhyng+Nm7xItR+VmM9xbqgtUsI3NeoY4GLHETz3eo5
mjZVch9/bMYf00396DqoSxz63kt2eykFwcAHKzhz5EhsAki4wpyu/VMPDl+YTeLW
fvOHUbcy+w4SiKcAWJae7GCLNz1x8HgQeMt7gHFvQhUAQboxLQ0cB9g+3WNeNhw/
KXeDGq9cnxAxPuBNImstTOLcOcz2GxFJmbeE3gViubK74fn1AStyBgrOSgLW8hKS
ylxJIAWUoUXQMZu1kvfX92TneiiY+XYBASxRPBnqT+jL/oieFqKUYWoXnF+gNWhl
xmJxOjZGm8bna7rzNtndMuELH1iKPboYZa1ByVULk+aQzP/rUQiSjRQuSSmy0D18
LEgxty/Cqp0C0CfonlXCIrFkxCPtHkcDag1oLMF+FtUXPoHd1alBQb6r2RJMUySt
xTwymkS34Jh7ec5A8PPR3CHjh+IZ9xJpq3DTjxr8ghj9e9pH5Pc4hox4GwOXS/SO
PwjZLVPb/wCR4Iq3YUV7R40T9ei4KwJswg+NBPXqAkJgUWcRPf7xlUPsMb6PEREE
otFPpt8mEGen4WVh+ALiR9fdIWsybHFlL/ZqVEWs9hMyLzF6M35DKPHJsn53ImBV
wa/iGEOONdkmpizSkGfCIDak0X+J9cRbrdxkoeXn+zLfK9iEkdDyUmBUyGTFb3QL
uc2Td/Q1rZ/3rcjp1TThwSBq7EbTvNoTzVUnZLq9fdBqI2asri117cBqcTY2Pfv0
hNpiHQk5sUM4SeXCf6wQQOyV/6HNUYYoP4gU6FLqQZfTwMCYK4sbiGIa7WUuGRo/
RYVzQmhLxXmulbcGn9ySiCT8FjXXM/NZKL2qJa0F0uSEIK3QsYVsIDcHJsxBVwvS
sRoLFRacQxrJGhDeiMxjaLlDm4+2whBBz2pleYdRZDc0EKHsxrU2dji+HFF1YTlz
SrEyS7quro0VPOT5DJW+mQQ2KUxhJBobz3QbvixP42d/E+q4WkQ4DtXbqIaBwI+s
aQKlteKTnU1vEiMUB0UpvWa/7sHllAVjtBs2kSUPn96op3bfUre+swSxvYeAHQIq
2wxidJRl5OxUMF2/ZBYPsz6xHWHVX9UAwI1yprrLgen9Li4jfM68ph//ZGM4VOH6
59RTIMc0hKMVHvwlvgiC0IuzFmth8F3JAsJXbeIq7hxNFpinZieZdOc2XtW8Dx5C
/1CUvRTTvv+49RGFunQgeqRpa4B2yxK4BqU2Ll3WSSYjq4o7kaFALDwM/Uz21IQH
HJ7vrRFv0kqGGkjqnhx3iAm9xRGnqn+oZiIf7kdo7jCZewWyhz9FFgIAzTYspc3q
51Mv+p6kfzHV1SAxIX1WMLs6evdjjCwI3JBhKSOn6A0MIDnR6/D4N6wvtpSsyoPj
qMNwNkr+K9welHH96QNLhAPobonc7N7lRCDCjXuWYJizq88wTPVfjA/Rzh9e1sUb
BXNPxyuviiy3qNteqbvf5cit7MQ9R7jzhkrqMj5TaoZEfrecC4VjtVBYvVTOXkq6
ezOVwJ0xjGYh9rz7SfuOF/2/1uOo3w+qUq0t/U7Oos8kDuYaK2EsuIW5t8YqbRZd
2l2RAwXzYlTTARjdyogXeqQKJbXZ3IRxfEC+1dZf0qS77RhcPMh/mLqXTeVyhqdc
7Nl45hMuP2aoeOOWILqD83YMul+m+g75270jDJR/CqkpAfDdCOrX/W5o5pZh2YOZ
1jT8OkLcZV2k46QbWuu9WJspeD2lTaCEEiQ1LQdnArWaE13XHtr2gO/G8mc5KYK7
FAiH0llunDigXzF+Dw7Eaf+OjxEWNbMPVYzCJQJHQAworDuger9ibwcW+VR2OKbv
IQ4SaHW7NJQmNcNNZ52AeClH6FaEnYcl7ZpsV9pOhMdb4mHgaTAe2Gu7rgHswART
68925kMsnJHJXHkYLiQ7ILSiz2QCYSKj9VYSrglMqMKgd6iz2TJzTreOt1Hu/XTF
Os0Im73J57CYRXIF3FeRKCh2Ilk/aTp9W5MlaHbkux8X2Md+ZtnYMeeKUyuvV/xG
ZR6eZOncvSclHZO2NoY/tlbnRSQJHpVJr1VsXa8SNkKIJgnrTiWLFoYN9a94njhH
g7y00Dpxq1umaF54+VTJABbnE4jge2xKbhkId2vGbLmz7TFjctkGQXZWYj1BO1Uh
mZd4WhrbHBSQ8to57i8wdZyMyxlzh1h9InTNXLADBdDUXo/Z98MV4CUN2EpfQgWU
NpXwn00NpBgI53sOrppUTYiqbigXVIZ4873CaqUODzdpY5lDKiAViFr0pKZ4UX/I
fA2Q3tPd5ZF8eUMNVYlAI2W7He7m/xJCnl9iaJQLV9psYRNH2gOZHMEqLvBcHPUs
UZ5k6WkafLY/TkWDIK6cM9uo08dwIIT5ySpIc566jhs7EhZnEw2v8pyKKnkYjh06
oU72xPiZ1gFhuTKXT+YDFcl0xC6wqI0fykmAU7g7R5vcei8fu3NctoIferm2wKGw
359qJNQIZUyZwo+5dLFV5h7yCFobT6Gsc++LOgg92nrvi9pekK/lO5FS+rTBKEK/
U7kO6e2RMob7B4729kakrNPp8/Q0lf2/HYE8cxQ6vUKW/1nV84xZF3cwrBYhX8Mp
gthtO34TLzafTHup3opkmx7ycNzKWlI7ekIMw9puzXtVoQayWmD/PSQhFGILp2OV
2U4f8F+1rvi0Q4Ix0xRa1SSv3SsiYfETKfgP7S8kHVYCEx+I7PqtK78UsNCjfSFE
TykPgu0URU8Md0q6uRwv4MjQ2meRBokTmSFYPbVjIXipNTAJvUg0A44k7MfbOmKd
ND50uMtrVOSpUdUFdxtjCZq8HlgF1x+K91RlYgruDdjIk1QlBeZJtP20ur9Zzfek
7bQ0C5vgb8loxDY3L04sUVP8yHZ+brBZ9xMWxDxzRvFU+ZQMZVYiB78ylKbT4+td
H9GkeQE7B/xp4rUkEwryJCHiIZ+X40tI7thmUpdPdEAP469EtIPrjlS3bxXIkfr3
riCD56BmiyfMAA5zk4FeSiFe4fpqnSnFOlIbq+cgJDwVqeziybWwyEr4QomxGDeb
dST+yfhhcm86yXdB406QfaQAs+OpR1TGxEJDdHWt2gjdCDMFC7XImNnxA8DZiWTE
jGyZgM76fNQw2eLHmpZIeB65PsBwPMMjAymtjVbwaEnx1cptmNRHlr5saXT4bREn
qxAAqSX20lpQhVek8wv+pxzdzuYB5Q3OLnoD/f5WtCh3dLahoXxa4pXgxv+eL3jX
OHpQtz6C3MW4z9vFosjUAUaT9tK1q538fjXK5y5bFPGrDr9pVmMO7pJZPVopOkGz
AegS76GiFg90gLEXNOZ8ELQ5Rip2rZEFOoj8FN8zBYY6U/7AefJZ7GWnUR/zSjpC
bMtQ4pRdsYoesRXrgsA5O/90DMqqBRaD/KpYfsgx3MIhcp4lG2YTBbeTUGeq4nT+
4Aqr/BJCeeOsrrDrMVBWxnnl3DjgFuXitEDrM6P0pP0/ma1YdkwXtzzDlrCscuiE
meDUfQQgToHL6RvRy8CZRBvPfv2aSpMiI0SANAHLYCPeoSVSAuP8zikr9v4qGF5b
amw96HI/I0vV2KVXZnf4fuRnsc8WvLPDlC0akkHaEEZlmGhYyg000lI6BoZ6rI+6
cOWUaMNcGv6C6CNFwVf+z7ruWLO+5Tg1IR+0nbn7SI3K4mobF7BGEFhN0+cqH/88
oOxb8x94YX4iruujCW0nlvHF/b6az6298b5OQ9IQqWHNWlLVKO1YuRd3I4fvC9dY
e1EYeLBVbYhDyeFPxkjG4o/bqV1zpYRoQiY0/FNv2w3GWzW+ZzeFDOAlrxpzPWeP
bZvGoY4XeXTPc+cGmWjCuwijtHXlyEYC9I9WvdYLlNF1h0LjKUz2bsyas5agZXAB
kA6wIGmr7IgP39JFrANG7IQ98X1Qgrh3eMsDLyEyy1fhy6AWdQbN2hV3Bsw3i/fF
8eRPQAUSzU2pn5orA3/1bIkFFIbghIfi89pmFIPvDzbOkZBU1qloM2e+j3rJ4+6k
jzR0kBdNxcuCaSAJvLnkZLvSkrjd80OKeF01TZfps045Ezh3xZH7XUb+li6c0Ksq
Yn0AgxGjCM7qothgk6wEw3ce/VjpMgnKSP/7DQmHgNIJCWwNRcKR1/ucqOd1TsYg
r6MfiujZYyeXdOyqCsVSIvnyXuHypsb/CC8lSqV1IJq/jvcLU9pUWKF2lDADigQh
oov9gEkFXbNiSs1k7F6h7LdXCoWkyeMJ3gwEfE5qPNqffDdN9jaCIau0A9UsyBIC
VM1yIAykCOjMsyVk4OQMa0IRRHGPnqg+Ig17X2gt5OmCecpM+fTABSoa11yWnJTe
lJCHa4hTZVPa2fm10y8wR/UAe2hy1OCUa+MctUOQFNUIhN0ht0ZURSPsdcoaixHf
neR3ibK5rrADxRlgNJpfI+m2OI2zeEq2wN9fsjzEVnagBz4DdeYx6IP7pxacKoQJ
bm+h4Tvxjipzo/ttbBL490340nbTWzJkj3tqyTD3xzpZRUuDziU6udxxOdFjnR4i
y8n7CpETxGriqZBR4FoV9aC+HDnAhVNA03tCceFf6c/cKaDyi/QqzcTcfZdjHQzu
cC3tHVJfwSIZFPg6xh5s1nUMEkRCyBxTy1hM+v+QfzXmID/yHGXBAnj1I++VnSEE
N7m+SJbrxkLmsLHVuMoIayBz7u7ybrxE6wycU7potw9zFS2eJp9bOkbN3vX5MRBX
qWD2GPnvnZFtNIpoy+FatX7U/y3GbR3C7smfAv41GYzPP7mwNleFBSuyHzPBPNHj
pyO/sdQnhdTsya0wL1N+XrURyXCuPMRIpNoepnWOujvM/5gfC7GaqjqRjlnnNsMw
ssJLaqC2eyuyoVmcRnPKPkpUYIWyryXR/lAITuKlOIPdr+Npmcx7iWuZrmGsdeBd
V0Fi9RNQK3IOqcleOi1SKOUzC8PBxlGY10TsRI0XPTTRK/s60NU0vgdmhub2XAdV
mhyfBbchoLm0pkroTJK5OJWwBqC9bzo1WKBOM82+jUdZYfFVt+4kikS6AbFEidJJ
QPsS5ZtQxrfeqP2Yry7kdN6u/nxdPy3xMxmLimK3qTiFS+FzV/n6sb7+XJAWTSVW
Xg0nLwK3JBMAiZnKnhlecgY8ANzxJTT6LAlHGTh46431yrpL0c6dnbQnklFCZy7G
b5JpLTcqOAtGPPvNVTgR9muevSyZrxHLh2lAqDquxWGopVL81sEu8p74tv1D+5XJ
6maty8IaYqrqAPd+1cfIpUVboxRqD77A7m0H52fA4PTRuwPYHN0k/cVeGkzRo5aK
HK2pKEh2HeJdrQKS0YGDLJ37OJ2nYSunDCtYzuTM7gPwOenHHLBnuLGv23rm8Qu1
vyUUXk1k25oxpF5yzPyseW09+rjotRckTryqZ+J2HgJQ2p7HqbRRYSRQcSovtcWw
4Y1V0zt9DXOV1FAqKMQIlXPEoBosI3buqFyS7OsArHd4khXbtJvleZBwo7kfA8Kr
ribUkMF64rWPkUf40QpLbTHgAi3ThqEyXt872Kq1WPPF33exCmYOX8sjr0GwXDKs
wqwZbJwpZR1AspqjJzZrhiONCLguNi/Aj/+PfrvQot+PqkzSpH3WnLxvDXyVPQo3
xiFxn/+06KUzZFfWC7jE2VmYRPkq01yhGQbCjM20193LlEK2lN9lIpJZhBIzPn4s
cbG7fZ9QZKjChqu+CQAXwRGWvxGPPj1PYmvwe2DGeZA5o/uV+nJphpfxC052iPZh
Y+pLzO4Q2q12aXV4XTWkbUUFjTH2ybGwoVxsfkC2IyeQH2dnTKhASw/ecUR6ByNE
0VIqDmROaVi0MlRVSsQciYwEJNHI15ekt0jrLTzI+fEMUSIq/StheOGFiVXqHqE0
BuJeG4pbjjy4esmi9eBDC0+NEPpEo2oS6UgERYpHEseRPMi06CDPFIUrQP14Q1/8
rd5+tyPSLl+pW0IrbJK7bHG2UkgoEKPbx/kK+dtqHWfjAVL10X0BuW3fx4FsDuJz
+84vwMp0AIXUc6lI6N+jNMDBIuxc+KNbhsA/JgGS9bHJABhuuk00l8A9qQlmM6is
vcYR31mrgppJH5ZrVKdTX5x37Cyo2ZrUXB5XwBPY+uGDXY4cDaYZIKEQpEVYldvf
EN4ysewWgDlMIb2XKXYWPKYdPkK8sZZ7Ay7/rPPPVsBPXwcsH5DUM2RXAlL91eRu
XlFTjimcCjgfOv8f2R6Eti+hPEMC6+1QAtCO/KA1sVdZmvEObo6G5hDQcmVTOLox
3/SDME0Y2NnzMzm3hQyOr4+r82ZJmgxXXkr/CnSDFAUBwrQ9gKbn34rRAauzv81r
ZhCc9uhX+tqTs+P1YyEThLOMMIEaXA4wrZ2nMlxCYYcTz5HXNTssT0lIIEU4DTZR
U3ZlMQe+9BILpogXnv/jQK/GdrNOivn4l9jLkiLZTEi7Dwi3HijvcvgEeG7xyJoY
pnq+SHFhNs4CQ0AYvspVeueNxe6qkQyiwfDvitAvaHGSw1pKNlWfHHHU9D+YIQre
9PpijS3RnQsa/xEswEGUbklLO/zFHfonWesZvXeew8TXBbJAYgOraMVgQVabeCfw
YstYC41jz/f9MaGGbhqBmTuQx2Pns1ldIzfc3tC9s6F2Ih9yTHcT5mZmOCeTEJWV
0EToYaaafWODLrrHfFpcERknImqHfJPZB9lVgmCDkqfOLBAJQ46+yab185iP+f8p
kOg88BcAM0mX67OONZqOT3NUDi4ZQR8NwZpxADP0MzIS+Am04aUPNJ9uEnHTGXoh
a1ll46BEqmQweCJs5CgE5HjLDAf/mcdh8eQSe7fPAtbcaoPKWNn0Bns5bPe/9EjD
Sd2cuXsflc/M3S6IN1ucBKrRyJ5H0tAv9c4ZWWQaT8ziKoLAILdQxb1v4EWuqfZV
pS6+wX7PZvR452fdR9FoKo6PoYu6ZhhTMRY9gTNHBKsxAV1a0EfC9gcgs75+JP60
wlj/4ciQGcz9vqQPHkfhi+Mr5ZeZoS41HgF1s1gNW0+kpaE7X2hszN6CucXErItJ
YfqIqbO/OB2URDZIgdwPiGHzXqXOE7dRIDKSax5hy43+jX7RME1uanUeuw9QIYX6
8dxZW1hqk6loXE1UU2Y5UTJ4EX7YP3LspHEPofRfrjPP6GfGp8nMWNE3HFRtXlyW
zAmo/CP5a8HK4N7aGxzjcihv3OWgqA/+zLJpl9S4CIT1gw7RqEtwA7Dqay2Lk4oP
QKQ/T56hpsHc8u/QafRzmslRIIQ4faDKPccGuqz7Tg5LRnvSlHqdNEEqyrgQHuWt
GvEnQA6JLb/CYFhj6mZF98eS73em4nxQ6NR6yp3DeE3PdR9M3VkPyjoNBYWp9JHs
nVXq5f60q+LguWTTDBPBQP+4ei3QQ5Vi9IObmBKetvmX+2NRHoYhnIBeClx89tHd
XXMYi6LrGQo3z0FiH4++OmDymx7/tbmtSyLdagk7m4ZixOK9AZ1NzdQvxgMAEkxk
ZBnO65W+3oPJw/YbRkmD0cJslwmGx3eu5v2fAln4MlJKLSTVt6f1UvgRzg6FufMl
O0lyBgXUEvKDofirHDXyL7AFEvG9aB7vcUbCDmcQdA2AWFv3MqVsOkGHqbtEgylp
nKzH/vUfVwDYL1FZdW6iSI28UDT/lVSNFIikq/fHf1fiz7Pki1bMjWWrgSXITusv
ywQ7SQiUOJKtuXWoRFvQs/0NNFqguF9vRdIYq9G/kg7SiYRNdQeO04cBiFVNvF6y
AveRZqyFU7c+WQfaj1LS2B5zR71PSiqohP7Euej1vj0vveM6ZdxOFD2CmPhHFX+S
O5sF0oFkVjY57bCjNrXh8EMaiuHJC95aZtusbG75YTz9E/jXQVhQlCvD3QpI7+mj
ACg1uG68rKM0nTMPpTrO2ca1dvYWCkC+XZwphtTQ2laJRHufE6GiLuFJ1xhiqROQ
FRaCFK+7nShYzBAM7xWYg4UmOGtH5m6b6AWL2KkrmKeo0xfPteUL9enUjUjfRUec
Pc13KSi9DCyrC1vyRrqK20omaKKTE5zUN9OLJPkHAe1mhV6Uz/yASWUhE3NUb4B/
SvUc0LKveP/YA03xc0MtGB/PM0tBinM4UI+GzzhnfGahIGpi9oTQgwNILSWIT5GV
EF48O7CP5yeZmyQMcmSE3PCuNXeJM05SydnHLJUjvtYXLPoAO4rf9SSb+FoLkXMR
POeD5JleRnQB4VNYIifQStREatGfJnqytPJwfKPKH0yIs2X/CosIIpotQpjMUFIC
LM1wYaUFCdojOf4CsyQ98Y+RFeOfwxbchnXHhdLXa/pwYEa3DRiKaGBmbHMHpdN/
QuDfyvzGlwbK3DBeP8ACjyknVjp7ombUmwSPtZhUdqmI/rSWDyg8WdHBjcbrKQRn
L9ONiAlhgz1WS6mhlcfGA0NEGHVR17twhvqqpPyenkXqXfwq4loV1FowN8mb8G7s
CJHs64tDubtxwDjkueT/ai58tKBCh6oTeDRCu2CBEXMQ8hrQR2PjW8xJGKkpzs3o
zj0sRaeVYkaxr3cM4h968zj0YOSgNbExcaqvrYh3wco9qarU39RAv620swT75DKp
xLcnx4Kfi7cfl5mByJj9+qNDbZYS35R7RmDuGHmTUwaw07CEiQgGpvSyURyRxHbY
YCnnoXqZB9SCjKBWvRx6mFKZg8ti7YcCyCm7d4RMf+VasS0OZTuFKzjlG4i/Fg16
7aSzonXcQfKelhNBtkKb1nomrDdeMAMiAH5muKNGVse36pgWJaCQ27JxaxZRtQQ2
6I2LiSFMp4rhrbzMk0H2z6L4NQDa+SyAftjHdQLyNMZZAAQuTtr8rauihhDLkE9w
iwrxukVkVeebfIAx1zcNOWiQPm8zVB34tsDrehKmlECZF3yUcVCSfc6yXsvfXSxt
PByZ4/Bm9Qds07/NKheoeMG+nK5US/xikqdQgR8+eX39+HvYB6ljTW/P5GsTG5xe
CHkVxMTBpHK76UlHhhx8gESJjEGDprOIUiDOZEpHzFn1ShCw4T3RlJkFlSjHMois
If7qXSmSKG6vUfM7W5XYmh7A7GpDf0SCksL73ZQoAzbRnTON5QaO5LnwUEhw6X1Z
zxF314nAde2FNMd+C1bkh6QAsbgONEtf0Znr6akxbDxyV7Tcp6ikYKBpGUqp7txZ
9afTFgqJwc53q3DydItq5sGxCK/vue7ecXcaoFSFB0YkLSs/MaMnZ6GTjEeSR6OV
8Z9TBTMWlrKs0AcJgXx7ItbGhtpaal8Jb+Rh219MXk9yZkNJPAgQ+mw/Jt+jCluR
8YbZJXE8/xxF8y+yvm/DB9gliE65RtgFSkzgGwT7fHPSF8HZ2soZmp39glPycsF9
4xTS3UEwWkgC8upEcqm4EhaX+VYoAzhH1gNY5xbJZMA2jk+fpz6kgX7yr1efFmt5
4dSt4UJOgQNrm565p6H07BlfzeYlR9mVnFBd8NQ5ov+fqalafis30g6MTtrE1AZc
yV/ZENS0izdXVlgnoumM/Yg/r4sH9q9rgajB7Jn5bTRoOa7ygweHf2og741icitY
8GDx9/G5Ob1ALR11Xgmx8fQ24+Bw93nPJS0L+/j792KenJCVADVMUIu5sYThb602
3qXLTh7uLp9vJZK8kvlXNBN/dyLQLuQAfPLeDp9vzpayoDnqEI8QaIYLktC/L2vR
MBuBU1DNhle8cjeNFgNeHl0nDEBdd6kwlgC+fqrk2epXV1Gu0ePrjOQoQi3y0Sk/
qf1NAYl8qUncHKYfmw3+WaidcIygujU85W0FIhU+q43795Z+CSHxEQTeZdS6+ZZ+
pRT/TWnl5taXQKAo2AvjdH43GbRz2ZWCeniwgo+eZP7o5TeQ0guDYYzBJ+nnMaIo
kpQUJMhE5+nNLEINqEwqoSAw2Zc3U1NvMj/0xy/zwFCSVT1HgZLUB1saOvKW4xhf
gwwgTA+DZBXFhcgxOVP6ZPbufkpS2QXBIXVNaEvVrU8XqZUXZIh4dAK7hPoTtsoI
UsX5pOp/noJYH5rsR1tL6wRJUsstg1+xLTgcu4D5obfqFeujQ4faponUaIBfFgv/
kE3eZcJE68G3rjvpltdYWUUeP7Xsok/OnX2Ahta6euEjWcQV9XrDjbxw0+oof3bU
LQzHgZ87TOEir7iQLUjfgdSsxfB4YTKWe89m27+U33qobpAsWp8e5J2jfHCfP/sv
HhLnZnW7EEI5vb5xnblbgmfqzw4m33zP7aMManZO2eqqGURAAMY7KItxgsjIqTei
OD3g4R+xIDPLTvdqsQnB1asoF4I2E2uIvhB+ClWdVeBT5sfAFad74eE4uTHz0fv1
c5dciZl8++oX0lRos7eG5HDzD4nUqieRnJb2DY0fde7VRcw1tXa+IufLwbgJ5frR
tboNokadANcV2mNxwk7skha1k4t8kn7Bv10DOHKYzIgdfsGt8KswJ1hx6ADp4t3+
9FwOaLZv2YftQSPNe655WYLxVVlBD9JJyJih3wUqHDONFz6N4eOOTgb3Xbsnv9wT
YJ8Q7hnDE4UuHRvvQKq4zbcDC5G9yRVe5Dao4h4x7uveHLCNTbSLJmeYORNUcNz7
jnNGDIFnyJeI08FskSJ2UQip2jtG0+U+0crCzQ23TuObG5tti24XEsTLTJMsD0/k
TjcSziY5obF9DTUYurq96pgg3SNQ72yThWjQ+wM27H7mfE9ncCLJ3YCf7v6DOKHt
c1laxYkDfEjhPOL/W5Dk0cetSvbNzTr7w65rfAHRBnCJZEsGob4MbUqjm+q7ur2u
UJKUHelIWOnBh5XxH50ZXCP7b0rsa6/zlDDYZBsaAvGMOODQ5izwOEYbgsej+qHr
IMtwDq3tDjgrXVZ85PpWGFZrFj/1hX4VvmWrlieK42uo6BIuvxN7Z9aekymdYMlU
9SPDGBQqTxOTMAGiEE/eZo6TTY8JyDC6ISJZzM3JdFbfcRJh3I/ccut+M7C+fe7y
p+DJaZJwvoeYZtUg9+DOdOr+vGO93X9JfSyMLaXkEzZ9e1v5oGgcEsI+bKPLOYJF
/fuL5SlSe/vX6e8gL80YQrLPKWrbjc+mUdltVzM8dw8Mr1o7x+nJ5sE3bzpfZS/W
Ix5q1BNozYfqbCHxOX0y6stUqGVyuZHvO875PDNY2RT8ud7niCjUp/SggZbgQXeh
/iSJ1LnS4TKUn9gHEt+SeG0B980/QoqqYKjiASAuha6LD6PE1mq4z54o+eJnzwgA
jvCPd94TZX6ptMoVKipB1ov0JPEHmuaxXEoLmZ4ZL8U0+aWPk87ol+FytS9aHiVP
0ZJDmBKVxDzGFJv9BuHPrM4ia5pAMIfNc3mWQbvwIvBaH5ThCmEI2VAGQ27hH1od
H+ljByHAOZNXndEnEeMq5eRqrESnKkTQaNT/dfy9R5worJlOqIKxRLnYbX/F7yqX
HyObJZl+zqxe4P8/lDECb6oR8hEK80wLCJDebdp5AzYY5uPlSrgnl/sRJ/y84W/S
so3j1lQG0Ar7mBlE7NVxeMRDpU7LnA6kbP8ps8UNgUtWebayCJqAgE+rEFm5HLyv
VDz+YoSuOUf9Iua5/ZoPd7oYu4XZHER/U52z2r/0nK3JNX4mR80fY9A83yH0/0Su
66wYjUbyNQXzQABRWzFyTgeCs/EKTxvC8VyuBXDq6W+Luk4Exc08sCh6C9NSp8cu
roXy+dd2cF29OAxsJRPk71cngRn+0/NFol8NnGYLytM0xLcF+OqFe2+Oe1vCMIki
xBtIlhMXoIKHz+lJl3cg9GSUYYS5ULwwvwN2gh92Sghfrakdz1x2NcTiy4Su77Vj
09YM8sdS5fpOgJfANvOGVIOOaLxrI/wWjcLSQwbGXavEptICKgDq3aRek8ivyWQC
n0SwbiQIar/sovRYTv+7z0ODWMVnYy9szT4RwxRtg0566I0LQTQNk4pEUXbPoVUx
mPHicnvEQAG0BHL9auHwiprJPwUw5QMa9DTJ5aXDEhme1aBrS2BSEnehJGcrOync
EwJ8EsuN7Z4PEZZ3R4tIACfZB4nDfhqwOLRLSGK9cVpXtLrNcEoYb1ZS0ukNmpqv
m1uLz3kPrg8IHhMp3jQ9y/ukT/HA/AsHHUI+QXLoTu0VNqZvHWZ8Vo11idfCyYdL
2s9hd5GxPimlQPngAxuYAng0X2uGgjw0FY30iYFr35fz2/Rex/pkR9wwuuiRJ6Dl
6MO/8Sd7QoC1MHrRdQGhL0TkKeK4qklTgFuUpsk6LVdxICciWX0q7+3TgN+fTnGY
rhC6s5XnLPJHdXvWmiu/YV5OR8fp9QNNsfy0MsBlxe0EdjMKf1FJbqKHjm+66Wvv
xFNHJjx5GhbousHRyhou519hsxEUvRSs0qSs85patFY16LnedvV0zy36H0sBTQq1
+L49rsdFqjn41xJIz/lV9tUD9/7+Avp8ac4IvV+NCD9xo50goXdp4ozn7EagJBKp
Vz1U1cB+tGohhPoLYrS8BzdZjPqL7JlTTUzV0W5q52YFTBnHwRSbznraPZdRM12u
WX8w2J4JWxqaYHBtA/ZTprWKOYWk9XWRrp5TEm4cC+0HVyXU/6ATN1qwrrQ6AMhG
8V4dGKW6zmMA0ASvnGq4KDaLZ/yjoplQrVZOMSDeQuSt+vg8ts+0ZQEJPb99xDP+
Ssg3NpGc20SGqXQc3jtxC3fr+okHUQ/KgfmO0mCH8r5ox902FxD+bpdBt6Dpay7b
DL2h9m4LxceOUzBuSaDjfVSNoz3yFyesw4uitDGifanSrcbOEjbxykqxyQtpQAH2
RpWlJCQhUjhJOSVyYx7s2U4f2OP9kVpWsJE6yDsIMuRjAZ8yB/T44by2e7QTf2A9
emSY4VWlBJ3LD4r8uKmzgvlqeH69Ky4ghi1UCAWjfFqEgQJIf7GJ0o7XhqtPWPrm
ypY2WndkG0jvdyHgz+9TSAx4ptO4DU+Ec4Ub90xqjb4ZCeaXg7qzxqOnIG/xnVJQ
zijhOFPDdyvnY1v3OqK6oIJ/Ogmc/BmAi9Y6KrtL7wj2ePEgFSeTn4jfevIDfx5R
/yEZum5AnrYFlAREKibWiPm85Ytuwf/Na2KCSMNnL3f02Pw8qz7a4PN+iS9tgHnd
MLPvGQTLA6Iu9II7/vH4ilfHUjw1jyumFn/oSeodl94Fi0vbYhQIJnX6+s4LcQwp
CXVt/sbR2FpDxwPLrGuBdaLKe5HWeHhFCCSYQvdUfcVtlNvKy0cbBySC8EN6alMp
7FkmgcmW/MhRfkCI8y3VvvtjFFNcpseCZXr2xjnqxhmNpRh1rY7U+E0v2Cw01DT/
qQhs+DuJK8gKZP7ArB2TrGueJeSml9UlritBXiVW9GxlHAGkw/nehvLx1F8ledeT
0bEo+QINvJbho1DlJxgWvSdfKROcvMJRWFyJe/OAFD2rX5bfDhciR5gwE7ixxipt
1Qk0ZAdGGh/VqZztKIJNpNjZbgjH3WlNkPeaqQI+yovp2EmkmCK+boquigedcfz7
DjgdTFk0Uy7IwLa2fmIHR6cJXE/dac9DPndFC51P+oVaXzjK4hGX7wji7BFOAtut
J/UoT+R3VjklCEbgn+IejOUwP6Az5uuuvSfM2pY5NHdSmrK1qjZmQOuQueXpADcW
qEnIxXv5ann9E9Ytz9Fos4D9aKxHGUnp3U2lXeHBPqKB4JIPMXfC0I8tB0PLA1zF
aJU8fE2GBXOJZXRDqcTkLOivLnv30UNOoIqjYUK/LxStKgR8zadr9W91eSBGcBnt
GBodr1u20sKP5iSJIu5Fj/kKunxru5Zke+X0tkWzqAra8YoVSNFFOR9AjMZif5L3
1NQEL2Pkcd0EKW5TvxE0B+8kS6yC+y7zO4O/2N2M6NpBiM24qXzifRJpub04jCVr
T1E1MUBnAJDe0X48wR67TglH2I5KCC/NDVMqe7m6EyZksFWCF/ZTBKCXsfmwlgrJ
wv3oWifLNEovxJOVmsoGiqOVQsGaWnNPVAkHXjJM+HaNHf+jev2UivyrkcH90H9r
5ITilCYUmNtY1PajeUJ/8q4TFSD313oIRc2Dib/D+w6iYZ1IfDoEzL+qCid4FPcx
/61HWcmhkJp+2nI1ZJFVUxPOkDNZblaKyO3MN5JG0JiugEbUCpqwa/wnwgKRhelL
QoqUcuaI6GUjl79p2o4NxpvZZ4RZlv7GAr1erY6tmP6MiE/q1FtwQNyyrd0wCEWm
nKTYDu2t4b80lY3evMNsBtOIT8AxkzwW2uHNyjLpqhRs29pjuPqjIyIUZq4Ym0UO
vrF2Er2s45bQilRg0rt9LJhsu47E/iLSXMATZeJpQ2n3SJF7YBdoNfJi0+ZNZAvx
Mortb95tkW/BOgInyTqkFYl4tyMnBLa6uiFC3KjXxzUIAem4HZSPY1zMBNALhq2N
OKuYRpXMr8tZnI42SbmxUWQEapcS9UxxC/N4SprV55au+uxVp2WvG/kWsIFLtsQ+
EVSZ8cFo/konEdp0O2rKfBp/XA6abg7T3W/3QJRsiaE3hGaImkxzcYXTpKu0mzR0
c2L82WwZdBFgoLFtTU5v9a4pXhLxtNG3kedG46gLaBRvbkxj+n0TTLCPfA020Cxg
FlOlsUN+a92u382xGQ9GKjxC2lc/hhG7T/6hH1nmRllgC3h4BroD02az74r/vJ66
Lmh73LFF3I8APAx0R5h4Xl7z985jb9lPmcWZ5d8S1Rr2KjEZalP91u2Wjeop7SaJ
fv9QAW3M3JtmcUEVIQpoR4OuFfM9n5CZDLQOYp10EGi0xY5K9RhXB4i7n9wL8jpa
uhHRtGIocTixA1ziduGHg3i0sV2Xyzy2W5jKX2zPIhc0WMSDeNs2Qvk/+2VXTSiX
aFTyfz37RWjDjLbl8VCmtVWJ1S+egA8/7vhN3FaIqK0Hqyiej0xXaOCw4MQ36fhE
GbDnGPxfRjl8cMB2oaPXk/8bxE7kqghlQ6enWjJnCSwqGFcm5w+x4XgFQp9JZrSB
iQTKFSrPpkEP5BgWluEFIacktwMMojnKZPXCV/FEpDnve3vncPrhRIAteW8+LsQb
vNMcJ3bq7yLZkfReOlw8tg5jRXx++n+DFJg8uZf7ly3Max0hkEnjfaqd+KFEQOhM
tty8UV29yPWL+EdqotuRu944+3qSM8U+ho+2Wl2sBF8MpLRXSDREqH4paGiVvH6b
GJvaGH6Gcsak4qwS19ju4o/M2boBp++rsxjGbNyTTeQS+sd4LXRIIvAMJzQ5jLK7
TP0YRSJcehkCMQVSfkQVbFPhmKsuINP10dWZMKLq3LmZk+RBIHtCmvWiIOPVxsSR
99SoeHeuw5nPi/4LrU+qK4yJXQD8wT86DQTi/q9wPws04MJDRS5+kjFPF4hrvOgv
McCq7uDLrWHLavc4reEwC2pD1DV2r9c7//lH+XrV8/cH3FJ4gja+YTn0RX4enkO7
rqBvjr9DJreX2Gx9AIMS+gdbFQo2Uf1B0R7n5bmsS2ZPLlPa5o8GOnAH/nDfhc4g
MrcxQFLOoBsScVKzj0NtlKgPMeAwO42sU+qTP88bjvKzIFUNEaMAyjSS62i8g+SK
bUGPnXdY9ZlShZFjsqq2I2phv2D0ub/1DeJUP1l+7Scns0VFjRfrnEY3fgWXi6vw
Rqp888whQjHdNdUAUEpQ4I+x51pBxhJ29Jpznofrs9WbrdFK5jfhukVATwFcqTv9
fDnSh0RKdPhFnP2eBCCssS6JJpgIErJ7ztBAB4TBle64htQIi2hJa6qcBnz9m/3z
QM2sS87hr7DgoH0jva2wTmsDn5GYNBkzg3mkPjkYPEWgV4K36e8bYvhHcCBbDA4v
FNv5XNfHumQHmyTgLsuapdWk1O6rdfl6WUCL/B7etlTolyfzg5MZXVRSQ1Qou3da
n09Aqlw0FvU1H9xQjZmR1NV4VhQH1D7/BDiQRMUAIsmgs8Zki3Ginp3N+qbPmAD5
QLUnHGBo/r5FTQgMIh0dyF/pX6zUSi/jHrKt1bYpK2uE9lIlZt+KOMrfA7deYm2t
UihoCS+B2c3taw0JhqPOcnVwVfMn3FqyPghcvJ7GeHghhysnHLtChuq5v5d4QSml
9O9Mb2QJzZPaTb5k/GBWcfR3UoHSzIr8IJTMGl7ApxLjnuRQIXrmE6YAvKGw79LB
vZF1Xv+mKJ5/m5Ysa+QUjOcqSP7X9QjirH9bBGMrLKkefO38jjxm9F4f2TlP9WBs
+OIj1eauCfPr5LsSV6tcUPnj5E8/1+PeVcF0AQUipA4FutLPO42ql4DKZ2mLXzPR
I/wcO/dsVjNS8D9UDurrMCPY3Un+40S8qTAjDTn02N1GFAw7nOWofoKg219qBS25
s6UiW0pSUVC9EJCue7z+YtHWJpYsoT74t960F5v8s555tIcO8seE6f+qV9ulnKKg
LQOd9n8/sTMoNMHsc2nkPA11wJ+5uXs6YiWLS5TPbc1p/HZL2PpsiIVspkwudaK6
ySp8nVTBRT09CdvjSgxHoBRwQfLKQsZ+vuZaYGWlLs+7aCsoqkTClSh7pVsle5nA
86suEd7LScKyOpuDLQYGgvlB97rSFWaEG5gFmNtvwRs4SccsPEILJTdNqhRd+yNH
IjQT1CzwhNEA7oBkkwIifWJItJI5lXiSGGQ0ZIuOcEQE8FkdN94wAbB8lq2lRHAQ
txgrGqdK4WStKTix30VwHrWtYXg99DODqB8b9ddZl/SaBkDZJMp35bGdmxLpw7ZY
6SnJy9vX923qNvzCOjeHMK4G3dAX8CZycoD+bhM9FjWid+tadJi4GJTkP1l9mMbP
jomWCLM4o7Z6DgMpdXqkrbrQS2HlZKWsyk96ATN4yNT8/5aG9b+WI8RlCEDbihmJ
6h0QbClReD/+DJkNxmFDQ12ayynStFatmoaZwfA8x7xreJCkGA3/biqlIm7v/5YO
MmcGyH+vWAv4YliWF0pQ8QPr/yjr+cNJAZNPfVjZih7p0xggyOGvXJb+vIBd0vD6
+vjWp2RL4kzfgvraOoTjFZjQS7VznMCIkD+eANf98j7YejBcKDfyOmFzXL9L7iDv
PKrPLXELgGVy1PsojpwOq2GKm7QfYCqxOl8JElQxzTOyTpnME4g2H4T87cp5XVas
zanxy4owWnq0iTUlHSlOuWTmY5PJpJ9qkPM+iutcLojhNfB3RnHZZCcC7vBkfYDL
DY8qolY+EwvuBRPsD7p59tMjUtob8TleEJvuATUAkyga3u3HYhwJ0c+7dUpXzYCJ
3H4Whg83aKKwK4TX24j4B7t4f9eGplf7n0vTpm+yUJbcGsbvPAKdg6Db54ZexsvT
iOL4c9cHGlLY/I5kQFhbi97jd42Nw23N4BujZzby5mfxT7xtWM2PwJjEwXgeO740
C5TRByn58dM5YPxMzRDWhJUMfmHwg8MuBNJzJBJelh/AUgz3aaVZxoIl07/5RvzS
JvS4OsLnJx/BqGfFPz6+6nld/2tKGUj0YVCLHsa0//YXic9vCbUoEPZ54DZLxrM2
Ywwg05RPO1xykBRhAXz4JApK/20l2neEEqCH+2q+Tzlnr6jktPACgBb+2wSyZ9Wx
n7ZhFEeQevsnJc/0ECRQBJBnYZLzLyTwLy8VJ2pAFvc50lBx76cxkh9IQxr7i3gf
RVonOKIgPKw/e4l7YvrFXl2MLFEVpAxuolclTNzp5fArI8UkQz6s6pJhGxXuOu8b
3FxR2kVxk9Ns1LFj9Plc4g/fFG0L45VM7m8t57r45yXH050GwdSXUsOxRkB1lJfH
WDL5/lPitoxa8NHpkMwuj4MEbyieu24QXIzfUHLJoZx+b0nBelqBA9uGvN6nywfg
vnDUsV6AdqU8YOTSQY+2I7cTLEED3AcTaSWwV6TOM10zRbXBjRm0x1RxIr+NYMza
kxcTm6aA/L+XNoz3q5p3b7R/oQ3lCmzfb6R/FGaYGUeGSbu6Yxmsrg+CdOn+4kq1
9VZgkkzsRsYpCxGpqLk10Nk+B8E5RV+dGZNPfrm+kGfR7hhi16WKfcifTMz0XWGF
G1x+RBIcxZdAYolmEoRRlR2yn6sk3N+epJigbEJYm70Kp/bQ5GBymuz6z6D8zZMS
8v/sBiCCrAu/R1bWQu2N2LkefS/FPl/YPwyiOR3UoYqbAiRtgOMCkbofBW13cbF8
Sl1d3mQbsZAY/lgWCsmj2339YmiNCjlsORY3ryep4UtqMcPaBpGciJIbNqc4pYUU
bbYFCO4q1N9pI2SN2KAzYPuNDk7ff9jWjvvKgpcvlYgygyI/IPqr7rw06XUQpw87
Dg1KV3m3hlmPkegGLhHs9xzGrf9xby/812stwv3Ycljbo7sHuD3mKbyWCKXmLLWy
mlQGUG7q6nFOyg0RODETTB6ZZtSHPbD3BFuChQe9lJp2kgrJKNtY8dTmjHiUcy2Z
x1WsJuE6gvMESLEWSwcva3RB8DXqu2DvN/e6EGHA+w2G3YdDnKabPtWB0SidMFGx
bQ1uAf6klkSEIweY2GsjifxyMmJ0dJLVaztW33LHYWjVYzOAS8y5VrUyUZRUMyX0
j2o/A7I/fHOiCJhdBNc7RiE6KTE4BmxivYoM8ACt3eiNqu26kl38IGcLP/hEBAxu
RC0ahks5Ml4RgzC0RAFSFZhk5Nw9WkIm+4jFKQrJXTR+xeb8lJjSgCJnYaxSq2BF
wVbIoTTdsaSW71/rdQ01UsXuQ+SqSt8MhdvULpYOtjScArWt5GzCgyENOGVJK34m
6D77LiVf2UgcObDpNX16L3Ngjs2/APN7FPQ20KVEgPSbNnqxCHc2mGW8U/+I+IOT
k5hCu9VjNJUFnlv2+r3npVOnykN5UU5jbgO5djMFAXqHf1WdSRCRH+Fa2b4XzRHq
yXNuLp6PsD0GtG84wzIN8YfAqR1PndYm26JHVsylcNEg7VzdhX4pwaBDD6lzxnb5
T6ALoUtNCX5ly2CFbn5uMrQwgy58RdMzOMom9koh7TMjEE4Np4qHQCerRY9DyLu2
mop2/ynjHTrxYjbFMoZQEYU2pbhjVm7CJKR65EQ3bXo2u8hUEf7t3vtqa+n1v7tV
49HuWBY6NQYk+R8AQnfG/s6vcSl62Y4bVPbHbrwUP0jMEe7BNmtSWd9Dl9MRRzpL
XfP/W2htLKcsO6Vk+Y8rN77BLgPKQW3xt2PBG6+d29offk1d0VjbfOTYUWKmWE9Z
WJ9ZZRicejEdOuFxIkTSAWSif8V/N8+Jtlbed6aykqMP1Xipg36tlp6cJ5xzfBjp
AN6nd2gu6Zq2nkcJDABeu1alSDbHriuQqUu5k4Odj1XviyFoT80ES/zy2tw4P5es
Ip1OLyoxRAIHqLliPNu+/o1NBPb+X1N6f8YDvrZggXPqos+hOxFr1c/yrMneocFv
oMa5cp55BwExqX8jg+eixAAVpUgWfacxdPvLz8hEvHiaSL4bR82BGVOHLqnzXYvF
y45tzHZ9AVhNY2cyHGRFEFC6ei4ftIEXdkfe+kHNVkmKMvupOxJFORYvcHLtoDpQ
ExMLXgO3Vpo5mwqHwp7svjQ+LbI/vSq0Er+sBjrZAd/j2VXG7rouekzrxMLI+Jh9
oJ6f7tVrjOvAysg3H2UgVRpnMpsWYmwO/o81zzGoDuItxZgS0r43ApT1KmFYotIG
JNUUHS6ELc1ZfDRQVFosFVLBGdYv65L4z7UlqfCHTBWkuQMpOuwpYpDYMcKgDuo4
/+QH20CbKWTnSWL1xkmCdtyTCHLQNOcSlD1SomyVN0MjwueUY61LxQbW5oc4pQeu
UcmWmn9ZrBpstNdcZ5OZTs6EkBIT5+ObgPsL3wS67vopM50Rd7O3nJHlp7BQYtKk
p/UISU8aE0PQ7unbX2G0jOUx+7lLwK6XQ0tfwxwoecDZ+vsV6n6RGjN7duDzeliD
8Jcc1sviPretRjFxkIU6COv0ENyxJRMqtU2/U4601b26PPTBFyEaFoyYYv+UCvCs
jLpOIvyIApbPpRQ0odFm/Qb3wVeewn9RDOVnIZq6GzmRcTup+8N1fZeeTaWzHOEQ
SWy6O/80SwU8D9ZkuLOjYvM0rEMoyZ2b4Gdr7uNikMq4TljvT+xcFt0pymgw/kG/
XBx+68I9r5ueTHRykK4CsVbzI/fFPYTtOwCLA5pX1+p6Qo+5dHSogDp8+9rlU7Q+
2v2YOEayT0+d28hZn6xkK1XWviWn+MV3hKYYvDbJ5KpUoeKmfU0334sxEgSYIfzf
Y7+JPVHZycFClGGpjkHuIzUmG60THS+cm40UbB2bTfKOhm7zDWFdGKV+k50op5je
zB+AE8d459uAWmwN12FUdpOeP9K5jv7VvPv6isIyzQPuz6zOW91Lf0TLi1k06BGq
vpGlwN+feLgFSmyD/znCZv3f4UVYZ8iD4MeavVslAiyQGEORDIJobz8ROYNf9msU
Gq6EqUzQL1WWp9A/VUJCtKBALlFsaa/zfmpyoZUzuk93KfJhkvhFuDwS1S3o4uvO
qT3v5iA0E7/JaqnTJBYWHkw9ryEijXdKUFs8P649S4sw8idrRYBCYdX9JEZCsHOI
x3H9b78hO/VMy/sWpw2aRvtlPZulsp9mYxXRFwuO7ajO3Z1UrLOuvGDupugEB8H2
lhD0CU/u/M5rRj3G2s5a1oHPU4yxQCdZcyEObEsWuOJ7e6V++EEXNuLeibdGF1SL
XqhEgcp3yhXCI8olieQfgKYmJPpM6eSr1nZne+fXES/WgBq/HNpjDmeIcrLtAoWD
E1gIvr2VLjvW6/J3Ng0rrMVQA/uHwst9dVl8Vf47j0aL/BUnAhUJde4uM/AhpCGx
ZmXdTyHv68hlo7HFyZUmN6MB5ycM3bpSHociwzWnGi74777MVtlbVWMhaG4jYfJU
iqpvfs7+JtbjaQz+/fzVoY8ShQ2v1a97brjWUjeoXCCDB6I9fRGZ5qL1QvWKArKo
en+ZkudIi5Uu5g6tSgPv+RVWzpMA/7VG7X0M9XEnP/AZkmk7vXCe4uBKWNhDwSk5
lfr/cBxt3lS4BKUzuZ267zrvi5f5ZbZTyf/5/i+MIOdnGWk5litdokMI5kjDP1HM
5YTyLcnyzntLYdmePRlHFX0oofoBZtEQ7S7BOcxx5M/qFivJfmrvgTDXfVcE+rUN
KiGcbMaxZcr/2ebGoTdAV7lCmb6gv2fGFWXQzZzG4oOm0pV5ZL04LkBQsPWZwmYb
Y2U2koB3BaQ+4EPJJ0D2zKRYe+LzVFP7k9DocEf+JqrCQZ+hJEQRHj/lD55qppy5
opafo05ivPMJlwH/MGhgPpJ2GkpRe6Q/iRpmWtFKr1gL14eRYdG6M0VF04nCsZZ+
NIfr5+qXgUICf0axFQAwpeY4KNEXvYEM8Dj2P/xYtzgfrScIdBG93J3IXLk4Kb7H
1ETBf+MQYJhDLbMdK2ZhTgitSEIjMUgooghVK0PGk2qDkJCADJFBYEcgL9w4wZwl
3sUMQWpDLO+regIU6c12XQ+YYwILRbofxfiHzmpM15Xt0zBqhTpeiq94XfFmSXkq
ShHA4hXf0DYUbzX2tSwACgisVykeYqEx66dYy0w0lzhIfygkqggfSy/uYO1hXA0Z
cp8d9ek5D80YeIftC3mT5NfQzFNH6ydlW9DEbqk73m5YIgyzNH9UtboH42zSt0zv
U1tRBmoyot1M5fYAbDETinRhT/Tx0TYh77rln9gby1gWTswZlfdm3dVD8glf2bnF
GbZeFtqsDgYraAOjdJEsJDLxUypiD3hj2KkGppXhZEYldV9DfFQC1BUV3yVrHxuD
HZzfWIRVQMw8zberhESNkh5ob++Ry078qRSiAuhy3Hbvq4Mvw7N7wbmD9569rmDe
xt6mAEnn/VPlrBpkKpZgNENvGsGlCpz/9SRFjaJEltksvaJ+9za152/qoTnEx9C0
g95IioSnDjmjaZzmUrlZfPO63dJuZ+b27/0D9l1AP7xK19d++arHpoPJwlQCge8f
LDzYvHCpRt3g1WzM4bo0k++W2DODzNe2fKOjm2iP6dQQOvh9thMXpDJcKWjDEzdO
5PIFbBVHsWF41mmeKX/VMtXl0wWX/+o+pPNWcJpgztsHR211VZhKa8DTBHcppQEF
FPIF/uhFQSInCL+p/mao/4vdNFv2d9n/1PQZGaNmvj5+o8yINoWs017Fc7WtHi5n
OhZynM+KPxdNtoXuKkrb4/kwPGxOwOvZ+TINMXv8I/FPwiek82N//j32R32yTYNY
hWezdWUx3soqEhM/WBlxtj4ETHCHlRMIwBgGhNfkoQw90yfk+ppSuOviCzNIZFzR
SWN5OpgGs65M/0QcIIOQrM2bcgeifrKMRi92XM7518DgTPs9MWV9LQDEI54ibx/T
x0fm23Y8lh9F9g+bYHuPn8Hv76qxTqvLvsTJiutJraOSfnl8EOxH3HtZffdNpmBK
MQmntEkR13hI81LdikomReE/q7EX65C9MkEuNo3InKf3AqTarcj4jKr5x8GXijiJ
uAWbmxdGxEclLB7JXlnln9nH7i+vE4alqC23O/LeLPGrXwe+NDNw3WcTXqM+iWkK
KEXvi2G+vrqui1wsIJ7RYgpUtx7Qqb6gV89mqgz3E/bYmqsWoKFX/thk9X8LZHrO
WqCOm+CjuasWEq73i2fODq62fdGNOySXfK0rAwZK45UgftMgQsV61k50R9szxvLu
qGbxaAQ3cI+KjEXbsuEsPDp7QDmQTznOxwI+01jmVzlq8q9FI672swAUXZNMa4ax
JoWuTfkzjL8VZCGK1sVv0tpzMyH+LwogTaqrzQJ03PDho2Ae30qA2/Pza3tm5Z/h
Ee+6cGlXtUMNiL9FybawMTGY9WVOueOKlULU3clVohXUMywH8am0UOxTZZh35xiE
Q6CcytMjDor48uB6ziLq4HKeB2mr1mV7T4Iu6+PkgneTxxrofTdTJ3qoovFdE4IY
lD9UV9LX6SWMiGwpvuL48lgmNORWxpcka+5Im9Fm3IQg5lvVrlw6NTt/4AH56bCs
6giHjaZiXLg0vfnq1A6NtB1sW/FQjXV79M+UexYozO15OapzR0woWADlji+ADqOP
dCzClbVrx/RzzZSnu09MmAO3dDYxfTxcjPDrfeIsoBskvkMoMCUEpPd5hekxdrzg
4RPogrTG+EBrYVBeVmzuBVr1JcX3ckXvZzU7pYWzcR/sv2mkACZfGdgtw0T65gP5
PCubM57CPAA8mVVQEbzf9E4B2kOxE744Cl90Zh7qJ30Urcg4Y7tjpKS0Lwf8ol7c
Q1F/b1w9hvftdltR/Z9xLOg5BzKGkDwjzMPqwkFHJ28biaSAZFIsiKRza3QrNNGU
Zl6ITJ3bhwzWjPJTU7PnJzoA3pd1WKe2rT7+0kfBD+0gPlpxpzvP2ERw3YvNJoR1
ZeoI5YaXFSkLeq8QvtCkhVmYU5YsRS2XX8aV8RAvgRTI8TqGQjuetlICG32b43/+
QX/LI3aeQA+OOazzVCKU7NV+Xto9QckqSorVcvIiS4d0w7XJ1TuFWLRcvt0cCTX+
UJBjHZ4vKQCU3zKqclsLN7F9rSXSrhiuyd3z5qDm9001wi73vzP+KIlyZ9HdjvVH
pWwsWiVDy9c7UUhQi1AtKH6umhB6NAUmSuLi5Krvcu/Ek4TIG2iBhzoa2OA9V28h
5KgGCOFFHRG5duMnXk/I79djZTSyR2PxNknhhHFnuCPE0kOQOReP69V7gq72MHjJ
IiIiOp/pVUbcuwOtJ21C9j3ZQ+R38b5xit/j+R4Yul1wW6xdBQQ9SpCSYeO9F1Dx
caWQD4UZeqOX5pNHiniTe0T0BuJOCS9wpHcB4808pCKP38/Ax2NK5MvHivCc0euG
RJ0jXnuUjlY2NGXXVBYmJvD5KnuVyWe2QORaSmOv0c93yF7lSPRohz+HzgoSHnCv
8aCa/CBBkxXM7VTTIA6JsMjVsHcccAxaEt7ae3e4bY4vDvkgPwKuK8DjzV1X5sv6
FZDP2FpXfGPP4cLdwL8EYpwlfiLFW3bFYOcooozfR2laZFMzkgsUbos1x8JJaJhU
oWnj4vFDTZMG8dssfOdw3CYr03oAgv/hUQYIgkCLZqdvyDPbGm0pmMhwyIfk0qg8
zzk3z0jc0eu42ptbkoDr4mRGFR44hnzZMgqvPll4A85YtWVOj4iGNPQUkOAdKCeG
Vktj/9/OmBTWdlWCRC2hedxiWeZocvTjoQByYz0kwx4yrHgvxQEz6/aMQuuZpxZF
SC9bv7FwRLhJvqvfoRap0Wn2B5Kycxj2OAV0hGWftZ8UBpAS467xzaPBfkZS8DGi
MQEuCUrVCHnyketTeQG/jYFNUfBR7YECipRkNSSnhUJFZKroZ4AclRCfM1cGgW42
++ovdhxzxDFcqQPvi3R1aoYp049T9kphylTog1QTvKS2+JWG5rii7g/TsEPa9UXb
HT5KkztNovXvDZxQZIKLgpW8O9oWhENWOVn7WQQRytz4an/1tstgqLGartOvKE4i
+pQu4NY9bvTgwe1C8Hkx43JxftQM1YplKjW6+Ohe5Sx6NZ3iGuSe1QPcCztJGjsX
whyG4gdhLmHUIapUQdN0ljX2GR5YL/J6kyKZqV0qqECPfUsKIVf386BBCL/gWa5G
RijW3YKzqcYlKTdyIiGT3ByQSYmUPMAbOnBPHMHcntgAOFjD7Xfs29CDJ3iAaXUY
KiDdK+8QalPJJFoy4qrKQ7Gu+zflxJqrM8wKN9K3NDJoyrgBvqzrcHtqsBqnTF2S
Ds4tUt7p/W9sFo9p/3Zyg6AcHewNtsoI49fTsCl5KGSRkOx6gGho8R+ihGX9Q+m5
RyuMjqiRGYnFPmbCLTYtO3vBhKUXjLR22sgrA0+1NTRaAHTJAQ6rjYKMH6Rdlo0k
DL8Mk+oLOQZEIhmLMShIie0knWNZcsZ1Rtmh8o5Nh9UwkjqBfkZjYpH07pNFHLpr
gX8DkxlsxPO3rO4ZimQgWkQNmPP/CjGZljNzHW8SSUNf7UPgGvMaYvbDfhksTNXY
9rDJfuZdx/ceR/MLCzdm8L4b0GoSiBwcWkwkKCT5XZWwxyLk5t805YesWGGY3x5i
0fI9/kY7YPZXbWYSWShF7i7ROjqZv99LT8wWv2EKKo3jS3yuIRmL6pUBlT+JQ3PM
dgYWW9fzlWSQVdumO4Nmjgw2/zl8XPIuHySooNE0UutTPCoiZgSfURm1lswi2Umf
qhPohdEPd37woptgzurGKmmMFIltolvURb4USRYgYJmeWyl8P3k+bxr5dn6wLWfJ
MMkULp/IUdouJJu+lwlNCRf3d1Wrc4SfC5YQq4MMVxpXSgNB78azCYuZtDVyPSJW
b8CAHUY14ODIyEn0yfbrOhBA9Opob8CpGkD1sLSdcERbDPKoAwBMyGGlyA4QPH3A
4nW15kSvINox8rUAERiQ1Lzw1JmAgIfLT8GZABUy8lpJ9eNgWZMrUj9xTEMDQi8s
BvTMRNA914XqcasFB2h/CCHqMumBtzy2IrDmt2BS/qBWDsW6WoOCHFUveGc8qE2v
olo3n+iQtXpVMYvuClO0hEpfTcMwGlSne+FgjFtyFJJ29T6KAdj59YOCYxipCLeX
5b9c2T+RxxwOxyFw1GQ1hSUZU5w5C9sZ9ZeH5SBR2EH87RJ5XGHDrwzJyHtGiOaA
OFn2UhCchB6V/vCybpv1yKUmsGVak/NEt7JRe6RbsrCcQ9Xffg8lr3JTAjbyvcI0
J77Mqv0aMtOc8bMQKQipkX/4bi2gOv5IYND2YWNMvB+G/CcKy0sbLaadBsO7CtoU
eVHbDxYkZs5Zw7dREIYGQAK3ltVWePeg3ksbKk214qCBQ/32X+BswJAeJJEcp95S
rPik/sGGIr+f/Sg2hPUzq2QzeTAD/RiFO41xpykZ7qWepxJY7JvuuQ6gJt1Z0yLY
AbxyyAvkmBZ8+Ji1aDZIxc2Js9c95LQk2ZbgJ9I2h22DqOowti7kZol/gUx/Z8IS
sycUdU9boeX3cvuepOdxyB86f8598dcbxPzIf96rFaDpw3t86oZ1de1LnU/Ia1bZ
hjEzTiw0MlxkePzFtv7TVfHs3eNMdKgjaXw7G91YnLv7SDkJk05Iyy7rR+V9QQ/n
6CF8f3kSqOoVwkj+VN/EuR+MgIa/f0i22waOfh5BJofdNSPgCNUS4wlAtP6mE/te
3BJbaP1WVrclRGy2OatA5ndY1ea7KEU5uRCQe1FzxtTz9Ac6REBWJMlabzMMtGAf
9JbWP3i6wPEDoUpXSD/IzQ8ZF/kf01kdFt+l8gJq/rDYTubdsz+ZnLh4C13Zz0k0
1zxNcsGn/hTrkd7viaRM3HDXbzRR8MFqBqmcRD4knax8UsGsSlXpGXhXFI2u7mAy
JBjfL/CHe0fcVgMVzpVEEKHcZNcDBba9FROGRK/kASPGRXnePkfKJDpxz+1zKdyJ
M6B/MXsogRoQ7u8OsqkprDnxWeVpTIEYgBYKFSt6Sbmu3UJMWhcAmkQXjlg6KBNs
7g2pMzx3/Q8tWpUUiRDJrGPqaQv66qSz/B7JC5p7sNRBpZmWFAPEXIE+F/MdPe7s
8AGK8/iYB8ZcgGBivTLFj9TyqM9Uw7FSwZ4Q2FsILajV8Pp1qjFKCeCvahgxYhh9
OllRmDIlfMzrdFka5Bxh6nOmogO+mph68w120opX5/1g+11PvWkmU6meb3Vt44A/
7xW1eBI1CDkoCS0wdsJSfshezz8nYHHry6GIpBp4zjCJeIWxltWgDfS2C274c8Xo
ZS4ZCQBd2ktDaI3y4CihB4yhWB1PyuVZSz733pAGsGrOtVv73wuv54UHAQmEoL5o
yXJz3F4o8y3VaT7JriAdjuPdm2Kjqe7LKtY1pFutuFAGZSctLlMAG0pcMQNnV0y8
fYpBPXjW5l4Ql7CpfGqTEKZgPUItGmPJ1aEd450ZbFnmqnsaxQGKWcvTBZNrYLCw
sx2o8wkjQF3aTdf+DFWB/a8AyAUI6Jqr/oWGtYV75dCmL1nyhqZSXSWLdX9F76UU
GVAQMBntjLlUUf3be0s/42ETk/+HdCFuL1gOBDqavqIQnb0TWosIsryH1eL3AT5D
zJXCI/25vBhmRQnuUabbDhXL2G/VApcNEvM/CIWk5joZIuKTVXT9fnS87V8zYLVJ
fKS6T2VVLihAvdh3JUuA3xU1x/II+hhEtQVU6YtvO1L5zPisSNIW3Nil+PfN+HSt
i9UgW7AWF9J32uiYXU9Uo7pfUjb/8mGoWbH1ASQK67ZOj3upwEp5Rr6TVnox6Csl
M4NKbv3epYTrYWDTK20YTmiGAd/zveAjsLyratWzKU8nERVRd1pn256KT6dXZmFV
wda7v8YKozmGJIWQAZBRl4qIZ6ZWIyxMuq1uTPEUa1cMiSpNZfItK1RZLWc+cy1o
Q/62HlfUzrt8Crew8ZXxpNUPP/duhYK9+XmmzE2214EgzZsVkCpzvM9QTkX8skU3
haqYPQQROekwcMtCZIiGsulBdxZKp/ye27O9E2LM8fHBv2B74l9p37TqXZHfoleq
IqFfBl11YKQvFLboee0j7yW6epjGYK3+KuB0RQzt6G0MdSH+gT+4NIM87SXY2vCi
ys37EZsGYdr11IFVncGLMRdIlyQcEPw3YbD2krYDYlJhiXkiPjfJo0KVh73dFZRF
3fgHZFT7taTb8TMrToWqIIy+wSAL/PW8u14naUtamwv7SV3GatJxnDNuzZtnMIhA
o+VK0bN3znwpFKBsTx7wR98+uRnK5GPWr8d0Dp1u1Gia1xK6vfW/cTOgdjKVTnm5
68rxwEcIDKZSInplSNZuDm/4C7NmVO68FWFeKMEBWScsvKTxYWjd1oMaTqlmVMhA
BqhzsPB/oJZH/vgkNIgS6ag3L6Vgpifrvl/YPBrIX6X4vWfcl2qT1ext/OZtVOXT
VBOIIqWE1/dm006DUg7M0c2n9Zo9WuEmhgJuNlgaXIHZeZd2frTFKFN31AqmKvQF
bpy1eP5ENG7MDGbEX6GIrjVLk0dCFH9091cD/phfFUMJoI8apss3iWsw2Op/t6+G
G7/G7r2CxL6NgWWGNtK+2oSOIuM40DvfMfH9oFBCKFc6dNqsp7bLSZdlLpkchQNf
DmaTnKLIoz+XnRJv9YthZxhzXmS8QlITxL8cYzxJBTfPxh9JeWrkYjyYz8ie4XkK
mK9JLNkAWwcs97JROeWfV23FsHSl1O34yxdeXq/3GPVECq856SMPcEoX2lJXI7jP
US9OWD1Ez725Hnn6sPRr0hjuK3/SZ+ztkJwGz77mcO3iKsWofujempgsCfOXpvk6
5tykOyCHsrRUgnyHiI/EVOpfg51oQAcwgTOCZYES4mV7DgW7yia6v8iaxJits77r
8g2GWReWgUPKldlXKLazQ14V7ljQka3xrlzQa/2m75S5LVnQ+j6AuQL1ijhhf63c
Z23R81d8MIhcEd+7X3TBbTDCF+txmaD/DWm6nqgc4JW/M1H0xWWI1dD1bzF+eorm
v3WXGoYVSAHQbktsTtxP9+1h8gZ1ZdOy98oeLEi6QqxG0yIGd3z/YWwY6RBnwkBF
eVii9Yss7zfuFEMJqyBpDveIx/F4EOH7UpkoRM1yLzBtHxFvIEpEIaZOoHLgUJ+u
auUcJmreI+PrjQ+WC/wpLRapifSv3Rf8lOq8k7BNIVsO9Ow4m1w5i3PQ1Wq5ToaI
3oREHcoV5UEcjyAjy7qNtx2YzOpXowhsmfzbGCYyYwMzdKPPF7reJP23ymFc1Trd
OwTabK4rig13chLIr44bqX4Y9GFCbNtfHdsgoxv6qPA6TdSFs2ZUYH5uLiFPQh4w
vAS7xXXxP1NO+UpSx6D3BW4eySyOudCjA3kZZMd7qt76juX2xUaMfVM77Qos3JY+
/H6YHs8xUGSU2pxBC3tnllWvSZZth0Tp8+5d+T6WRSCP2TXxIUKqE+PmJWhqw/mn
j6CDOW5AC8q0WhISmwoFgN3kDJv6TOTe8csWnqFoa1Ves3kLkf7Y1WZG8idHGTgV
DT0/ajEscgN0OAPMHH3yR4TSqe7M8H/CvszwUG/loF/PjP+P4MKpKjHNdHJ3H9RV
+tOYvfyEmfXRKZiuQ9+nOlvHhVRH3nut6L8YagzR1ixZTkGAxfLru+e/KOsVawrO
XcyFRlPF/46y6qth+POqntt0fTkgCTLktXflFAXqkCZWjXGQIquC+pwNngZikV39
UQWL/sGqWtlNyqPL42IUD8mfjVA8e3w0goat29k7kgfhJJH8MXaj92uAyz3r0Qjz
ZHLV7y/TY7FuiERVs7SUKSgP9HrIJotdfpsu6iIHkZGOYNhg9pCiFK+RWVOQpNom
7bs4JdKfHHCoaTUQpO8mVPF8Q35dWPaHn6UUt9BZ81Eq8l3iEe6h+dDG/ptdW+wE
zI61uQ2zRD/GJlwHGpkkNVba+hGD0BOmzm56dsQngc7PGWGBiSql6EiXQ3Is08aF
jpz15dJddI276VXa/kBIroHKLmJqywI0i7dv0XGtmvBEa0Ok0Oi1r5rm9PyG79sQ
ondqgw3Zz5ir6cL5RmsrpbGGuwbInwijxw71U92rzABwc/0dALVwZnGcoAhdIlFI
NuKwkwfynq58DpcNqjWBRGRjCFBJj9m+5s0ef+ROoIIImEqd8VjyztfzrdYdriUB
ScM1f7b+PbS0vfMfaotvgBduuSkE3WMfNENUbi1rZqfG/wP+CR6zg916t0BJnPiX
glOJQptKr7OziEFUQd27Od3mVIBygtAtywxMPR1DOy06/mnELDWLqotlwMSa/1nP
DuWi0yn4QSLbZ8uvF3TC1m72AJFmcp0YXjps9iy+K4rZg76SjRoNc9OnVNDX/CwS
GWyR9kT6WswHmHAyMsV7bQdBrsowaQsZjIUh3adBEQw6rmz2BqAaEM7n1U/6cN+v
719pHKSUhvBWs0WwRzEhNwqy4WG0FcmRMAKsEzjKqyafPW9jksO5CfYmszLUWSLk
mdm7GWBqBaOl9nyJWzDiki4kMJFuLN2K3UPtHWhV1FkCw2q94kfvwXRYBusMtzsM
plL/BaG2DTEFyixEZm0fK6NlNhAffTjjVZnCduyEtrhpfgUpH3HvV4pgaVB6mrYb
N1kQYcnirptw+i/Y5IhjSn11Wft+Ix3iPvOdWiHNuqltS0TTkdAPGrSC1wQnu/NI
s0eC+zintrrg2c7Dg4tikgO1g4v/G/1k7kcMZJKlDUtm6BzJ8gcUK/2mH4xSMdjK
bKYP//yTfplCMKniNlwIi5zaKQBG5cx37pUo9edHLKYYuIz7jL7kzXsdQKZEBSu+
bkThAreX/NTqaoCoTQVDYxskutwxGdSph/U2gTE5Bg/yPwyg/ddVM/ZS7D+qjRdJ
kiv59hb0v+NDk1+wKG6KSgtqxMzefzVE0zJ20iS5wQllRQQ+RxZ6pR/UF1DQmvdO
dYqncSvinToNFJq7MrWldQq3u61rAYhi+CXYnNd+bxLs9ITuZytaXXFzKI9MZjWy
nAbexGmtruulMPDDPLU9mlUCMAppvPXnOYHYFfnOIK7hFSIzqrZw7LVy3fUx+P/v
CiEF0kgBvfopDQD63qfOh9pihEIzXe0qvR+X3V1aTYVI0PAdtbMSZoQZuHvIVRu2
YmzB/ibF7pVmS6EaqGmxEiXxCNWvlFhkKUfv9ZRv6EUjTaFBX8YVb34NEdAZV/1S
OBM3fkMJa07U+X67IwmcxF08SP+2OYj2uvzVJxv0PYGIhVhDM/8KqOyQpR9XY5wz
pAbksBHiZLqSgaSBxkJpBZyJq139jHP6yxwOnp4IUA7f4TiPi61k+PG12QgnKcsJ
FZGma5Md6ppMekOo8urSqd1TN7bED09b8Dr4VbQdw/sC4pDtif/ZGzpdY3d5d2Z5
9/sFmrK3tpHp79HvXR69B/TWQxcU3AYcUNLNhgQDH/31UA/g6LpoCtHO1F8p+BGA
v3g8HK95BgMKl8oJTiNYN1/qqUTNaXO3yfbcZgmQhRwIlNKsSfuaznazCVHetPWW
cbfhAVwOMJhkVqoTVPuec13eBR0Xvki2kPg9M9RDSJpjBi4//anC7nZ7WDeBWjdH
jSlHzajkpc+evWmJ1XooVX+i13SKiErKemmhv5QPgM8IypqkeUIepvB03iz8q4Xd
aJlUXhjArcVL7pxusvT1MnsXrxpWU3b/oK7FbxClUf3aNDx0pF8ySmGmg99KpAV7
zmuX9UnekXR8/GmFrleYYd4s68gUTv45uZ5iLuZzYIh8PEaktRrGF2pq43S0dmOR
1HiTzqxZwbDnLp+nQ27jD6EEl5+ysFO+j1AtpLqYhiRqERw3Quvbb4BL+9y+Dgt6
en+0Y5VQagUwnH5UHN401b4hJW0o5WeRYcdStc0hObLqmpab4dsME718wx5Q3kKf
YYB2JsUxMFIYK/Y+7luhJjEhrIkcFM3lpHZZNuntSR1KM3bNoG7tbHGsrqiC017N
zga3mS3u8JR6bYA6TagahW06j2m6UZmCxZUa7MsT/idpCfP9IhgR5BiM9ZPU9Nv6
jCrjJwQYXu97RMPbNFneIqNZlBFk7wjSP8UpfzRct/KOrXzpeFCeQeKXx2e3aqMI
Fve34T0kycOBX70VPfJvqG6TAbPzrZNzuxeMhByT00lR7YpK8IEyldlUH0csIkZQ
tJOlOjxxRpLG4AYBD7FRQt1jxYcZlIeRRTEfYJynsLgwIXC+/IYcBRjid6+f5/Ym
0KWl7PshR2zAtVQa0D3iR4uNh82O+Z/X+jU5OJgtn38baMXnlVpUWUcp7mPW3G+v
nINKyvl4+/fRujSD0U4RURaAq6i9j1Bxv0LZ+asfVkGAZLYYXlfqXpupTDPq+zSD
InN5bPq4dtS21+yMn98l9Usbbe64fFYzfiPW5KCJI/qzLgdMv2//yIbbLFaDxfpp
eWP8/t8OhXb4OirjyYDbkrrfy/zsmDtKlPSORsahHJORvEe2ihBAm9qkv8/1P+gl
Y+UrmoceIrHuzpEw6JHRe7kYMKourh/9bElZqsawQPy4D2u5K2go0pq7XCVnw0ND
Y6Tyky+q0TfZnusFD6xgBEm2N2QFoAyaST7bBCdAgklGV6ltRy98ubnJbogCOyc4
0ShpnR7fuyke7KtGGLLHewfKXFpIVw2XDWTA2eQLnCin0Pb94b+cnn4tcfmS9/Cd
ETg2ZuhaZ9N4F1GvdMsasjMb+GRIJPOsE+g0EOkFItiBUF+Av8Z4ECX7MEvrytXD
gS+1GTR5q07ZGOqevVvPkddI6ikTwApPlkz9GVE7NUShTWqay7DowhwShnQciT5W
arVLosbMTaBLBTUT4Pw8UeQOxdUAqxCgUB9VUIR98gQwDXEHPgk2aqwCkkPrv73X
yvbGvcBbuPvfDnqJvy5RC7VniBLjdYNROr3kAinTUqLMXXf1KiTqUhnVU4ZZs3hH
iEZi/fVFpfifvndJVTvpFmZTJCsKxY0X+poigegnerU1yAooW6Plh3RukI56uPY/
1RwwVL92oan56TZmtRSdwLcFY6qG1YiPUZYHyFXucFv40wDGT9p+jL9e6jHoBhfS
7+vqXkxNa2qtfO06Hp4Z0VYYyriv+axPBK3cIhvRy4n5USgwDGVoyH89aBep/Jbs
9nY2kLdNWx6tQWppdCUzb/aYQi06KQ7VHQKU70y5R4PlM8LzXzJPdnyQEAFj3fus
r9PyunZIE1VPpiMs5LiYu6F1SYjVXQuXK0afjf1NoIO3rnxTdPCVFfTwYcC2AH7u
Kmu+TjCNup5As1QTEjPyamjDUI9593BQEer2l56UTC0wZdufisywaUP4r8tFQG8w
3RhymXSvyx60ndDBRzndHzTWVrs7akfftov+wlkWpOUlYc+AKVMG3LkEJRs59QVN
mAQOI5/+wNtSYbJfIiSxCPkDLsJx5FZKQ7YWBcKlST2Spnr0FbdsQX7jaaapEBp7
CQuBFrQT1dRifdSdPjVF9mi9pDEOLxQTSKOUy3UNJaJ6SbM0adbCL3tPwlqcFOL8
ztlXAlgo9mXHxj2uwhvuS8gUi4M1Fx1abRD9ZnmtCwngou4B0Jn9OqPQ87GjGEgd
2xgPQUTweu3WS9K0U/oEcLWsSgKw2QJjmiCOY5af2bsdw6hxaX+l/UUyf6mRHzOR
kJp3ypbQzse41jRaTtmPEdkwNYKyMggKgrQcVyMaqRz+DxavvHyxKo2ITvDrQFdd
TmjQziBWbASu7hFbvXUO1WuX+veFaBOKArorD4bQOeBC8H3JZ+DeZXZbsJ8RKRcy
VLm+sxU679875kBqBFlufUEZdTYyQVVJV6H6ZBrGOIQyV5qKfHuofzXe25fhhvYK
6DhlWfvDHOOXdfDVR9cM+URXmuO8d7e62RLKAQbncH1DTzcreH7MlFxqHzIzFa3f
PpiBoiAKIoi6UOfJJ2C9ZwaGsfKJAm8F0GyLtempM1e0lm0sq90UeHq89q0v7irU
7HvGQ9GdlLx8c1mfiNwzkoCIdVGq3b6QaHWWdyP1V1B1BT9rLFGgKcvIi1vF+qRH
WkCQ7OrBqzIfH/6D8y0G1J17KL8a9szJZ/LZExGb7COZwBmS8bMULhCUTLrcejMR
KNq++yG6g9GgEC+LDPakVi8joaAHkQNRqysIyB3LgcjubUGbVdWq2ANgd0H2v/Os
UOZyl4sauueFYSBb9g8iOf3DBMoQO7DNjV2oUT/+rBRvyfMljkhI+g55qyU6VJuO
gHBqyq577Hg5cuMgJF68aZL1y3INn4bXapSigTcj86NtvUZaxr1I5OLgtbPbDM8q
dxyXq1fQA7HOFmX8WN1p8vJ3FB2hyYz1Dn64QI9E4DDHX1SkqbvAd9DP+3kIke84
3iwM4958uKtpoub10a8o85Yv7jRZBVYcu1sc+NxMB+13WGpQjVW6JtXrmVpjZXBn
y99x+9QCItmK9UIEV6qfQzeRt8D0iHkVQWxNPe42KOaw1QADgnX6PK+ZaXAihQGw
Cclk6xceo0W3efnmVpzBS7eRjHFUr3aEikNXKFk0/FpQmwZ/2Kb0AGag90j3OZ0y
Im4WWicx+3d76mj0awQVOkI5dxmfJ4eCqvJT9fo/4SUCmPaRUeoNdd55CN6bnjvj
Ml7Xsk47cjagNFbD7temo7H/0d/R8UMk8jpPSe00w12GDxC6MWZNu0aBN5xJaNQP
x95nLoEpL7vH4SlOuD3M+uK2Ek9zCIwoeL6qr5OyHmARHcVPrBEGAVlH7x51H1Li
QnJpZ6ABDpptPxCWWNmVsjyJObA9sB5nEZkrAAM0eSUZjMhh08NuH2o/U/krtyAd
1lmmBgnb5iTrOPHyOMvAjX55hQdDrX2zZZLFk2wAyQJxQi59plBhG2MPTJXAhttf
0mO/QwMVVCNw5WduJEUXFLIvjvQRp4cfZRRbxTrfiHN89xtcTQrDwyjn9NOGqZFH
HB8WtoLqc7Gy+Fi3I6CjLZWhfpjnvZYRYW8TVpS6ZoE1GJYm6QBRZR6kKt6NqXYq
HzFt5m76ztndOEUkSiYz/yvbnmVS2itaEWrEDHIRu+YoBFXVtnrrgTHjbAI3H+Fv
AGResE8CXBNo1zVyDiaarU7nEC3cU+hMR4Z3dDu1SqD+/nuEgj88HfeQd6eTqy1S
nAxZKc6MAQFh1DhgjzsXzk4SX8lhJHIKxUE2XbhcRjhgF9XVAo2RtkJ7td5g7DIV
JtnAGyLoFlPK/WB87Fw2z2D9l8W41Xw9rVbWk30athRSawVplnaVCRREOTozx37O
WPvc4KFbQcZbrIdHYkjva4ijquEm8GQ+WtIbGE9qQ/PF2PyqjStx159sELSNifsg
vho7kusWmolJgds92IdjytmeQYzZp/RmyMZCYzR4ylvT5vaVPS/oLtR4K/YJN0VU
+F8GzPfdSW36k/c7fFG3v7+7ZxIHABeREONNYSUxosoSpbwcsYhtIjur6U2HmbN8
rNFQKY9tItvH2IO7j4WbCBnLGyUhY0EUQziJYg/76BoahXs3Qlg3iMpuCSI+tMuR
wW2ozAgmJJxkfaAgRprLtpmqxSDiFSP0+OX5H1eLh0is5qMe8FJ1A7zCXr6+kcy3
4Q0oRp91OTOq7BXrTq4gQCXvzpZTJLAsYE0Z5C1scEtgv3CgCY0yBgpNukyIVkWs
ZEJAFLBtKzCkGVHfk8Y3MVnXx9JhCbDr7AzQnr7MNvYuvYCileJfdvd3AglvuGQM
CxXiCRz10qJzWWWrUda6b7H+JymYZwer/eteXDhaSidGqBJ90BO7jMr2B5A27lwm
0cs+Ad9KjHyVtmzK7lFjMsfCVghIDdsomA+ZvzjV40vu4CBri0Hs4iZgx/dmNqKo
0WG/Tz+OptZ+Hg53+7Lu+uJdiIcPommvTZSFT2Zcrj+0Wtr3ZU98zj0lSmZT7Q8u
TpeAlARx4GM0hd6meQozlSETtyBiix1g+SIJp748m+5Qy5Cqzp1+hB7eQhV+3Nga
AGkm3SSg+O+zcT0HM1UbglSIijPya7a5tzIFnMTslGwZixjG8J2L26Gzhi3LnYxQ
kiyt71zUIRhdSeyF3tV94i4vfj+CyGsoJpTzf6RjP81TXgDEvv4RE9XmpC4Kl9tV
/h8kCRclg9uFqx6zLWADTBUV3wAg8ELLR/MnpRY2a6tf7v0Mlqlb2lE3REmfKL/h
ZwVL955f2zcrAizY9Spo9T5q50clGrh7a+2+Bok7w5Nrp75zRlibjBHZ2iFOPXxy
iQTjb5Gzhg0ydT7i6BhOHI103a8TcwdiiqiqTUmoXzxD4ty2Hv5byRSb/D8NvxRM
VNxWCnVf77Iq4NvdzJfCSCD62gSE20KnPb+UQsyfIRojuwdp7XjGoKIQzGG+p/eN
tFFnxp1X1+F2oGPvshg5rtmO6qQg4FScjeXRBLDWaFjaE1xkNKDw3FPKiRhGr8hs
stjktvrScZOcI0P78dJOCNX20vRHqoZQEe1tVwPU+OHvvxHB5n5Ck2uRVnOF0xR3
a9IgjcHwZjbLkrL4uh7dRqx+vikwyTrd8dyCXYV+RVwKFhPFOhq6T/lNtxif0VUJ
45a3EbvyDY+MWfXcmNBFeZXu/MLNUU4lfexoHrmIIwQDB+meZr/YEbEfG/dzaQef
1YZUMaehaWVh8ux91uEj7gqlfC3W75OJeQFQld0RYTTo4X8npr7n9Wz43UyQI+my
9LcU8nyRtxkj19q+if46LbqLFjXCg0mnnHfEGFS45vGnkHqHoOAjXs9gKKeOHjUg
2URmBmCEavkJXwe91pmu7MGI023z3yHKkdGojRUjzgV8BklqkD+S5Xzf/mx84wvJ
CkLQuac4Ua6xY6fUlJzF6BrN8UAu27H3nwODVNi0+3HVCru/ZcZZpWS10F5euOF3
maGtFL4qBjvMbkIh4rUl9pZwxTvdJs8gbo4PsWAyrvCYjFZNDcFDLj/m9I21oWp9
Dyr6pF7V54BB4Uzd1E5/AdcdK7d7mmCyfAwzU+FVQMJmcmTxqgYNipfotLExXHAc
1w9IMX1i47PWvtvylPw+wqfhN9Q2/8BooNYM6YyVqeDDrRReINZbMMPgB58Za8sU
2rJtRphTMGVScHIDKmajv2XlJDoriqT4YZoWZpoPTIO2KgVk/kJ9FjmpXRdrxFnb
ZvjKm2r0OFuuG4sPhfup/NwMl81pvdar/XDXyDm5O7lZwz2Xh4I60+XljIFlCqLv
1Yxb1d30rwaL0pykNuQra1ezF5ahlTjerfyON/igwk1pAs+Lro/6WbynZrKUMiE1
/hSOdvbPiRbIXb2w+scjWV8xzTQdFLnYnGoUDLb8C2p6dTSzvThmVU3JwcUP8hVo
CT2yrRO+Mnj/UGn3L9taSo+eJPzwnzfwNcw95IK86sVWXnEqGfxVbWW73kni3s0b
VO4kJekV9e4MiQwtBfm4gCgpGXlrgnvpW+hCYjdbCfrxC6XJDLBS5fdRt62pE43a
13isZgEIBBgZCIgRR5/NuKevsewAqGcQ6QrnkynrRj6L2NJYrlFM+cDfGDUN5Kwi
vla7sZoMtvvRU2RAaUvkqt51Cac5kQO0Pl/sVvLv7HrYRaEZZnHemrP7+reNoTOt
7UF/B80Wsl3uHizA/VoqjshgjK7HhOXK0ymBqahc/ymAsw3C+T299lb3dBrAlAJF
/PRRH1wIpwqQ/yAXRujG7rVhikJao7R8EeOgjKTyc/H/ntRpNRr31vYQxMAz5yEG
cglLc4tVTBSTYc8bcxOlrSl7woYuGXjlkRXIIKaCqrvq3D5MerGy1E3XwG0Ixdl0
EQxMiHj0EahQRoUlAbVpvpWvg1ixcTizzBjUyO0Ad+ZoN0K4j5kr8NhfY6Ft7M/j
BTygzqYu+vIwMMpHCw5YGvhaCzuzaVG7SDi1oSPHSzLw037GUKX+aBFSvjCXCh+X
Ek9U2NPcoK7QKZzJTykMYAiIbSQCPBgI8Gy+cQPjTj8GGifBcIogyWWVsGiEJZ8C
uKNiKzUJaqrj2quAojgNO8PlyLSYCNPlmsLeEmQVH2dd4vkIYRIuIovJOpStZsiX
jCLvHEOxUy9UoFcEedp8d2lTa+YwFw7MDgIzTcEf0a3jazoIFM5YzPT5gdytyi3D
6C7KgRZX/sNQnWIQBq3xGXIsNX68B+EPa+jm+p8qExRrp0hXQlXDyS6t0judK3fH
D3vBqy7axkPQNYYVXYk4Rqq+f9L2AH05I38fF+HSz4kD5jP3oqmv2PX8ygwrkElC
UuvpCJX7m/N+/jeJ0tP1hW0jIRZHYEjwvmfYeRD6xP3Xyn04zlQZup/3z8rqKvWl
f9njF6D9f5FNbP00KJWwgZ/N6Bq+E63/Wl01Q1BaOOcIaOUmQX5XjWTtsfSDj/MC
Rt9kfb2ZleQPGxDbp9xHSo3HZZ/i2dyVl+TU8loXRexdFAIyqaTP3nZRBSnnKbcS
aZZ0Iibzhnlt7UWx6Zyx80J7xBuz/HvXyGkzNxZoorHFSokMNVBOlfxlGuSppTrJ
22vRuokb6XLGMa+TJ5g5OE2YTveREf81ix9/TUJFcz/tA62mOcOomA/Eg2qxuaWs
2X3EBKpHCofxfALSRlXOgsxSQUFCQubCkTVFumC3/1jKEPVrwd278Xp8Nvd6BGBM
F+LTPdSvUcY1r4OF/OM82GOZ1fLRUuZl3gQDh9z4vX/WIFenyv8Kpy5RUgqhrF4q
8MWGT8RX6m44rKtCn6zwR9w6DeXFnaLrFc2CXxGtZEBuXoNq9EEjdXGEqKgxkq5E
hj49yL8QA+mLSVemWMq6m5cDQqBlJ4gb18eOPa+s3UFFGS3DmelIEtcpcIQ+Qmg/
qasOX0t4VH7A9WpZZOE0BkkIbF7XJxWqlCiygA0wk6qpETHQ+j2YHs4TtB4Yv1Ve
lFlSry/YtFRpxfb0wlS5H0pNLEfWgT780mP4l/GMi/AaIcsas0ILKf0inHxcyB1B
EYpac+k+nTFOFlM97+bN5yEaXq7VQxDXApoylh7rrHG53PgPWngBjihWjmX6FEWo
W+yzpdamxttORUMKcOwZeLaHjCkvEbnPFTzYMY+UVNuenS1x84R7Gn99qMlVPIqu
+I6I5I9DnccE6n6NYj+yZolfw2Vq9Cu+dclcxp3xRhY2Zuui2tUgzxtx4bSDgGEW
aCFD0GTVhLNOVwa3TEG+qDkjWLD/1jSJBErERcLfKKdXGLal3AnAup9toEO1u0X3
whwfmMKv/J3OOtuwWuMCqXPI8mDox1onByCW60ky8FduFaXLwthpsPj0ionWZ/fZ
K8vAWcSOy05CyVUdtP0kaO4mQpat3jiNtEpyHL1uCs51aLbkc6lVFUOQZRxrTyOA
Ou01G3yslIT3iHoAr5So6L/yjzcsMx94pHdKaWEdj5O/MmOq2shTpaOdtQ5Y0Pbt
i6ebJrO0eMVL6A2zU3vpHiB652R6BRPoXpeK5UXr8nSZZs3txZae3VQts5J8C9nb
OceAHK6b65wKRHyxGQWg9e88i5qf66SUH1B550XT23lDSCkD9kQssFPnNok3TlVZ
gOKr6WT3Mg69p4QRaSQI3GQ1HO1RY1YatwON4PVEYkrVT3OtrLPKKoG10DJp1Fom
UVcqJFDFr6Dlcy3o8xL8t3Kp61sgjRC0R1x7Q0+Egg64kw2aTqq/Cw2f1udYVTeP
N6+dIb9YrT2KWEjbx+BGFWTmuNMkCUpHmJcuuf65TcvrVVWO/x3HGddYFQKEgcL5
mfxSdzI2SHm99AAZl5vVoMWtUVGmQ9/Pu6rDJu7iNEcZY7u501Dg3lHlT7keXZvg
LStxsG/BukigaqArkQdKDxls9r9GfVo6EI6+uthgW3ygQ6Qsy5igXe4rkaBkdeiD
bfaN6mpDlvv4Ps9pL4OXMGpCQAlNTZWilwYfi+gQW69WYdUxjrm+QURBKa9FExKk
z1k4T9NxUaUM+DmlI7sGKXMu+5LRd23hrz7wsazA1VlJDyuUTI8ucR1Xom9JBPO0
ZRH+P6J6Srq2PKoy20JvTsyOEkALuXmV+xUovFjxOX2k73r3e3vVmmtjjcA9Vrua
kBhOxb4Q501ItXh/fWhBfmoBUF0waJv1mcOb8gB0Hg17aH++O66NIrhN2pkRBtV6
+YMWJ8YB6hVqHKOiPEx5Z+nF5AXFADgGC2pjaGwg9vSxxjNtOdtkN2h7ZH5cu4vd
IGwVdUdoT6laUk8vdZH1F0hscKdJD5QUE91wrv1AhKigPEWKAD2/uNiDUVY1fkz7
awO6BY6Wtx06tNee6YKdSsj6ZDBM5dCUK2R+eTeDTuTASsobRp9WViw5uHmTCK8t
f3QK5My3RxtodqHaGQdI3QX8h7V9jBjW1eTK7I57z4Hb9b8VNC86Fu4CFZp/7J4J
4/RrmimkFzbZoNhnkQE6+qx+ehE9/f2DGYX8vNvyJePaGgpTWR4XlpRkYBeU8/cL
NdKTwVDgEn+io90nZrtAiBYat26MCsGajaAwmE7Gkkq/Mfpy2+E0swc0GGfNDEP7
w78PbWGtuLysR83/TnYDqeJ8Xj76Sw7b5YmScHeIfjnuDsM5g8DJKhd0ZX4b8uxe
JV/YbTIxGtYupbe3FECfnLDyHF3T7HRetrbBuCS0nFv1HnDwbE674Yq3ZB4KT4PT
Oj/z+hZ3iA+9bnhVXjU7eihgf40gapNsbdSqi6gc7vrDVPWevL++qwVJRZjoDyfw
YLZRerJYQ5fcvqzsaa0sTtCO4Ic2zIQMM5ARCRr64OgIVaudAC3J30GwtBy/RTDE
zfqkAlCqKfPCrwWzrzf9TbzDqPIeszjWQwCvbFSViDEX93FvJXP8cYHZ/MKbcWxg
S9+yy6SMc/9wrwKm9Xd3qlRvl0sn9OnMeCHp5IlGqeAhHzn23b4URffJkrHi/dIH
3CeHTh5Aa+21CucUnv7R64mu+O9vV5MTbofxgqKwYor76wa0kCQOdbSEITdMfNrx
5Hv8TlFsdkG0XdjB4B8khm+BfPNQagdcEWIR1QVxS/P1JFCSyUsKmYn1MVrsrY+Z
NfgpRHsY12wVKW1+3258/Oy3UcHqadqA97PDggcLwoPHZO5adDr396xbE0r/oTZV
whNgxEIoukhxYK+di6YkqDGLkCJLm/Ck43Qn8MMuwSIoSwZNNm+ghiBcbgHZPycm
C6qltkQnquUVW+Kdx4X9u2HPn8Nzz3vTEjqOEZ24zeKA6CbVxSw2W4oyoh260mEb
ZrXjeUmbhN7qXmKtVAw0Jkq+zjzY+mreClJjPHJT+nH+6J9hSoniwneHV6ja1VNk
pbmKSJA4swcBh35HzI1in45KQxnCSJ1Dpjo8DrAI4ntVX5lRrzrzflKgFhew8uGM
hfUzlpIyn1NigdLezasVlMsarhKBTP9aw7zThVJlZ3kqwLR0MpNZHJWCcY2Exn5W
xV3Um+1b1roVZhIM7K0OzdogpQRmAYg3jXorBpsuwPKSWgQYxuxpWa7p2TOsD2Zs
subxObqQIGtGTqS357n0zCzNkZITAqfaEzZ5uCPpqDMmGQT1aL7P2u/7YZBihRUT
hzuH5t73Z2ruwwoBzfa4AmIqxNfsQXscvztKkUZz2ZmbBi5bP+cHqwRqbz3B3uAf
JwQDDY+RARjIqbrgitQYC5OulwiaaGfM8yBHjLh8DF8yvMkcTKq0g6RPpX8zhTBC
QTF5UloQzx2253QAJKEMstkKpcnuKcLPCWbEylYaqO0It/ETG7tkslUHXSPAkbSC
z6yzvrA4ZLIeJ0SarObvUodkn1Gl8W2QAyxl7Q1bUV4dwEN2oahuHYoYWaJEDJup
N0f1CdrYSAJl1hKI9GSkUuDszkgtw2Oh9P3FeuD8D1pDJagTut5tJANiuSwLYQ5w
UToezHZ/tvrqcER+k01C4uSS12V0vMj1qBe24S5mvt1OWdQByzfqhpeOoJMhtN7A
cawUd4Ah9LONIvoYQmCXJPPLPQKxPk+RrPXRC5yRFfW4nwq3X+TXjPgRqW6MVJPU
a0tR/O7A0iX3cC8p8XHIEt+9WCrAQIIkJLctHuM+TSK7qON1xIpS8x59tj+rx1u6
9ALZ/s8dVlU6kaC0QXMHNF5MZ4j7YL+rF23dmI37dAvI3YjuW4O7x3sLhXHu7VfT
Z8AaVCdXVX0GHBxHZ1VhgJ0irG6gJaAeS1aWlvlbRNQzjQ0uliZpIfjobVyA82LW
V/3b0lK287yWUrKwOHS40Rb1XDe5TMaS6wNCR+SA5U5SIVJCfpnyqN34DecWyJ/O
2ZI5zQgmz2HNdtlxkNOjguYh9rlzgSoQuNDUE7in6IfnVRqRJPkjxa1rXVDkqIbj
LJL+6oDjKxiS4xUK8sF+01A6ybW3DGN4rcg58Mpnx+0jzkj/PsWN7hNvO9vYJs3R
YB0W4Dmdy/bvD8lt6Bud1tGUG82QQN7+cpHUfXdn+BNxibxIdNBHSSV0hZuhY+2z
Yk1tUh5vx1AnOA7tRnNZjjjVydhz5qp9UQYD8VlF4TcO5BFdTPszDq5+FUkN1MiO
VWXkF4L2RAS461RZrsY/ybs5Faj523bBx9zjiyy4xlAGeZMjvYBCVurKQQ/vrJ3B
zj60yY8Lln9GNBYbfV8ZchRiWLc0gHqy4rvjUU3vyfSUO2c4r4+4kCNQky7p/n/d
iMANcr6v7tZpQgzszIFnAt6ajpx23b5cYFwxndoOBmPtTmzvdJHmvFRc8BCBVTJr
OeCfkHwvljfl8NGX3Os1eqo0ToS10Bicamx8eds+3+rZwyQCgw8SxubFFqONGoSh
Z6g7816qqwQZ+aS6gTgvhBJYahlSNe9UgEK53b7DaxDzH3A0RVO/EFKHOMZBcSH8
lP26FzNBjwxJu4Huj6j8qLWT/VRy44UA2bdSPLm3vfqLAF7JkzRj6KzuoJjSQMhL
WO/BrsEM/SJZHdg5IBVSzfqc17x0gwS8ttmSfZh5SJXgovFXXGCIV2D4WiE9MIMy
Zl1+qEfk0pJ9UDbnFJEFtXNAusKmfFEIeHnJ9ByOUOovg4e4fd+hbd3Xl8J4SLeb
k3/k/TX6WVau2sxUJoXZWNMM8/t2nsb3FwmuJZQNW+tAkn3wcodsAmH9oFFFg0PY
i+BjPLmEqQjL+wxrSaisk8aiHkQrg+34sI5HnW2lFR4cD30lIhZ5BV6qzQ41/zup
bCjFP2KaSEaO5dcwc35pu5yzwGyondJbsV2iqIPlOk+VJ22P+KsBT8mOAr4KNged
nKzEQFpbLOVhvm3nWPSiNot259b0sngWJMqiYq4Tei7L+uhBRW/D3PRZsQJRD+uY
Rmqvy0DzaiyMl3bVKWzKSJeAkJDrXeukSgR+xtsifcjwWysp3vp4uiCIzv4Pkpr2
JT03o6AO7QkYB/7pBu/eug8L85rvWGYlkES1AyAqJfVytLvys++N+ccORk2BYhQn
YJQZIX3D8K95yp+gBoTibwfmkpn4hbAKngjGLmF46y9UIRN02lbmvdtW3rkYNM+t
jIDVGAuIUVDEKwQgWEA4oTLBeUk9e/i+xxlRfuDCo2eDyRakmPF9qmK1gnLn9WmS
4q4psHIdVeugaWG+DZwsWCjnDcCuZ8D0Bt6dAmm5BpWPjub2WIcYMWqh4O2Ux4wz
7EyyObnf/KeyKrxaXkbnIOxSwor2RWyJkSTLAC1G/otZhV+K11DvKnIz9u7eHPZU
nyOIKoQ2QTzrX4o34Ghg7Iz7kmtiSGbW7k9PGcsfJegwfMByRsU7cySH8CQUjMsT
KfT6i0LXffaoVPhAVNa7Eqmk8picNs8HQH1an7icWR/pddAmMo77n2Zayf/P9E+1
N9rhHnkc+YhdWKvnG+LkyRRjzLv/nhotVqPUs5mHVtGRykLKYejtxM6i5l8IbPXR
60UTlOpMYyXEUv9d+QiGpukb8vvUlu6w2L1MA1GQJU7nJr87BHfZ0AtCtlD7kZTN
Vu25NO1Pp5kcNh0XqklFSGIeZamiE37RACcTbyGRwJ+WqRJ+r2CsYwmLL3Yopg7l
0NbiztmupQurNbrCqrkg1NiglbNGpdv8JhK+1TIxYxZLjV3q7TDEOCpikvaxAmjZ
gTH8c6i+pFCuDR7mP+bcBC5ykNFesWxA5QtE62kmF3IL1QlJJtBvp7qeWK98xxYA
8gEs3xkSyGHTiNhkakWdcpzKFhH5dXezikbKlJ/7EjY924oWu2pFE3RtpGz4irdj
ZI7Hx/gdN5u6MgoUkdI2kF0JmG70/HwAeQa98S0Gbf+QnF3HSPiHmNfVlzqBuZpW
r+mWC0eMoBbPjT8X48xPg/3fu9o6V/S0dLw7IL6+6DUdhNmvUWu32S0zRgU3ujzH
2LXOJG8QVj1u51ZBs6UbiKxbwASE2nZnl7Bky4KTy9C7y/OsL8wD7JLsFslnOk+u
zas+DflqI2cJ44wANy6l4YHfgrykNlSg6B9a7+a7qyjbcxintUMFE1HCk3jpbGZ3
tj/guH97UMMpCu2Xj5EM3c3SWvyRy5wJuKYq5PX+Qe4ZNXmX/5EBkVs3Ky+6h3Nc
3RA0PnQIOj36UT/VtHro216+ofHOzeybcn7W/gMsO+2OVYq6MR6tB0skkm5OqmfM
JK5Wr6bkiAEcdR26yvopu7U62bimP9+M1ll86Ga1836rHBiekCiYSeIemK2MLqLl
0ykcBKXmKPOxkuVEkCBVtzknA1wglWOR6C/RCejojUPCiBlg137gqSp1qDq22s1t
HCPvgNHC1aT+pdLhocAkaKXT/4ZN05vK3aMleI6MTqf0tR5nm+nbQ0pjKUmcBa1L
URhvKuMVe/19YkolQRdaLXY+7RqgQUUy0oQ0ZLM5ATYW8/FULZbf3MKl8KjrEp8o
aiP+OppAMpdTPff5n2IOtz79jEGy9WZWlB0VFgQMKptRNwE9VSwNf3+BIXx2mggj
IJAoRUWSsBn8gtAbpUF6rM5rnkM2mohNKzGX7EHP0GLtIuVWCEKwXcdlHXiTjEH7
jCqTPifxbSsrA9m5Ds6TofpAFNIr1eFjf8n/jI/3YAg2J0LMg17zraOtiKgDzGYZ
BASo0G57OEu5ZKN3GmRDEl85FtSFyTnzqIgv+wIaysYSb4+TONuQRFkfzkG9wWrI
8MsY9IRs/6tVODtcLGQoGmMNVKhPfZeSPg69p8b8N3YVhc4hBEoWPqqe1R9khpAQ
cf4DvVXV1SvVSQyiJuC1lkgHt8z8L0TNl2T58/dWRXpWj3Xn1JQAjdm1rV0uzvY8
dzYdpgWhUO6q/rLLXmyt9xu1L4oi+Mb1XwSkVp7Kna1lYnvdRYjDFvwi5oXoa5wG
/+VCCVOXjiT/Hk6koWNjD/GaP1OZ+orTCqy01knKXrcPjEJQpMFWUPJRDdFq+VNn
Zjz+k7IzQFtrvL7nX/Php3IbTQuTidw79yeRA6MdC/8xSwXXCJ0jDXffrt6dQh8t
m3EHHbZbU1IKSoHgo83usrR2zVVJvlJWfmoWgFgF0WoqfZBZh7ALqGIf4XnI4qo4
cxswM3VS+qqAtzw238aF2jGoktyNaJKkHWumuhZVHqiIEZs8Ym4vL8+K7Wy0QTTM
7oRrmPyZLGlTKa+KHJOuwxB8hn3NDjYpKSqQzGGLsS6So+EJl5S4dLCyMTH4ds1i
vLXPX5Hk2iINyWM6VHhfIBJxBqGlc/Bi2BCIHSYn6y+niZsN14s/yT1/7ImOkKTE
PKCkZR/POMLftZ2sCazgYG0t5+72272nVwrO9A62fAnlVrhWp6ofQJ7kxsKc2rr3
X3OJMvyCu2MCXD3XVHWP7e0HBw305wRh32iwS9+deFvfREYkTDDDE8lOIeSQmwpq
EyCCRkenr4mqL8t/2J291ZKudls2zRODmwXUAiYa/Y0UgKjD+n7Qx84xiCWTKzR7
89KFSILetwdeCDDxOUX9o1wOtIbIllcRD+9yy4pUG5o8OKZrVRZfaDzEKHcqThVy
G2DFHnVnmGdMjhQdwJRdvZhjR8RfbBLV4rJt9LUYyG5UfL/avvPC/RGce6Z1UC1u
hxkFIrn3pgUaL/TUdNk4pT9jUMBVouqlzNeXaA7OvyX9/cOYZqZ3dX2xT0WPRnXR
wr98glwl45NP6Oty1ucbYGmO0kCTjCxU9wklfTSSH028Y5og1G3B0P5/f/OjTtol
2k+gCtdxvsdDJVRpxbcVYoST1CPGWEifRyss6E2aeEspmYCyFsf4iSPleOOI6v7M
iAA1p8eiqXjBnPgbGXnCmHQIUvPDu8eHGujiPvCRvbKBAcK9x9og9xQMEoW5uY6i
N0okv5KBmStP87ja3H8YteT1suUT6GQuXqyhe48eURVuM/9UqelJD7kjql0fR/uJ
Zq2TpHqxB63zTqVse/q+1OPSZS9ZyLlcPWC47iRufyAlyrgZsa3FnKYRciZQghDj
/7sLaR9tsjOxv3/aB7os2tFSF9SLzYfpUeFlvWhn2341ep2/+BR8YSR6FJYU7vSB
DKhG+n+BPz2Kjax1T7arb3lbKP62oiuFKMY08pOasOCzB3d1LyAR0T8EdD9gQuCl
zX1cVbi+WFL1p4ppnR66tpsmfwzIrpCHne7N5qam1ZTeRMHthSeDtp0J2uw2Lx/L
8QhJn2TaJMuAcZNVyBc6u5eRXjUI3z2B3dH7cDmek5exEbkPAtWk8xe1K0goKiSb
QccN0y9k8JUAj139KE6wZQZwCT+0gtFFaOPtAAdyC39ZGQ/2qUWOYP4nSN4loROn
TEaXHG4iyAbQdvRhAKAgAKb7CwXFoS7Qj7MwaPXT7LBxVhdmChqmULvu7U3RdWtD
C595MiIcQjAOXqlkm1q9RzZDXPKsTTprGI33/LV5WMBoBIv30Ru/POOUKF6XLpXF
F+jUrg09S5CQsIhFMdGXj9OUlEYSEqW9Dt+W2Mtle/9cpX19RVk94D+Afq1zKM8n
PQfShImhAydh9eis9pZnLAPKwHN0S4fZwLqfrNzl7CWwqNVAfWDfnJ1U7WBmHRF2
LsJAgLvueA18SVLxl401beajPcJtmRf4jyIj9lZl2MapGTPclIM9cqOb0LqkTLS0
kPiPZOj30j22n4tFiB9YiHj41Kt1W4diUNZMMDeHz2KWJfs7M/5cd9Gfxm2jsQm2
EBu1VcY5SWZuw/2b2unG9awTrIruHwnR07lc03Mt3+1FJ7Zevcv0smRvEeJhMTiM
FY/Te3gW5ZrmvCwzrp7SlKoll3aqRqWISA5WgN2vZ4fryRaLz81+kC/zdCm8Bi+A
g2MJOyZZ9SeujigR+qhhedcLmegScNjY5u78tYZAzxbiA6cfdB+DPnAE1jd+nNag
9BtLasDJ4S/QJbG4RhrQ2nSPKBcDgBH6Zzb/OhUCpYbipPezgdOvl4lr9TQoqf3V
HJTNCgBXCQTAoNb24d2k78yOmYaOrR1YsDQce2PBsPMbN44zSKdYlI+xvtz9No+N
NoPyn3oiB/k3QFmmZmXLFmNkNfoFny05cRt6fHVrra1dkXtQ+ZiAYSZWxEtX79mA
RUh6tOOnKfnOjOBfNEKR+lJtpNETQZi8KUjXD5Frfi2Pyxq3lXJfQwjtzptUqtIu
DMSvE2kc6EE+MpKO0UC1jffTR0DSEgW2PpCbrbWpBcsGeWfOc6xbCDHEvV2iX90N
nRcxnwP9d2ObJ+FT3bDykOXgVnYJAF4bmX343cLWT1OL4GuYVRUSN0FDSCRk4d7N
SJ7WuxlGKJc1eu4H53MxniDaRXpMmrRwWfeHxzEvfSA24AFw3nA8y724V1JilSEV
BpWfG7ndZOLv6uC/dqDqxCT6FL4VxMWg8hHFdU/kWD58uYF1j3jgwxLXH2/EdxHF
Qbz0EQ5qqxBHY0C8JbIdpwa0O9y5C2rixsUO+PIIrMsSWTjg8kUvvRWBIfEVgwQs
L03ShCoMq5UqThMc1aqTyc6D1LdWuoaiDddLwiK1NTXe+sw1UhzWz6kfTagFyco6
Y3HviWL9A9C4arkLo+9w+GLzif/MpF8pOvXp43nHfSpJCND9wqdyFCTEhZ6uH7Sk
0Ha34y9x3Q5QKwJ2HV0vCf9PALvdjtCI7DG/O4NsYddPZVflxr72MRIPLa1sg60h
XhjyLhytAhgC7dPP0yk3l/K53vu6dDnEIA4ydg+XG78aQUUbMvAr5ek/Jh64A7vi
xF/dwHOtRHnvxeNRqa5znx7YXP+HZh3TvLY4N8uaEdrn1maJMcT5TenPCU7H2w13
zzWOT3C3qeXzT9xQcBZZX29wMXlkPEj0XKwsHbT9R3CwVFT8F+12NPViOUJuPH1P
34i3DBDRDa+LgMJgzAsljmiq3nQ5o2lBLeEM4TLFet24B28rDCd4A6uT7RlvSsPT
/gkUT+5iCntHG7SnDlohgKP5QCWSSNdjQJrdWxABKcnWQclqC4ClLyWfoZ7zx0V2
9hNZgaEBHHERu5ehgO9dFpWko43hWu/WiqXVGWdeolErZK+OB7G5yNZ3BQ5D/085
kwkM0tbL7TlhyVH4EGHO8TbZy9V4vmxu3ohzzfzobsht6owLm+kHQAiBCZjjTmv6
5Rfetl6aVCVk2ZGF1rf/FbtqNgT9XTQyOa6Gj5s3AKos/nrWBHDu54T78HFrNc3E
OUkIzLR2cYzMUQDHKT5XB12GWhlOq4wveveWva0d+tccuqVePzkeEKX2VPXXiX9W
/4x+gd2tcmJXP5mhA8582oJAHKXMebgvoDq9yAm21tu1W5d+1o51tDTFH1fCRGCq
Kz59mnVEL4i+6logeQgrpH1TDbnyccTZxosJFPiV45mTMR3iKI0rXjF0sQG4hZQh
qJl6g1mPBquhtEe6gYoJJXomUwAvMcwFBWjjGShfGTMZlE8+ZkDiCpvdrgx/Gmfs
n2kogfUVk3TIxipkEgbj982jtzbR+CvTL1UEMmRBgoDgVHLtJyqy2zDhJlGwGjvb
mQadACZLcwW2vImeZJst9jVfyKyTj/XZtSatbRPv+QINyXzT0ty6sAn4okm5fykA
gZWONyyYgStMRih/yJ4V7wIC2DYEt7dUDGqdKoPTD8a4msVunsUsDP9p672do2ef
y7K2OjrDehMhYRPWFK8p3Mwu6PFvcu5P1W/5F/f9pf+4VQeB+a+WUPMUutUyhRbj
+qNov06QtUkI8TWoxdw9qvKz3sW856UtDAnuil9spJqYeVzIHvaS7PvKhObVhqvz
Ke0VtMl9H225bhHwD2DpXptUKpMk0wf3bZ6GMtnO2zr7QxQfOZzfY37bgBXCD5AR
d03Hk6rGQwwjmnEhrlpqlmrJU3wwjIUVfgEIGSQmIFG/hX/aIFA3nod2QOjusYch
K2nWwPSoPNhGmZXtCvfyFcjP4fiHf86mi3kE/JSkRtNawEptvhzsa5Pb/xm6lUgX
x42ZcLGMtbcEBWz68sqLvqvq546XQ6g1adNSjgMPesmtk6S3XD8lJ0QK8vBe/b/k
8dOPuT1f4CSu2KjubQJYjavYSCN//i7/B2mnyoyZ6tFP2Z8w3aR75N75TApIBW/T
Ma3gs9RkQP35g8gG6wjOf+oyWJCVyarWezEiwo6qacIWyPdKhxYFqwU2bo9w//7P
kMjzdop12a4MVv3bxj30jTK3G31gOhXt9UjMKrhnXe1gmYnm+a3S4F+Uuw6aRIrM
WqawNH0+ozCeWLMN/X3T1mKUodbPpExkqAh+HhvwfKJ5F4UpwjiwlKBWRocqkeMx
Ao6jlCcMA2HCBlgtxFTVYGvDzDSnpUsuG8VJ/uYTQtjBYQVDF5slHxF8+XVb2IWg
Np/HPFpjoSDEGOSP9xWmnnYry8KUuu6QDUc/XVAN5+mu1GzrWExwSOQssbR/pw23
9x5rzL2nNo02pDtvlwFpbb4Ok2gEd8WOayv0yZLVJMUrnlEJl54IiHoMnHltt9jp
w0VjVT7+P117oOFwseHZ/qUmwVQEiuoMC0R0UnFf7/Qd/l8XcPWFxGe9Es6McLhD
0/Hju4JqB+Yror9I41UhZQNi+KZYf3Ge3wIz+M9/iEnsK+O+3z/PE+liHBPyBhYN
8Os/SImPvBzA5FWXuGdYjZl9Q6IIXn5yaRzv8vsicrtg6P7wPcMOI+UZs0qqUIRP
ZGOmf6lZxO4K9Y6kMTiav0QlgwmrqTXQeys6Oo//ri9UdCZfbYhBtm9SdW1rvQbF
X4FVu1PyBW8i7P/iM7s4/ITJfJGzxk66M1rAY0uXa3gMJWfQVtTJ8HgUBYNGgGXq
ElxvKABSWrheiPFtnelL3MtfZ7LYgsPprvY0CPAJ3ewPy5+L7HLO4I/YChMXFJov
0/5B8ffZUqq0phucUaEr/ztjasPGtKpCSzliXgOUDrx9iCaLJjxsnS1ft2vAFGQD
KcvULgtNGzm5EY6b0IVgD13DfZOQ8FlxWqqdDMHD+Zb6/Kgl4Y3MbbROoFQn/ZxS
XlM7A1WgUea1jvpRbGME5mmWRz6vCYrsBpwfv1fR1+DlY4K001PCXXA8SH5lywVi
iph/IrhzKyrRtQ538MTB01Pm3hv17NWqrtAEvSPmsGb0KkZJvPh55XVtHruOiywc
/6D8cNnLusAIe6ZHocO9UeyWA/pCXxkIFbhNfJ2OKOR7BwIrhVly9VrLndTHqraz
QlKPhg+7/eO2pY0Nz8TK2CMbA4KW7CR15/0wVkksLOC1Y2OUTm/ZbzitshHCaOMO
eZeFS7KmAylOiJh/9hNuvnTWBGYOno24U8YSNCY2nzRsTDs2bchvHzRmwByExBec
3It/xT60lGEf8wus8Mg/M+jiEwEjoWQqj3YzHT9B5G53A7Fpy6uZzKiQxZbGmImJ
K66dBgiXIT3jwHrKmBGO2MQFzP1JBNtEap27xHsEaPYYB9npm+mboKpZnqLgoWTV
U1a4qyyDuLzvsvd01yCxMk9m5tQjPcTgsm92l4+roYW1A4adTuyfkK9I7TgOU72j
98QR9MyRBKISOCfEyyQg+wIkKjcH6tI0eNmX6QT7cf544VGg0CPeQbmpSic+SfkZ
Hh3kQvREVz0t0K2GTvJV9qjV7lMXEkhlQLB7dI+ZasESzqcawIMV6Jdmdpj6S2s6
zsUGv5ZZ6b35EEzFdpGAfEnbFNFCp1Hy7QMtWmiws3vnsQSLamzM8ZeZtfpfND3I
1bvEyGbO3AMfqPmI+qDZEgft6sOSLaPRQI+gIcQMugDbKyso9cgQOMrMaoOFGb6d
Tm+63Xptp0xvPsim5zERPqvmBvwkir20aFr1HaGWGkkUrDVstmszi+S9fSvfqmOF
1Ln8UWyR8qnFUvmXMqpzCeX4v92UtcCAjX5o8yFoJXkJA1lHcW+/09jKyKReHA+f
tGJ9GbSqbmOx9ILMyeAQLYJC56Gx/0mQvqGymK4rQiSPCOHter69/G5NL6oQ7iQ4
ebIpwdo0cp+CC2FQMBLzEkl6wUe7Hdv2KUPs8xQLN28NfEjtOI9//HrNMAEpP4QJ
ZnqPYHqDR2UQpmdXQ8TzfKaDdDr7eLUbQ7vIPeZKbdqu/WobPE7A2oj+JsU++Ewi
NeVU1ikW10/gxyM6PSX2RJme4Gxg0QZYaqHJUl5ZUWd+iAxJwqATSLSPnCC2MjB+
gAA/tzYKhYm3fL0QNqatIAJq0QyLN8ZjZsMNNGuFyGwGnZlU62bALlRnZrmgwaPw
LCX4GhPMj0dXAlyC4VfngYJDqMBNi+mZba9e0oGUDbx7azILGt/iQxeu5iM5x9FK
RGA0we8WtkpQiE+V+rNVXcWEvZ9vje2NN5U5UosBAVGGq1oZxpAVPikCulypHG3M
/BgtB6wiWQRuYbnkQC8L6SIfuTgvn+QXEbsg/alSs+iA8vZKBLmwUC0TSbp8Q6Nz
Sa8ZdnUtp9s0ZgUtOBpZjsTbtQzSwAIOlZXIR0ntjs/RSoXMkmn7Dm+zJfiTS8Rw
CthFMeLS87ZTPH/G1sOAwRTp08YLcHXgpG2g1tm/fwVlca38x8Y87Y8TkGEWRr+e
EVZna4ak2GLN8RiMpPYH3hWUEqJYqhSzQX0RIHmH31NJkMLEW4QWF/W3YdhZvEss
X8Ri/YQ4WWRARalpoiTxyerYsgptWZkMKpbbv0kD4/6KybQsiAF9Ocw4NEVDY9k/
fTk4hQVAsWN/2iYc7DgDwkQgJN8th7JL7vMAYYhguc8yQ8Uxlps34D9GrbQsHEF3
2c/yNA1dg86Iv+BKUhL9CGOEo5dvcHrDexSfNl/QQhs+omlPzmteATSLLTZBngus
06QpJEgDE4BdkPcd85i9Jk+IrRvkQsgGucHHIOvErFZn5JmJYy0ZFmQGeswLgIRX
VEDqwqsNJkzJ0y3Xw+GyrU+q1G354QcAYsz7ybYo4IEpXucxzDay68RcSmjY1nu6
OmBMnxY6PwaHO48ttdrtkDpaGU/R4dA0v2UDLl0+dH4WlcT8Ui1hFUUr5Gr8p2Uc
a1wrUgsK3TqlPP1OPX3FrMw2V85loJDdIAmft4tZlm9bsQ3Ep1iaEp0OyhclcK0x
mcQo0LFjMWRB4NUzJceoYrwtr8gFg6ygfa/gKtTyAm6OUkj/auI9vzFJenoLyVkM
langgIBLWvu4Su6XZnvqq8oulSKT7GPrfV/PGT97iIq8iETw57lVQrYv0IkawiAe
x0M4S+73N1SZlWhgg2Pn2mjgLal3ZMFD58Gnd7zPCQw1hLbdP36fjoEP+zdR+C42
nV9apGN+CNA6bjC6+StPnQAPfHyd9thqvYjdNNOMkdftmQ2bfvDcdh+yld7gX3yb
PsruZwpZVINYng2R0Sm6BM8j0d3fcNKwjWgtfDXqgnfF5FUFDrVv16o+SxtLgH6J
9pJvOq+3/W78PJWm9rdSmQnSgY+gjPrnMOqzjBpc+sQvhBSudHK892wg9hcgfNj/
Bp3fF2kfT8Ce7hEkQhwAXv6ndZ2I//N6WlOGsABRTqyCh6cqhcypd4Mg+E6xBFZw
3YsLbwnsJ3Gc9X6ntD0o59AKtxWY8/h/D/McOBldAQ79eotdkWh5LoTO19keBuNt
1T33mcWPUh2twny8raRSEz/k2He1TvDlTUyZN2fVmR0X3uUTJOdgHVAygtbduMIV
BwLjjvpsS8u38xgvDIUDglE5X15nYoH7lnlVSlT1S5igr6kMElqEsdvj9KGezKxy
JQgH3VEnMlZO7aOV6nyHyilajLLIuYrS0NAnTPj9GOL9OflujlMxPOaTwH4ah0xR
gm26CdM+LLRd7+aZjO2Sssi8cAJqoOwDz9DCQURaxHh2d1fvxED96G+hEzw2ITxi
BIbZHqflFUyrMo6ci2aKEtAnbzubxuooljyCvsKkuGu0ikLa+JeHA/DBdh8QAqCD
SaZB3ahFcvYW8JMG99ppGZF5m+auHbSiu9SP9eTr4tid0YeBn7zgtX2oe5bNAGwY
4nQaxFlS26vxv4Dy66zdiHU2EEGCB68Ok3/HnWbxN+hIw/H8YcozhpcfMuwOMpU/
KxI7SK/0eeAn6BcFyGHnpkWrD/9J6xc05VtOOvLwpKS8LIloMGYhkdC10DFcrDHf
CJNA5nwPwMc0pCM1sW9bjhCNgUntqvoZElTLNww9YR4NAuO6PKTujXjzQIu9j6B7
v9VENijbtRtzWrAwS3k7CH84QWTaKY7CjI7G88nsAXbrokKwd93BC1uiRgO94em6
iJd3t0Ix3x0AwVd1Mc4oXtGxdYJ7cOS1w2HVIwAUQdowIm4nGFRcX3B0I+1P2jZ/
S0S7hNX5e1TKcVe26tbmg+5ncS9xGEHlScs596oyZJ9tWGlghHjSVZWwD+wnjuBk
5dhjLyZ5gzG4SHad1auosjeYKQEj1KpqIUohzQWlMnVLWOR9E2cqC5fSZNUVr0aU
sjxtWFZoYfO3iDJZ91Kx/CDD85zkjxKI1l01nXYA34vWr1uNBo77Nw96GaDJEbmf
EX1agZvWnv1qarmc+hlvwOTmWChj9udQNt2WN8sThFT/NdKPrMPUdk2YEdhbyKjB
wGjp0Xf2BSlI0/suE6H2etKKhqEFz52Ad/LhxWp5Hx6RQHBeIfVcr02qyDV7leaF
w03UFmvcMBtA8+ZsfEr0itJHRR5tNxBGVokaaJsqEnLKFUwAP1UYldA6OYPJSvqH
zK5Wu+uVqHr0803B3AuHVx5oR+yI4qY7ZdjstHDxAD6yo8G20xVKxF6fVEKi0jQK
LDVB+y9grhsCahqhTpr7bOrKQ8lp5RbPK+cu9HvxrhFj/nLo4Ebs95DXCY+GTThL
+ZycM6vjnr8nPt94jOymhlAdm4ymWefz05abQPZEzFcoZR9auUXiOThcc7OrnHQo
vIfAFYLSV9P4kA0Lx8tk7Tjewpfzr2/XByF7fMmOtKnfoBavyjfdeWlEyf93UAwb
dEe/X597PAlyxJa8p8kggs4yMSOl89IQhgpGAspEMWGe1ppUE34WyiOUu5VKuG5G
e31WleguryKxLsycytmv1Q26frdSyY02CyKoZpN9etbLF+jhkvXVMXu/E4td3cHp
cnN69sfUc+O008C5mFEjpBAVxZQ902BA510XeGGgrEVRWP91fAHoqERYXundaTFt
IE8ST4F3H/RSHNCGmkB/gPESfYPQgVKQ1AWMB1pbfVfnot1gdjGywXkGSQGewHBi
dx7QQa/nbvaoa+Xdv5gaA5xmP5twjUF5Rh5pLh4jgRLKZ8/1jFC49N8Gq2c/nho1
Sjg5yAJvrGlspnqPGMXIM6OthSO9QF19FymCxjrYdpEV83eJVB5nGm2RbcYsNrU6
sxcZGo7gwfYbFVqiAIjj06ona7/TLYTovcZWVUQO3D8p840MOvUrdDm2S8m7gG8h
UzfIqHcVFgYu4FDKRMA3uUjcX+wYsQhHCBZ28xqjoRTqZbvOoiKhStcIHfGLU/Pl
xHmEgW8bC86fgRPQXXwjDOScNReAOeUjp0fVXHR0AO6cC4SJrR8XkyNgp139pZSj
sDzQk2ldbFewR3FzZIrh7wGuYB1RIqxXnDsFJejjO5NA/3DY2DxHaF6Aa/Ousqma
NcgqJAwLGu5AkAyMSEwyb+ugu/DfZc9rUb4TPHsRHYq5nWqkQQcVzBTjWpIH5XLS
UpT6sF7pWpnlVpEqXiDJx1BP0ZtZgDcgKW7OTuBmaq0rzO/OCVf66YK2ftlpGnPq
yPvvE0mdVcfEdqNgd1aCI9Cj+lk1hU2m1vBSWntTPp2BPbR08UIRC7Nf+VU2UOBP
nE09XKK5Mij4CRH8eO8Zpv3P4W3DyFo6XpM0a7tehfBTf3M30cecpy/ufGetKTdO
02ydneShTDuieEP4zBanH3a4yRfGCF9mCJ3JcR+uBi8Mj4BSevke6/7HZSOiDh8D
Vy79w2Zd8sxpUo+2dqGWzxInbNOAeCM89nZWHkBm2sAJMwfHFu0NTP1UluKbm5Jp
5BIVY4wkoj91WRLc1KTXidVDdozo2V9VYzxsXtABxsNXX7VzO8FBsjdDqOCpQzQM
34pyipDIXtrh1hMiHErTo4wspC8VHMjAXD8NiAWpnRdCBCsq83a9zJKvCw6Uz1jz
Ner2fZbeNwIDE6BofzYulKrlcqv1dYZJJQGvRTh8o6oePXEDZ6moxFng+tWRnATN
m5k+6Uz0rLEe2pJJ5kdqlc+ji9C1rs5Tn6lJ3npPRP9/nN1wLEk6+Qp9Upkdlc4W
vTdzhZ7VPsK41Mgp1Tg74zoXocZS+PpOJzf1jBoxnkS6UYaQtOdF/cGPMuv4B5Sq
2qTXGJwJmqHRafp2qDHVbVASPBEtuRduOLPAlMMTEcks3uBRKn0B6zAk5ghmW+V7
bAfye9h9THKCMlmzHpmYbe74v9KWQqBugi7w2RZ3IzuNKOZ+UsoZWDflJYhmHxm0
VGYKvQHx4t6L/dNVHXjK3Ev0E3LLV8cRa+WZO0JT5ANs6S2kvPRtdkG2rmYMR00z
pcIlG96qaHL4x4n9pzhIwkRJM0wkv1aGCtoVyKo9kfCr6RScBxpwpUG+X5Gb9aaM
h0V9o8lNrookg37q6c8b7I+zpct0SYezm+RrwxwdgR5LcEeEjTBTNTWZZGRJR6/b
iJrOg079OIOuSqtbMpZrOhWmCO12Ecejjn7MvjDXQfbP9TYNNXzVuQYZbCJ4YTvv
yDUz9JKuNwzZ8yzbaFnVr3tp4sGPqvvdgt64pKUeHPRZRsfRopOSdRlQDWu/fDvr
i8dAils+NsFU/MTZ/l6fkRio3+sj+nt1qCDpJQTjgM8BQTW2r+qstSINsp75SmKM
apspBNeczykk3ZjI1iUdCTMObbbVZapBBbK/Rew1up8KLiNKNTPFU7Srcm9Q8E5w
4zbGTZda7UnzRTNMdf0Q9PO7Q+lw85TPKm35lNFzrFkMJI13WgOZCrhAcKHJbIrg
bKeDXCPtPNZQJkuC61wIrnYwaSEINhSSwA9jskUw3qHFHdtss7uy9qqG/ypygxQi
ph4awj6kYqAQ1NN9P3+Lh78BqfEovty9F9HZGBrTlH+4Og+yRtj+hTCpGFWsdodt
7xXg0tDYiR+cSHWPd/6OWexjpVDn/q2pRQHxy2m5f77AXITtX4bYO3vXsd7yVEWW
r8IqXmryC2vFrc0rmrQQt3ah3jhX9PtHZMaaNjeQcP3rxxSpf14KdUfjZ4+EUux5
ydrlCdkVHOndfmvoVQSrGiXdFtVSJ7WOLGrvefqsaptHXPk35wvdbWk42iM3Myry
XAYrbVv1gjCrFLKO5HILsEsffIt/hcxBLSnSmwRdocIsaDDQu1q/8c7sS+ZUHg/G
mcdz7MfCE1J2Pj/DusEbuJbRK0Ka0f2ipEg4FCPgyxvgO1fQdTcOJuhTomON8GJt
SPGVhWwE646o6dSgakP1AGpjP+Lcn7PYterJMtqaNtMUb+AeZ+VAVHm/xL1Bm8d4
D5KlzM0q2EIoWbJJQLh8hlAXfyHGNvxEpjc3e2DkqkbqepvgBjsUW5s9DVpZIad0
nEaBbFeQIwssCW00yVRetb//W0Rb+xUeQfvJrahiOcmmPuWWyg5F6KlDUEGfosV6
RNoGmBQsouRDjCEYpRwDYr/o7Z8QEDSX9YtE7PVI7l4R/iHAZFqbeAKhFVP2lcEJ
atFdIKKB+acidWg5NiUb8N9D+KcYAoIecCffgloxwMK7lGWhgA9vLso1bHCWLZyq
QO4sySTTmqh3fOlLWcuBixZAs0b+fvXmWc+pwd0z5ibz2dxtwNnFM0iQNr6yr8mX
U6GZvXZxXtR6l9l+FDCFZ5YyaC5aA1SUnV7d2Fyw7SRmnNbzRLbpjhsI2ddoNw1t
mlZoo8au21tptW4iT1qwfxWS4Tnc8hJokAV/AEOqlrxGHxNHogD/JUspYj9PbvH1
LIpzME5h8uEUzitvkmHloTK3RykYUTIraPeULYmhzjX3WAYxTcuwoWEKGMvS0pEv
sUayskZ4kS1tSxcL33W4fAd6rkZQ7+jJbWdHvhWTJEKxJq1DZ96OrW9tD5CbFQVy
I7rIu3VetClW8HRy1uSWqpdmP5HFgaYwLNrdHTA4FyQzOjcGTlKzpHOKLvadfbWZ
r9GGzgUwZbdGEcFZvwDjLLzWX8fqCT6JKYWKZnwwZz4ebIbq9EMdQa2vmiGKKJMi
v6r0PUET/MBSG1J8UsLyOoDRq9rUycbOyRGoiC5v35kg/xwy6GnWarS2RNEsMYG2
Lnz9cujSiJrTwHkxnAObdY8oc/0Lm8nzpUSDcO9Bwsql4N2fL7RLWqJf914eWSTO
W6TcRBZ9ULaf/QW9z6R5M4BuSz4DeCy/jQiGoxFf66iDaKgxdBisPCHHGTUE/3Uv
P7DLq1iTC9CmXMkkRNcbjtbm+L112Y6SGZbHCWzU9hQzhkBxxntZ8FGfps7lMZic
myGVWq7I2kbK3YmI7a9Ap65mLbE2ZzGIqtQsLusxi1hVghusWHBRBKBuwINMScCe
JJFu4M0fQs2cVIfFXkf51jj40JxnSSI6HH5lyav5AEcsuUWwQgwcitZH1DAEF/u4
l3fbgVVAjwMuxN/Tls4Qn6yGDNZDurQzyVVF7IqlfGfCmTZQcMzoB0sToAjrbR0F
JBhJc45BrN/Iotz14IwVZ5NtMu/qfUbUglu4MAu/I8aV5bDCW/L/0jjtIAKrS1xS
x6mt86APq0FLETn/xiWeZoaMbghIa2xv8yZxckpl87muGS4O2ly4P01EhcG/pYX2
XY2QLzIC1TmCWf6GY4OI8RBSchGtgPq9qJ/xBH2sT5P1vpfVdB2Q/78AcueZXCy0
kB1VYg+LXO14kQGdw3Xgc8DCdaIVskyCJ+Zj3/7mPuM5/p7VDY7Wpu/HPo5cNZCD
wvHx8WBVOSFhdNKPmWrbBGI1w5NDlGf8iphGEvBBCPwC2dA5Fdo1Ih8ZbCpozxSp
PQt3Lco+Fit2pWogH8x42Uks6EbOUWSersI8tRYHjOk60NZLkfozT7gt0Las4k4Y
aW4boKTuvHceTJLZQPFwVQ+dC6mYR3Lklshc/pzQ51vnMvXfm52P/2wfLsBiDOum
rCmUjE/6R3byjtK6iRSD/LLtB8j6rkB17Mumi6jQVX+/PwOJS0V7zgKNpjvx6SGa
ZNrFxCT3U8Ov582APmspjxFz7akGGz57ltPtN+aSO2HjiP74bMIR6vdIDZYBz4H6
4nvJEb33eOmBz96lkWfNqmVTmbt2PLdyEmhcZ7Qu6gLqtrKD1o0pA7ZYb41xY8yx
C4V1atoJ1eErQ+XW0KoK6Pi1itSukOp+0k6tlZ3ciFNp3VeJzoFKqjIq/IwzFCLu
eqo0Nc39c7wwzRnmJUkJIgcrBGkY1fCxKeJZiV06t+BqkxbcvHoanBsX4TaVXiFU
W83gbYa6pCjt8a86Zy/nZ2axLEBf6ej9FgdFunfwMkfWdXaHsfdyare8Sr0zQ2mr
jro4ZcngIOrR5e3n3jnwWrQEXuyhHifORVrqsvtm7ZoUOb9oRojtpctP2jfMKjQ3
anOWjxyV7eWR/HXlm2bmuvJXuyehTxYhugxg/0AapjLEAyI2n/GNjiAajeIPrHzD
TFU4b6KhN6vB4s8hRmB5N1oPp34pImGN8ElJLGbjkJOgkegtMjm4O/pc6QYYA9Tb
slDNkjmUnQuonF62DTpNwD+CG5obyPZX9qlauUCMOJ8E2n6AhXFmhHuu9xH4heol
F1kNZXmaHkv4Wh4Jjf889+epwJZQ5/Fug56jCYO5hqmdEB2TwJA7zQRkLVgk4+yO
JSKtSnfsKMqRnB5tuW6j1b15TIPH1MwtU+VuXHvZ3nntwUPqof2Y3DSh4oivOT43
n7Tco5wG1rEJZBvEHaMP14puYmUNyUVgaBiy26HDwpry997IVjx8DvStl4xpCs9Z
HDaANCY0w1RMlm/XNyJUN0Z98cc5WXiYEA3CuFw8xp+ulGJCiN6JIEpbe6yvlHHd
6mRa7oAhCjC62OvL36XPzV/bCYtDInbxi5Yh58pWcUPcIof16fUNejBn6uCWnaxQ
SzQ5jqD3I1tzO9F5pUv2qznExHbhc2F+cX7BQgRG8Cy+v2opb8W/Zc3TNKvqoBLH
yzMp8q9Wx+YAbR2BQKtJl+NH06rghfuaFS5TygM63rLhkBnLGt7PI9pGmpLoPO3c
aqm12CRD2Baenhr88UynLUBkPsEZpvms6LwdAS7kbIuRmtZp1GCMJkQ+zQL7U7G1
RngUlFaoD18eQZA1ZCsz7l/DNTIqHcwnFNaWc+WDhR5a454DB1Zhoa4TckfKB2F/
jBSYtRSSbqn2wlC9chX4PVkdicAcWjpCx37m93xtiRZuLG2ntfiNJLadKTj1Vvjj
zCUu6q84VcCtYykv8uCa5ujnpmPytFW4ufn27qtp803KkfqNHyBR1miU/RyCN5ou
dvsO7wCs3Y48BtiRmDV45KnfIlVQI05G3qftPPBwb6efp7+WSasqUAwY55E1jb7u
cUZNxC03roBhhewR4lAsb6MRL3jgtgWbCyF4X9tzVqaKhUtj+hGFjglQPD557o3A
Kk+DekVOnINTVRTbq4CjWbVwJktx3UlmA7RdwkymsnTFqkZiJzMc8FBLslFg5TK3
1Ndfk46eR11AOXrhR3lNn76lxySQ8VRS3mHbIwOcyWoboFSUefQ5QSKaEv8mA8YY
6ihhmrYW1+OltFe2PikXmUw00lFMbYmK4KcrzIxQAJewE3dAjbLjY2kcXLnMP+3O
TUbLhX6+OJ6Y8txniGzB/5dMiGRXWEjHv34sX8O2VqF3YA9wdDF+OktpYCGfmDNr
PT3SyMJhgvjBwht7/9DwULjdDbTD9dqUhu8Z56YtIGrXJCky42WO1xq039L3ASix
qisN0Vbp7j8a30dGeCNindgm+BdygTq8cHzGC+RD0IDaD3Un9HPMSdFelAZAnSWp
TSH2ae/5RP4yZHWG9K0SpHB8eT8PVEZjx4O3Z/OpknOVwSo+W5a59Hmmfoxq8mrk
DdLaVTz8HR0aKqsWMhHvBBWcMadyMRyIHSAGoQTdbte9r1tX/O6qLv9YCQhluLgu
oHV1Aa2AYWvNn+A2Hq833xQbkCYs5YLauqP/PhVRx6H8/2QXvsewArtozY+vIPbd
UAh5V4c8BuYc27Dk3xhWBJHe9SIWl925uEp4Oyt0QTbydncMzTSQ9pGixyD/+4C1
Uw8vSGJT223nB0O2K3UjcQfZ2CUZ/WDHdBAmWHM/HCEhUZzZqEtPPsqfI9ogDG4j
6V34AhEuhiShUrPZCOOMZpQ0nEIirK0aRaldRcaRabJ7Vu2PDqPerQ1M1dQUGdym
7QTRuKXhoS33yv4HYFa1t2AfgBfCOyFIcgy209YsrhwvcFh3BJ1EQZypPFWRmkhp
jOwOhTf+jKsQ9S5PRudycxaHWSDEFxLyn22mx0JO1RC3/N8mH34SSUunfcbq7TqP
TjQb5N5Cp1tK06LkJPXw0WE6mJs4Ru1aWAO1GUyxd3VvK5Bu+xIaA9l1wEnCo5nR
2l06dHnqEnjHpWfYIJ7JQ7/UvHYAX4OXrk+t/MjlJd9yUHo52wJDB/X7r9VI4I9I
9FoJv1FbOnB92lNgTc8G0k2deFgg5d8+herMuOL7nvZ4QOPHnTsuyuJQc96mDoam
N7e63LfJp4Tx0Vbh/I7/MyDDoqPlRrqN/OBfCN/utWYxJwgWx65mmWjzqeCWf8VK
TfYemIiTHzCAdYQrRhAPz7suIpbeiscycc3r2KuyURCnzSNAB6BQnrLp29aGUCi1
T+p0bNWPONWAVyoE23AkDAai7iCuNAI7EHFko2Uo8wMkhl6W3oa0Vcg++CTh1L46
uvBEFQFywIdt0su23D9yCOZEx9XpfIZApLYavrz6kNkDtZnWPzyTIENkYIzZlJY+
GO8VG3BAbo5ZdAjYVojWXdkuSI/8m6xTgStYPVAJZBGbG3hUfsGQ2vfAZ3KTFJkN
astwL6BfXMm139tEnyHvfuMr3fP1bk+TCygG9etkpU87tXXspWpyX7kjDsK+Q/Zn
w2hG4HKb9JzPXZttvit3esFOMft6rJfB5h3yxWqY+5qOC79pmTP86pdcbGtWwXOH
Kuby1Qv8WGM/OfvqO05Fk5bq4OdQSZ2A8HYhFFHNhnaM97O648AVu5pzr+MHbnnl
B2QaqPnplBX/UiINR1mCiAz7VUej++wky6lhXVcYhP2EcpMgTLfzB9OopAVrZDzU
ly5t5xEL/X7/8yP0BTFC9J50y1NIc5HLKKdUXihI9Z8lNZca4oHHuZNr2izkdzGi
sPyqRnlF4Puk21qLCLP+TCZDjmMDU2PfcL+A6WWFJ8pHQcE76hUx49q3q5hNxLs2
uizSbZjfwQ2rDtqYqlKoJ7H4VyhaqasMdrau7Rcpe7Q0y8vhjbsn6MVBnLqm1x0T
0CnO8C4AepCxEQRRExJJGMdgniWDXsZdyoSN759Xl/1Bd3ahlrBrW/NCKuwQW2Kt
EvcIgyWMBd0/PyZWBtQ/tPeYc7KWEzHKH1XxG7t1kif9HGGTrqXizh5XsdsQwa4x
vOy0mqqEd5Z80MUKFw88umZENIjME2Qd+EVs89Lh8v6I7/nTt6u3Tz2QXtAzI0mc
BUTWyIkgpquDHr3H3ZdqKxw4JShJ7hC8ImAmMGy8x9OIh/AUn52EXPgtbuXv9GPW
4neDfZaMaVNKQJlL4c5W8ocDqeBOxTJFsIu7LasWnD+JEV+IhDJycja6YOw6xJWd
lmBu+7XJ07x01+J2gePKReFLHF6E/TVYSu2ay5Dgof5wnH7xkfZXUdfyViIqaO+N
IRkSMm2u2ozqyDE4Q8RqVCsvzQy8F7312CP4j04b8TX9rJLD8OfAZLX2MS/2ayOW
gGcCzDKk5HvhS8brLig+Z5BSXYHboDheTwbvfwR2t29v1wRNzuTBZeXwybnhVKMx
rYxK7CvkMnWnfQetLhYmwH0ORHsYN9xvYRQkqYKWg8Xpdu2VnB/2Z8neMQ0k1ASc
qYPj1QjkSxWpd/5NKLJHxmBi8ZB1Mo3emXFsWFFfikuGS6fq0MY9bvyGP6ld9qMM
L0DKPAQ6Jt+AfX5BctPD+NEqcS02R+FxWKlLbZyqdf2mxxnQuQPeg3la+4MDlxea
pcLl1cTIftxiV0m/vOmqo44W15MEr+rTcSGmQsjt9mogeJGc8avt/ws2apJj3NXF
SCzXEueKIWFnGFItDUq42UJLZBXstdWVFK1cCd9ubkZJzb2WObSfzk4XUfnzIx7+
PEks23f3080d9mzQrP7ZzeShu5Ll90QqHkZ8R/3oi0Ym4BsQ59STodxZ5j1dOyJr
UZ7zck7l13+Qun5vHLWi8ejvFsCZLul21vB2qFPa2wLdlxHB3mxvpv4xsV03bjWL
WrGwWFHWQ8I+aG3R416TlQGjCJdmyIltaIWjT09FhLjXwcdmDSrCNxNym29+gj09
kT0Xl8ZilS5B8I9pjq3+N21KI/9l5Y63419ObilrCK7YEVxYc6JN18vOVz5TcQeW
4oDyBjgvgKzS6I8kSxQeCn5Tb4peiZEExCO6nHHXeeeAWXduRK3uXMJBWcfHf4yT
RvIObjSW1Mb0yHUbJOkq2d3MthGlqhckr7UUueuz/D8rdqfdPEnRBNlJuObDVg8y
aAv579mbeDL5yEseBkL1iCKGbtSGI0bf6BQQHZ7hdnITAYN7g1W9hI7Wy96GRXjN
EF8KX5g6kiJmY+rakGkP9M0gAUljw/2dW4D6A5btTPNJLXwMJMp0xqfD3W6qIpnb
DRsd5+zd8DPzGvp+26GOb8fP1zOZWiJzqDlOKpDmjE5zWN+q3irGj7IP0iIRjAt8
ClWdy++hJWuqASpdh/9OAwvn4STZ6H83jECwsMD/HX8O5NCTTtKD52mH78Lf4bhR
x2Xw6kuFYHktm9+TwAam356VdMj8+V83+Junqw1doogrgoeCuBKmemIQJFVSQqTP
rMryviYCY1++AWRmzh0TSiryH8YGC8Or4RHdvF+tYWlPvZ7bDTppeWt7Hz5mGIBS
9yiA00FpYRU0Y48aOZ8k4zc55MkTM4+Ou2Kz4eT1YNOlzoE2VT67X0LKq9adJUsx
GAfm/w4SVe2PxTWN0H7/AX6ZNA9c39/FFdiu3H4ABevp3+fnZjuq5gfYFRLqW7UL
nPW3nXCajdzgBvaLj+N39+mWInVQSB/NpqUEAPn1se8w0OVZZF1rk6y+eAZRdRgc
YRyzaYi5OV2Tf6NHNzZ9ldQC1js46c/t5vs40PqwhljInM8VzaPwJoX2Bxcm+2qE
qFdwWZ0/pAZ5IOW099sPV0BG+gdOU6ASQdGPehK7bU01Tm63ACC7ijsJVIWlImID
STffcIovr3BrjarZYUxCmuDDj0+gQIY76huQY01PUdX5H/ateQw6Egj1km3G7LX9
vVmlA/PFx5D6OmZqUeUOzNNUBZFJa1+VLlJsK/Ygguyo1yLMO5QPlRjrpNJ/X8wi
Q0gpVQ5aBt1PD/vHcgUNVoHHoXq5R42dnrt7ote/O//j9y/AMcciJ6vRU5WTbGzj
o9j4bbHw7GyjgLDvjH8s/5521dpYKRKcNAWTwa9/TL38MnpMucuZgtRBlL2XQmdU
kl4HidHFZO8w4pAP7/8hIV5es809er0a7hkke7J6ZDeTaiQsEgLF12WsUCttAYw6
Rn53n2h2TBl1cOs+U4RWX2r55xYXra5e0uII/v4UbbFsw5myKEDVDud6tSFiFrJR
6mSH15CfeszenpAYhpIHYWrysGSqKTlzRTUn4xbTwCcIKz55ObTntkVlG5BAb73y
z5Evi03xWFNqf7SF4NRJAuKWjMZCFtoIuoyT+oS5nL2rd45GJnonydioUDXl6WfS
qhcODC7Z0TRip72O3A0xCjq0XuNpWDC+0pSmJ6j+JpiIaEaBPTnIVFssQAO8Hapy
9Y74GmnAsQPAJOJZ7CedAWoqKOMD4T9RiRaOrncn9CS1x5NfcSf2Duq0yNiAs/I0
V7TyH0Lg60CChK9PPMP3vFs8H6QgeJJPItRo51vpDWEoB9dH1nBJZeL3mD6tk2LN
wEyqTtVAv/4XBDGvf7PlAW2eGYEmdsifOudWGW38cexA6szJ23jS4U5VRcIH7tql
60jz5vziAHsk4FUxeFEneIfbGnZWNqy6Jx8JgqqFmiyH1yAiLOIBYPv3PShhKoSx
YGqBODdQt422wIU5xqFcjQnvDqqhxN/vilvTXI1PLB4Akd0VORnzLRynYkDyBc2X
8Cp+Q1wmp9xteL0YvwQ0rKC1LnLr889K/ZwGq0QiNq5tbFV3a60mtMhUQeNyaXhd
Z8hIXrXD+NkA4t8oy+QtPvRlvf8zxHtu1dpnE306d0mAHaZ+UZXMw6omX+3ZnemY
DT/Af2PcjThLK7znUooJzepsY8bL/I1m8KRBCWpGzdihNiRjrBISeZQAxuVrJ/dv
hHn8zYN21MRCZtGNgi0vhDcQUbWJv8h7sJgHpMyGI30HAb9bW4F/0JsmleULwnY8
TtEmV7W7i1HjoaPTs26tCyEbxPwVp7HLadAe5Mzm5LFm6BdajXWgB8k5ch3FhI/p
NdKXJE3u4nFi8HLc/TxC+yVb0ugLtUzncONfT4UJgAsE8EfJfGcwi7hEkI29I6Sw
z4aLKycT3PCxvzIypFgz8dKKmpw7SqU9iNJgQ3o2lb8f8LUv/BTpuz3vOIAK+y/R
MjUNCs+thEPiYsPjoC+ZsgbChjg0pnIRQ7t0K4yRZMyNh722XscsUFVkIpguixz3
e9SlRSBVCBmpYMKP5lmc9FzLUwwGtmd3YIu9dny5Bu/jo0sJNpoRvwbPhFGp3UjN
83hAH1OHmuRT8x+BXGfFN7EttrGqTfMO9rk9hFurscm7ilMMURCWSNkxoUIP3e8v
f01oOX/AVv+oipIldsGy3tGRbX+zipDd5ht6o/b1SFfmM1VOYF26M/dndLaNYRxk
Ch1CAS+jZlM9G+u0Mb6tsKWbz8XsqczAh0LRpGUvppOZ1vTbXkBMZ2Lx/FpIz85U
kOosnCV5ht0jjUFDvjuDgne3pd4IVlCiNKNGdM1tmZKQT8KpYC+Kt98Jf5krxe8N
NWPL+P2AgghWWJM1CzYpLahfnNEe7Huz8l8Hd58O9a14mmPyka4dt/6+JnlmyPZr
9rXnalsi67Oi66ECEmJvJJoYVjo2hP3nrfREvQBD8B0o7T0TMCUmI0suhj+MIU9f
HJ1szRJC+fMh+toddwFeWN87j1VzWvL7lpoHsFeV8UB5y3nelb5HwLK+A7ugqXQ5
5BDVKbFXVXR6GdLefGZGaSLrNRVOT0ps2CNp5pc3hzu7OWdwgbhVJ7A/s9FMRlmq
d/W/9gcwIlOI3Jkoqvv926mvWRFwzBxHA/k08sNVBSofmwSSelyF5tT/UzwPM+MM
nVm9TWElMKUTZR5cP2iLG9bofDbbjsDmWk6qb8h8kFwpZJYdZdrJPe6SBT1RqmfX
cV0rj146i/jq3DbWmpDt7KaaqD2u3ooR6dHTYh31Ce7rykumRiZqKvHLT6pwI2FX
m4bkiif1RPd815dxaE8k03I3kmO10aXivwjnD5cDn8VS83vC1C0TKu4gKULOqyzE
N56C5O4LgFMxh8IPKFEnrQIJgRzAlCshuIKwhwjWF08Y+aHP0wKe5KqnjphZv8Ev
HS5XK8Uy5cf9SSJOhNMVZZJAOwmK/sGDyst5Dp99tj3rltcSwbuoJxOZ2tLgizsP
EWnOQ71faxfEjKEFHNbWkP1YC+Gy6/R3yB2uxJ2bzkK7uLATcRStEK/98TKRpiMC
lCsqdYhWJRnhAsEBnVWABUe0EXEGlFtdOznQupZeLfSsRfywOq0B6FTQSubluSbb
dIYsy1ooBB7BRpwFMEoTGi+VUi2OMwdbkTnOsbXVzIKvbhjiTItANl29IZXfripR
Gk2DEn9kw5YO3ymVKjZklkz5j0gcEZFJLd3wuHWErqu9dVat5/EeLi0NHVPtfCLh
Y0PSeH4+muO61cUIQvzWehyJS3qzZK2tMhi2JfSasOPOgXHebv9oFX/cJaz6Fim4
l59cNUWb8X5Mlw0oN8lY7cqpivTffsqE4SzTvUVcT6PhkSt3UJsXkvrOgSLXAPC/
Se0zrMvieEetU0/LUbAONaJYXXJAS2DpON64aQNr+Fa/yBxI8lBVKyy+hGVgMb8+
mBWFjwIkbtF44+dwBz5xA0MpuWQZwbYkYpgBNxsHshH9rYzZXRSRs8qtCg902yBA
6vYfNJJZU2g/EkL0e5x47MFKR+rilaNZBdmt10EQl9I1iAFlj7ZXj+Dv9PP1whQi
Lqcao3Bh9exi9UPIVxhmAUUZTOJmdd4EtR2KvzXo+zBe/TLHCkVcUVQI5ak08KnS
ZYEHQ3heqnUCxhzwEmQ4av7ka+lKNAQzXoYrz1jnj2ykfoGOS5QzB3vg7k5j3Nh7
KLPTjBL+oDi0vfQjZ5iVo2loFqMNbaGcgt85AJ6d0E8Rwc5euR2CQcG5rr5GCSOi
6rXTGN3s+iUdEIRS3TvpfZ9L8FGgAc/VFQydOEDCOogVXS92SetGt9SGyj52CgTE
uxsfHvrF5kKvIdCUX6RQrnDwsWRrTYThUqndX0JP3eKxNRhB3eN0so4CnMd4ue4g
AbqxM4WutS2XtQ/29NdJGblPksS+aoUa6j8/hj2v1CQKiAjzQpprhUx/k508Ezzw
12jtRSGYvGojr5cZC1rqyvyGRTKABfHSglZy7FEQTk2KEZ4OIb6SxWfnDv0r6cHt
9VlRiNjZb2+d+vm0Xha7ZEUd61xVr17nqmKWwT2SBNcwW7149qF4oRGz4uZQP4d0
5AW0RS+xa6gq9fW+UNEUsw3tkMWypPK/HQ5zBBelbwBS0rPRn9mP8i7jGkm9epPy
enkOXRza195hivSiOVToY6Vkqe1+2rRWaVAxxi5JfD5tVO93spshEvBglBqOmoXk
A9W55fcOchlpkhHiAu+wduVqmTcas6+Iko3cPwrVR+7A7dpRgvymg2n+N2X71int
9Wmg7QZcI+ErKUVqE86cZXxOBaG12N8oXBWVhiJ4cqGZ4ByOvbGE+yNfn8CmwWzt
YuBzOATB4fvh+Rlk5kNrHAWwz5+n1YNc2e5Gk1cPExRDHy+Q+rtsiVc8t2lWohMr
Z0mpSMvbR8+8DXA4+G20gavBvszXL8ABoW3h1r8G0GFnK67LjrJvXxv5xWehofTc
fCtz8mJCjYsU/WdSr/ve+HWlHCcg6Td1+2tM/iO721hlBOxEwUlTBKq+zjoUYi7Y
D5/SqrqMbN3nSGqteMZv2rv6TtVFwOMHqmvQ4CtiNFDXGiPWfqUOMMBXbIKZ+IDJ
EXQCPoUPqsK6L05rxLguCqy5++QafVdcQF21xpjWhR8sEF4DDQV+QV4MiZAX91Uk
B8+tuKkls+rs/1TsXkjuLTx4SiYDSy1WymReOV5nR2ZooL016SDl/bewUfygwDLM
iJkXX+eU0a7WwOc6os86iKrZzPqu1cFb3Lg23L2zgdmkUDpvXmCT4DesNinND65m
YlNIiShBPTquZWu0C4ScUZVzdvQlEaFj7Tc318fYpAoypIV/kTH77sRSXG4+l6U0
8IE9cjeHisD7HK22CaqghXyLWtGTQivATWK18P0MyA2n45BXhZLFOqeqKV56hrtO
qIVblqSlQLh2zYFo80Wg6UjulBRvnJqKUXC26n6+9s26gc2X0S19LQ79joapYl/j
ucnyRSZ/l84OYEEYOjAAI395PU8SA1b2xeeSuVwiK1D0WOB2YXxiR49TDFuyUEaR
jsRlG7rIzDoIcO8NnF0Yx0/+xj+MlbgZAsrQOsnhqvJHjWoEDAlq/MGx1VygzRom
ZakKmA7XwwCnpbuDPyIeps+uotWnqUu41BzxhICSFqj2iP+OEYavBJq5wb+Rwfbd
Gd7UujeMcQ5ewRkCGKw6G8FGBpzBziA9aITfqMUZ64y55X12zKrfKTwQza4oZdda
4W+ShNshKqaUEb7C4lmd7U5RC5XaKkrlgOggwuQF5chgQ+HJhgU9yhB8pJvO9P7H
GgLzfa6WIR8EzT3MXAACQ7kuvmezzJGdJLrQv61xteZc9FbN9NCaDSd7+s+p5mX+
hoLeO0PdYQwGdBnDoknxj5PbP0FwSZsejkT2j5Sc71aXbN7zvMazYcZ++sOPWsfu
FDL2AwBuV4++erfYjtNTKnnbClSQ6SCz3bpQem36+ytBWclAI4t8vy1ZcbeLhqlt
WE+hlqFK/DUsJvweHqL3rvWlvn6kus3HUCvMGXZFNEW4LZ958IWg0S2f0OLwiEF1
zXRHRwzKeSp4ZObCS+R1PLGmbAILBQNIx5SKpy2nmdG+06ci7XoFM0wp75+jbvhj
PHXA0/l7brvk5PM7naCvlvdVP1GSEZlf6ATaQcYeBeZgKbWLLKaSERBSSuChwMEz
7WzLNZ7Qza4VBAOgsdlbSw68jNsP1dtZTgDG1atipNAWP5xMRFrge6LXbxEGYQCq
HeDZHNints0L6/OsDZLprCkKrAh0TSb3wArtMwY4qeYPqfDAYwIPFZZZkzAdSQat
eX1V0TAt/SrPMzNxEGco1bL+uraAvhb4FGiGT3KksfirkklxkvF1KGkLw6vx+8nv
fgqpiPY/gBG4HlQsS/odurLuo9OTMQQM4EFYNeSahGFMfUtfA3XFVleMR7Bz0mny
FxsU1aChqQKMCBBYcRhFgjEunXNBB/Cp7VUgQYV95xlq+QhvgfQOXz0l2n6Shq/v
5gvI/mAvsaZIT1NsQ29Wnp+y4IhGCqi2A5mr+rTvCrkFwJfX8u2Btd3+yJ7fNrxu
wvnEWyiyNobnqDKKfkLNa4q3bsyyED38hkgA5e700OKnzWisZdszf7QnqqPbuhMn
kOz1ZrFtoT8YBHjIpKv535gTLOuqO3AMuBsEWN0p083hb4sMm3DaWVaKt6/NAUq+
P84Uq566CCp5uIpawU/Am4FN4LiQfVNK+74I6Axg52QcQ7G8nULNZNOypoS1sauG
lq12bjI1pr8JeISG03eI0N8kYNukTZPakGTIswTc8iFlVYsc9nS6IoGKtZtGBkw2
1H87Pgk/MVQGG0C+vIiyP4Na99oMlIPVDBkhBGaIrFopi7Aic9CnyDHNiY2ZNtAK
KZsd77VZna9mE3OPcTu70rn8j+wV6Q6sWEXCKSsfA3qdGXOhfbuV4PsfUfgQ7xBy
dBPsEEafAj7aycfP4gfA6BmYmJYddSsuASxTtPuAYPoRRSvbAyoiatnEtTTCBuSg
GknA5pFHqAAUlnBRQIJRU1tZbiCvMIxid9fr0aL47Z5v1tzp/+mYE8vgIfY/CF8y
wQSFhEkKGRjNfxn55QYtSoq2vVdovP/t9JrgpN5LRMTDVCcmlSE/y5ITX0h4nV+a
Nti1Bn59/2et41dbeAIkgZtqhwyWc4okXYRsLWDoKZVunHqntJ/fuDs9vU3HB1Sw
VZ7KBA9H8Nlju7YuNjw5QB7SBmNlAPpgvQX/SetLomrnVc2M2Ylp+pzkl/KJ+sdl
DVfLUGXdhQEVP3nVmS0KCWhSI3M0Xz5cgcHmix7iGC2l2mIPgd/BRrYajxtRfMb/
ii5Et7BbEaQSVAGm42ssChyWqFcnzyNEgMODIXSYY5u2V1rXHpNJWMItPzAFyO0I
xmV3/71wXbUrEiQI977FPuCI7yL9/EI6EM0n3Dm+o5uWtEQNVa2UC1ipnu3fiXu9
mbHWAmsqMJ5X54h6EuMMPMda+eRnF56VyExEQ0FJ8j5BjBlnVQu/YqQ4ATx9CXYl
8XsLKWN4gjq8P+1ps5FK5gh3s9UF+2GO0gPgVFt/kWPx6dLzFBl7DKYbL56jW/o/
GA+hZROTmv4lWxNAzh4jtqF+07JVxgt4k8LNsITt83iCl5YzgNHGJeIK0E2LrZTz
8UWHuZxYsQYI+ZimUzluZfSpfE40uHCMKP+BZpbBL+xp+kX2jIIGHGIvgHnbji5+
OjooylAYMSsSbR71I2KYXDuV+SA8CVVdVEFuxYJBfL0Cp5CrhK7zvx5d4B1dbla8
ZmVJ4Nqk2OnNpi35k42R0raeKjbtcweUxHdV89X3QZ2ahHvp1xU3UwbgNEugca6H
tkZEk3imaVC6WICeR01h3diQmHzjp5Gm9CTSWz9hplzCSew2ydokPBedl9xgr5aD
+Ts3fcvfCY1dxGu1BksotY/7wTZ7BvJXlHK/dwhODQEFtdUOP98wN2F/Zb5GMlOB
qc3BUQ1ysi8jHGThu6nJm1IogrNkkpWL3ZbIZT51j8QKO6dY6ogWBhsYwFB4I4A/
e97ulHM+qzB2IYdtHqeIOw7r2Ex7jgGjEpvEcwlGVLoIWuFVbUETpTw4i1bNazEb
wlcYohCoiDceNNShmqKjE6BD8lNetXUkQoQ2xSz4XfwvO+mXsZK7MmavVT02X7/p
/er5MKxwnI68ErbIEV4BEYBXx95x2FK6yOnWFFGig/dn1myAUNrYeNjb9iyGPkBq
JD94JJq5+S42a3fEyZZDhrtVRwwBbH84cCsU3+vh+A9GpjuG2ogryy91Kv5WSIOv
8IqqC+qVq+S34tp0qQrmg2qxacYlRYEAfuh9BzX14iER/arXVOFZWCi2NmOQLiQT
HcDr266v2vM+4u6ff+VRaUthq68Q3C+2czRmHv/xY5jhRmIobMl/tp1x6ZJkGBmJ
x8RH98oeV9lE/0e+FnoWNX2TPmKMZzyPbOzFP0V1BAAdQ1YAdMV4oipfiGTkNgQN
z0TAmiDIm3L4U0WRxH39tBGvwedjthrFkv/Kd3BVQTe5jaECeqxzS03OyEEHYqSr
GiJCSzE8puxek8mkH82BZidXo47Tgq/JIs/NWwWMpaUerGQ8mmq2K6QLZqdjsbjC
phQas7hexYHVIzXuwkZdKxQRIcnwcJSjcwtJGU7075GYIPK3K4IidrU8E+A8Woi/
fyH64sJHFT5880BKRKhY8pTnbYtwnPO4jUgp0yMuFqX8m8v2MZu5py5WAqKGmfYl
nCRX4dIiG1XZ3Fo1N7ZwLNNUnH1m3Itl5P8SxA78kV01kNAYrzHsnQuuwEJ5MdQj
66vd6o97MEq+3jbdPxEJubLCpvhkv97UGdr2QZOOlpDdFAfuGrEH7K/znNCK1QkU
DQMWIfkrdSMlxSz8At1ytC8GMIgmmfQsSPH8yI8c6C7YLqTLINrZpZxoSJTocghA
Od43KcgC6lWrfZjP7TWg1c4QQxNvMuDJiWZBY7RgXgoMnaY0CBYmDbM0Q34RBCjT
AHpe5e7Thh2DFZaQrDh2WS3ZPBFIvBJELOCUe5FtV+eEu7TBOqb105yijEXRuDJ6
r5/5z4CXMLl3c3enJ3dFT4hkkNvbJbvf6W0F54xLhDF2G3JJ6+I0xpahX2ia+He0
o0R4BbEQ7AqRCVdlUc72kV1+Maml3lDklRHm4TZfc9XgG6hD7nxx8R2e9Tu54HPD
LtnGPd7XW2PjVyNENd7FNhVvREUa1W51GphboS57xnVtjIlyIvQBZlh1MjVKttb5
cW6JGgmrlku5f26gGnxh3PMPuMtzHLgluUrBFp+IIfO8we7LVmp4+z3n4fzYDb1R
ddVye31EmFhBLVvZ3E7Yk9uLugHREGmBZPkY/Yq+vfryCtoyHxj1cY+Vv/xbWW+N
D8Hs78d/FM9JTwNv7BnFudV1f4nrU4RvRxkzKUd6FCMw2JoIeqgmM5VfUPMG5DVb
iCbysssmNJaFrCqWCZ4z/a8mv8YorZk6HDY7EzC/bC7ISKuXEM0jWjubqSmU7DTl
ve4XM/VbiUVs/Ks+6JPObI4Y4A1zMBSbLuw8rKUslcVhHSh8xf94FN+PH47QgusE
nvG7Q0TIpF0iDhAqmmZxqhblHd+XYUygNj+8Vgixc5Mx5HuhIqSxQ0b9IztOWCj4
+SV7L6snPbUfzl23hhNUb410YIebuYRU3bvtK0VKmp+UWyS71cN7D6qfP+yQm5bM
vr6WYnmPkDB7WaKIDrUfvATxRkAoH7387s8f01Zm1IV1bvCkng0oGq5rwak/9DTS
CR4yminUbRNnfDFXl/zt4Po3e/4AAtG1rAkxgF7uGMxiNcVzZplemSoRMx/87+9V
37jHOx+AgWRAKsiSQLztN6Ulo7dnzR+9rh/XbjvjNTsJiAih2mkCWzVfF+koaUzc
qXfPXG/I5pf5imoikiEE7r1HvQyfv1IbBLggsy66K4IOXstrlkn6FvqLn889V16s
6KTZhPskWes9OCxZ72M49rqajbFpYRR8aFty/5uyzNbw4R1vLK69j563cw/lKvFw
AHaTTdxzntx3CL+Mfoz5obw+zdbsXVl09ZjdhdAvTtHPJs2KN/FCQYs1DTi/OSH8
ZlM4tDx4zmn3BLfwPZUx38CwHtpRHKCmvxSPXsxmtD5b7vudfuc0xv3WnUw5TCrf
nGfy7LtDsPaZDPjh4KqFe60YXwsAGzGzkLamwFhoearGcGfteZL5ZImh/Z7lr+gw
1tWyiND9ZH0fY4kplHmhJttUoWS9BpWk8CjIaio2lcXz6U0+n71uOVerbTyO/hcC
/aWsKj4yR93SeUhw86oh4+NUd8NY0h9Mq7Z/BdHXFH01/7EUI9c3AfjTuWrS3f9a
Ub4PZMPFSIxJEV8p8GjR8eS03e4Tih1kIfHT+rV9gcyGNYo2vLK4bM6FdVHEXYKt
AwucoWnUgnKaYRw/pdxIXMjj/eIXPesGmqaZmKORj6MWSKMt5hTwZMAleE4XtC00
20EXRNPe5RUUep/B3NmrO0HKqPV2a9mxSZ+zBLLduv8NaJF0IEYatKoYI4Yqs4t8
HMyQ/JaJKU7pY4Pi8YNRCXbfq8LXAYKxLenpVHxZnixuAijL+tTSc5xPxyshxRqP
m+fz+9hTxtIEi2SMcrjNc/M7B9YObnJT5wCH3s9Obstd6dKiSjtWO8ZAueUqCS1/
CXwdKeSnYEFBC3GZVLCd4dMZbDmjUzJIH41ZuV/FJ7CdV0wGniXdT6DYr3bOd0kF
EMzlmLg06fuChZwRHqqwaF3WdGeFgCXPukT5ZpL+nk7ixAkslNcWdF/hrSYlXWZl
pe2h5dl675512vjrNAK4YX2lOCQefcA/9xAUwDPAEC0pXEQDeeNqfbBgK9Tki9id
atgzUewo80mvxARuODF7k0ePNLFySjF+tQuJkwwbLhNVPih7o9hcwFg2fczcLTko
W0p/112JP+BScg61BZyMau6190VPo+ws/h5yOpvbeHNMyBVV8m8jt53gL4F3PEsT
RtIQ+EFnQHmf5L7mR4CCt9ubjIUS95NSGHXPnXa+XHIGJ+sV8vcw7ACjkhDQUOSk
wxMrK6bUToU15T5Htosqp5jGGXSVWseTyi/yJ8joi2da6n5vDmdnBYqZacpLqoxz
nha3lr4uYpA9R2nATYTqDiQYMOdd76dic7ByNzfJSSXsQWQAwhHWDekxxPSO5zHE
efkJz5vXOZ8dzmWPxXqhFiCFFwKt87d4Pnp5M1YXanF18ZmxQOn6vICAaZIL3Ul9
bqkdun1rX7WAQhOi5LdXQ2CNRXy4P+O1E6NVS2nsZEiirZKQjbVEaY0nCL3uNOnS
S0kJuHonyq7oLtS7uYmsNCj7UczoBWHnskH4EIMWbQro874a0/5iHqP6z92ONYDl
B8CpxlyEovQLm2XJ1n1uSviXwLZrhGWHiu2K3LGvRW3tyTyAX0mD8rPT+zJdKf/y
9Tp0OqVOK1S2glA92OZ6b+e1scn/iiy2P50/LXhu21rqDMITGeaMGz1oxTwEdRG3
xoSsEYzp7uNUVHvpbMcNZTVwPrHebklOM4dPfNUBBXcw20M5wtBNopOJfLbLr6Mp
48yMm3gKXMh+gkoJyFC31i772xvEg1mebvkrqYvZ/iFlH5ZkZ9cf5M9FKvikBfBO
iNXk9Kkmu3vxnrdvp04d5zHCs//Ar5OCt4A6f19RdwI+t0j278DSevTKR3TP2CjK
umU3ZUFhnE9RPaQQ/xfp6aYTsYhDBCpfC5QldhyHOEP+fWkk9YufWPYG7zDziGCo
5cT2T7UfrlGTrN+Ui+5ChnMVriyonxumCQ/0K90Qxnk8Mwp28MWGr+chj23KoFmh
JpTCsFuf7F3hfKLslKuyW88o6gOR+pMarMou0ISdiMiXiFQojtoqqDXwSptQqhhQ
i5ceZ3MiB9J3Lop6gM5kdEvbDAZycnPzRspRgoyiqvuV+tMGQaLLycmSMs3gu6xy
2KHT81+haY8Xhtub+JSL4JDFW1aOrjMoNLXgyK8qHnL9LXAuNiiP3U0bUY22ybrR
4ND4X2Srydw7Wi6lC0ONIuRazhsUMSOL0gNT6tjLCaiSkHQwy/9Db8kq19hemVRz
WHzyS8Iy0gMu9ujQLw7pj3+a3Nn2xT9fUTmrZm06a9pOo1f6SX+GvyvjAGC3Mwv9
1dpA2adQ9QkDz/Iykaa23X/cVqfEZsOfnkvS0+O7DDplzM55XE2NuRWlKH9m1dQS
wzHkam0hnvWNOmzpBkTIURndX1EtO3IJ+7uEtr46NbmVAe1n4RN8ZqdS1KUMB3+U
1JCx98GD+OnRcGZslb2pVoIUJGHVLJi/ts/D+lNnhWSUQjzkvI26ql5aOzGkQcqu
WQ4jlkC7t/axfyQmqjlKpI4mQ4WA/nx4QGXBDIL9vTPoWECUGSa3yHYj2fXay/aG
j+/qiwqRwnBcfdC0SZdv1yPd5JdkvRSo6rSMr3QAFUI6FCnL3NoWc9REMpOjrFuT
a1ARvo8Czm08mPNzLjsk/7QvasjxI6h7z3n3UEfmrneXn2zFLYLHiZBP1j9Jsnmr
nEppoQDFqIqMkCMBtOI+af3J62MB8ON70WFlzM+8yAynIx23wWe2CQg0DCvAm9Hk
c0a3xcZyHzTFWPf2YRH73dv2w38e6BgbptLK8/UNqSxgLzV9npopa9FoSkr/2/He
rJe1wmM4IEQtH9ywQHmYYIfzxnwfmJR+Dt7dPwGXotlO8eqY0al0AUv8lsdZ7ciI
BVd23KUAnP32hNYBGhABVSXQ//e+BXoy7/y/1dSwh4lc0xAkztV5ay3fR7G581IV
/TJeKXoHgCKKpuUyOYj6qhYSyEPuCvW0Y3ix52o29bPmha5nHZWujvnataUqG0nO
IEwqF0A7vVOJhXG10R7w+OIrGcOZAzWejmb7Jf2GmRxBxCFpDkvS9BMHwotQPIQE
y/tiPW0SKcqlU0tNqgWEyqmmp7Xu766rYPNBlkqjS8pllVz6YsJjekpenM7YSSYt
rN8rSM36EcBX5xiXRN+rueGOFf2/3X32HPl7YVybjpFxvmRwuTa3i/qDn3FW8D40
MLU5JQEyEkIwlmJqqBu4xxAE4W9ZO6wuK9sm5NsesvEJg7+56g4R1h0X++clU2RS
4dlHOtrgBucJ0cIks/MidIwGEXwW7kgk6aD8ku+xySbzHlz9s2HFkd9vQONefSlG
OoSwRS5lr7r2F8jynXrAohOV2DO4tp5PS8YUE7tPziLkJYRhrcuMh/7xldd0EhlS
f0gHxYOkXF6SHUQv9MU23ll2IzqrlRwZqh73LnXnTQmbUawTbSqJMHZJG5IFbgfT
tENZXtx+guHqLd+sE2dwdyPpZkdMleOOnGfARkyqQIhdqswbU3Rw/hHqziCpuQ99
iOXNJUOnf1F7Ps67cLDgBXj0yzs2rjzCscbyl39YomPNxwJojA/ldsHpj8kqPoJh
0FASxjLFd2DiqiCLjBSdJI/cOnM7VgiZzRkpeDGi1jx/tyOmUqJLV1+OdxkDv7XL
5M/VYp1k5wZ6LJFHrrr7vLqpBqgu6GDA2++VfaNCc8HMkpDenmkOSqniuI8229Y1
BsmPpR2NojwXMvTLyZfEjc6hl1kWnua0/aQRDf+pYcei4D1y9aO9VjdT+wIPKik/
MDI24/vUyfTDhp4aZkT44nXWHcH4HWfb9Ga87iau9Aor5zDEIJm1r83X4dhcIpiz
uNF8btmrL+81Az7xvnVYEq9yxHrAVMA66Utgsw/ZDid/bJG5RAtqL3291tc+4Bcv
XrSRHzFQlCc+4UGafpYyeYPeXpnV66Y4Xn8Yeb8gxHF0qy3efsexTbSlMwrEB+ka
oMXKVLI83SQhHFfNKyxFDsDJmfsR8YEGxk0pGx/3nXZfusaqqIx2jD/1GZW5UtGr
x6yqXz7NU2LXrXBi8mhplGLIbS6fsKbonjXiQQhXe3L2OoqoxaEg1AXwGjjNjDeN
ENufv2eWDYX5rGVOiXr6q1UqVZdj3/kZ5PRwISjV6CtVXdSx18a/rBkgmxvwtPHr
Yw7IBq61yR4cjHA+Na0kQvxu3PqS86rVBILCpEXFgcDjMctQ5gywIlbx0utoah2d
uBz0801ApMRSjRZrirOxlMDe1heyBclygkSd+NIx2VzGN/Jb/TztCYYIU2E3WjzK
7UVAAW+HuEGcAlv7fA6uwIW3kXFsYNgkTFwn/NWNwuBkvXg0XboFlTEl9Etl4Lwg
izui8CMO34qj1AhZX2ko1g+IBmcfumB5LnGKny4lBHj6idLVf+75G7hw94j0f8b6
UB/PcEL6KTtHyHqtHk0PuzbQrsyZQaF1XSBbGrrDa7SpmJTakXf5MHiUP1FQCQm5
iMAe6eDmYzPfk6hyY0sy4zARPFPz/iyfA7eEgKSckgzCm46ZHvcoQoY9iwU4bUks
vyYGMHh1faMXhv0l26CloIlUY2Rug/mQynskRziet3hfrbRO9gGcjcF1eSm//ZrL
LDMc2HFwyYzuKTK8u+9VduNvr3itZXUJp+Uufh7IUoWfHo0va+QENns9TXdxmuKq
zdmKzsfty1PAh0WZj+2gf7TfIVHwhGxbEB15nTL6z0vij4ScT59N+I4V34+/E03p
nWZ/p8t20VtHgYqAW8RLjl2I8mYhQ5EEGENcQ8i3Zqs+F6pnQyPrq5z2tk52v3hP
8d8l2XmST8HoM2ov786KxR5GS1pDMfRQoy87g7DfbLcNqsh9vn5OxqLWDbeXwTU0
pTuWb22m7ZUh1z4qhexbk1EHw55h6OSiiHThIQadsI5f1SY4JFVaZptMkvg4H3BS
z0tX1KqgJExUOUR9XfTF8hs01P9r3W7NQMDEemEaApvt5DfUe4RRZmRdREjrt2dL
TAVeD1a4lkdv+8RM6+IM7lJOf/iJqgW0sHi5aAbrqAkCl03XYY1dUGAAgcE+OGuA
ssUClvoQCLHxp5Zi0dvKHQN9KDRzSHx8E9NQnSNzFKkpENwjZDPz0d5Jv6hKAfwJ
1irUQ3F25/A4oMjt+DYrLu84auWEGEchY3rjbX4nKsHJe7AO1wlPzQGWu3dkWhVk
ItDlcI3PndXR1isYtxBGz+t+fauyy6QxJLR5byxyZe4yZtpCCZ3gQHpr/Hq7PQ2e
2zSCi1J1kFiHZJrKIz1u7ydNhfKWf+yYUlByohNyxDCz9GgtB49MUp9vESQxF/1O
si3ga07WMAIut8dDUECZWxhuaH5KHg1PLp5IfTcNCErE8foJMxJZnuUyXdmjGYrP
SktW06/kS67X/oEKs/mfYibkuAwsoMcQYfPd6XC87YOlUeACWKXjmyaklpuSdAhd
2ScqA3UTF+anTqQjhTznopTOQYklls4S3EGAw/ILEGcZT4lRAvsFytATZuR3SiNT
5XG62silOmuLtNOhcgQQp2WkoChjeW/6hO3SvILcEpgvQUwFA2P/14E0P1m7O5Yl
LtO3DIByvBEITYJI2etv21tWVtXQx9dvECKlA5ka1eOHG4ZRTfp6djo7t/VmHRuD
BgIcscG+0NgCDmLGBUc0sOoZCRE3jBglO+EH9c7vOwSxRMK4ZYC1tO3HXe7GSAMP
RVZHb7sQtELvEM9xwXB/MVRjYC4MEp46wKH4y+7njKBbTyG2RkEyKZelu7Qa8e4v
vPWsxgzUbT2BxulwyiYvtwGLmeg0E6E0bpovgtJDkAkuN/FGr/1N2UbRh+xHZDNU
7e9PUTMFow8f4/C2WDqfkN7whw9M79iiVfIxzWCkQ1L5YA7+v/WG6Udgc3j8/U8i
6EEKFuL78f/4FU1E9CUL8roSLQ7aAKEWw93zMWWO366cWLtIJaCXAmbgijiGJll6
9SXtqhxUzL7/KsVpyEAwzbiKwZECYgPr7e8uZxRxMk4DbZwij4PJXmp+r/QODGB3
IO4cqIEgImkAk4aWBq6pabxZ59nVqgvmtR5qJTFutyQJjbLi/9hHWeFwhjjS3Aln
O3fTggO23Njyy1NQGVZ2PBsWAMt8Th4YBgOU3l78ZLJEy5vSYHo8kcKCaMtkebjE
31gxLFbs+nXOqM0uy778QsIjPhRTFMV2njPA4ernyv757JDQtly5+uOdhYZYWmHH
RNADToFM2OOqKbezbiXagYRW5TYTdkXoMKeOhKnCo3P5X48BlvxRkwee1gaF9cfg
BtaeYbugyv/jiu/5tM3pnJtxUWh3+S5xxsN/t9zaBozRsTMF5OGLD0KCdrrz3xe7
DF68cFPOnz6MmszEhV2ei2kZzYziOFdjUukrVyOQNnTRkXk1LHxAfc4SqVqglLSM
g/MqK7/0stF9+i+IQAy+PudHxyy8OW+J3HMMLshJ8hxBwDTwgs7Ok57EW173Brxs
v++COWyWqhOUgrDU0wwytqwUPx+vLmKA9EL8Bp2KalwzkXqbPuG97PSi+3nYUgxG
VgZEjrIHn21JsZF0bLUDEnzELL6h/zkRWMZlBTiE0A72vcbFKcDMy0UoJqmuafLt
jis+ZTkTNj7yl5HiD7h2e9S5RjqVsn7PIp2iTRlkD7DioecL2YEWUm+7tGyh01Dj
9EDV0F08dNWgzru1UPSSRQww16RhsfLyOg8THZI6vra6qdjogglF70aHpq8XbakZ
7QoLleLqjdh48ItDjurVu0wbTRLOZ8QbqF0SMQLJKGoQN+0XyLmT7WCHqQ56WRtR
IWbsAA/Nq4I4X7DMgwdXiOxTB4Eq491nL8CqQ7Hcz9j63wFTa7zlQBGyMFInSCyH
Qp2nG7jbvKLICFwhPBsPSXa6O2SxkcFnmBl5zdpAamX4jWu5Q+lE26pm7deFs2p6
jqGBjTkxGi+AagjtAIHmUx5n8BmkcUpS0m1vKr/R+KEgk3gCwGfvMUri9de2OZSx
hevBoq9IDlqF0grBHI9zEwW6r7bU38+Kygbdw66xkXEJUZUZOsbcdAbo/H57Zwxm
GGr55xncF52KudA8gqEQHqFWXmI3rBjX1zan+VqWUmTCjXJ7s0lOKvp/toS+QzE7
ukQdgPDlj3+jWK647X3FsNehtBnGB4EB1gdOakq+acd2g+doWNN7ual2Fh+3hse1
L36zpP/lWgw7hJNLQ8VYw7KSFfbZ7foaHg2o6jN+WiSm2wMdQUGChIwqTknw4BTs
edEtYEhneuQ9EyPwGQ1j7WfHc7J9oioaSOQzJnhD5/E02S1x0EUarMcR/NVA6cx7
gonLU2e0K9ZrYXTfv53o4WWm0v5S6fdY0Ee7alMTcnr9Rn5v+aCfB6SuXYiAaNTt
Gzvw+xyQ98f3JlladKLRwP1TWL1cbdT/xw5KOJnNfQqMSgYKwcJJwPEGZZFovewD
ZcMnLX5YvuFwWTPsDH9mI+zUtdxhcq187jHThg/DVk0xOSQt6IrgkwvSP+Q2QvdB
1SbuP0XjLn5YvMdRWxUK2ztnDY6URKEn1dWGyRaycYWx3v7wfXuoQ9CPb3s/wYlf
v1yVBuhcXmWTGAk73XLAoXmc/+zkBCDDeN0FWcmX07LU2ZSAK6w0PetsRY1+tssM
+oBdpBK4qeQvff2bFrR8yjIDvGkzud6Dudfv/aeLLOgmP26xP+cG85E2wtg9ohGz
c7KuSK/U+w8bjisRfpE5H4sIHS8YA5nEth6R2M0RZ0qcdxwiSB2lBsGV1lTDvdL2
yOu4dKlka5qaQYUb4BRdISHviiooadeLid6VKtlHImffSlZhY4NNuCm3jhT0idWE
MJZHqGY/3P0xVBSBRiBeYbIoVjr+mb+1f8g5lMkUFkbxCEJbhpvxo3ThhO3W7quB
KdyrmBYAfdO0t2Zg81D54DC3Mb3RD9yNxRMD6qjAZPdtTx0ED2/H+S3mw+2xjt2Y
11Sm+RYF0StlL3j9x29SaP8YE5DcknFZi4Ns3V+z++i1vkesYFlTi0FK29zep0UE
jTJ8OJjO4P0bKcuadjgrEGyZRV84SZXVhbTuYxCvZG3r2j4SaieJccZiEropKmjE
9I/Ij70tut+DtFUZ+OcY7RCjeWWrTkDAjRVQ5cKwrVepBWOjAF/xoAAZ6ONiAQpx
Hyy01IdnKQr9BtZt7qxmPUxYR/lAauneVoc6zkp2QxwnqZUnK7v9dmRBTn4uLaZT
T02aUSr020s/a/solRboi4zE978jtxPWbLqUJUwMmdC8WjbiBjkyAFmH+YhUTVt3
sHJAK3EVRWgclCLtPOSoBHSNJz2YhdJu4OMuQXLzjXP6Mh5JBeQBM8+Q0CMJFcWF
G9sUrx0muxl1XVNAK4WfaJeafcbab29/fXiuq3l21U88rKzbcmmr+T14iUxkyacP
20RQ9FLaJqr1OsJN0GzhJwGZN4mIBlYyhL94l9MULBULTUe6/0u95B5lE+lZnj7s
22/J5m33oRwizfmbM9jKlYA9Gnh7/Y31um8DmqiUDtCSJyJILJz9egILwspoTOQv
H0EPYGEOA6fch7a4ziYAHKPcCNFqqGhiwoblxlVwNUlMyQGbYfXDVQkQWTrs3awW
z2y9xXwgKu6GrIMQ+TVnjVubKLDaS8/Ln/RPdm4uTIG1KCxaup1Y37c1XkYfz44X
SKZM3UWKCwZa7i/TS0cqFhiqUddnwkqY8hiG6xOWjwha6NyUSxd4mOVlGi3H2K6X
j2wJk2dQhjzwcvrbHD2Ekl/eJ960HWgRfHdAy2KrUWx0MCTuyfn8XgZHocXymncv
cIkP7+d05xkfeM0NCXbFtLfDsAAnf23d7lvZ/8hHBVS6dCE62TKHQ2OqJ7tuD4FG
cMyjyc5hbzLc9R/5mHqNRTFq6cIDsjBebSsYEOwPJ//ktKhkboNGwFJoNGomzSA/
PkhNy0hPb6Xinc+Kq36S1phiOd2rAxsFL3g9IYCsX63KuSlKJwpzF4ehoHtoCaRR
oabosTbE+18KDdqGZzrR7PtEo36GQ8YVwar8Rtl6ZHhRIaGHTvRqp1QSSwwa4lm1
s6WRinCuco/DsBcQcXIBCSVDC4Qo7iGGI3GC3IOj7itAhz5N8sS1cR2hvAmhV2bN
nOnvBi5BSZSo/RxEzpuf3iAIt+/FUFp7+r8Igh5r2E8EbY2N4dT20VCi5vKOx1ZM
+RpoLfXQrduSTv8v08LK9UCYusfNsmpOHm1s4CZh+s5K+XyqSsf9/8BCko1gVmUF
RFMllByRam/ejWJMHjqsA/BKWll+FPKuvVEDHauU9DP5Jdp5ZxaRZdVvLprj6tTY
/V6xeeOXNtKGLrip1IQHlGLl9fK8PsPLLbWvXg+yzDCUO5VC8zat4XcMJJMtvD3l
tE2pN9hJO2DgyVnM7WEqnBDDLfY4vXOWdp/65awVGgBUzqp2seTPvRCwec7MSctf
IAR7QgSjeqiJdqRRm9xutkB3pRTqNTRSmrATI/gJpfcCDlid//SmjqVCh5FIs3rB
MSqzJ8kGOSsmH1pwgEaOhDh1o6+PmXddyJrTjVVymY9KeOIm8ORBiIc4XwxVabuv
/sjaDUY2hVxqOwv6gkmJbOXkRSXrngCdQRq6YnM9Geqaz5yoCPgiTP6A5wEuDSoZ
0NBJeXp6NtSXG03ysclxzcZKKU2auKBY2mM0jg9rsg+U3Mhrg0D8YeA9D5N9pdEM
C00aht8XJVM7QuZf8qHiWekDW1ZQR9Qf7Vx2le9AMn3TuSBt8RjmSMFn3eJQmXlF
d3KZw1HK4GbSdXyevCa8s5Nb97pjeMsecImIBOrHVIPWmVKDu7dfRSd+fbstp5RT
C4krNpNHB3O7vMAvktHwSruQrqFiXXwbrohCpi15YA5LqoIFFLEYLrl4e2RNnsLc
lMx9hqumptRuyK6Rb8ygbh9gDlrnq9l64rPBUoaD+nUD1gUVGRpJm8L2cfv88Hel
HZgIStIY/240sa1lJdB3AmAvS0b5NHXADxPnqvHe1Wo5X6SyFenGfdu0ccOfK+HP
ZSnNxlGkkJyNaNn9deGMBO9O/hs9c/Fi233djHG7/OuALABVPkUfkv0KajjY0ZDd
Np4ydY3qZsaQe51h7tf5Zqqw8Z4sfC+9Tyr97zSVOzj4FQpDCZo/Md7UFXCUzQDz
SwZZAWj3rzpQ2LzFMxLvRnnw6/QwMg4ygxgdbcVyC6Ui7xo9jEyAKosZJ09Gu1bq
dc/MLXlpCsoEt+gf1i90egDKj6EygrgBUDPKq9NtL+o2tnD3IXIxTYVUkAh8QrsN
xxph/1KR+U4oNFg1o9eIN7dnEcCm3XuiCsLtqVmR0dadnbh1s6fksHk16UKvYE+o
o1v1OidoHHUIRgW0+XnTwyi0NrEtsTM+1Z+yqBVN/i8yhba8Wavi+/G/t6IuAIXP
Eiz/t6JkRJr3cG99pBEQ4CnmFotTbtsaPeIBfhQgoOW6HfIyulNIJSVQNXo1z0Mz
JGPAFE8auyQOqlG2dlwu/teu4kzr8YNjNlsVUUQNGBR3xzkdlrN+RFHJWufLB3qk
qpTz3derU1QLn0P1x57r6hZjSjkgRGqAIJSLAmC5IW6I7L+V9eE/urVOnKcaPLYk
DF6QB5nQZzewWsjmy0uxFqxohrUEFOM/l7SC77Y4+dXq91vHSlyRc2mFKGf+fJkO
QjUlbjRgbDmgJrTGb5Dv8EehIjEkdKnGw4e4lx/nTV6K6gSk7HWcVbb6wqIB18GL
RW7Oe9q8RWf9TzsYa6F4sZ8e986OfF0nkkjtWDEKr/WSCiQrQmkMe4tKo1lp++QU
awvz9N1UzyfqseGSA6BZtTzUNz08kIDxdEBC0XVwBnuf+dz7CHMSwa8VkzqTwnap
ain3e2HqWlWFhTS0SzqpogGTBpbK1XN3mYLgkQOdxJSVj6LPT0uYf4F3XcDDJKES
SHwqyBys4ZjcPNN+FW4D9G9FL0bRD45R3hSWcdJuZ1fHk008+FBaOq2ucq98ECeS
yopI2uauTI3VWgYXnAaWws9pzaEHSE8Fm6YScwwbVh9+fpbIT4vAfa24tZJGG7Eg
UnqkkvaL6FVErxWjD3XobYyATt9KcQm5qzSFKRKIwycXYpvHN4Zi31hUeDePpBy6
l+YnKxcmeY7xm+8hoV89alW+b+B2n+fDUck+tGHRtfT2lmO4jaYAttgC1n1VDQSC
OF5FQH7CIueTYWDP92o4RD09gbutCMvj5cXoe+cc0TaYRweVzgUghHS+vuHg0LUC
tiPZLCmbpuPKb+bxbJyp1XQO9Cdp4WPpTk4jdZfuiZshYADZb4bhsh8gSAjeh4mS
v3WahCdLQutBXwfjTULnD6HpPtB7AFigdQVGUgp+NJk30XnyFqzl7U2FRFfWPlb5
iOjAeCBMNBAMTNzZvzvX82Deq1UwmekAk2bB8hiD7NRmDN2SpMjbZzBuCwTzjorL
GCu6w0fmuBC4/EsKvADd97qoWtlyoym1w8Zre7lzmUR+aHfTPcRfJXHrBkQNwp9n
Rse/OaJSUrYLzVhWh8b86Q2XY3QSUVFRUQu+hwVlFox9nYOMAfV5HqbLhenyenP1
dJAHwBTXXoGE/CMdUy3RTQfU3kES33Sq9bNQOLjkZRVTJzQJATdhdAsSYcnN2wDa
XuWbYydCetHB3IhIa0pT9aIMOT13/W0DI9NCANhHGBa7UB0VsQTF1gOWKwOV9GVs
lF1v7O+vZcdehjniHx6LT4ImFNH/19cmx9lWhRiIMDyGE1Yyq1Zrih0Y07E2dpCR
RQ4mxNzhKdXXmGmNlU2/wI8vWJHKUc6EI1T/Xcfl+UmOntJfcE5lHJCG2uqFjIly
tZWKTOgRSVW9p3/kSzsimhhqBB68I7BU5tdzKBe3TcVm6zLv4yCZpyhjs5eEmiBr
D/1iB3CkG3o38BqXGgK/trOR2uXXMgVHYonX2QT69yIe4AEAxeZ9SdYUMM9Jf0eM
tLRyAdfsovoheHIYapyKQ8JTeTOLA8eqSngMy2VaULq5wx/ZPJOozxwDTjrQkGyf
PW46f8aiUqK+bHlk89kC4R8yUl0N7nK4cR9x3NVdsNLsEnPt8aigVKXXAYTw8Foh
OpXZrxHEfcmcreLwjW/pTiBZqJf7tvra+e83SZv1T3ffoincj8OWI7sAiTTbLkYY
SuvYM+ZF2pArao9GsBBiZ+/CaQrlyXqUF1/Lhxrg0wtiU6mv60aJWMVPulF0+AxA
4KG20H4IrvXGKYYRzJlRB5/6CkFxAnaXiN8jjusYXmv5qt5J78OMFITCPPdWG5sg
mL/+nCvXT6RvWlOIOck4kmqfR5ZmS+/nMeW7OSMPWXd2KP/o0DdyPlMDOaN9kJO+
ORY+OTMqwH2uo5/PY3gzhVKr9WAL3YCyc9pcpPwEFXAGmiPaBVEI65IjGHn614PD
gWlBVrnlaxK2lMw+s0Fi00Qgh8CzteKd4LjtmODQMZ0hYoe4xtzdK/vObvvgNx5x
TYOBFr5YhKspUrTBky8ZFFGNdU6GQR2tRci3Sz1o4PThxu9r9aQcPlMUxnT8Oke1
0FYLga2UD9Z5uACKIlnNGoojyjgw2GFF6gqlav70nF9tp6/eojssg2Zd275VCC1U
+6V8DfZwJnCuV3gORPsTVZQv4qoHJdF1KSU+hayS8edZP8ZcllBYIpoZI5AsfQ6A
riICWzXYFijL6QLJmDTRb2sdf9gh+duIcFZgHAUHfE6kOJAIgYgT1qYKrCmVcfzL
M39UHTqCJmqMOTk6fXNsqjpRJccgVfK/wLUh+leVpKHP/ZceHDe7Shn5Wuf/GzZH
u1NNjqt2RNs7BLmV88UA7WPPvXHpFBDebz02nmJrOC5t3/q4Caca/u3egdD5sOoa
ktMH9QJWnr8stOWB6TMfKAHnpRQBTe/fuY3oCb+wJH/ZZNUJNstoJAXOdgYb+udJ
Oy9UzRNvnE3+wg1UEBDXb1YmJSALZCoaBWNvR/bzn4Gh24CHUBT2iNHNxSbPTfN8
MKJ9qYOSVWg7ZmbGGzbz79wjMdpKhptDASXdabgqAn6uJLaygmdYzKW+7XnW5M69
uCHyCC6lMDjPyv6Z+s5RiH6skvvt0A6pPHHpM54iBflbPBj2HVQX0xEaS52C4MDp
VJbHfnt4EX6mJpi6qf9CUcMaDbT5JQrjhiLEKyxqwpY2jpKjh+X4cQLrbyoBEo5T
AWzotXc8fMGX7pn9TZaj+6Jvd32sDzMi1cpL5dp/T2ssr/O8aUggOEFJcWSsT8qx
9zYh2r6FGTNWS8jwt+LDOos6M2oke2Padb7+1DXhwyKNFFEj7pUkn/XFbB+Us2S1
c+TPOBZ0m6BglmbDBZOGNO2NDyP+WoDchZ+LFPkggMj3rpN6EZgYKJ5JcyIxJEHE
vVpJwX33zlbiCRBwTdq9FaKIfGYG2AlWi9KhoUvehCRObYWwDc5kSI0kQav2dbd8
TJj6rekvdvQhtvg1Q4wsSBt3/5t8eZTvaIdGo2wyvO7yT/CT9qIp4j7uusomNVDD
p70gowv8OJNR6qQeVxLEJXHriuAfA0PmsfJskDtd1xk5FL8Tvsz15fMEyu5Zs3T3
MC8nD6/83DS2WDKZRgbdG5YANuc2YwLfDLeLF1JPK73FaZWYXOvw8G4nE+NOK8xq
hRCN0yUYi90xQWc2tqxr06FcAqyU7oaRfusEg8jShyJ6LdZYhv1+uTO4vpaov8k/
uGgswRJkq2YIIZ0AxTAFuh8IDNsesUGWv5o1K0K4eolpDuWrGIW0yuJ1Mu5/+2tC
gulFc19fHNsypIdrGBYwfILYqPWwjziG6+5qa3gyw3hFpZdn6A9tj1JwldFmDubW
Zden5S3uEMoKkPRby9HfU9InuwRweXOiu3vMIWWzarCZ5idDyMHZOByptoRzlBmh
8xDloqUwLIgosG7C8YESdqjLvGLpJ7DmXN+Cuh0SA98pblA4K0QaI+vFMHDzIvdu
M+B8JNqw7crSOsiZQ5wedZkkCqZLqJG/GWPguUgAgLrfGLIDYk9yi24OdjjP79Wt
oBYclohzWiwVeCDiyxjCXceFXTJexOTt6DJJvocsuKCn8sfoo9AvlTuQ2bdGsyDj
HAwPBg14+OuGciRGcC6wtUx+Z+sawhs6Shf2dePCf1xHM/S5acNpQRJJKlwoTNyY
anb7SZF/wo6C3m1juEN2wjiO32db0HGWgV/9aLfTO/42ZMaIkH1V0+F99DAyOeIL
44NvhqoQyUOzCrz8M/3+EmruSCPZJdCXJVTcBxYJcFuaAmYAbwy1cvmsURFH6rl4
Shj787HaoIxg20Cn/fnKJtVCMu5sWVc0BsMt1nWcqkajyNZ4I+JF6PwLCEeL4Fb8
dPo1kb8Y83GiuVXJd25fLTGFDMdyIsEBO21/fY2ejH7ZulbBI+K9QFOIYdjfKLEr
PpSE4q78NdVFGK1RvPlIcDQqfeuL3ERZPtsFtQacDsnyxPwsgXLFgOpmg2cWO5yC
JDvMtH5lt2yqbSXj29Sdvq+0Vv1N5rBOknOkqIPT60PpCEnQMKG5+uw58GrpdNUf
BhmbO6S3bPXIDCUX9mFN/yZIMKtouGcDj5riHHA+kLUIhWYs0I79N3hG6LLDTbNG
w+18y1NO41hmLIzGV0iBPItmK+I39yq5Lk08jtZ+NMQv9Qp4q/GhSrYUldb5PIiU
CtsbZ41fITj0Jx3USCW8s9YYxd1Z6LUpJUG5cAMcC4osI6/gyqk+35Xn3cCtuT1s
ryONNfOAMu8o0c49VwvNL5BfhN1QCsONZCv+RV5Whssgn0hDRetVT8bfSFABy9Bq
+HIQ+g0bV+rZss4iXN6bee5tylb2a9IeDvqOLHKX8qOIqpB3G0AN2s72lVCR77NN
13L6lwoSXvnvpI9UTCWn6fSEW02PQb2ABbtokx2DEfRXuJFOBa/hGnhQ7qgm343h
LX/LNKTA3RJGGvCAQ3rjVa3PcLo8offcfk+/nIvhkooJfW3CX7K6tBiaXK9g29Ft
KwdGXUaec+RvvrWegvMM9r5htBy6WYOuxmDc0yZoXpBar7teDiuSFoCrjKg6TPXS
Hj/jKZ+onUYtlVHjuZd56YpXndR7CTTQcmzOrX/tq6DPVH4V2fdJ23nLQIUC+s+J
J/NjTvQW4kMuDF3onaAjkRqfqUPLwownIt2M83cx9yU8SC1rrJpZ0z1eJeQ2SvtN
vBJ8ui2SU1vvUjWqlNpZuKtA0uuWwyR2pcC84D+3Q4cza5GunKO211o/Qhp/7ZdE
Ge61tOAHZMEfzGgs2IUSQCzS1igkxQLnVpoRih1ZH6LPUlne7WEG6N1kfykl3vue
ygt4YMMVwwyCR41X1LSczs7oQHcNkhL/tq53oKm1SBlKev25SQNxdpCDmabVeQB3
+uqOdufid5eyUR080omB8CojmYO2p3gZWY+N0ipNa932aRZGLa1Zlk7LxCCncvzg
3BlUdOLkFamcXzFFhp9qYoPGU4cBMBwWxqYMRLBnRWFpyjncHJIxrhY0R+f77sIe
yKfQ1DJBEVmz28gYJS+7mSCvg1nNlueB+cM1L+QfF4PSwKP32CxI4Agok9SBPQGe
5CnnXgui/HpjYdj/iRpWsGgpm6NMUY6oLd1Kcp9ZgEI0VqqXtL5PBxdKPf8nLy72
IsBxP6CJ3MqoHFDE3gsIQqcKdmEAQHsiCdIiUnUU+QAn8VnDyY1UFOL8/A48xT5t
j0OaFSj9oEkmLEkz1jV0ewXMxmOU0CpjJ3m0MnrlMjeMUG1QwMCBUk71/wWkyd8S
qei9Vrckv0hmlL0Lt/ErJUs6MtQHr8q3/ts/UOrBqO111PWhJGJE9g+ftVaEQXmG
gEoD6CFW8rSSdRxwRev3CQj+nBS/lUTjD6P3jucrODXTQ3gyEV9mIDm828JZAx+R
eLYeBifRGuxLv0h5OJYCoObM3JLAE+R7iyEBMYzgdSzBDOSX+Kn9fAPtd9uo9PCE
gXXgjdQsJgSK5N2q6tvJWG8JKVVZQ6/IzUGuRnrjJtoDWt2CqSZFzGbzcc8iJlEK
ApEPOM16rpqFPckb33B5gtxzcU13IPqEizk7ucydQ3x7H+QO1+ULdRs+lAo3nuy0
AFgbHQcz6CtB41jfW41j7JRxJ32G7xF5crM1eGkckZxm3x9gemONmRqsgIhAKw1F
EmB7FEvwbnqo4I4+Z4A2WQpuKZhKfpTceJra0h7KWd8+/j/sb0TL0S+vorhlH+4/
QzGBVuqwWXNmmse+Po9eXi3IpgU9AG4XpE+GU25ZKw8j6Q97hvgaKas224tXcrpI
AGiZbq1DAYxflDO1wl7D1oIQKf9nLB5Kn4TxPyi1ahgVDMTeO5A/NfQ+mkCSs2DE
GQWvWzYZiWOKsb/GD/A9v53BO9TxHA2WLVgJwQKIMaCf9y6xdnNPUxsFMkHwymJH
z7V3x39ksWxlBH9THnyvzV5AenzouHHc7rJ8ThGIzo2LYISBf0jcBaL1B/HIJhpu
QoYL8G2hJErISu7PS26cLCGcCJExjAwOIdIImlxWygolsEBtssiEJBXnsCFfoido
nUEqCIg7CX2a/LO/pS6fKSMPE+jDYi5GbNgG3MYDe6foIPny4BM2HRQIUMtPzE32
w2mGHVrqtQ9p/FZOK60PNQFCgcCjO30zcuPtdZs7J1+3lPQh/8LDx63NKAEXcO3n
lBCmPO415GAfc7Lqu2mRKoKs7ZpuHZgsElXWFzbUaHjN8QjivPML9qxeP7+J5nsX
mEdXnP+Pv8zeHh6kROd6BibsjWhtke5xZjqsQ2QO7ESa4lkT4A21EJhKUFfXYD4d
R55+SUymsV7i862qL9a4oLBpJquMEqfcUxPzy/F/I2OTEJYmPHWqDIDpxTLnp1bh
biGhIjWUw+JUVrMRvqeTYAusSySUT7dg/Z/ddOj+tUwXQZ2HlNzUhUgm53fX85At
w/hw6LEAA2b9vD28YF8fm6fcVADx7jOcovkRUY+P9qynQMvMTjftnQ2LE4E1PZjU
9YUkQzO1T41udpkkIMLErJQDq66OQIxC2tM3ZVQmK99+uXLGvFtACgyDb9HQ7EgI
nlYyGpUmOYsJ5/EXpyZRnt041gl11EHxDwCBo8spz02LFnRCYGQ4/1Ac9Ql3Yt8f
Hi6nyrpvwTUDGji9DzGMoQoyZAwPbbKa6me6RhQdS+/RrwukF48RVBKT3VT+80P9
TBrUfNHVNEU1rrTdSERJEmJ/ELxhHPMN3VpbPCiyWB7DSL48ysfmuXLHd6LH+3af
rck6x36rg+MWytmyT9kV8hcCe/3ZbgwYiNzcxGqItR6k9d1qLaLlCzc5PA3ITNRH
YBydVxkvHTx2vC9t5E4HZMIgNaaGBmBD4hB0CQeLmGB6hw3ns9ZtE46ArjlWpDLH
0fFU5mN+d/PIx4QmgQTg6bNQjEPr2IfRgYduSHjdaDCHlE46yXKw2pi9P0Qj8ROP
c7oZdIq/RGkeJmTh5ilBS2iFQxoCiuxcBuFp517SluHELTtjKmFx7/tLS7QZV815
8V+y4+zJmwlYz1hFOzso9D/gpCLPoIJGiS1SNAQni0Y+mkoIo2fbMzPpNuCJQu6P
CmeaHRfo2jBu6bVQNiGP2N+FMkSIyAMIMvDDXxlipuF/r1CaFBrcFwu2MDZVdHA3
MPoC1jrOVFzQ6dglaDvYfppooUK9IaP8bPiUV525REhz51QOwWxPFfyIH89QdflC
EdJTFzWT9RAVOZLQZINXx8csB/mvfOuQzvB8O+6oEq+4tPDL2tjbS6ouQ0p6uHIs
K3wd8PgWjwChl1fkJKVtwH/OVZdfG5g14xjGjOxjf1BRskKXG9SWl7REgQ25fVI3
pWv31Ia3qjfMAvYMSPwRpVzZQq1afv3+YoH3Zqw4IvfOP3vhO9xWwxB2z94+QiF5
px11t5lDS9aqTimRkzBsKyYTqQH/5ENw2GhhCH+uftrxmcM6SEaSQdL12PF8jvx3
1rALPPyqJoLiLnhkbx320Y3BnpVm1P+jEnGi9bW2j8jR6hbrQw2VcCYdYjCuZ9CM
6Bjni++14EPGKW3Bk4xzj2XzW2gsE1LnZyzytEHeUfIGr3YCR+UK3WsNzRe/+x47
4vhi8NqxEEKvaJadV0pnMJzZc0mDfIS8XAQS6D1/sBbbi3Msb2ABq+LpjxO2tNFu
MbSN32Sa53WZf5tKuCAusjg1Pm2YAIXfBtwdp7rKX8rf6ns2tWCxzRc64UWYHBAD
ofuR/sL54NTzRwBeM5Wd1OVs+6+um72dyE3DVYgba2XAgWbHMr2Z+1Iz0Zjltp0m
3lqPTU+Q4PTgswC7L11f6Roldm1hFPDlOWKWLgEAW4/aAvjOJmHYDEvQGf1RiLTg
9rP+5NWzD+8cmMlhw7lCqCxEE2lCYZ9vBQY5qKkG+N8a/uasO+5l42jVE/GZSVVf
3sncntV+7obTIVVz9aT8IFgler5aW8lGynymF+sQIiEl4cguRWVwSA24JmRvrMUl
4wmK4RpuBzvn4rXZa/oeUcBAoZNbxHfGFCKCqv0CTaWwYSRJ4M5MWcKv9Ba2PgZ9
RqFgkT8MsSP6GmtkGYekdG4a7iUlyoDsnxah9x+Nld5J26FsVGZmbGk42MZwGHxL
G6MinpKYL/Fv/6miloaXn0HqqjzUlyzbHz5aZjmfYjyT2xSF8XgW4klJ7VyTsxzG
9r+4OzU9nIpnVD81MLrL8K7s/BgUMLHSS1LXvMeTNsEpTeqz+Zdk/ecwyFHeSffP
uZ7uWAGE3w2ftSnJk4rn/fjqzLPUGdfJ81YGovPqMCD5LbM93Fjp1NBmLZ6NrpGt
+jpIpEi++SDHOn11oixp+SnpxZtuv0MbWqzIQ0moOTS4ACMqVcHuDtzh8KFPhEfm
n3e07gjw4BsO+p4dJjh++fGkqtXedcS85ncwD9dc3EVFPQD01EbsckcfDf2weR69
BVFsUNaOhT2z8P/CC0xUl1NJTe9Cjklru6qbsYMfwKhZIl3iCkdqerFMDfFFJ0kt
hjg0Ge1Ut25VftBrR0kMDznehjRuNTTmS0vb9zNZfySVJjlPANLc3FBLZLhOa7fd
X3H2fPYVMaO6tOTNBS0Q6w6fu1wPuz3d+7deysjGaqFd9Wm5XC0sQmld16fPGeyu
py8YHFs+DFVxrRoAc2XPfpqZc+VgMVGO6JyHOe+G9bccak8qk79ytd4zqeSf3ny8
yf61x9SXbMSNEE6xkvdzHk587cnrv9yjmVIcN5qaeBQ3zUJrz8+rRhBcRJnIAZqu
fHS+oUFwBBuBewDID2p5KVMwyeVIVml0bV3rCmD4XC1WoEIIti+h9jQd6WuUYH/V
zenwZmenP+qsb5+hUUoqpejlR7zbKK2NV0HKq7vreD1ZbRhVxbLUfXWrc6bg+R6l
dAaKq7JnzUTMjyCt1yKB01aMmrtENfqyrWtjKLUszjZpq0i7RX7ugG7s4IwmsE9N
kyvBl1AA+rTguZIdU2lKEdDCn+ul/uHu8I91h96K/DRvF4jXyO8rZrFxcvxkUKoc
/wWM5uZS1BoQ2uOzKA0GZW692wacnHZdlELtGvVPUSbAUm6srus7cbUOQIrEoO+j
VcAUhqbP8sE5MIDZ5N0wYDl4eBsvghXB4LY66UO2k26xyYgmLM2HhJUrOrhP0Ws3
uYmUTYOqBOhk8A+3/OMfucte+bnijIO6q/qnDBBqYERN9um1haHe20BTwxX9z9KC
LOHHyGBTVHSjXz+dqRO5DoeZ9yc9nAiSlx/zZrA3DGtvykDwJiN4Wdr8FMGDJfwZ
vNxYTIZmhOWVqAsCK5eLuFvVAF7UQR//LAsmfgPZCyea5ONrq2UUPrQhi6gfgJX1
ViFwV2Zicw9B/PWprfOc0uKNMYtmjmN4OKGGeqltpy1tuXs4LPYbJuH+57TTF1k/
nPAQldwgwzSd4qhwZ150l6SqJjZ0WOUCEKcQHXQknJu+l+eWAnAge0zr9gy/tM1r
ccwT+HPZKGntvj0+S/tu6PwQluw7ITw7O0YHlyWS/EFBNU634Au51Qg9nTEXPlIS
kqFc8KY+BInP+bhAPNO3W9UwI8biPMhUdwnxVnwxwL2iZWdkXp43JpiSBTHmUAXy
ADx+YdnDSxS//jdk/hdglVksiNoUSF0XwQHUPN+gl+2cqu8BtQeeoOoZlbuyCdtq
3xq868baUshKXZFWR4C+FHgmHgpEgH3fZYly1+JSGBNsXzwIlXnE9K+IhlOzKhjk
qBBdYIEyUH+tigQBny4MQW/lauoM78Jecy5rMmtzLAZBTu9BOWJ/oVAKI6UunapE
xhHT+zTf8zXyF750x0SYZrx5sGwRUJCJqGIHQ/7zr9xgW5qYpmFMiCq1CkCLOxXs
ig24a9sgrwUV96FO5tAujNTVvYzrOT0AGaztPvdmfwCk88OvNgxS8W7G2kCTDoAq
sshCZxyGyx9Ngt77dAbVus8jpHeczTV0bMNKG19fGaYzS9aJG7mzB0TRCgkD7e7a
d9QG32PW/PQs/xqtlf49kiRddyGpYSLimmAtpW5BWqoKu9YLzChlWWjWiFuQaFB3
FX4gjC1IxUnE1hxlo7r6OndwmL5mkQPMItqMgC+SWUmmwmoaGzgYN2xvwqYATLH9
1NHojTZ7UyRGa3mSzaU/6IpTC/IOPa4/p6yMIXFBdWAnxFdLMdXtLFWv9ubkRyxN
ufD7E4YRH9aK25gAuAcQwguy5BSDb8Sm5wAYRhMoFKEeg8OdF00BnU86+L8qROIQ
2Y3TOknQNK6hh0DMi2Wj4MEa+lzxnY84O3JFtNBJQJAEls/pGUtZkmOEk2rpohyq
6hK2Tsqeej1+YBiDvThJtGtyToQNdBqxKtic+KhrEMA3JztvWTR+h7hhsXUd0Moi
TPQWyVzUH1m/gC+I0I6b7e/cqZ0/vSnDmw36t0Df2GweN9uCapUk6jy2ULNPyL2w
baYDZMTOkkTG5fAGJKYk7JrgcB3DEg/MK89UzxgUUuTmxf+FYoxdEnxK1UY5MJE8
gE6ZJ248eWM4rmk6+nq1I9vM1TJQNaFjEbn+Ci9Ckh/ie5C8m7rYnKHGsoQ5K9+g
ALRfA96aIwe19+n7unNk0sm80dJr8XMIrD9SCU30Coh5ZTZgC+YE0sgNncY8i0m8
MmBvfl4v5dAvc0PZpSTj/GrJqKlRxo+1WO5JVqbRN+5637LH9L9NXtTXS4dpXOt9
3lrLvgJNKydEQvzgC3gE4LGnTbkVOnEp7sbkhJSYj3cyLkJofyeep3Dln8Y/jek8
cMFHas9uoETboCqVJ/O5wiD9b2yx2L5mjZ3pVPU9vpCStUPHfl3ikN7idaCGU36j
4yAL8anETnA48QvQm3B02icbGnpwJj9bhINRXivOTpjxkG6Bj9gltII4ieHcV6fb
25C0j/N8MqUVw6q1FnPwOL6QI65W6YLJpfubXXErSr//hMWhDyUxKm/httxqPWVU
yuTuxeP7xnRvfAWT69vIhTb3ozI8A2nEYfhmTh4mRBMFLAjcjEBGYQM3HAobAbHS
Un4lI1sVjV5warJwi7/LpU9E4zAhGHtvhc/d6vUTs5uRmZjlm7fu5OVTb+RwTz2+
wmLd8ryBfK0lpM776GMhuXsDwtxrukCXBnJdUvDZda7WuTa15AFsyP7csbNbtFL8
r+Yr3YbBN8rJ5EzC4mN5kl67zP2CMPzjlpHapWv0hnis3blZSz+3/LE5Wdcyf2vN
yYErLkEMeS5yod0CaryQPVaecvkrXrK97J393NsuNBs7zIkNfPpi4DODoKgLhe9o
7WnlTIIZyQSLQteKL88TY67wiFp3tkYZimRaYP8AMNVTuaxhz/crCrECf0PP9yWH
3eeFjkx3gMC3CMOMa74qanZeShePLK5Fc27rVaadwzWarit5wQHsN8jpiXR4opYn
HYtuN2wXTn53nWrvJQf3vEp0Zx2uCNbaaFlyhcX77qg2Oyacfct2b5EDIAldB9Sv
D8/yYRjWK2MrNpI39PYktNBCbb3Vfs34m8MqhSXkYa0THOJE9XYZsk8QnVu8/TTb
D4e1vus74VYWbyAFV9SN8GpwkkoIubr4EorWyyp0g0UkZsrUQfxLKYTZgLIQ4OO7
/3D6b0awF2u5xxcq74Hw7OLNv5ITbbWdwUyfa83cFbgB30826l9uiN9CAtU/2C2k
Llmrjq36/vXDj+B5pke4p4Olbd9UiQIcCB3u9X/uerpP4F0pG+ci5mpXl46m34p4
CdzEuMbWP4jO0TUhtMrd2ll47QVmSa2WwUztgcOmR+BqyLAIhI5weB4G/IxtLca/
OdEKhyYPUxHIRChqAUWFWxTNUjbLHaQPFxYaC6T9eNYlRLA9Lq3KG/FEiYFZD6h3
48ZLsYm+QZuA8BVh+vNl/AdlPE/MqKNDLwbYpuw+jhmxyI/3V4wmUcIMvt3vIIUZ
cXqC47I6dYIYRTAoClixRcJ3m6KLMXg7NpWOsQrgNeiXYyqEL0Fz8+ZZBs6LpHUd
paaGsdTxEIOa4tOl5m4uvN+0/je+mus/sJghiWSLgFGbOw59AxHqqC4ONqk6srYW
EjC5yb5naU9f4VPmsxvFLfX++nyYeQxSXmfaKavVB/t0+BVD6KUathhWMU8CVR6e
jRFku+T9rwk/ZrFqmerLEmskOjElEcZW18XQNgzIQPGz0Y6gFiklykYEd/RT9AOu
8dPXtAtwMnCaxMBihrQkb1vnZu5BeEDnyX7dX524nKfYmhzq5ts6iOVJkterlQ6Q
lPWkuxrx3tzJjnRX96nvaOPXV6ym0AfFM4em9ZgJiglvwHc9tFfP2Q7Gs3udXsEp
dHiE7fuENZn1j2xNABLv4BZD3kNFHLYiSQTvihDGJcRH1o6YRSWmx9kcBGesweQa
22YbTWhOIoyc0MpCzjLYq1ik52UkZ6x13xwPLOmn8aEV8c/p1Zwda+uZ2skRX9q8
moD/tyyrkHGUOBACMd4yZg7N2CWS2Bx6x5MDuzNAeenENeweIxfaaEO8GwmR8NKJ
/dxt5F4lLbs2GnxozddFY6hl6cCCzAGB7isw3vDHKh6v9nCgILDsManOdcoH2Wlw
StySp9Tcj+d51iUdSYMtOm9Jr8q15B1TMeh5r3zAFsCQzrxrRJ6Nq31UAr2lz7xu
G2emnZBJppSKH+4sr4ZIDsifBr97qTye1sc/HBoKYYjOqhOu0uYcX4eSMxnaIkeT
nShJ3PY0Zoejk5rK8U7o1Nn6LJr1CMvWFCX7zkp4HBPw46tbYR0f7gg/DtvoPgOE
RxluSxAHvYlgYkSbb1Db2OWq0bELtWfdGVA3/m1MifZtoV3Bbl2r9ZhxaKI4lnts
nyz+BCHuuJMqREevhZnlNDSn5uKYKfgSQQo/AGT1T4rsE7YCxSpi74bRnFqyyk88
LvExAjVjrufhkYviqAN/61rNsnzzZzq2qamwxv+1ZAUyFUgqQFTKhl3a1oERFSe1
L8OQ+A2K1bvRlb8WHfIitNBk9glwLkx3k/0nHB1ayxkJ1Zq3FHRqp2qmbInLJNkM
jQIkpmjTaDFmIKrmGUpSzW1/ELGun3yIMAjSd7NyVYZ3OrG/wLLM9ZJq1LOMZttN
7aamdc5XFrFSo/kpC9qRDm4SemJsaTmZM9bJ8NhGil8hxQYBzVajs7jfMKqtB5xK
TIuCiKBLSQb2Nj3zJal8UenYxdxNSS79AsApAF1RjwMZuNdHSOhLSjsUv0WQjsAJ
yBTXOArzZTcy2EBBAUZAqXnW6ckApWLcYqwv6tthvLdsft4FN247U8M+1fVNmxKy
cOpdqHVtJQyF2ZkknNPJiYjrmTZPrnY1wuHqEvZac7hszxPpo/URrV+io6bcTr8Q
oAYaD0MSs6r8/c9ewOKmEE19wRtY5XJ9R9zHuYzWCSTRIL+kHOsgj+LxpDWK4Ttl
mLRh6NZSRnk13sy0CPQHanvw6khZcd8KB9BVFOVYTP/1zH86xyL2jX1tvJFa5BII
07gyJnE5Nsu3L4qKIOKSmDNfCeHKivll/9GGAC92HIGWW4Eu0FWKM/j8kPlTJgbG
ouRig5YdongunknTWsP2a6FnI2UX7hUN7gMo2FsfUe/0yN2cNt7+V6oCZCkAVD/p
0ABi9epzN/+fkvXDAsbpVE+W43AwAhReNs2L3CUr4epKSU2Pk5yEUyxxaSL9l98l
J/zkvP1OrsfzVu7UMzVPjkzWlWiKZldW800H/QDiS2GU/7HJ9oYVvKw58+M6PnWt
YqR4BpFlzwZ+YSPsRcfM2meAzu+4ArErZRn+x8LXeiisMgvXGfQ5jKwevYX0c7xY
xPfR+u9a4MkIAOUG5iQl8wCZo/zeyv2JMl5Fz7xnChfO8wJzXIlHpLzOSBJFzoXv
xkhmpkfz80fJ2o9+qr2L5mebbj4aWH4q3IN/6uo/Fh6JGcYdd4dJWzJdegzVYFPu
6D8jNufQEuoeyeHK7YvYUrO6gMeqgV2yiYcdKyalsp8C2WVYyp0wq6/MZ8PRGBaG
eM0f1ufdvKiu8Ua1v4BeQ1Nd8gkvNOmaQwueIpN8zRqxT9DsMpPAZLKsUHkhHwtL
pb6oaTp5k9ToJRAbjAXgB10v4A1g/E7oJmJ6S4IOT6AHxN/Vjg7sgQfGANRpLb+F
Bg5PuB80SCDMoTC3Zf4acNnEizhq9NITrMrRbwR1gXdHzQFcfYSX8PNtP6Gia7BS
YBqlxMPeBvBxOn9iVRHr0TC+xi4cCSLdJTRm+Awkh8mlBhG5F3H3vVVjrxsAToBW
gqpHVhXHvG5IftbPslhuowJUlfATBHR2u3HUNxwkjRUA3qB6A07tlZ3//DYtcWKa
2RuoxkQvPASAZGbAx0n+aXpVgDzJV2W7tScUZ/5QI77Dk9xNehfxBcRkU1TP2u/e
wttDsIO/iXyLjk7TVOrO/LpJHbR1zv63+NrOwEOJWOb272OGa4av2I94Le2e3iei
EHsIbHpPKakZys+Q/3s906yGG5MYyfUZ8URBT2um1Tx5EQ3+yzsD5vva4/UWE7AO
Ji94vSH6KRVlvsPGyLe74kKE+QguS1AYhAhsvac54rzSqDF4i32X20a0KYc7DTOg
riduF8kii0M9NpfSNzFR8QdQJ1oYfQK9qSkSL++CXrmA9NtPfsvQejTgAQtNrKP/
I5+onf+IvMckYBl6Osqcl3gkpPLu3oO1n3+b826btKigXni6BUQX8yrvXQMU72B5
PPEmqMbQ1Jfg9d6JzVBSzIu2kcD3d/pAX+FT52hUWSGI42sUTDFW5esImqPy3697
r0tZ1CKgVSQCRErTPe0hhW+yD4Kuld+5JxQr9zjkvpH40Axc5aXCBUXWcI0G24Ec
Lhc9MhwlcJG336OlVPekGTFNs+d3OKQLw3YLDduXZL44UqiZhqe00GGkruAu2FE0
UhTzrx/Fwl81ROdhdReArx4fPdMEQsGhMip3vPC7pcW5O3Wer7ZFO8luKvZpwYvf
mDZzz8u6ERFfkzNllbMbCN9a/lsZjCbZfndcEp6vg4Bl23waMK+svGQTxY0ESbgi
46VJqpKbhnAhPSE1Hbynk+ldoeGMnZM59nIzT5m88pp+bsTLIXFX4tSYInBYtXRo
EnDAZdSxXVIrEzMh3F3F38dILFCQ9AZhzUAjy6kx0EvR2kPFPNgz4uRXIxNfqXbi
hs2BGVdreK5kt9rb9GW6+Fi/8ZP3GfZdC0xQOJ8ln0GldGUfG2hsZ8bPML8g44bE
WmtapOTOPnoOmLWvOuK60cJRSMBBb/nLwFmMSB5tSNHNAotKw3J8i5iJQxkQHOUR
JAW2UR+EzBGGze1w1Awejxcg0HKGzTd57qalWJwYYB1qkE0Mz+Q5gM1D7iIsxWyq
NAMVhypu3JrqGabpkIr6xQjdhVPqbrVeovVRlz+MnOG66A2JckHuAlO4aLh2zS8T
aQnTl/KLUkRItIVN+2DzkGEk3ePEdc3BtsMZXKq4alE098lMifA51yrvhmspD2W0
ipItOVtFWCvfajBwLhl0JXaibxQvPcT8SCPgZ5RauqNyVIaFedxexdunEkVTWRMd
mHlWrd+w/fN63pUoWYUBz8ryBeecyCGxGdYg15A8rdLL9OFs/xj6+Z7+miiDS/uf
fY502Zzo2Mi45jDQH+t2ie3FG1j+gmICUnKThrXfuQrEj91cmEwdYcKSRVAJA6uM
ayxu00btufB59LoCA5B5GX40WmBdCEvMEdq4elh7hgkwhUaJynfAJ6+ulNLpx8/c
Jvb2I0qV9kDzPG2otqPSxJv8Ll57BZHlNdXlKt01HPrsIXMzlf0A1lnkMklVfDnc
tmdmC7I+Yf5nX5oHOLID6VDscuIZMDiK9Z2xLN62jKj5ZRsVrxtHq81JhFmJPoWD
PrKUP6btvSBvZCyUiebnzcjD9ZJqfdnQ3dj37RgWjHPH/1+WlLhR+acYSqEJr5S+
jjQPQPqrIBNRDQZ6NRGrKA5Y8mq6U4ODv4l1DrfRnbJ92O50xKPCcFmwydFJYf0T
Z8PfOUcBGStmglbVyCf9inyHqn9t3M59waUux13C3br2ne6NFaEqpmMegknr6h0b
i6cWBaP7snAzz1V+GBfHBDhGy2sf2v+F8IWDpbih0yDafD/ab6X8pCx6/ZZ5SnUs
jY67ghQb8RlY71t6nMHQjVXQXEZEOvfrRLc5ezoZm7d/eybN/CfVSLbwJTIEGZSz
L6JHDbIIzOG+tQ66YyHL+llNPeSFkwX1ZaYWKi9NaBVkz02iQpEoqaubckD9SjLj
L3jQXRBpIHfIHJNt6mQNCT2Kx/1hFQU4UKobuBnipCBgYkykfXrKt1fktKdU+2Ln
WoKGnjCfgWHjnW26c3yEZpeSdB585zlmQiywr0MCBx9S0YxuIBtRjQscIrf8gW4v
/ID3A42g6uz6cji5nMx1SQ7oMFSJTJoAHHIK5wZIcbbRPTqfb4RjDUPlDryc3RaG
DZxOMgfOrmuxVHhxA0tHmt3jC6/jF8kuljg/JqczOaTIk4NYHwgtdVDJytT31etx
81uTU5lDgJlTJJKYD0avrmPBiIh2xjseynUMg8iCg7FxK4osHXPiZH4PRbF2FAhr
nf6JIvC912zrg7xLUtBYCjmM5MG0jQ/qIV0zYBuXKQeX0PmhUExjVrCXfPp71R5j
oc30y6U0OGnoirAGBEYzOgSV2puC7nYe7nib7BizesrB1ZcDh+XkUnut3CZ/yYAN
yr7WqgOlWIR9qT3oBD1M7Taz8jvlLPf5DK5Dfd53JS1XVlt+VWC+oAZGiILM3uBZ
vCYis5gCUa2Ur76PTu2mPZhRh+P5MYvI8r3TLCNHKIMQAkAKH4bkJTw8RY/2b3N4
6gFJsAMy4UmjrWe2cUhHIxDr9ZDC6oDpcD2xoUFx1botAwBWe2cBfZBvtCfzkkpx
MBVQEifV+5CVBp2stLuiU1Egp3oq7+Mq1oxLu+jlI2CRv43iUMsAKm1u4AmhexBj
onLHMoAIPpcs/H4l7crsmBqV2nGyODeP3SqOB7solaqP5J/oZ8yEGjw9F4ZZhcpM
Md1PD+hpujY3ZFKwYc235SXo9zR7HVh5EMu+krZI+aahOfrKpAY0+7RwEn5CUlhd
HaCYTUWdnmZ0JNscUuj/bMuNYpbN32je+HVJGDA7WJNRb1SC1O5p0guOyAf/Z88x
83x4EbDomZC9sSo3yc58iGrjJoyd8eQx6tXmW9c4MFpyUW2PiW0FXlIwYXlRQg5x
mPoYGVsdGl5MzpDW9+WwzeNdoLhIK5GfeBU1ZVQSbclA7ZrbLmJQ9jPG/6aR7sCl
PgJtMQhERRklB8Uk2TWw7KcXai2S/Ugb7tZWhVnPBiflFK8L7HfO9Tj9+N5ccZ16
I/aRirKOuYqPcZb8PKdt3jOsNizwP7zWsW+aiDbcoZ196etn2hOMibhsNwKHECcJ
MLt7m8KyLMiSB9RGd3rtpgnQ2UvdH9Vwsg595QKQC14xrHalecWLWOeT+V0FXgVx
UM7bRnEQYIrRThl7lkiMmerA8IKW6dVZAcqYyhowfgpSB8G8L7WfVwp7fEBeVtsN
4ZrFfxS+sDgPKqFmEeysc2ANpbLZ8tJv1AcS64mBBLkoOFs0LQcPpHA8hQoyCb4o
ClObGTx5fei8xydEGfwl7zzm43OfUloaxxFIdy9PPKZWAoSBAiWTV523oMDhgUkX
5Ej+at6Qarfbsj3W6rc0BpWqxkgDTfkej1abG2/+EvZmH3Sn9lUDZ4eo1AaOzZab
lP7hUPXRL59pQfgJZtHZnJDtQK/grRBEEMBSU6a6inbXiV8ZYKI4CwW09q8k6rp3
DKb6z6FLp22U+sCG/gZe58p9y4T9ecUsXEFiPfuJL79pSsaYeCBOy2mRfqBrGAzg
NGW38VY20IMz8tlHzrlzB9V9ve9CGLSKele5XZyk1QCWU0IAm6XSzeX+G5QHHxP6
UCuZ7hs8ZKFXxtuc4N6U7U/wDzliqGAMi4Y8W+NQ/2R2NodJxx/vCrMsaO2FBQmC
8zcAhDk7Hb6MY95uyo/BeEvWcjIdS6/l74VxTGiYi9r/WMNCXFvHdqsTCtiE3SB3
dKcHgW1UhLp/YnsGY97G5Qsg3w3y4On1hzFi3QSYmH/lfgaDO+IZ/gv5323JtsPj
NnuD5NNgF0An/iKMEhLx6eF3I6UocML5VDqZjUv6dtX4cL7P7BChEJpw1hIk5xY5
1B33BHpPt4N4YSiIe+R9yG3n+9AQSQGbw5qfbF+wYQFuSW/9ayTOqciz43kSqZzO
BUevFTEPjIu4U1qj/+c1ITL7WOlYqv43h4l52KNt2ZMdOmvOkf7dOqWMu32pyrdf
MRJj0VMUiv03QOdnSkCPdHm7gHbNqIifJzB37jepTluGxsJTCBDwBF06xSxUsJ+U
2PPOM6IBwMKseU082leP2pTBXpG/NPUugk7akTzzlRstlxzRVckok+bUuEOsmGJT
IYLJ2KgKC+FZnl120NEkRbcFtUzWhDptBZZqJyd3Xoo2ylMjnEnmta/ZVYMNTr1r
ov2ctcK54Unel1rjwTyc9KxJETgn/iP0ip9DKRfkJ9Bw5tTvB3wJoKfYrn4cX6qR
EGFh/LUuDye1ntCvFi+eM+fPJk2j+VcmBGqvOd4MU+6nIgQEGjPVywMZ6XX0zQcI
u47xKmDAKXW4P8S4g6W2M5QrPJPovt7Di5fpFRaMNRtQuBd1DaOJ70gzR2+6muWJ
4pGkopENWSlS/UWvCNaUNQtCKgQMAAnlukbbw0GML+YL4ewvFGM8eVxT9IAqB8EV
ByvjRA3yxUAxnT6PbSQZxnXTReBA+nZb/FvNaiMbGgfZSzO+pR2i5RfC3iPdX6M+
lcpd2I1IeMlVrynUcMSZuXaiUjmVIvz3nujHEsU2AfG2VMeep6NHvzvqgehg8zgk
IfcO1ID/pSyuLkBmPmTit6kKpaoFvYjP4nU7FBfyaqRpRjfEAhp1oaWRB1KgL4sB
ba5dE6UPAsifLkOj6OLED7/yOnwaV1M7oHc3/d+jPLvJx+dvyI6iMeNxIbdgQ/ib
W2yxjRiEn2QWOdJKTc4Kf8qM+W43nZ4p01hLxnwZCixAfoKxCvypL7NDMqMQXRT0
WQ/2/gQttCbFs8s9mc6pvC4/Qiz9k/iuq0nHwIn1cglrL3IHGx/AiD1ey2PfpncJ
eGai588NaM4jNGPE32Iff//LgxZ9T5yHLuqouz6niVtgEey/cWKe5SqHkCFY0OUi
YglQd41aDDmpNUYGE9WWB2l0fxVZjf0IXfjTCgeg7Xv82qNo7qGiDTduDuu9lLCx
TA0S1huJ31tJpeMi2VPSLGJht1Jul5sgCaXHNLyIpYoL36Fle33BSHKh9pgNyFNU
4tCoYXjY3oh8n7wZnTHv8LyGk/NLwFwMAsv+qBdsblrq6zsjd963Vaec3qe7Sz3B
KkiYF+wQGzE5PPM8HWu4zysZ2lJQmSYmXlDammw8DqC0X31ho3z81HbWxcZ2nEsz
sOIK1nY9dWmG6LmuspLquLftUGe8LViN6mN2M+p1lNaoim3LxJU4VfuXrq8ellSP
Sv/pqnnf5r2HEnuxqgPflrwQrE9gw+lqYkRxBX8gJipYanT9/aUBdgtyGV8LGdIo
5ojsI9/23aM2ABN96vsTl/kKKxTVqlWDRuWuNFl0gkcv4/R7gn+EEAQutq9dt97X
kSQL3vR8fvIyghgQcumgF/7XoYMdAZN3fdyHqc0J/cVLuUypBfAHu5AboTo/BooI
3/1vOuFitZPJKGh9vdr0YzsHmM1P9ddl7WZZozui1J/URsHqvJol94ruQhj+NI03
dy/wys16TKwkv4IXjH0IaC8yt8fD1kGuzG6UTjRdcsbF/LItu/i/HqUELoUex/qk
sJK03PmbKl1bxUsGbjXq9eL/TMtc014DP370jfKAECTVY4FekoNgDdSph2752dFU
NgnJ0bldQE8x+XJyUQU6x2PZTViw2L3oX81oJKEGtvkwcWMfcZg6T5h8wtaOneyt
LpQ5m2Qtz0JDqx2nIv4Mtgq9Hm33f1KLV8hcPqq0RvHk3+WZPw7BCwVyixe2x/u3
5bq68cjNolLjVdFRflwBG66Pj0nwPPUmnbAaqcT6gEditppwh+QEELXyjtaWQCrH
QJSsxManAXSnFmdyu1OdIYjJzwFezwzIFgLM5VwEzDT0+5I/NBlIoj5VeXW6pQZc
HBwedGbJEDwA8GaKprzThq1cydFssm1+gxp/dvmKrM0RID0m5JjBexf16qKMbYGO
YYYdQ+rVB8ehOsMUL3imApnULXq6zu2VNC+YMj2osTl9n6ZsKRv9VpLLJ3SIFZhI
/iDIU8MUwT/o1351XBYcNCrhfjzn/GrBcAsRZQnGMajXQ+wywX/EHJ9NoltRc/WI
DIRxA8dkuJvrU9jYHqJzaVb9s+C1mv78e3nSaQjB4tvCTLHUiNiKRC3LOnzDbMku
tfl+5HYTefAMpb0Ga0zkT/JhFbnyNl285RZM49q16TUHNtkbbwJbl1523sbdInYa
PG4PUVDtnKTbKAuKCAOZBfG6rvQGG8yf/8VNoOH8cxBnqe9XAgilDO6FA6RUy+xh
hyFQlx3c28THuQ3GCTCPM3wErjiN51za6dgfQg8ZIOSM0Om07MI5t5Utt02dIYCO
q7GXZ5kHNs6LAvSPD4LZrEzhwLQlpzJranQogSJcfLYGg2t3XDsdxKMNrKnQUjpa
3N8IETXqX2UZDH4dM14Rn2Q2Xz0C49bojgYSizYNOZSZbWDR+gY0LbvNjPaYLrfI
+HiVwzbaVtt1tBzdpGDiwZWS6IkISdTnnSFyPythPYsHrTMa/6Rw4ykXj12i0XjG
3NEH5XXwicYE6eQgJnpFSM/EfPq6ptfnVxYdRNJexl6dfOyyL6is9LUUYA/Ankm0
9AN1XOX3ez+BpH0aonvjPEFhKt5WNxjMQExbXE/16pomvuh3sB7YiWwuukW/jKgn
6EWFZ8szUpUkilOx5VtuigXfaXW9vJxoGJorIiC6pvbdlYBFWBl/IJohm7tfHMSM
8UVONydoje9GbS29MCWc/MOjkPWz/M22IvVQV3eb6j3r3dsxM5ip9gRw6PLst2/V
TnhrzWq7Sz09RCkt9Q4pcWti4UCbS1ygOXNWYxu+4Fp1KF//5uVRJRUwxhBXyKj9
67YrvEOdjLEDyEPz42hpeaiwRYeR6CJx+lJf6OsQJqI9+eHkey59PneTvEEit94s
XlvPD9TAf/PBYmKq6ei/07uMHoiNDVsgpK54/4sfcfx3pr+ri62pcFG8rvcr9KuJ
MOxpeIm5wZrKtkzKniGsCRNkLoBZwgJwLxudCIqikuJGjokAP8yXpsACNkfeIkZ1
9FzDOUoQdiOQpNwWQdh6j44jFTcHfujqScPwZnM48jGpMerFyDeUVks0X0KoFizZ
Z1vyWf+rskFcj1k9qwaQM3fM4ObAgpJS5aodhwR1x5xZtuYLqoFLKbdErF3RYuN8
S1/Pmrj52m2xcRb+kFIT3e9+9+Xa0XJeeip3nUsMkWwGm4UPmbY3XtL9H6LqL9nK
/ZWz28/umVZn4xUr8UiBuDqXJrA1TMTstzPkqhhEfJv3Xn5UmENJqKc35omdeYLP
3bD7Yr6QO5xOSbouhTu+LZjl79bBE9pMUm/yPFebQ/HJR0fwggSfSgGl73yT+/tz
vJ26y7eK9xn6rZ7HAoHOZEDjWockAlaq7BjMBZkvaoNV6o/THMxOByIEujrAQ1IL
U2ebYh6pTjzGjn1P0RffW/gsyXQJayL6aiU9/k9MkWXQjajtOk+LMjFH+wWSrrZ2
dqIO0k9Et5qh7COq0A1/qmG56CeGMFLKhM4pCc8a5200H1b/+rtqwnIKJ7RIRFqr
Kn8KBMDVbygCcZtzfdK3c+bLyGqbe3GpTwJ7w+bUwz2NW6N/varUjIPSxJNbR409
2HE71hQqxN99Ewews3V3vloTmyN4KvTQrgIiP8NmamYu2p7IS2uNL1WpYMfUwQ50
iT53Gj2bwRMCX+5kfSsjPM0ZK/D39eo5fvPAgCUvGSt3pFKk/DOYB4zMnTN5ws7+
NOs84Wz3oN2PKEdJYMXP6NRDNJwqpXF+WN823rKgKucSKq2P7P9mW+0jBJ0nNTUs
5CKJ1h0DGALmKSHabGJ+oOF/tI3+SQ6J0v8ukOVNw9FIRgJkrEPs8N6q3Mkk4Z7B
ZZJOvn5dYdQBXjPtt0DPZLSYlC0YF+uxJhn+m7ALyKRk+UcrN7kbJIpOXzIr65N/
SjRar+HNJ4kdzrGeYF6qb+rIRilh7jDi7JAVbiw5AjWJcHOhaysfPs0uljTlTAix
JqnAzXu7DyzNnz7axarHMW9oHqoyIs3IDcqtaWcK1j2YcoHAkOnZwFZUqY1darKd
1LJ6X6sfPdfOCyqO4O0IkEXE5P0U7hq9PYsJGSeFI8tjng8wRTffGVH1/e3p684U
7PcbS8AUJsmWt+/M4iYubYq4AbUK6dMsK7mjoVrN3KqlN/lT9PUpfjsnD03IDWm6
J5EseyNqTzjZZBYXA4R+rabdSMoCLdClsPKrAnN++EGA7o5aZN9ozGVN6Rj4tgtG
820xfiuwe3jFsLjGUSqpL5QoGIp73PlosWsW+R2E3hus376w+OJSjY7c01XYqvvJ
7xrpSmJHn6Lp9LzX8QlEvM9kAm2QIhiYnQO/7Of9Y3v7jUJaT9ZvnDqVT28gsIXH
R93v+SA8ddMy5hXacDuotqgNEnytelOy6HloK6TZX4ivGL0e6IeVubO5cf2kZ2fm
rvPZU/TRsk8uk8phqBGC8tpDfXuK+jMW+Ngkm453KhoV56q0lSwxnLQK7B0rTr52
XzIHCItpnNOWT9jpBFpgV3OLPlusiYYn+FuaqYEJLGgO13nxEDaG+oeTXnGpbw6B
SPhATw2/hGP60j3nVvRMifwRO6aIfBI+Wy2JgFxQD88GxakRP/lGStVCdmjKCQD/
FOsE1xIZZ69AG7pkjx9E/VH9B8MmCDAoAqp397g8haQNjm/t+Rsajhcf619QUdwq
HUYrywqymv18NRBaVqiY//ESrOYfy9IYn0sT667jYJEZQzIgz+vr5AWSvUpIr0Ba
72PYvh9q923eTMEhPfpcnHpeoXlOFTnD48p8B+/Se4XSw6EMxCUgtBnclpi1tCAr
ra1hzBF7RN1KVNAxmHJ0nx7caVcgPqQHdhziokUj9eI/I/NXFth/+D2l/uvaLOKJ
TI028r6vT0FOqvogL+MUbZUzpe4UNonHRR+oTnKiNtKeX5/3fzG1XwCJue0nZYaZ
e5jjsB6Z7mc161rUuhmv5sXbepClo1nj5CvAywmomy+72Al2ocU4XdPRvdxQFvxi
n8pxe83gJf17QleRXw/PVyJMWajjy9PHQyjOy2sVtv7cThxKQcM2F4eFb4/chhCI
rY1rlFfHSmxYAqSTtCx5WWd/oiKQ9+De2rfMGDlzlipyBxTIW3t8WRe/D1UMaEuZ
0PFTP4GZW9XcLRFO3GMB40KRl2t3fODi9mgeUAKc3hngN6/ZG4dOeBFOBkpwxdnD
UWia96GAxvknjUeazNd6U2oUBOFVYj3pqwqGmHlVMgCTJFzi2TY/azPzFe1cyGHN
2u7j3jXNMlqTpQ+Jm+b0nJE+bt8/dSG2CgKnqJSGGU9VSk/hmoghWBaSYWuiGRF2
0pyFO7xz34XDQ9P1By0rxMYuZW0ambSWRP75gekIynv+l/VwvRvWGxRxKg5M90t3
AXHYW9ja+OwAsi5bp3rs82mMIIxzF4H1GEQ99wizuWwuZ/aHwuv6BrCCQGlOI9OW
bfG+Ol6pDi7sXAcz4xYdzwiV7TM5NL5Dm5dSUVO2Z5vYLMnJAat57Aj3Xup3KEyS
qKR30PlkVFu7cCXEhMnsw5VHR1H+iBt4myOBu0HwhSH5toFbYUmqH9cWE6fJlo/W
Mo6k4nRXCYHolj8QyWNzD8J8UAYwMRki+nL4LK5tN9owjx/A5Cl+LQbrXdbWO1F2
kZQkx6vQf5uR4hQwxHeR8hGHJYqrlDDCPeE3Gv2/wo6LKeMG9oJlWHqXWjOdKj1h
mj1KRgZ0MT8wwCzpnw3n1n5K4Z0z3hoIb18qr2+QvjbSrrFnZWl+JhWrLASYi49D
cQbNwfOhVShgGT1uDcxvFNEkgIsE/Qrb7nLqcln200QJHdOiUdx0eHVIEC67m0LY
LHn2GZRltVRUfW+XnkEyG/BikbYjTq4tge8lmxXKSNj0mcq1d6f3gXB0lvna6jJn
MdRqesZL4DFMji8vxIHHj86taGsUUOLDpS5mZNRF7gUp1x73Cq0GetvDvqMSCYIg
wRoZsW8OBoMqR2kzgVXDAJDHfC9fz3xfGtYTXrOOWFXthcdpgHSeNrvp3FR0CG55
1dAXf/vBqsBC/7llX9VyBwgvaP6lEnjZaOSZ1Pi5/aOerCciGAVphV2WkBU2p0js
rXWAkpzyyfwsTZIPIw3HTf/bOPKPGEulzw/OfwZBvUvRbY9xDQfxJdE/NVxsPSoX
rqWnNcntvKfpe/FIVWiuMc0797lS7QreA1vIbOGwR0q78vAUL824R+TSKkcIZa9R
Hcx4eofGlYgIOCYLXNnlCc350suSOw9MHaM//tQz19k092pngZcJlQFKQMm46gg7
aqCTTS8lsly90wDf/8B0bfmvdnweWO6kR1ykVVTsgfKxbM/wB7mQqG5NrH0Ota6E
+ANdkrkuCk/DafUHsRdNbWmwA+xs51j9QkVyZqVpg2xtLzW7fYc8EHt2AgPP1trN
b/oH4FyaGFGhdZ+JN3gXS4Zy1mpfMYvUyOGzKD6I+Ux7paSeDN2/0m/uYNu+qCB8
XbGBoZpuMCcM6F/+6bBg2MzAl1d59psFbxW6cF+4+vMHx+PKYcqiixKe89SIq66d
WqiNE9evAqRigUmrXmfbHmJ47yVkmAGOtMhtPFtrI+pBt6a0nVtYFkdg7M/1AuFm
LnKQKZnm+D7t+fNY8pXfgZwCxSt8l8gzyivJ4XEJ/bkzoVIbkjatpvsTe5o3xOu8
CPkg79mPN0IDo9ZGBSXQB9JSYsGPqshTDmMloaQl0mPXxItJ6n6JXmMa53PyhbB/
KkCeHpPqtU/87vMq4hRToxRViBnj076ISizKvJzdqYD1mA8CVKs1xEQhS9fmvStw
njWlCOfhJKwn+chTO3JO9LscAbjsaDaPXEDm7mrpJSi1EONq1cZz7pxvafImhq+j
dLvOXWPh637iJx3c/jgZL7FmSJ4bH6rwbpGPXPLqHgdsbvPPrL2in6hRXD0riDes
00ddVGP31WdztisEQr3N3a9p9HPiKtidMHDATSqzf7FsOw5ZYiaoN5+F1sTIJ0ew
XWdgLLf342LkTAv83cUtZneX2VFgxmlT0QITdp12aTsaGB/1+Zl46NAprM9AznKj
f76oDTQEAn3fsMNUOBHpDHuergDV5eP+3JsEXQUeghVBZSm0t35bTngFqC0Coa6C
jYXltjD/ekEGvpEFiCQkIWga5niEHIsJWexZXzlLVsH1UC+9DsSWyTg3dJN/Lj6C
CJddN3TktD/xzICc6froX8TJaKz5n3DBNMbv4EZIf4GTQm99BQZqVyLjgmSw0CRN
0T3XCSAFtBIBCuhqHisKobM6nXPaJu3n70KiLdVn8Ta0/4woGwrn8XZx8i4hnGa8
pQA9EQnvSmrsOAr+zgVKl4HosENvLpdoWsVswm09JbeRenVjmPi3y4u+MW2gF/gy
u6V4CAtpSbbFkKoiRXTuFsOvkOvaDT7nRb5IcfnSRfauxC4FFTOp9AMC83ElI1pl
IcVMnpuUjggrmMtd9xBXO+y9+i541IDRK9ZoC/NXIiW9osWJdcdt7Jd71ZtnAFQ9
yW+VvL/iP9UPVg71SrvnOYbHRx+3KFwAZFtOoItumnTALJS8jY1peJT9KOgHB+Rg
Sa2r6TfC3HIB/A0dO2zFENdZxAtP92MknQeYt0KUN0GhLfewcUyNIrocOQ72II7h
lbn7StGxVTqtxr7OHFz7XON4JbbaVHDXrbsYbhbEHBXx8x67jbPlCzkPn82XSMjm
jE5Y/zIuwoObbJH5F+IEOm12Qj2bc8rkGHxiha5bNEDVY1VSRd5vOBtHEjWXD3DG
Aci8LnBekGb9UKuhQKqlGZKB8T1j0Cx7agE/mpnw56Zzm+dsyNCcsGZKBBg2+qt0
al19EfIPaOqSpRx37gyepxm4K+O2eR7AJMXQMDaMl7ts8f/cizBwmGGpU+7OgehX
KMCE250HSWa/KMhYNTWXbFQ7okM+EpClHgdDcfjoXdnxCRSnoW+LAjEV47kf98FV
6aXAvSjwoETwRExtPfOjsYl461gFph0zcK12J9gc18Doi2DEoY1P8Y01lxkIN2JB
BcePUkNSnX4CbjPwt8+gp6AxekAfsNCnhwhyttlQt8vmnwWWOoi6VoXJXLMVPfTV
MNnT259Yr5RmnNzTtgL5cSFAusS95iyBIc6vA8mdBFQnpiuXB5z082Zq4WxdnIcI
pNHVOu1ZrsTK9ADjIQWA1TV9r2G1q+LPN5EzrUgOCFG7kvg5hBTiJQnv+phCIDV/
oYoiKEtaLeIHFygb2RDcIGl+cs9CWFR5vPeI90SC9MI6mMOyCcUGaqn9gtN2kWpi
7ug8IdIIsaJtIIhSwNQ8JuwILo6WiFhn3q63aFDMrQ+Ez2Nl2q3rzg7fJppex/oT
8SvIR5e5w3NGbUZAFWtOIdySF4YMTaGBHVHWW5VDBfb5Jn3A3C3tizwX5T4bHRd5
Jjw2IX1RZfy5K5k0tL6Y15rLlwNC8bzW53GIyyWP8wiBcx/QCS0X6pe1Kqb52L81
8yUneQgjTB2Tw432M20APAkZupYUGleaaQRfdCeB1oED3N8OUg7cEdk2dnBpNC2F
ad+Wsaemzvnx5VgF7LPMTpFglrjycEMazBlbJ7oxCGtxj/4nURvj4a8SgDAedBOf
N2cgl+t3qtKe67RRi/X7ioiCBj3Ya8vPoqVtx/9hk6nQgkYoAixGTyfo+Uoq9ho9
ytSIsGVSZ2UFyL23QEmLNXjYAbKnf9vuVOu/j5QHk5mWGNo3qjp9YGDXNMbxwBhu
AxFYFjYhcQUUF+oUmXpDoOAWR8ciMvCYpf5PHV7GfTHKYDeuT3CKUElDnpZUgGte
CZtogq9aPEphc3Jgz0qitHc/l1rSm8GxjBjG/xqy8xMcGf/4QzjMkUAuCQlfz4hn
yxFvdtXbHV+Is0Qw2jo/2oud2TDk1IqOKyQZWaxbcwMoLLIzBW83elYrMMwTLAC6
6G6NBLuF+rRmpdPOnpiU2oGVBRVCT+OBrh4CnAcok7cZWZT4dsKcy1rfCLYQfhlt
tpOwwQptU2k9yx7+w0KAXNy21HQCIEzktELKPugWB/vIpP2gaCmILUZyQuyZItMX
z12URBiS0R6e1b4lbJWpRm9dxgtR8n7Kz5cVx+Wl7FIdc1XoVdE23awtjck9B8fc
dGOhukRuZzFbO8vPenat9PpQdWn9B5coPQbmrZvCulJ2veRGdD18zbjBweLGgPaF
Tpveh2fhu18vdXQCsNPjlGg+cVBoMnIEseiyVlnTkVTSEiPGlqtBzbzAquksn6yO
vVeeBTj9hpNf8kK46Y1x5uXAVQmhH+8h2Tl5lJsT9boLT+ywLCt7Z+53RqYFXPMq
LZ8IE7yoSdNld4PXFO6+iQwP48mFmBT5fz6Hs3Jkg4dtIfSgTlFmdz7ww25R7TTO
Z1BNYJRwUy2rWD3Y8+lqRXR7Y371nb/RjX2OXyPM2V8lQsAGRY+m4plm55yPwJ3d
lWOSZIhHvJ+i/ZcfGu1Px4xOcOYX+I4h1M7+yQcq63gtIECgFAeoAY/uBq5HaI/n
WOx9VJIiktN2yNG0b4SQGtUW1JWk09YXXPFlAfBUqCY2NjkGEixhGi2+Rm3nPJZO
qut5NELBQ6HOO0Nym+Em6rMPuYqibn3in3DhtLLz+UBjxFWV36a0MLycU2Z/7/PX
WecMi4LqbCJJM4eXBKD1OLnmozgRigD69ewiYWrAxjU9U0KrGwemltQ9JRNHg+ia
+9yRBsfibxs3BL0KC2Zhi2lAl0n+rAjvKXeTKKxmm+jqlF9PSD9dSmo7qa1p87Jh
k3VFUqaXEuZo1ePilsh64TNY6G3uW783kpDhXMZedd/ernWfYVuGI0SIkCtHlUOu
GH+DdSnw/XmbP5XKKlEsV5NVT61y6Px8cQBAWFRmevDKfSq4U9aFk1ftUC8cpY3o
5sBKTSVwfYuCP/wYLya6cAQQxLu4BOmVYa8jQD4lx+/jif7U3/Dq1c3N9b9OBJ1Z
7qPf1FWNE5JDwhzPIgVf8GfI1sQ+IuH25dTqXnhz66KH5yJEiQwxnIr2PIOQLw4F
Q7rk1+bNHPhE/C53mgkJMl0KAogqEAUQgGJrnX5qm8a5nzoHtFBAoKQVs+pQttMZ
O/TcKHY1wKVMzOe4XX17xG7RFxa56FV5mY+GTRPWLjCO9FgWUJp4eInk/CR7Hzxi
tpA2C7YlK9io06v6Pur0Rg9W4e+CtF/RS4H4RAYbMo5QSfculzMpBbKuLjj/JyfT
mbJPjG9ZORt2iarYVUhXCBHIbHWVoO3nn9iKSV/S/ExJzWOEghcyewsNAb1vPKyn
MG6+x0ml17lTqZThw6bSJcXIUmPR8juIUOsK+pyQgwYqlgt18Y+9sItPTsE5P0BK
g4y4dx6e1I9kt41fg1qfakoHbpeP5aK6ckhiRlKbJh6jdjoofkZ7zDjORQIjtvbX
HO97yF48vhEiLE7PCpLt+dEiXHt39XEKcZt21LKcWoUlUzJRFlZzYDaxSQ/msWGE
RQzeAckaUuV+7vMc4w1fHvaQjTkUVVShppsdTDvVF/rxHbeI4SV1IZDfo+00k0Od
3Ur0sstfLE/NQAtzlJjXR5TAPFy4rTGd6SLDk4zObTsHohoawvqaSpYT4dZLM5PU
seAK6d8ySz9TTIsaNYxE4hKakZC7IqpnzkOj7XRLsLXX8jn04fiRE7t6DHaaSCpT
fe28qn6AjUJ3NWaDvAyWo+9w85CbOZjKvD9AmxLxgTpiL4s/FR4Cyy4aNkgA1v90
YImG3pEvai+S0TPTBukLRycAoDYzvGQX2ZpOsWoOeReKWxeRLTn9HEoCcsTAj377
KE83WKkYuBK0p0dU8FpS9lixqrLRNtcPY046gSy56tnnx+TC+KoCacnLhrNjKfvd
ua9dhi4v8YRk4HHrSoLgmLVzfmCaL7tZspUNAZTwoLc/2kwafhcXdGYo+VDHbpx7
0i7WbNNHa51qaut0DGg2UORACl7Yy30xO5SDpRGEv+FjxZFjYCg2HtQ+Px5uev+Z
aEm9uz5zk+34n7FleTlLDTUlcAKVMZb6lOvUiOLcMtGjAL13h2TSoFKxEMlrLC2L
/5jC2aiq+BiXhADZro0dLV8dE4JrzeujBaajbD3LLsz+9agGSqjv/7LfypeLyEGv
PevdmdBNMmcRg7GFgcq4rIkFx5NAForHl2f/UuL2w9Wt6jShGHezci2bum02oEb3
MI/wBSkyMDC5zewHZRvVvEPitkAusgce2wBuig5Kaq5Mh2k/tM+acjkhBuD2eKR5
R+0SlOtyR/WAXTQYUAywcXtosYcfIwLtorK0ZsZO8EmtcOyOAVhAO8rqhdtcsJSy
BZ/xtGFqaTkOna4ntpbWz8hjXstx88l0/yMd9Y+HwOl5y+Co6HZiTuIqvUtsZWWB
zdW0NOHJboTtxDI/NNaHQbsn4pf2eM9OLzHjgow8EaRBsy5nBWdpbjFw0CWShAlE
yqkRQ03bc7Fr1tBpc3IV5QrPgQGVQxCAK1MKJFUYLaBw2yCe6VzMyznEIS147iKP
kL6qmaPVGo0P69i9k4MQsKW/GX5RCNIXSGm6zdm9OvY6DuxReHwPQUXy06TmXRKd
tLZgsO89rAJtHb/JwfGNWbkLlMYw1lfM+KVKvXko4+kLgYo8ZgYw/pR8qO8wad9t
Zs2Y8+FvE41MvAmKY4qNwl0XLir6O7jDVgdXJo94NRZ88552kHXXCQ4CwF+zRQZR
bDpUnHrwVL0AoMX03w84Z+uTvPI5xP3m/6nHeXkCD+6oGHhdI4oa2Qzc8d+k/RBh
DWE82WmVJefr7lJAaqBwRKTMhmKkrVdLcS/acLM5Gk+mOfMe84y7gWXbqbvsKtU2
mbrwC31kr9IYlpPoyEt9Fu27pyBeaSNXmHzNojkracXf1w/Tvg5gqLLpif/0jTBB
AGIg9Z0hCGw1FiqNeZfHu1Rcz5Z8tcB+aR4fzWTTJXhf9o9iyjvlrrcz/pVn6PdE
gHFyDDcG6xq9Hj11YosUc8gfjHNKDHmHD9eNQfj7n6+64jDTwnwbXbQI5lHnAFDJ
O4afhr+dW9DEeypvqHPpL+Yp2v302HNk5ISrpuqEuOn2Nr3+L06Ie6Z3r3RTEJfU
I6oGUUN/F7Ickd31z2oKxxCUYtRFZRYSueyzSs92ZbK0VD8TCvNjVaMtisUPd/RT
0tjW81iEkoY8FOcc4ubdthFUAIvdTcmz3dKT8KSQbFEbYMYsSGxMD3OTluzlg+Yy
2Dx4eQEzO1l6uLvuslpFJ54YE+z660aHFWe//oHUmUGOJP5v0SYh5K7ub4C5vh1V
DyzxISm8hwQUrouOAvQTPOaYTQEEO5gXYqpHMpNNTrUy387eVsUr/2zBZ0oInvG/
t5lLn7ACvnUdbFPs9ohOIfZ81BbYr+VNRqWkBoN0wux39IBNjhGhsYcBmLoQc8Rk
fM3rq328jgt9gP7liNeWvvC+qGFasU/Aa8kumrE+sRKPxAn0FE/O+lkNXg3lShRW
ypTy9rkusvp3N4f81RCFgqXXp8LAB/EnttAEENurfSMh0FZWMTVWjG9IZCWA/usc
4KkgKVnwYbUCatHPf+GX5rQJTcS4jgg6XPCyBRTqkz074sA/O2Cx84wLRH7MT/FH
8+FPPzoGCfJl9pKkuHK03w3tmRhcnVOjKpI8M4wp52AdZl2Vc2HI5RRtMSSHjBn5
RWNcCYtdT1yR2PX73Ydh+SCGZBOhjUEjV/wMH45eg1JtGWcNAh1IrXaqQqQu/7sO
RjGhf6oknsVw3piBpCBI6O1yH2o2qzMZCszEIeg0ho6jHTOrUUb0Alx/mw36WhQQ
Ja4jpm/MkTTipWzTOzH3eGlUW8Jdx/klmhU8qIZrffgpnCsUoyPN85UI1sQlsYuP
oE/3DKnu6VKEIxJWwA5mSrnihnGyqSGs3BtqX4Lwwvx/lLXEesAWSwjHo5meD0gx
SkH0E+uoHJqDSlJQ050oPpv0almSUmsrM305FAP0jK4ByNOlsATMfHkXocs78Cnz
dY67ZoIOjFuiyefC/t/DT12IfrJQen/E7lyK/HQW3Eu1OtI1sly0JBnQlIOK68/S
unrmfBr5s0bO9C6HGNSZFfE5OMKbAB0F8Bt5P06y7iejGUAQC8YmNZq4ryRXBTjG
iKYLDQwBAIHfecFjVx/cr9dzua+numTIRTWhL1QGWt3z2b39WHgHvAutYcGRqDAR
G8dcRTBp+8dA98QDgnxMRe2w9ReGcTDi0EfA9bnC/ZJF5YEVmxNteRUFRgC/pVLX
/ALuKN5CUtOpmSkuJ6a68B4rLDnxIIBF6RrbLaobzvEAL3RdqxSfyE3ZZHkUJ4IQ
V0ZVQD2pM0yNkpL6rh0bo0NclgCfj+nojwes32Jp6kax3ii8pnuA8kImsy3U2zNx
J80yYL2gPfla31IDGLvpqDeHNoKh2a8dR/RhHtJMQeAepO7KGhjwAq7fnKs6IjLj
tjpMVEO6W9/KYkgow/O9iWFmF0+j7KYdrp2iHDxKR9imgY6ZhNm0Hr+2lUM6aMuZ
BXFv+x531ZeYHcxBgfdpP2VuAxrPQBrBlT9+6UV2mAASUJ5/Z3i023vR0bFIY6E3
mIQh2hFngvT+HkKmn+CDeWQV2FQMe1jnE5IzcBVbJY96ZQzhxrVhChhpy4hvcruo
cvH+G+K7ZTzHM6OoyB4lsQcWyMN0zwGB2v4Ne6dT9xQ/36Yo/H9Kz/+RqgHG7dg+
KQfHGwZjarifg3h6QaHuaRdyPs5qbHT1uqcpg4/QTyo3Gf+mGycgRueBh085mUSq
J+6KXDGy2mLCnXYZsx1CNstacAZrs0hQuqBnrajFbDzgm/mYs571ObOiN8uYMTqb
1MItxgVh+tNnFotFl8YkB1i7abV+7RhVb+l4zRDbDnuo7fOWssC00xCS+qCfYKRL
M1RkUvKyEBQRjKrCXzIVlJJONTDNP12Wqy3kM9eKarAC168SbFL6FnK4KTUw3nRL
cKyDYxWUPDLXMELgvrlOS3uOFDo+mqpkhRWxyYXcTCob5fwuSUeUIrbNwS0EDRvO
ZAE3mq4yWH/3u5y274u224tJ+MNI6KADGHZKwQoI6emTpMOpnJYoEdvGkVl2BCQP
qExRrJxq1MDYRuy0QmORP6u9Yy8SCXfIh5VOYiq2Yrk/hTSeL7LoNarZiaDUQ3Bs
xaJAuvjGTfd51sL9ALw7mrDJTMcsNzL3SwRbKw+S4Di01Ua0V2tKjwbDmq/iiW/f
rqA9Gtbb04c8vUj2m2H4tYWx/KHJX+TC73wRdafu9vF8sIphJWZ675e1sN7ot6/e
Qw7e8fq3UZgUElGWDIgfH+cgXrP5UGyelQo+LhFFUVCYr8XTF7ZtUUeAXhCmwrX8
KsUhrWm52LoaU1zNS+keLMFPBPb7gi+0km/pjZR2/09gmBQblegQyzxhn7CSkLqk
vagiA/381EzXFuseuy5gDShBss9SFTRSuL6mfWHJjBFkBt4IVX+H40710h04wG8M
3UkDFVKf9AzCPbGcQV6NI2jYrf6WmtkpoK074NUD0He6lCHzTny0/A8gsxmjK3nB
xTlQ3C/wp0zcsqZ9bGIsGdMXdsTKYaX91+VwJlEWIjTxMOLWzg6XbG5SxcHTICSo
nPxOHG3RuERK7jtohYtgoClq85IN8OjBHFUnf8ky3IYU5yo1/4C4tz7UkT8FgWk6
KBfyFzxUgmgrDaiMbHDmxHgLA0i3+8e877bhnSFvB8UHv1euwMOLnSzs1U6zkcwq
uTjpWIJzEOJd80CdEFkJqZZmiZm6XLH1K9dBezri10l385u1eEKwp/mEbKmUiZwZ
g5+T+pUHyJ+IbQSlxXatzFy3XEa5LnavXDkK8mBIZkwhPhq4+rhN4h8c2BIv6QBz
JcoNJQgg3oldElO6IBhdHFXjXKO4G3baZmh5f8dlpMYrsNeI2rAZXmILVvJxD7fs
cPSCp6FFaIQjTu+hSjnQWNGYelPBLUlsnek8EbsrSm58oBugGnlY6EmTbL+2kvkv
v/mdIzRm2kqnzhhv250rwm4wNSd2uIoYlkegnccRbHYkGkgHK/0beePGGgJXqJaz
CrtaUZTFNLrUVX+ZBwoZd52/YFivH4LyEe/aqrckQ7bsZceQxhQooPKjXgcMU0Rh
qv1UGXTRmhaVnrTeJaXhO+tkFQIYRH/Lm1ttF0ZXBtAOfh5/UxQUxA1CQgyTnEFe
UXZi2/R6rnweytCmDcdjbMaVfedftfwLFd6tJHGABhPNJ6/ba1Fmt/lipUWSDMzW
khAJRuHBPCiGZ+fTAooXtyK6ckx15qvy761yDZu6SXGfrPSoVjpZKF521bwJGMeG
VBkIwu0A1+u7VYzaZvqpdr/6LlUW7w0KXpHyZ+idxkeL1IjlV+gx1U/FZubLgMcg
dJSkvwCUoo4r/4Ftd3gFldlXjm9Yrpw1rAj2NverYNM7JQRmcLZbKJ5hWNq9RXJb
0y2CsnsCBhJBdhLibluzB17pIIiX2nYaCUz1oTEhfAMM5qJozfeyNABJ4GjkBelW
e9UyKcwyc5MK0+4o/7aB1uE59mUVPxn0unPyNCC7wexrH07nGsuNY7kNVU2omvtm
c7zjVLo9Xcwt5ZysgaNXjNUJDLmQFmZB73Nhfld9jCcjbC3u4kzCWmLtHlECqvhf
We4XAsys6W2mAYllrL4X5p+iwnjdQkMnifwwKJ5rW1ejWg83YjrraAsGxxu23R09
Zvdq0Ayf1Scr7gH8DryjIOIReeBXQXEYpYrWqG5FyW1Pd3hNu4jPjBkSDdSbrzs3
WldBvYfuib7BucIG916iK4LTfQfR91Yg/BB3fWzYk8PZixhw9UwVVOhW9y4tm/sC
RxNKJiwD6wJHAHcPRB9UVqzrx+a1Oi2cnF+Z/FPDxGxupxIXIyKIRXECUxjCTBUx
D6kpgxklGH0D+Yuu6IojcgOayfOk9BQ2lBQbqjtV8xB4vHMSJhnXXBJHvaBNzOqA
CoiGLT9c6jwsklNAmt69IeNAo9tWB5M1Nt52jIPLc8wvoNW9JrDaApQs5iqlRBWv
XEWI834iYHd6m3i5UBf3JDDZUURfESATRGdZjT5ii7u/WNw58XuaCzfgRSxOLHpt
rwxqNgtv4UMdXek1Uj7OLzCeQFD6b6D0o3HOB0iIrV2eN04Ri9scL/467lAhiYT1
1GvWoz8KmytsTowl9V83/qpP/61UeAUokgCILoA/8arkAA4DATbXk/BlCZzh5OPx
fpyyx9j520RvbVodVW3GPeWZoITZM+hz69dWBNcGFwlNgmtfHj0Mh/fDL/EXoq0t
h40QanalDWfcsHz/MSltSV7HBAKCzCLrVjyGLqSNoIzH8HuTKwCenaR2DVs6rGtB
bHUEVPnUtDnuNnu3zXJn/KDOe3rR2sYqKd1QbiGxERahnR0nRPnK8/AKqCrnKc6a
+Pir6Zx/fRWXySzpAy9mq63Y86uBLJKSo5KjtLS/bekUX63IgekN2rDoKO2LdPW3
hVi/k2aHrazVQhhUkIwyZZpSG0zRQPtO425w2E3xOpxJiQ1ZmJxY2ws4zGn3n38K
lOV2y5TPYtk6XTPqDvQgbPb8cFwrYQh7+C7nDzp7vLEMPFVIHSBOQUoScNf87miM
8Ukpjo1Gyhc8PRcf9rPG3Cy5bbqVFvXUXDTP6yUr6+e/GwyA83KlJyuBSra7nzUy
pCV49R8j45LtWJq1dYiOkUy2F3AnxNOyVA4YLQzdqnq3qg5/HzPF8DXyybhXzb9z
LYmERTjUhMP4OD4voMIHGBDxD0r6kEcLZSkSKlmA2zo2UerYvWSNi0XyNDo0IOXj
uSuwcBfxwCkQm8cTzDibta54HXmuoZfJBN/ykT9N085lRFEGntSCD+BADjbhXuRp
hSHM3Gfmi3UuNN4lft6GUHbtEcfN1sAqJzaglf8pxQSfwQGNtnDnRA3tNzGuPPOq
ykt/eObN6PhYa0qyuK8AAhUQiiLn+UcOKqbLNii2iE1QHb2AFm/M16P8q48oXO19
1nBnopZYvOSgL084XD1bANWPdozgA7NlpP1qofSmGKH2xz8BAMVuDDjSiQ/5twCa
yQvO/VHNrqPOou9tbcuQDZ7o6Uq8ApbwqTcbJM0/IF8NfE8Y/w5C5NKzFeU0Zcb2
l+jCdumqe2PwDeAi0V8kkyVXgw5N1FJSKrqtsmFQ9uvaRGBlphb/AJ61uHj2eBB2
wfaZ+OGhgfS2uaslhNFs/nb/PaDmi4ez/iBNk4Hb6hCSwAQzAJbAxI6ix8MRVavO
Ge4SCk+uewBMLa11Si+9hsg9PUqZFYLuLBUbnIJkfxQBT2cOLGV6jzHJyz97Haqr
ZwEbrWw4s9iI2tW33CiiOhwML15dr93sI1vinCLEVWtLVZbVvfsdbmNbnRfVh5JR
+5OIzi4RwR8OiQvtDyHchuKTtjBB6P5tuSpz5BuzQCP5oNqWKDLb9bbrb8CyRHIR
EX/BSNHwpPH93ClwjUTyKSLIo09P1odg1O+kLzL9pD0+M5QD+m5yeuOcn0DnDIy5
0vribhHihNRHN2/O8D8Z1k9RK9/kkECx7hxYHfB74mDe3tYF7bWEKvRdim7iA2yD
gwqoshKcRMsbGPmn8WL/Ay7d7+mtsMhHT4UsTGHFL+quqpjSo6QRrO/4kvdPbr1A
mNYmZaHUxalhIuMOIOXXLee2RgeC855aYSQwc1f77gweaK0jiLJiS6WKaWGJS0EI
pIhzOp9BHQXPTon87HVd1lFWpgvYF6iFTONw6MGK5/tp7K89tee9/MNC7dHu5PLW
m6ayUYYpVH9WIZvmlp+6c0k+hzN3gqMv+ASM45LnYK/jDI2bMYYiYCRd8MUOU0ZO
g9URhO/4LJo7eTuccDy557hON7ePd+Y7Sa+3I+uKHHQUfqUVsncwlpOH7uh/XnYY
V4gdAmKX3ldB0x1KeQjBw7ms2LRpjbQBQdDlH+3Bg2MCdb3oDpBCRiOxKIjrlyW0
TYIKj7ibnp9VRbjylJpfi/1C2/foM1BNReGVA0zUdFBRvn4ejwCux58aFfGSBtxE
3tfhTx2KjKu+z6hf4rIkrRtBk2HaJ/dBa5Tic/WDObzkhHiCIHgB2SD6KkBfpzH/
Wp5HsWnSjbvHvOtQvF7oh4Wi+82Unm+xaS4vXHMh2fQGOatKueWH4AKQUq91kT6E
VEWbxR8nF0jZ0C/vE3mb/9AKpHd6TFJjrFs42Z2nkSFtZSgM6Lew+VRc1N+0+/cC
0LTJp5Y8wRdRJjOC0caY3I8l+W9t6alak34XwXXduRZm6gECfP+TszMCjf20qXEp
FCK0fAeK4f9k42TNFtdhRhepJDZxuL7i6K1/NP65SFqCOEQYQFXOAn+Otwn70hHJ
nS315+kE9aMZVQZ8DRokzCknvyGhgDu016W71hGHHzInX0603K6EJ7qsiK14wBEk
wivrkfYWGq2Z1Mx9u2ll5fS40bZvbR+I3lOUHzEDOs8fCsWURjHz5gmw6IIQjEIF
spr5OFSuht8e5f3z1cY8dPvxS04Y+VJR/QYuxZeYlsVzJcbTzF4cC7kYKUjMXmOJ
5ZPwg+tcrewdvKPhnZ3gZkMXWPYl0IltyjP75WoJ+TKW8gUdo99hopVlgSdxx/0v
LCrAufU0Tig0Q3BMxi4C6VmFftbg6M6llL2VsEigIYHEfWn+nnkIQYWG1avHuHJX
VFVuLaEyfcLd0xg14TwnCK7k7cqc07DJlznZwkZmzOVBFmd8fd2mHtK+WxDWxpf+
g5xr8FP5DqVQZ4hTvCTOvXJrFbg6KjrbSlvJoghAhrtx+JEWmLVh8iMwDaFi1S17
7NUSB6tbN3hxK/fy67WkFdmCWqfHcSqBtHbpLeVhfakNxYetYmQvFECnQpsCA0U/
INW5wcgDx/3J46kSTpjuGieOBq/sf6aOeOZa6bNmFCeit8go0GbBtyox9+vlmp87
MH4Gu1xV3e1U71k2p5ltIl1hDd/yDn44mxEL+pvCHVdEaf3+EObd5hMqN3ik27Xy
eyfp2h9I3MkZCwsrni/BKRq60CHsX44uQ6kHtCk1ZZ7Q/a11tv78N65Q92+eAHuT
AKhUbd6q7eG1XDaOXlY7WZK25rpspjOZLUmy6wY8Y0Q0DrQujt0asyRXQvO0l5Px
XcMYyhyG1hX/DljjAoSzxfl9hbJKb8/DKx9qRps88SVSJALHOzp/I7T/4Tv/VB0K
LftsmWUz1aeVVj+9PlmY30CMWLyyAwFFuVqpM9eXTaTT/XIIXSNMdq7OVdd+FD3M
AhLC2duA8gXUnZLBWKQ/0fFGorYfxhghC1TQidiifL04Eem6hwjMo4BY6WMP3FQQ
u669CSV3jx1dDTVMZDF4qIvMu8yVGfHZaT57rDLKoblnGjU58zEuhUgOFJrVsp/L
USqdFUINyQmF/kmkyEC0Iv13M4OFA6w8899kqgnvK9ggB9rbJBBgIocjZT48gAub
adYZwDHc4/nyMHd5FGMgEu++A9seGqvr5RiQ77OwqaD8cbeGTXMzzZVAnnmdtP2b
OcZIZ9hy+oVFv2TIW3rKw9GyT+ZF72Y0IXUkbJ+obD0Q43SfRUgQaVaxIpRgxsIX
RoqIZqCXp0cFZ5YnBFhoqQrfPSHfttZ1xynWoiD6y7SSJjrfD2YBSkr52HZ0KxA+
T9HERLlEtBeXZ2e11wLQORnO5aKtff+DlRblSEeYeexaX8aQaWokE7/tgzYqbShu
wq7UfBjuhbKtI5zGJt9tAuDfAcORzjUxHS86NFW0Ws7IrmxhCXc/teAzpX6Tpyyj
oIxJcD6OhqxxGXuwIKzlUu2ovXNIxugeU26C5OGD2/TrNoYFO4275RI7XaQyNR4R
eYV9OCSN/+Kr+0S5HhLiF2gyZZMLTkvYlveFTFOETLbnLQzUeqNaM0bMWhxRhCpp
6YFZEttm3GqAnlL5c/x2IYvD+lnWl4pDGSJpX/mgSoJfyfBgzJZUfY6peLqLagnR
JeIWD9Bek5V1OHLByat8231P+BwyVZhve3S/XCOPTi3j6jE477yQycZpJw3O/Jjj
0lDhuUlXThUuQ9/Mq2gdoY5i8nUlfgSN9/T2OeOsM7LmfG0AypWfjjV+z3vnjAIs
BH4HzIjHXuooGyAvT4p5jtnG2E+XCk1tc0wVMT3ftj1z3EFNAjupdum5K0ekuNLp
woIQuBdKw2ffsdlVA9HRoftOr6pkPKhgvz9KhDFox5cw+lbhKhRrI+fTmV7HmsqS
PRsvvqeq9SZeiGSwwuLh5+uKIUY3Z7cr8tZQq/UQwH8u91fJDbI2WrgxXsgzFKZ9
cdppaCCxFUCPG9M9L18zwf7DZYEi7aIp7TLmq1So0oDNG584Oaz/NomAVPTldQe+
Ox7w7W0WfwcKXe04JzMkqtr3MAbrVMWObRf0WuoQoZKmahwKYJBf7txezuKDRYpr
ekARWHdt5wu/AFB6APZeIlKvwhbdW9KRIUHL0GW0IkDDLbKfenXqr9QCQZ6NeL9e
HFGVauNWqxk7ulBhBPgBTOO3dme6BohHjD597YQKL0AfnKHIJ6ETlbHHoquV8YZg
9nXpKx4M7pY0ijPy9H7OI3u8Yo92cMq1AbAHU4+tx9/q5/n+5L3I6GixExxf0/2S
kRhHfuvE2mbHmdY78kRVcFOu3Ttq57TP5o8Yyv1LMN2meNnOa6f9xCdjudrPrsqM
+ZrHXwc8V0XcVSnkFD5fNxGqfUy7fc/QHD3bqPkDXyalJS83o5E/+mWtdYHFz/Gb
qImPBBhUUGfEUjZNEBKshVjN79DVdoOBdpXiueRkfOKoKD4KTO1Cc2dFDM+N+xG/
F0vR6nHP44D0eBfymVquu7pWj604+q80+i2wgYnXzsgmZ2B4NSzaqZh2dtTyhp7J
aa+kg8f//L7yhZIdg5dG2biOrHRRN3e+Ii9AMfslbOwC9zNPUSKsPdKJBaNmgP6S
ERKejwEod+SH+Ux835CCN7ORQTkzrVXzqDrc0LcJ5zymXEsgeqyUY/xk4OPLpWGb
oTp+SOumBG3b5jIdwPpuuo73uk8Eu+03t9khh5F3tra6tjOAoqBcma3Ck6LI9kDY
dMcdPAhWXb/e2db2+rkQYteE/lqZ53vjMp11F7jJ08xfPQIS71crGh4wbHTkZZI/
10yvHv/azeX4i4aZ4tRz2I5y/xYDIhSkctk+quCVymwY/AnuSweluNMQarBR6CxE
liOh+ki0ymb96ukG6Ju4Xo8Y1fQJKKnnUfyRTXVTMlyKfEWiMUI/bclt58va2Emx
B1PeFUr/kPV/Wr4rDrsC4WH5x+W8so9TN1KudvTyk2+m2fq2t4fAWl0gNcIJPmP0
rhRTc91i5+Xp7uSsgxLTR3VIXJS5CdcQQrsAEKcUJW6/6xfGMyd3hS/14F5e8i9I
MCDVH/+rc/VR3tQKWbqDQ38g0aQBKxInym1oVWqOicT4Y1hnhJwlzzrwubUeqrgz
bOt8ca9Clwe+LC8irtMGCKY5N65XfdHOsMSb7715K3QX+EJKLtbhfnaB0i/atiMk
amsuNFgzAdIjcGQdH7mDHFter//0168PCwJ1KKRWJbVaX1MjJwncfwe0vPTABYMA
2bACWo3A83LzBJfg2Dng1bB3vx9Lvhe3jZFPQZfjhnMoAcoC9ikn+nX6lRdIB5pj
5rpdFnAnLNhcKY2LPXqxIfUmPKXpEa57Ta4PVZ46j5IrCBvETSKo1b9yNJTPfRNC
3cwXFbVOr28KgTJQr5jtIuxGMPOGC0mopsv6HYrbgsWEsHfKdT1XU0ST5DqqpcOf
LTBuX5VvgW7vY/Veu2P/efpcP+5I6cLN5Y3QBGT3kd9UZxeieEjZX1wN/r4zWW0D
f1Ot/VLaVwncrdusJ/utwyOYeTipmOAL/ayKDiNHG/CN7d6FS3vxcMLVcWUuiib6
vEkqQmgJ4CJpbuoiyubZCKxHeTN1BqO7iz3RZP53RcKozZt7eg6fMJzAbcy6IlXb
miP5Y0mazVpDvOK3U7ux7dTPFjO5sD+sPQpSy8ph8jWtwNx0FiFayvGcXYlTgbsW
+rO2UewTjgxkfQGv1qxJOO8nLZXPltQyti7bT2wfcJzI7x6l3bi+HUXxGhzk85H1
wQPMch1dT/g+lYTCGs2J9kZ85Xi2+oDinoVZLUWHZ0VX51sru6Z1vKkyMJ3Y9iXR
B14jfN3vtBCexguJ4cyEGwd0qC8o1Lgoe7NsfjBj8f3MsLvWAsjDtXEgBOmGvlnk
UtfrGdu1iA6PJxHwX/zDDg75G5yFS7eEFcG3Y0rJxkcEAg/CSGStTp22VG0IEQ2O
ssxcTNSisU1LQXE3qty8XyCwIGftF/YFAnwqb8e46TnTx+Ej7AHQuf0j5SQP9Fqk
gNmRYXlyu5B/15T/UP1yPKkzHxQC2y2CQHqsC1DSLR0k4h2Ek7mjO4Gt5/c1z+Vt
FTMsQ4lLg0vkdR3AAQ3dFCusDNUO0GE+YRpyH3LMGeFQqfyv057SJu+W47gULn0T
UrOxNrfrgvAXxAAMkDRvtNzDHM3g32bpKUwOPWPJ4tIwNrjjOOJoVzbRUIXOl0vl
05JmkMHW7krmpTetjADSdA58hBwtgo9jbmrOvHKHvyk5PvdL6qr/qe0dJyh6TQ/E
ChkkfrjfsBMzYPmzh8En/5C7PgQdbn08UabGtq17Ct6qMoExVAIvHlcEOtqaGjK7
UoSG7/EXhAgo0asx4g94FnaEs1WIm9duMDraMREBXyHnhp6pRCw6wAzWNigmMU4G
8EZ7dBi8XqX8DlLxrrhJeR0TrwfnMiBNWPr1okV8FT3IGNOYEaPshF2Fq5ATM4wh
+5GzJnz6lGtaiEcdLCepbiKFET09g3VDXkx24DoUF5rG06hIKQaU0HQ/WAEzR+oC
Z3/7YpfVFT7tihJQRqv2stYHRDoVbLNdQ8cRZCFbQHVCKI1TBZQGdBDGbvLilcRj
UltME9gx6siY25d7id536R65UaEz2MP44ffB5pGvpMcCI5gE3NKzkFU+gDCjWpu8
ct+KT/pAeEnR/nDWL0FEuaFpyB3ncTAJAfNEW3pOZk5bg6cPqv22geWr4V2SHWuX
coSu0lWJqy+rRx+ooD10RzAvcVvIJj5LTJXZ5xEfNmOUpX3hHwH6jCkbknC4Z1w0
PWUIoNKgsZF2DCXrwT1KYEcs0ivmdlloy5rrfkXfBZ/MW4IIJRZHhhu+pf3/+O78
5rZfZmHUfgmKPCPabJrxhW7+1QQDsqIvGsmzfdGeYwLXTyDrKI2x2BdWhJYlQPi/
WcOhFV9DB/JNCTMJP0FLX2xzf8Mcap5MVDo3gQzVGxjXC1ZdNEet4uhqx5c9ymHV
w4lktkeZM4EHR2udtAXarxItz0OHsdfIF4j++n8X7b+et3RUQjB5xDl7aWqBlo8n
FqYe2/JfZVAgLonFGRu+hO6DMV+7ZHKeJNUzle/+Pk695jEh1IKVXcwbdl35SneU
1ei/OC2ZEQlJdKaMbNQqtCj1dc8uh534njMRj2p6+o4yFh01G3EJ+6Hf3FmOIJDl
PxlZdePSvABXm6GlPXqUWjv2B3pLBExIbjpBje/E7BMpw6Ozjka35lD5lex5AsK+
vuosVpf9LlrZFltzeBG6n1O1AKMHOLw981s2A3f+bgLqH1jn+cj8fIUQidUqd1iE
SQoWlWR0hov9XeSW9XIulLtUolY6aA7PQtkCtWvsTfHpinbwGjwqLbpzy8YS1PzW
HyU0UCvw6a8uHytFbeuXP3aK0xyZwBYpc4tCa/G2scfJ+odBew2a+XctzbiAOoFm
5MFXhNkWoj2E1a9+mF5+P35JpO1lSBnJVq74V/9DMCZ825nQUgbdy5jD54o9MflC
kFMYvvE2pWiaf4Q3Z33YMNRMIJ9zCgOrc5at3vFZoSNuYoxwyBQluh+StbJWK4tB
owEm+4TJQy8pFd9RurTVwqQ8sGkWGeEuf3Es8p5k74Kj1XjKK88EP1hAGVXBKl9n
YHjPd7LHasbFS/wwfD/qGCC0Ts/xh017BArt4+B6RRni0wA4IcitH4A5xK1mTHiv
5zNh2hRbGDd6r8lPQ+e5lkCZ8f6kSvX0NOt433LzE3gVPN9OycKBYpqPxdHPRFa4
xbN9ayTNZfbWqvwXjjmPaViDdBWNlRFuuQxf6OGXWieBrt36T4Z1K/URfA6DeVOz
pPppUgr5mr+loBJ1Pj6cAjqfQ4BTUwx05gBZypMHRVgkXbA+48AlZn3Bs33+guE4
6PKx3hwrxuaqlB2fQHSGPQbkLf8J6qCKbrissJ3Ao4tjlIhmL3JV2KC0xQRqrzYK
tHcAuo9GXlblGBh9dhQWInwEkDLr25Nzc7D6yxK6pUnzBiTyv0iXOLrhdXK0rrVR
n88SlKVPvI6KXMVARsVDpgk1sB97trcaZOV/0dZvRqRX1jXvixkPtHDGlcEyPQlS
Y34nhw/2z9adReHC48sSf+Ll/8EeGx2dasobndOlNnrCQF9U3t6wtAI5TdL0NprH
lJNMKUzW4+RVgitQvIooGPtrYER71+ICdcSdholOpTOGwIQx8f9ecDllpf4D0Ed1
rTPeJWFYyp3g4nmIOFJXaiiBAkhg9Crf4gDNPZrW8Kv5IRNGsvR/pqADrDSkdq3G
lEifEMdD+gWoxHWY5Qy7I7oiRR8o8RneQD2COwDoxiIWIHqoML18tQkPxEHg6kX+
EVxIPtL6usrz4dR4D9haC4sz8p9+IhKkF7ND6Dc/n6xX2FqLlM8W9LEkpmfsWB49
11OpKgjVPoD6wO1M4Ac5rO1j7mk5GymG1jvjXxqzzPoO246nj8vz6zVPJaFhi9xS
qWPWZSjtkPI/k/mq1LJb6uXJOUZhT1wGxWJQ+jjcAltGNrRemrJ0oW/Xz3DngxqH
GPtj82iamt+p7aXSPyZ0d9WQ8k9QsGuf45D527THQkHWavWuasqbFUykoyNQve+U
9YGPsJwsfLusx+i1SUJrCETyivzwd4MdqDfIRuv83touK3ZaAsw1xUudUpehtPRv
nPI0n+MO73j8uC/9CdglzCEWNENNLZd5suOEjaDFLCWNXI98eCaJKk09c09uXAO3
cfMqWLm+qn11KLX3HOtreBkfd4A67JtHbM/Y6R/J/WrHym87sEWML2ZJKPWbfQld
WvEUD9818v7OzL8kIen19hTjfN+nZWRZJh8pLuZ8Ph8IhOtnbqOcLbvaVu/DOeUH
l4yEsg+rAldAiJA39Up55JWNGcpdGSHY1tHZhi3oPe1SeoG7FubFfbHdbXDE/x1e
63n/g0dEhH1Dken2xApd6wZOFVfwf+/ks1o388S3dt2Q71g7dbth2FdHzfz3JjmU
40STuCbAN2sgvs06x6W5xdkuNy/kos7yZntp12o0AU0iZ68jWeJK8jMNvR4vB/NS
lmSzftspVJezcEmaxBbgUF94KTfZgv26pO98+WYjMN/kuzH4iL5ZKNge1Vlf61lf
cnAgGHUI3gplkta+XMVqa1F94k8PqtabcRD+J6eb8CinHtU/6YHXw+UACMD0NdBI
EnepIAl7/RUpb3xveHqukB9Yugt06k3RivqsrCy2XZU7dA2sNwIH4SgeLC5YLMOR
PO0Ji1n0CZRXWyiwzyE+YPK2X3ZIGiy6xbaGqeOwEvF0mRmtqHVNrGqNUG3l4Wlr
2qhZ6SWCF7TxOdBsXjPzSJhMTaRe+kuQlrPZ62X7l/oOYNhsUiYcmCE3M0SzShMG
huy+/77A82VKR0BXnFVCVXLGnpCcaS5kHyaxZbkCMHSErMT6LICsM8DIzaLEkyT7
ghY0nKIlzsOXI3fwDlTScRbkzGpabfb4ZoC1txgyIS8+6esSoMD1fOYZ0PcD1AjX
delameik75Is03EhzeRqbR/tLD4kqCF+JPTzTLIfuE2hMIQMJsZWpLwrcWIiLIvD
yMkM5dcw+TvbxuSb2fvJSyTSJN6auDRg5do59bNjWXwpnl3+OUk3tggBUs7xySDt
3fkgquAOBUPl3wpI0a4MrJSo15XGQRv4xc6DuGoqHn6GZW+zKMolaLsUaYNMdSgu
sovvemXVVJP5nvbTSZXvWRs8z1TmnwQeXnxC4UR4inmoSP44ctzxK+S9yUGeyZGY
dL0QON1axbfNTnRqTdMRzXxT1t1fttZCKzhK/VAbe05IkeNLAYGKRXruDLTl8ZEM
meIpxwvl+c+YLVdy2JTDmPHmylRL2ecm8exy35Z3d/k2YRThLclZynRY1T2jGPNV
pmsBFJlSM5vRquRHygsN5ct5gl/k8njy0Nu1pIDHzfQraZ6h/US0URx7+dpUu5r6
FIQBL8DcR5bHgSKiCu7zPTLXDJT5Ajgq/zQPRfGaCaJh7Mn64pQk7q/aUggZXIyR
Pwd5NQ25FYKsKtM7nBeWE8aNTKVuPdgzb6gUcQDU9NOt4uq7eGQdFLXo8zy0E5Rq
KSw3aTHPJTtAIJITuoE/FMfNfD5F56ZTonprUfBaoBAczPihuw1O8gOKpulVVTmu
tIngPj6we1GMuj/qJi+fVse207L3Vg1o4TeSLh4jkVM6W13cNltKqZMGVQ2Gbv3t
eh+w2PCS2QULtvTUPK8T/zYyqs8T6LyMMkv1fF80PJwtKXWXpUCFavk2phqL6o+W
Xo31lQS+B6pd7CkXRaEJ6kFdBHh8G5/OmwrhGSlTpqqCrbQiu8K+7LL+Z8W8rBlx
GqnwqRRrBPoR+PSZMldZno8Hr5wRFXzIcVn+lXbASc64d6QPv0YxzD1GUDLYSw89
uafHB8aMd4MODh8V4DIYd4eHYcwUouHPZ5ZPQ82KmpueyV8dmwwb4Iwrt4PxabJl
ZMqgkNyAxuDFCs/clOzlE8rRff1xOeg40EYr3Tfn9vhp52iKeaYln5g4haxPXUOb
QpsbUXyWOT461bpKgmQ/Ba06fGoYY8AjZAMvCKjo6eYQCRU4CKng9PackhN/qcgS
at+O0O1MP21k2L2KkcLf8WArRDzxIwwipTJRzQJ0mUnxcynRrrLrRdEtskQCroZV
6EExleBV4kb0Kj98Vu3FlBTfGx12ASnxTWvxuw4mN5hom3tN+bU1eKBOEymtGk1J
VoG4gqPgeaQbL8A9CSVWSlxfn0i2FjBKbxkPaaxYqEJ2hnyK2LiMLTHH6lOB5SHL
90EOwvNSoqhsqZCEVq4DhGMqbP/Dtxx2JCJsXxJqk+/hVH2POkwhzWkMPWNMXDt3
JHixfnABpBBSqVcPvb9DhAI4eKqQzg1ZZDS6zNOOofMvc9kUB9mTCINLy06bfd1h
xjlQ2JCtmisj1um1nMcC+eA427nCZoTEgNb/b6B1QD7L0yTsjZt5yWbKn5EgqKaZ
o6uCMvZJ9kcXruDDzt56+vRQU145RCM/slgkvmK1TdmqrLWfuUoTBy0jBPTwLnoU
iocyoh28CE4LzcUOhymCYiDEiTqAFiNVw3/RVPLdcHikbLb+fAkWpGrkG8E8Ojd/
kKN/3H1Nf9H+kPtGmkizhkWy50oVG+P5UDoTuttXVACWyU6a4G0lH64o6R9hncBb
/v68Eo2TUC/2yhJNX5S2aaI4Ku1L3wORNOrFZc3McJHduLfe2SJT0w7M1Tuil65g
aZg/tgGnycexyWAF5phbhSvrzFqysZczrz5omw5z3OYuKOaSLRVgHoE+DVFDpeQn
kEDHAOE2rHulh6beL12g/gAO2lGl4H+lpblXSar1qJ+sTsQm2Qi96NQCNOh18P7f
BD7wgDV5yxjruDa4oKAkZVKEypdJWeFcqagj6bNC/zVPUUaO5G0+pNV71T6x+7ta
Mjo1d86BWvR1RvDRlkpgU7KlGvmJLCQDjZLXiugCo/pV9AgE58A4+AQZTIKrxRtw
kKYRFtn8Bo3I0k+DF5WW3YntOjMBMd4eNDSgDHI2GAQMb1gHVItdbqqFKd1ydHBd
YdZHEcSHiNIKITdFN7uMgUqZ4ORIV7S3QTdN861g/PAF0HYwHpWUBRkGWMLFib1i
1hs3fNGaBEUoVmYDCsMeyxoCVS+dU45dmjG6Hnl2R7sb25Ot0Ce66zDaEHT2yJsE
NL11V/uYKFdKVemt5gI5GPf9oPFpDL9Ax5xG50GKbVnHZ/cNq1+Jq3mJBhuCWa/F
WnCBnSZ+Pt1M9zJ+D39UlFdkz2lEB82MLGwcfXcTsBGijmHwDlphXLnsOT5qajSf
THRwwnXdXM8mhU+zK4pDZFSxTQsWKhXaM52WwOloco8315+r14NvF8yh0hG3T8a9
CKhOfZNn5XR/a+ioz/on7ET/4vwzDBYFhf+Fhqxpmbte5h0qj/GVPioGB5vsirTj
3yVdrb4kV+zLSNpAudQ8nlqnPWaSkLW3a+7u+XlgsNNKn9vc2wauzKP2cUrI+3Ez
9DuNITSO57Njtuzl6fmSQ2NYsO44gSUFif7dwIGgYh7nVatYbF9CGvYc74+v07gJ
VIXw2ghlquRcOkCx19XQWUGg2mEOBHtoy4l1m1KYJnlk2fRnaS6MS/tZMCONroiL
k1XDoPsspB26/xGECprIyTHoMV2ZM7HLrZ9hoLkh2NCSqQYxgmx+3I3DeSpI00ad
Lj7QvGeWYgWRIdnX/9T1g68zuDsCivRkiq3QV9JoIeoe/Uft0Z2Q0gspIsMMsLG0
jJfFuN9uschm/d6D1Cs8PdKylKlK2qfJVz5lnWLEgPu93HirqSvu+feVAedHO3DM
Tq9nSZwDbYsyhoiklvHx36gm9G4YsLj1vCg/pfYudDMfE6O5ssLLHhbHH4dhZoy6
ZP0U60lkDEhTWOOjWGOhVzoBNfaCE8d0Ho0RmIkE5630YhiToWKCGD6l0hPDCSj8
bvmV3IdUH0FeZMUgqw7LcL4Hu9JqU8GQBsbY0ei4Y1U/CELGpfsKC9UPWiiSABck
gsFVZX0ZtL9pmvpFH6Aho9mgdJSqPk3rurlwa4BLqiB5+rqYZ4FWUjVV2b5vU1AN
SdCFUdbppjeW/3tsvXMHcCNaf0hogD5df2PPbJ8LX2HW4prgmXZPBvsZ1C9JqyNJ
qWfJNet20MxwTgRD8yaFAhhKXtRqpv+UImQynoIjFHZsYQUJzlHavnLtohSK1Hg9
H1iDV2Ba1woSpc6x6DZmWXA9zwA1f8HI67UT56ttr20/iJfmDQT7lLZfSkSd0NM/
lby9HYT1scgJAmrxCLeFf2CjxqkQPErIAcLQ5sTpN+55/2qwaOD+pd9P5Rw2phc7
3twrLtk/Ts6XG6q/qFjKQ81os5/uZWR3uXGg8IVfyvCw2LRLpyAqfp7XS91V0nEw
8z4rEfp6UZp0SV5sQ+Vkq0UukpKA9t40I0AbCJqNbzn5MvsNfzzdKgCi7GoQluTd
OXX/NgOtk8x7vN6FnFiNkUX8OH+gIQl0itSKUB4L2JWCfgs5hNc66nKCLeMZKMgG
j9w9QAH5/6KMHGGboZCK+vSUTVdwIWT/vZK7caC3sJEaHpskPtXIs3W/Vs35Mlb0
XzyVlNrCGVTArrLvrK5Bi2/rKJe7eCy8EDWyvK8AeIEcX1CAK4RL2lqhpGbo9SLF
bvwJGF/RaN1awUqS5IRX7ec+vQa6x3RMqqhapg7tpU0iBBwRsF7OVJ28B6Pj5vgC
j8woTqDp6lLT2W3B9Q/e44v1LQAXxHb2CBI5sftW7JqFK39SA+elCWfZoyvIRmyz
gO2Hwqqv3vIpUdshTxAIHq0ZoRnRD9aodTnstuIZkK8CIt8w1CUk5X2s3Nf31PSj
136mj4Iu+oqhIVsPWjjb7fYtrVQnQ9VIzc8mxon4QoUn2bwEo1TMt2vAh4KC9dsn
7SmNsO0WSeWa5vc526Lh4XRJ1QFjU9kHsQh7C50HQAq97BoxqOp6zq15bhhHFPYA
QT2lPosQ+chbaMSfR+VmVgoyxNOLQV3tAWt0S56ojXdIJDj2Fyui51NwOfZTOAjQ
e2QfjqMPzQjkFCea8xGKlT7nPfaRfpm5lh59C6gzq0AME1YaV7rbkQZ99HX8IstJ
Cso/+fbAdsKdqugBXqAv1BPFPeRAF2SGeDVCjpy+1nqadURSl9sEsPrSwiQTUAT9
cI+LXr2NRKZebWeupLksl5JyRTxxu66vwGHF15cbxHVwbBvqATbPOBlycl8H7f6K
jZYfG1XjbMLimG7pGyrAw0EZLddxla4kZDNpI/nkzvFlZxKjiislNkZ3APcyW/zU
/T980qAeEGbBxf3jWe/5l77cQ/Gf64pzUqiIMt3xCWGtYB9J9vUKCNxqpEUZqlkW
L5Ng7jx6Vlx/sntx5noAEvMu1YhYqcX3AS4P0gJ/7kzc1A07zjX9867lMRfBrbwm
hTXl08ckuXkdoA6IrlNBTFiCADhPzPO5ZzDG9ntMYuDuJdSbCpEoxf1wL5y5U1lv
rSZjdJdDuuoYgZlN7aTkh9X/dC9T9+n8IJK3DaMbKoGW86PffF3/9VZpw4YJ4lzs
WPGclJdtmlsZkdirU0C00nYcNclbeSUYOwqjI+GAabGsyrX3kS7XIbVZPxZLWqrM
tiL9ngHjeZoXScwZsBe49E2t0eIbxDqFMvcpztY9U8pDxu10ifJiJh6F6qR9649i
qmTyxfMjLz1RDvM5cCUy3pT42hTuE8IYdrwwgIHIiylAZKGcNMM9LdCO/tpgRXaf
weNOdky4brjd2jdGm/Rlu/o7CrD5XsmNg6s19BnF9m20l0ozrzqZjg/3RztvZzEe
YSrwprbIv3Jsofm5tDBMa/siEszRn2wN3gYRRGdi/gg7wfJGnuHPObfBQufYrpc0
X+zXmO+DzcvUkOTJtThzU/p3DL730ADtXlIpbbW5KbMc4hKn/3UsHPkRQJNcssQ9
HeS7ziYJ4HsciTZW0O40xquK1uOu49wJDrMKNtEVpnloa2gvyBMZ49URTl03N/qO
qEmkbUbyU2/Bo4iNyhDtHuAF1C3HnJIjaLxJ0mSYT2ivnscjY5xlFar1bSrcNM1v
ikYJSQ7zI85eIUcdOKkCA9JQevbKAXySPV1spB/hSf6tcjIMOp8jclvDGu6acgNR
lhFCAQvgAF44WKAVOnvKpIS7V6s0YOnl6hpGnotqJabp76ISQbjtGqUYWIjawswx
9Zm14GLg7sJP57oZxDa7xzAnp5Y7F8WcXtojp8dH60wtSY51JWbRgLyKea2gshFC
trnU5YbwbrzWM4e0K6LT3936MY80DUNSwPNrQSWaMi8sBQhz2si/nrwWU96b1v3+
47szP8hvDv8uzAOoqNdM05bG/VOJhUgIBxKvBdhcFNxkCnIG5NNkz6rC28aVjkKb
smWA5WdxzWpI/zh/+4TVRSt6KOx28nuT33JRHEzMTjwQcookF4iML0b5g0bK0nAS
pI6iyIrQjXsDI3z57exwjIO5dKpnt22iw2N44LCGY25+ww697Fo1RIQ0XrO+ZMmo
U1bgDKID95yt9bAwrQNnhup+MNAFsbEtdWtzPXJhYADkDMjnB5JsX3PuMIFK9CM/
+YsmFx8yo3+CcOOC52W/MonVr0wX4UvwtE12JOKdTg2unNp94chS4tlvvQuPWVr5
9M4sPSMC+nNiinr6BY4f4o8UXcIksnPKzMhIceKQlLUSPJIRc3GXh1L90LSzdkYV
fH84J8HdYjae9CiElOQ9Lkf3kS+h8GfE0gnQlNWCi/nCqjWQOV4v0WBXgOfxGdCs
74ezuYnxmX3e5i0b4LmocvMiGKWqPqb4jga/fFDVMppbfiaKM17bcxxzA0YioYdd
ty/LgjUEQm/AxSgwBwKWS21tRyU5DAYuwsddvfF0FJKV9r85+CUcoyfF7burLSSO
b7vqdYf779F4OTcFKYXL5bpP02+UUI4j2+uBqp+DMbY5TuuVnXCq/5TjqJflkOR6
2R1TLXeuwTf1A1Ig2FFIt9OY8aHhD1DVpZmdaJoWE+QghgjTkvhky9YuPlkW39Qv
KvEATwCrmn/DJNH/L7+JLTsHiIDEbE5oGu2eQq0QH3aIUTKUObJZjjLTYm+wgA5c
ScCjnVh0tcd8wz8aczcgkRngCGv8O8jXst0dWR8CNLMO9Av6q/VkMxFhGC/0ki4d
vFqI+ORheUoFzlCIjynCb1WyhG2Y3orJyskM6+V+mrT0vl17xE0l67qwmQG8mYma
6UQngY6gnf1g6jVO6yV4Vrr1f9+veYdzybrhs7MLkjAysvGf3F4o0v/YVy5sXRu2
P+58vBfIvfcSvIMnejaJMK55D8WKQOO242/7SRWmZ5FKLM7jkOPs9cdyZ8HjC5dX
vc+iCalOUVgyRhHwDHBxcpyDCb22iW7Os+mwfMO8Ty+RCAmYXCFZuZyZK4iCngRR
FLjtuAl7LmiD9bQf5s5wLIS9KBNflDQYTOPEACr4aTgjAWl4mYOlkCUacfD+LtTy
+00zNe9mVAoDa6XEPEDWDxFhSaS1gt3DpyhfGXsMqJrNCSqIChxyCWNfGNQbBTJF
v93Dd+0v3S8m3UbLACODGRsvSqmWB5Iahh15BNf1AVEb3/4OjjnqgUVIYJZeO5pr
Sxk1xERJA7DH7i+Nf9R/TRKpAUdVIGM+zQkW7S+pAN5URYjSWrPdpwY041mGqswI
GGlGb3VQ3aIWAX0Xb+XGisJJ0gdZadqBRX+4uQ4VLicbpfsVCouOKhezIL0239ZQ
qTaCdziWm2YH1A8ZWi7TN56j1Ion/mn6hlzKpk6qnxD/uOupVg/ySxK2YiboA3pr
UPECyyBf52o8K1ATNfSDzYLQfqJ+4wzGEHKERYJ4CdomeerzGJaxFDLcp/42ERgj
JfUStQ8TcnV1Sy1pJYmaXaTEKscOZZoQwgq2vNyzRoAzAPGu7UPr4b4VYynyWtge
xM2CdVjGrvv0k5mqNPmHiUKRdnnlmRqUKtFt/hw5acR/EaRpqn/Og5BE/177d917
nsAKj5TMqGPRnI+gf12k+Ge/0SfB9QpcstUxGwaw5fTizn0PRyOsHF84GLwrmpvS
ioeTb+yPxkCfWwMNsZ1iO2++0RLLfFrm+DTyLpByC0nPomoh056I+h7lb1c3/zMD
TDjZn2/homIVkqXVBlhPvumYY38O1ukOlOcrI9YFWW7+23Jbmf6L/NW0BxsFLqFW
KtUmj+rtiPkqWrkvKR0i1+hz59sjXcZnQPnV+YkFhQ3ol0OvpAzZw/1BP8JZcJIM
QwvwA/mYpuUdQMMnpKjzEK5K8VlhY47aJffq4rMHIvEecuqZQtSf++N8IUob8ds7
9E1Ln4VFi2yjxfQ+Rn+leiNkZns8ylOp82cgGRWS91FwP/nqeHgTQU0BA74XlpnL
A8bobiccyJYqgJEmPnlnBsKYMvaY3UfXJqM6Sw/GBsDjHVKDeLC7DUG9yERuTvo7
1MBLka2O7Do1dXeszmp1+pv2N3UF6IPagSdwcSNpwHVMJkM9+NWhZZkToOwBAaKH
YXsm+H+UKJfQinkGuuaz1P5Y1B7ExXQROFknVKRLPum92DhUTOBpm8NFzvhUbMyy
oeL7pFYwwSDqo+5gxl16vACwZg+2iP7gWjXHJF8pV87iHX65RByCqiHyqt1jktbL
mSHWXs/lFpXIaZ2C3CbjLLIkdiecgK6oE7ocXtfGb5fPGjhShHIIUW2WbibRe0AI
vllGbN8UBtjI22sP+azVNGZBdtFdPRk0nLzpAtqP+AaerK6SIPMk3sLkUKS00DjJ
rPFohveqMv/sIK4kXeIlhwRQYUU6L3LxIovUYjPhEPjE8eouz/ktCO4lf5CkA4pw
AZobr2m33AbbO2CAhqVAKbwFmo55umWLThtHlCAJWmZqYPbL2m9/7A9MhLOUL3uv
+7qv6LSu+tPdfwqE78Aa+mefuWqVlcHD9Aegf5154UktcgIseQrhOd5xmRAv5TIy
SNJ/Qjpennf190Jx97ksq4x/Xx61c4kwsHDK1MKueBAvBZJM6dxU/33t2GlfjO1Q
09nIQujof5S7kArl8l1gxCmhy3CYOIhHuFtiMATnu0ujB0XUUr/VAuvDeaYjmRj1
yLk3x/HufWRUIqXQeaKwTjZ9HyZpFszuVbmAcwAtw0+h9bPVOnlwhxiPd4AxTsp8
0oN6OpnmcVbCQLK61zFjXD8c5hGef7JMzk0LQO54fG+FMgiWA1xudKvsia/UJgsa
YiPlIsBcykQitSBHYnEkM7i2NCyP7V2mBBYXF6B4ghy/3EmxDKUXNmnE6c2ejuM7
yhXvBUj68RFdZ8A+PsVUl+vg0MZilero5iG0+4Q86fGyVT1powbvFVkG1WP25bFr
B9qLCRbVNll/X+8r6WRXfWPJCORbxuePjbt0/VPyqcuGp8GYR29CCMNm8A2bbQCS
2U64wXAXFSpijfruoApcHf5staCp0f29x9l2zA2JM06MWfBe+9A8R6YlBN09ZC02
MzVWBrbdS6ZvuRbDRidQCDNQqHcrTvPSI//tujdwtu0on0u/ATLVRiZ4sAvOwVup
Vi2tuiAbwoXh3yf0dtE7++VmRx18josC44lj565jFh7UT3izihVyeJynS/kA/vZi
RWIo+7/JwtFV0+fZ7cHnjB93iscxJIHaq/27CmEw48GO79J06WSTQAACjv032mA7
dh/AzQwFDFa/0EedFCvBU0Kmxtazx5f9ZxY/zWn6peI5s2KSSxl29U+CaL0hTutz
KXCLYZjSVxY/FPFfHCcYi4nbnSoRdrolnyl8tw99WVZu/ud8PrS0FyGNerW/8eve
gu8VLAdXtgrjn2QkmPI9msxuik622OxDHTb91z6j1agwtyPn59yFram2HN34VfJr
LeFXesdzVb8RalTu0GMj+VTz03yReaGZQQ7LrCHPQ/rE18/US8lin8EVvPNKBkZf
wPHSM8DLDwfqeS5fHQJg3sOg8j/fhrDsZRskjzS1wXw/nJ3ukfooxLhxXAwaD+6s
8kKn1L0VvAaZQCtu8/vDD1aSGeQo0ZE/EQDhCblZ4BQ7gpAeC1RldCL07QoFWjsM
kuy6YnWrRP5NNDYWV9fVcM4V7L194WO6tVNsXBufZAtaIVgJ0Yag2lYoKF/Ct0AC
3Zm8OMOObkLqktVyxCkLFkRgZwf4Ojo42p8bs2Xjw70s8YiQwFNQRUwDUT8pdWGA
CNQYaEjDxc/SktHq1V5/wBn33F4DEvXZxWgftlOVOKjf9QSqMV323IR9pUVq4ywR
ouBJPrbiUAm4ktc//OMfs0AM75hrOcPNi2ZphxJX1EA3jnlSqspBU199akghQJWS
ygZ8xfvTvwPmN9qJsC33Kmm978bJOZcJa2U9ya+FTQygAp0xUGaHHbKVbewk+uu6
+1srBYmjhX3lommEkKLrTdoIPkmGSGgEWLjTd61x2GLmz1F8dTqbtX1MtMf7B/ty
CFJ/R1EPazLawB40KBv9ACYPYT1Oq/X23UPdb2uQmGwleqCBbnGQLiSz5d6FjPoo
4t3dIqxYpLYvWjlfRhKEiV0Z+JDnDF5uOAZT6h6uLgsDsOs1QNda5rv+x//KGBe+
2ur9uRl7vQJK/4aoRyIeWUlhXlT8XtK4RtIMwazQra5UsmMvYqMVnbB1QOhOP8bA
F2BF+uH0WTuncLQTGmOnpMjqj3wj/sh1Y/S4R94dDwR5Kt0uXRFoue/JAKG9Y5ID
MGUmlNX0h5pwkt4y02/ASlfxNT5GiuLQHohp78SaReX4KgFxiIVOa3+xFgRQUlUR
lq6pe+NvWcZRqNfWfom1pYl8EayTDacV+MpEDXyKN1qZK2S0Nkmc5/k9+b0yIM/P
kfjDbq9e1CEqIqHrItrg7DUVPriDBuRlZqhCGw8ehbJiiE/TBAAImWFzfX1XOn2W
1mQ/BmkM5xVEIe2NBhdILPm27aXa50pswNh9mEo47AZmxI4Jll2Gk4ACyBPfuiTP
+fvNW8Ky5OgUT3h3ZesKXM2uEwLPZLxbNo+Ss7kQ4VXeg3ZlGr2wVD4MZTMohsk2
9z/ZbGXjboGdA+WwltG18lHaQ7gF7y35WYUCFnJ4Wug4yYRc7L5EupmGi62kd+AN
M3L+mjMvilBdcm2F9RQNr2W7VfG4YAcI/CgFoYwcD/vxj/FNMq+W2IAW3kd1hI48
2nPbqnn+j4PYTk47LFvKvVpdlzOUe2BbZpsdKc/0WiXPoyKWzxPaHPrzW/jeG4lN
NRh/tSOOWNOMmXcDN7nYqx/5UEhMgvFeUBnAJJ/bREdLSl2OWp2uwibyLQSbKI1q
Yc5rm0isDwFBoHvYyp+yst29Dnu+6uwHP+6QoZY6UYIt20pYPfc2Kr8CDL8i556j
2M8hG3G2ib3DyXHlZZgF8wHEK0bNlFekd0IyLQgEnMhhTzxSlzib4UJcwiUVsRAY
mxE4ISD2h2wImCfQEGTpjYbtiS3WrvF7sQE9fILrng7J80qmcZHcNEw0xta5aID4
XC6n5f0R3TaBKmpjJMUc6MMSu3Sr0nt6TrjQN8dYQg7ssCfUYtCJOamjAtK9SWPe
CBz1c0ffFK1pDozMvothJjdYj3KUueiBIvuN4bpBYybHYltcXWHQeBtu6In/0AFP
hDWY7zM56JyWJAnsgQ2F2nGpDZuN4aKWuQEJqA8G7jCetE1KGF4omI6u6ibo6jeR
0sHBllYaN4BwdBqVDDv4vtaD9VR5LSkAnFL+8fWC71vukDMNl8kJwoVOIUkqq5YM
+L+4GxHsGzc6KLDIZh2SdaCa0Glv/qmXENGvhUM+9hFHY/cDNFC1dpJd0JNUEfDW
8jvRrKtyePE9d5yw6RaqXRWPDSyxuTPDhGtm/Tr+cxCl2l4yDFGjCtZBLs5SZ6rg
flhA+RsFLcuAA0o5F8c88BeVqPbUErGhtx9WMfcfWVcfLwfHB/kRET5tm+5pBIrs
23DBpZyL7fkANlxIzzI4/O8oX6mXx1NRWH7FI/9bcIYok1Xg31khHlGW+9X/e0L/
8QV7cnpjR7Zt+Q7vwTYDuH8979rty5z8q+EfC8AGkGmuTGp3rdBAQF8lcgrZRWTR
e5eZGL7GLnUffX52xnOkDB71cd0XHVKRbF6c01xLaWRSQrNNBqlH7duj9MjkcmUK
nKCSflDf+NTl/MSlCruwbsmhRe2vyHvB4wVL8IM9QeQhcUwqHCUFG2seMzR0G0H0
ld6ID91q2Eyz8i3Ch7+osM3eaFpPLsAfDW9vR9FjEp5cAtpOvDN1EAKmCl3DBx+k
iw6nqMk69LSBZINUyueRuWhZsqBcoQfa5DEmBoLVHCG7ZI9r5dtb1RRLg1owpp4e
dMFNlgW/rt2vx3lY7MKydl8h6WlshnIefFyTPOT4ZlxMlV7GppN0jaah84qi4fs7
w9nD1IC5hr0/vQGV5HVthBiPi25pLAxlsSXacgSY3nIi31pB/OfiZgYfuVBfoH01
4ub3bDR4Kc7FDCjWl7xyiK064kLkudBUpjVOR5FjNeYoNidJ4ZzAJ3Ov4f2d+2SM
kRtxGHbOA1YyJECEPcHpLdeEcxottO1z1Wdb07tqK4DoYRZKdk49ihO2gSzCCCJY
B42qs+cf9C3QsFQxw5aeh01d5/AHTSl5rwyRWkho6fwsdXL9uxQ6ldjSyzMudK3E
uoRLCP6ufzfyKfB7u65KSGB00aNdbDvhCwe8CPFn6BvrKj/t5nvKRCzGVD7vxVdv
rBOXH/0WkNM/un8NU/cFxXkUb8nA8lw6v+7XaqmA8rt16jUH+uK5UBlPVVnU6HxE
PDO48M+xCM67U17Vp1fYG4fWaUIKmP5ubXYi8681F2DQv/zBDf6FY/xPbpd2SM7V
oBP6vAVLCbbWv6pZWUAppEwOw1DORMYVOv1416M5+Y1mA2Hy6+UidxK5aNICVicx
5uNnfeC6qY4/EkKUvkLk+ByRUufccNeR4C/XCU9//Lpk96eBcWUu+uhasxaf/O+r
c+QepfgzIwold6rWjaIVryzmMu8iHrHi/84agIeJ/YgxInh7n+T6U6cbWHzcMBhl
7fCiCGweqSdN/lJofStJDfFgpJU+psppo3boFvkqhJByqnuZH7cVv1PpeUB4slqR
dUKajR51wAnPtN6di+v13oNDgH4FlZu23AFnyzxseati9gIM7WpYwErFs9UzKMc4
zRcH6TToXTzUEb3Zfd2x+O1m7pfNE+eFvshK+MdjKj4jyupdF8nwYNoRwwSvU4sT
GZfWS8QL/VEJcjtmlatGhEc2Vg24xUWXWK0lcqXpkgEGGEzalN26TetBZISSh9nh
1VUVJS3Ypz8/qpPAqA/B1laPuWSsu/gJEgNqVmUHul4y7o+5WPgdG3lGrlsIllEo
jQ1gyJYkacns83d1omIuT1J2XJOym250hx3h3pRz5BwJIl3d2TMfT9bHasTrwlgD
bHLMuYIgqWzOmZQ2rfGAc7MKm+0U1mmKuXKjf87ixdkKkhjBXAeczPPpwtAWTN0L
8Kd87GeuM+PV+36znEQMW3FQfkUrwcbFWgxPlHnMu2PdvfjIgut36/wSitDxq6K/
tjb46xMGQ9NcdbM/cFYg5l8+OnA11hkVhyjKp24CWygxb4lwnRt+H2EU5iyqWj2R
au2j90lUBCmGfXnbgMaUnDQxhYC+gLiyZkMYQzfj95zJHaHRn4geg0QCk4WkOtLa
OD6WnN6uHpO7L+d2h+CsYRId0mVfWLY5nl0cbVD5Hm7DtZD3puxtr+EEw1Mzpw1N
cQ8Hg3vxvWALI7QNDw6b+gcGm2zqr+uLVRMz5uW/6pJUc5LGNip4g0isgjvUU2GH
OInMk9Tcmg56Jek+ncTP1feJcsPSuxQZHAEXqFYhBvpai8Wz2thb4pwMYzJfeeHp
ZYi4UfFaI2C2SafB2sPZzBKsIMegJWOd4EG5jRRKQWUmRvWrbquiDXBH/AMo02tk
huaWySjn03R0Zy/c8rfSkJgdeuyZVg6ZBUfwuCBvJjWVJp4AUTNXDYgmEh0YKnvl
ehC5UNDdP+bm3HYik8OaOEHR400CLOZaD2FocFTnAgOlXXFq4USQzurZQOM8veTQ
B7QXcLGwEr5VWRlMkyLrRtYl4HEf3jG76BJR3Ml0U7SBzr/jktZKwyc8O+wpf0xQ
/IeGcnaAfkVUknT5WUZqZfNr9TdVpFAXUF3VD38fZxUigmiMyvb+uCL5cbCHmp5l
G+F1rxwG79o4U232EjDceO1RfHCkwsEhdj8qL5RVpbyVg41YSjlu+jEAIqTf2m0Q
pwHejnlYKijr7X3XuRDzkfeZfZ5DpaJbJSXp7jyxdGTNQkj1WOo/nrKkBQm0OoTq
tExQW8tdEpjJvJlfHe/hOYWAiZh4f/939d06yuePV3yObAS18q3A/+jSIG5CytsO
1SOGAgALMTjtVlzDAR4KsYNxxYvYwrqfj0xwGuUdfnfQQFvFqmDYhTJf56l6H8zA
Q4ptcFkNouEUCyEN6R0r6bYdLgHNXRmcCmNNYg1mlkvwF8fOMiAcPrCcyAv5iuE0
mt/MBim2v4o30fXM4jMM4bWOiE5B+JTgcjmf9raDIO83iDeiNvXgLd+SWrykeqts
TLfY4eXUNfjMVmdj368BJrDxt97hZlnjneQZoiIBxJkfAaIwkoa+kuRrZjYBiVDS
gyJzGTiIu+59nrIO0tmTZYUJifJIe4yKnz0goNvUk8LXWeV1xJD8Dl3bPWccqhUz
QLV5ib6hXQ0LCinvdY1lWGIf/yehqujRAyxtAhVbeNt6LEtUiksormRtjC3M1NSI
Ruej3i4MumQGnql5nqrBs5qMom7k/gCx3WQoGqVNACuYTPn+XR2xtyJYw+bciH82
5kJSEMxyPS+XTPfi2jJt92MD4AMhXFdLhQy3loH60ct0KX2TmxAsvS97Lm0IpwoD
f5k4a/210d/OCzVRlWAXR2AhNxLCXdEFCSeD63n+tnylJ9Ce6qjxlLwosrbu200b
0fVcPLVeK6rdtw4poRjZfuQ29al8pl7jXYx2/C8HEJlU5vBtAJBkPupHFHZ/bL5f
4kIDfZJifw1fFRydJmf63bhgIrYpeJoVMqhXVS9EsnUN3SMYRfirU31j9hlLTj4C
QILPnUEaXFHhJaxwkVjs7pz1J7j0jQbrKXp1wR5s0aLp2wZ/l9pIEagZzaAEYNBw
IQYng7cM9HMRo8uLBzf6r+VDnVfMV9pY8/RH1F+H0E9zSdDQPCLRVDt1+B6HnFi1
hygfl03x0ClObSXLxtscMfi6elRobQaDaYhpLALsifsUB83+yrgcOz62ProuUan8
zkPNfOByf3MufjdnAWn/Frv5cb5df6zFeq1XjQ+A928yjwnbYts/rQF/lQ4VNo25
VymqVlMJ+GJJG4YdBip5gc5X1FKGVsJ9/ZjOX6wbh5XdiWXubqL5jZm6zYErRnVw
6vkPo1Q4nlUpGfw0ptOsFmVLu77nV0W87/EoVvHZiv0s6wj9jYpQ7ZO4qaQ2z6G7
u7jvjTF3eKTfsy5J0lzPiPAZmtdfkacCEpJLv3D/CufZTo9cBM7HEnOqIV8mu6/6
ZDFIlAtXBaSYmgXhTDO8WhBW+S1iy60xwUp2Yjg6wqVCTjj7++DCN+3p6KP2mgP6
slOMK8lYicqYdOfqC+QMNLYmpINkBU9TnzV9xvTtlhxb32In4ifsKLJhnWFOl8tj
nNcXQJ5WzVxVgyioObnbsnBbs16G0FETA1Z/QctsnHe/1g3y98oBHd8e+xJl2IQc
TxwJFQRN+ezoCmorHec7c5NWc6iAYCBzy95+2baqQo9ae7y9xlEakZxLtjJaauCD
Ll7tsJr/KqPXzlviKdPVmewE0CZB/31RqiW/hw9IpBYLCSPvF32wCq8bbixebwsQ
nASUpWitIDJXyIpCYnocsLg1iTDyZUit1Sf9zsHvNyygG38UDKNZ4KzfPGACxwVE
SVD4VY7u5AcdA5oj4GQeBWZ/6rJ2GxF/6o5jXduF2S750t17tee2ANoHjLhNOqii
r8uREVj+0z+Mlpz2A41FlmI5oUAJZQ1c33RcDO7T7tsw7a5SaNZsjPXGePObbztz
W4wLmNdbtzWUfBPx65993gMj+9ZF4vnmTN6U/Jcjday+vnFTnDEf2b7gncXoPldc
l1IxOwuMO1MnrlLFHU8bzTaVidTvdgSQln0TMfmO4aKxaNajaFnwOCypFObJKOHC
rUIyHOSChsecfq3fS3l5p+sQpk5z2dlOHW9HKDq4B72JeW9RfpIzqzjYOcUDiezq
B2K/BfB5c7T4CVsF9hIR7PAEjS9z97e3NOyjKeDTHK5CwUriNsueDXVX2bOO4gHH
7+Qd/iCpndZI502zVPiPE3VsirM4eigP6vofqmBc/T5wnb/Dt98tedC5/9k90Uqo
WPevcXojyFa5pkA9ceX7N63aVMFEYW9ghpPsUfrwnLPVOD64PoiSPe+no3gA2h6t
cgKxLaCUad6e2MK3ud+ze0cyFXhnTm+55XUVGa2+kb2NBTom7iLffDJzXCYWTUer
anb6s8ZgRwEOaWMzQn+guCBSraYyUP+RhFuVUdtlwfLD5wjOtel1WWJ2LWZ0XLYu
6pLzB9rmUcMMFX6h2s34B02gv00x6aVuRax8s3T/B8G45l8dI4FkzxbGsL7JBmCw
nukSosobM8X333MTkSVDj+/GHmKPc/WgW2HosOnxyf6KRJsywuFKq48c6t3iv0Ys
VDfRl38AMWoxQtLWmr9IDcs3v9lCtAEnulyW7oSYAvj+2JaOIt+ZV+KckqqQxmer
Lh20f3ONKOdp8RZWzzEHBwSVQAz+ueANKhWbiupoTMzN2bqO0TADSvcEjYI1jvFK
cUVLEktg032YwqQ/g+oFyX0g2+/TuSVMA22S+hhGoF+pbe+SYGO0LhxUpQb+d9PA
61Ws3kWwMqfh7dvCIgtJoh54I0wFUhwCdobnAz6a0dCcv37k2OtJcXxihyUBXa4O
DZTr9lwQu/j3pcWfRunQTxSMZg0ZvBUCHn9r+oeXQZrATbiu7MXDMBqwKHOHceTc
Cu9Dnqtve+/RkjPUQxiGBVnAIaIYrNUPDxGAtQNCbIFhOoaCcuL5yu92K/4T/p7V
Q7lhIuR01WIKyJI4jZNZlgnoyQXagt5gyeikS2ZTrzis+bIeBMDMHXq3a5vo+mvH
YGbhzAD0kYhliDPYT9T7XK+iM43Ex+UM+tMbJ/DB4c/RAV0mMa9DXV9PiEB6qz2f
rhSkFMnqNXqz2vv17A7zzQ41EuYVBL4TKUM6lwvCFPISNiBA6W7e/lrFBYLMGN/1
L6zAvXqpuCdcGzYP2ATz4C6UbAG35ITwA3/r3VJBp73pTRTj8i19sTNio13lHWeP
5YvL5serh2nSmG1DZ0gwiiCyK6Mh3zScWq9fpfxcR9qNH2B9beycy1tjO/3H3eDt
keZBLnllB2zWvNLV/B7infI+L5pZyX5Sxono7ckh4hGAt+oJVxtvyH7Cw+fVWfub
d1ZTWC/A0PXs5ejhDPAaLhW5DC47HFjEi3dmQz55aMUxl/SOA1J+CAiOVwQ0NoEK
akR4Vgj70+Qlw6Og+XkaWMbAgMLY+xEcxDiNSoSvm6fx5nNjN0asrDFow2xGyTUN
f9MukvLCKt18TYDhNxF+rR2YKvd+yflYPHHy0Q6HQ16UdjW+pZmJ4r2lkGGT0UEN
Uh3QrRd91TGmqMBz3ovpDUMImHzJcAotJ4+FkLDWvIb9sIt6ukvYLrS27sVuLcP8
+ARjSKWl/tKIZa+f5w+U4JbpAyqELT/TIoP09iS+n+07jh9zGJ4E4b6da96hAtFK
p4V7txSjkJ0mEmioK0ciQETDcH7sPcqtvBAOR1sBW2kRUgPrKYPjc6+UMfgWI0Ab
HYzosoIBr29mVLDvbBzR3/NutnTVIr0GTcewyYgbzCn9cimr5N/URccxJVl0Rx3J
a6XF8nH/BQafZeL5r/Bl8VinDAbsxHoJ9CQf7Q6GxmHpU7q4HwIOaT7KzhR4fpob
y91Q9xQ1rCJcHJW0w9BPI5vJnaYu7Fr0iY1Wbx7Poz/XTmaTW5pQa34VAkqa1EWo
swioiCUmPO6Uys7UyCw1X/+PJUlWIvsycLQ3B3LOl6BTtJ2ThGCYB3CuG3Mkxbya
TjAjFvTxxziB/Fhf/B/rOr02uQr++8vWa5bJUdDjhBLxUbX+Z81PUYPBYrUMBJFE
APzL3vnSmbKdDEII9ezDGmpYVGlzj9XAYQfXghtdF1ITMacrr4QjauQikuI2egFk
WB/L3D6lh2B4kDYSY7tZNH7Zag4yT9BRTne9lEJwC4I4Vv739we5T51Aw1h8TBYo
G9oHqd80g56daU0icQCtOV5oTGp7nAoP26WK/lPsEX7kHjPY/CCVs8d7LfAtoToP
49rFmF62GemRSJNPRMcEwRla+3X7J/au79uAsD8+7Cg5u9nSN6CABvsRUbIdSPqM
y83RRcPYcECekIuerZmVPXTJzOBs6Qkwo2yGnOjj93KdoFXfegd2WUfVaoHp5flP
aS8cxiwngCRNBl4vYuEK2MxlUacZVhoVUGgMW35mNsRqRBWu+U47zTu4wJANHba7
qgnD3MgVV58zX5WOY0p/5i5RvjA328Yzk2fbSINmuNloTlcbjbT0Kl/I7ZkpO0he
fziUyXz+bscUum00e6uSKqHCXrodoxaPl+miS3AxdQGd9S0M2c3moYMHc2nakxRX
x4aM7F1YGO6szcxSpQApSgau7xE70wLCFZmDRWF57lTmT2gIt0vyF/kwf54hOhBF
RsVIsmfhrqopUrOA6n6x4fCeduypertrivCrpeJvcAEw8Fh2QbCtAUDjQfF6Irp0
cIXIIkQPis+180vZnwVFFKn7W+myPxRFovKsxEAMoA/C+Ell9Ic3guhZG3AVsbj8
r36ftXNnf0MpAm8ksTm+IajbzpMRw1GkLsab97Y/CDYhwYYzL6Et6EQNpvL4jWr/
OTdqkY/kxI3YsdOiJPHoEj2bMsnpcOR6i/ZmK0NvUO0CRbOFPOiBc6j3xyuUjNtv
HO0zh3gDa2gtEVgp3L6HJuBUkHJPdLzf7U6fBTYI0IDMNd1GE4KXdxiDYFGO+bD1
FRDZv52tONEwN4Ro2eY0UI/tDCZpqd/feilHXaECu8HnjDeHwc9Lpy/Upf4jYLmp
qiJA2mwZTCOH7roHJC/zXeq5gRGMvHIFLmLuHZoSAiRTiS8dfcwchohVR1VOn333
iGaXkGGAmsP/XVZSv5mgEbRZxU+UL3aOPf6ESnnAJjd17hz2QKgB/aRJDC6tK/VM
0sBGjh5xtmhdKaE9DeqQ4pr9MAxvdXEvZeh3NVV0b32PjcUeIp3kGsoFJgjxw6MG
e47zvPin2EFs2UMqrZn90mjDGRv+XXySgA+UKbbZnC3PbiuLm7INeeFFay65IxDt
BrCSvq2wUcWxLWtk1/qwK3Al5qfEIXxr9+lcGmGFP3qggdqQ0cAZ3E8BiMG6NBIK
dD1jqQESc6Vj4COBh6fqpa6cbKx1KKL0GK+/MscZWIzAkBIfsGlwqlpvAoGQT3Fo
wNFSAdia8PzYywIkZWMnm8rzFifJo1sjBZ2/Pb+/yiWZR4QxDDIfRmULl2Ec9wxm
nQbmxs7JptVSycg4G4tA5/pzbFI6NgkHZH6pgZo+vOhm2zErvvxds6G1XZNhdBsh
yUupymRzKrL1UiH1Zc2E44Oh4ulg0QGI0EW/tM8qr9xGH6FXnRfcdDIrNHMO0kTp
RPneJ0eYq/UnzkvzoAn+5wKYnB0O7EGHIBSlJYRevIPkumODQD60Hei7qeI2mKsC
l2o5jTzL9a83NyV080p7XiMdXVgURtqxBDV5mbDZEYMTZiHcWobMDVnu5h677eTu
vEMx06JdgvBizZR0UwGWBmIfsTw2hXljzCS1WnkkgeYjP2UFIY8SlJFIbUrYCLG0
Pd8LpJxsBmWakbFmRyrZdi+qhgjsweXoCm/8FcoQPanbq3CCIMXA+p665F8q7eJu
YZxbb5bvORN+TKWHN2YusejEI1IiEYVi4tAQHfzdmjYB2X5AKlDCy6AaqnxaZsXe
gvFzAsEjAhfshYzCbf2rAtqawi/9k/CJ+WVeooqCImszBPdCzxoYVIpwMUVsDbUJ
l0IIPBolmcWgwHMwVamk2oyJkJ1FH9zTnZucq3vKE5RdAJW51lTY8OPWWzkI26Pv
zknG8X7N/TYey1klWX5vb8OZE0k2OtAp8Qw+6fkx2wxtNHWnhKVDlyNc5lXKtlcm
jLhRUqf9c2U+GdzGrNoR4nhBRKVt+NLOHuLeG+1L5oHC8QTz/zwYDlZo1Pv6mYvf
Ep5TJH3Eh8iDlTzwzEx5Drb92CdajFhcxmlHkjG+CjNPLQdC6jXLQohKVIHNJyaT
K1km/0FQanWlWeOcqs5UlOWww9MZ3bZ42AFIzLnaF/GVNbwmf5H4KK3ICGq86qKY
VQfGYeAu9KSSts8JGLvqtHdlLMDqVsO/xKIHHybS7XkVvMfSFfUDMo8geChiBgq4
xGJ1vtTgdnYY0uHw9qyIGkaw3tJGenVgF1K6JlhGgai5Q+hcWzxP5sTZpn3gJFwk
eY+pLW6vQACicnDE482O1TsYJtX3hONO9lPhD/LAm7mIDPQ0+cbIJR9p5AwVhTp3
fFpP5qnXe6Ei0YjnYC48YkUdlppfb07z0F2Y333bkIIO01BSyujADP4MAqNR5/De
qSYyVBTiWf8E8h7xLM4NFintknWrWFNmfPYD9I4bGEofiSGd2t8GF/qn6slLlNd0
dR47da03YwgJBLSApxYDz6sPAsBssHYelWQSIHQvabVp6plteQU1GtjsXTc0Ly/E
f8y6Ss7mhLENo3ErFgPUfndhBIkiGTFVWV/W1OEDylP4fbvRpeZN5q7o/ytGU+y9
VSKBiC9N00C4G84g8h7yf7ynJroVLwWAMKwfZ1rgLrYDSyOWbCE8IBF3bEoPU5Ik
HAUWBFlxycGr0wwmLFGCZX4SszWY727kmY1fFehVQ7AY/kam+w+PnhQLruRxllTB
RqXayWtJGdSiidaHeTiOg3NTa/9c5PEDS9+2iFpRVdoCqBwi2PffjMoTVlZbgA7z
vfEXXOXdSAR4kjXDtAWcYYdIYTQVgV+3SMI5ak2IiUS45qlLgrJ0OFXuH+BC++uQ
d02bfGpj2O7pLwiqSIVBQRrnZqdvlKZ50PzyAaptZ0Ti3NcxrdSUb/xdUz6SkUmm
s0uBCtCAfmxkzuDz4LK/HfOQs9k5rqGVVLlhsasUwMn2wwmXAo1FK2GyhAZFnPft
6mFHVe1e00OQ84j6wjcn7x0hw0Of5l7IZxmmWle+BIAoAQNB/JXzEexzSn8dcp2C
aMorwKcwJOZ/ft9vMfum6gNRfDVfV/tjRmjwTA98WHMd+YCbSQdJMUObcfjsUzaa
mCVExO0y/2aLwV4Dti8wIxxpIYrBfAjihax0dvPtodEwc7KC/YXsgMP1BzE4AKQX
oiM/kd01XChV5uQdUtUV3AJtA6odqWH0gfUhY/Nq7xFFx2Jw1qVlOLFiUnAYZ2vT
gZCukjTKiG9+9hdjE1qwaa4MaSXMN8GOMXN89D84ron59ium8oMxlay54WVsMVyR
fgK9oc5sfQwWKjW6mCH4VvY33Wh1HCykp2Hn1bUJyVjRs3VBDx3gasueiAhBY87h
j2TVkpsofNwdHEA6nUxoMH0RU3cOFOSNzmvY6WxOgfgfonNGH2g4mdy2krxbXRQf
P8hN+i5GQG3h78ydnIMDzWwiOXj5EGm/5j9HGrSrBtbbOAUe8fc/1Es2FQQm0NnT
mnEhkF7K0sXg/6VEVdmmoEv3fwITo7OlKZyNIzDw1QMDZJlPCnN5sG99Binfv9Sx
nP+oa/5CkMNYgi19KF9JX4sRPqExdvu77hyEYF3sTvtcnshk1iwr1Y1tMyzMAvlZ
J557tVLKvd2JpNqHcfUY2Mr4c2B+zVzyF8hfSI0yxxNAX09p2dYu5SVk/M/KTQRX
CfS/Yd1lRjObJ38uPOHtF868wysoSseVs/uBuzDssAkUEoOHWEyppnJo5JtKe9na
Sq+Rn7cahyQjGHPxUnnolOKmBfiQZmKZfgD9x48QNNHNHDjnaapA/wmrKbWjVx7y
eIy5e2khlxSFv6URXtUOOaNTRHKqPiTIWyXnQs9GISamKrKiPXSKLkwujEWKHScW
tRG0AUjY4TByRA7xRn4L1qLDUo5D0pJqSswONQJLhF6tHeFrrLBqxz5FuxrFf5AD
ceCmj873wMpHoMDnq61CzZbdr009UR35WReeNmTlMnsAvGz8uXUp9+5lZ1XP8diN
I/3XlVZ4G5FQztTAoXScHtHGcOa8WZGDBY6YQ9pLZaVNls/TjpaSU+qUqGMMswhZ
AHnjEAaZ3MqZGsU25PSzBc29pZ4CXXj2o1MzICXq4Gbi1W5md9ChNeQWwASPtrRJ
mVLhzfJ0OfVCnx1id9nMWVEEaP/vRqwLJaSVybPPqCCDm6c+L0ZvAKkyGgjh5TGm
duw+QtGjfs9uEzvOAJ1ICODZSaryEjexBc2sIaeOwhDGoZ/qRu1MZ7arXqr1lUgQ
39LFKQXLR4O1BTQekgf/GJxJiAiEmGisA7xvcFyBjt3Cnx63Cl4UBP/jVuv9fv/v
fhgq3cgZ+w1aqDoSUWdI9FfTUiQlJ6xyAnNMW/b7Ol67vbBDXYXyI1XhPql/oe8n
hU65znDS4/aZHxR9UIsdaqbRj1HWygv1uTypX68a+SygF/V484C1uh6BlmhqK1hp
y4tQSe5gPekG5UxRXMNBwwGot9Ic/1jefk/sHUJ6cqlzq8brcd0Kintz7lIIyTzm
xnpwo393M8ShN0svWfWA8laYNFWjPnihTlRwTz9tl+WmYMbVpvQNk5CPJ0StRnqV
8yd7InMX7ID5ssFMamAopcOz+vMdRZ9hnUiNUuxZG0uh8vOzsoiIQ7uJhf8NujwA
SW6kv2uOWjSQ+njUczsu7VPG5yUU7VgRxyYmKDVLfXnEGnOWoSQ9dH3RHIoYIWLD
UWTHkPOjrD8Szi0Xc3bZIg8qtrkEwYH8CojgmUGl6lBJ32cAKcv+huxydnxDDCAZ
fgFjg/hof8yhRnRqhftZJ0vZgvoUzbJsRco7NYhKT/xG1IvrQ9ILfFy5dCIij4lo
0Q4eotTKzMj6RRk25bJabjx3apC+b67AVsw3RaIXuBk3CGoKiN3kP/OYscUDFh9N
l1DFDqET3YyjXXjyy8NMWHnHensh9eok2q+9y6tv6h6NROFz2jikXT4KeBkgItns
IFOC6EjUooUW0AHLSbIi19fb+XnteK7+BCOvCIP1SSQ2W1Lcst8cxKKX63h8HK3o
zootndBamF89Tr5csH/8mZ615Y2Ng3rM+gJWt/tCV+etU8MYSUFLYSpmE28mMQXM
tLpV5AuofrfKX7rvWSWnj2T+9qciiTMc0TGmC6aQuQhHb37XJ66yh4YC7wRRUUsa
KX/ZnLAcSJrSZ6r6u92D+1ViY+ow/ffbtSRZ6aHi9Brdqb48WOgzWlVLMQ2zaafy
eHWy/Yu0PDR3T3A5Iv/81rzNEPJ6Xwn9hL1pKvRfzcuGMDuw6VKEkn3p5Db43C2T
FjaoTKBS/1+iQNXOfBX3DS665HCrjN7LDWxSb2VHyyVQtu4GGd/PtjP0lHe6sRU8
4ONkGn5FW/Plk0CqA6rRHjU3sUm0+rFq/of35BB2ZRFQLcg1qhOlX9FUItYbsbXq
OpOtQMMb9FKBMRLnDOirk7cfPRfULdyFZSZJ0yGLxk9YMmAKXPjfb117Jg+1LRQH
MnQjoh99mxbLgeaggHlacXJgHS2jkkpS8Lv9VF5MvT5a7R1Uk3qDc40Xe11nCRKq
UBikcUFJFR519j1JmRS8l0bexOR+YL6VRtSNXwZAMQOA2siEkvZ69P72uBGheSrD
14LPJhiRfFihlmnjVnu+S4zH5VGgUGtfT9g1WJC31XqJNMm66oNMJeuFyJNikHB3
QYs0IBW7nyONvatHDCQM6wZTYjsWYH/Ljgymq4vlPeism10Oi1qD4CI1q0m9Wdzp
ITghHOaxVhYHc26p79dMEbBrXUoK2MEvaSboDUMTLNFWbcw6vb35+IKxk0NoBP78
LfzpgfH1EZ4Qk1gQ6kfZa8coiPEKHKlImkCfK3FdHGKVTfcug1z0edYdS1JgWxeH
L0z163MPIE4kzjdhzc04cgl54N/x9L7Q9towq5dGmogHrTRw/DDJ4jFd+HiPJhqC
9CmiS0rtyK1anplChiUWg9LU8Vbujv8shoByfnVpMX0Jl3NfqMlgLm7SlGZmlgDT
ecFedyFkJkoiRW0F7hRzc+WKTzcWjeOFNHGkFf9vexcOCI6v5gNBUCjyNQIv5X8J
TIpw1RexIlKdhlYy6uM9lMwK+loEN62mbsiGRvrw00kaGpkf7PjKyNKou8Vynbl+
uuR9cIYTM2oUpBWZhnQwWHiKP4iO56F6s+mq7KJIzNMJ6ZAg2HHbLMFOZ5WOtcyN
VXRrV4tOV27ZXefhCDA1sba/HWseesEQRQaGsr453YPOZ0+q6cDvElL21I+Elx6K
ULMwEHpLlhuo8McVUYCjYjEHHp/PZF4t6YPhchAbTXmUyDO/dGKiIXWrTdsSvcZ6
9RxEAQprkwUpSylRhWQVX67Z9MSe+VkhbY9RkHcCHUnQrn/SR5DIotSbPUsVgsJn
7chxKStLc7UtP40HQFTfbjb5DA7nO3Sh+epwEmiKwU5611yag5HaL2C8cqQlXoDo
tHToUYxZbUnd7uSsTDhFF2WJ+dPSn2MxK3EElJ2dPjbty4nZ4fsnVuGnZ6enH8uf
eU5/PXdrLt5hyXZWE1QUDAsEIfG04RdOnLGDH8HmmJxNKXF6buDrhpMChyI7fByX
6mxRhLdjM3eub3escqHwhZVFqwpwOFQfH+bQq15atiPE/jRgi9n6+jhxSLdSJ7bA
2f5rE/WKrjtuOI7pJ+G8Zzn9RiHIViOAAHeB+3PfsInnJT+iI5QRJXqifjZXh4LM
fjtzxKBC7BMWR9AgQTz2T3MM5aIEX2UO3zY91oho/jo+1JTnKCnQuvBKMn4Q2Nd8
g7wmjGVX0Pqi9MblmnZ32I+o+GR5G726cxPSyfNA5l/iEvhPvAY4DWOI8e8YCdf8
Hyh0xCH2xAgWdrkhaJ5+l2EeGeh3ACxF3LCwtZh0VAEKEv+elVd7sywC5lSYblxe
8PNdtGEnJosUSdvedpcJIujFpYRb8aaIWwiPVzwEub2tkp1YwYdc/vuBBbIVQpzg
zIU09cMO8yHs7zJZjOGEkbSnod/rMWMPxPguGmHNBZ2gb9lT9dZqMTlSrnNKHRgq
7SP1hmu6KirNtjIb1nsHdzAjYv9kKHgpH7w2MAz3dpzKB5DrjCPztZGzcN/HVPFl
As1ppbquFyrQ9C3vZSgU/A2zPyASVjywNzl5FW7+E3wk47CIeC7n6U/Vg59v6ttu
RdKHXq0E7e63u8Zy3kfzsj+UoKiIqUe1JaNOXVWL2XPo+42QCHUInYVjq+scDANk
VoMnLcUIFjp2+u6bBLO43kFtL6isO/egJHYqN0av9t4JmO9aR23P363oTyoTjHqd
+ONr539jE3VauhHlX8umsongWNcB29xOzKZ7J9KJ3W2BU1tSFWvSlCDguGvvrrYE
jbiwBBIpUOgFjD8k0OQYrjfiVpafAKPSc4vCRmL4uF4igt4P8yN5zQgl3eOTtqdc
EEArKl42QOkEOc9nk6xLdLIQHHd2OlzdXGGOfcL2TYLP7oE6ATJAMVCKesRQX9tq
Di2kRsLYmnP2IE8rMBii+RtVNjeIyzGQZETJB2EcjDqtgXYwF3XBfLCKXfhsUeO/
HDY19Oj2uqk/Sjld5EPl0L0sQ0rSN8+i/B7Bj7VK8lZ0WGp4yBPUUevsurOaGjHh
tU3rtnx2r9FmBuBSMA60fAYOgg8BlkxADCMyv1tgLpU5ysB+ZwbuRR6a1ghlPLKC
mnXAeeJjlrSp5robgbuTR9+GAKs6jwYYp5yTVKBIv13u8MjVM/bcYnUVYDoVs2GO
LWiuUxu7V/kRYr+4UahOSKaMkzCmMjmRr7sPMiaAverskFG4iODCpa2ZsKYC+okz
UTTsQQDrkA6eSQ3Kle0PiWV81NQJ5X19L8D06D1HtkEZHGhmLKavy2Hcgh7odf5m
uGGRPaPNA9TmoEcdVUPu9PW0+J/xpu4Tg/gw48/2WFCW/KBQphN1fIUKd1hoS2C/
k+qGj8L78DYnz6R7N15zIe5x/IcGn+Nwg6E6XP+AEPlUJ40UKooZgS8zpqeiTVWF
uInti15oEgax/dJg/kKDcgTu9FSfsz8cwMjeQqso9zRQDj7UKBt993U/qohrG+XO
xLTIgCUyyngJcD0FN/EpXSsgcEC8J8S7WUmqMvJlpNwKeTthhz6iJUGe5mYBXTOj
y+JtmrWyYNOD9j0kvbOnmp3G5DC2l6ctNTzI4hQEhcV3gph3udYx8FpTE3P8Udqn
r3Fu1DlWESvFfUCazm6XNZ2+367y9uZR2APgBpz+ysczTJKPRCLLIw+egDWnxXVP
pB4+MtsEZYc8F05HvEyAugMYAsX28U0AeJZGRUEfpxQUSmnRfJEciJwfQpLjLjQ7
4x4GgcTW6865W4T+FK3z86HQ/BYUS7t38+Bn31WlI64vJgUf1buevxdqKYuX7vLB
ZYnrUYqlhqCAwZd7/78VrBGdj2An6GWmT5G2vrCgYiV/OjDh45DBkDLNlR46HKyN
HCJdZ1M695tU2ynw02VyHQhITGqWcpifDIHCrAlkhDJxg+TQsp9F84uYMvVZQsc1
KPgQkvIPbu581mTOBpg2IKlvxgohvr/U2G1p7YEa0/68Gl12F0GljAEBAZK0sbAY
BZ/iw2awBh+MUpmDYNn/lKOg2oiT+mM6nR08dDAg1SRZaTdt0cEMi2yDuhkx5HHM
LmjVBjvPmhHPNMmfgBGogORvDvQlMxhWmjxaMt/WmAJqoZhwONm3wlxj+XEWH7Dv
r2CQa50yW1x0wN83JY1/RjiQiKKGMICLDIy9tEOTmJLzbzCeplmrwJjNNb8PC8vs
ZoGhkcYDw1g7For5x9zJLE6QRZ3YuIyCroovUj5twVYBbuiDMA1h/xHUEa2t1br5
1S/ujKVwWcxE6nCjMYfwdZTDClUuynCbr0cF80EKi3Iz60sFZpoDtE+jMDnOM+d9
H1D7XwM3DBQlnDC7s1GJN3MbCjHwF6ZcenQ6uCtv2zS5aKesMQygjBkFj/kfli9/
pxNxI4aQcHVHM+9m3Jzkm7pNfq/6HER+qTk2iEZYuGhAa7ll1A4Wcw9aPeP6RXuk
YqecNf8vxroKoUylEy2Z8HxKHfKMoGJy7kpe4/V83iXVvZalIttLaAkcVFPhpb7J
ODX1M/DuDv6SRraCywp75m6Pd1t6URkZbjmZp6SORennA8LbY4Ao7mxzDl2j9xP4
hIgtL5P1RRFe+TWg5szXZB7fEaHu+R/PdPkZRNgy5aFlKOe9BFK9lp+e2oLvzhIT
aRkIn3/ru6FuGdxcbmQ5hrQWw/z1XDeAEIjnFBZYxy8zse8tQue9bkMll2q7bUYY
eZub6r/u8JwMRKVtTzZbO0QuqaXsZhYRH4YXMfW6BKCj9hSlhsBXBpGSEo1k1kGd
v4fn9u3y2kEwZ4jeuYKfEZnwSY7orw4fOcxmmpop/w1VFIyyWWkwG/M8rUQaR7CW
pdJa3INf7o+xNTRKk5XEi1Ld2Ga0lddCnKalqM7VVwRS4NyjULsOrhvMo72rSXNr
wlk9yLkDXYiimWJXSVr4ZaSUeZcpFggUouH7WorxdTZ5O6jECRF/NazIBMF2uaFV
3Q6cll1GqFP/GhU+NrLoT1IP+VBdJh1xymZZK8CGgd2vGSi/9UX9VWdt371Cia9Z
HXPlEl7urUtpsDCWdrUkSRl28DCV64A9BTMqbrYHpcNt7N5F/sY3qFuDDGVbRHaB
WotXl4QM2QO6vacBrMOVYeftTZYo2X0ooT8uu0+CHo3dGcL0Itlx+o13DPQtD0WK
XX0G3diWtZdL1BtMU7Sju6+ppPdVGX1L5CTB5ngZ42O0IQFpBtjiChwuBO/tbhy1
PtqxpgiJdaHnknRLaJgvG4jVfPCAfB1CO1AlJVFSVjIVU4HTrXdspv8/ApG8wO9a
JJ7zxNLCuBLXYugV5avjqqJztXo7IiowvBXIcXB2zPPwRuaENxWZUxGq3vo4Gxp/
rjCyRNKcOABdVseu2WhJloMX4LiS+XvPmRbOFXPEHUFN8XtLmGYrwvh5VUieLgss
V8k922d125kv7h9XtzB0m5QahWdKCXmpHzzLloeoTU+TdTy4hVZuhWvNj5iRyaRX
xhXuV5ZtY3nAn1lOGRBX+TCj+Cy/L/J7gdnNulwx/8jf73QTaZg/tCUrx8OntqlQ
l3P1ela5HlsD1unm12rrA21Ga9b5FJda6uOrS5h6YgdyIGvMm6LPQZXAtEZjvWRS
s08VKGVgbz9hI7cyE8/6yTEITqm5jDfLYyNqqldo8eDDc61nM/Tgy5kjoIBYh9DZ
b85CXOoPQe2uQeYtL0tn6TEuvPkGBwW5RS7Ou5LnsTh4O4alxhieA226Pe/KoP+G
L4BFam1Rm+fynEfnpJqHhmF8CuoCRkELRjw2/Py2q1JJVhF/AG+fVXqnchKjsDkR
ejzWWxTAwq6RhMikJVqj205bHUIiGM64xh/XHvYbdIp5ys+Rde7G1GErcqvS71vG
rA51omfmHFwFRFuOIjhbgnolfcE2as8qC9Z4DKDX1WJUg3ChdrA7KzJL9uM575Ax
ePGhj3KqjzDSWwgJhLTYX3iFSPy9WZSSKyTrHq25Vft6MTkoxKrNvAMDdXe1L5cg
EMqVqLIQVKF5WyQIUgBdC474qPjlu89fOpoJd/+fmdxXpHnwz6DHNtUqF0vy+LDy
LFFlVl95mCV17Jgc70jVeXsQiNNG3z5ZDbbdolva27AQSiZilrpluR9BEu1HNsno
jLvgmCTuoZsY065rleOFRyhWzeAZVlRcBcEPlpw57iKNWwHTI9qIm8tufuQxyv2M
t28O9Qkg9efgWnPuGeiQ7HNmiQz5YsnDfLIWwAI4hvLGpkG7sGOoVaCYUk3ztfTj
OXoc3kj5d9CDdEN8qslI1+nCNyPdcnt3A/r9VHH5DcuMfKgrh8DPqUQymueRAxcH
wp06y+/4la3Mh2tLtX0KnuE54b9YmtvnfWRvpRJmJ4lTJ+v85HTicT7P4KB3i5Vk
XlDqsI6vLd21f156nyDCz6+Ni2oC7tfaJjnKzNbhdFRMHHpGc94OT3WkonFrcDHJ
+IgMamj3aCe8xTvS+iZtsIoBLyalpOsqUkwNGspoNYUa3bmgKJlcLNoyJUpDEUPh
VKC0M668olEE6DfwXxVFPHNn1qTnFBmBu4TVXWtJr/kWGGZDxqyk0rboCrgIpgrB
g20YfMR6a4f66anG0cMpzEf1klgS8c1nwUa5h2uMW7r1Hjmp5tWuHQWljL8ZaAKL
sGQilPKoAcL0VwKz3+AcTsdc8XtW2Rhabiuuu9t+0iGdiJzODVO0bWCOyqUmzpt3
O1shdBu5N+8/c8xkFppkDzj5WFodFk5yp2CZEuUwXIaB9zDcg1xvaieiGmaYZ9Xe
En4YehzOAxRixw7LSWL/OwbmAA8RHJW6SuMy1UD4wraffk/N73/PatM8yxYzmLC2
BpkyUrc9oUyXA2gD9O4ltNdRiY31nsoaP+VFd1yChgN3l6wozDnSdxXvXtiWUcFR
A5ccQul44oTRigWFRwGQ46GceB381Zx2es27s4ST+dBnSTa91quL7KCsybxXdVy1
RJaYi4/yzf92cQEKbulWjA4NEdmqg9zO0ijiLmPxn0/5W3lLQMzGsomuRtT4nvW0
3X00jnQfU8t9PX92d/XIuK1DO29pdxz90bDaKZceaM/esWuUaIlJammxejEFeqvI
/rSId3jHUL8u+yuhJv4j7W6d0HF/d7cpa/8tEZgbD5bDpqOdBQEL1cGmeUMZ/3yG
AlbVBQBShQlAQSe1GxDRqFFafNW6cUPlb5LOAphGptDzo765ItygwzXNt8rEvB3N
p04xo/0OhmxXJvNqIDqk5ZSMsok1gdmGzo1Szn8KbC7oMm81CqlPjwH/uznFnPBu
9N+bkMCZXACQQL6eQCXZJtya+WXIZuAULeOoWuD/084DMRwTPK4h46kUiUDU+tY4
hP2b2/QskHLbH85JT4MRSU2trN6tCyJKX01PLn6JQR79SWnWEStIH5Uy1N2YRLFk
NMDMz6eTzTA9Wb4unW4xm65jT/tUVt3EO5o/Q8vRkYytG0CMTEdvreFRreo/FBzD
pciXr1tbFK7M/lSGvMSVz9pTc18ngbhgH5/LuRFIamYQEbZs+89i3Fnw6tLfzUSH
RqfQ0H+paJFXH9x2rfD6q2zI+fiGBrSVt6NGoB9Iv1aGot8QMdgtfia4aAjYuS9Y
Pr+oafzkT1Ugu/xzozOwavogmxbgkQd87Z/RpqdxEJtSPHHg59/QmF/ZV5pMpuvq
8pDZ/vd1U8zFMfpRGwNXmAt/oQ+WSfiwE9feic9i1J1BDohVJInJemFPlmVpahef
oDqQ1E/vcRYfz+2EsHhM31qEIbVAblX71rYGdtcLmI0cmg29CVYYvrZPIKLJ3SkJ
ifzOdNn0plvFKjIEliBKNaAhldmZiv9uiRX+N5P8jBMt6UMpHa+H9kBTUoBQs/g2
S4W6nJMBdm2OcLOC00V109T+UPr7zjOB9Gujwjtg33zbV5yXqp017snWcDzaY2O8
0mCfqSTLl1opgd48pfgRejPj4rqZmC7mAdu69Mt3Mhq376Kj58wk7UsWiB0/1dTa
tyySnWbhzVzMZmwTT3yi7fvRqGLEHgemI7MVCGJCQ4sl4Zn1C6OVxBOjo1dN9Udq
C9x4W3NISQ9aUoloEBl7W6oqK4VYqNYEv7lp/5rmHI8pxeNcTZzfO3O1NvVOUkdB
AhgVJPCyJJplYF1Ft0Bz2mZP45kpTboVERi080xKxYEZ5zBi7sdc/2GZua4rWGx8
iVrPNztaaxaKnZv3NSguiTjiPfqOMIVSDNpgI01THDIU3LCifk/ZN7gWdVq/93qn
AVZpMTj/FIIr0kUV/m/nCKq5S+sOUmHpHfumVKdbuQUqqt5/3BHVV2YDGzo6QcnW
BcGB6fUaAjHvYnCY4lbITkLlEZiSqI/yQM2zCOFb9l0YGtoX2P/rQwTTSnKKG+aI
XoJtRIdhZHI31oz372ycwdIvg1Mv/4QhXaYZphBBLKWegqt9m03AnLcE/7F88N4E
jgjLgBfLWF0x/LPKa8psEF7ZO2OMT6lOcFrUIizz3yDhNHixw3C5EIVCTTdRovLm
eW3cY5UblN4YI60UwjDcUnVEEekrLdCxPHvxC7f2sPSRoufkpE0SCd/JkiVVn1AL
fbGFk2lYYlZfm1toyPerMKu9cxqH+WdGMulbltcYDBLvQS3gg++B/TrSfVNX9HCk
GDh3Xwp/zhmDI1jXKX80t4qVfWIj3bxpdPiz5NAkSAZCEMZdrLLw4mTlPTnHURto
5F/TNrBL9FY0gQK30uiHWZi46RdZ07+7rxyPF8n6gveABWtpL2fhyIcdlL/xFwYQ
XLw+tAvk8agm86p7k1nT/pXlzZZ5Jr4wajVL5venSBOcgxkAcDZaSNVsjzF+KM1D
E2Jsg1nwGsN57rbMpRvDg5/ZtsPtoH1Zh2DOVrJHeVlbUmyvO14P6gPqSzXfffuv
L0ylxufOS5gecC+qxTke1sIiZdNyg2XRr49FzRxdmfm0grEASfHZSnbZjyh2ZsHK
PZJde4xH9KktSY1u7QVTNEfbwf212Ruj6zEHFjJf3JkC3sPNimzjQoFwif7XMF7N
ZAq1mKwGC0BahnG7adyGl2zGat9QVE7oLt3IqVgjB1dJLMtLt58AeM+xGgNxKRC5
QlRwfdEqOeAyY63V54+I72tqRgcCzbMhTeHzhpSaq1ZLRBV6ILu11tQ5b1yEJPc4
0iBEnFv3ovy8qiW//ULZZcGtT2bn60/BSGbUbKdwUHNF0mBtgk0epV4BkQUZ+A2u
EkDqZTpkZKAWC7v9c+fHp0vSJFHiDcEm1m4YbeQuMrFwiLY3BLQv0PxEaXZKPWvH
D8dm6hWOxyt9EZ+xUEGv/tRhCYka0aJRLdAdGDCHqRZzXUElCX+ToMh65ProGnJz
Akr34v7Lpn4ufIwpApIl48X0lUULr3PYynz8rG5h/q+0rihFISx1ZzK/AsXASg9W
qe7+jbQdBgez5kSsAhTBk5p34272DNEFilh3ZH2t0xv01ffrL26ImRQZPFXPY/jD
K72tL7N+8E5t3MRF0d1wP1MIm1mGofJaCacXSuoliNc+y2Gel1ngRoi5r4pI/yxS
eFxu15ncEXKwFsVfAe3Lmu55heqG9saEjOKJGXOWOZ5mLOtAb4cvWi3U8PPAlO1k
WKWy/kXJucGYH9Lp7FR3KJGNpN8in76w1zZVSuKwPguPmEYtux8PY3j5Zaro5YAt
Fc594JRWwJX5oT6KPnIjhZnhYJP1GTKX9YB1OJfz0gx4n5Gx2ZnzO5Qr5Xr+K+mS
a5PMDgqaDHCgJwV4KPRqKLnbetI/yrIwyKyBYCjiZnpEWSx3Kvcs9urkwTBOFDE5
hfng10gOR89HX4S42WmQXhjkdQycAPWEZYFvzIl0Xak59I+SDYYeB/z1wm7GqW1C
bkyMRb0nbCTBSiq6IDgyFzB4UsLUMeYzkb7vlcUFsFcA98o8FcmPbruoUZ/8bnt+
X9G14+F2nl2GmWJwtYIMT5K8D8cm4rHw914E7P89I6r92XSvqF1bvcu/2TNWc+Cs
34f9Ip7RMhKFB/6MScrwGEWI1ihUB0u/i1Dqgzv8ZO5qSISZyd1uqpg/nl0ryqHJ
Wg/r96v8QX2+bej/6m3pNpVYJ9EBv7RG+D7i05lumN9M/CvlYR44F9tMFTSmTTLb
O7d/VwgYeWATOWjkFzBxuOrLtoaceTnMsYFqi3SVuV4f/bY1TTCNIYEPPkTd0w+Y
huw3Wyyyyb+yg9VcKCFH7NRDUKqPzPP1/MuisFodiZGfSnHxTSGjyvqyMtSaV+q5
ZuQu7u2AuA2zuuFAQi4OcQeK9CodIWxddAvWiz8ujFrEDDg4S6FTg18HGAh6M/+o
REJcv6YaT6CO4JNFLeY7BlCqT7S1lnyXJq4RKkeRT9JfSC6L6wN1+motSwFs+77X
bLWZ6RTVsTEfbjJGWKDI6WlzhZlxNdh69W1ALUM/6URNwUd95da8YvZH75Oo9lAs
nloo87G5DPmFOrGRCGfdUY7M50loblIe8Rsv/Fq+MOmSh40qt5QpFUdyehkqNcf4
qjcCBtGVFCN/k5s/wcQAFx/LsUHXz/z05tU4WJAZTqIt9hc9e4EBMlfMtE7ohlC2
W7KJDfZks7B6OjWu4TEqhCtlJIHBb+/FS0ZPhibsxjhnQyTsJi00KzpuZ3Lx6jav
2AcAYZBJSbi26KW5jl9+JUyh0RtXBDStm7R7QWnPnmaP6jT/n83GSeKgqoKqB8mV
Ga6P2qDR2Xqrp0yBN+9rACAv8C0FmzL32/GOv5AP4oOZE4GSsQbyDIU/Zt8FRkP5
oOl+CJTogq/bc6xMeroBq3K58la8xq0J/ArEv1JgbL19aetOWih53gXqAlAKCsRr
051fw9VCUN8mpyKkS4q2LsBgkvjjwLBLeUXdguLK6KCq1jwZ6UKTSmXQX9ESy5+n
NWbxpQLjbNDYgkaHIlm6Sz2bNQxE+SuMStRl+jJ0WOnqbvRElWetCszycUPMb5z6
HKvxrfm/Ek9+o4ikblTVIUEOEDSeaF9B5/NNUHeRix/g8UxISgABSCF200OZ3Aqw
EK4vmFgxH+VqiPQ2EmX/Zi1lQ5dichRbLu5Iesg3tUxuJ7SbqswqrZY9X0pOvcez
rrMJ8Lv7ih9jN/tZs+/0DTKWbSgb7GZpWXoZtbXFN2Ck7w7XdeQfAYMgTpIR08w5
iM9OhusjRhjhZ9Lmlyyw/EPH0VPrz49CdieKBMYPMLU51ZUxu4TA6JYPMrNxxAnx
MCrr6JcYZFJuJbayWsoGpRgwrVDOL/2s+Be6g4zByVMva0pWVOTcwTmJzr4HUqLy
Ur3oDgOmwKu2lqZxBZnD5/b9gGnQ39yfR4pNDPo9AC3WP+TIMMePSmuuhE+P3Py7
Blmshgt7N4LnG6Faiz1pITY4ezkcdPdsOqajvkCDAv42f8/F+ZlE4wCAO0UIymi9
otyEFmQsIIGJFj8hsJwnYYl5jRoVHdQorNjzlBansNzl5MyJT5dgdtQCWLXzpNkQ
0tkEJlQDEA/6Gt5WyNeQsTLZVi3WtdoOl5JhovwP8twP6qez6RnVUqqMaNAKbJvo
IBAUgXneLsHoNbD/+eQkjEwbZ4XTfyVD45VuT3hBEWstRsHau//8GODi4/utlVYY
d9/ywd9a8uZ/o9D/blNJnIA8S1MCU31YddHoUKwnnzkEIutKI7MR+fHqsHcqBjoL
S8xlRwJAdLBf2f4T9MAX1a0ZmIRWo/8rqdCzLIpE0DCDfnpUVzqlD3RVQ2KioYoM
udAgUG23Cgfq7IP6XSXfvmDfqkqQUwlnxc9vIGZbG1qWkotkxxK1rsd8gGkwWAQF
fWBF88ITE5Xzoavjij6QKnzQGDJPNgUG7SX0e3hc/zvhQ6XnIrMJzIHExPxMFu07
1I5m32h2CK1dP1ozaTsM9xrNNN17u/bCkIAoFkkRjVQ4sF9peYpUM6e9dU0IrLU7
wnEAIf0NcNS5RVzo6Z1KleA8y8I15SGpTuIw8dzNr4vlcCVdpxSy+kN6TsFOddpD
PvJ9tSa0qtYv/fESsejrUCbO1o8oRzWK6EBVFIbBUXQFeE500iDZ4K5PozrPPK3m
RkbhOUDUjIJlShzy/5Chg/saLJqBcTppk3ZEFtNTTE81HvaxCYWJBNzBf64L+m+X
ZtvYps8NZ9XhnQum+mFDKMKfPXXQz7o65zigKVsIr54RsWPQeANwx8UF18MlyDwQ
g0mARZ6Qx1/yijzDF+b+Jr5k2M5iyWScos138KDxAYOlgo8C8Ig28dvvMrqUbBcz
1Uv5/GAXPUC0/CQj7MC9tuno1+Pbgc2lswjMkaMCt+V1knwICwrh1K6v/qkDSmaK
gpMzyr/jr14uQMAEqaudiDvWv/LjK9SaLtzql/inOePMWZk8tETZKgmsiqjBlpkn
eqI+xYTCpN2G2zb1qH+1ZDfkM26DxusiH9q1ANPEoTFEZ1kjQK+zpVA8cBrL+Ulr
4ciWrPpmnbGPMaHMAhrLdDcJoWhkFm1K8HdWEbc9cemMmy3gTRb/jG5CZKMrDQ7k
1FtuEFMMJFgb3yBZ0Z7JOwThGgodmtG65+gXyvCIuN/iZW1W280Gpq0E5zXwbQHZ
q27oc0StAnsnG3hNTnnUTvBFiI4MyNAPWonbFBiPxOlyThoaTLTNMlubgSnGIMWi
skaaJVBMIjpm2yM2/aEoJqM33TTHCXlSaY9Uq/KBYwb8bODtdcs/RPhRPj3HsUWb
rCu/YCur+1U+d47Stauv9MJqIi5n+tzZMk6XJL3qqaBeyygYwADFs/17HiVYPyTZ
iNj6z+uA5EjcMciznUCwbmxG6+9p6VVZ792HXMlmHhcVqKMLskgOzzN3GLV6NXoT
d8fqPzyGLKJCgX/4gK4m2vxwHsNLOdiOIivs38m+rHeueuy6s3Qugjndb+aKSsdG
aWBcXfcZuIJDoWxDihXU5TMATf2Ar+os7f7qR+x3ugsif4a/WYXHysF1kxjGmMSv
gQzdJPIp6O6nSfwVSn9HCS0kUb/P7ltbIE3ne88aPwewWVN5gGREFgG6B9yiEyJZ
zLGQv03Zz58oxqdJ/BeTw+O2tafJb/atLzQRWcRjkOOlNphlGbxqck3Ci+aPLAtj
YQjd2JVLj8nb0h8hRjaahRNIpGV6/KDl0FvnKOtNDqeULvsFyuFKEd0r76baPDV2
i2N40+JqRkrlxM341MGSmOM8sZ/RMF/ddD5q8xgTq1nD/rq0J8Bb7aEDIcy7VEJw
YxUohluGgq12q0fPeGTXPIc7t0keoaiRdtDjWHvr6anDzyVvQkZBOgRsEPdsvLk8
vfktycdfYlKOT5JaJ2xMZa37Ory8cECGdkBryzWP6vEK4EgJzdb/Igk/helRGWfn
hM7zNtX3dd5uwsSldqs7k5w9TIXORvUTL6RNK0X/ZBeXmf7fDf36hE+7PXy50ahJ
hrumpH8q7soFF7Mu0qo45gr0oKahKyNziXrzS9rD3YD/xmMtFYzCT9ikFRl1F17l
XRmPcoqnGJins7y9KNlKyfqAbx/IHOu7/SR0P7CRtARHmuznsCLpQx9sUxvgzByn
EdoNUFILPDpzHgAM+dY8SlymhQj67+iKPWpmjbSQJxdX+Dtv/bzwGLZa0UP3xtmY
iV25F1f6YsxUuSA9NU/zTJpdKevhintTt894NbH/hcC/6+zLSYmctpYG1TyySJFz
eJPYWMREzb0VXOYHOQUAD2nbanNdunmr4lWbgZSMvIjDn8bDvlrwj/cXWhdb305G
Sn156be0osJn7YXAPKjjuOAQHrhLWD8zlN5TROQvWzF1PDWKj9fGc+s0NB1p4n10
BhbrgMtn9dC/K4jOxT7c5xMxQOxQ9DTpcAS4Glechz9bZWhGzafKbeooYLJS3yGM
SvgZzLLWbjaHoCEbMS+X2GXFUlBmtJ7EFv9D1+rq3mAwO6vpRD1zYfzmo6Ou1NBM
YBC87pJdPwbIocXLtNgIu9okgjKxa4WvcdLIMHkjjvMIV3ieUMeeDtKoTatnyVKf
WuvcWqaW5AF3QJVzOrdZ6MOG9lKQiFuQg5I9J3dhnGvVBgicR/KjqZSyJVdjdKXc
Q/5IDkiKdZlHI1wmJQHYVMROesUvcVXcXVL7JP22dSCHK8SCjUcTklbKV40JViB7
t2sq0AbYv9r4iaXcm8QVkblH6TzIK+Bi09iwVnmwQyztuSg/jX4GtBP7kvIbmj4V
IJAJwCMw7QYJjtcDiLSs+Qj3WIyyQRCCgrATZyb+6djhGm2Yo5p8M9lsX1fegvQ3
EPT7kR6KBn4YI3eqDFOHszmqIhU/rdPZAtQ6j4h/4EHMjTHDIjlwhAFZ8RCUgnf1
HwEUVGd62JGYKwTA8fLWpk+fxaXN0dlqYmgwIywEplOaS0+SdFMsU24/6GZ/0WNe
F6leecADc/n2mhw1/D2brMTE6BNCk8B08D4Jxly+hqxHwjAsXFP0vK6oDOWM/Zw0
taGh0Sioql6hrvkFPC59nXxpcm8RJjNQV5FaIcYmf9+XOdf9G0VZ9b7N5n6eWKo1
QPKuBXvUplrFzbL9x8bgVhPF2ph+PU/2hSR9uhO2YLLNBTBq1iDXcmQUmpffDMnN
CfMG5HaF1SdAv/rP5fZArY7avHboJtYctxz2M8Ylm8uITVpj2Feqxbo9vOpHCW8C
yUMdxMnqeWen2VxPryY74i1hW7xF0mXHUdLq1SN2HgV8wgeLZDS6STdcl55ThZ6k
TJOp9BgTjsiQ6AT7BYQvddmwm2LMBlO/ucB14Ow3xIUf8RZGAHJdqipMNVfh/k1K
hKKz00xve3z5XnaBPPzoeEA6PR/tY5O7EN2lH4JhPrV3w13tDjD9/+C1XyTE2m/Y
THZ6dbW9e8NzuOpjpim70WXo0MykwtwJjJpJHgEjKVpBO7d3LH30gkbVwPqqlwAO
oWU/cBvW1n53kQf/zEV9i4Gnr7EqunKp+u9bx+brYQbRRFs2YBhQfZrCalvX34Um
cjD/h8SBD1EdtaSuN8Odr73r+rC/vMHqHqudVyHLyTgvcOpejsLBeRWOrXlBWs5b
IB/tGCPWRs0WfIrf0YPaJUGbU3J+ap9bsoZdUpdp5ABQ8qSM80Ww18p1R7ntPnEe
I2VkUObkgI9R0MkxKjeA69nqdztLJD05GtVAqCPZvGGHuyisBgpfPwWUUQf02LyN
V1bRN/eiafEiiYoD65AJy8MV9YiHtcrEIN1cOf1WgaqvHytvlC2dqDf7HMriALa8
YWylmEj9WQlWp6Z0ykkf4M/EjoTL6pFW3WZHRMLpnwtHA4C/lFnr1a3kFJss9XMc
rqn4QW1NGbOOf7b5QVNLLL3OmYQ5mSmZII1VDPfIPKnlRswM1LrGfCsF4zfrTK4p
VOuv7wEA5y4ef+HzhpipLonb10jWFBQ7XQD4RXd8xLdBvDNDpesI4BDUynSuQSuZ
rr+A2v2hcGIsiah7MUaG3DYtM9ZNB21mB4Pwet7pST1WAXfmeqtY7iHodGRaXcn7
a9C5lcFWYyoccYUbJb5kmu2hCHGgtSHoaishf0UfWSSzkJw7hvK0XNeVVVwzBfiD
JMCLr/58Ac7o4r/Erb3iRZ50AFNEKZ4FRy2aYjtsBhJV4Oe0B5q+HPg8V/ovjk/L
J01El9MWE52m05McfRSlfC0ygyf+s26w+rcFNTK3Y6z3lXf9Z4lUHKpjlJRfj599
lEu2y0/UyIX+5b0Wo87KLUKlFM3VX7HcaysqqcjWWYWqPubdQTadKTEOmdVw+s1r
39GY8vGtL9GcdPEIwL0k9pjnxvNFP1AhE4DJUfAKnFSus1fqja+h8ZCE9N93/hdD
YumoRviyS3WOY4iigfmOrYPTMsaMCZLMRtc6XKfLivmQdvAdQWwAJJdT3RBFO38n
p2iejPRBVd6DGWPzp1Bgg7wS+MhNBn0H8WWl1AUckScloDxQKiaSa8KdtvNG5uPs
RRyoZhv3uKh9+Le7bXoLLTNzXpCo3eyJBSH+SlgIV9JUjQ+yhd3SY4N15VrBzTXC
gaOxylOwym8ceyCvZgw/K828JPL/yw0jPEffHH+i5uIgi5d8D9tsOLkckHuL+Ist
8+/0oM9IyOoAdK/Z8GouBfQCRGK5NIL3GmnLXX6JOUPHofYsW8FkBolZKlrMqFOK
wWHCs5RtGyBbETbfBLCfwzaRgPqy9sBdgJqbG4pzrV/mApP6i3/b7ZaZ6C49TqFO
/mXYm1dWqnnY3fdXp31lvSTOfwDM9uAgz8MiihTOASguoT526lvneK3/1xqUzbFT
jZTTYlv9tH8zsqIMQKWq2Vo+JiIbmqxFzjcLHBnKMCSP2V/0Yb53ijf9M72CmYaK
qqy0dvzjj9GSxkvDLZgMCTPz7NfntjqWdvRaSwYARJypLWT6uRamFdMhBSg8HVXe
mq3YNLAV1cRw/yaSEe/jUXg7JVLeL2E7Rr4u8a3ZlFMw6OKl8iAosdr224gdRXxP
C2jL5mnwaGz9huXperNYut6h1H4bWxvUHSO2+FMWT18RJx2niQunze/r0kh3P5Ms
VNbDeMfKUb6rxH0Q1x10K3gEOjtezoGqjzzCYRqIJstNcDZdXmHRLh+v+RmVUXwE
nKK+54HrIvf7btsVQTy3Co+HTC8qnEmz2QEnJQZsLlDplkUNg/CwMbfEuO7723W3
kbqWMhp9jg0ADQtWXj+OtuFZ+X+7SbX2tZaSWzaz/RKKauU2OoB6DHbJ7CuwTXJ8
Wey4yR9tTCpxqBu1/Nx8Aem3Xz6RgeX31H6pfvN3RcRo9A2WlBd68YzL0ABh8zwL
cynQNhPJ2eCKY7hJQDGvUGoZPN+lNxGQiCS/092nkfrjWEwCg52R/zExy4CGbeKq
iioD/a1ReXM9oSFfL8doGGyO14kSnKxnpDPl0/dMTn9mVTHDRQ2PwtkN16Etagtt
aVIEYG/PFcTMlhYhmSDioICoIoaS/z1Xxe64OIUVeRm4OcU0AvcPG2rbVExsr7wK
Lwcu5M8aZpCN3cZF49f/zxhXvJyq751H+E37IrvFWMVUlWgCa4HwdXCQBc0yVIGq
fzO3pnE1jbAs0UZJb+AQUAHUeDG2bBzAMTrO8V/eMBs4b8CkFIiHwXm0pDJjWhUD
EhwRlXuYxFZmKCmtNHa8uHaswjwiGEBWSfICcPU1OU9hV2voBfGgTh7igAfBWs2c
VaV1/0mhI/XCJo3chrQcUXjuFd8HCvcmGQgS9ERDH1ojDy4BwEMGAAkTSY93mT/r
ufuY9WlhmBpUgOiK558/IkLckpKLBycVsLKocduMDLNZCdRhXRjbtEwukJjGXGwV
C0RoIZCYcvYv48plCM0qTyUozm+E94ulkVV2FBJjAhweig4TD3J1YWcCsG7+E//W
T56vo9qGnP8HDgovB98CHZpRx07Xxz/rdPNYdCG3McJe8QwTT/PD2+sUdhtuLlrx
nnRLrexVGjob8IdSym0NPptGco4dwQza99gwaQTXjLaYNqvmVZd62kTrPFnMv/cX
vDECAJyPnMKdacuWNR2fcP9ljeOXpW1QgHp2sA/zjZpqba+MR2UuvyUHvMV5zCFG
zbQ5PA8pa0KesUdsPPEVnizMP8u5NrxOqzqJkYxM3Es+/53h+XAlii2Gpt8l7wcV
kZirtZsmhhvATGCN9FR/CMnjtMxbyzFZTwnjQ+jFppI72PzzG0MeohScIvSETvpX
DFa2IFLuHHDjooCquOLz06WiJnCtAH1/udeCiXoHRC585W2zcV/7XKxanvIn/N/z
ElFtgU4YBtp/zAP7evczoLQYmFc2aiqX33WVy+8QgTuwzuZdf3gC1fjNdboFG3Cy
PnQi5QlNZlAzxC+PXha1arOQWFb9CX3g5YlUTMR8yyRmt4LHMZyUMYJoXLnIxR57
Oqzs9u4mVbk5PwgNV/Dv517NJ9pdpRUXkRVi2zr7ORrAm2W30AnRLQwyMjNuYBMy
jfFlcphbET7pJ6ekrPsFwvt14c5O7G0VN1Wd7QNoqc21eJsmer9A3is0BKbXUJzy
VnD4v/2Tuo3NuUhwwa5xUFlG9MQN0r2KZYdQ1lWguQ/X5b9REbp7DBgHFfiTvohh
b3r5iLwXwq/gotpcaefNo0XaqL/XnagvtnybwtEUjfLxxnma0J/B3HLeClQAdn6s
LguzOy3U4fVgfNoyKJPgqhdd2v4f5ttB1F3LZMUIqN/2YihoE/azEZG/0BmsZiEK
3ikSFHrM2+WPcoUVfJoelACK9PAiAfWHgllenOknaMnRCnx+hlsQ6JEmKq9CwkN2
laggKu0NC/1+yRyWzTFOR0qXpOMbPj0yfVUmGdJ55XLgNCCJA7HEBsNygpWVvd8P
TRIk6lTE2pnxwPl+C/rs2MvsS6fdMATj39DF1438+50FDSaOfOx1mrKCwAqihIxO
f82/cKg5btzO6HSAaRYp48964Xt1swxL9d2JRrNaj7eJfyamzXxTNYtbr9uVn+ol
Mu03K1rCMopHYJdzpP+GpCH84MvMPPJPkSOiOnPU2akfairQGRRmiJBrB63Jw9gg
pP8eCHYCxSZHr5gNrv6wtXqgs2ao7U2SDIOgag117Twg2xMv/FpSlN+70gMMNXPG
O1tOq4sTYoz1HX9ziLiYPLYD+SC5A279REKz0gEzdKp99hZho3OINeBpg9/37a5e
OqPxJ3vJzOO6DuWsCVoyT95/gSQsEkyYOkPqKqwkp8t24K7y5TBMltG35XQJPjpl
rjO+SI1SuyWH8EXCPH/nhnxXiN10wZofReaD8t9ByTZdle9VsfxBOSHobodVw2/6
iFKdP6J/GOfZmz05KODVrqrTOdIbWvWdtfK2FyLjIjhQ5vnIJUzs7QXAiD2sP6Jw
a+3kEzNxG8I7x4FP0thpUAJz5PtMnsQqglQJ4wMUqnxjlc1xOJXLmJCqiNxGguF2
7m89A+awXPkhCov4wCRPPWe8hQ4uEXqs5BTANShxkRmpX4ioZ9uVMGZO72BPGw7H
SyxcyGgt0xmy3uapNsBOXKZU+sS+0J/JWRebM2QBhfcK8gQh+75sPUaQ8eVtllXs
9aF2RNAtC7tl2UHWInNjwsXZ4+V+q51Mv3ZRd4xNTVhWWZhVVn4rIssI0IZFW3aA
IBYkKKv8cZ6GYQzJFnvVvBmNntejGGzCAFPOdiRl558Xuub/20BjPNGuKinW6k0o
lW8B3TD4DdCYmwnHOwABw2ncwU7qyYitnyDaS/aRu6Not1XrPyrAecSjaBs7rduK
ORXxHSZUUtx2nRXiUo5J0RQK9vgz0NLKy3PERtBFPdXXllCQcwsaMz8xXD9B8Lrh
gy2AgG/MfMVeK3HwCvLrBWXb2PyyLOQ+0cSEVGO1zxrW9chNkfkwbtweEdM5K0os
mvfZ1CyvxYKkgegapdNzLeE4vmwZcSP9V2GzAOxWK7+WHOiJER79vXrQagvhtXIL
zN9ciiRU9kWc1J6dOdV4Ck2PkomjHLrBxyORKECKd93GwfEaZendESFlElqYv/M3
myB8RkEIijlg7bISUOA+A3Knh5GKoRwqloM+L3V0H9XAXYfxZbJjZpN8Wu4zYvLg
NqdUbPPdmAWCL8srLqhde0GgBsLSSiCVpR2TR16RkNvwT91X5s2NyZXsBJAnKNXH
XxzCMknjcsVZpsf2yzQC/5iXADqGxIYjkR3yy9q9WiUaA01VU2xl2KTSjF2YFJB6
GCPlG4ifcDTNvCQbDXxRZYFDEixGfSXo6cYcC0P4C7RCg+N84LN3hXdDiMHn24ip
oVaPu8XqJFIePbnDYekW04xO5v7pBje1gxb4VAtRr8hNhUVD6+GP2Wq4SXgWYqXX
EKQoKgi2aHFuU/jxqr6qgFjGhNbcNBJMjQ+u6iWMbqx/G8n1rpBgwFAidxzsqY6E
rKU2PmuFk0EsrADEsn4bSdNqoEvcbzUqxlx84boyQmGR/UHRWrarbFhIAg2Yaxc8
Zf0AWWaJqC3z9FVhKnNYDFIfMxFWkrkrIol20mx2tfkImm8ZxucYP3AOZ50tJzqK
1FqKN8TReW41o/8Dx5UHG8PG2Qn8PZmuxAFvCsLDAJX5s/tQgkI9VyYCTyXVWsjp
rJH8l8dLUuN4OLUqCADPLVEsiVkfG9Nn5+S9mzM7Sj29I4KWJg9DcOiAdcHHmUNl
pmaILJ3cobsjHYjq9VZCPKLp6N9G9Aksjl9SOpxZjt8drl2kowk/i/7c7aZvnm8f
+bVTgj78BUKvy+kokd5VlnPoHVTS6WcHsjcB6bctAd+3dN82u/vQ1V4JIgGwgVoG
BkekGrGQEEoEoYbfFBgpFLOS1djmBr6cPsQmNmoijqkAlkrGAocp3LRtTVQFBewT
fpUzk7Q9x65FDB/Lkhq+e0+KcILSzE+VVY+PTWA13mY3TxUnLNPvrQP/MPdlZCkV
LFFcViHYoEG90SLpCYmg7h7NscBhZekOSE9Ys7Teu9tNMiVFYz+ifgd3DnURXnmy
OO1ijr8K3NHUUzoeEnar2/dl1d9ouRvrFwz67jnPDwMh2J16o7z013A/tHxZeX1e
2DCBEvJb5O8wtgt6U7YhGfP+CsiMnS+j82VmeuAnkb6fVrCq+dnj1lilAsnDDFcc
35TcayjGvRRZ+yg7zQANFg8AQV2lLAxJWL4mbiy8uSo+AISVQRfFhh7ejet882sW
YsRmTcD+wMs3LAoXqofwMS2tTKBA9994BGFLDhC777W0H+lmiYDjLsneMALGSF4H
NeJxGZ+B1RpDpORQw22R1xHwkORmXIycjP98NclH2NBqrcH3ZCgLeJDDX64Lpmet
M3TPluznJGNzo2CUE4zomBrvW+ROcqgaL2zgl93V6P+ssRbuOYVqqBTjcwMLBoPO
wkCPJL3ZMNJRWYE65UY2C/Dok3KnohnaYjfJKZ6z209p8uuETfvJPUhrSvJRwiCz
36LJQQtUB8PUIKlGW7NX6Zr17WOsbfi4kZjIhqoYgqgn2ggiv5+GosVAMawGZrdB
dq/+xVsaem+I5kK//r3gs10D32HyLNZ6vq3RBtT5wbfv+MAirBMfxsFstnvVxjyZ
lhEkKjGEp1ihrePx371I+/S8DAVVKj+od7uts3Bnp50TrZ+XsmJG5l71REyv+5BP
za16O5d8ka+FRmnv5ahezW5kHMyqTpvApON8RbiV002TJ7qOnRhet9ogFOV6Z+8Z
NfmY6EhqylwVe6RGXlxoS+Ra8KR5l8MiZPkUIodIt9c8X9hqBhbTBD5TA7Pe7lgF
9FBkmaG8QjgAqlkyboB0Ifr39MHP3VFSW5vJJBUwHAYV86chCt4qM/SjbK4cUeLU
qB9Vo4KHhhpaCKc1zJbEH1PO/sWPoKFYV/HY3GJg7GdMqKkDjP8I7I9nAOoKeErr
DaYAzRTfrljc/Xlx5rYpzGu3ycXDDCaTABkBjJ+0PmWdt9yAkvJ9o4UU7Ti3BiJl
4wg5fnxNScC2gHSmM850wNEj8TifS4NFBaP9Z+x3NDorW7nrtpLd1zzagYno/5x7
3loHiASnEZjyW3g5mk8StHG98P9K/m952vjZqiMnEyep8psn0QLc2EXsPpKbHPRz
IRQs3bLr1xYMoBq3dLFwK3o1CMrSlJpBep6UMjB72DLOjh0yFvZcSNzlQVKr7Hcg
TScJXgkD9T5oMHwJk+t+nihoSWoS3I7Q0PAdP47t9n7O9ZiSsI0eyDnwl/a7Kb4M
qqS5t/SZ/BKR+/WjucAxP40tW+lBfYaEjEs4N01wr72hCvECdDgVHJOLEMlfssz0
NxyoGyJr2taiKiQ/qlT1pKq1N9UDBK1/4RSJdv3QuvdKDmA8YHxReD+yLu+qQbJU
FPgJJ14qquzVhEtTmWFAIxXzFXPeTqFouApsDVe+g2i/ellGiNIsd//jWTKtHHlH
Z8eVWVZ+x6kquYQ6S00evVdnIwp4rcZYzct3K+YLCEQU5hQUG5ItKWbyzayPa68n
nfpgW/mHVP5/4AQ3EO0InWRlg1WcpQFlINezNHjZx/jolUntT9Ig0/3Tv2a4RpzM
TlVsvlBkCYntJk8DsnRKseBQ0NYs69l8QVvuwcpQXOQrxCPyM2BJvZqpWQ+y+4oI
WKt//HwmRAZVFJ7TpvIpkLJBpcfRdsWjDneig3q+SwEEUuQIa2cx7s96pk4AQbds
AIn3UYB3OLwmqmFG9dgjcDpJ0GLrse/Q1BNPnGyiWH7mEMMBsuMtTx8KrUSnX2p1
VnE0SUvOC2HM09NPKWtgm+3+DtRkPBw6s2nlvOXYWVqCzCkJbmvJuRfpmCIJZHPo
oOJp4M8Nmh7wwrP9sIBSatgPddIYxipudjLqzyatufVI8koAPe8iaygGHw4rdbDq
6FQk7i7j1nFxB6nG6p88P3cgPwzkoqCDVQ+Y961P4SFwx/2azHzjRpjYVEVuM0Yu
wAXtISmA4qIfL9fQuR4EvMeS6FoQ4l5j/4DQTqcX43EYQSSmeuVMLVHxwR9ornha
tMdqFFlrpsJGQOojHSH2ENGWPogrZeqNl66ONBwyyBe8WL5/WZdQrGPbdV1zQmr5
mFrPDL15bTnJZvkfw3Oi5adrVkI1AePbChB+RMgBHLbHqNP5J/qmyv6oWk0H38+a
h/ZUZHRhVl2ZGorJ4jL2rWo2E5yBgtnVrSG52iGl59/h/DcLm+dc0jNAoddN3eaK
Qj94mzvjaBpRJW0E9k6P9XYC7XcJGNXEdJXJgZWdDn8gpm//hi2lx9aR4lAT/emr
8Br+89/UEQv5lSJ/VDpmYyY0n4VwPSu+JcBroT7bNBX/fwkFYLOMSNrdbLmsy431
Gx38JJnrOATAntJRiLSjoZ9VCaIhMMAUchZd7kp2nbWOPvHW+IEtsIx6B6luNUp/
JA4PxIAWR4C27Fj9p+PXarURv3LDlRzGpjQZIQAmV2+b21S7lF3HnJ9Xd81dByb2
MxJiQFFVDrD8b7t8EMb/zTpLkZnskQX9sHXyPxB2WuPJ3tdXVp/2+KcPzOU5PChz
5hJGwF163ciMixAbxbf9nwhSY5X6nwv8+rrRbHWUADmaGaERiy/3trUOjScWCmYH
Oi9VQpabMr5isnzDgaXbasWQKzguGGhVxuNh7ipHLgCMdqsWg4em0P3TFe54+iPv
09D6fKmJuwpSwazLk+ulNTZB+kTmJnBZPbvQGkxYUF5UrSElYMhHQ+vaYdSwGyQx
i0gr2E8Zsfs8QDTVk/5NVjIIXHPog+0N0S97blFPK7S/1LSatGmeK541tBzwk8QX
wFz5RDLCNGUR9uRC5RmXhsqdbFWRU+OI5m/OiG/dR7UhhtGuk5X+65NO1zu/siG0
08sDQ61gw1Osfr1sqx6FgR2ZoNQxEVbnZG5IEWBLgXcy+f1FEGHnw2Xg4BhaNI5n
NvFPohg9nHRzJCMH6brbKqX9EkEk+MFzwyj0GJW7DJrlEzJk8mSIt2Ww8cd9v5UZ
NQCUOe7oXhZHq5AZX0Jvg0nhcqK9HNou755Dmw94V5krQS56enm3O9LFSsutNUYB
093DMMhxEPUl1+OB7MZPXXp2W1/Xibpw/9slERgQSVzLbm14QdgXSx4oY4eIAl0K
J5X87DqTSBFQv07rW8Ld+gXrAU01nuRvt3PfltNzOY9cMgc/c2j4FTDE2ncbOb4c
FrsHuf2lmwmSaGuoK9iyae+DAPGk7oXg4v1WRfRU9dOtAo3TKqrNoxVNSpVFvQpZ
1QAYUmTZ+kCBjsk0Mh+qF6htDc36u5wIOgEHJ+v+wa8wNZnnWGw1jgRBNDWeAowN
LLd4HxwUlcClFXGYPBVLcXelO1eyBNw84eR5VifmteXfe2Vbyx2g+4FzuZT+Gjy0
7X4gu9NC7C3I3czWUkFN80gnUaI5qjAAq0KBEJDmQ0+ERifvzLXstd5RqEempTof
eAAUYHoYg2HRBqQI8GRVCE93+Gw1J0iIKph/XhfF5vT+vogpWRvpya2wN4rMRQsn
fC5sxDKR94LVTVofa8fqOZM0khl2F1o9XdCHmM+6wSqP3xAk5YvgGmQyGXwsns5z
OTbUQyweXilQfwsoLHQN1UXLHo/yIt/mn59Wn3hJUTXkB6kW5F/DX/q5GqH7TSJj
GgzHGlBmO/w4Ozfnfnh0R495RYo74Z3LYype5SY1ylSmpMwcgOjP1R7rxPgR13r/
6ihbQfNKDCHbn0BXQcBLW0gLF6abW93ckBHxcQ6Eb98XA/1/N6uDOy9TeT2JNwll
ZAJvwrwIfDARCqmKBsH/zB11XAqRgOCp3ReEVHWD+KR6yJ6seNZdAn/duWA5F+/K
psvo5cgvf88r9H2FRjBf+0pU+Q9u/XqZo4vvmYBG5xIizsg0XF3GELL+QaF4RxgH
5FR6HxAdBMyeQgmCGUZFVHCrxoG+PKfjIojhgfNBfudj8zJKFeDoBw7R9AXggNUg
ttxVXTsvVfgEMO3czr7RQGV5U1x/yXSC3VCInGhE8IdGGOtsZj32QuRbeiIM6rpH
j3bJ8DSbEso5m6SnG50/idMIGhtxnJu82XYJBGTaQDjSfU/AQXiUSgPybHnujWkX
PjUmxuHXdRtL55FYFpNaK3JY/krSEv1b6zUi0PRtE5lJ1K4NnA6bD6nqq+fjZtqw
dR0hnTG9nLU3wxTL8Wp07c/NAMcGV05klsE6rzkTX5JnOh1mh1D7WCBfaWJJmyoJ
36mV8CBsMj8UIibtzNpqC0TQGYMmWMhLSL1YU16M9byOg7Gz/KUhiw36I22HhRGC
nbxfl04XPDnEoKYx9ooOIbM9Ekk/1Mz2oOx/+dO3EMPQWnrN+2SjvFC7/p5KpX4C
13Xv+TPPXL0Bpbo5YlmS/IjdAYgaOfnM+HZsBmoltTdsSmHODeIRyrEcVTNAEjSJ
3kHcqDx9IllhR36XebNW39HR+ZX17Hr0QbU6p4BdFR6fZIlrMIRzhEAO+lYphuwm
TUJcWZmhm/3veuqLRVOVDHqPM2vHWtnEYLibKaROtVDqS0WQht4e77SEuqXO0xx0
tE/JYI8VvlLFpMjnijqz00o6/FUBkobOskka52+MUBqFUxmZJcIyqzMR+yfBWOY4
02meOMuwjtXJkTp6UYKoHorDC5YBDfn7UGqf5HenLglTufwvVLRwswY2rKjGGfoF
joKav5UNIPkNYyupluRtkFCbMvxr6gagUoRmj/4Muh7RU6+Zz9wue1kiFz/XSw3j
AhhGYdFyntD6URBOyv7gvjLkqOdsz/m3dRaLP76SfzdEZqvAl8l7KXHcvbuE3qJh
3s4XgTvx8sJBezp6C7TwIpuSUnse87NFGy0lYcbF/RfyOvFO4jNHmUQClhASbVPE
XZsktvlqeqi4kKCmp71l8fJs01Q+xlLurSdwLBJ9qnPMiHi0FtlvYqtdFicKts2G
ZxKGTdsMUSMIX1hHJW7+iGtNmx7IPrNoNWGt83pBh1ReA8RiocVyWZ1uc0yL46W/
gW2mRMTmjYL8l8sgp7PXv8//j4t0jDONFHY92NWMtz4tBLF1Vw02bgUL+mvAeQ3O
OhVpz4hpJzYDx3c/mseGBNETbRHXmCnzS+KhX69ZIlIVZ9LGv7dg9erO1a2VPX4L
SDiYe7VzT1hdyHaM+UgtACbHcyyKKDUx+G3KT9qq4e3M10U87Nqt/FpAY713RWZ7
dTpvWcXA0t9xdBkPB7y3gtUAtCwBGjP40MaABCPLeYmRMs7weSjUeuTrr9Z3L5kn
cbeQd1bfl328t6OfGC7kUAcV2HH4zUwOuQlQ03+5KZQhqnrapZGh7eEfWThmh7UF
QsH23bkWl1qHzCOxvIlL/uEXW7F2DczZdek/oBvS9pNdwbiYYysJ6lrfPQ2v04DP
MzXPSbS20TuMl48zIGyquQgJR66+PCJK+7kPmNqE0q8Mv6YPtSS2igxK6UJaa3eU
Lac0x0H4bOiVDfmwG91h4w54lkfvQy7H6Qsws65PB2zhAhO09akwiHJXEFUCaicM
ogTgvwQEqjkyQQj80qnwAn70AMUAbAoyfsfNx4GJYXxlumcJQNIrQye3Y4ugfU9M
zmsCeKYISEY+59Y3hsjjyNa+GhmADV7QTwp0lXGlVqJZN5Q6DaGzdcd1xzPEob4B
j2ecT+cSLf5snfkegtmV1Nd5xihdu+ybYvy4WkaRBQwP6AHb4rxJjQTlGCZE70Vw
/yLzFSifCVTrMX2aUE+7tWM+BLkfJcueSsmexwpkDNUuMHnhzR2NfO2XvcSPbI6h
zGoJdjP/5L1kWERusxW0JgggI+ASVMV1uGzhJzl+B9Oc2t8JkL6bikuG0DqkIuoV
nRrHTq9ady/t54aR0zCRs81HWXMw93FEN0md4xIAG6/Oy3CSbr15GTstufHBMz+a
pw4BJrbThPf04vUfGAN3Sm2e5s1htlhpYYw7+9UWg0OYN1Q4IxreS8bj48IT2h8J
Qmf9MkRdjW1NfIRBxRO8iFwL2zaIX6kgylqRbWcfjlPTtIREiXubY/u8U7XThP4x
4X+3PNteL0I7T+3lZey5cpFkTmx6ldyYgE9iOckH2WlIkg5VFKovas2kDtCqRH6r
CYGG+NnEcS4dAI4uzZWkUE7tY9g4tvNZ+Nl+ORJn1FowJHCcTvJsujeBmyszgeNL
L+W5v5RnbV1kFi+6LQkd/rhHmO8VDQRm3mhGLclMgqC5B7lh917MuYKf3mk7qiBz
D9sRb7/gTwOBi7c8UmAB251iar7PEOnQXT0IWADS0jUxJMKD7j9+Uba1WcEleFjF
QTJoQV5n5w4f/I+UkrCW6EpUat8cpGZqoIOtvUU9x5wj2Qms7M5SxcwlVf7LKkDF
VEJ9+mHzfQ296yaq2fc8VOWy5ylutjlgj3GFEhEKZ+mpMcuoaIBVRqfUqLI/hXYB
0ShxZ4NHaMyPCVeBwBVkboVNjl0Bi44ZhfghXQJ4In8Bc8V3yZaUmj9GIH5v5qJD
RtKNA0VyxtW6dWtEPX5i4inYJ4zqI7ljirMgOA9yOk4yu7MHG94mL2dTgwRP9ia7
rwFqNE4aCZuD+eFONXyj0wQTjr3dOl8nCu5nGL/+3987GBLRxQk5I6In9AHMDo7u
9MUViyKX8q0DFb367hgF8t+/S6WxMqpjFnoYvbnFtwPYoSamLsulB+S+SAo0uAMJ
ut6xko4Ju4b4SRMISs2KeXF584GCeQVlnB+F6drJrZzs0J14c/ZMtwAB9WZSy1bI
/LbTmzh30Sg81X7+nugAaRbUVXQiqyBGUQWEGdJVT12L1XdK86PKM4xVrRkAVVpY
9EOxEhK/7fwErqVdKO4erwrV2UgPTt2oJyDhBhiRwRHlNpyG7VsvJ3L5LikNmWIX
5BnBWsNltvMFuW2DRQLy0pXkF+xfgjTZufbgU0Ety/ZsjVKoGFwcKaBjpDWNAsCx
qA5YkbZ/nX+yjapYod8rE4mLZWVwN7xZ80TWqdTtZ7bdcyWi5ysDOOXLcFV5meY5
1oMdoT0ug6wO+1OGcYBl9MBFk2fm50aeZ83xYw8B+qeFFEACsOwERx7NRA1BTVdo
O8TqWAxUXnVOr4eV4u2crsuJpexPpcJPAtZwI3ud3v1tsgwFWQRJniMtG46j7+eU
IpiBsWmW8D0YTxi++cU1D/JNSsW/R/DyNu2alP9DjY1a7m+03QVcCD5CNvb5a5jw
dEVAYwLD2uwhI+d83iMbozXc4uF5kGEhBRBWs7XNQlYNxki/8Az+ngG1SBH2iLQK
97g6tj+A6e1Zc9C4gBiJ2i4omlgd4OZljxUR37UTA1bjpL/qImKA4ztU9w61wdUm
Nx6fcBIk9ppZIVw7JQC6YTKkTzKtMzSAFjalTzvEp8pb8WytbAb2q1y8YQsPSv86
gazuLlGABQhmSrg4VpLyW5sSUms+DYyJDL5ZvvlyYKy3o7QK51WcfKxeI7UQ6jwA
I7YyGV1t72rkLhK8XmfEODTMUzcQn5+llv4bWW3D7Y4Evaa1gLuw9R8FbzoPt+f+
/z3U44l/WGIf4gNEVbRSfeG0diN86o6b0tyLNCs9tTTMZ5LaDp5rw0x3SApPDZJd
OYOKp+4+4qI8IrVeZvUkXSJcbn8RVrm3TFLe2gMVDt44+cyzU09ILLyej7LKhDrI
+11wmBksW57GhR30be53Zn3o4w3W13aWDd/ujiCE2/Di4HZgHuh9wf+AGbNoWJki
V5NG3Xpt5SCsqj3NCZP8h9doCr9wT2xgs/XjC8rlQQHAUbUfYRZRvOop6BXb8mHn
QA/ttgr/tRtYO0ssziAM5cdW6K6NlCIA6bcUhRTvY/HVuF7TaOSt8AguEW9R6DtO
Ap1r+ZGjOT3SzeLCCyLr0RQfNC88XiUs5CzSae9pw2Xg7iz/6ghIXwmW5qwGZjS2
PPOR4kPBuv/UEvTssykc4OLe4ry4Sp7zp1pKVIQhfo0E7Uz39ImBeK6ylkMlLRGs
WugDAXpzkeIcYCYmhYbsfxL3CsnmmF1NMDrSvJilI3zcmMw+sHU7Iqe3bFatl8Ma
MoI49BGE2SnxEqCaw6xqoPMIx0omYFf8sqGM98XfVauqutC0BPqjfl5ICvoGMjru
zkj45G2Zhu8+q0qc0Sei8kZJn+IpxrbZ+XjEFP1EZmD+K1TyE/yGMDcXppMPNgNC
4oZW/johJp5FJAAq8HSSkv8KJJeSebc2L7w3bqQkFTjwiyo96QQWhk6NVfj1tpKP
NvwEYYYCOwTzCDv6oFPMysmgYkUU6mTd5VTSHa/N0r+J2+uKJ5/omHiXAYFyqh7b
e+pfxJ5/aA/euRthwAx3+SYlcvRpQ/y93UfPfWJU5nAVstSpI0C2u2NCcltXfvxp
62dmH8+eKIu6eE01KVxYO6MgHxB9M3lFCeezJGSJ0WobKFcijN3mMcaGtj/4sEsV
5Bd4NVQT5BE+DePuth7MkcQbth+5Iv9os13HY0xJ0SEOyn+oOEWynKev7geiayjf
sslCaSfXWhJ0QXxXo2rfmgUUH03ZqQ1THk6o9tkxs4RyztwRYNt7h+4hgHmszd3G
lMDCTdj6x6676zCuOPk8lyp3+tzRmL21fqIxxzdMsO9fJjAaiuYgQBoIXpm7zZlB
zD5e2kbS28OGcfFtpXbPoQJyUZRhzh/Su9BuvC+oZ1qLJT3Kz55rnCBjP+BAEHQ6
kDwl6VEK9nYJnaH3tcJ+fmEXe/pOJcngS5dy3Bpsvi8iKmFPDj6/eCvsUK6zsFHn
rTcbYvLDA52MsvNAKmaIjbR9X+CrQqX7fz4feQTclmcSDqplpOm3lCb3q22PEcBd
BEalb/Ej/d7E/9PssVUylq7/w2yXhZdwhHl5D46WCmVeNELPY7338ST1StL2XEXQ
mNm4+kAN4BryWL1DuICerSmWQtYNyWR/oJBUn6a3ro//KG/YGkZdUGydOVn2DFWb
iaBFq5g6DC1grbERObBjAGBhTCTPTFlV+0lZZZMDoh3cdYE2DAEZMk6d9bZlUPma
DAlHJI5jsyshXP7sXbhHtonLZbRt8CKY6Kx4z/hSeNBY1/Qw/OyQjitPCFPdv3EE
APjOLMayRBCJiqpjZPLwBpyc/FchGoVkCEFKxWKbQJq5RnMEYKz0+DBP09BiVI2I
xMYgUNreVyper7Fowz+7JKfBWQrjD1LwnMxpIdrMa8Ag8BgKoaalOlHXR9hjmDbc
U3FKLyK7mOXJCWsh9zmS5GJoxPMlFrcjzQXXTmE7Sziyk4e2CZHVNs9nho3CBlHW
dGLGnTESJKz/5cpRcoMJwCl3hWFHrKdWIy1PmmnncoffzKoKZhSwerxcGKwA3Ya5
aTMLtPt3E9qFkmckDhIft8SEpy/0PxFU66GSh/WJ5kK7PvvY9n+w8wCPeFRZWnOB
YPVRdYKkTAJL0JyMkCeZDaNifV3hifrpxTIEZhSNtHaQcMHxKFvupNApJEHTk5dl
A3W+WqMoMGPqhgMxZyZ+2SF3ouzy4vW7Xgj6Qa2RincsDG8cUp3bi5egf5zn4atQ
IjYlIH6kDz0iLqMKpuc1ZjOt5XQbZzjN0yw0WZ9OwoGDYffYfu1M9xjuAkkHhghy
Xu2eFDnaKYaTdbZwfoL+UNZF/RpwrRrdZgw8oKlisHDkPTDMZ6G6IbEGpaH3zpNI
tVYLE9SJqPcPekQQsY9JNXFyjUVNP/nWyZGhvaPjbNhwUZqnpyUx45krzM1SuGKt
S17KIIaavUP1a2/cfzzjw4kVAKfAB7EcASg0eXBgGJ56HOT17OYC0XSjeNq/4UJt
ZUek6lhMHutRy6pz4Z+9R2Jze/DmyaJaKDHn3nOLFyHfSsLTVH+UrDjcbqb4Uwu8
knG7Ko0FcjQX5TUOoU4k8v5pnHetuDV/F+GmWHPzT1V2stGttQNR7FXSCPXNnn6L
o0dHKqnADjOxF3QzrKnMGlVN0OF1+BFCnsr9CIxBiBSjnVcjRNmwCUqcZJwCm9Mj
IDIkgQXzbJDxLurbtIAzYvfHYM6az2TQCRyvzWgHBD0linK1CuLKz7VQ4+kz1E0O
c5KmWkN41N66+ZS2WFpj/S97CnuKa5V6ZpLLgs87+EyiLa9iKxhp2FHAqwEceA0v
fQ+HLCf4g0ceRaW27K2YqvTpAJgCd712qYrpNO93+d5UUrreIaRWiDHZ7m4m1fKa
Kru+HfdU0Zwl+0V7cy/P8Y3njXBzNxrwzIsbzbC5rgKPTM31kvzgamP6m4YNHzw3
Haydh4s5HFbO8wuwz6PUC54IGntp30TCjZlwLiluWRpiNVK5VGjs6Tv5/sYfQDVl
00e4WwOQ/xROmGw2J8Aj7ya+fc6KrTyTH+F389lWlMU6UsrqFl1fk/kgYghl0eVM
TS0HGaLjYc8nSiArTfB0n1mryRIOXZpSHVarFF7koDohB43stE09FQhbSf/zUIG9
wZA+s/CaYWAra6aHz8vl8D+opwwUFBZ1u4CxpVdCh40AhDu5JoHeExY40XwMmbec
76+EfQX+W60iLAqYKsk5LX3rpuuiwr6OPNKI7w8mnQPd4URDPRrA9pfaSCm0to4t
N7G8Ea25NRvvhFrdLm5gX15SySmwSVE+xff8Ex65taCT9yhAn/4w5A4+1uZMaMxo
W/nPgdZAETnBfNfVDAI+Hr3nMZRJu7WwdCOCF1PPTZcj4hkAS0h0C7vG/rwSnjF+
mkFcZq5t3EZi21KIghKLcD0bKnOMPpOkZgY8bPLzShGYNcKAdVYvJ+oF15P2e5cG
KGyUVgJ+rPb+xavUbAfyyX9FaGi7yJzfDgnb1ERjBnkse1Zrqs8DvXYLI7QXSLsh
4ua2tyEMl6MFGY3FpcK/q41EMBvu5oPzZP0fEu+aNotecrYVKWjMUnLlBqVeATbC
rvYH+5L6l0TLnWhou+j5jbMVrjkICjmi4581BHLvmQYtu/7j4YjlN1ZUqyhhieP6
rBFOva688FxWGz0hCLQbFg0wC7hkZSbaAF++WKahQU990V8nG1UN6lLJeXKas3iv
8I3Is+rFjQz5cojhaPit45VYbhTsKJ/metfGSLIISkQvB3cohdzkuPsDg1bggBuI
Kd5bApYJ34dFheqRhZQMTQzUMtVy4SiC+gOSJZoUK+3SnALAufS1V0/GMCbn9mtF
qmvAE/kdTU5TyOVNJjbFS4JrQGFQaa3WyBWD8Mc9NgDc4PhvyHPCdTutvC8/oapU
xAsWRcXO2Nxh0VlT1GRoGhJs5mYAtxYnmf+Oq0i9eN3ewmFvmAGuUT+hhF3YSQQR
w61hF/1sB5CJ0Rvcchsqm2QoFU23Fpk8QiFrmcq2pf7OHPOo1+pvGmjB1Lk/iyuR
2ppRyXoutLmyZYgruB/jCvqSgy0F5BSu5orlNEkytOJcZAdLKB2BJGURlDKlD76B
9TfIOvX0wxddVFWRnINljbMCpOXbn5b89HgQbx+wh73Afl9x22Giv86iJZ2/l3YE
Ur+lyT4BpaDOUuT6o0sP3ykgj43fwPtGQmbmvezZ7+/Yzy3Y2cO2igYwCTAo3Wed
vAJnAsJhMkz/v2pZ7yS4XNzs02LVoBefroOJ4sez2O+WiRZPhM6LDjU270PW99Ea
YPmjOhkC391n8wTXGVxw14zgrp87pq2wGfmRis/t14LL1ceGst8hou4wz2nsOuKO
cbwiLzkduSFIWz9/N22SVgvdJqxo8SPJNl55tTtWog1an0N70BuEk5r7xuXQ1j1R
pP0BfB/itg1eF98VM6hmlMJBUGprBK2SI13N8WTDW+yNtgYf0FvR4fQ3MkkQVxoE
mZLS7LMisbiN5yDYv6oF8pvj4LZCWdz6vXvwSThkPZeEZvsL25pYgXBHlGhptSV/
ttl6qbOmiR52KxTN308YO0i2FuJoDQt3JeDBPLbuMhbE9a+h3P0nm7KviZS6X637
vyl752KzN+UF5AkBO3VX4eQMx8w0YpJ5A6l1qzJ44uJYnvNt3M1t3oscxLQNd+fW
gxHmg0M+0Uh1dedzyeRNuT/6Zgfndl2iNaErWuW1zX36MAOPzoL1QQOkyfFp+12S
WVfJma5iWEcHf4I+bgSVFFRu5JV/cZmAE629p4LoRHMxnX0sV2ihJy/rb/GSB/FL
2J4yO+9KiXjSnMBOnO5hip6qzJhzdIPc4UjydphkHnGOOqRNALfwwJZN7JB5cxZt
/d0DwCowkEz8O/RUPAk3FdsVj2/Uc3ou0B6DiE5MUeAgdd0xS+Pmss2Jyu8WNJ0A
F9jyMOEvk5m+Qg2JIfMQVPAbaU2hEZaCn8wo+hOCRkMNWwBiSCXn+oYKsDvSLfds
Ai6Jg/emd7gThB+fH5wuOjRdM9YGIUojQvA4fBSmcMhF61kjj2RUWwNk5dEtuSg/
vdI3Ub54dQKmvTabd6I5IsWunW0XIsoQ08vXiAOcNHoOXGmTLExBdF1k8Q6N6DeD
/5c5Y8VblOGSzf+etXsCb2AdRldkjxUAoX2YkOjSeH6R8iv2awjBV9pOVG5I12eH
opcHAlqFnVLOX5DCuOxwZbXpkPbC+pj00vV55xpDng+5Jo+CQC3Gj2MA3y23GBA+
pfQ1b9pYeuBwj5FGBhe3DyYwWJEqo5ghfwQjwXU1rcc5lOXF1400N1sQ2J6gJLIj
FgzlijljXtW+LKmcgNDE2C/U91KXyshSv/vTwyyeHze2j4u90hWnC0gXQSCyM+rA
PLDl3cCrHRp+hK0tNTkiIeXD3B40cV1NvaR6HXiRLnbBpmNSy74Vbf8bYCse2f08
G3fqjGd0vKVkTYmSPGMB39xB98TG0t3HR9O2GFScpomueUH1cTLoDK3G6P6p6BvA
S4T34i8x/ORNQYuucn+7NtrUOSROkECU8tK8iBZKLBd8BEFA9I8kCnN9EKprbPyY
gvGDs/YMVBLxDf5fbUp7ImOPL3Z86weiba0kh2ehBeYMCUcGIga0BF1xeWOU5Apq
933kSndWUCJk7rexwwFRKQ2CkQRVa//QzEzPSows1Taxwb/P4BQ7ADiFT6pW8nmQ
/xHkyU9biHQ557sJ09MxMa5d9ZMxujfzUS9MUqq8xLokPGqtENdHBXDp+wSo5oyP
P+Bp1HWx4aFh2eSaZVf46/2206nF8Fa6yT/pNcppClhgj7h16oqeA/zpbuQZCC6f
tQjQ2/VED0+up2i2Jq4XF7FF7HPpUx+xA+udwE9JKHP7+spgvayXdzVmx3PGqKFc
HVxUZnXWnszHLpr02Wvr6kPa091p0YbNLwz30nnrchaazhiTt+CyW/2YOLUOUo+1
NbZPCFAEHV/pbOPmVbGF54ghfAN4hGcfPLXtVcsGosf+MLLr0YpGvVx1KzM3vWsc
NdKLBDqB4v2WqC8bK55gx7wBnR9HnbgyvbAjxJeSAaD9es2y2LDp0/A8xChgW56Y
bDXFkZ4pf9QxdPObiLeX5NdanGfdbhFlOjya0seFCNZFYOZCZkGlASYveUOKtYbs
HnRYA0qmYEg1yP+Y0ZuEiHVtpjPPCS6M4AYYbXh15IeqSqt2cWFrxzICGfpVIq7F
AjWqAVYfmALgkW0Rr3JJHq0trXQqP0sZrFRi7Luzq7zOq+L5vYFOitYHDGJm5ckH
pG1LmpPjujtzmNnKVrzbJvfABzcbPmSe2wETbs5APhoIBRq0gPwFnmYhSXf8Y+qc
MgZC6l6klNswfoEHRrSCwmzo+2eZqCvAuUhJ7b2FMXzS5wm9qylOCUz6g2zoueoq
e2YETk/4BAw7h/fYOqTGdSbZafL9xTKA5KsG7wIYQrsmIZRjeUd+3g+uqyMn5R/J
69hZK9c8JtjKcdrYj76zmbPvpMRGBQw40k+CphA9PMZIttrxlDlcRZoeemV65WvK
iMSb0oJEgKF7szDks+VTZMEUOO+WGSsdiuX6uYPO22qHQk38QINedkDQ96ubfOSE
SrpvrzcCIHJlICMPr7ZTC8uVg05POS6ii/EdeJY075M3wWKs2jC6ZxERNwZXWaLB
UUFl3IZrCqUJ0ugvLZPxSF2KS4+FMecRuDXVmXknbnqx2V5aIbndf3JLZnoQ8qCB
W4qDTOvv/WHDZNASfa6MDB4Abs+acW5ycL2MWiW5klRJRJC7qiHyuP1caNkFF6DY
H22kIpsbZFBMxuk9ukNPGmAaBG1vn8NDPuXk8pe+pikYodXm3H/yBG/xCBzC56Gx
3lbRHX6o6kSjfEz5G3phc0USEQKYt/E6u0C+BUckyZNZ0yqPDSpCzkhS2Uh2JLdf
DYGEatVOJzIPTMlGnJ8tPHtW45FtupEYhMuBLveus9IoZNF0KnWm6hbtimkD12jt
S7kdtYeWjzVoXaWQsAdGpY0NzvfNUAmmGi4h8M4gbvu323w5VZW+PS+iM/rMw9AH
Aj4AkhO9FiZ4vmN9aUD2WnY749eLA7a2WtF1NGHWfIqslwG7IxkaQvWwCDRAn1f7
yoC5MdtI0VBsXxzQX2KlgbqYOkBWB427QSseOLf/LgwqBn6Lz3EUsof6MYTG4EsT
9AbZ8apSTrUT36NGuEaMsFmgLxF69Agzfe3XuiQ5+cctAEpp5pgzImN6UjDlxv2g
sVKU0ydEg7yE1n8N/uEsYc+EhlerYl9N9ZnRlf0AQ6Wz3GGn1k029SGZRk1wPPUD
msoQsQzHwkKeuCI/Kd3IOpTIYnWPgNhmbbGvkmU51Ev+JdfWfsRxZf5JCCJ/+jCu
x9gFwvnG7vkS8PLRkYSd7PobzUylZo8sMxtsY4zZxtIVlzMxaJMvwgs/Vw43Kuza
SmtUt2v4Z6U+n2nICzpIkjdohsrSV0ddATv0VgLGwVgNQdXhtNBtt9xLmDnbUzQV
LfNQH2SvqRhYtfxhTkWNCgvksUUpaGC8gSW+wBulggz25jnnKV9zGE+sDLndeoWJ
Fp+264EgwK0O9grN3axyDn19kbZhUHZOsrod8uVBSw5o1bdhZ4eQw9n06cZRlCb8
dQ1PPzAGrUReHbXLKZJgJnQ4KQske99f0+2+GAIjvRgilZi8Vkc+RRv1fzDVhR8A
ynIXfdyqTqY31kEft6JumT9VRx5DYq9Ap0O926r1oksCKI7p2r0vsWbpt9MKjFGo
e+0COJyPpp7E5Ib5qv7RrGzhTVJ6dA2+UZSijnHuX5psxIe3L7USe0jluDzmuyO3
mYFaOv7FOJRpLSAUKxHVyq8u9GCDY2yUyD4MVd7+Izah4prTfvKiNYH4OZ2F9Jfw
YTbcYTvvNBOrNpHkN4uClfwBnTlxhWkf/SJ3RiZdNiK2TAtesqsGYygVGIveZKli
Liy0ii7yNhCKmpmvXWG+fnbyIadIi1zaEJtndZwhM5sEWwj7nUZrN6Ay0PqnbOBb
DRTCWAavn1DLy035Hsgg6FvlMHNUDzQKyna+3BY0VQtWPzL1tvTdYSUQ38RDTLu0
K1prY7LYOI8AoLEPWgqgrs3RkEeHnGwysE0mNGNKQT0SMmTLQzVukAzuk6K2WLLx
kWqwLoNZKu16PMlDEqdWYUZ4C1xDoSXphSVyyoR1Qualx0iopW3p/0phG7xa6kwj
kuFnF9MCtgg72TkUSzmcAiHk0wGPkSJxnACeelY1MCrZOO22RBiKvJFtTzZyw1bj
5qfvgArFRpi/ATvpNWLAapClGQsBbib19VKWT9DtiG4PZfnRFlXB3q2egXtlNCZ6
s2HvWtdz8+GYmcQdFkJN8te/ltn/huSGYN2ksgBE2uVVsEzLgclKWeqI2OaFi7jk
LNwJYWyLSqfJH052Ule3sJa+619bVCNudukm4x4j+RdNjCU8f2vYcwv/TbopF+lR
atlzIR7PWUjD5bXiU+auzC9qoENSQKQ3Uer+jCCawflnLePzFf+VEK7Cqd+isdV5
DxO+fmWv9rDIFGiEQ2+r4J+wd+FEk2VWkwmVOeV7itlh1TmKAsc2WsTigBDZm5g1
ZQ5tn7B+eZT7xKafvxFLNjEhVXx+EKaC8CdciXTvf6CpTHcJ6EOSk+bvL10Wq9Gl
CHQpojFP3zG+PvuvJIHZnAgBzEmJ1kEou7FiW7aJzB2u1KkQnDhHbndn43gD2lnD
VZoWIeubyU1Of3ZMkkVYIo+eTvQ5JlNuU2czqWFbYza6zibT2S13IlAOaVbGjk3Q
zjC2KcuaZDzpiTsCKyOkGK5vXLoyDCmvcedg5syYsR3BjPtt8PzTsdNXA3Nvk613
CXSSTBkxZ0LnSYSlph0/RQirW6y53RyiTYgkg1wy42P0svDbkdyt9MN7b44Iswjf
f0nCxGUXBHLq6kWVZNnlplyl3yQ30ppsXeZJVX/LPEMNURC3xMaKObm5sViaFRBU
gud8YOZXPUnAIfKyNCRLzvghWH/2Fzm7jkQU5nOb5GULAf2+lD+28eP8BevEgh9U
1XyBsSfhj9sMb9rEawgu/mRk4YrNVP3g/ckBYaaSzfRd4J1NoPn/PIpdpQt5uKho
iL979oCcYOW6B50/vRfWO4KC5ffhDtPA5wx3wf6QAWQoA8mejT65AlY+nnzVSFgC
F9LmM80+YKjAWuNe1w6TtRD5DeuMhspD1U38KKcqsV8lQG77tryFzss70bf86y1N
xiVlG206t/XDbJMtVBvfV52FismhnY+NzbpY3sFD89UTuzUZMlF1r08D0RnRFnZo
ei84U/YtFT5Fm8EAdxSkLDQ88XSLTcxTAWympXpf73y42FTD6PbN1DXitZhM9mPD
KXBriUTiP+qSKRJ6WEzVY95i5HbsNrF4YWPPTEvcxuhqWJQFzvtCznuuJ2+94dbv
3YUBA6UlWfXO0lmc2xXSQDx2MGDA/fZuWObY/RxVvoInvrik6yq5OlzpH6yTkw4d
EYcknPsR/Kok/yzxVmv3HT//ztE2WsXJMuZW6NjzT6KLpI+g0CeSgyY75yJ/YHJg
w+5QnfnG8fpC+fW5hI6t61wLuJkbgCTeU/iDke4NyS4biLhhtI9qu1X2RJfamYM9
FlXt2UYueFBlMGw9D/mhkbuHnRlQmuOfAJLx1VG0UrdeWP1WAaOB5JgEo116RKOF
gBPiwEwOxPpMJnZdyRDYrn1W6+L7vFSEbIrgvaozpROhnOSsR/4fyH5cyt9IuRGU
qhSXRFBMaKCuhwxaex+m+86iSACbQWslUKLbE6mmmp23uoV6RVSnxzsaaSuoJsxg
qUSR3SEdrbrU55Dt0yK7b2KEGbWwLr77tt5VjOP4jeSQuuRKE6NtHuAsau8uuYS7
o1BJ5k13Tc3ZqjdcHzjES9YtZ3LvOwZsPtp6ASY06ILq+vn6invJqe0OVqOrvGea
sNbXzQolcziGZ51zYyhsWckACLHiFb1YCDXu41BjDTy0V4G9dqag7ptdNkthxsmO
oX8MpRzAFm9XXU4J7wbNUG3CL8rf7rOxjFmXr6ujNavi24KfcPFjLLjWG9neqg/L
CSYuOSEaLMTporjuymf+5UuJn0g95/mNLfCmWzj2oIJ0PWALkd0/Obr4sS1xHCKY
DinyVChxnOOssFu1TDI/ZipDpGtYFXMusu8wF4nTlvGymdYr4CQRf2r96KI3dj/l
OUsvZxAuSKdY+6tTL618BKN8jICPTLaDxt5QxdMKdfvUvfxzEfK8LzWMQ/qTfwjr
WTbriUTy5w2X0z0HVRZtxaqgEYGBFcNpiNR0W/B11HYJ5tWyZU9C74T0hZgdrWNU
eYS5jmZqWwmbklqvhif5vvjlvv8wZWyBGEn8t2h45FWFqvf7vFyilqMJyUVkevDd
WPedUE+GysO6nAuUodx1IafALdJLAoKfxocWEmaE1mXCiZUkfw5jZB8loS/Tv4AW
LqO9lJdOk+NxmtLRxEj/YXXmCzDFCDNN3K5p4C5pk+xtA9tcf5Kaa2ufU7SxvL46
2chK99VGcATqLS7/2bOfdsngf7upv3iVlcBlirrYbFjNIpDuQ1bef7DtZjmsd2uS
jl2EF1bJufeVekwivHEvTpglYq9RYVXY/lH1pm5muKxBseZZhQ8QNJvLrfjo4gDK
UicEz/o7+A30ioy9k1DsK5dqCtQRSxlodwfEGjsjGnA9MRwaHxvSj9+nBwve32Co
P4DCpcP33WLEXksBci3p4BmFpwWoIllhk3fucZ+LfmBZihp6H8XnEDnCDqsMlgsk
xUzORpLMNrZwKY9wiSncnerTnzPdxq0zFelR11sMNiaK8vaXUKGzAMhsiN3UW4vc
oIPS+kv7bT1CZdtyu5CVOdFr14vMPYu84PCfUYryN3TcX/Nnr6BacQQw6cZ1mDHP
s599WBkz7jp7B22kR15LhRwaLYn3hsAkEPh/8ZT6wHPVkAIsZ6XD8ySc1yJ5h38O
vxtXFGkgz69AvEd/ld3z3LJ1tmru1d2qB7dpDt8yGrKBWZXFApStB9Iwo3Qtknj/
S3riwC2zSXbCZO3GVZnUm3C3oB1Qui/e7BbvrTuAVC5A39vDxQx+0gJZ6Toe+/yn
qZHkjnMxMFBD0rcXXr4SGqxPpZCKKY6PiTzcpg69Sbhe6HW+SaM4XQe6RGx4U93R
mK4jBHvfzwfgyWgTRpJFRpmGrxseDrUrH/btyImal/R+/au/QZPDVYmGvmZoa414
UqT+SPiH0IOuk1jDbVKOF9jrueIXawPxHIqg6MP/nxtly5e8wUZVOlY5BMADlTlK
hg9+CTXjVUl/nl9TGHKaUyvBLDqSReFvYmhQuqRs5Kp2/sZq/uTKdcDrarzH3p99
GBQEELDOW+a0324eUwRthnkTq8++iO+MLfsQv89Jl6y0bD2w4oRkUc/nmRk8ktlk
0AOmOzVAvj15BJ5OHCo+VWvm7DYE7LJb0FH9XwfUSpiBJ7Hucym+8wfCulthf/Ck
zEDVvbqq/qU9LSj6vXS3tKkI0eKtE45RsEN6TDHOkbrCt5qDpwFkJR1/DxYvnSib
o2GBBNDtCJuXrZHsj4XHRpGJMoWT/k/ziAXoN9rzYTFRZq5oeGGOX3YMGA3C58nY
DHyI+W8z6pPP7NazwMMSKVYpdjTTaa7x5WYAqdbD+BD3PlnVUnTiz3G2uKLEasoa
JymCT2Kja3+3zhhaJrnU16V7GNrVrQRbg605XwHNRrRvfC9DSjqj5B8S14Ba97FI
HyfD2CkGGrXmnId8q69g6oe0B2a4SlKB7YX31e1nFN8ddmwIjB5j7hU34RlKzeKb
ltMFMIf0Kt4fTIZE8JJF6Y0jvAvOelCElG9nGDNfn/3HM5IzDpPe8IkKBOBj0jgz
81Te2RN/UqnV3K6dSpOhVGpbXH7PU39LXAYDNMXM7TFrBePdyJm83i2HIS6uvomL
H/8GQvWPiauk4lpBjUE20os8YeEBH4TLyoqNHWTH3gO3pQWmW+08XG1ntpOOr65Q
T1yxNVVixMn0qaxroHcR+/P1ZRm56fnYB7QdlVLoSifEzAlL4kMIJu7KtYzWZ1WM
gNSwNuZGXxQDkeofL3s85jHIdEZA+21G7gPKyb3owajiR8kPc17Vfbiha9WvDSFb
4vB/MSw+CAsS5KqN9ZWAAHu51sXU7iDWWH38ahqFGwwVUQ4jDngQypVF/KNVEI4I
+Y9NvmDbKIHLM4g7oNNl0M75fwxhS2r4WojhEQAf197AudQrcr1+7OuJ5SKRL6pf
HY8NvLKjYHCno4vPoXAV1xlU7pV3lXy3DjUaXgXrD3spjVkzrfxnaMgxsqoc7GUE
MAfj1ScFK25bVJxG9bqqW1/uAm3wOKvU/3czDnYohP44gxGdpLm32sBheNnRLiss
ka7u/PsppHWSEXHfwa2VVWYer9vPnPH7MJC9vtO4zaUFefnKuMSFPTelDXBCrpK+
wIwigmyAClbPqJZ5JNPFvzDTjz3LmFKIV9NgHREMvG9MF+FpdIyr7FNaQsIKBgUV
aiQssm9iva8SDH9WN+i9E5PPYcKRN+vh1M1xg15Et9VM9il5wL5B/Y526mmzhcgE
9LOpNLXWnCIjwFI8vpVeen+w8PlWusWIrUccdOyIBHRMYi519lvqk9UftZEbNgeA
Orw4hJpflp97zgz3WYqBQ7AWizpxEcfW8RnIa+bEOSHbKFKStraXhPIpIre6eGMI
/gBrhBIZu3QoOTvT75v6rMeWWgMZitOb/OCA9CFx19ftffF69kGzatLOnwhmZjnv
wZ/oC0sPpRKdg5gOT6jzxPDSgJHPn/ST8vdHAqK00TVfeAJC1dBU3YZEFg6coQft
72snjPZlbRpDKzopT+M05Il2M3v3F4s72VhGJnYvalohOgxv8UZ0D4joQGtCWyU8
nYgCQImImHmozZImkPPOLqj43JijTFofK1RwLlZvC0yuHFsIy20EfafsLDPzKOVZ
VZO7fJjqivMpiZSFZ4bvtOSJ+xRkTib6sbFx68J6MPJOsujcL61wEUitxouyaOI2
jAIWt5CoJoh7dJtXcQUpWCjgTpsvERwYSBru3ARzqSFQw07h0Q+0b7KvQ0mhbSiH
k1Gq4yeM4Iayu5StLG+gZYQJu+tELvrVcSa83LFpWjgNrtCPWXmVXFIo195RK0ou
2/L3+vRCw6EbMcZVnHJFDMWgMDjSDQeM7RzkBqFBrJ1DA/AO4rnL9uPzvmslKvfp
uQsZ2IOT+lFcnRC6o2cCWUIEo01CM9IZyrscJ/ujBl/lom2f2/8Cp18Nsj1FcG65
HU+yR9vvwfvp02VnAsO1pyfQXQ3l4Cb5mvg62sqNz1L6clWRkTl8LTRypq7QV6x5
alkFphwqxpac3j5kfTVVW9ENwEbgU6LK150ZK59+GVLtMenoYP5ouEo5vEPJWyHs
hy4k36T/EEg2y0mi/BXs1/imNpZbPz+dmNH9yvbq3nmD8SGEhAWz1at1NlKIYiHy
Srgb6bA9vuk7xUyyGwU1mdXhl9mzoe8pc+TIiqbw+UwTQCgYccj8n4Nw3LRf4lJM
1NjJnXxV4b8R6j397OP1VNL1qPhrVc0CHCKbUYX5bs2aDKjTGHRaFmN9uIS7Pc6X
lwyRy8WLO8Zcfzi+x/x52fCoQcDFTf2Cq0ijM2okCifiQWlnFV/Aaj6C5D+Qmbhb
TELhfmY4PtHMazDjkvOIEbvJQ/z0Bfl0sxpHwcb+5iX53rWyEfapr+U07UeSezgI
6awilzOlz69BPNYy7e+r01DBaEEUluU5CcXuQksfrLYj6xMNL7m6prAHtBU1SfPm
FOJxauf2htpwoneep6HDQxfR9dBTg/iy45rj5sonC0D3sVrn7jnR/K5TKr45ZqTf
52R5Po09OnM0K+c+GZGniZV6VmtJLMCeEfZ3SGYZl9p4hk+kOCLpF0ysSzcngMbc
1W8HNZ2bfm8yQwyg1nMJqbSToR5fmgc8qm9s3Sj/cHSvq7P6y0CvxVQMtyhK/NoZ
Gp1ARuzvtlKhgQJRdQneqLdhkuE6lmy69MzV3W8iwH+eyF3GnuD+UvxzSuQmsNBw
Duz011dMJ96Q5sZH9MvGKQXE2Iu3kB2HWQfv/bFwsAczpbCVGH4psNqkQraYhg+L
dtGFVcyqZxA4R+o0W68c5zasiZqnjWG6i5M2dIOYnjZUyHNRqpy380GFe8Cn2qEg
EX4DSjpd/zERg5xYzRM4NOtrQ7RBZE02dCO3ksGJaju+n9R+aqEVcRs+ZJQhACg4
8DVHiQl5ScKm1nGAQq/Rs7aylA9Nd+ynVL0PU354aW8hfBivWm98b++O7R3Z1je2
a3IM5e1uAvyBW+bsyVu3Fhqq1qLq1rMjbU+5Kt2fSasZT9mNnl8Jg61OMU56nG7A
l6kL9jnXxv5JzJwLrgAxO2s9xM/m5VZlsDSnKlNqgCA53HhdDTIenBFI4+O9KDZX
0me8PwusSSE0hDVHvh9cu2Cc9T/LZPtV4QiCf7rBxN5L7zIcqyu5en4HGTTb9gLI
dObCJByejPYRjg3C105ratkVhK+9khp6lTfKPTn4Ld1adu1CFwYiK1tnh6v1ZBrC
O5RgATsa/iSIDV4BLNTDLLOUnT8AIY6+Tqk3j3CNLC3IV9NMVwTQjMIBeB/MYr7T
y7Y6CdDIkHZ47/ssmKfGyYLeSa8sS0EbujOfVFKUrscd2SL8cAzekFo4aklIQwJE
HvQ2tZEd/Sxi28dhHUNfq0WDRf8R4tpiMCE+P1gjKIepwgtIGXGu1FQphnD/7GSC
ZWq6mf386pT/3NWgzNA6C9TJZ40ifXAnihgpYmkQYVUfbAfzA4bA44JRvqD2QDNT
DK66RHtVCdxXT6UgONDJp98Ke/Kn+BvgfGKMvUE63OSoFrBivuzmP7kGw9w7HlPg
zbBcMDNJsJKNwnRQVDtz3zH+7tJ+yZH2TBSjpzwoOUt1ktarS1dVQ1XkcBfqmxLc
6sdC6YyiaA+t6l22FLIzcVXy2g+NcPCEPWbatYyriyWSoys/vNoqOrP5UJtXE1Gj
aKxDHzKfytNn9qag2ZjUPrZ5tYTGbSNpVcRs19HGdr8Qb13nqesRPrG5+ec9KmiZ
4CaRnvn7A97ZzWjetmonfo9+VoK5AXk98bsSjaWJyarZOmTXCJomGRvcoaILpgkT
C2vZcE4KgimHyaJAHha6JgcLF+tfnIdi9aU3H50UhcgUmwgm53zOgSGsUdOzJbBH
UU3YzravOFKdCkXq1yF5423W5bO6N6+FzUB2niI/spYdzc4PQpzMwurXJB8ZvXtY
PTS6sUp3uX8+miYhYqEpcMPJFapTt5clWaJPOeDNY/evndd1tSM1ogoIsd8zju5P
v4cLqcQcr5tYEJUn2kHioB+bXMIob5fk3dcF7Jd2OQ40aRRJfmUVCRdAhDTUs9F2
U2ImG+9/c0zMI+QmBlik0Jbgy0Z+nsjd9MzamGfKh0OQdzDXPreIT6faqc9mYUlO
Lo/H5ufcoNp96n84PfVTjp7UtuUrKoDeQ3FlmsimHm1LwxTZO9s73YhOBrSPYCGq
tKaHqBqvQqiTPQIZGgI5uANxT+SPd+D7rfPd1Ijets7zFVCzWudYf3gknfXaBAC1
FUe5JjUHdiPfbzmvd1dz4KyeHSHRsN7/A1kn6XJflIXb5a5WmrNBJm0XhkYd9ku7
VYsLzqGgq5wRnU49eFscg6HKU8lNwy/3apl2gK91JKz1nhN5YJqCmhl6ax3DJieI
o4q63OpTEJAPoRToCGCxHnmScTQjUvLTXv7jeUoFI0gqB/icMws0QgPWWG9Ie/A4
2dCYxIz50ukoyLmJZNfkMw6wyMJUGg4PJPleJFATCl9FhMCKwTTNa8audAd6dxWs
2ajZpToD9yUeQz+yCS+5ErNFGt6cTPN76+wy4Bf5RzFOvbq/4PHaSjiJ4dfGloUN
ukbqlaBKzr37YMH1Dy1clUaN/bG92YqnIJYX+owmX6y2KdjEaRsjkWQpxR5IobJ5
6M3t/skjunOP0belEV5RkpZZ0anoGVHmZAMRfFLT8VKhY+7by/ocbIpF02a9cHFL
KGBXv37LPec3OYNwNgC799mjXF1UV1sbKrebBCxL10BYaXNaBWBdEaHMs0JcB4lE
hGVmFAdtu6VSNS9AZtSVr2pLoWy++WkMRa1eDnpUiLRHYwI6aLUnr/EQRf8ekZD6
V1J/zU3+26I+8ChdY38Hk6G00H2ytElTn0sEBS+UO6oG/J6TcWBLApQ782tZvtrH
dR/bRqzbI0ur9aLbTLXkA3Umw10bTVvw8kFcDcuFuYTADUI7BLJFu8LkIj1oYQkE
BZNNCafbu6bA5lcUhWHKIhHKyDJEa41NKOH0EiJihV10QHysrmiJ2oi+JLL8viJf
m375hO5mhZdyFv/paJoEx2CBZOU3zaAVUiTnG8kloJsgswMnNBRCD6UBH4HOv0O7
mFUOOltf/hYpOvmUbdxes2Y/QaCya+Eb/2kZJE+Q8kRN05R1f/RSJqU9PYPalVz4
p+J7pqa1fGTj+2YSG3MyNI7zCqSTLyF3wC0u9sMCjjJPbfSu/yErcLFtzWoferQG
LoLYHguWqtwGJhoEGQU0GHvWdhJA+7sZsqDnMt4UIsEHwUZaFa0C3ZTMBRF746Bk
tH+vZw1EeIy4f2p5j/Zckv76ODwELgH2ypcMBPc+UMSpdXzGDUX/1PRUC0yfC+T9
OQcNzW8VbcNj9SlZTCIPNbyaSHhyCcuU8WqlLFj4UJB6r4Z6QO1wxeGiDvC69iQ2
gKqB7+TeGwTS8TOQP6uwhnbcIPOFaIdNMXUMcQ4njLAdtEzBCa/AaV5EFxAp51eJ
/Y5bqmfar4poGWQ5EYq38PRyqYBS4Ql0cwOj0uZRMEGkYCb3ueGKMYuOUmfr5o3o
QzkbiaGboQ+HDS0pbI6BQH3QXbt1hQEDGH9ONjwKifBUVZRlg+6P/J9tgXffhqhv
TOJTrbQbcPrvTdZvknLvC2OMXEWind8XvAwyK0Hjdzm00bRaxezIUxL2FqCJsDSe
5J1h9KGUpTiJHUv7Iv6wsufnmBXVZVDGO3sC6U2+fIztWCqnRbXb4ldUiK959asx
pM0qal29e0fLf2p2dUEZ/LBtgeBmGs561dT3GiNfW/aWF16oPZOdAi4LJETVJveL
oFLL72DHeqXwtHiS68DGb/WwUc0YrbteaUlRx01Xa46Mw8JZ0uWYaSJKkJzorgpL
46+me/kEyox9wbb9PfUx25JABc9gCicmCKDNEgXxD4AeTn4Bt9GfpVb15JI6LdFj
/fsr0g0/n/LNzDb4oCWjuxZQtr9RZw3FYxHQ8w5b+XVWr/AcKsLz601kuBmdAjVj
rZNlK+Wtz6Xyfn/jN71VaPDAwKptx8WCwHr3di1HJkP9wn/m2AHRIaT2Hp5nPSUx
AKa+JN0ZLDfr4JtuYDmQpbCvFVej91h1BmwswylbCzU6iEhhX4c3IZ2xdrNhFuRt
HafaHgblNL1owCjS4S8rb/JC4GRn6yOmw+o5KfU0zANV+VjN3+AHW6vbQuNxUGSj
8zn2OLX1ajhY8dUwuH2VV55NCYbMVHlxfRpKAtyyEgc7zBQ1R46DqjdrcyAv/d4R
te74U3NMQ1Ic1byLpx1TSGFneUbyztBXdNdj8uY1n0mia15ucp3Vs83UAt8Z3muN
jcxfjLF3SdAuTjkHl+nI9E7ew0DMdsPxeAsN1BoNpqxwxWZFruSV32TI5+YMk3Qc
+CPxG3ZDmfn3pvnf1NtUG+SXS4e8vikvCyThfSH8N0lkFdixzQ8viAC5S6w9A0kZ
LW/emMlzZ8TN0UJsaF2zVTHheyEUXKXw4hEuz1q7M+HAaRqpVULx7tSrbQHsBD0S
GUIGszRJK1AlYrxKwEhmjtWAUFY4NkeABmRApsqfPXSh61/cF0JwPfTTWFNKkFP+
okigbW2YMxvSAN1hwFluiGk0K7izxCPjqriM3rYtFDLUJ2HaQTVq/vw2rEAi9GgV
Ydrj6A/KhdK1lNAyTxSfQE0mASvA2/3muPykHmwzfdbvgwthIbMGMciqcWxj+ruX
uUC8ffNXVL9+Nwwvf6KwbACnVGIvrYXv4lMQsMH/Vjp+dXAOMS1Oo4VX/oX1f/hb
nwZwcjQN+o0hIaxBajvLf5orizozLw/DunDS33VNnG08M46vOMluR1oUT1ruggm+
sSJfjtf1LHSnAm4mLkQu+zKGPflGEVHou4l7Gv449Dd+vDHQjq2xT6uf6ssNctd5
24IQevW2t+HsDE0PT9xq76QRh8rZQZRVKkMqZPq3ULArbjtdFzWm3YseMh/up9kC
wNnooNX/ZUJs9H3yQ4CRzsc/77q4H4NjDKXq6YIiEeOWIYQJ/Yd0Y05hmJGi760U
/hxcKxUwCj3TwpsTW3BpPwY1mM2CWNT4xNm9jGPEAYTEHTDFUf3j5V29H0XdWi9P
Veywk/j+K0JEGHcFfRPc4ELSFkGJXlweHTuCBLzinvFsp/6alAtrw8t+vo/PQwa6
W5xviWNo41p3i4BxQgorY5+6uw7dkkFPKocqfweRrURCPqHFr2xMcwQpohrTXAhi
19v6VaNiP+l1jGpbOKgk+VjUDGNn3l3aGKcM8fflodZ4uQdGh1K8FHMVa6e0gYPw
nToayAVV7Q+3rhsoViXe7zqNK4VC2JfFdxWW/WgP1+skTgWSCiCglOU/6LQZUGRE
RVSL/6KaPw4dHUoaV36RZWkaKsa1O1cmledYhN52OMzA+Ri7K39T7Lwpud496h+C
R2K+v56iRr+AOd5Ri1g3sRKTxjy9FTWuXVpbOL+O/y87WQoiQMogRl6/TPBJyVn3
9Mp4vHLa4B3pVboxjBrzuuoofYjPYj/4G19d9UCKSQkVcBuBTiImJNnd2k5NCqmQ
umNk+EFEdxFdtGsb4BxtLSjPuzcsjHO6vx/1z5oMSe+PUslE00eN5LmsTWJ8UNec
DCJJzowfowV1LE3xURzBn4vPmj/l+3v3JW6FG8Tnee2NvXwuEA+rCJU3bQb1LHxV
qvEASnvSMMFE99RVCO9pTRxkwiBl+pdf4z0BHBKN3YACbH57SEvDr7KTGF3wksw1
aoLmQVmyxjPZAc/66QM63bxrdpXlz+u0KJFGRr4yvXzr5YTIO0M0dfiIdh65v/fr
+mWXmJfjDr8bXthsem5ER0F1vUKgrZcE8AS+rijBa1EgVsTUX84TZND4g72v1tNR
1haD8ki4co9w4jR4O0+ulXAvwc+z7fn0mEpSSsM6ugitjfiCc4f66mQQIZD+5BYy
WjlxaXJFkEB/z+Y742iLu3tJoQ/k8fCOuK0L+NOC2y+PH55xCrVpNnE5cP2sK4X8
gr42fdEhZyWNm12duLeQLQfXWdxA8IreM5Ahfi32EMysbnP4I2PdANggoMaFYKFW
DUVVcAXTTPX8VIK5npeXI+/IZHeQgeuKpvMBbZ8aTT68Fg+3homvmqIPbNAgc/KC
rknpDJz/l3Jkpm6ZKDWnVabhH0NBO4aegyzHg0pEQaXGVvpigyHKRqJje5gT9ev2
8fcimZYl92ASVkQIq5ukIYJXItVdhD3fvqM3N8+nPLJvgzHABtPowAkfuPOW98+1
kzrZjZy6FhqOb01mPXknkSOF2dnhIK9rWKN9q9ktiaRdFxBw2lMQqd04wqnkXvbY
i+9Qza/YvlGq2eZIdLq99wF2RleLAxMZz2dF/q4y+bDikpe7o7dFRGp3QAAAO27u
J6M6KUI+ywqEsBAM/N9iOHv8C4SY62iU0eFbNKEhKEp6vAx+BpsBOm4Zv4qCM7ve
tjNFLuUahb7PpHP091SXp3akF/PIby5XFXRqlxBf/Mx1Z9muWId5NgcvJUa7crW1
FEdDK5PBFCYJXUVqy297xPnM9a7RlwIn3Ly9uJWDJCvW5Zm0lo6nC1iBHd4P7Sz9
G/U1q8KS+gp67X1ZUuocMTGDc8ckxY/uYffXAx8VyYEKWIJtlmDvwaG68/J+m5CH
M/JjewcoJLOLtMpFb4v9Pq8gANBgAeqFo29g+Z62MQh4xlzAy9XYlsBG+M13jhLz
VUYkWZlli+bqtGi2WhD7mC/Qsy0t03skaQSBVmlei3VhCB8QZgKvwXofNu+7zlWm
kWzc3XvHQOGBPQnXLuiWk4cj4w0PWHGto4Ja23R9rrBDFO7FhT32nbuEbgqMG3/C
j+r1E+veFPLFF8TSI6tH7n39tdSDFzYySrS8AgCC0fShXuzso/98WlFK8KqAcrbd
UrfHKO11d5/7x4MVAfD0bI47m2U6HwlVZ2ZhimxU+HCFNi1iNuPs98cx6FoJvu5O
0ArIl95edYdl0a/9HhZ6jIE/c6fr3ImFws+VlYwc+1Ish9cL8uMmrQRlsUoZEkzN
a7Pl3T0jurkkBeo4B4UJnfSBSbS0eh1fo8NWWk7mfvlEd/DkuTJj8n1NsiV1D3al
671Y/dvDqUUA3T4V4yZfyQlHz3VjzlVdiM16UOJbKTE5mgA53k+KinclJICTb60q
sQmFNhRbfmbVsOr1xCU5VrFhjoYVcDna5J7sNQOC6SR3qSHLRYPbzKDYOmHzM7DT
BSJqV1jf8w2w9ckG+C96hWNJTmKr5xr/DncvHKLlZta5ncFxXeXEhOXrMEjm6Uec
RynBccRjdTc6ZyG54/Qe4kP/hYEjr++qKXRW9F4BuwRuFtkAtkXL5MKxIjgveMHd
sbihTWFcAe3RL0+1i1nsiSnG1b9Y4alKybxOoViio+fgAyTLWbHsSj4yywIUcf2f
vFpAASAlBa5fGYRy0SmGHAt7kbeGLiDhvb+QXJagl2fswC6kZaT9g+22a2gPgV7e
/N8gPz8zmMnFcKQV43SrOtWQ+N5HrgqZY5EjSiAx4+MqifcxikydvHR2Thg+zudd
K5Vl5bcAXZqM4LJJsJhU99VI8F8tDfPYLWrIOnXNa3lXXC2rovK3YFipeEBh3+Qf
1EIRKa0KRnG/BEKsHIQHeH2BvfBOXtPZj5k6m1Jm6loAF5s86LBkJsogTFWdooU5
sEaTMINBQXt4Jy52qzinqiv+PacFvDMz/FZJG24N+KPK+N++JCAeO1scOtsjR5fA
ciUQqstqKheNuKHPmOCRwYlgBLs02FQnoMt+u+ZpV/yvbdwp+R2fJIdyArHf5/0X
XIHmDsnqNoIBCMkhkIVm1Ud55G5QUnGUkw8uumKtprgz/xHGpm+qTeZJrzUTiw1m
QbcuXL16sZjQXygD24qwRaJCdEndyvFKaChu5t0WAEUssghrs1vuoqoEYV+y8V+U
5bxOv+WdXbuLkDFJUWiVFX9L9Rk4cE2VUSRUed2OoPLPPvxZiddaxwpi+yRvq8VG
3UHe1XpDv5FBTO4MDvOLvd3+5i7snZE2MIjCTZ4CDi20R2E4qUu2cnWrKkHT0q4I
xvPsS05ULmXrgUXN+0gjSl25Etq972wyI2JfeN+gJDZY51U1gclvkMqZOPlOwf3B
bR/m9bi0A/QSvuX8wyBbM5DaNFWZ9Fx6/400szr2Kn/HVX3zdv97NWPr9qLKLuf4
uYtu65/NrOwnZhMBPDN7/1n3ZfysJtE72FQ8s0e5k0MpVz2xBGSsZf57Y6tQXE6w
TcU8hE+g1Qs/NTSfOW514j6n5243Q/RS0CwiJNdYsC9Nia53oMm87Sj3jq+vQNMD
IQVfAZZyCugjczgd0PO2PECuKWPKp6HK6HYPx6LDUqoIVW9PVkLKtBKqfpxcjpan
dFKIMySlhtjrjob9JeoA8m+sCAAjwa6/so7YrOS2gO6Z+n10Hfric4dRx5pkby7I
X8gsmMIGWJ1LvcTYjpn3+iqEy+cQHIRnHm1Isu0K9V0jw4syYErZ9JKFozzq/oqj
oy2LQ3yFr7Dy/BeSPB4+acxFAlQFp8+dIxwNJUZoo0Sn3pL+2wFYthJSkzbYIUI2
v6iDlqxx51uPbgJ7ulbs1qyRGleeAWu+PYe5+1wm9V3zEygBuoj6d3O2kXyI7lyR
2SheHa8XGm5ssPreEBuiHfum6BI+LEaxwT4gdTK6yOnDj6PkMBgb2aWxqEhOnzQG
7Uo28LfJXV7sjtnZaJ5eva8QgVFB6wLdmjJic2FwZxjULcsSdcbH+Ez1PWDpOQEP
EXds+vp11VL4bzaxb/DamQBiZbLSw0kFg7XZI83iWCl4XyFfyrxEQhq0lySJTJHj
JeyllAUBO4Jzlqltvi38VYc6q6H35pMOszbDZy/8zWlwQ9UZE8Gknw5K+1MPC56J
IOCc3mrVyGkI/5Pl/cLzeY88pFw0wPIq9BFKwzYncY+joRLXa2mFclMtsUuRU5mS
I4JnTfLAArmq7ma373dRbimUAxEcjm9ZpsW25Gy3oW/T3RzZoeMDcWiCdlR2P777
xpPbGYDNz09+GokQ1pycOjAfpECEDIdRROnZjSVz44gbR8tz2ucQmHqlzsG0ZC/0
SwKuX1F8FQP+B6lGXzF/O6DEw83j4x6XHq7R7NKUvJ+JEk8dql7/Jz7lh4uxAFch
o+/FzLzF3Pk1m3XuPvTjltE2CCl2Nq6aUZwujQ58bjc80tXYYIfiOKqt/zsJjxEF
7cEokrbMMyNA9F867Pb5AY0p/dh4wX5E1MRYeVXO+/pveRixAZ61PKledQ25pB6o
rNF8p4N9Af4sPCvS2xnReCLOixiSW6Tldz8xM5EcyxSxX2R85vMRJbm4nBrBvtH0
N4hnjnvDFge6oUHr2NzO4jDWjdAiildecgfRfOtFPRdfIETfBdLbTq5avDND/6/G
CsJCkH9y5zxncUDklcPoHpHWeu+QkRfh7s2IWNuJ3RNgY2Bwq2VGMwrr+glQ7tOb
NiHcg4aXW3kzA5abCv/yr5nomBJ5Hr7uB7kLf29vO2vY8kLfzjbt2TzCypmEgEM2
8s1mGfQL16yO+2zcSKuvaMcKMITpP99QTpYTSuMSYu4QcEzRHperQPUSx387zRU7
kTXC+S12GJeamElbJmULy7FBb5xJoJ2F99NPls88zwgXy9yQjOX5AjV2TPqoC6Tf
bLqQkVfR64WJFUkKcp2lf6n1Rzbuf4Oz1TWJ6cV1nBiZTeIn+5s3ew6USydW3hOO
17c2zJ5iPVWtVTK5uq8FBa3wSJZ0QAG0TcAQJubEYDkvaHFGCZK94cUWxUBBdAPl
00GCttyCtxVqgqcrqhGyegLS2Jp2haZsXxsVMcSZ8Gw5gdd6DogbvFPvvTxse2XN
rlyUOYMERWIq26rJm5jmsWgg8+X4GbgAyZp806LzNAPSdTBogMPi1pvdtLlsDkgu
4pnXEnbsPztW5yJzXozWJK6rHhqGfm4X4KUT3PAdT+98p9/vxy1S5lYweX0A0i8j
XwA6QWflwDx28aHt3PAOcSsHoiOUgm44f4c3mkKyYNFFliX2rFKDWqmN2a2inMNf
poDT/6NkJdYMTCdBQ+R67U2eXw+KJeKPrM2IcF9BTnkdqICzN5CCShqL2iblDD3g
nVFAmdYIf33rjGEnzp2NDD36rfgtXbaTns5cAJ7sc7JkGDmgqiDa73PTdNA8uGG4
fhUf+nekv4ZTRKorf5D1BPHVf2YqFtzsCnUhsKQdcHyC2oV0Nxc9Xdy8WoTSBDrN
x7KvKctJqHY4+gGRazRPYoaXMSM1y5rN3SmphIzu78BsGpUWfkMiQPLbDdXwmx5h
LGDscqJcDIK/3ro4wXe41ST5AFcEZTPbW/LXepUTr8lOrjOOV1Xb0Bjqv8TGqotd
/g2dvkEF4fC47StcQVCai80NzlhYe4JywOa2uYCk313k9WEcmuQvkIk6U8TCn1FT
Cb8z4r2LT/JYcdUhTCkUuWNW2uRPQvn8EtVmpww/RJFqGcAD8prHyUFY+v0W7Z53
m1xvlHbUdMW7Gl0CbBb9mu8r5lRWTgKFtRpS1S9BgYpYor6SO4AUFGFl0vIGLFAc
v0e6aGlCgP2qhBcTR5nxYWd4LCjsEwl56qC8dIs28FARc1+d0vohENiEa6OkMbae
3RM8/8K+fS1SVnr0NYCY7mk7vUz2EJwrN5LTjNu8/5V4hEmQy8hbT1cNm/gUfNP0
tn5FXEQairkm9XUmh6aghXWVm5oiQm+f68A82XVGpTFDG7Yg6zAF3X3/nKD73tvb
vRcGwA4AGP1MrAmI7TGkY9pC1D7Jnnx7Wo7fPXvaFQg56Y3vz/Hw4C2oTVj1Tk4l
i0BHC3ezyM9s5BVP6O9neuKDl+lCOJnHZ0VOSB9AeG2yVp8j+g5E6DPZlXYcq4Ej
yZMtZx0oSHoAWcaBagRZxYN647QPfa62pdsHg4TjjfvajDjMVLbWpvrEBjh/FK6U
/P87q3D1rbxeQt6EL3pGn9sES92nDo+43Js74eWf9BqApll2Z9YN4rLwuG1OWdtq
/7GuxoqjpgM4LJgsOQ0wIaTaoMJ4ZsyDf14lLwF/zXd+Y7uRgsFtXcIPOEMzpETN
abYj8cH94/mBbtVwYOOBSpnLoXTf4a7yxY+4DKx1jBS1WP56U4lRUsSIIeXNuZ8/
vP2lgT2AHtW8GQt/DXrQxpLzFqz/Zu6Al8dZFqevu3Eob+lmcGwJjlFdhaXqecvS
3WaSX2CNff3aBSLLFNehqIB5LBCy43jGxikqvSUnBYbB3dexP6JvsJBsbEwMfPX7
nGL/BK7OWyeOyEinJFOh1J/hVENX2O9M2OZA8PCgHoja2oOym/nk49x/sF5pkS+b
FdfpKhtPdPNdsIcN9EQsRQ9bcGCxB2BQ5ZJ0OfWDNCx8fXWPCRzF5hAiazl3RWeN
F6VBxlBk5mtL1wf2ZW9rS4yLDKZJdONeq2Lh/k7AwFey7i8ENmfE0pYQP5n20rBu
S3qsLJ3rcWLA2irEAql2FFjKcUPHt5HigVs/y+QFdZSGo/ywZjMykl0izg+c8JcV
qHHJkU7Vek4RgRJatwIawYuJyC+tCoiD7kHlyUxeCrwZ3rO3c7EDSa70IkVbiqG1
Iutnb+CuAYWk41YlIL4D/YPFcQeY9KPjHzfZcOqlhKSLWZInBTv/JF9MChThND7X
I8k//jBah5Dur4WkpsLHkydJaC7u3NUxGFwbXxUNxq2zOv2Zy85oQ9cDilOPVlQv
838SHazs3m5FrXSJ81FBtb2bvV9PsgmROqK/0oRFB/VmqzIw95sE37QI493NLFWK
+jrfJ8vMXAIPSm7Va5pDU8a8iruAQ8YnjCqe9qaCLdVJQA1AV7WKhdraVz81hdeW
fr31H9lUBI/Vt7cXwRYzxXlF18ZBFWlXZMDhcVFv6gob6xLr49zDLibwLNFj3Gus
xUlfcFkbizU9bWvsgMNVn7RARnlGwMykpf46CL0wq4fz2eWuWXAhN+BrM3nEuxxZ
qa/agmSWbJzCtqTGsuC8tpVZtc/Rm102HeZYxK5ZCiqhV6DlRy5jtx2dG5ssE0LY
QXPaEkOuOob8sLhHxbY2Ux+27rT0w1XS0TspGyhnf3MzsXl7O+eFFs8TPeRaMKVi
sCGuZKsM4BugkQp+Up9cx39waJoZ1TjfzDJ/H+4QmvqWiwcqhn+ASMmuzQcHviCo
ItSYwHqbkRX4dBnWp/hkprro7KgxGV+zIj1PXr++hAzMLN6i45L7wluGUTN6kQ50
AVPUfeyjEo/BmrUertLQwCzBad+P1tiYWgll7G7fli7EQG+5CscIJ7ejax7KOpnl
yJK1Y83Y4OFZTvZXRynsKRDIm6Kef9bIIz7aSsyBdBxJ6K9EOJqDkYOC0Lham2f4
heQfepYuaHzHzMBAM+tJ12rgp9xSHzNHmML8iwwOcEBBdqYKTD/cuxUAlFTfMAee
dFeBAUnmcNSUOXEWyWlgHPr9/+voa84lsTTv1PNIhE10YctYpGYzxWh61AwTbaeI
2gi8rpKegE+1ClxePe/voRUR7GYaeX9VnVl0rVJFDFfjm4jAcOzHGPDnT8xc+q8Q
EqbQGhdwlRC4FDs36Joy8TTd8veTow1ukP7gN3t4FklBsP86ny7Qfgd/RAR62EsY
KYcLS8SFniOKbEaHh0k26kUJSwz93QG36xijtmbnjc15PQ1+SS2RINJPm0UPAi6P
e9WGlcd2Z6MLY776HN7rERcyrAN6iKbsPavaA0jjw+6h6lhl7yYs0uy/i/qdjdc2
INkdGZ8l5aa7veAbYHZ/NRQ5qQ/aWTdSh6wC7csKjky0fMFU5PPkddrM+8wVMAq4
mOQeXaZhCIVWnwRWGaI2AwmIJHud9Kcx85zr2ajE62ffKS3XNZ024cgcZktjX40L
ctu7xNGKqmUuAvuQzSscxvx68h1kQPozoC88rVYgbLVfJ3Rni66YOSBeCfBgVTEC
jT1/HYE+0UEV+mz7PMxvfd12YQJh5girIYkhvkJ1v3Jtwocx+znngXS1m6mItU+w
s4R+JND/en7yn8HEUiD4PJWypThajTFvMRpF4f+rtDge5pznLyxulNqEna3nMHSK
cOZJJwzuM3Bz/S0vao0xjrp4L+DIjaW1LmhJY5aZrLgDX3S6szljFD7YRI2Ke3eG
a/pkXFBcxc6aY3C9hRGM7605XCNOYZwjStXhRL3bJzXB4Fp8Ym5ziykqOUunrLPM
nCOf1btITkhTH/pmoSV8vw4ZeKxL0t+qI1+4ll3Cgi3bELj/OoVtETbT2Hkbwm3v
xj7mNjLAFc6Cwl5EHn6NKdD+f0GWqPOaXoNCmEhAa9KDIaq0j37DV2pomBmpTHtN
++ZZRqBcXA+V0w6NMEWCSLHE1OTkKquwr7+MPMrTuTYsioqoataP728ui1tHmnAr
OZsymfdai8zJdC3PkAY4AwlxHppaXfXeavZyPUb99PNQOMBVhAWEUeLKZIiSZEFl
NJ15I29MqKnFS0MzVDV3CRsZYbmvuajp7fEkQd07zgNQOdSuij+nDunTOxcam/aZ
ek1bDZf3zl7OZCsQZ4GU0xoroi5PAZxhl5C6XJX+XWOA/N6fhXghMTdjXbS8164J
cwmh4RSDu5qyZPRLfuIRusBr4utnwGf0XnCrzYGkb6wRMk7nfLYfcwBMcrd8Gj5z
cd7YL0EMQtItAxE3XZE7CFh5yFKTyB7nbtxE3IW54V3aw3yqDgPsP/0MSXrBKNt0
E+mp21EEKYAtiIgb1QCgn6Qla+yphQNLzkQk0erZUa4C0uDWzaYucRES7xxJeb6V
aW3Ll5IFTVrDt22eIkWKhMYHfMIrp1s6cuW9xkfdTdhKT8k9KnXaWw5T7IhrSM4N
El6YnYR8BgxQazHLg1feLC9eUum+16Eas9Zhgec3M4Tw97Nr/pgjn62+GQWWqCIz
QzcFjTMQ/KaOsYr7tiZiThAxj3PJuBKBtqTxnUnuLHqvMqU31t6jK2tbgbe1Xfyu
mWmTIS5YoWbs2Kmc2EoTxqYQ1Lf1jcLGP6osyuPsZkPbfS7PBiXzdnM3FCiYYzKj
+nHKN4k0zBg3RG1d/dwOwPT28f2dN7Zrhxi6LqN22VQoXxj0yrT1mJIkfWBNub5/
ajRGoacEiNEZLNderGzAEGhJwmzNrpycPv7K3ztCLuMOh2dgB86VkpzCVZQWjFBI
AV9e3qXjJy49nygfn3rAPKXl6On8xqPiMdnE80J62ObACDc99eTxsivkSJIbw4Uc
mVjCFmj5OBMBV7FkwcoCPBfxySHU0oIwQmuYBUQXeg+Wrt06E1EADU2e0+5N1ujH
0PskNeH1lGqIg/HfpnYVTqK6f7H/VNz74eNpu4KyiutkAwh3NAFm90jH68WELg3d
XJSYWoz4Irdxapn2+ePhX1FEpgeUukxoXfkvuAdKQoU5cFdUwvlxo02UjQP9INbN
9PLkNJSKsyppmSKJwI/PFIC4FHWSfxNArVhR4Sqy+zOb168c4v1INL18FMnoXCww
IOHAwDrtCIpJHCAXlLXbZbMxZAZPmudtYO8bGvHmhue5EYKYiXpYsAi2L/sJJwlj
Kmn6oYbbr7VeVezqQMHk96abwfo2POblJJfb7cMN2KOP/R/PXY52TSZpgW1+m5qE
4LKk/HXNUFzs7K6mTu6XayUgioI007WSONVktA2Jdf0XVWyrtcX4O0SdL10+6vcy
l6cMndrREn0BP12mAo67a1I7+5uKjkeIY3ocDSZyJi2DM+CnWiM06ZMGgbn3daSG
G5hdbcndfl9h5VFTY017Bq+iZc+BhfTmSjWQFKw+KNVe+Bw2K811wDyq7+7ywjWK
oauPv9DQtX5Ytf00vCoyE82ukvYl3S3/05U0p9K9ROx0kEf2U+peWQOTWs/4ykPr
S+fI1SUnQedyePJMPqS0wszkmUGOVP/ofWqCYwXEnbwsC0CsmHPYarGVyNZhRjW9
Tl/+4mUrkNbLppxbfY/eOzsUw+L5MRLVBQRs5f/kzSpI3RcZOEQjnEz2j2oIwbox
oV4BuNHdrnMFqO71hbw2OSFqJY66LBVNZaXUlP5c4uftyZfUeWxtTFSfhAXy+daY
28qfuyc3Z9iCP4j/pb/PL9y1W5GDFxjScKXlAu6+rrvvl5qeL9k5+cY0d4OI5yQr
1GqEv4n35C7mB1HP3TX0TRXBHr7vU76AZTIDBxXWtxsNo+dRY4FxjPxZBTrb6uoL
Yw6O4fmpDjAID2CGGdPDJ7SPw/f0ZoStirf5KjZU2fxrrY9a+v32VKyHzQfOWsZW
7S4Hh8gzNTYRcMi8h3/8p5Yskob9178l5hpk13ghmCwkAMS+u0mRKDKX1BRpRUYu
LP9WstoWnJNu6lOZHMY4qrICrTNFiWgqUn7S3VkyUJyz2U7Eo01rzpukpKT2qFB3
nda4WD86Gffh1X+05LXdl/7QLKrWHispWaZKB4mocYwkJeDqzqPRIQBAU9xJ0hKq
alxgFvgcgcpte76y6f1K7DnyPJUGsWeCJW6oFDP+6RcyymbsASAAWnV5ysJx4wgM
NfUkZ0ZR3JSHfjn+tKIzRfpchqDIDLpu6V9uWaEIfdtf7tb5shATgtgzRE0mkUEN
JaYkQVcoh9W5AJQs1lVIJYhL6e0RIyI1Rd7Zo5Op/70fyiBjfZ375vPGB4cRdQPT
CpWPHq0TLOmlVdyCkZYXn4yoCLNqYezY2YsYAEzeTCOVYHM7cPFvJIoelDNPUnYL
0TMZsS2LoWrxohz/E2AuF1uUVciNMKOSbrB5/6ttf3e6/mtQwDrbERjleUu3lP6R
0pIoR/EaIpIrxLk9XV4ugkiysM+s3oDofwZ8ezVVkz8ArXO7oAStdWZIIK9M7KTA
wURPSUoRS/+08+BSM5amYfd3s/FxuiDMRPmE+NQwmSM51sDhFS4vY22lbbYeZ194
j7QuszppcBFRxI/nS9Z7SNWGe3QA/34tC6UOLYSjOmlL1K13CiyEyqn12UsD7lXp
w0+sHJ3AsABv6ZpP69QtJOdqdtVgFshnPqwcJPzw4LO5YfTiedUvuFXbm2zzMzwp
NXk8C3fosPyT2WDntIUpYoBQGONIgQLUPc2RTIZRXltLAsl+mHYN/yzSlpoOovTE
DdwN6J6XKvdJAgjvZWsJpNkL2Z0WRCv820lOurTQpHLdJ2S3iL9snhTaaw9wUoxx
a+fCPTNHL3sPxT5X06Gpu/k+R7JWWJRywXGeOCZLFqq1hd/zul7dxx6T+r1fn7vm
yr/nfxwFSMIrnJkRLSbSMGHbM5zI56kZv/vIFYiTac3/SRAOgli+oGXTMIzf8tXS
r8c+0pAyIgaOJtLXmvLNt8Rgb48JCD4E8MVIMoNKtpIe6QcmRvLp/oB5gXYGTpA4
xoymnfjHDwtW5oVGNS/deoF27yRjKolq7+93qf1WAcG4BzJneraWvqzPe4YREexN
px67DQ6KcG32nFvrg4mKy/Lc4FbSeZpU2bh0AuHG+Zzo8C3xKKoPsvOXA/lUixAP
v+uNf32dCnOz+fLqI43ys0bfqZr46Q4QoQ54tvml6wpKxgmyE6i6G1FSvNw5+THt
+uz8nQGtWs4IetK/NW+8bj2VIE7q650ZOXEj/H4QM51pRIvUfCFT5hZo4RKQxRsT
XYVrZ6RBAqkXgZiPqln7zJAw9B8UQRgMZ5rbb3wQpWiUsBm9EUSCJjMvFLQeEpBO
++oO42XwRo6V0OXoBQVEWh7Nw71/XHxhdM7BCPeY1iqmo/Cw9umzsDCUcy5xBcbo
Ekv72uQIK//0tb29a4R/fJzFlwrqkrHncNBU3u5b3zERBgR2dd6cM3+vsUmoYJnH
HpM7A+wh4P/uA9narNyS9cs7gT4RFpkjgc8iDvZ1HV7/cQiRo0y1Ol1ffY0pEqkD
XxFMH1Q67VB6y50I+JEOi+6q3JDf614UPHqlNnVTTk3HeRk0ArVdDeL4skCIsHbG
UpASCxvtz36jycPc40efrDY9Ao7Oda+kQMqsRexBq/0XAQJCIClVD/9VX0P65mXv
tjp/gfgir/1GmmZjaXdb0hXO+Y9hojj+ge+4pB42slj0eRbgY1jBGF6yn2jWO38g
NuXBYXbvj6/NJb5t16tTQHl0+5Ec53YmiTsaDUzXOZQ38R8QaK1xHcMkFgMe7x6D
57g9eglJcZEIqOlmtukDAY3W9KAROsx1j2lR5fEFz6z3pKAtCCVTVyHkQArhsul/
LaMUTZ5ntj2T1b1RlkiZOA0YFhctuIE4TmMxSawV8cvSO/rA5zVhlJtOoiKwKBZF
ujKhkDZPcfhb2HbN2IcdVeADCv0x2eC/DITvGsOwHwCCekJ9v8bi48AKStunOowt
73DfVYp7NoOaZQlaBEm3krRdi/KFEkiMj6Bj+oK4KS8y0nDPfTvXqRrIqqiml2o0
5GPyyAeqQ+SjIrnT/2GpIo69yY2jouiiHdcXf7t3pitkpsfyW6MGpnQfWO9vPUky
ZIKW0A+MpifUjr04PZAi+YQVCzVh2YZpJvFDZnptlui3SrutMOyVhZjXNLMMfFdF
F0Hzsfvu8f6YXsTyGRHHzkeXa1KXGL6+vahTl2JmJFnhZzA3MkluwjrKez6oNlL0
NpTzzIT4BLwe2XyDnupo1eYnDJw9EMvv1MqLVh478bCph/QzxWRpNfepvsBZw1WE
YGaKHq2Mpg7Px/LuyRPlyGF+PlNoy/SzR1KtflpPgP26tzxv5ZBdkuAfzmtZ4mgX
VIfmZbKb7gZjzhUjuHU8t2tPu6tqZo4C89g2OYNC9CoNshjtObD9oDWLrerDI6tg
feFYyQ4a0MF6aShfwFfyd+ZRcULPBVVypRzHyaZApeytb2n4meexFFUZWwjm55s6
babuZ4seG4TnDdkejzctToIxOEesziKvwOuUtqTBL3iCHKjkDMIPDYXgRa9bMEzw
HcVGS5pS4n7Sub87OfxU2GwcEPiFMC4uS7/7mBWu9uBzZ+a+DdApX9RcJvEd75aF
LsfQEzkeuR1Q9mc4taxIi6qG1fgrHxsWJmabPVCECQn9HyOwjFNA955JP5qUMus4
YO/+W4czlPWkoicdwQijhp1qjqXeGLsqoQiUmxvxUC6Dd6rTo73DUl97+Ey+zSnX
ZUhfI8Q8pHjRI8r/acdn60G0n1s/wJUb/mbcqHf94bPTb0hnOfZjY40JbSpkxKeA
IVMYGlsPOOXbu6oZbhUGixHI2mwH+mo7NVYEAzefYh+rpMfvP+Dksys/DgCgXm1B
F3ubLKWL9CiHRpwIumqdR4LswnpxyIdDPYUBlAR2iQsLQU+lRpgQjAnTYo3RQnD4
gGM4Og5hjuMYAhNECqd6MUZkMWiBaxtUUv9zVygbTwma+lDbZ1DqORCKrTx4v06X
uZDLXpz8i+rL1SDCzKnmymDI92/6MwBDyNks2XsRKEFV0fceZ1rNRDNvZ4CeBBIr
DfCf1SMjo9jyxzkfBjWtlOSHQxgvRJ0UeKdER5g8CH2+xnw3jHzkKJq3R4Wv4zSx
wRvnmqANpfsG5O2ap4A2zfqYGSU8cJ06P5XNmU35bG/KYnz2qj698Afct/PSelSq
l1ddjP5AdOiOo6L3tDWobo5oxEr6BS35+FnSnr3S8/7qsxYDlzmbUpATVhYNLCsb
ZtMQYzHpL+nbER7yRQVNoYphmp82b86VPwtThhMXnbDgmvsOw+i4h4UDTJPdVRJH
6YafumJyZaHpq+AJlpOFWHCcKEZnEa+j8shg9pM9AVerkd5L0VN3ahL5YNqtv1mZ
xSOEcxNFZes/uSpjQxzC+HLWhfo4b6RR/PdVvh9R48tUvYV1ahqaJGGn/9iJWmbh
/xbvCq9+Kt8mI79tunHVPxSRXjBU5JT7O1uB8bsfp6dtvxL04XLvdz2jDflcigfc
8G7h1gyUmAHAN0o0uGBizPKWSTTvPGMjiBCmIFU08yc+4XC89Hm8GFj/vJXGP1Ff
msAfOKYkK6DAWt343jaq14WGHZjDWjyjxrLFFp3w/xXBW2LLi/sFx+t+HVFh7dIa
b3iAn4rCyVsEbC7YXTJlRH5DqMg9EomLr4fgNkogocxep4FuOycCTVzlcMezUlRy
qO5xHZrK0554Hy3lNdt+Z4Z8b29QDd90Zvjm47BdQ03OlrzPyLU3scBIXkgzYvRe
kqym109le1JjAUgn+5Ukx+geMAQp3AxmqSC0BPsiklUkIB+xWd67+kvo57Y7qeGd
W3yI33Ht8v7Amju2BZlAp/hHeFMOrc0Qmh0MeYyvil1TPvcr09S0Am7SeDzOsPuw
MMUEMQ0JqIpz8uA4zOOagUTTGQLsaSX1P6czjDthZp3v3TfrE7pJBPGRaNouyRu7
MToKl1a6ghgTN0E4K9q75EWOU3ya674U0+XA/au3ezS2TGbyIVkO494Db6C5XOrn
iwosZ9PngfaY60YRJOOSaS/Gp20IRl6F9S7CPsk2BIGonzVZUQHx2F8Nn4lnWbfD
alGLH3Uz4kXafLy7paPLG2KWmV1UqxL8XPatAdbrQr6HcJUP7S1y0xp4JiIZCcvo
nJqwO970Y6zFzJQr03RvgXrjKCAY5RzD5O+jU5s7geBnjo54I25N8ktQndsiJOSK
rsd87t7w2Gc6XNv+bMj5mpoW0YJX683TFv47lZXieuSaRu24yMYI0QgDEreUa0tx
AESbwe75JlDNS1eOU17vypxqJclOTHTLct+W2T+1BJm3vu/nX7WbXXnCzYJgXbOL
YMWi/yQD+J6PUKIl54IHcRZtK1xuRma+KqwcNCnvytvPrlXiRkJOVatgh6xrh2sw
+ptIM6o1CYtesGiP8Z09ULLCB5s9DuiPCWYShf76Ft6pbQTpVGFAL/yF2hYvnBql
TWXzGZGpmP13/NuQTO+/BEfUegvmmPu6Emp/xeARA9jOsOb2Pnx7aOglSv0Ejn7a
VkzPZ9BRUf3iUfaEkcdPcnMSsCqd+wFT62en2+dqo2m3lRku7LYR5VWkImokDFG8
2gnDgLalHcfjm7KyB0ZA0rYAppenoy8Oa+2ZoojY7T2gDddHg6c4rlRCOKe9r4cz
Ed2xBHTUwYNdf20p2XEStedP6W/YZnZCECa3ikvgOmMZ7n04zQGiUIGp7aKxc86b
R5slFnUQS+wHrsHPlp0d4hXrgJys5T7nAMRJn4xQ9OEoFN2E5F6r27x33P/IHLk7
KH21ZFBRqHKMBFLDsBAxrW/STlYaX7JUCTM0A19aUOADfJ3AvRrNw/b8dk0AScQk
KScmx+MofmtWMD2OkwipP+O8St5ngfuQQG37u0JhCi0z5LETc+r/bCZHol6t3aYz
cXQ3N586Rw+0X5m8FaY4w1RVydrcv5kgpP/VHRTDcOyYvHIgiONE3Jxb450B2aiX
WV3kPgyIExnYv4MDA3UI7Zd0N7tiZXHBteu3NXVD5JRzQkZJk7/sp3Xtb0eCJa7X
xMke1/7J80ItLeVpsO9xnOv/Q6lcc6UzVPwK/N73iztGj7e8dxKrFD52rqjbEjCF
ddvfWlELRNMaFKaA8QvCFnBh9lORyM91x5fd4tXGZ3XPu/eODiaPJHk1rQlAMdTt
zRTLtj1vineqZ+xvOX2kJeV8L1zecRL/fJ2J145gFjOH+CoKfy3uApDy2mvPAGWl
qUhRq4fXct+LiGDbTi5MgurFOI6LTAaDVIhCABFc3WvqRw88jecu2+Kt6OB7oxlO
wgUsVvo4Q4/n9hZgzuiKML80CXhbXtDxf+lSYaB+czTlBMZQLI1JAmCDSCqMSn0o
ka1iDl1mH4DVW+3pkmlGEDEn7dDLVbqw4BJCYmaSCWQlDXTIhvGXv1XtppnVIv63
N5uAFyzAcEfqsxLzVFIzLBR84XBRMjHAgUH1Au6NQZw8CUxOXN6ZKg5sEqT1JHJ8
xLT5VT7uIZ4oSXYbD4UmykBK3+OCLV/Vxl7G9OYO13jMg+yiA5WXdklbhvd8x1oc
6oBbSNVhWpTFQxJAcgAUH+JHiUNCrhFVYg7oVSl+tmAVmQC7h1doGCbdRgywivVT
MrNWQhSxn1kakgorB6QvrherUiOJ32caWY4eMDzB1s4/00NWfH3e0+OJEzyH+cu8
nsbVf+CWU4IuyiuTd1jAcwU5LizGXGzuneFSqENd3hW0lXQVT7DapzzCHM8XAMSt
5beRWde7+yTZ47fZ2VEy0YmwND06CQELapYmm1WCevUqGEDVv7DOWbdPgfsPcoPF
vNbf35fsivg3T8IBKyk0Nre3gUeaxfv5jLCiOiG71t3tR1t5iofDHHc6JUnMemdm
Kao9hBvBS6SKj/0G8iUlBAMiMl6uHyEGjvbC/SjeJsbzulJlRJXoxqrKklK73uwG
rNLA2Hl6+zA/XgHIxsR8dMITv8AIAxT9SM1cPBR62Ieqd3yMLZiRAYbvyQQWuoBT
x+6aznwcbA1Z8/jeHapyI2Rwh5QK8oKNQSyfCIbHVgNNFOd1O/xzOFMQE+FR6Pb5
N8k5ZZkYZXFuI98LEGvtWpxtVPEw/1DmrpjIEjGKT/ZmsGZro1tEbeWkW8WBPr7W
cWSDar20F6GRWcxPGDoPs+rkFIIG6C4ke6855xkHLFRojuNPZFksZlnW8id4AV1l
IAWKc77fj3ObPFhNVkuKWkJsBGOEu7TbEgk+VK9dqktkPZ+1XU9rZdo72BZZURwf
xS/dDhnqyW9HTPc8YEZiFrEE53AKIQDx9vCt4FEKFEAIE5eifkp+ldacH+T6uW17
JVygHFgoqgpZqHXheYrfBEZCTIUiYmOBk9nWoC2+9l7HEUdl6zaPkP4L9xOgdmiC
RBl7XD/QJCXnDsAUVzaQZ76MRDrcXUicStQeAXTp3aRQBnfgEL0hMkTx9fLywB4Y
1I21wcjPU/oIPviJCEAJ7lCb4X9YBWieVpk5mazQD1V/BN7FMxvkLJjrwgsc/Ric
dNfWl1dIrdInR0kAsWCMyGZtRR0JySDe3a/g6JoQyVSLQ+U+XRvSNcvIum5Ut9TZ
BYldaatwbYl/CLwZo3ym0dktK+WpZplvyUs6CztBolm+iAH9PWHgHJGxKpnZtzf1
2yJneaypTg0giQovtBYmyCk8u6Xqi3W2/xM4KInWuCKIQEWJocDD4DQQqvvGmI1a
hRAindQKfvEHrts8h5a7uLfIwhVUqLhrf8qywKJh0eRpRxbV+iRCnAQ8gK1NBVEo
jEh7Nx2d/JZbGY+5RzmUFs3wOg3CGc+ksZv1+Cg1OIcxq/8zzbgBkpNzQ/trW9wb
3L8rM/uS2BqyynNZA2oqQBNW/E0NI4QZVxEut6fk2/IMLNA9gGNpWkHMG9GPvVAq
I193UCLstI95lbPoFLmLGGC9mx8Es6TnP6cFwZu41WwILGMrT3cVzDuOzc+mmEH+
ztsRosu6GDpMUf79I2TDSZrIORPk/T/QjD+Bv3qPvOD5NghlpoXJ1ykuqpHyIjfW
NUatju9NWCOUS3Hv7ch/N3ira651F/yEfEOskcWjKjOFQq8iKDKk4Ax0tGBZ6Rmu
82tnM/NfkqHwS4x5/H8YE9X4lp+7i32OaxuvXq92w96VKaKuoj9Z99SiOSmkDh4p
qLCRvTshAb95N8cW5pVasZKVDwnjkVHy8k8yUqiVz9bQhBW0g16WgKzLBSiPDH7v
mOD2jfJW3WTouNdkDe44Gl5d8knQSwz6ccG/b7+EC4uityHONzbbPqwWmAoD1UpU
BcAJla79RKtyarXKhatSL0cCOhYjeHzKPSUCDS9+v1t+7qyJ9hYeIk4GghpiI5GD
QOE8sbxkJBezq3a3DMnVVbRt8lrPhi2ZgnoNLEvVd+gPBpIoeJmmBA+OIyOQKxSQ
+VyoZHewd61mBHhWpEFwNZ3j6WW77MLIsA73WDabGFQwPqKYG9gYv82EbPXyAhrR
a147PjCL2XthaRU0G2eEygeW+COqOFWY45emtpexTTLXm+tb13JNoap9sA0e8qMl
bGhGQ9S/9D3Xg0h4i2AaaVd59Z6/AS4TA3ccEBLzVNS6SMAk3elStzeXLqfVkbQw
lhRMH5xeQ9CAxwbCOyWOIa6ymFn7TdC59yXN18dmjT6sDyHh9wMM23hIRdv8ePtS
HvI+YODwQOIblMZKDsiaAeYwCIo5kKhT1VmCDlTqQ9Bz8oeziKfhc9vLmBCHmDLW
0F0YVO4DKXhfgfyHmQr3+M+6yc9kAc7FFgRzmFIEZBESNCFFgLD9ddxgGBnv71eT
dLbzZsTnnLoTZqp1xhyiN4F6Ek3ih1RwE6r5k0ZL3pab5vUZRABX+Q42aZIxiwYx
F7mPC/Lzh5H6EVaCt7XP8Gs1EbEFuTrIt+yJRMvXvhAhJgg4F7wX0U9qOFhujV2L
fo65wrQuws9ySeN1MHr4SGH7fFZ/IqMmEI6HLnCar9oqFRO5+7TP5aKsV9qJu7WQ
/+vaUymZ1M2CmhXcTrDvcMBwQgNnAxafs/IR8xxIDEYugdp6o1EEZGOWnCNYJrWy
Dj7k/ZnbarOHTgRhloEw6Cespdg/TE3MfflhUswNVJRLyxVsHPZefeAVy+SVveE5
tDYRqEO2kurfYP/+EoyWJwcZtsm/koECd/asZ3ea3hmk+xp6fBECl/JSD/jue7CM
TfQ+AJAYOq/koHuPolw/ocHq7E8VELZKdGYLamvPBUxVKtCDWt/AX9PeuBokFuc3
DpYJHkPHbsn8J0V+oaooRmKibrc2LoE09bSpJuwcMqScy3czXcHvhlcPWq3k3yZG
KdSC+IA01anvjszMKGxMxUXdegqkpkHx+zngsekclrckuEM49BSGGTRnA5o5jSLX
ImZkjaG7XEGyWCXX0iHPCOesBmawVeOreNbg+Rv8YBfJw00ML3QBRGk02u/1uAGL
EGGQFZsnON7uO79sWNgftJ8AZsOIQ4woC+WfnAiD4e7KAh+9tspUB+Bs5CnL9/L1
zh7gtvH5WINZ68lPigDLHFn9J4gECjPJhiiBs5RCfdJCcf3m19ypbuBqQAbJC+Le
apGZqMtETVURutonkOvyXpETbjLFg36cSTGuhg0KqnUOZJcYWJReplg+FQ0LOMoQ
+A5GHQ3yJdlVzhF4IQ5H6tUuX39nYJpx2PqHRamfSWvtOBouGvtewurSJN++6z56
lCQDtLsogBd2cqvRzbq7VgTbRyZvdsrlKxmeJjpHIdNRrW5uIDNzYuHkMIoe/19A
FvpIUn5Dm37D5MKlOkXwRShQz5fHu36XD9kTf+UKJh8ForMXVX40rpf0mCyYKa+p
7ukc0b+V4xWHur5yZk+4g89XUi0S70HankbUd8nhJ4aj8vCo5MEPTX4t0uIpdL5V
MGoHwOgsHaPWIQZ1FA6a4tBGwG57T0FTbDzVxqTQrRFN//Vqy/6I64s78VTR/aJy
TdrmEkkzA0TeDcw+Q2S87Yu6Sxdt4IkV2VnPK/ks+HBdF8u75yA6dWKMBG/4vGsC
LfgnwCOhyh1Q14VoFHS4Pf+HPZaK+zY1z88GVtBRfo2hiK16mB1FTqYLdA9xbPmK
mlaFHrbOZVI2dSC8q3JOanhujVhg81z26bI3LFIv2RnLNzUhqkGXKPKZIqG8x/6N
BlF2mHY+4rzz3zoADF3yuHjHX7hwavwy+xuzFw5UYR5Eykgb/eXmtlPTYpZsoSxm
6qc6TePSR/eoYHWOHJuiEPu9sQCzI4E/AZVwS56T3y869bvL9pwza0gN/EKeZZlv
B9jGoQsBYkUbbABUHpV7ppP2RHZfeW4KJxRy8nLaeFNrg2M30bMsYx4RecpXwbO0
H0MC4BGU3JVjuTTCqpaIro9xdUKxQdeCo4lf9bR/ikSbjtCl5aqvlTgfZy7uWG2D
s6S6Q2iMarA+DLCA0yLQDkx/zT5zVj4vjrdwPwqVnoCY3nOq830hTK8pWjP0MJho
qDIIusLBCORdGyFdC2Fn7FVXf0n7vnbolydsSwuYlB8BRqUfD/Mcz+bog9AkPZet
nWzRETISO2RRj+emhGBDK5GErqyKB0MukbvDHV4Jhl6WC8mPfWfV5XMPwUpaIw3W
Byd8A3y731HPWQ41Pml0A2squCwFITh9DuQqJpgck70NzTs/+0LzrK61vPY27aSc
r5NUh+faXRd/Ao8p2K9oPWmV1bQBRBGSYM4RG0E90qqKIoJLAq/PADGDGgmxF4jf
eEEGApr1TXuH3W9r9TryUvREo76XV2i/jeFzM+88wRsisRfUG5MVe/Wcxc8wDMRd
7YJ514x6dYa+HeySTna1Ihgmru17tPDiwqAy0IYCB4AQkr3k8T+oe+GsfnF4wRPM
ttTyv8zqd6FASmgL2umgT/QTgpgwxXz765wCe2XFyy7htQOm7BGRPhvv+ir8ayR+
vJ91OJq8+R6CnHDO5pxqPb+ANR5LeILqZOV9O2QyPzviuI5IKGpjbNjbyt+g6lpj
A5R+nGvY8OIhOMqxpMMhbbh6XZG+4laGxXwZ1POKTTiW2oxS9iGL2+GI+zJAkZPJ
RJSATplEb19YJuWdydaEANS8UvgEoM2ReJu/qcSCwJQxfoeYvbF+ZjcYPUXva+QM
UcDwMLoE9HldeW6i8bXFQlyk7vjXPyL9jAY7a2KEkAnHizotiEs8DTzCsZZ1piW6
ifevrNjBtzv2FSW57gGVnWzclfQxqORSdwWd/k/BRHueCR5arDva3mt2NmJU8lvv
we0vzTlCGYCftx8jqgXJSwG2I6+smBm3S3W50qD99rHpJkHAGVbmOs4kJGGHLgA5
Hsy5zNiOJqpFruOiXLnhZXceGYwwyr3i7KlOcQt3qWu0nNt9Y2YmtbpbUCIWvIr8
UW6lrA8PyWw32+w/9rl5/jZULKjW15AgYxFIkHX9RX2iZKY6mdfRkX048SfjMnFL
gEyAFML9lc6snLdQXK6gRuHbWmTutqEi5lPZwtNXI+VgkaQkjCXJLgwdCNjLDxOV
C8ESyhCrQMwMxKY1xL2NQReLUoiVjlmMdLGg/6CQWW0/V35pH6x5QZIN0kiJ+XoO
7mKzkbbrMY32QcXoC3lKhpyajNs4YCUC1CSTXwl9shZIONrArbzQppCnbAcYI/0i
6dehaeMeEfoZ5I6fAawwI+q6EQxuVn2Q+ODmBeLfq8mW2FKf3PFQ4Kq13OqT5496
FuZHanbTLzveodPIjy0TE9Tl9IV4FaWZwO/dMfrJV363Vr/89dQBZQw7/9PO1m7c
e16JG2CfLpNRAdNzEwVa62wNhFMYTlloeJ9UksGLbDM8r3Ht8jW3/4MYd2WZKkIj
rGbzBbPCIns1UwiiKu9pkhv8mG8jWx7YiEHaO5n8GCrfkuzcwE9J3YMmiO82S66B
R2twaEcOQKcZkRkhhSUuFt6Cwc6tegq6AXNxhNyxyDCAE+m6yAt2WrDq6rkC0E7D
dMsSiRrt/r5ZRSzzqfYqr+PG0EOZJql+gF8h7mDNQ8VYRY6XeQZK7K0cvRRcKaBw
DQBSdjgbqGIT5iL5LnEtRGbdVFgHvqC5w5WHuTHanbYcnpgX8lO0TnCf/2xNEvNi
TbUQJZFkQ3+6/xtuzP0854EEacWIVmI4OP83cU51VC6pSlkKj9izPAQwZWQPT3dO
T5/jiYSODSM07jBWhn2GiHqtHWBv4pFBgY2zC03DPa5AoY6J3AnBKWPo4hnzbVa+
EcltL+0VmYke6/TFhxWO+Ans5adhzY6n8UyVOT3AiaePoBPTq8wkATumc4OfMcZq
abAzP24Gqm3wmTnLDjMW9rmovNME52YqwTSfZGeNPDgf2H+12uYg36U5P59fJvyG
L9Rn9cinlHjFJsxl02cjagj4HoMBtEyI1Hq08VBoLkl6b7LnG5n6fiA+jimOGRns
to9ECI4vE8RkpHLenr+4mFBU+3rJcuzKtW71IaCTIthYqUAqpNvQB/TahtMpQYuq
1d2WSjL+UvzYbKwWdLXh2b3siTuV3F5IjtFhbQzHnRSafwDQM48KlO6ItSYY6e8i
VvyiYyZoU5U2muickUIJ7PF5Z9BYXZTH+WKDoKDW0pkCJdx+NekaBNGA96so/FQe
j6CQ4WzCD7kTMfXsUWvR3nKrdzifH7GT9bGqNp4S/2+6CmJ5tkylEQZAbXwHr8Bw
PNomAKxp5nkCeRozhU49is8q1oxcGTJrudwMj85mzTpRpbnxQ26mUxzTZAXBInCI
eODPxVgUSb0+y3H8BOJZYWEY46YZOKRCyDDrq/38gfIWkBAqWdBG5gVuyNLuYULU
I/m+p5x0OKUT9zla8i1l0M+S2uk6oh4il6Z7bMWGn9wSD1+dhYIBaxtysnLfHRfM
eaQEwkJeHR2d7vAMRjTPsLnSWPPVeGCskMuDk5AsJOx+hrA4v2S/n+LT6xvrKUtd
DfcNUFLW7hZ9iETrIeBzKi06Ef5uCax20YwTpFEaSv12/IaJIJrifl/ZOhL0UFZf
CIlaGcLvgXA0i/pzFEMgsGkbLgVRzhQeE/bQAqYTly0i9lrdWW0Qq4ghU1STfvAG
WZw6Ou1eeG9lskwuitfvENS8bf9wmsgaBD0rTXtu7+QN+I7V1kP0vwD3NkqAMYlX
PMSTOeiLEuEarc5Ic7gXPWSFKYdQxAm/jZguyyLCGMQp6wp3g/72e4Hcdj/OP78p
ovoNPr4QHvXW5l2wJYlRdFE5M3Q4f4Hs4o9wq1/09Z6L8MKgIMtqXHGlmS9QEI+v
7kxawP5Y+wL8HHXZC8bdkyyAs076qrUPZxmPJFUSHTiUOjARVGuLnZeNa7wr6pbN
9sTIDsM3vOMo8zNJdLBzQLgYhabNXb8FlpLtZcYPCgve3jLErkGxFq29V3FYmBK8
ZhOOGS4iLvgoAQjyiiKIemKD68ZUqB8xB9WkfhS9lKeigcXqAdXmEeuA95casYQN
HbA7C6f/Og0AzzH5JitAQvs0JazETT1Ay0H7/GrT0I2v4jX4WezRco/eEV8JNjtl
MrbFTPrhl90Y8ODtsCS5X8RB8OoJeWPqN3mmso0u76bx2FVjYT+xflQrZD26XiYl
FoSF9OY+L6slwNG6YQPoyhCbF0bMCbxW6Cz0GFx6ELflhxpWfekVdQmoMC48WC8o
eXGA7aYwUsSAjRNsb/pYPzJ/UbKSNPmFOH74JAkhah4WcF9653pn6+KbSG8vWCVr
l1257ymcshxs7sdQU3ejVs6q79SXxu9CN598pC9wW5PF22KjDrGiyREVBS6GSyQ0
OoF+C0nj8EnteEvmXwYnjqEcFqVCOBcAMfBxDPPfZP2KwuWsKJQJ1XPbgfeAHBK/
117Au+aA2d2O2CKc+1lQ3OsekPQlu08ZV/WFzeUfb0Nr6jEdYkzv9hWoqVv9pZvO
uXYzMBN7ZIruypM1unk2/WiBmmDAv1Xw/NvhjpcBCRz1UECuViU04ZuXsY/KfI1H
aphqzBvUsE/zYyRoeYI02Wz3Of3Uxs9wESFAbm5El1gWsxSfZDVgMPQlWafYV5MD
wB7rGBhVJBKt0gynQ3R/xU3PNSQsxzy66H6qgsELtiAghxV+xb/DGvBno36TrCCq
IFOSnyJjN68FSdJzbpvMpuQvwtfg27MZAJ+3DNSwHXYl+PE+glz4D8cIzuq0LsO4
EoJegYFAETvyURfCh29ReJ7SRsvVNNQUvYyn6lVG2qJQsbY6K2/z3vy6zYwI5CL7
WB4AnC1OcIRhiidK8eP44uJf9GyPfnikjGfRDDfRkRfn/M6130k/5bJvaA59MLoG
58tszU+FgdyC0S90Lse2+RfXyfHvqRsmjHSbzm9vG0j2gsgB85s0vSDwRkw6UAUY
hZkzESzDD7aWi00DWNSQoKAmlqPbkhgH2i6ueNuQ++dq1EkOjfNBNQtJA+bR8WDI
jfml3loJMrALKOBOQXndTQxaO+mf89yE2K1rAmoqcdI+xfnktmUvms2Hz2a8LmtO
ZWUGBOLseDitH/YR1YHWst2XOztpvZEJvpcikBB6vUfhBwi29TeDJABN3O403o/O
30oZuLfIbG9LaMWG+rzG3MXuK7thxCAv9RvhzIMqEeAL7Dsvb5uYOQGmePtCCAda
XRnKxz4i+GOtFFxEpzB9jNj/KHNvBI3pu3eCZtstthVyxFHs0snX7uKBDFS5ZbMH
iFQM8KlW4nhDa/72RDuAUiUESOP5sEbC8tAzl1maj28MLCFz3+dlOxVKfxLHn/+j
JjCiJDj0qanbGNu20cE6bh9BpY4tVfJwi7TU57OAuhhUjL++FoSxTkF137AbFdRJ
KlWQhUYfemkJBzWt0pue95ViULs2KUhIQhlsK43spBbJcho4ymaiJf6WsArfrleL
914vuia5/VO3IUqytiWr7OKEhcpCkDQZmcPQI7ctOUxc4q03YUOYpWxKIuQKh8Zn
CGOsZLyIin2cbGDwCYppTu2a+mQs5FLdy7n5j9Gc8UXOrXPecSaGuBv20PorwZ6H
abS2AZ0F0LewTf84LeXtUBmNonVythYTd5juMohGjz9jNpBsdOmcm4GGHolHjqrS
dY7RVPOa/vf8vrbeB8EVBaGGOC5aHmK93EHCfkRDjnVp6f1an4dsXtYc0GzWGOyS
L65A4avzKAJTDfLmioYozwnBR5gglNsmncsPYkvRo0U5DKyw+SgCTSgsbd5Ed8Gh
CjJ8FWcO9ton3SX3CiAYPRDVFtkSTfZLJ0Inwvi9drMusTBWrHH23KrbzB3kCklE
MtAH6MP34MBW+yEEwuNxRHL0HSiAWoAKRXygIg6d+P48qoeFgmTHJI5s+DhVg9ZJ
ukKh2+x/A1yA32QiHBafw9O2yyQ9OzU8XuYPvr+TE7csiMvJ6atWDdWp2LqeFYop
C+XMZd1WiivAO8UVkbWkyvEy9v4iZ000rpUqNfLaeauu2kk5XAcEEV9I4FRBLc4H
irDkvG+ONvNW6xgUGcFqaa0Nvcv+WDVoMJyf8mMt5FuNMc+KXPfFtJS3VRdIRInd
HYpZhvVUDdwtUsYv8+GjIxhg3X/51ZR6h3bvCBOL6FXNi52JOFemo0AzOAWH2J0t
SX9zGszOQ2aJyriaFM4U9A6Pr/I5+N2tNRX6LZ/LgOhm8LBBGGNlSPVTQZJAQAgh
Xgy/dxd5p/axgUaDU10Xke8c/ETp69iPp4WMxRUxKDLigFmAI38JnpcCfANs3qwV
uzvfhdMVEM/2yNyWxV4CDouEUIRJUKPqoI3+8C+unXEX55hWTxp+7PqMVhgWKOZs
vgFHVtIJhZf5KrErntELtZ6r0IQjz7oOY5bpCiOjv9Yq+4EAo1xhiecaO6S11r1v
u6miohNxWql3/tjeP1zXCixOEUZTNhiragwPER8Ut/OKIDlHrBLQDW0XSVovEHkH
I04QtPsGoTHlXght9XXslGdKgcX8TXmHMPtoKMZoQJynLw3d5PFBc8GtsTAPU+TR
qm2WARhH/O7SWgqmIjogW9LuzpTQvTLQO/xVH/R0igesJNmVS3NeatiFcYvN4dHN
7QYplqRb94etF6pUxhI8l9LKfgkFzyjNGqTKmdvE8fRcjW7D1qmeL7lqgBBmo69X
8yuPZqi9AC+Qnd3KWMvhyp7OMhBS4anuQDwC8pQx0RvVS8nRbEJC5lxXx/5yNUFY
HOYGoNFgObXWRj/lc/nacvwfhCRLje+lkXuSmnM8G1PnVH+LOfBwmMzt7qfZ6/pd
+wS7kAiN/Fbv0OcVLsUNUGiYCwEbu4BghSwL3r6qDREz+rPjANYqJ9e07WQi+X+g
Zz//1HCjo++K+p4gu8PcfunE8ET5GtjeF/HZZvV+V1Bdm4jBFDIeAs32RgxsbC7b
MY6zKh7ssOXED5+8pFkFvm9jnQvs5GlOTphe4GpVkaWz95R1MYMvlnHYYTWhWXQo
m3hA4+B0CMVaQ4C0l+siXs6plJkavIImXFWzL3ZdGqZc9MPhxEYG3yBH3UFqVQcM
xeHeyK4EI5VOI9X7SbBg7BGtfrwO7cQBCl184vIYnEW7agR4rloKchDc4/PHyzKs
GDnToqbf3W6Epn7qHl0i5g9zkIWmMpDteQy2fsUXvwnVU3ds2GNtTbOdje58Q1ED
s1p1QzvroSoe9kur0ZqXJBWIg8pk80NFst2gIIoSXuB2x6O5AtXZ2HsSTxWFAhNl
e2JdfhLXWxQoG6Xzyse2Y/BGdYq1croD2/eZwTEFAiBT/dfLOnVkuEuRVWQTWq6+
odSAxvYpoMM0riclxUdYx6TlBl6QNIcPvqVJPBsMnZqk30iS6FrjM1ak/3iJt1OH
VNpuxLDuq6CO/L1Del6jO4LHyRlKyMTTwBoLbNnKgO3Obib6fPjSxVIEAE45scYY
NyyhB4ozgl5EMgpRNBiGRxizz1+VSZVUSzRa8qx7x+w7zDdVuIpHr927osdGaL+0
aZq4qlnhvqh9C5NF3p/l17OFYveLirEjhOCoJNET4i+01/wKAwtCFXOY5KGoTNcy
ypdGHF6kmuj55f2npAItiTHULuxc7jc/xUaNo84DlXj5nc2g3vUz90gkkUfW+LwC
KzhfjyT/++o3VioGF7CZpQcCQkEjCPBF01Ei6YDGV/5FBYWZoB91Q77Rec+ditUi
RBkSphyt1z2dIC1apj+WFUyrRIC/S0+FPhKd5qTRse5kB1+R3GHF+dnRx/0gbV3T
SftmgtLBC1I/po0PYMewh+/BGbe+9rWaUnUqSVojGc+Zwe+EzZdrZE5T1LnnV8yL
/YmyxBifcA6nwJl6DTUwPCjqOME/h206oxkYPCVUxT9U8fAtUVsLXW5rblKUBZkE
ofpMNn1H+fMkUv6Qk8mXniCExCHeOEekFSm2tFkKsZzOElnR4AfiL6wEb1Z2y0ew
AItb8p+4hujeTnglUQGwyfPn68zHqGi37YXozYLqaFgudscZLfkluGLSVRRPfwVD
jYNwT1evIvAWG/bzSiDOYBq/0cgcELm2OHT73Z/XHtzxEvptxhzLI9vMO7TY9eo5
s3VQZSgR/tFx77ND7SItWtfIxo7HrwtmpNf61YucbayXG5TyYig1ylLdtBI5so8D
o5G+8YIGvvoGwik7DnCMDXtHjXWolPEvBXQDF3icM0+8QZM0u/7a+R8lWxKk4dTJ
GXatRdWL8ZSGazvk/Rq16MrZGFyeQv8jqAiXy4ffUTP3NZfzOBdXbVfd7vQD14ux
4vpGLw2teqDYiCxA7w2ykpcaCPKaV80t2J+H0Fa8rYVHuNKE7xqs38WJEazz5Q04
a2qP8TeyWDZN92zT9up8zwzc45bTNLuSRL9jW1lV8B6jnlLM9eQ5PqtwMb0LLgdd
roelVyWvudpluHqg+t1QxFcM7Q5lRVFWDdxOsaLjDrDeQ6K0XiycIZA+mSII9HUW
FTmWt5qOW9UGKYrsh//y9vUBVbe6bGUBE5B7eIFafYyYk1l04oastaLdOB5Syc07
JELP4oPjssc4AyH1Fpjo2hvowCHNH/qVfYsB8h3mOcrGUznq4auIeKUzHuOf/HRi
Mdl42Ru0mv81nw0IB6sMSsYUGluCaD0mlESeg0CVe/4IA6hMFrNusDtA2li3hI+j
VpxPtOoQrUQn9WLmbK6wpdhbCSswdAcIUph924xvBen/r6kwEkzNIl4744c68P2q
9CHHreWwH12OTxZ2uMfK2E2moI93+YkwiY4IQC5erpjjhczrrjciRPWWXkT/P/nE
QA/TtyDVpdDIjtgbxVQ5OA8/GKZ+o3N8yivqSqN8hHnP9WnnFbELuz0vX63gWUHN
/wQJm+TbWtARai9ahRwoOqFBu79Qqp0BJSFSeqQWCxo7uPCsfbKs/1nBUIACQkEj
60G85CGjcWRFmUft9u3AeCT+hngXEfhVp5QUH3XnBx49RLqWdafsKexZqlkFRuVS
PEmTZv8MTkd1rW68Up9HkETud1DUyfekE1wpk2jPnE9wOi7EBlymbazPCHkFYX0+
0yEcz7eg13/xPNu2hyFFsu4W4a7sXfzKpmBZyMbxUOGQGiO3K+9bnZPbN2JtqSG6
ocxHPMtPvP+RTcsG812DthBSeYvqL66PqJ9YVSYrJTj8CDgismIO27oO+Ve1j4EC
zWKqcoeOVP8JxoFwOk45y/rta8LZT/CsOYOlumLvfu1M7pmWxnOt0BJyldvM0A0x
jM/VFGSGmx27yBxBOrT8DYkrD3z6UdunzMV022ZfW8L0YOfjWSpNMbinCbTMywYI
Tr6XElOY3h7xRNvgrnqgXU0Z5+aVjZqyHxxEF3LqT5rZ0O2rQq/uVzjVEVu5QvMK
Odz0xA8t5EnKr28b9hN+HJglGv+bklfmF+fwg1kyEqjL4MeyepZaGLYSr37nghYK
9VFq08rBbsc6+phMweVXuYpDS5dnUq320ghvHtiiqnBYKcPfAV70jLtw9Vi7CfLj
SnnNhuOB3jBhVtL6aqtd7192/a4072NxJ5E7Naox82DhzUGgwKJSTqY4LuKo6si6
cKhEDe1o+BXU+lytN0ZiUlvP8CQsxQeVpd7/lPFnGtIzjZpxMYZJ9OeOp82qhzmm
eSloxbrCdiNOfdp2QIJ79Z7L12N7q/kzxufuboxjVU3Gm3S437jIfic2aJAkYu7N
mBu+YjVxzBcritaEsWMsYkyGiYwlvqnDQ96dJwVaC1Uycd/Feg5A9WlMH6ZIi1eh
iAZFid2nOB/Mt3lSEpErRZ1wJSJ8yGVjHZsGq979q8kY4obg8QvPjfGyR5jhJKCZ
WR0u9ydVvnHLiLDIScHYccANvkc7oaIFcyd208u8He5FHhNy2iRraHwUptAJbgM9
fZNKaz4v4q7gnoow/YCp1OkNp9f3miNioAhCATAJrSq+DPBTIi84cUVzGnSfdltk
HL4TCswWtNKTkRv0oXvSNYYmh16C4eGmzcr+gQX4pknZ0/xqGlbitC4wf/MT9WYL
88hS6enTy2Rv3lHSWboC6elHDqHs9BlzwPrzQjaDwLf1i+BeD6ccTGacPUjsWX6u
MGUjgQ/etJJa0lnw1bT/JiFEI0OzJwhZ1Bo6RK6xUBKN2rTVoFeC/2z8DYDEboxv
o3WIixfZp4e6lzU1BhIDqNhED9RP99YqYWrziKOuyMNAubpj25R9VoPPM3ACrgMg
d509z1rK98r8tgMc80Zr2YRRFhr0yVZTs0dt7nLmyx+MhoceQ5vQ1tL25yDWPGf+
vyIIGif/p+hAr1SterEq0+zoJWufcadrkUs2A52ZlVlwl1e9gcIZQ7D/iPW04nHp
IU8naCN46LPRVKXiaLJnqLzTmmwOzpV91/BIyIEk5crdUUZDV4wsQA6tJzMELByk
VC1EkGQ7wOfyRjF1rk03ZYaD2Z6g7A34gTCMC8yYii8jvrbRytiWayTwvSO9sVzB
VdupnGxTR/MQE1EGDqAU1PmbqfLkmGTxeMLyq8SCX0/B6WzhEdK/KcoEx2fQSUb/
82c+twE3NyZN/bfRMhauhBu3xTik8fz1ZCkpqnbL8Qdbsh70tV5tLD3MSi/4BCWY
hg9Z6+d4J1B8ANQpvrzV3YQlTDcKo3PPG898m1tOaqWbQ8FnFiqKedV9pZPmlKRt
W3JodeIb3hKJ43tJAgF9ALXSFJ0ZM2uiOz6Ma+lOmMkiXUMQLb4SPcwH+a/HRuDi
k4kpNDSQyg32uhgAeg882BJlYjDjlzs44wR8/Vblodalpl7w0mlH0tFstuXWv2PX
3+mXcTNTiK86Sgzh0GHwENzuYTXjaaI1j6R+2GT9cQ6uRlLz4HAL2Y2/DpF1LZJ/
crqicF2beAr+ukxO388/Qrzv8Uhg45B0jLFoEHQJgZp9t+Yl3EQ142Kv3DHLOtIT
BQZVEokiR3QeFr1AbtGIvICNc5EzZx+ykLJ3fWiZeX/qbO92JGOl0qGzcy/9eKvB
L4pqoarJ8YiZskPiNO0autX4oNROmZT+Mo5MeCXfUsirAlcS0FSt+X4uoDovNmtW
eFnl2RzTxcfexR2soyOnMkDWOMFGnbab+wrcJgKHz7GJwQHi2jhv7OqCjZtthclh
75YT6pveq1ohdyRD9VHmr2ea0yuW3ujEPfx8Wq/+gTLyijGEiv74HzmG6GrOCwPl
JRU9HnU0yRozeAldCHcuW3zmAZwmUhuUbJazb1mmrwFr69tOyJy19bgAJnnHdcKJ
7btc0FElTEEpDtXcxfl7boqm2donrQYzXkRIlhP9t21y99XgZaWV+28Tu/5hb1qo
MrcBzXl6puihk1NF44I2FvD/4qMh0YgVgio6RbuHSTF0a11LPUNGJfNrnEzm45No
c57jR+COqbqo3ObK8yAZ9ENDMCcO2f9Os/0jACNyhMf6269ZoYpyMg+Zzt0mmc8+
3Sp1PbYqHedEOan3vZq1JrKbgDPkwFucqAHvSTIFJEErX2mk1YeCvyHzK+KB3RGS
vdAYcs40DkBKN/wJACWDbWg6s/e2myU1dhV0P8LBe8cvPwSmrKaCSUHV8bRt8czV
pZ/rfhuIaMBM6eWd856Ci/SbrfHeKqK2oUlbnoIpmK1CXPfmEygOeKJTPFeufGms
wCxjxqoR1Rt0xbU59L9G0vQo54zyNhYuh0bFXsxrLDmiSB/3IjIG+jBsZuPZOvuS
dJ46fyg47lOfky0gPth5k5FXrRPE5sjzyu9r6OEjgFzlj7Ur0pdvxk5t92HxorQ5
xrb/UwL5v9fif6YulBhRwHc1jmrk35gjIR7wTuKvwgxNhMM1sRC3AofgkNwB8Tee
ELD6a96OGYT+RERDtUE2Jtp8vcY2q27zTe3wn4HYLonDcJPkmmq3su13pj4H7B1j
DHXvvyer9VZN30oCujCL6nxapJGox1H45637mXVxOtWAt/ABwL2YoLm9V9fmv2AM
w9MMEzJWnQieHECdoQignFY1kh+MgPnMUalAIEuvqogxiqsNaT144lL+6Am62jK4
nawrgcSLPqNYXS7JJuP52ITStlcsIQCT/KAvfzM5tYuJ+0edWVlc3pbq79MLjwXC
Qyw88XhAguo5W8WpNBLlfYfMsauk7wbrefk6RgCuMdwSbXWqFgCf5GIZBppB3sB9
QC2Z2/dHVLFq1bp8MAm4rQVMhKa5RdPCVCqGgk+TCj8LOGp7Ph6T3dz6jOwTtXIN
5S5Rm+j6wGzNGyQ3vS2XMXLmPJGt8RaTFZWFJgiWF0E9x37Nh08Uh57yRSXWElb5
BTFcT5ASakidDqSLg3Uu/a+qCEfpIiMOkesr6V0s6j/HOD2dFvsP/KB07gD6xVFJ
mlEojRvcqWHT0O5mLUCGvZ3bV3rd08rpkCiYxB41a7ZqB4xOIubfF5mmSXgv4uOp
8d38PkK4sw8zZ6Roz7U68ioxnQnVqgypZP6rsdPaVSo9nLMqyKshcS6CbMEQ6Skm
CXtX5HyF01C1M8/RjpGpu9bohvvPbgwxm8BmaRjOnZdFzfhSTATaGv+xNn9/i7xV
DeoxORgxz4O0HCeeQk0eBg7330MhiM4mSwOpJdpb7SaVrsuy3er8sRIIUP4+R4QY
MKJfTA/XmeMsxgU4w3m9pq8Ehfdf/YNGXJkZ7b5lWpSkNzWwZhPgcxYKQd53SEaU
1meSbcQHq/OwGZnCcOkaiQ2R7aQWUCaFwcGAHd+itjs5QvEuG1/GuhwfyBVJECGm
1j9Kh6GpJF+FtNSSU09hCGKdR2u/uaAllZQCKWl8//swGiQae3ZcCjLbSNJeD3XD
3a6UAg3rRh8J9ZVG86gRZ4CrWWLtwuaBFzTr7YaGrnWdtbpFlmM5TZcw1ajanVEG
F/DjRESALYCBEURJm3RmyG9NATKJsipEGxvKE5SI2cMIGiGLJKNMwX8H0zzXSVth
vZGC1s0JU3KyZ0DMHYsC+rfCYoEGOac/zfXOZjXTwVHbyafVsr5qvnDJ7+ghQMpZ
G1VT6LUZTzmz9+t8ARY8hZjHj+tImaOUzyPX11l9CAWur/QLikZAVepSQsfXh8Qh
CSoqMxDCSVDsKgF1ZtDhbdTO4jiGBjNDRrcbWhh79TehmzcuAsRSrO4J13kmBfPW
vyp/KYFVW3a7dIQls5jh8MpjLuQpq4dWX0ehpW37xskAMGYY40IgLruCwGovNfFd
VrQVy5NcQzQ+u3kFKpFIkp5HXJACB+5Dw6Qi6ZwpobCQjUWM4ipjXWK0a7SGcFpO
kWTELKgUbEEqqRI1ZKXqOmcFevOEGhuKbSCof2qhHKfHj/Ync+CsJ9skYlRCPlVR
HsC6VGVxeqhaT4WUAlGdQFhjAAet//U3Im22JgvKIt3fj+9LUpnCf5Inara59PkK
YqPB7y1gzr2SlWMKqgNyDeFI+d5uqZKKDlwkw5z3+/BJFEG4RHtEjcug9AIqmrz+
Gx/liDo3LtVDuRukBrXvpMrwGlIvRWiXfBBkPtCWNnaM3iELqLy44gU4GKhZX/8c
er8MRDds0thlO+m9ERcfgP8BbDPs3er/khk/7xSDVa9UnaUq3CHT3myV5fyX7gLA
kel9cy1ZtqKummgB5uKjBe5C6ew1dzl/cCRxPDdpUayhxflV/eBkgFEzQM87di/x
zmrnhrIs9X3xd5FP7iI7XkSvuw9F0A60uQ2DLEzuTibPeNjV03TRMIbuI/MgCx6w
n/cRVYeg2qeThXVwQR9dWkxzwk9hc0hXJNH0SG2fgAmptkoIgHauSw2SI5fVUlxz
f5cTRB/3Ps6pXlayuT9y4F7b2mqvN6NwEV216lt4y8PGxK82/BWZkIvS0bLchaVz
XWCbLUACRTTmHZzGwGnm2qI2SrYDHwOSTYM18cNrEMOryD8KAtdecARLwoztdX76
sRmh+A7BByHmrf9cqAVqaaMNvqvMM3HwnD3ilLpNg29oChWohWHsZNJB1N13TxKc
KGGDUuMVuxy1xX4s6hHn0lM9lE/GEXf7gGgDSs6ryU/xciaQtDcxurPcKW2/O9pg
fu1ciwu2kw67kw2UZ64qn4m+io/yRnHlOm9o0V1Z8z18Imnv7V01KvNbwVt3E0X4
VocpwfO6BMkgVOb0rGDYoC8CDOjIaZxCqZNY4Wqjq5KwRbOPTnZ3qUT9TcNu4JB/
gbkKw1TrN7AZhKFvwlFWH1J8x9pqRFP9Yro02zIK9oImUxWXDkQ+CzNx1Xg/jtV5
JSkPcQ3+N+wLgLj1YFrR7Ke82eYgoue68aov3bPC77Us23XEel5Z0IAaNE+Psarg
BeecCJ20EdhrH2fNkMj3LS0YCBcfOJJdJAAWVQ6/RajrcQS9BnVxGxQJ+ynkk1vl
3jyxmzz8j30J6e48itZdXvbA+eHWgsadP/fEPvx5LeMYmj9hkrpzPpqGsUPzD8HZ
uQYtfcNy6JWiBogAdtzH0R3qH4IOYp6faLy/5H07+i5vGka7UOw1ttyZAOvGVaWP
e4mY90EqRTNk/5NwftX9YbYsdzKEbNWSF53wf+rbjRaRWVYyEL+gFhk5CHMoK5Ss
VCb6gkeruB6X8nvIHS9Gh8YwawhyoulMezHZ4MIvYNSmlIc2+cSGo/HU/mNyaSwc
jsu7kROKgfRVmyAzT0duhEdLIfQ8ZJoZRGpFAMrUFYdpl0qjML3VDlJJxF14zWkL
J8iDMuhqilu8kEVPNT4/kl0EmCGAEQRlK1ovrmEJN2+fBNYn2T6v0Um8kzYMV8OC
wfGbiU4ZlH3hEg6Gfyhnysk6Vg7jsSew/6plaSW8RPVmwmvR642G6dErPWYPaO5u
+OYvfbytXs6JeWn/RrhU5iBDvcrUBP6eIAPci35dyudV2QgzW4XBMXhiG8KuCqro
WJydjPit3M38foLZo/euDyXq0F9tXk0oRWPMW5d1RzNidK8FHKedk0vyii+Rb0LU
H4pVjzwcThuuatCGSO/vSVbOOr495ujJD7jzjRbt5ckWvng9Zm0PYcs92rb2WfY4
43DDvLwx2FgxNthYTpCWDxd3cjuOsaAiWj03xeQLfzonegeU2GUlY3NZBAiK2fhk
SzfSIYckgaQCkHG8JiC6zWZ1GvB70FH00DmYDgO8vXsfHvXnHEE50IPRcAr9lcNw
xdw1T9irCsL1KdAxmR2aLvbSGpwuixP8nXyo1CcWJWn3F0BixHe6RpO2ht4GEKrL
WHXpY3fDZfpdTM7SJATleOgtq6mx9Awlz/4GOHhbtEoCqqT4E8TTSka5jE+ZpRtG
YoxeNv55qPcAkSpUxzlGm42nG3oZaZzW0CLksQy4yAfYZdhwLk8fa9oe0nxvuBow
teJJ2w9F5GI8mV8g/4N5arjVWNy+32DyI09TNrWupfoHNWK7loUShd89owjVUQ9l
mcre6Bgx4NlBiz3spAe7OJ2x9kV7z4RLrT9alIwP7No4mntb+63MXbI32Wih8R6v
FQ5DfZqjlX6ow0ZCeCe6t/BILkf3cQHIWS8r23t6KhQMwBzEkcEvs6gdC9Ti81Ar
aK31iZrPsRnUTqTCqYQlVWFnRrYFrLqMNBRW9W83VQAQE2Ze13W+ySePmKLoICuu
VyaCXVMWSiyStNPiQUTUImB3avEQQUymls0EtSTDfvQ4cn0mGXGu6bE5RSJ+FT8s
/08kXstecvXgcPGxi+qppnpnXufwIQRGq3KtN61gxKgXQQaXnjxgmG0j7ipvI0qk
taYYMwvktbGy9xIqS56ZQqwL7llXXY2K7gEnLkI2wHwVrFcn4HCrsg5TiKnnrH/6
5EtrOFqovWWaTZlG8bob3ZjG51v5uCBjEEyJ9WpddB5K+ikKN38AhHdjpfVFBiRK
+UBJojU2K2Nf1hTejS8xODLxUTBwmeoGGcyNsEs07aqWA9oDcaRc5QcGtjATTWtB
bTWKPH2xt3DewasQiqWAL/fzYanIttRc56p3JZpiMQeRQoCYQHtw/hm38g5nG8ti
ng7NwH7WCE8J9gwdbwOkRLv0vm+pAXFRF8RQdMgGVK7xc6bqNnP5P8/Rh5t1kGnN
fKkGKPfQJLinqy+JPIk3MNG8PKE8NfsA67zhgltLyEP+qvXA8PD3fUq8NoSE2jZB
OChIoe9vX/JpgKIIb+Htx3oj7DypVD7eoXvrQ0avm4DI5AhN8wV22Mk00nvFcKFS
twF4HFulD4BCDfAcX5vmO7kaH00EnNKJWO9zos9sj+NduSNOJgrRTVVAQtCU7uR6
0u206LZdaGvTZzRfbWBJoNMzTOH+E7/xkF5LETP3wdWd1gT6aqAFR5XvH1lZQSEK
tpPN4HH9A/+X0VZrr3qxCtqs9itjYU6VoVQCfopIh6TuwejEFiWrGYFhL8AOq4aq
iwfCH+ifx/uy6q7IvwYD+V9stVvmbfxIqtqq6dZ+eqG5F3PEMZH0OHXQRlHQrWyW
nLNT7DCGJfyYVsU2kmQr7uNrayBC3ojils+48jLXroWAg0gQ3RKqGzVrlOGQbKu2
xOVh+RVwS2NsSYPnCHUVR3S3YyrhE1YohEkl/QtEurJnBJHYzxvzf+uPkzIsWhAa
KfiDkuFC42dsbtBQdIr0E7+HFxKxx5GGpvEXbhKCfwwA8TZC6NmQ2XJBvIGF/DLi
RV1DB0mZwHUReW6dtDYEQT60jQye73IpWIOtTR4XnGWJiz0DE1cWmF5hiihvYF0p
4CTIn+RQfiZnD+VUqmBIro5VQWT/69zVowBf2PBwwLf7hrruroe398vuTK0F8w+D
Gy+5v0ReMiF43Zy9KjRwhYNeHOlwFcf7HIMErtbQT+sBTfoPmU0Zjd4nenVkuew1
1mb+vwswS4U8GUzZKpPCGGrRQ+vojm5ufe2aES4IcgeGnLEmnGJzuArW94mQLM9f
cbt1Zrv73LKgahIpNnorGtAik0bUhD59tiaRR8h0O9DEHS+dn3uW2hloKMrZxn5Z
nLsmRsNEl0HnYkvIjvtFjzg6lGjAOdFLtmhljdbOdZJzwoTo0NdUwSH8fTAz4LuL
fokRq0Ju9t8ZSNJLvWEeIkXsYQqwPt69nORAWIaDyT32IiDa5PEqe0A7t/C4aFkF
hGERKInPCWnLBLVbTiw24WNl0s/3hlL2Wl/ZbeuMtrHYCF33k/PzXommx5Pu8525
IYuKECWIG3om7DelhYHIqJkM7F1GaMXuWy+0s+ue7iR/NwU33d7veoO61u3Y7qEG
dyiRj2kSAP2YsMEv5yDFi6z9TS2rHNSM44L8ePjbwMSjrNvRiTzHR7ltMGW2jLUK
Tc5Baz2BJgSrsKHMnTOMRyAryGE65YN3Bzl5wNOkkoMSnK6Plb9cwGjFnLGfaHey
qKr1PYf31pgl2org2YVn7JdtxKleEIKFjhL7jWl9UnXQcpWNNBIBbSglEw3q3hwr
RjdnEHp+y4FJPCpZ5FSdGs6Co5gb/f2p0zCm7veBJmYMh6NyD6x3y5ceX1Y30kgz
djnA45wAFSdaHZXK49Ui79z1gSRGpH3Of8T3Ej1Lt05J3WPdUC0xp5KwAtVe7UvZ
Tj37IrjFvCMaFTVJjVyAWwrIMxv3rexnamTcpFs3R8rlgRWi6KGRF3W0t6yAeo3I
8NGPJT95L0zNCgsgt0XLHBQJAGhVzFMpnvZSVIWO8k6mgGBjtXK9ee/bnwbyJIAg
YGfhKhjYBAyq5PKEAfCRTkNonXY0RNoYmPEQanxqRUvXrh2MdprAK4Xzw+HDyyqk
/bGlkZSFUeHa6Q0aSlQEkIppdQVg4Abt6x4NnxePR57pMBhtQc3Hksm05+LtNcLH
C3BvIrHs5P1xdiElL663Oni66B3tcxMKqhtv24RLDaQh8PXAU0TKNKlz53P/7BJH
zuVZrsLnJvB/GFK70HOZ0fwAJ8Qo+cGeafEUZtNEpr30BpqGRyYl713KdtaodtVy
CdrIKZeg04caX2iuAMT3Ir0DOhML5WvlqvPIfxiqmDE7XhuIRJLZnUDpXzbWlsQo
nG18Vvt8dWAgMeBfn+pRAWu9jpOfMpBM1KHAEreTC4Z1bqCPWZcPYvBguCqNlo4L
pE1FRsncDFgKQHgr9LLqIh1EiHTww4v8GAFsoEy6Dq5wRnDXLZIVp6PUnSVnyuWI
z2kGBlWwgJWSh3c8wRE2e1xnzAED6jXV8D5erYM3nnjBhlVU8DIGoD/+NsiP7dXB
CtTrP4hfZ6pmI2A3JGwKA/2uOfRH4MPsLB5EYLT1RzPp98ARPg1zwOx53nJTTFNb
nK9JC+UunYnSOMpFR1Dr1lUVrb3c95ugSZip4VWy3TQ/kD1EHpcfWEecfwTouuzP
qr0HlJDyQhox/RleSqV/TCshIS6ohNc156tN7N5mypD9m+V9kFp/DC+HGuY1FWew
TwZeLZO3xR8Nn4CayfEaQaH29v0FMZGe7gutNcw/jFpi7Wysxl3Tq2h4Dw6HGGr1
po5ag2hMfcg4Bgr+vzKWzz7BJly6P/A0ZBqmq4bLFACh6Dwt1pIqSfhM7JAnvUAP
uvWjT1qQeZe+yNpBB40l+jzBdrbSVZmmIq/4uPz11NVR+rdyQgMyjnuIISi/UKbu
dfrxF6UNNPCYLUj1t1tvmX9Du+x9le5v3x6NFcvIa572dIZg5pD4caNGul8YNujk
3K95xB7u41zvJC8Q/tM/cMehlCiabUoDgG8kdOQXkMs57sm1KtiNTdJ69K1FAAe4
gDbBitZCQZp6Suq2WvmG6GM06OW9W1uEtgmZEBCXvxz0Vhw97BIAd8q5jZimLr7o
B+0OD2vFvytkr8wr+atuh03leZzUXSLLa/SWEc61sld6APps247Dj5L1kznLE4Sb
uzP/pFl4273sgWYcXk7nuDUzUp57fE1msC3eligZF5kwkr/evVxOriy84OEZgyWQ
6bu9EQT2ug6KsXuCv6iaer+3+z/Tgts2Om3vUSNLRw9JxYGruaTd4FgI/Hwvy2xf
RjsdziZyCU1ObmSl2+lqNCd6wVfMQi1BVaALlFtXHYQdE1wN28ydBSkaDnM6vQFb
JVRZ8RyAtaPdAUrTEgkermouu27EJ4zCW+pspfnRqyl45rCGUUeoECRE8cV+avig
DTsib4GFmQuK5aqpbDYHCAOJUgyHZ59fgzEZmf5vqzYPY0tlXLMj94jFWWZeZcEo
mVhsZDd53gwAa/Js6DCsaHMkWo4f7c4X6VDUP+Me3MYAr/pTu6x0tGXmUIXQMQim
96RXhphPrrSiDGJ31Pl/URvOfLP5Zm3s/SvkthQ/Iyp6d+Ewm2jvOsWwDLJzYRZp
J0PBWw/JQRTDPj3fqU7sMna1W1TovmXB7pwMK9bu1NzbmONMCTlYvjBaMb0lCvCH
RdsLV84KQVMSFQAUKqjYzCI4bIxcJOmMfKn5Xme0pjSNbHHQLsy/XEceBL1pP1Cb
3+chxAqv+JTlTyHqQPmN3PNkfy6FV/PdXUHdxFagwOJuag9+Nt53Dibzzceu9ioZ
jdtT+3dF6CI+yKK5grLLLq+Np7k8rvipouozaTkeMFu0nVuGKEL3SftO74x0Cmat
vwQM77KCxHHLbh3EH0EzLd+btRcTmbrsW59086nlPTTtGtOyIXDbwzZhsoJQ2oK9
ZBl67XB2C7rqXRdGQh2GG4LnH2YOEwS1W3F0FF/WfLRYBHVmJD9YaiWXuiCQKQ55
lO8lWUtNj0/Wj7cIGKuUfx5fIEeUnnY05ICPrk7crsRFLF48WK0DriAoZGdbRfIk
xaB5qOUgObR3WmlHGRnGvPvZnSf5pqFFKWW1+6hdEAAwZPAQzJKL28q/MUpbfl8E
2dhna+bHQJQHOEPlfZvqxTH5Wcodv4Uk1GOgfLXNkrmTcZF0kCDLrKL39LDJ5yze
HGk26XL/3zhtKKNJHiSvz0PQItYo/K4iWK2PCALon8yzpnbawkh0ApAZqPmsy2uZ
cY4fUhVUQrNwZAuRK/J47lCeefRmJcZW3mPqIbYdkT998gxI/Mjf9TBluCj4ypNw
RL4WisI1Rfq4pZWfXWamDWrbBCHPVl+SXcimVznRE8zlfoMTKNc9196dNzafan1B
hyeq6IoFe+hIL/Xe4yoy/wfpU4FPcRwF1nipbb3+ZuArW/nb7OQQDwjwde76+1US
/ER5zD9h2lM3Eg6i0gr/4gYdd8dRv9ytJB2cbG7SaQomHz0C9fKkEBKWvl6VRiI2
j9WJroccKBMBmZBlw6ew/C7ErR5GtFKKsJgGKh+BkERwNr9tLjkY0JcSUnm5NoxR
7rcumPLYW7xU6HnAAQc0BNjT5vRqGiKujWbToQU8+3WqZYzHLjYlREJh+iREbt+M
7F8XfgUUPog0JGThS8gqxVkhJwKyknRa8UaE92KVHMyqKMfBXozD3uVbFn7g68Kn
PtgFc1kTqEtt/PjB2V7I1RuHUn8mW2CKyOqCDD+mJaUrDyXcoxi8sF8t4EB6IKU6
phfUu/iAn21XHXEZ63kaJlJWSzuy+a8jSSc/VNlxrXsvct2hgsVtWDREcT6c+2XC
Ni9lh7W5VE/0Llr9U94YE8yZOSPTaPlqJ9ciXakGBFZY0/4HMoi05JHtRqI/V7Sd
6SjFKCxbWp42uvRAxwLOm2jn3SbYdkTIF24EqGcHG2CmamEl1m9ROBvCLpfnSXKd
jidx+0ffyaPs6iSGipMxptXG5HUQd92CAsr94DWJckrWPgepjBpOA9xeYdcVZJcR
dbSlF7y1b9um7+tzTbYWzC4/xwaJdUCS/f7BV28P8rG0g0VedfMfmqeFTVm72vN+
/YLKgrCVxmbNt4DCezivfnyKw2uDtQ7PayAK5mVbsuN7Lc0wK7U29r6GHDu/eaq3
edBPglaNWjXFdB7lpihfuN0C/mAsHwbJ7Bc9pgm0qyoTMfiHmBqOSsq/LNLe1YXB
Yu2Kyp90l9MvdG0IWnMcPJUr6lbHH+gnO5V5Y6WYLp4LU5f7rGPyl0b1/5y2B7ZE
qpq9lzuP2lwkVDewqanSojxJ0UySGP+lV1sA0LpCFuakewADeahq9+BG3doJaxey
GOYJa0DU2qTsXcO4iE7PE0cRIRhKl9hwKt8Mi04YiYEES2o8wXWrOvclGRYD7Eq5
UYXGB6WGB9S1AKRu3zYHFGDDR0i45TB75OF/r11UhHKr19rcnL0pEj8x99xkA6Rp
LKPpwXBlUbfPEp24AjiByXiP61oHY4h4vayftWkDFBEDs9DvHk6tayDHqHpuf5Ws
kgsxWdgZoUOTF1WOGzCIu2hlLbauWwbQYWka9zlg/x4WB1EybcmLVbjoP6TY0/QW
Isa5Qkjp8L/nvs52G8xhzh8Js03y47j/drBODHHyK+n9XQPaG06JxiYsKPWPibxb
MB+n0cIr2NRxzVZ2kAZC7zd+/R7/jklbqNkbBUZ0ujCWsAszmwoxnAhDCIK7IS/5
pIuYinJ/XMlzPVV5II/zLa9KbjLASequEIYkRvKJPhJL4/TopD00jEOTi6Tudb3G
/4Pr5lkyKUsu42TbkoE4l+maW9zH/9yet+HmqYIDGZQF0k+EehDGJZb3B5lfgm+g
0qQqu9KGW7BgBDCnsPXeWfimaITyyjLYd/It6snddrf7DLaXOG7Qc4Q/KmqHZijK
/eQW9OvSWi+ZLKj57ieE/jWKaLxFOA4DV7VZfbR90R7wFWqXjCbGDzu+77F7Nnhw
Dkru3FL0u8xwif+vcorHx6kHBFJykX7noSYfEB4jt3dOBKm8yZyfwsMWn4N0Pmfe
oD4T0S/8a3SIpCn7Cw/DBhzR5q7d07B+HSkBbGIz9mKWH5HgzMi9h2/fdW88Ct+s
W76F/79iujPboVrosVSyPy7yS5liUD7diJRCJc0nEVO4EL4trlaAFwC+RiZUEnsN
W2a/yRqeZf5eb9SrF6ikTI1NWlE/riUpMBkdHqhTXDsWTpP3jWF1C2UJsll9g1hf
eYcFysiNugysRawqlK8tSlRrGFTFQ/InPDSRRvJKM7VFvEWEy4icQ1jhT4KA0TFH
oSMw6cuopvnBJrk4GsoeCck8T87iA8lpusGzY6W4RAyO9nL6otdixhRhrUpelcbZ
a3HaoQoad6gorFcDJo+X2KQ/kDJ61sbZ9Z6Gy7ekp6XXqlAbfRjlUXdnQS1y+aHe
+701nGxF9u/X73gFTaRb0rKeaunl7QWEIVGK/wBMdNokufQ0Z6rJD0xQ6INi6ZQk
DudiKo7mbvvH/wQJb9qg65Y/XicW0howoTv8nzWufW/wHb0O1OEyLZzKsonK6MGZ
sIoG1kwCq7sD72UuQXcMlau2sitnCtkpWKNhWkneNfEw3NEh3uIdCbL9INlQ21jq
MHWgOefK+rFYIENT+ypplp8owCW4It+DoLVN/6KXmgCbw5K/06mKoQ3vA/6HyKmV
S2gIhvw7e1O5ZnM/TEPAs9S+tawqvzd1iZJPgYQXAWX+I/lsfQJ3LTCB3T3FKPeX
NLrourypHHqSKd983m1jIDs9qyOqtPysBwOmWqq6hHj8vLnMD2NP7xD8qswSvtNi
9Mn1yppMQWWuPEGHzjSpTyZWc0TGmaHjm/klOoWPCeLmklRfhNkdhiFdIQvoNz6E
skM+IirYI22nugs194i5tOjPDLkoDTye9PctUWgVZ5h0o2bEdMBYDY4X+HMTufwW
2JrijV8CgA40scj4hNRtzG3u5/Hzo05qFbjGLzDXZA5PrRC9bIttiU5IQ/k1nxp7
JfgWSR7yODbEDPifghn+KSdGy8rfM4uep+iwVNchndhtJaGhcJJzOwn7C/iNYksr
cVRblZcnu+6mu5ymEgpse19+t30hDTDq0zdaR3i3YvOh/Bxy0WxUhTAZuV9fHene
RsvH2cL5BhNDgZ+n0xe6IX5uIszqWvwBSPs+5+1e32R3vA2joH+w4G4msv8xn3/y
9C+FU0ASysUDCDF8z2GZmUME+Jn1lBYeSc2GMw0z+kqXfUAZjFRr/e31T3yiLeLJ
O694bxGI3A2TF1DFXCpQbi4/oVLbggif7VSShd6fjHk6P4w4MWdMgkrraWkIhdbj
UdQju0M5X0bbPrf2/IVlalmXCUQxOKVJpV/DWmuRIZa2vXulAV1mQRMdEFm2fsja
6n6aHDYM0PTQ0AIUBFAnVBQGQ+JqlQmM4nDI+XCw1RJRGJy7917OKijX+Ad6UJyc
89d7qi/j1pUWUE4s0YhDnznOw4KXPnd4cfaSeK7xGcY5Q0SoPdsc00fenl4+8OQD
xQ+bnNLnOcKUqB0TdeUA9JyVilNWSNLPJIXwi934iZTJPhBTnDHwQIKvnt5VVIQP
lOgm1I63B1/e4HVgbcIZc/ag7OKQQbjutsVEnLOv02FGE2BwlodIlVRF91+XNET/
8DgaXDEfoaz3uu1gbiZ+lCzS7F1KedX3P1AQauusWLUErpHqXPTQ7rF4XnSg8Hb8
KhOSP6/WzHyx1TyZ3ihCEO3JSlaPl3JVadkdYX5hH0govIOHvSm/iQ+gIRx0t+1G
yvcrbD46zgAa2NbPE8DNq3ZJWZD1l3Xq031ceB2YOjFJjqXRqvTZk/ALkD0/revT
Noh3BvZXNCoaxfT4MWC2eGVaxaJSFxLn8MesoObvL1oXhgXiNulo9dWQ5JM0r//7
/wPgcCii3bI4D4/4n6cPmlzc7lBxJhrbBuQa5fVQ5DR7JUXo+7stF218kv3i16SQ
LiuXOC4gtbKwLrWcQjZBNOgHm1zxR7Bz516oai9/OOlVWGFL4y8OtvQqjJz/1Twb
eS7KXVh7z21MxCzm4BfGqu/wKuFqmGGQPCGpA4IyOq6eAMsPFFqzPdMoo+LEJBjn
IKI6ErhCHFmstW5VJjcDyKZsM4AFSsHFTUlFeKbBN9JeBo8NPo4c+EPLBfzGmsie
iLAMQnpoGe6I1TwfbxUR2e5YYqlZFmKYPUlEonlxxilmhLa+srRvS179xuR65U11
rtWU7oDa7lUWPWRl4qpJlNM8eUdUbqzlRSewuFrnzh00nY4PR2U33SDSk7ZpU/cw
tTREM2tOMbZXAdPbNJYqK8xrddp9o8vPEHX52cigI2hF3csguW+RUEbbXt47rZHL
tYxuVps2JODolsi7sXD0eZU8PmJdtbkh7IvXs2njry+CF/WN+mm4/toJE/xCwVlT
QaWDJvQyXHPK0P2v8B87AsrwbrcN5oXdOm+G/Ky8Wi6YACBJCdxjJvzANVhUBN/Y
Ys+BS8qz6U5BD7ehWwfJ0Vayip5NBaUiR7HI0hndQVJsqrQ32YjCKUKcO02msn0a
IDyVJsG52PTVOX9VPOeMtCwtNJytHt8f/gLr4dOCdshBBaMwwJ1VH1K06G5mvbYk
4sSAbvMlTpattMdj6ea1zo1xvSJinELP8T2K6PFfcdqWMSi7Aie0F7KPmMnpa9bk
hjpy1hq0XtyQkIk4N3xIXrPVAdGxeJE+xH6dOQ+VHCiLp0oQeyZPzxCYT/jgE1bn
8NUlKyPe8yKWHkQTUWHdMU3Ey9MIeUJYSPx2WgEWHwHn5LXgHSccwq/v6q56eNBU
mNuKPkfc4IEXHfRW4T3JyMECMVFeExC0qvu57SJTEFBzIHKXD32BLFxvNPMQpL5w
5gLp7DygCUOlckLlfpeD/rFOUikGW5qpbymjps84kte6FSWkwWKUiau95NTMVjCp
1lJY1dCfYMKm/NjVhERVuC65dJ2s/AWqu23q/eAWsUVdVGtLSMh3IuqzMTOLgQAR
7eyYAzSE2vnxB58UlStr8V4cL6gi1X7WguDYmJmp7aIxGT8J4KG0+O92Q7bhr3hX
+Y5XcxCU9IMYZcoGpGwryOI3UtxNyOZ1CCd/LPVmKTo9ZQcqQphFuunFwz3ekTgY
yhj8NGgs01ykKt1mZyAHkcGmFyCdQhQWsicTKcO7y3jsNlNVBf4yMyoScmJ3kg6H
qb/oqqNE/lUNH1DddALbs7kDWGipOeLekhtoEk/YCaenAs6OmXjlWFdf8635LeEC
vv8+/z7bybi/aJoOWjW49r6hCsid+czYeFMeXUxXN2zKSO6dmBYzlMDfTYIaTsqz
gMCYvqFJsfNHpFXCsWoLct+BtNSiwlGC1WBwfkLlH/KSkgVTAlp1aY8Gaa1yV7ce
H5Mnx9LgGuhbfCJKDElgaFReb/osjKD16DJfHf6UJpUdDEVjVamSjwfQ9MziEjjb
gTbGCWggxegpg7P0UfLlzFqlTcwxTv4uPs2lDXpzjedE5+oDwML9bHepA9H9m0r4
//qMGSa3B5k4sGk21dbzo6Z8wdMcAirrcyFsolTpCV61T0ULOSRgjae6tM4N4G64
8sPz7+eGoEeLUMyXoZqXvy24z7w0V1KO600DEWs8IhmafFCxSppEPc+8+HdJmYvJ
7e9zx/JlBnPNwDTH3ZMvEYHiYPH1JPt4JvDfEVmw1Q5m1ytSPeM8FD6K0wBuIRsb
u1R48Ii31Lq5KlFb6eq1W7tSHve/Jqztw7wubCY1fLLvgPIKGnQ+zpxVz8boleb+
WuRMzFELRFqLoOz198OansQuJyIcVhwF0v7CZMUA77GCHzYIhbs4a6YoMcqZgF4L
i3WTFKfOZO6TS+BcLsjekp6K4zUpIAvJhBq4YJ6z9DGFQjRiZp42dpaFN1P1VMTm
DggXn6F2iOP6+If6PajxbOnv8gp49Nqogb+SA399J+ofJzlAYvYqd69G6pM8WDm7
TORPVw4A1DQ8bV4UjO0wn/uSNl5QLx9D+F4pR9GQhM/AndRp4nd/0NLI8EB18HNn
G+CIVR7wKXTZoj8v7OvO69oza5/IX4KFfr/sQL0rl/RTUFX3kQ9OC6fufP7psq+1
+zTofmigmeHJp05GonA2d4PuF8U96v+NHQ2wRhTcN7CYbUJzWPmZynqwdjjqpvMy
1QBVE4A+HwtoeSdxvXxqmD+GMBhiSR/+3HCoZt4OnHNa1TvbRbzuRaSca30jYzk6
eJgX+UTuOfhmwO2CV2QrVFXfuUtIbNO3S1FrwKgTNXZ5f3JvKToXmsbWnYVicGIk
5XlLLyU7eEoXEgXgEvfqWg+feL64/NgFgo4pllSx9khoaeQquSBbZi+AnvJUToF3
5tWr72zLEFHp5gV/1jhq8CoWfosQrzD9jzc34ByQo9QdC/JaChbSU4O5da5g9cUi
B2t0ABvOdjh9Bo4iv39TVYGXo3O0oJAycSWj7OZMlrxYJr5cvq8yYPZHEs2tvm1P
qlieni1DmX8jsix0LkVOx8m431H/S0iJSi+ipWCb//0xK/QOHv0Z3kwfAVoKAYTM
4nVeOcgRZNv/ClaWkWgNtSAx+uB2Vjk62smXGAtqY6M8A/DZ5hllHJEnccB4H5tJ
OwLcGOtUvikeVtl6bkxa73K0lAyf5kSwH6N2RXuDMxiE7+78pkYEAIfOi4+taaog
632aDRH9KQOg04fh1DZ2kf0L4VqCD6iT7dgPKEF3yiyFk3Lqa3rGxOpSDqjtpxzN
2RWpkCtWG8aUMb5v/VU45fRWUfzKJooaoD1tGJnxvwaY/EyBfLnpg4GYjczsbTE8
i8GEDaRyBMaRgJVI3N3hPfOCo5sBiTKu2byE9i9sz1eXzV305OxbFetxu+N1uJOI
XEKkwBTcr0mjsCbKcTsxPucypkUST1XH7OUZoSdAo+yGUg++tgpRUe2Ky+tq9dvX
6aGZpepZ2t/mfkkKj2D0Hkaf74akmoSyF+bwXQSr0BGcGnFK1RWIbPy1sXGZdE+k
OpL+DshCpG0K7b35qYGLS6nu7tQ5V8QO1CLimug/k/52Wbi48+DaoaP7TEtI0CfA
FEVbdiGXirr9Hg0quG2nIihX8eJduVaxzQaZka+kfZQJI/aYxnQHeIQz2NAFxzP6
zT3qIabkui+xmBNS2s4nrroTMgMFjoUSAgHQbY9fGnQWj52xFmuG/rvzo6Ybzgy6
+cRWCAvdXHsZT1cnFuPre2kbgNd6PQp4RDlTFCHchXEPXAzuVJDN9bxSUrpWhgw2
UEkVx4/KnZy/atzmyGtvIHcSaEV+el7VU0ze+OXI0NMzVnG+dU0ZAaPOI3ptOQYT
gtFPPV5pKCj0vtLIVltweZ9wk4JVb/zDUTA/AAtUEaZIhaCu86IWoSlfuLtRIT+K
YbVd5XBbpBCiJrcyXtbtNCO98SEAOwzc4gxrnImkqlCNyzq5kY5ElMfjCYepcUvP
BvK0i6u0A2V1qkKI2zZVw8WoivDUXXZuD1g9tvhXQ4D7AkhV/nD4O4hEDaoUkALO
AWbkuu0N1yR4Ao0hUKJqxVfI9Clb8bst9BeGEkZ0Dh6ws8SMLkTZfc8P3L9JSNhQ
cNNLlig+9i0XfDMpWpO4xsh/4wW1f5GoYgrk8+1iBvKFYh+bcjHI0esZUcixAI1U
RfSJdr8CfU4+H+aw5tTWnBoH3dp4b8Wei+4Sam/1J0ee3e33abRQSN2xeBWxjSCD
ylSFzBrhcZ8Girmajf+HlQYT+uTL5klYzJ+sBarz54C0vZjQoJQHsUG4RWcUr+bY
D0LM6mx6Yw6+KVaGwmNudGyZv24DyovpzoMKFAedKSBWeCk/8YaZsrbUnPnmb76V
izLyVhvC/G5BFBbRq2C/iR+hh89nWC5pO7U/rfyFAGkupEkedIGb30z/bhn1Pf5c
fazN695gRAFIDeRqsjZPDNAs6z0zFxAQYlH1Ly+HYG8Zs+xi6eLLJ4u1P5AgAxqD
Rl9/tTByM7KEbgnl5eXlUaWXiKmEPRz3mYSUXmePRHn4jqWV159LhvvSEBL3Z8IU
5lJe8ZA0dqw8yQ8rAbDEJZ3GI/+qZulQhg5iDDNCzWqz6jYTZzL2OTJ72pTu0YWN
N3kGkjF5WkF987DxQEKVFC5e78A0Vv5dilUXrGEagtAf34rJppAbZluHviDBW/Io
rH4IRMQengeJ2aRfBBEBO0AYbjw16odv43JCTt0Atj6wiiUx0ntd3Uq5Ky+BF+g/
qQni2kZnO8Yib/ldYXoVTlA0jDHfjf6OyWGNGoLKpzdwqZPSMguUHjCJ1HbfcH1l
MXl+DugvUuAjGecrrjcGS14lI4OKvgyvA9BY/VkEXgexy3xWG+7YOLeNvXdU6Hrr
90wLembNs5OBs2IctZ9DOPetrVeihl5rcGqing5rD6dO06kWiLh05pyw56lYX2SA
864c23ZZ9xuXaLyJ0i7eIg0dWwWzqYh91gHPNhA0nzTgr5LnuULrRwrvffuWI1l1
oKRLa/nHYaVxt7LQeggFde0jmCaeCW/MHYfAkdLrvHkT9uQ/NIp+PosybHdS3RQy
HYK1CAhBL9bvQytupHCn8x+d7+1geHFtFZ5H3N5qI4ix5sTtZl8enEsQ544XdofR
W3N9H38/H8E3uXbhtpyh2v7z4hBybEJGspA2LARYa/r+t65UaLubtT2Us1nX5aib
AymY8rBlMJ7jGjizADUFCwvIq3SbJxtGoYnFi3vrjVMBakBvko9Djpk3NdsijhDj
88RYS+UbmZ9xJ0g7QmCD/sZ0C2EjyWiMX1sq9HePjVqj8xsNFnouKUHfhSXXjSrX
kkge6Ek8SCaonEB7/YZy1KpDBW8SZ4qcUuMGJ4gKI2FbnAWYCx/bE+psZyuP4TYX
wH/hQs2guenmZ1vhYYWKYDS3sEuEoEP6ICQYGJ59LE0ZpXpmallUaG8icayckWN7
RfYiP2Ng3O5ghA0IYLfoOKpcfa4FyUfiW3TL7DjL5foz8TN9s+uy3YTLPYKN2pCs
3wL/4vMRVxDRCa3YXoa1/zgjkKnijGiyzIQV4iIi3vStJW3b6+trNraYsa/GyO/f
oE14+6SylySjxxrnqzbM8I+c2wwNXN5RRyoO4J94/NslMlCbjNQQGB21Y9bQItlJ
JfYCvYJtlcKsSTFXVn09QbJ3u2383ZI1jDITk5qnuRL8WvOjOd4g3KDIa6NqtlFv
bkLwEu0sIjnIgXFdp2/8umik/Wp9TS2dPocqv0bh1v+3buyHK4s7Y1PGqTfTNJgf
v3EUOpxT85OdYsKv7p9yJ3CGQttytiqEIoilZ3l8ZCIahMLmfO7hyKn8tEwcoko8
wf335hTEb6dnlu8JYqzWb9+KvDCNV8/E2wcJBozwAVVpeQjUC6eF0CF7UJbYQ8ZI
BcYk1V1wIvPi+tVH184H5o/pqhQss3REYxUcuwzLVHdokuLtXMTYMGO+5TGt8l7l
9REiCK9ke4l8nv5bIGlF7YXtfKNUiDexfYbo4MtiXVPgvtVbEkvfmrfEukqAmU3D
6mGWgvRZWag0Njwu3B8LJIYJdcXVFGG3QJQjz9U9kFO9IQ0nCs5sXR6frIPersnf
ZmsKRlCbaCfCcoN7Gnzt6zJDSescuHOj2I2Bh+f0GMQB3UIlBTyh8wtwe1pNn8gd
fyyu4oZofRZuDQW9mCuk5nwF7rXPtLysTSawWFEzCrmnEzaxPy+wNAZINAD4Lq4f
Gu56eNt4DmeIImmiGsjvHV6iKHk2EfQAd/KByuDCPg5mNr5QIE23/X5mXIj4hMid
RNyhiJkiUWVujcpEFLzhQpWrWcxrcRFgOw5C+GTzJonDYxT1xdzhEfzUfPLt12fq
YWlbPq0Kpb35emz9EnnD+YimoF3MDcVcujuBT1UUsjKYnfLkn5eduztGF6Gt2D2c
fzGnmJM93IGxwgegOWGXicnSUuZJFpPQ5GYnEc2fIN2bSdvUTTRkxSZAH1dNNXMh
Dr+bEeHklv3pqgauUiJh7FrAJVSwXbqp2SKO37jaK/pCYZWaUwcOv6JofLmPRtC+
v3Zem1r1XyIw/kUPYtiHH3CEuVxvYCd02fXRDNrYEY6rTTdax+VXMs+7jnVBKfwq
s5mYASI23IJ7SLWMNitF56T6epYPbMwy//e43DX+wJIG0qVK9QF8Or2CuYijgMiv
EEXuH0CfcypqFL4qGQHuCMAgGDJRL0QlubbqCgy7trVULWL8XLstL9E5l0OB5VKC
p3reRS7Qsxva3aL63gN253DNlxIjLIZSA4mBR3jYSLOnSfNjF+pydIoG/TO2ggNO
ugBcM3Gg3Z9nfnTIWQf0V6MQz94rCt8L6547Gevj2zSI9oR6wctT2AVRyhL8M/PU
kPjBTXevro6Zhl75y/XYQrOm3TbRefTzdtWKBlSH9d8xZKU74Tz3GWV5LIu61ahu
8y01kokNzsrba7SBdJYaOAnGlJ0yQ5SXFZbRXmRz042FXZlhgSra4/e9SJl5CANz
wOhig4WQ03eS7qHfBHh/GXcVhWk65Z/7xeBRS69V01SIIWtwfTjwyNg43Tn4cnIY
RO1GZd0FxaYF8ZJMhpIjX4xnl859Vl3xQx8zA+L6ICtdSa+pO2o+mQPCZQVAqbwg
g/w89Ja5Go8Pbw+tQc2sPMFVdB7VefN0bP8BORkOlLmvy2zYHXE8sIMQnaHnUc3C
MpWGtmbMAJd40+hrArjbttqhZ+d7/WwASlAqgCIHOdj6VV6LjBD6dQVZQueaMVwb
DGc84ro3fcJAR6COlhTw2WK6J84aysiOg01VlN7I2G5JW6drZpYkJ28cYQXNsj86
9eRwq601JzTJRleCR6yBmI9hxP8+1IC2cksrsVGyVeS2pQEWPWQhTZYVZyF5Kla3
Xy3RHnviuuxBDugjJZUV9Y0D0H6NaiRoxz2rafON/w9/E5QyOyOdnQG+aKIuouCd
7SStse7WjWrJio3UUQ+Zc6lUquaoym7vPG26egCK8Rh5wkS2dgkJmcxCQDS2zFBU
o2RGNHq+wVuY/crPIFwvTkIA1ETTb11M53joPYbOKMaPvpcnC798x9qrob5ldIIx
V7tiE1j4yz//S0qBYiO/LnvY3yy1CJUidEWoeUv1cd+HhjDZZP9e7fQTieI1X+6/
6dAdmZFS7qbwB6DSUV992uHa+Vp6nhtaL6TN6c5ONGw7UplJZ+IcKCTOcGRsCUn8
iarY/PiAHC7jnpjzw8yiKenhnHaapTDwVqmXtNynJxEWJW0o32SlY5mafuyASbey
NjlYn9JuCUuMMO/ShUhnTtIGfmDwNWMgbUwZZjNoHRILtnXK3SRygKMbBJsj4uS2
6GExHySxBbhSFp2qMWEySM3xlFX3NcWXVE3JtTXmxYP2m6hZNY3/iIfvbmlZuJYE
YA97pb8tT9VR3ATlZPgpoJfcFMZjGtjeg8+J8UyoWvCmfuPeeCSTuTrv4UyPY6gP
2NrwfYnt5xddXe44gtSY/Vyn+OiIU37RV8BMZmpZP8qq/jlGGRXmKGFOBgkRBFvn
sdkXYwxKALC3Uc4dVFsL6kZXO+udzKKGfR2Oyi2uvN8WRi3HhvHoZp7scX6ZGePN
bTMvuJcPOlb3DlWhPrwGL4SvvAUHi2CrR6JDrKe569tZ4TkT8gkegVdJBke2B+/s
ifK3cPLEFGH0YeFR0i9YZ+rPRQG21x/e8sAvOd6ezTUJmZpbQaPIH0ugcZi37ett
QJ/v6kDBOIm3iVboR5LvybxiiUmg/w+9nVRmm5LuAWM0VsJg9M3GPszJWn/JfLG0
5NR4FCQiMsdz/qHomXv2ar1RKPN4HCF8kiX0yEclzNDaqMut82KCthEFl9X7zliB
+WC27vxCkZ94OXgzdBFeOwW0iulYB+6NdlEKLBOwFUKrz5Mreo8zquskQcNWlpnk
hXKUhXZ9BZFl8voJ9QoKRA4Y9KfgZNN0EvkRLAiZWwVgAN7ue2/RKKGkxP72rzll
/gCZuKz6rm6ffsxcowiq6DdyjDJimE1WsATV1RHHxiznujg39PD5uvOT5hJvDvAx
cbsiw1BGZ/jXyr2KC8bJsoLezGigny3kMovcAEOk5J7rrVZqsqQXM2GYsc/vbwiD
IISJ76lm4V490aIU4fH+eGdz00bD8kZyHSOmloXUU7uvXfVo9mRBxj3sHJR7hBRX
R13RfbL3quVSDpdAeBShMrxHsViPeTkJMR9L39nPBxNwJxlg7lZX6sVtUJxyE0I+
Wr2O1mJNLRG1mEfH67fx7qK9ynVNWwxkebc+Vs1fetcbXO1DkdZe/TpI2Vt2Kkcn
jV1ZGqaYr2/MgkGaCM3isT/1yPNd+XHrt2Mtq71oQ1kn/ybAZWx5vY2rqeG0l1X/
hbzburRRIf55VflejcJ6eRNdFVVMhjcfDx7//OzyvoEw2Q+3IvlL7vf1oT7sL/W6
OrUh5QKTZfuDXrnSaegydtN6fzp7g4wJniXca7ziMEh03BuaRObLwMSa9YRt1GAJ
TIY1JjaIqMrV5ZNsEe7PdkfNFYPRFpvn3c25/bF5L9P9Nqy66SYJoNhhDB0FRhDw
JZtqcP/JuAxIMf/wfXBJ80WMLL8hoRH22+Pfmypkc9Bdg7XdbssSEG9MZeTyBjZh
UflZvkABefnidaBnQYugRHlm4Y8R/c2Xj8LkoYhC4E+Pd6xejCZP+hPtP2JoAn+x
iouYcibmEEbgYYPTfkLEPGY+qFCweAFiDt5wdJQZMKVTIegt6NJowMFD+JrLa5bN
iVE8FVmWugnnLUrHxmAxqge6yhLFRZVYNqIbIXQq9a4s9WUSGw9Ej31M65tP3wDv
mhJxtib91aNYoIYLhmzJo+SBgqIHK4VXNE9QfTGK+Synh0XRc0Ei0NAbNVqXI5jn
bPOHCkNu698BQ1NLQqgj5t0ItoX7EtNwUzwbcb+SpZRt2IzUbhoHl3l9RGsgLfVy
oFUOvDfA8RCNRqMkTtiQIXowvknkT7e+8VauHxPByO1MPaxdvDCsEXrT7r38qE1G
1OOUpybzLrsNaMvlhiMgaVT6XGw8DFYyYo5q2Hvy7y3foVQcrAwJKu7fmIP2Ym53
Cu8qSj+4fGoMTe5QlUEUXPTh1QECyC6SyIQxxE0FfPvk+OjbU2eTsagWS8C6x7kO
dp75U2hhUGlouy+V62Z9iEnQqRwGqW+AiZo6XlkzJoxntSOO2LzLwzPqkgZpu4qb
Dc/d7tP8l707Nnmt4ZdBpQMnlnfE+n00SITK/NkR0m3zpTziIzoG5r57Te5X2BCC
JzQVNK8cvtLobOAizm3gFmTqyVPsZYjFF349jE7JW3SfMSt4+IyHBdefAAYp4l/p
wWQd4BE0i1aCM2G5ruwr+e8S2sgorlEmQRXhAhBTb2WN61HksL0pZaTMk4WIgcw+
r4nFYFKdMjNd5oyJLtHvg/QAlmgM00sUeNLRiVToMVc1KFQd7MTQgLz7WuplcGlo
cF3NYl4ECBHRWBabj35FqOFVP5wuw3WabkMsM8haWC+yscEyhfKQucO3ARTe1qU2
quvUhMdOYtC3n9xgLO4qsUhR6zp59/UdSnqglyboaMuQHeGqCFxuH3LxdKaYUoJ3
mEfuiI5N7Q54njTGTeGvxoJ9vBDrdD2VaSoJaVs8mOG0vxQ3ksvFMAJuriRZKr+P
9a60Rr8oV5qHahcQnJtD0P4Vxn72zq8T8LOFVtu9y/iE9htFwjWIu8ey4PbcF3i6
k1xlTwUziSq0BPmAwfteIhKA9vxUdK+ReftiFXUToRfm/YKfQmSvSbFV+QNKWSCf
vpx6kX8vrXreuTmO7dk3cWOfp4sVdmm50mN8vjulWrO+qxhO6R2yiCfANHMu6PwI
5bXZhZF98UOIDbywjCZgpJQNBc320gE8i4ROblxDPP5tveYf/xGmzZEDiseiAcNM
tb64PyauIqPhRA8exKFlT3QVqXVoXHZ/xFE+U+JZP0cL1lnkvBvSHFPSrb+N29yr
GrngKfvA77QY1OhHpxJWlEJrZjjtNcUGjBld6kNOsygIbUWIVKaxkzRSJgVXkMaL
dTSEFAYho19PwvQ1yr6HKsqfMFblkSeH05xbchsGo4eeG5OmONcErs58waIn6ZBF
QTktzKBPBItpvxghcXBwv7Scfdx2Pfn0rKr68/T48joxb6KfShaNZ/ib9dP4uj9O
jmjv+3QsfWLJ0FChYGpC1XZVw2bQHvQio94e1daAEtd2DG/X7BIaAnz9bx4donrn
xKkSSKsSDMz8sHz28SK+m4dKXPUa6nsuQM+X5M/abpM2p7KfwuHbIdmZRpW9ipJr
XF46vaN1j2HbzUo1eb8EdhgoDXdAOzCHvBUS+O+b5i+6AS4GLRWUyogCL6fy4sJF
nNTvIlfWs0bf12Y+QfICnJxQyoM3kXsOoEKCQeXn0iXCd1DV4B772nNZvBpVDeXY
AJCdX/10MrfTYFDCuAMTEAwUPuEBpMGkLGp4EBXS8STEzORjv/FdXqj5E65iS5Ur
tdtsIOjaWrgnSqO6OsjOzBKRLPOIGG3Ij34+SuMXWLgKlLblFZutX3wOyXeqxaZb
dQHk2o7EsY+TQl31QiEMEjPPmxr6ZtkSd9pR6NF/H4GQxuym51Jh6F7TkAg+D5mo
hk+1SDH+4bER6728z2kbt6yixv5uCovXaJcqt8gnBN6EMFmNZHs/WkqnWPLhNiRC
Hq9+B5pAvVQM09AXLlAMgmj+6GWvuXJjw1t3q0Qj4g7C5+/eP4b3nDL1MjX6Gexu
SzZpqSb8Mz/Rd1/ntLd6ViWFNh+S3FaXtwo9QwkXZ7scKX0QVV6AuP/1ETY8Vfdj
MsIRiVBmMdQuXyihDCVruO6V+PrPmc61XukTbKt/9TS40mDqcN7v7bZLf26DpMDy
yHqqGSTWgpIa7PMWT+8EMFfpxZogc8lJkiurVHKUEQLwguE4efBgrldIaGoH7c8l
vHT3WIl3ovHlM6ufUF6WJRlYBp6YVIYtd1ZOdZobY5L3JBRgK0LG8nDOPQbkHx5U
wZjosRJNRj5goDQ2oQCAV8vSCVsbPYoLDK00/DRiHgI1d3pKWQe5NDAPUSn8MuTT
gWMXglnCj/uNrL6CXXrai7Ecw59i6eMzadqHivq5Tap4xE4d/ytjCb+EIR19fPx8
oe+trx5xk+qPabp5B94bQ5WjkInham53jSjDvg10t5m/u1fLygpa5+T/p4gyRtDs
hiTgx6j5AOJ1AqgEyuC8jeJqIJM9rGUYFZMgpl77l7jjyUmru/4lHL0osZJfqG+/
A3j+tuOf5RR/4tqUKDEvZdvepNez5ZBTxalqT6OJMP5HHrg7pBRkihXenvWpsOOr
hg6GM/eeYuLK/tUbSIS4tXpNv4q+r3upjnInAEssKRC6CMudwj5+TK+dR1XGD31Z
c3g2CZZ/4TB0IMdzzkFo4YW7wGeo6ohZr/F8egijxhPPU+b4IJhNihmUsPGR8Iw6
reFz6SpyuXpO7CFgf1tSwt9Z6SNJP8fykEv3XI4eKk3nXGmTjlpfV3+CVMZMBTdF
heR8oDvBYwLOHcSuQbvgU8tgoamWk9oQGRwplIWKFXATmgjLELmSeEltpEBTiQzl
8cDbIPyTL/4aomdkjacXCJIg5Ywev9YcDeBcyw9Dypl6p21phXAi8ZTRiCcEXDtd
pMOY0fXxraQSL64ksyzaudmzRw8oCwqG1jaMs0VC/XqLlibbcUAN71QyI9wyaGns
2oBl8gYqAJz37ujw26F9Lp8MLJKW6eeoDqn6uTpUmueS1822yRRpedf9UVyiNQbJ
Lgyd4ECAp8L0Omav1L2w8s6/oQ6GoSjbC9+o9VEMNueunphBaJv/tN+ouleyi09J
DV8O+Ap16dgnxQEDy7ve6qBXwmFXUVhzPCRo6++u0WEWeEEH/cq6LIe/4evSEwIQ
tD1+fIkHLwcLJID5n5kLedEADwnyE8p8fTipVXEytcAEIWFVPt85syMzRB/hp5vh
HAWxgDV5zA0JOPKjz4VjRX57Hpd3jNrZXcuRII15ul79pZC16m8Uz/nH3munEIjq
5cltM3XhaYCz1pIFa/L3nEJSr9/hyangC5O9pNtbL+10y7AUmUiBMfdcuGo6KPff
0s7scnaCCKr51MVFEh2Y1ZBlb/MyFgQvFosA0gWNNxf97qtvGGXbmSTpfUqlaB/2
qOoITMQR5h1K5E+jUiqxpLzdCehxmk5dWg7PJgs2eNlAu9wAwTBB5Dj0GYfYRm05
mkPS46Se5pfhjGeuqNicKhhrq4wkdX7XwCu2nEyIeKgT4WpRBDd+R/m5Ta7fWUi7
r8hZKeH6wj9jWTViowVQ7n/Oj+xDk0PM7u9KqVWpzoDHVeLuhB+bWHedk4bFtZbZ
A7Ic6ocJAFsUcKkSHza+wL5sWClIE+7INNSRJsUyNyJeUg1vNEDoXlOKb8VvxQ0T
g5mn+/2iAIEMldLynrgnK07pVHXifFnzPZYgVwD4i9khX81QbN8vKt3ki55vp4In
QFUhZw6xL/tHlFfz7ag/Ay5Asg9g/WFgben0hEH/Giblwzke6qnryogPykVnjSiR
DU49KPH/nMnmW9nENgkVkLroMrEcuSJB0ILXGZP1dJSvojznxpgf/p0694hzYtki
iM4nJcu9iILorj81PVH4ckqmM7buO2BfKXJ8pmSnsF5aEKvnxD4JEJU6/06oX0ZI
fTQ/ZOl50HyPQ1SrQjaDpjri3mxs/5+5Pu5joktBZWIwljj3uerEs93yH6u1azlw
YYHczvIxlJ5ipZkw72Ms/j1R2RP5tAseK2EHPgXc8X0JEfNY3cTUf4sB/yQPLj6e
OQeTBs0mEfVpGCA3nltw5dxiQBOYpmZa5hZ2mluGPIrQL+PhuaGe64h2EGXKktBc
wqMaJjFiCbvZ4QAs8/OO/Jt1cOEP5F3FfLbb6dTzEFggVpARz28LeYjniCXbkHON
9WBpYrlP7g6Zk2TNQv9mkxLvM5poJCXjrTvnYPVwLUQyfwoDUExTkOmo3Mlqstyp
hpwYM2XGnjLmDddbkrRhR5S/xPWCPkxqfqyqau7nwJ9RHtZzs4mcroGOTX7JkVyz
qZpCzwucubI0QNizHYDkd3qcXhmJga7raCZeSqQtzr9nYjPBUkYH6SPZZgypV8p9
PR39GO4iAtPpzuCWTk9auH3jpkHF2BL0QqMoU3jLBQTaN9R3hinwKIhhcbqMovU0
PTN/qgADcdMVmWnWKWCEfSIzwWuZPFh95fu/8pMYt1AT+wMcBxtJm4t6Bnoqe5d1
ZssTIOr1otqaE+SkRpNKkENaXOhtaitIF4b5yuKEJX4h7bBAI61cdm4XvCD5GQdW
ZyfIO6Sb43jPR0HUXxGMHxQkXPRVBLpag2seltIP/13I6popYc42mwzcvjW5M9Ae
K1zQvRsYL95689rRkQfdPBgSaaFrUsRWRhHtOZabfe6a5mgwF0Q+yw5HKG58hNYR
gbE2bETk3Rr/qDrHb+P1oraIlMIaQO3U941qqpefV7FnT1bLzt6hJ76mIXeNx7Jc
mNzJrxWAGmPKs79xEM/2N8t052lbNLvSFvxMT/CzDjJE6CpFit75oKwr9yCcwK7+
X+9rH2QZ/TDqZXS3qRJ6/vM1aqaSt9MQm4FNAAfTx52riI49oF9OUP2JfZDMVwNL
ecy2om380ZVDwN8Ke3Z5K4uA1yWD4gwamhEJxQy7q/L8RZ5W448lF3juA+3k37y7
ApuwbJbEsUbHA2kV0V7Uv9/65oMtrc6AZR/6GH6BBpAY3rUUrM4zEEJe/ObXQF3i
qMN/h0+8WL8iJ5aCpT3PpU6Jh/+En8jewh5cgpSghaNxRnuOANq4uDl5kv8z6qZf
4HXkxWQpjWsp9/HjWVm/LhYq1lc2v37gYzLyMUf3Kz1ogY12i2Op7U25cXZTCAUc
j29SQm+MSr/ajAMc+n+Gn15Eg7NfFYlvMtGEBgzHunnD56upj9sOVEk1+zuE8M9Z
vYhTuKk2jFmXmC/7zFsXFh09k4t4I8HLdlsGpjtg5097583LB9hzZHANNxaRdrUP
T3YgXbSXcisgh9xF9M1NV0cw4yIkLHshak8Htz2ZJnk0jiojGpVhcWoXQJVZOfJv
yy5YpqIS3S8bvR7T0BgSXKQ0Apyk5IT26hDfPm6Bz2m6xJx3l/d4oH5nJlhpJKSr
X0QvzztJFd1Ojkc6NSuemnYGu+5r5WEgPJf0tCc/JsFeDGu0iwqxrpHNvGHQXhHJ
mUhpxbl/EWbW/Vski+iX6+RLm5k4mQC8ZDJmplBsgu+qWI6L1Xu/V0VbxVk6xX1N
xsLHktrNkrJGQqbWynZGe9WTUwXXVUy4kfqPTgyivyLlAwEuVS+9xbqwMDHUAlKj
CXFyMljKyrZJ9ncYNY5qzGHJ7SJYRTMFv6JaHrMB+kiGuZiTCXK86CBQ0TzBiJFk
xbDtZgbmzsqNsC20W60Sz1WMNTovdUBpbiwyb6PNJKmx0FFvzBSM/HRrpvuHoJOr
umQEjsZHwhP0WY7RLGjOIiipUsU16z0UqEaZdmmnZ9hiEhpDU+N8cUqsOM2w7JMC
erHXuqgJpWRxuMwK9hvdZPsyXa677FkLdnn7rgueptkfwyyZLAAGXxbqbXg9plXI
/+tvqAHbE9SPgWbgL4FlAMAheJseAjYxDpMnF19r27t1qSpKa9Gb7WMMUiG19soq
81z5mRzQ+3WpghYQKuzpIfYyB+Ieq4rGlwLagqubCFOFc2USFP0fM9E9jvRDDkF/
jJNuLzjP91H4B+zPmYSVQ3mQJkPU3TdwBiIU3MdNiMRGMOJvyizVCggxIvcQcO/e
hHTZ2SNhZgmhPWDJUMU6XPkUzF/leSoghbtqaLJC9tzdDe08pDsnzTcU9hg0vNv8
n7B1Kum4Ri4Ee7oet4VM+fuwsFOpwLz/s6Pzayy7xHZ7ZSkbBG+aSZ3Tk2fDObE2
aWhbOV/07SUdMfMAiPsLf9iSnMVPFHz3KhhjP0GjUZ49b0av7BhxSVUJzG95t8hn
WNkVckAYBzaNveCFAko+fvcdr1eEM85aAm1PJeUDmZKIBZDalVS4fHjU5oDAyDlA
bEb4nWBuLhaG3kbEzdIW7DJ3ZsZWawTjNvpj+7+5Qma4OItdKz6NQTNGueLNIZG3
i/DpRrPpKXY1U5TOTHqmmHpeo7rproGlTCAgeTwKy094CgjDFb4O7TFoe4v8u0Kl
Jl1u4PeX6qugN3adrXM5SFxNdhM5l6RrbUWo7sHIkdMuQf+YWgZ5fDUGIzDL3NcG
ZVnEMud2zxUcFcNAsUq2gP7thJDfCYaM/6dvNSIYm5w7kRD283U7emjivlSYEZ2n
M1OUI6VYSAKdFi3yw67HH3pJHF2S6aqE8Pwxztp9Kq0HvO+FLhMknJPh+2gmvJmw
Hd8z4LIqZoSqMcv33JAR4iBza96MMURFSiMLa02jh6kPqqwEGGBRDULNcVVvnty9
FslhEOkad5JRP5bgGGjJuwha4S2rFtfAXyUlZi34RSuWmKH0gKSm2C29qy2LBkI0
v9tDdUJ2IuDDd9s+DrBw8IYxLhHQUahR1asp2h+HGqAhfCP1nmnHvc6bmhv5/g2z
x2RcyRlaO6GV4gR0641DHzMV3pscrdWXK5g2QrYQBEK9NpN3RaSnAbgDI7c3aToX
MVq2v6s5vRRUJ7XYad0kZb46gFh8xUimcvlm+viFF4UCf+rrgK51GWpdiDUrvk2F
NO9EoE31f7UGyLN7z/qjz8ZnxVO3zxFwUQE2JL4aGQaLn+fT8Eb+msxitQYylRz1
/hE20Ptrfhq5Kd2UtgeT1U986iF9ZPioaUxWkJjvQhlLdVD7XsAiIOOuoftmC5j4
srXR/nzAiQXoy0Q74jCEsAhXPkW1JUTDSFV3j6TI21oBeLgu88GzTOggGqAq9PcW
9r4mPUf/fie8wQF/623v1po9COrv/58btj7Su9MNnufROUkZTp5TUfWREQ8gNoFa
6/6cGdNdC8JDf1TJ+Z6GIhvBIih4/Y3aPMTGy8RhydUbroTnwxQQ94aOylQqG6jS
DdpN93InrTQXxP7fJnbSjwxpMsWPdF77FZUrqDtg171EqKfzyrZIwOLkmBcxZb3u
yGvQhm8/WfzR4OL5/csn0ENRouNhO+L/gFiJelo3H702odZN9Kxi+g9Lz8TWCNXF
eXKKs99+GkO3/qk0FjtoRHeNpnPWpf8kSW2820NpukGiz6atc0a9Pz8yeJ8/9nQQ
Jg4Eueltp51iOHxW0AhVzCmdmvt9RsIdFvPCnqU6Jpau4h0nPTWXC3mldWHz5Qot
mnzlIRMpEreMDWvoISnnSs9FHIdScdB3OOlBNMVfsPOXNzucq9dzNYScKCP1TnJV
j3A9tsPiY0Y5pA9UmjaUSNo5Alk7iSxGjVSE6yKKxfBT1Qk7GD6x8SuoJqnaH8/r
iSHxKyB27xfrrwN3SZUppvSpr8WAXvRTlxfJ4SSHPogX/u1841OWh9fvD2PUQKRt
jufLJntPDXtEuOXPCS9GUttJ19w7luYNJ+8k9kqv07Xjrmzgdp2326xrDsYB3bWW
pI/+XvfCfS31Z5SzS02rXb/S42FbC8v5ebfv2puSf7fEFzG3BCvtlTzCQzi6SQfV
KRWZe/1ZteY0XKY/mdLqjtv1lcaZ+ZLvWSInHqDWkddisfijeiyN59FjVJW4aOGQ
+qJcvjJNi/W0+ntAWbfA7rtwtfrG/io6euSSqboGWdT5Bhdj9ozxurfl9qo96suV
WOwD6doUtsoVTTsTUEphw6KGQdeWW6UkaeWWO5cjxMj6JzVhgIitJ8OnAcQSyLGO
WuwX0qx5ryUavSYBI8AQ/exmZQbC3F+r1GHDU8RyaWsn5hCvjbSf+HcpcDpaaPf5
YSgGN0YeHUl7D2MSVNKq1TPjnFmpJrH/hBht1MQKnTMyZgBtYDGmfxqhZctHBwai
ZuQmLwC0wzWpuMPzJa+3uq2Ug/V2i3zu7WTD59mew0GxfFb7uqeoOqE2qgYPXw7w
enzue11RtR2vnpTnupY2mxDLv+a6n0cb/x9T9F3atRF+AGp/TIgvCxtC/B8DYTv7
XsjQMLJqmiyI9hHoFRWiykKr4vlQC4At7KDBtWXrknTrFVrbEWaOa76/Ut0nB3ci
N6K7ThUt2xYWAJvxY1vGSHP2ZfI8oWtG+Jz5jFp8xZJy6/shn6OYcNFPF/JYNOnE
dyh7museS5i685/AhiJmSe3bpQpeMkVfRB+vNMVN/OoslBlmt0pDER4WSgCgnWUS
GHjA7qeNFTmV0mujJ9g2CJQBSlUqBziTjkotqg5nDktP/49o03+tsgl83y4jS3Ny
+tflF/tpCFB+2Kpm+4ax4I5DE+LQ6x3dHYTmKxb1qqNA+xnuVJFleZTVXhcFtcqn
AFkyWCNTv41Uq29uBAtim70zhV4F4rF7NOnO2hn5yFTltedXa1rAIVlqWXxx8h11
gAVFGAGY+cmHW75aZNSGMhAkN21nESn/Ta1vKD0aaXxCbGApBn6tcNXA0kHMKoJe
GLg4aqvJj+NfG8jkBcHJT1WytEXo2f7Bs6+lws7IpBGm+zFbzj8pPfMulgk9aD5d
UyEm0u3hON4uopHt3I4/mzUjBSr9RIhwhEimjHVwUR9/j51uxgBgcjXURNMx0RvL
rtq/l+am8xjcrQmlPZ9WyBbwzAATEIUuQsXpDPC8tYFxR7vRUPQ8v0bFtEiTb+Hb
vDW/4aZJaV6bxGr23qdo1rjPKNGC2d3PY+eQEQ7bqiTUf2S9oijrurz9xbKb1BDM
02A1yzZnKOMa98vpUebNz3lN6t8QpF2HDO3bvAQVzfJyEfHQFntaLkPfZa2ql1Lb
DubdjQbqP5iM+4Qa2ISfuJkPickt425ElM1TT6ql/93SHI1xOTq4OHY+D3E6n/gN
lpp8AM0ZrGmVVm7iF6kDE7Uu886Jnvcw1N0/hodETLb2MsgxPkJ83U1acVcHJHok
Xxlzuo7zJx7BhMV34zBOOPwCgLHecFBhqk3Iy/ZN33BPnHlLX0TjyYHVNiV1Hoay
t65A7rSKIoStVoalG7W5nNdTd0G8QOOtn6LOAHt8EUbjyJ8uBbx6V8paCIlLaVh8
SXm3H8Zzijny04HQchVYOZHQKywHphC4K02rVEfutd0WL0M8zofPeG631IupWaj6
C2YcMqLYwUW9PsJcFFRiCEkdjOmOwZW5LfMvbGCNvrQEj+UDPVpX95Qc+4zdRFR+
reJElqbkgHvcyjnoXxf4GVZNjt/3PXHEJTj43MS4aA9lejKGVGmdihl5wZVvdEhZ
zqeWU0NccOlccOgTwftTij8B3+C0DFKyunE3GSwDqNzug60RhJJt8EOBo9fcEPuw
0V6OkyB4wxw/QDgcFH+l0Jx5vCEbHrLjEkUSBy4VgIgMERkj4oJN8QWkEaZyvQRg
Zbnnc4XFV/edagiQa9oHJI8B+P1gwaFGrmtumZ5StETmew+K11CY9Mc+km92EWF2
EiPqGX7BlAmXDd6G0m/ci5PcakCbjzmKsxc2xdZZhqUhLB6TWdTKqfd+JTMLqjei
jcte5uCnLSOMjbAQk6lK+S+Tkq9ZgoBOO/6TAryORJG2Q6q43sfUlByNhmfmDm99
0O4wh9ca5hoja7/cVngLlr84QINPFybdxLxGrMFaq9RPmQjieeqNRtHk9unUgxwv
NXYKcSSbbbxsJXnohBE/hoYONtMpYWlNbEB5FUYhf6GURI/lskCkW98i1GB6q2Ro
erqm3PJ5PlXuA5efyKjp3tFePL8PyiurHAMGO0ZcuIMCSKwfBo+rRBxpcaWUZJ4F
iHwFhhd1RMH8bGVfzXbv/Ob7dwmHMUoJ/HUIy8iGzoTn5xJDfvwVJu+gXJDhX2Pc
9DRbqKclt1Booco4IOxMx/HXAyhxh+YfzM+KfmGZVgwzKZlrXA46KzTACEwJxhIb
33hOgy5R58Y2FEjYH57NBvMJ+A9ZQTdPQqhNCHS/ZeaXeJ02MC6ItKpki50+ti7I
TG1i50KwzIKsOcZWM395/UdfiuINKvyWGKU7KVSHTmP4BkiuTw6S5c5vLvnfYslH
GBK6JUVhbSvzw+q1CGN0bG+/P6qBsy9m0GSwAFWMqbojvzmz5MoXwetDiSdRePNG
TtQ5PzgzMoCxBo2HzcUUgDgqjyvGOWmMwoKzaAPSchH3HvzJPvn8msd1OUuA6YSB
nRt3LrzisRiJOB1vTBVOTufOnU8fb8UfIuBCzWnOp5m/yd9we+lvF35GLltPkOxg
hwreOqjrIff5U85eGBoYxnxy0xDuqc0wCliCcBkpIhg8Its5copKJBsjofEDp5d9
MAfWjdDm1E3vhvhkTb28F5BEp1gQyoDhzL7XX6dLSFoM4QX5G9+V7hdgLqDVSYoQ
MQ7F73yaGd8jBH83V+LPX5QyBR8nxejRAB/eacfQtEmvDSsoGIvGQ5R0cp6p8EHu
qFBCtBFiIZhhjJIOQULgN5XFBnT3K26gzFvnaSeKF2rU2/sZX0etyx45zIW3209L
vwWvYafBl7FmsDoXrppirnlDMsUq3+THBnPXu/kJ43fmEmn9bU0YJ2s7cA/M/wmo
xINozVpNXkcCK0FTfT9P5sj+YHemV5NIMDY0PyxiKpwFq9HDz8zfW/HQd86wDtU9
kOuQ0hHVPh7L+tqFkG7/ypR4jVdLX22etRctkdFO18Qd4g4QW550vM3ScqeqIrPD
soleioCnuwX41dc0cj8tnRjsBMyvCWIW9gideZnEGZA800Z4DosTbkyvgo0BsTKl
reQLFZIMlG24JExf1LSqIMT1CzBaWsgAUTFc+yg+ldc3V0SqcqqWMC152PgwcjE4
DYxqGAAWUSEzX0FkpCr9D3jLgbRT5zXjkvk75aDQYyZiEWVZrWgwtxaodD66vOaS
OquJ+UxUm+wp+4dGucwpOHCkOMxS7/9x4UrVv7CPitEJn8iH0Pgg1nztGVhINEBV
ibLtQT0dGNAdLIY9lmwYh8VPq7SWikWXphzRmSsHmwuiSI/Zw9RBhVquu66hAeKD
MV8g8FH7p6cM9r7jUNoUoUYkc+EQqWwtVG46JR5oV1Fq8uK9Okcc1oVnqx1lcYGv
KahZOTnNwIFJJ3cbVUFvkm3eN9d97ohDhngMOulzkgW7XSpJ2Z38hysJWO72THLf
sHlaXCfaYId7NlBdXOTYzvgE6N0n/UHT4zulZ+LRnELzDkow92EdzB41peiG4FJJ
5Yl+9grZersEl1CQ4TFqnMi7KQhe6GAcEckyNByEOfRhipsF6STsgtpzdB7iE+t7
352G/jXD3BTFWNHngQKBisn1S5rKqssVmOZENR2IL1vF7t6x7R4kH6/QpTPf03nn
RSJspu2DPtjSfIqx05wqSlZUyWObjn9VyHP/VnTFFsR7bhOAZl829MlZFniq6x8x
5hKj0p/KN5FhtYsocRSPVQrygyl2LTAGKR6SQyhi/txWRb4TT9c73/K7NRivxheo
mMnnlxYPFLGTp13fnFJkEW7ngJTgfgpeQPk4W227lzpkcxDaIYR495ZCWd1TiJAk
9b/PKe3L0DkrOXT0rv+iZWGiUXsdt5fAbDQFs/0mUGO5kgCgVE2BQi2EpOIF5SMq
QawPJrHPlOgC5nUG+xNM9PVlzE4bxuXMV9G+XNps1dR8Kjz2pV5XdnMX3STExE95
QfVzgipt4Pce5V+M8wnl7W39oTBTyB7FRyQy9YVnXj8aP4OYX6LsEb6dcXuvuZVv
wC+BLCN7MA+omeDQTteQeprZ6vuKMU6UarYNguS5oSVQ6b6+s3dnhRZZlLyX9lhJ
GiL7Ien8AwQ0xO2ghE+Bt4UsnIU3i2hbxAUeDWwhJ7uGGIH/KbKeKGna9ezfqv7x
JLcrng+VsGJhpNUeukx0Xbn/8uj3Tl5lZPE3YKeMQBk+Wv6Uca8BV4RLKECc+5hO
TdLqc1SEHC2XjErpUMc5vG/jXsMYb2cFv2lSXFZzb0FvhJdfaH7E4YshDgUk001Z
w7W+tgH+D8ZfbP2ikkZXvAq7JQxvKeiHamAmsKOLhiJGQEN+anPXUgjd+egaSqah
e+ACER0Llo3Tloq652nmEd1iw5wnGSDFoaWDdXGZL65Eic8SfzZsc2tm7tNfhAPr
XAySzPBmuYllT8jug9KU/YwFuDV6vxHCS6BiA9vdZyNGQIKm0w1fUAOxMXutkdfq
023oOxSGTuoEJC0DJlTUDydvM0fx8FhUVcecFy0ChHX0hyVSOVpzVCBGi9OkYk8d
+XF6Ymp/9UqU2ofNH8/ALu1+4iaMMX2QCNzRm0L5C8b7BkvY141mvpbKeXYzXvN+
BKbw0Tyo3IfZJLsRcHE+lLHfAPiEnSkUpbed7J0NdmOu01Q1rGwBXBxneDKZ/k55
P2mBPOliFTsm5Egua/jO1JdE3+Qt0zxIgHZ/SJ+QRtMP1CNKL/3I4nsYjszJiLnx
AVjzoGwOOic/L0qImuFHmIgG2Qv7SojDoqz61/OjtCD+KruIvQy8l51nyULZUV9n
NgqLFG6ULNrVecaEMKWP5ENTfFxgur2r4uWV8ugBIqH5zaXglR5rCqxwpAlHFO/2
wekMOqkZjk5QY3wGsI97v9NYRCv1oU9ZjFib8zV78aGqqANzaEAMgaN7k6q6ZZix
8eFDp3A0zyZcksOP0sWJOMBRs4JT6sCYMPvWg+9SO+G8Jd2gj7TLelzQwNA6Qkzz
qTuIvROjgl9HZnw+Tis6+gPhyKmVzLnSz0toCyLRrM6JyWEhNxXgS8vlKL0vhIxD
pDPs19NwXSBW3koudqbvQA5B/feKB4g34A5YtZtPuPnJRTbuHMtuTE9xeaSsRjYU
GXq8UHPfGNl/GhNfchM1tMmiH7JXuJfXa7QWBKr/HMKpW9imts6cESGlLGLo3ftw
kc7Aya3i3jCK0PY+8Bf8jjT+/f1R3xjzFc2ab8GlxOCHhQHfQln1x6JDwPocuzZk
9v1EcinBe0lRjoAmW7wNpb9Qq8WIBYHPtVgCQHQvk2QYHBIJgiYik4HpI7DJXJZs
mKEBIkkFb8HgMDrntu55CeMY1niEghJI7k8+ZdVHi7bO+bM7/CEcOJs4oEFOVrJT
FWs7cYfRAI5BqgS+HOpPV8bh5AaxNNwHPu5PKAw904ZDpaUZnm7XzNtCbLMAU8p/
ocs1qcjsYKesoYaXsmPIN46y1g3YsPW6gdExDWqZO6aD5XiGJjVfjV0ii7886jJ+
553mvNpcZattiHL9LnT8+n+MllUgQ6fPnh4KWpmavUXDg+B1HYMt6ohb9OnYoOH+
2G0y85n2J1gTjsFlNBscamVl86KzSed2lq8o21DZc/+mex3tvlWBcPtTaKSoJT1V
EgDwiV+OR1e4BVEfXmZbhdHLGQnK36+wCWJYyFc8sbDs20KpntHWI1PSvlUSNQp4
hTQq1MS4qxN2hlOtyAdM8qrYMpYljzDfv4UfjGhcambeYeFqQ1W4uoqth86yGKi4
Xfdt2POAwPqNbg8FSBFNmNxiSlkefTNXk43YQOaVbOf4fpTGpPs6R4ogveJlczCO
W58IPZmGQO9ul9tMuxEi8pd0Q+l79JZ6rlQnceDUb7A+0jmXbjclRwGH0/1NEg3t
WsJ7FqcGTeaE3rpw0bSTMBxiO9kCKPW8FFoCETihO8uY0kMcT5WgkBcWxXtj3I/P
2LLWgaoS1oJ0jlWUiXFkygrVrkudePKuO8GP86MzN1eXfUXs3aRn2qKS6wDyzJVI
dxMZZDAhs6qz6e+87CPeNkoXXDSqKYciNnv3mq96EOCJKJwMVCD+CyR3boRlpDah
lZVC0njmGuO+BgcH+Z5XsR8oTMnTOzOM07IuIGcBQK3Y4yhnpCl3OEjm7I2RJDaV
6JxG/V0ZpUVBmaHVnzRJNTaihSpaRVF+53BYKFPScfo3FC4nM1RH/M6mthqtcC1J
puibuyuh+4zOAyVH3NiDb+RMJ+bjKdsP6gSx1WUJpZvvW5NxbvGRewAedOgSBulI
dmgdV6pQpXurqQP3kZQvXp2hSbJoYeZYKUMFp/6l2Rxe1dPmxAwkoDRxL2w3cW46
dEZdkMbDrdWfN95bCBUF9BIsXnqDwR4ygm2EeUlLq+m1P+AK6qBCqpCjE0D28GO9
Htxcxl4i741Ns8XGoEh9UKWViRlfqnLNbSHJhMT2+BBC5zexwX6vURG1kIk+Z9x3
uUnyiD6CqtcWx0x+UyBxr4H7SFgBMe3JzwGJ8gfNNgJP7DSv7K0iUuFXUosCEaLk
rah/MgjLTWc86+2cO9FQLtZIhiigUgUWAV/d9eEqDl3bCG7sD15UcVsImOQkuSmz
KBjxjlQLQMZH9VMOfnJdKzq2/FDr2i5zdiVTSfBtfbxCHTgKEHPS2IrVy6MW8M0d
gS0K2VfuNjLhgoqsDHi4b2qeF1bGX2WViaQPepXuG2RWjba4XXamABU7xJfI3w2m
2X6vO2Ky6t5EG6l5PXneFuoctI0o6ZOOq7MAgto2JjZUWkce4atiRxLFtvm89ZMq
C9yMYcy1HvcIH+6ac7hHBhXNE5Z0B6dgctVo8vF4tTfkf6yTgBfXm2QcC0jl5BQu
K39klgxv3oOdMVfVM5yJ5SjKaQmpIzRrJ/fJAZhVDEoQrEtb4O1keJ0mHLWFt57A
iG6Zo6g8XPqi2UAAAATNL4ugA//ivgfDlW0q9haAtk0Isy4Hd9oT36BHlbWMcxZT
4LMY6ueby0aME5beFxaz6YI+zNDpukDIhwoxO2YlcXONVb+De/SaYzKLL27vzMeG
ApxVVMCldbjzmOZ/yLQyqHzxDcWVzlJqDLLL2FNAFIPzJZmcaQ1jDD2qS05a995S
umboj7ezzmhkt0ADwSK7/2z0jjO00kiQMv7BdVKsni8SElBwCXoCybLkbYjW4UOJ
JWSk7WX1cxiDwyOPcRuB2w1IWaBkbimKCq7J/DzZfdczSapZ1vZTu43/xsPXlAnY
7QCZcbIe4Tpvs07pX8Yaq2PcZlXngC45uLJNVKT1gWk56cyA96a+v6jc3a16qEhA
jGuGP7pHzIpfN195Twc3QfU8KlYLDtTA1N2slRXW8ShPZx+nrBOdDPCMdKD7TqGp
FVIJFNH4a16yEV3KtdCTeZKjZCB+mg2Se6D3RWj/a3j8rGHCnIESuf/SIiH1sBMW
hkBK5Qq75i+lGNBG7zBPLPxsuG9ltBtjxUTx5cuJYV/VQKmOFnPKXIQ6pi7x/9Ze
9lM+XK8mel3H9CflHDWgpHuLN21ZHbZhx+B5f7LKwt+tvvk+6WDttQikZaejuhCM
tS4L6jUTfrD8x0aUfHWASAhtbuC8IV8cf/FnZka+KMTpyLuvaBiQU/EvSput5kWe
RP7v/CvgQMw3tAx1V+pXZxJDIy+x581+kKPU/CTA896HUzwL8CjUG6a2olhNcFgw
SXqMQ83DHJxlHHjH+oI6Ol9xpVn8ZU5KfS694k1jN7Bt+2r6tsCmuyYAQHu4K/a3
1o2hcqZ5AbqMiaqgJtSEyOxlddKWIJjVVL8adNZIJU8PyAw9/6jcZAAaiLEhZHKx
I8fIaCLXJTDn6Ci9PUlWy+Dn3LBdbdguCBgH7FCLlgvYsXv+U2GF6IhlXgPQditN
w4UY4/kVgXfTy5YiQGidAGEzDy6ZtbDJOuu0xpQ1hNb4qtNJq9wA8HLWiLsPgNNb
uYleig/fZ0MaGYzw+XPf3igydIauos+rqIlmgvmz9JuzAR1J7Yu7mxHzunZcBs0b
/cKxNBvGtxMXEvw1cVYciBZnEOHpG6VdQOjBHRKdY+m3YH/Tkra49ucxg2EbsBTr
l/uyIwwTTeZjGZTQMxPZcJ+Ly/AZpEJMAQDzikRnY+0BKocCODWP7xKh+lu3l4Iz
aALWTY5QQRhYQq8hQlPbJS5xtOsFVljhiQ2VURlWXKamald/5XDLGKn6TqJk1WdQ
5Bhu22v+qw2hxyJaN/r1mUF74wHJdTr1n/uDaaNtc/5bC6iYkhYgMmqkmyhhZK/N
MkcKTt3+BrJrW/dU5oe9ie0MvvzO/VfKqZIJElI4vO6fJZOkuDETvsa248pHFpXn
MNAjyhtfGqSP5JkobmZyTX7o7Y6qEX3FkgNYaxSoEyz22BcZnmid9GIXDqRPWPq4
vfnqZxJlARUP9UsjqZBdYv2Vy1oKRaN0otI6YDT/SBGsP7ZWWqQzwLwc0D+BlIh6
xCiPKSKzNOXTa/MQHy1t8QF7/D0PXafQcVzhPn9iOSOEQC9ZdQ/03Jzy+Wh83yKY
iXxFTYUpUacZvOW9um8mXtbHS3f+qKg95NjMDAFk+bOyyvvOfxljVIBJKCuIKXrn
Q2zOds/2TZmXLL7ZTQYGVi50y3BxA080DRJ3mJo5wIR3kl11kmFaWH86fZlQB/g3
jC7UEGj+mUE4i4655pbXs2G8qKXiiqBWlmziVJopORmEcjBshjHJPxaybexJ8dOE
eOnqzEyShYhM7Rt2uGRV6SfTxMMIW3TxEqHbe98tfA+G0ug9nmVRThPzKuXw6KUf
6Mg0cp/Qer3HnTWpmdiWtQq046PRg4CWLaCMNDl8dW89dqvxrScv1R+SvMGXivQ3
ZRvdgh0mJi/4R//2x1+c4nsSdrx3FBo0apf+LPbqcPkCKvTdyDfxx/Mu1L72omJt
qlp9g2XQTKS49RMXVhA+OOSmLQT+XP6G13xxlVxlVubfLuYo5Nu9ugrskPydVUAu
Ox5Sb2hv2LQsmA/YAhXnj9BEFHm7YUtg96sS2VYAf+LGpO2C7JwxOg1fZybLfbXH
NKJ9jTfoYRW9+aqwwRdicOeGeP7Gbc5eyjOLAZ7e3YIiI7qf6YiOHrGsVxEjDRAM
YbkmqgcDH7MTaD5bqgduesf0pIxw83TEWwtBX2rnvzamfHDGvOLvJ5CmzqSQ0DkI
5cArJsyjcmUfbihU2yjLHhEM3Q9zZ+w/63Ov4BfQqeP7xCtxBOmxOXs5mWAQlVWW
eYZP9M5/BW1L+eWFF4JuPa23vSik9gk3xpOVzlQGBLUjCoZEOOdG7uAgMOIsM7wD
s6/fFwL5TYV2tzUH5j7IKIAy9QgoC0gS87N/lG3qVs+A9nse4wHfvZLaQNpq77Oe
3vhVlckpZwNN37Ac31vSrNAlVo8RwDyvbZOwqevt+qxAn+Ej9LJH5U5fY2tszz4v
9UDL+L//+QXFA8222TPfjJ4YyOFAjzLQo/e8a16vq+PR6MIL+LbNmXVEns7D5DJO
VziJanFm3wm3qMuHJI7Yan3aYY0nA4jf/5ObKhntH7g6S51s3ccjim5CJunsbxkg
77BxUhiKogjHO146qilEqXw0mI2JLpo1uNaCa/o9ayeR2RuefoWkAiWrVAz284XW
kBtcSWkRCtd1tRqI+38XHMsJp+hgyLIDGnolRkZ2kVQ6uHnYO5Euuj9SO8WSMx7n
iw2+7D7JGAcbEZjmIyueLyECCU91qRFtvaJNec+xCawida1DEnGyM4WxXSbxwutA
yp3OI6fGf7bElLNNIYcXQddUu/V1odD3z4S6SZQBTN+0rZsiRp/biMZMo/coxu9j
tZsDVMyWuc6Cdm4PbrO0YImtQY384NDpA8F3r9eZwCNwhoMXQD4dw73Cn8GMzORM
M42dNLSlWIfe/xKcHefo/hYATDjCjUHFDi03/C9tOLfctU+ifA7Cy6SbRmbCVbC5
CNxCdSV0GMkUEkt2ChvdNjE8VUszzmge63UFwW+uhtNLfe+P+y4n78YJdGFGmEVd
UApuy2gOp+RX5McgR7AMJ5SlGvez1iwhJmqZ7Xu+A5xZzi0e36UMb5bdEscJptw1
Koe2twpzQysw45WGtoYVbbwv5WV2DaRC9vWC1buoQvARvRcwBrhFblNHUOU+iVq3
nxGuRrLlN/35R9VF0Q+OwWrjEKojlLf6AUQ+LMrZZJ9m/OOhCs+FUn92GT12NkIn
2kj1uozNdLwaGXYLV1YVeWBqDNu2lVl63avuFNl6EsBNZcqewM+pB67Gs3tzXZsv
iqzaL83f8kddHO61vynQ0JXXPXs0xdlhSBgTYwMeYJQ5Cpogu3gfqPQvVvhyMN+C
dSyNDCNyg8mtNMTgDogJ03S2dnvsGZ+3wv19lFDcsD4Uk9lbRudpxmnlPAmQUT7S
Wv5EhoZygHy98vLYEdX2VpcqcIlYu4FoR40PibocDLTiC5eQb445Alf9nm+3ZNyM
sAwobrYvMYhxkuSG5hKofj0yVIolJTdgeCg4PKRwTFXJKIeJbLvrmejyAjoa2Kdv
d88NC+P/cATMSI61TUKdESKBEWdzZC0IxnyIPD+BIm633RBuLhdwOiEjLMTVDhL9
IjPpxcEJ2sSqVnWsrkgIX6mNqnY1yzT1TZFNSUD8DYt0RFTazG2hceNwH5I1i3EU
Aq7WrarYuhRUX/tqwhwIa0/BdeOEsUInEVS8gs3kpk1nspV0gWlSVMHkRHU0k3Tm
/RspVd4zkUz/baZKJoOpAEoqwLTdm6GiH4d8jswqvuvd+3FRH5KbH/pPxEJ5ROiM
2QDu8iI/e5oclapQje8+/VqZAAaJtROkkBO9zqrLfSv1oE+tUTLlVubgokNjLO6g
KsGOtcbS5DTVNyDWalakvFzqP3zg2Qo9BMbfdyiaxW7/tUj7SqxnJAUI4R1CAVGa
LNRxQo7GkHD1L+GqNk9PrfgWNz7mI1EzFGkWdSZ/v6wiA/oIAOM+aPNQfofi3/V7
8P6A9L8onjGS/PvVEJA5pQl6PdgU0xRSKfeKN//bp5LmL3Y+838L4+bvJv0ky6Ma
jodR1IVlEKWTvya59ZfVQZSIipW5lrcw3CL3NQicfftAB8/q5lgW7aZnWEoy13NN
h0qajP7aBwu92otapEUJV10AcGoXZB/id5KQKxWiLKUYWpYU+k9O2/4y7+eBZ6Ca
WYN9pZfITGb4l3S4r9HxXomg94ohLqA7EoGgNYr5jIno2Uvv76HYT9t55+rMjfJg
nCaz55yOzJfuYrRIk04rsJKi4Q+/XlGyHxMwFse39Xgwf25REtwWGhU/rILGu6D8
IuV14nKu7lQl/dzA0RL78xprJhrp5Onof2cGRU1EyUwuuwD3agWkAbe2Thei9Z1G
25okKpl7a538lAhSQVHEBImx+mOWSGk97n5NptugE+0ASwMF7eqZM58DzXQO+sl/
IZwQBqc8q45IxxDWC8nUjKDZeKFlLtrzv2pSZccDcIkFICNlKv+PA7L8RCTwp7zB
+P/qsD+Ek03VBUOaX7sKV9X9lTw6WXLJ57O+3XvL73zj7ypzqHYYIm1QmY+KZ8FR
N4bp+aXkSF+s2UYz5dttd4NE0mTYoVqMNKVsz2H70DioB4wl8TgdmwZR2zeAZLcy
7+EziFUzGCmBBPyoImDx2Q2sV+hc5gmAdNusMqKGQbJ0hYk5lVLyvo9EbdYrOwc+
NBK4KVH5W0PCKXQX43ISF0mTTjrpdWHCGxNluxy8VXYqK3qoEp5uzjamTa+G+zg0
fbPrwp/yuisNxUnH1mTQ60pA3ZLZIeRZt4kz3Pa+6WI7lIhcqFkiwWvoYPJSNacY
stxwO8C978ime2X4q2xWsCFZAQiIuAKgUBx8hUc3T+wiwwJWWaZClMm78/mBCOIO
fSzfEDjAhXxpydck9bThzS9jnNanxVbJw5XCt+v1sBSfIcLrOj8vCiO3YEW06E9s
rQtan3p3T6JDHeV2zevE9CQkRXvazG7EPP7+KygKb9j+OH+7TmZ7rj1ngvyguQGY
FgCyHyr7KgrdNaj8R+3cgi+GhyFqcVvncQJLL0LTK7ScP8ZW2FC4aLTgFfmV3zYt
jQindOtZyegWN4peSzfKj2fc/08R2JSMqDTR5BZtNZGsx5fkl60rG6pgv57wBW5n
ozwQ/1ZvWtHs6RDItIVBkrFrxxRWa5wr3LLM7WtdiNjggA/YrCZgYRGt4E4na1gu
zqij20V/x7IXfhPULqaRYg2I2W2RRnTdS4SGml3Huu/Wa+sjP1/EJB5ywXpvRd1q
szV7gJxk6n+LFkWcH8rRgWFwV3tdW7PalfNGoTenBU2VnxuE+93IR3oqvwWkHlHL
QwMKdmPLZEm19YT2crBxRJQwPAcpyMqOcd6+d2VQSzdgPUfZn2IW/FsCk2jGrWf7
jXTSDRbkuKCeX2eNX4p81MPMV3H/FXxkzWuGdV5EZJ4ymQASnbzLebZveD+oj0yO
klt/9UsL1ED6Q0bA+YS2hJQu5C/aqGz1sfd1bdEjYsiNNGnYPBWxn3Unbobb+eP4
GsUKNgaW0dRpoq7vyrCTIL5zIFgSt0YXfzo10iy6dthAvxYl5wW029FujEeMPVRL
ZX1p/LO6ZWueYS1dDnioPieE5vApQj9/oRPhtYveIDmM9yb5skr/Jy/ZTPJBSBDu
NyMWRuNawiMuaLi0h4vDQfqDPHSJfduyrPstkeRBHw7+ymNHtR4hMbIze3UET7a2
ANiapX3mI6+yyWsFwWDCdfvFhJYN7M/ecQBmF1ihVIWqGJ6YSsPkeugdvNt8OLka
lgWFLz+LrpjLCkqSudsbSDkphcUaZoIRcPmNkmUgiTF4ijtTu9jKj9niKiscB3M/
PaMQ8R1X9X1H89x0Qq+J4BLp4qmkD5Tz3x3ddkhmVS1Dr9Fmbw20SjgcvEq6b0kW
zdMSm+NVQbepNfv2byyShlNJu7qVUsJS7n06Y0um+B4aICdTNXDea9FXC6Bt2Qiz
NDd38vKPjBBdyzUG2JzX4fbSyF72srwPJBf2FiGgFsAH9sWHz6B6YkevUA3BMrnN
e7LQfAZB4enhxL5riPjamDHE3tdiMneYDclmjO41TV/0eY/pBZj9e29L07OrfTOR
NB2SxkVBucpHoNfUT+/mIsDCdzMHMmtxZNOX5RGBItBYDTLBWEfm6FQVbl1C1UGh
GfkVGTCUrXKReye0uMey4GRrNFrC8eVoeeEXW8zmDiRRfv8chuZ7xuJP5ukgZiPl
2gE7FxyC7JI/zktx+GAci4hZJ3XEnQ2E/AEWIOe4f4DOh+EAaMUJOUKwXgZ/Hobc
G1mVj5q+HGUdXNn8QlxgtMa+zZGfhsxCPxhVvVoWMCfmW6Rr7sD0isuTPV9Byki+
SQc47roNeU2uWS8i7VbwnxD0VdDzZtRbpF4Qumizr+rOvTRCJmMa7FKTXSLGjoIU
GibuPpnqNCOJwuiZX4A4xbToHyX5sIW28YzF9GKnZNcA+X95wZbRg9TuWZmD7wpy
2kNEWquxA9fBObUqFHATt8j4Tfl/zH6WGZ2rM8cv/IV94AiTTSQh/gFW/HAd13hs
fPGeWUvk2SvToXDZeLElraH7z2S90Rq1WElsxHOjzYkVG3vulMES03LznanYU8M9
p3cOttE0WAyAUEleqY4+HYWGlGEy6for+/N2sYJseVOGPndfc3dyW7GmSjVUfodq
L6MqidvmZOLn8WNX3u64vVFfCI/Uiz9W2QmR74azKdQv+ddEqH1w3xQxjV7xf8Uj
doDvSNnof/eeD+BCsR2d6DhLPyEVm3eqnPFLkpnsnqgMQfrx8IQlDfN3xWfoeNRJ
ggvwbDvTLSUN3WQBHz9GugtK9Qw2v+tHqIJtoM8d6TCaXQ0yFPhHiFZ71kUQqj1a
A0r1x2jUC9G0VF+sM2fVk3g2MmjkHkFHiEwWjcqyMnCdX8a2pZBHcliFb09Z+SzP
WOQNWDmd4gBMxhjIwU5Hk4Ortsc7VV+NUDZNTw1JHs8fXs++ahW9X/8OSwAs964H
5JG+A5VYvzvF4YYwSgLP6NcA1B4txPy62+Atn5p53sKKAADk9v6kKjVqC7gG7DnU
76Rkb3jx5OBsTeStIbn62f6MdM6DH2FFdkka/XQ6axZSPALFTlu2cN67UOhw0FU1
EZPLp2L7hqfFomdN9/7eh1tQmA91M2qLsK3q0qquQBAa9Uu0+r6caybukfbkxQDn
enXh2ii6Ug+hEatNsQKC7mxZlPj6jliBuoVCS+X3RTzV5BgQ0ddOwfK+l1ufVCWU
yaS0FIOfAt4UFuMP4RuRdgjGCum73E/qpFkMelObrcrAxCYRQMqR5eWzlhA/XDmD
lQtWXl1EWD9HK5iDrpU56VAGBy5mp4mYbECmCbUAFdcQFEw3OkMXIciv4dmg0FAo
brUvPjQMkEMWljSv5b/4RgCjNAzi9sbax5G6aKi24xU3zM2J5ERjMfE+tsd2HOl8
C5sWc6Ldi6QyOw91s92qnaze3/HaSj3HrDdTZ8nEJUgJZ/xdq3erZFNVH16gpPCw
YsHz28YYNtF7msIem3Zcdqj8cs99SEfoV+gu97KlA/Cc1M/utw6ReaDkat95oBg5
uPLXc+zTDx6nCpPup23Zrgy6WfcD9P+Fei4yaUVOJLm2fzuM25evXEaY3mX3+rGt
Ivk0iJ/hknOQ6z0phdBRZnPBipe/ZUezy6XSxZ8/pCa/7ScAlJvHBE6jTkivK8q9
kYfRITmMJky9pWbAMFKY+J8w+j9pTlRWn55Hcgnq2RnO5bySxU1TrGPHF/+P2eX9
2HTlWVJ9AYxnqF7xW3gCRdfLhjaY+QVlmfVWS/D4qH7UdmN3DJo/fbf3ISpa1YnK
P7l42jQRERQWnEpZSKxnxgeNAgteMuGJqB5D+MD7ZVFWX6y2wOiJWyotTP+JI7rK
6PUh39X4Vf/o/WfugHxhsq/d1VNgfRgimAIscelN7rQEjLK4znnii5vZwS53UTFc
4Mn61f2PDhxeNo8zKwTIiju/qehtj9vq8grsXQuxWAfQD3+6nHFBopPQ3Hi1N/kM
zgL2rc0pxMcYgGJpHL909SiGSEZaVIuvGxTVvXKdQLYOYUXn06BhN0BhZcVLs4p/
DyD98M6jeRwkH+47URdDnvjHpQylia93F92U56tQF0Iwy6UKSkfNqSkKH+f3wbZ+
bXb0FP/bP5v7ez6+8Rc1+KzfFFVZwcqEl2t95Zp7P8oeIkCvcRnpR3JxfEGWI4kQ
4yHgit87mfvThwA+V+HDQBTx/4AueU++WwEJtVHyfDSS0tftKfA6cdIHYX7FaSVU
HLOBkGOO3/u00flAg0UCvUH7YzSVN29PXZFLaRPoHVc1VLWvz1OOHGRDImfcGrSM
UVYtnVrMaI1ycNEWyPiWorSCFi3/xnHoADIqlm2n8GZ4+W+9jEx++QiSzBTLA8JA
nSvcyK/YEOjm4poe4ln5pMypxtz2ORtKBPurf3wCAxktTKF7/qEExS51iBNrrYCH
p/REiq5nYueh2xQnPPBLhiTcMpe+mAZtdmXu+W/C/A7jmPIo+qo8/ZwyD5lC5Dzb
5daywcfxVJp5iQEzt3OkJbtURQgHC3pbbmtb+GF85K81Ge9s8f282FSYhVLC1KjU
0i0ftjjLejwgsICtcV4he8vYl5RD+JqHJyjy8n6hy4qin5tt3FwGgY84p4kCmzBA
2/dzyK0Jy2786ir4kqriYpn9vzBK/AYm4McqJ6WhIvFfir30PSBj/dau5nkNe5Cf
vIcUbc65LFseoGzdAOPNmFrE8GwlIi7o4sGiW7HInTWl9hp2pGqg3yGxvKoHcW01
DNuHt7beIguWcwuRsoH2HR1KeIFQdWbGUmNFsn4VaMBRxx9+WlxP6tIkv1qGTWEA
SnIumpV50K5GRG1bmVvfyHxmXqQFmxzXUZeqCpcAoOK4mI5gYos+Obd+eaGWbEQ1
FuDtoAI1Y77ijgyW47eDF+rzQEo4ewO/atOGBeQG91shosdj4tP7VBaXnlS5/jqf
pu4hn7Mkcb0iFHijx16CJo9fFllbDoOQ33KiyASxry6Hb6b3kmDKLUEpfC/mMWYw
0hjZ/eykHnbbZ3Wjs95dkwhXAztLdxUxJ9FtVyZlf7SYeXMaYLW3FMoPU9ARm6wu
oliqXZpyYJ+ZSTfRiY5eh3/hN/MYiJWZdbk/eck+n+tFH9k/doItpztZVqq0OSf5
bp6Ko5I/gb5+OlFKSMe5sy6+cK4j6z2Fx4kDtK7lGD305xvow1rLBTMicJn9L6Ys
cuZ5DNw44vHWN1W+L7zFz06CN9ZjwyMPc+bY+buGiaD6eMK8XMJkB+8YVHmLJVxP
5YYuYuzkPnqh/ZfEcIGZkoCdS1na6rF6U7oEJgEL6RNk1tKcnnMczzgBsdFRK3th
wVl3lUHKQXzIrrf7mO40ZOeZ4PjBi0NsdckoRdQ2i8ujq8NuaXRjCFfOzvbD1S7V
dmSfCSg92N7F/SvMJJxVNvx3z6TN7MWwCGDxU0Jfsoe6ICJIOkZKDkDXw3S3/tkq
q209cxk16cXA20nV57gW92MistZdY7aj96pxgObyC8e0M2ocNTOiiJlzJYgCBLJB
7SScl4VWsBp5Jw4vDdyXkbfFyfbAMwyQkJzpz6/wGnDQo2E6il+bzSD9w6DMkT0N
q5Y3TrEJ+tCR21ylVd9ZovVLyWzPM6Myh3fAHHm7ELRZ3Q5JRuZZQnCD9TlLLgD4
fZGMd8VzfNU2qYTiXopFfV3PuEQSWwPpSDwEsaU4euqSw9sz8uEQtjgfLO8IOXsy
W8XFCAU7atYzWbyeZR/65SPpeXlvtSyBHNb+I0l4roCogPXJH0bBMIb1r912DegL
V4VmHVYMjFkaOqHk+ODKkJviOIeYYkxOy9Ph8g+zaOfeZBoLbjY2vcgKafayiQ/u
PH+2iKDv/hSDza34srHbHL5HuDZFGHyniJyKzx7Bm8qDq5kEJuEoAUv7bHSaNEsd
8s7lr760HDzHf9FIlE/lM9vi1USo9qsoKS5UvNcpT2Pn+9pHzZxSi07Y9YP9fkAZ
RiA2Y8YSx1Yu97nsufeIclo3gpSEWDnC0MaxkxmODhffBt7GQ9185bFj+ZIK65rb
IozTh7Zs+Nk/vyabSn98Gst+/ifYeTfsFgdrwTFuXVVITMbDPYjsCjnC1ezz/oCl
rKIwYa9LQahgQDetRBS0HhWib5nQ29zzrM3BYRVBN0kScerQKXbQCv4NyKP4Acml
naLugJORkwJjcUrdxx4sBxNSeAVYL+RWnvopZUXJvLejmf8pWuLHV+E/HN8uk4N4
qWI5EabzpHeshHgl0Y9JghFzu/IAaHBHB2R5ovvh10J/gtifMdzlVj7mQM/vp+bR
ahje28Bu4hX/lKi12dfH7pU9HcKssoOiigvXd0fHnhoksijjSlipAdxnfHN1WUqg
vRNW2Yyi+wuvPpX7OS2mO4T7G9yWOoJB/2G1ehQNeAjvv62cGrXtp+LQHM1R9stl
ctb3PJSv8Kc6/Unjae6mPThA83WfcYy+W1sPrhnJUGThPjNYZNM1UkPacL6cHwNQ
R4QYi+LelmewtNU58fTX9fpuZQNgii6tTydC6XAMFCOQfDlEA/csXRprn2/HJbUb
CMN1tNgEjxEw5JpDxdIcYv7fl6Wwf+RLaO6msNRCCLZ9uzK3QwD9sxYDoW2fMt1F
mKEzQWW+YqN0tnwy92gQxVqjStyeIy9+PT1adQDmwRBqHl4cN6hP+VVg68b2PDzi
wuobNl6vbx4VbTuS4JFYSw2PIKx8kDzMYi9VILhQopkLHZII32ey4Aaqg+wCKxqk
0Phz7pCXSv6k7OTmnV0Tpx8PkQaDfWuxJdEHPiuQHh9ggB+GJs2AGoykbH45Ouww
1feywLEY4KsAIQijyg/PE9QtZxYNwQxQ44sjHf8FFevnT29+wiuq7aHHWQ0gxt6F
4wXnEGBVWRWxX4ErzBXnBPQuusil4QqhwKdc2kPn830pRBrlFbRZV1w0mKsVcWl4
c2oBLbK8OMlOVzBouF7lWQ1/yagkC/vJxc7gFHhCgxVAkjekEBqON/2AFXsJkBpN
hGgjBqF4yWyWzPdubt/GjNUqXrCujRQwffoHOACwOZVqo/9RjhBI9Lb2DcTpAT0y
NP3Aqooz0zgZ4BaakEtfd8Kn1nXH078mSiGQ5v1yjM4RmtwhhPKMFlY4KAEooJ6o
ECIf4Tu7jXwa2z+Gg/67lbfkD+RET9vegnyRV8aifvzf9h5SgLGxc6/3+jOcZPDE
Rm3f3xPkAh9A5D6khANIhWYhfmiWLrPO/qF/CDJmblyavgSH22jWAxGywcEqxJk3
QBUXTZo9UZR3uOTTcARfSI0vFm9MNuYSmeqSxNo4Yrbaxrw2QVyZrnKxAcd3g0zL
yc1BUzsCFESyrENiLLb605qdbMHWRLTd6st1XqOPHIhKUOkf6x5eShcpZKi4fUXA
qlX1sbjb7Y2OTshr1SkpUPHlIL6zuUy6fk5okgtSrjC1jXIFXRhEChDv2g8N2Ab7
qJvBzGRcNWxX9SJ4+lX5FnSsgmNpO7LJrTXFgu1m/2R9mq7zm6XTTW1Vn/VE3jYm
linavGPIGr6nHdjwpp8aRTX/5ODet1roll2sg2nM4+S8p4S3kUWuEsY1uO2B33Z2
8wBZ3bRQsRBlAJ5hO+3NHaF7ldI3A/j2lkDpNJXtwjTpd8Ls8RtzVZz6ec3WqDkg
3dIM9Ev4qOTZsUcpfpiekAhpSbhsUi8v084bFXCU5/E9OIY02r3N8Yzg+Cq0jHZl
HSZrxIUuhVxjo1BlTp95WuH3G+eqSyTOiGSE3SyLj8pvPNPz3ovNRGc0TbLU4ni/
iTbkM7uG5EiBNPANOW4eGA9v8x3OEuB0jtxPqUS6xHrlzh2d1VkbXQ+Vw1CiNY2Y
yv0FBbwGOYGIlIWxN0RAwyR1IZPz1QRtYTjhsLijdVZawUjApxIA5Be+GtreTa4c
wC+QPsx8m22WPRracVkk4Pu5IJjA9nw5fdkEb1wJNErNMkM+le12XdY/f6lgyMwG
8H8yS4gJec4R1LEL+1tNptKlzX1arYdVcny2NDKH+be0oQkOf2Wigc2p5AOocg3D
zBqC/2KXKLXqleKIUlnwlQancsYpgSktbMwRNW67yChKZFV5byvcOhKIfcpeniQN
8TM7+NPIYieF1BdKVTFg7XVCR98Py2luscbYDubpkT+bfpDDiGo0508Yidmyozcx
fAMhRZMH+qv7x5ZT14FCjIIMtMTkjHUAqmd38qAz3h/zy22LfzMGuBMxrmkFBK/F
WbY0eM2N9Np6Le9XH8mbHSRO1Ot1Ay2KR262hCU+gRwN30OG1B3ZSAUZ9/CyHHWQ
ahh0EQXE0y3KhhoQ97hvr+z+PEE20JP0pVbLGCBFCuh6/6TyIk6546QR/coTvV2m
iiYOpu+cDsTFsBkqFBi8k6pXHUx+3qm7imSOaw8nWbqNNcZF4vl+aQLXtjkM8dMa
i5pa5+L1cob/0oMcQ8m7dMHKqbL9+YHp2i5UHZFkpKMy+DLWQsit9rLdm7AQ1Bvu
8y4AW6J7aXwXYVNxApw+fw/P+Al67KnO9yWdyt8f7D7kx1ZFaYLCBBI2joIMbsv0
OQUIzLTov1laV1GgblRbrz0STk8qpaMQF7SSuKI99XRrsPBLVIx8ciQBowmb7bw4
Zgxg67HnkO1AqBFRLWfc2c1k1z13qXvOuviSUT1pavKLG9flbOXsr+BPbDVbdwIw
bBb7SAt6dkR4N71l0S47rREx4ckUXo0NQ4SP2hyCq1ShDH4k5tZGNR/lG5dmcd3j
UKhIaUFrCpCSAzsdAfhhJzQIRBbkLDEtofwllG3fPfY5hL1qDUAUvP5cKFbzKMjc
0Qzw0jXhAkaRYFR+HeuYUpFrUCJReCMWIjnS/d0nlV+Co8hBbNaRTEE4Zs5iWbIo
jHrG+tpTQCggv8FyNjJUFkyHaZSlnvMCWY+65KmxOuXAkWSYI9pxAR0uLE/qWk3T
gH4oO8NrOMSvbh11T/oew0pNlrtCNGNXNGYmNkDc3zNnMx79klmidwRD0vBs2pMo
WHW5sTHSTQfGz6ctB3zGht9FFW3B496oEU4azhSFolhovue+G9wCmHnaPvpUhOZe
CuDHFTPC0axht6WP60iXpnLs4eBLA1r+2t7vR96zWatBYqjMptYJQiSViLTzf+OM
sVg4SbyRIjRJx1FmSdLjMYPoN1/MU/b9NjIw+8R7MnjpSPZBZY4g1HYVL4yMWpDu
1raUYYn9ga06WnK0KTQfivQgiJpXJCuis2CpxPbUQg1k2zevU3/cCIZBZSszRMq5
HfSWoS2dNg9dP1acWVpZeted8Dsryd+2jSjQlA1KrA9c4McjmWCUoacIiyE/E4RN
zW/1GaTYqF98ntSula+X7NSx1E1mWQkPmqKX7E1KRjkoEyj2c1/UKI/oTbgMzk59
T4aviE9r+9lpuF8meBu0JP+PInbaoAF/wG8qPrRdgngemKUvw0O6WRMUZkqRvUkj
JDc7axUGn983hB0rg/enyysUmiH/IJDpuiEYx8D2UVG4gnRq0x8cbAJBF8LHF/On
/Fad14+6ac9ltBO380J5RhYAZKT8gmd/fFky39q9UYlSWYYUB6N5tjtP9/faN7R7
ExzKfiGf/xI/KQGyDW1kyQo4mXp+HS5VhplfSVO5zAx8JkOe+Mi3JRIh66AcwQgQ
NbZyTwVMRCoUu7KxBLl+WrfTtz1QWXHvRUMUs7OU2DEbL8BNKi1lUUAVKWujNyzk
v+iioGJsZFvZNgdJDZCo8yiTyCYOaNz2//6XR2n+fd4tQyXBBQlF9YeiButkV4Q+
sMdPS+KUui2S0/mAa7JVAm8eEPoR5F7E1DJM1P1yY1ESQhUKFgTVfdTBvIsGOKa5
d61hgnrWeJQm4RLdxT30NWQNb0aMCggIShYJzACejPQQUTcynGF6tpY9p+ScFqU8
NfN72n5SJvnjBWQX9g0EHkwa2ybQ/rO0KOhHANqNhfwf1ASX/hVk9Eqd6gOF103r
WZyPaXeKjoZI7X2ti2ns9CFdvVVEklttXLp+K1YwWCp9vopQv4Jx2CMtRIVqsOLU
th7K1V6VP3Io+/KWAGBKEvatG8RJ7zj+1yk9+lLg1mvUsAwNi5bquzCDoQ+saC3s
F0IKu7oQDI/KxJgFHVuuUZ7s0zxUKZr3iHMdef9WHhxmq1iFDARO5BnYfJ1lnsf3
SKqF7mKfP846sk5zdckzLmJC9dbdy2tw23kZ51VJCl/cr8jnJ/z9UtnKm+pXcl9z
Mbu4w3CX1tVqCH0xAZopV9j+nGu2s7+bQ+BVf6hAdi1MyA+ouyMb1R+knCAcaRqf
UWwIPCdgBZmVv9ZZ0A+pqM4WCIfNOpZfbU529ORIlHbvvyZ1MNOH4PenrAzTinxw
G5jH3DS+tvFBxzhXJwqV1bGBZTBYNPYSfuaiCMjjqKggi+Z15CJRxb/MvcNpUetr
pr3dkFGYuRU9E6MMqDX77kWIkFsm4h7epDHeZEGq1VoTSRELBOVDxmkYjSV3qZaL
znu9++CrR4ekn5qJAiBJ3Jr6fy8ZxQex0a0tEy49joF0pNVav1aH4NRAG90TFi6v
vsNb0UF3O8V4Rlg9WIsMui4wvLVhYkoxbwb/CCaJY3fFZXYR/0FWBQi5E0phExAK
LAvRoPcjbbWbD56C5fDqs2wagMu2TdCZuXiEeBMPA3SjItZZ49ljRrT3Ea6ecEEQ
5USNZPDdMknBTpqgSnEyaJFiIeHGXpxXd+XhzRaEppreYUoEGuawUav9jD7jiHDy
+AbYVH5FSihQibExqvBE6YlPxZpa/u6Vm4LaNQwIYtmbCQgnt/io+5BV4LkWy0dQ
V5U4s0XGmvHrhKxihdD1IQXGVylFXFVSgcZ8tCPp5XQ3W8r8eDEvirvE3mIXCsMp
g9To6j1bByT7868wPzmU30C3gAdC5rKohVHdKi2iEOY/m1eCZUE1qabb4v1Xcg1G
uLNDml7bmYWPSpw0HovD/0gKAdLE55Aweg/Of1V3XTZtKEzz7hhpUdpO0UpBYfSD
CHry6CLg0qC8jOPMagJNYulf1nWmxGcVtSyVYnzvKyV7tEQ6qrPtn9+CPQ+xXmSa
9BlmI9rsy5GrTHv3jx+F2R6V+DOhBhFPcVWsZ7ZenTlNUS1+hpzFNIwmsLkq7r6L
/XAhEdVi4EiuqSGhPAXKKRpDQJrNxGKlDH23SzuALqiUb1FP1clGlr8aF31xhkHX
XeErnQAmpONfn8Aed9oAiSfgTLfudl/Gq1DO4LgvlcxkZoNZqQKWrXjBKhaZsJqw
qeOWWnK9QoSCkqiCn33WJziI5EO6T+zNpfxY4UFpETMkw0drsT2ZsGwooy045MTt
3+d9GHEgbA4bRuM0AT0/64wYw6jNswwUloCO5ukoCg1Ji9Wee1NHc0gIMmgMQ+BM
0NNORBBGSFoU+PsrZ7eI0g4WChj7hH7YYLKJLEzLWAs6bW5FDEh1727eMtpL8Z8k
+MD2QwbVgOzEykLfIptJIhfqA9MFCH9fWHgAQA3dWo1/qNswMF9p8yx1sJbbn3qJ
ir3QKXepY5n/4Mb8hrrIx+DdPq52vLAahDGeh5G3u8iTz1xU3moqnn8C4T52fa/T
+chfrW4K+XDDaMzMZ34r93RlorlzqiplOPuIo7xTq3Qg3o9MUuYzVJe6Wik9+xsh
xjacBikTsH+5jA7BjBmGAh+8d+4MPdxmAqtCiV27A8ZVnAX30FXO4X5GVKwIb6xB
kMj95T8ws1ysPADDU0du0+hfLxiIjfE8nyAmDx19VK61g/tKIv7/ZDn3W/dhKHHv
0dpUfYRzuwUzeFpURb5M2b4xEDy3vxfFDswL+U4+hPcBjsIEZyNdeXYzmWs+EQBN
DrP1ApqyjUv1TobsIBePHELjhbMutXDBt71n7wPQbT4xZQpjvkgR76/FxqZ7groF
tP6in72AQrcP9rJrhufDrv/fuYMGO8jGLD09y8komwjAKGxfFJ8K5PsXQ8gtdRG8
mcvxptQInvxhefJc5/sV/vlA2y8gM+UCa7ZPvZVh68+0h5MPmZ/oEY+/kNprHtxn
ySSX/v+W/h0Uc2vV4qMgDUsfVBdiSs2SBd53SCXL79edef+anmPBfUFINqV6ip5L
Az3fmd53214XBQZuoDKxYzq1z75x1O0EVz003xCwO6n6I6hjHJ75Up/ayYB7R5kL
qTD+g+XMpItO/hRVuhl9UZxFimrOCwLNLWin55vcdMWq0EtBVZPfZrlJ2UfmYXh2
J+2KU9N2jKr1fvZmlBR1RLzKThroHLT/A+rZwmjPBp4hIHk0nBFs0WTOvBQXazUq
L3wRBDGVR2u8jvO1J/vmNXrSpdpZP3H1KsalFVRtxRLVUMV0Kveoic49u+yQE3XU
ho1cAPKKusswtea8XZhFqpWS44xx/SHibOEnxi+Niy9qLbENuipNf8l6NU3Q1Pby
eE4+hKf2GYRkQbyWMtQmKmMD+6J1RGj1I4aeFjnGkg3dl3PrACnqb6se6vhYFSyg
i6uNbj1dvY5qgsqnONponSVRik9G570MJHBMTvku9z0uJ4eLlT3CDeUsXqQIhBYA
EfL1v8xhAqLoQNKtUx1a8qJRCVHMZYlby9YOFKXwVJ79mooyKIg0Ry7vWhbYwqt7
b4e3CsgsbW2xJJ7FEBalyJmBjM5vO9n0Ysfop5b7YdrvnMS/PqJVmZTUf3hzVJQX
QS88X0DmLxJHZDtoidCz1e+B0WHOPawItepZk3quFV555Sf1CARJ27QzcpeN1/oL
wH/bWroumIF58z/X68WfJht5iNrIImb26Tdf62zJ8YbFdbgx6+gmi6K1RqKg0PON
OE0hscZAc1j6wNEK9juicaaKeDPpBb4wRA4EgUc+oRo4NB56k+m159LUqBNwQxix
6/Df1PeNp7ew3T3vCDW3z7HvbDbL2NHUdTnjM1/VGAwj7wkg1/hGreNpmVKTIYTL
YlYbvZx6jN8dePcPNfjk64pXDMG9NdmpDDwtNBS8HNNmuVKW7yfji3A1ZkWjtFB4
dwNQdqbb0cvZ5dasPMQlPPSTiliQ7dKwdZAgW/9L2KhrgSJTLL4xHkEppWc5MmP/
nW70kHlok02GVZqjLaxqxBls1mHf0Fl8GbGsuGv5f3UIXn5OaEpsK3WlDUP/Y1dN
1VRM74kA94cRRVriXORw29NPVOZyNe4nE1k3br4+PyTTKCBR/09yc/bvIjzu8r/L
KGUNMjlWafIb0xHjXla5Jq0bplwk5UIt0iVo037OxahepuN2sVxRko2mVSTgASA/
MV6CZ9DbDgIxGNoGL9zAre9YN7qfdT0vuIXGxqTgHK2nO0xMS5DapRuQ+IUybxNY
UKeIpkftHPkcu8+jlNya3W+2iPOMKoMJpd6omwXF7gG989t/RpPiw21HVb0h7oJp
wOK/obbEErqPA+0OuW6AHjTRRahbs+GVbRv1cJWRDMRb0XbnZVa2CWuy7fnHdwij
5YCL3XSds8xoCnAweb/PBVmoKpX55iDvM0sKl4v/ukSfRQl1+TMqW5lKAYHiFuJM
gJ14sDPOE3wITWLS4V8CNyMsblNyPMMxaoTgQj8AL5KK9q+ddxQSqLtObkQ/B6Uw
nMKVrqm224l5R4v/A1ahzBeG2SZPCO9jNg/+SWVr3FTV8c+nkYkjwOBDafsotRgZ
cxllxWBlCYa/s/D0bd6Q94NJw+SQSI3R2ZgFZJzyDpayRQNwJT+5D2rMIZM3fEx9
0AEKQhEOCztvzz3S3SuHoBNwr1x36gfKx5dsq1dyqEb2CAuCepnNCctxVoKTQsZC
/xbiFZkDL7t3npMjPj5KzjoLciEFVjABhp8rAdaINdkzHqwopuCD56FKYowO+n0/
ypmMaefy7ruaEVfV1hrB+O7yP4fgY8yOiXOw2/KTzWKgXTCmwIojucUeQagn6arM
LTiJoAhh4KXfjEXSo1wm5LKoqrQvEX0zzcimCz1BF0iR6yUUr6lzykzZEQciRwGi
M+4L/Nxb62y4BXYfEtiZTqy7NO8u8pZX4BSNn11x2x89Eeq8Ojh/v0+duuDWE4QR
AljmCvb4Y9T5Qa37iPc4085joQFwA4Mfced36NrwdnNo3Ac5KNlgglYpIgCCktZc
sWMXAUjNTfcKBezapr/7I8l0jJFHDGQT8mtb1Hc3sbf8qqop5APahMNRlxSwZ3bv
Kk6bV0+PVYx86mzyFGMEzaQZ5OzWc1oNP1zSNsl/Qn4GJmqxErSI/Pi9sNjin7l3
Mcw4Xafaqt0gzdDSXoT7QjdYwS2p1vVrPh2CZPHoxOZF9b8+cZgKzn1maagDFgOg
2/j2ZPw0vfPBKDKwK0mXakv43J6NegdcexwNHJQtMzAbi+P7HkY6FuKMp+3TfpsB
P0dRdrhUosusBvuWAGI23NVuKmZhLoX4wweC29Wey4nythFGIrEnhhO2fVdI4H0X
m3gzZV/mHmYqA25DT9OqfqO1qkU+xilAAI6jTUoT11kX98unlgzntAOWYoIHJBj1
clFDE+C7Ew3jk70Y5pd+ejZSgGokGE0Sg+35q6vb8YzWyy7q2mjvMYBgrOaW9mi7
/FKvV8Pi1StkHqraNtgmQCqsW3MgW2PmVUChGuxu0Nv8WeAr3cokCKb0XPKynRym
V33Gar3GQL417/wP6Wsucw/n5A4s0PYfBtZqJ1hK5/zRy4cXOc75UPWOaG+I6IOF
C15reRo3vxbj3bN1G0bRM4+39TYp5c7HiDlisVduBtnJOyL8DRxNkcSxhfFMBXWU
VqdIrsRF/Xc3QV1m7SMwx9RCKECuu39RF6Zw+2rUJQfSS/YKbpoJ0I8W3NzEVABu
PPx99GL5s70bjn/BdjZ4f6Fp++7g3USPKRl7/rGn52FASXWaleAj9TBp0q8AyNnp
XsM6ULvkDJkvNKzwKScXF87vv2X9zbhVg4MrdXlPhHJuA3Aw1TP0kZY0qLn7+jME
jv7rY08UIXJfRs1kUPsj4lfmnOhuXJaj6Gi79HNWJc1aFIaAJUKY9x+SjwUO9cjk
arlxs1IYOF2To+JsTCQrIjujmrjOEciVYlgXicFkEUKZZCIZuZf0Sig4JXtwG1y1
zWda54oJdHL8IDmA6I7CRBIvbd6AFJfIzq5Wi4YMr2Rg7Jx7sP+7kQBf7XEKp6pb
8+/Pg+JAcmSeym0PWkaFDjH+J+/pLTNV5m0//wF4l2BnGiqxS3Yj03Oyyp8389rx
E7VbhZLv7ZfIJj3nQ9EWH2QonwmJzhPWAALznFjLxTJylokB5/P8iFSR4nTXykAU
OLTaSrSblN+oJ0FcPQYjn5wqQxCY+3P5Yv9wYPIkDhwQZ/oJPa5uU7zeXqEu3Uvu
FG+XcT9UR50NXXI2n5bqF7XR6lhS6yH3fa5MtPg0+AwthWXy00vYohT5Soy8FleO
O/9SaT646XDEFyO3vi/5QSJT/4KKKQfKTZxHRNo0HiGP1NxRSE0qKKVFaeGPk0tj
LpAszzFAwKxGYHTI6YylrmMlWuRbyhf1j1gZLeDE13JuVYI62f+oeqsxCAjmazz9
oc1yRu20LcXJmvIiElliIas90+vy/UJY93Qn3oohWPYspdlhKiHtX0b1xoMtZX0+
seaC3w2gaDEAquBI86bqx6pkkfVOuut55oLjwlQdj7PYpd4xg/jsnKUUw/gekdjJ
pPmi6cjcsv2YiIfZWyWgqgcchBJkrYbtwGMPSYAuXiErKSyg0BY1MYoZKRpnYSWu
NMs7OH8HKZsDsYijdAZY/+Q1xpBPZMyQ/W8WMKx9X+iFSQRqoJXOLAUs+02atCvN
d4nOk8lDRkrKmt9WsVsXCy8eAb9bgOWU4v3U4AxI2xNkOt88uHYijp84uDLfQRwd
l7c1bFK9/FWWFbx/F0PWUINLTr4RIx2SCNJUeRyBNalF84gEcy/j3XtsSJ+zpqsS
KYkXl/byiU6UMzCYeuSSTgVPjqASM9AzyYCiNTVJVm7ZBuvsffJBOufQF9vfabBL
QJNLidSLpE1fzVIYcAaAncPJQQBviNQPip+a3NvEFrmjRtVLi3/onOjOvMopnIjC
yvv8yH9rfk7GKRQpYt07BbGcb0BCI2TFP6QlcxkU0eP1ur7QTBo38hCSGggq3Ca2
6Z3lz87o0k5SKKdeTt2M6ZkBylLkmPlmM+LNLTtD8jA0U0c2VGoIKHwpjBf0G5vg
X6CKGopO+V5RwPAA0MsPLeioi0g0ps4FgzC0Bh9W8xF4AUpkqGSaKEACZsu7cbPP
Xf+ZriF5iFL8FfEo1C/NhdFPd5mnD5r+Wnoi6aRCx0ZZh4I+lwfVjtjB3JGU5Z3L
6tIG5OZWuUtdVjyMx7IIUE4SaLQXhxQfv7nmGbUalLFOCKq9VHVJu7GHinKHio7f
KyUjXZf+Mfn4pMCSVBS+RzeA6a7H1n6QiDLio4GiRtam1/K49Xvq+lT3T7g7Eapl
T9zW5TX/KZvVBP3JH/YHtuvOAahJOZbPwgPso8yWC/mEW5wgHKeL8jaZxGkaDP7n
MPRAWT8BMQKDViEXZEdP5MhGXPnsC1Fc4F+SN7m+/6h0j0VgXIsjyuULZcC3XM2E
E68I8rq2P2c6/FiuYNsRHn+VP5IGFmtRue79phIBaj3SRujk07erMD1dRXRgnYLA
4bET7YosNnafFM7mofz2DKevHbNIeA4t0rKk1W9sHljtaZb5/ky8kWcTrb1ick6Q
YJXCKAyceaBopWKmeh6p4RiR0xUvtlTNLF1PvIMVCsffjmVZZ8ourBmjHbzmq+w6
STUWA37VPHjnLy7q9gWXqdMTrWR7FtjHoVhewz/27G87pZ/M7/OwDfWbuVFcH46K
B8URJHWPPK2y0E9xVDNPlrvXhWTaBq19blviM6JjYWJqsCMBEUktoiCl2ZSDpvvT
OP6EVjSEqnlupCLmO3d26uJQFH74ufGfLtiJQz2dMyv/LOueK22vcSGQDE/kTiic
V+A/D/fa5yk9CcQPHv/mVCZScxRxhh929SNTbdIn2kyX/v6AjGgzlmmjp4/kwTLI
2gn9xA0OQxgHzwGtRnVJjXEjvKQrs+aqM2viEIqSqdGb1J0Fk6oI4CvRhnbxFRg+
ATDhgz+Tr3cFu5VgjOlV/qwGB3BsXDxVnvwVe3dfLnMzFb7STiMBL394f5GsTdzB
GZM5UpNSyIt2jIDc3T15CKfUNKkZalgjEPpz5RWW+WVkTHZtdm2hsmeQxy24qO/r
11t5CBYja3++Ui2dcvDtBIQmeukjkgeJbgMiKJw33cSgufIX/qEilkWKXmyFffA9
wwbqEKCCrRtDDDJcZROOSnrOxikfuztFUjtXRHRZg6uV1MJRAjSDF8ML84CfownW
Eaid7E/WMJFCOyYLnXbKcmeheKPmiSp3so5+HicCjvnjyo5Db8uFhW5SmqjDmvEF
5GF+9c+DNaA0s0ih29KHGdQ7mSsPCbZi9aP+I8AIz/cfLNRqfVD6o0DRkbkKXa6k
OYPOR1ZxTTZ36umETE2RwOh7kUZTT9YgOJs3QkStDnkmfcubdZlr3ulhte83wKzG
+4DJYetvxcjJ6a6s0REQ1RDTmuqGNHL5/TND14RUM/TRT8KXtYxnzyIGIMYGZ/47
ZvUDWLum9DdPuPJDK8Ddz90AGFMYtV62W9ZIbjO6R4I93E8yXt8WzgxXvnyMJHuZ
Y2y17dKJAA0uleDxh8qj1KyftscsLr8fjzHQGVVDdc/vcwePDBTp8E5J0qKoL6L/
DITpJuAspXYFuU9+B3Jpp0HvE59rz6NrZfXOm3ddZfPKIBTAQgERofcBXTvJgx+P
GGWGqDHQafH97CYbnSJfm1w/IGcEgWbdfpXmYmZvDjOuCrp4t0WzjPLRchIaqwSS
8erBdYBVTtDzLKV7Ak7zlfQFbdeLFt1KA8/M8AW9vAwYMB2GDoke3W9HslOB+kQX
y6jTMVvd+Q+V7qf6p5Bj0b4H4cHntFC/hrDJZXcn2ctfW+KT3rnm/MVZk0+zgp3e
u98I7+eNUtK+tyQhgM0UqhoL9v9iUBF0zswxBBQc3adK+Q41hkrlE4DHLOH9FjyQ
sz2PQr/sE7HTJ9zzOCv/J17pDG/sfKy9VQThl9Bnwr+CT7xPLG0RjH/qAU7vXiWi
cdX1ezXW5G9+M6MYQcunlcb9pnvIbZmPgTCQyKa2yssn2TCPbDIxz6Fg5Ywll4x9
YrqCLV0N26dIxV4pUzKbdxhWY3c11LZ0oCTnWyZU2vrvoX2LLhCJgqGrzU0fkc3R
u2g7sh1fsMp3li3P0rLVXLU9eRYXogzFMq+xOR9+eQWUdvTyj0NXq+jI/UhgLc7o
VvzkpdT5s/ih309jbYfoMpvid0cZEkSPd089ElaDy7SXXD3rxTC9FdXf3tFY1Q3l
LIKJlfY9mpSe29KY4qJonHbiTn4yr/MYCgkHniBaoq94iTIuFjP/zALPbTqudP0j
ZyehaTgsj7f8xP6x8tMCLoxKrNi3AiQ5Z30cFL+GJs/DiUc5yCBv9PZJQIYJ//kX
KFA+xi5WXehTvJBHSJTFPBWxefxlI8ud1URiHRJP1pNw7Q/emduzaA/kueiECZxD
V0ebuQryFN8GEyb40R9Ch4lbgPHzGF6iDEa2ymR5zDFCvw5Z/Xim1EQRZreWJQkD
2Zn55X4/a5qn+GTj7ldvsig9UXYwwN6aG/FYzndb4v36TkxqbutroLWoCqCgQh6H
/6gIkJ5mi5iNBRKuG1FaBUhAAIK4j1GgrxvOL8kQm4OVdbnzjaB9TQlyOFLkJXBY
QEbDoRBtjV7L18kaxlFinntjQxsL8dBOPu4BxxyqMw4LskUtRwHz7M8ACOVPWBud
Tud5vLoWR6h/xb1M2ZuzWKhUDuO0epLmIA89B2vBAPNkot1to+upZlS0jhUIvblk
eUOgoz9cV7o9ilLtZjwz4ZP5QhdiQEc1aLpaSTFL8ZtnnnwViuakAlbj6HgC4m2s
SmX8gLH7BS/khA0QBTG6Zf/ggwNkAAUtmVhWcqG/xh1il1TBcwHUGRGXWioJhiMy
BQmfQ5mli8yZc34KAEUhkCw2u9ZYVMp644kUllqNO7rZyMXjUqPuugmr21EIq1Jx
3Fez2EmlwdhIGknKTpQoFTBgOlpJn53+HrgJif44knKCYY97tHN0m6QI/ekqRDud
wSUJydkrQg2xUSjBS0aGacQVzIl2Oz9KqP23gk/OJ56kbiPAL/P140Ds/TLiSiZy
5QJsAW3repKMw5lJytU0ck6zqnuO+w/kAmcuZ9C7dhqmtHuFBzR/alIbVzWw8tk/
XHS4c4oEbZXK2qAuagta5tMsrLzfmeoCHBueQvJ+GcBuDQykea5krt1pI4SEckhw
tQcaZ51KEulvHqwa2xq8h4+EwBPLnpwrO9WoaaJ4zQbyoffhy1zzHmhJmadDfJu4
l1i0OFVvL9snLYnzMXDWF5NXl8CkBgzR3viFrNUqE6sIeBaBvhjGF/zAB9r03s6f
KDAM4fPrJ6DildD57ZXr8r/VuRf3+AZjtPvz3F80tqcpftCnwHyQORiVnEapY6mw
N05T5tW0q5B+z2M9QUBwu9LZ4JgEk49lKOiCGsdiodeTar2PH77Q3iG6U0yf/6z6
PdmEb6NRUn9S9/IsPEovOE7ZqKwNQvvby3xTeDEqADAMOer6X+RQULdhhkEelTYl
LEi5uGfjfGKO67NE8ccOqH5bzP7vf7aHqI3dLHLJjcbJygasVBi17nCFuRU4R5pQ
4TOsyMOC8VinR4DvCmxYNJiLXGT16UdsMymfs3A7xa/kTw4rd4PzJB39Bqqj6KXd
10V6onkM8eMZ4kdwW23E0BM41w19yYNSwaDSkq5GFxZbfAYZ8Qwvzv3kpK7N0+R/
+hIoGlN/OqJmK6uR8qi2xt7Pf7SOyCO4Pbs115Ymec3URvmuxbupi45cipZVJUaJ
sOwnc37dhwZ6Yj3Og4BEUUk4Lu0S+xfPhh1dxh4WrTXL3lAAGBGTZhzFtY+8RV/3
KyO4F8IQR4KV0mRLO8hBwPPaIEE6nqmDyBW0nRr7JdlKxkpLYUuecW4loXOQ3Olw
SRmgWJPsctMxF2jaVK78EkOFc4c9sN2IIDczWjRj3Ed9EkYvxn2UxNl4TuZnf9GW
Q+81FYpfkCIejdxa3hVlgvE+p9cNs5h66OdPqhXBF1pyJeRazCxn7c03ffILlyyY
bWHufuWPUNsPo5VNpBoOqD1SKTdsiZCl4Qbk6ugowetJTnBdvTQRgvMIpqpt5cSU
qrGtgt7uwo7407zYRD16O47OVVV0gbDnp3NJSwnMTJnPwXHriIo+lvF9GxBVkHry
cBsFR9r4Of53vEEot9egPCJwkt9UqLlHAvbrsYGkJj6spb5+cKYIcEYKczKRGcN0
m3PAf4YRHfawiulV8iXEubSd5mFH7hIPnQlotgh4Z4so/HXzATCiSoRhufj9TGJ4
ZSbjmRZzIgTBY8ApvuTA/z7vJBObOhsSSd5SG/IASSLNn0G/Mnc9044d9u5gpyzA
OBLhorWZLEC2R4NXW1PoRpW8qSSrwew8uYym/VIQg6BUJ7r8iNKtaHYL102xlUs5
QfepI6mO+MJ7Cp+lEZBZbrna27SjkvXwV6IxinwbYsY8eT3VudsJtGBKR48eT1KS
J7+mDTrmD7B0shsoIGcfgbxwXC9sA3F5UWqQH0zK4syB18fMH4ZlrtCM39yQekGF
4VllmlV/nZIporaK0wgpoEXckhrD/6RmNnf+Bmg/NLp9xw05pDnhoJcMgjMZk8mv
EaRbEn/jsJd6Y/VurxUsJfUuPM2tab/uSr05XB9atUvCCZk6ph0s1budDnrCYlTR
zCnsRWtT6esMEM9hzQQBgj6Phaz6apA5CQM0uoAV3CNqWSVjMGjdpZvLhKKnxj7J
kq8vgzOLOW9VWveByjDUE7x0s71xTWB4STcPnKwy4FSA5JzkZGnPmgjBrQC/CR1d
QUC4NPCgh+bEGLoMykvwnQ/4srwvfimN6eYsUrlFJcF4YpgsmE8wQlVxP2VMgdmH
vShRtYS+NlgNbig2POFthA0xOce+W713Ow+r8Rs/qkbXCc55HafkKmmP5lFWlmCr
fZlvHnPJSnB1F+ew2U/HT1sSd/WyPwxwwybtHqeMnwBLsUPmv6MqfzC2z1l4dTYe
/a2CDAb42ucYGOHoPN7dtA4+IBSr5vBtd0d8cnDAqmTUwrgTb2I6CdJJ+2kPPbCI
6ENu91qQ8tGD8aMvyIsNF6U5Rx0QFiEToOesEhWfJuon3dMDMBMid4j+CPhsfQqR
gin1390WeGTTp7soFRXY+FcupIAki1tYIMJizossgw0BjgNJdP7RE0VGMXt+3aDr
BE4SnhdYbRAAxzw/rkA4DzaLZ53N3NHaWFgB+171TQxb22daYVTk57l61u0xG4Xd
wbsO+IyV4xOli5BuntLXSwZ4OBBiWs3oIAvts1OfC6C2vuXNdx4L0GUMiImmn8M/
/2/B/pWCXX+zLf7bqVOJkYrkQpHY+XsVh5/7OwCivggp8CTfYiYfUt4Ljgmd+NPC
BGLKEyODljY74Jx092ThLTezGh01bsAXdYdA86U3vZY7bJ2ZgoNLCYuIMdK0Y2kE
5MLTEkSfurfN1FaT7qFSpEtkDJfI8M6TYlF96dMshD5IUF6hezARhFT+ZWvSTQp0
O7H347qnRfG14IhYydw+62CpGEmVN5ocu48zdIlRn8PI0y2MAyHekDzqYyQjuCjb
4dFNn3EB4hpnDHnDFYAfHvGAfMw2vaUubKgovZrVzPUEl+nxAx4gYboCtCnoJAzj
GH8JCJlm9mOFhq5pIKad/crGGM6M0FogJLan1PHqYe8kO4LR8daelwx+h4wPK3oG
v8s+J3IqQozCuWKhl87D61KlbRgptJRQd76Q33U08gUiG/WtDpM83Ht54fOAoSLK
emmks3iCRVaSq21wtvGkHTH2OsExKdkK1EGSf1PxpfhthCXlNzfGTOisnR2FAq45
wLgswGgueZLSnXnbfVi3mLTmblWL5cGIZbs+r9E9VGujg4uAChQsx+uj8JgnOsES
zq6hjulCWdDOalyFBuvKJKhtNO+0iYuNJviQ3/WUxYwNcQtm87ZzV832mDdAuTZ+
opKzQJNw68MjuUPzs+E+dnKbaYc99vnMZtzUQWeo8hw3LojEVOIeX1qSD6hlgWIt
j0qmhD0acvm87GtlPiRarmnwo4lZfMXhyp3sVnMjlN0mv3jtctsxPgwIWEyl/anO
8W+uhKv1mz9mykYVQgiOiYzIWEGGLmjouDK5uv7tFdbzPiMW8mQrypOih/a54FUM
Tcas1FZFnYa485E/BIJMCHdsRfZgIpn6KvevoSjXwrtneMGZmVp101/od5g1d/Ig
cEG9FVLJnXWHThDj5FWHrpPdxe0uKRrCe9ODQU/GrSA66eMjZJn5RjMbEeU62UGf
sFVytymXCRlon7i6kHqg8kfQj9QQntwFwZUDmEW7zW4/ZshTumoRqZhWd0iMZKlR
EPGHKBmTavXoyokB2LJR5jS3plWmSnfd2O7nvzZNplIEmDUUg/jf8gTWAGlPzV2V
6wDNGSdiv+dF6qlcTKoj/NQrGMo/ITicHaBNQvBxyGBnLyYe2BUzK+Sjvh6UuWHK
7h8tfX4xZQsOVxu5TM+ChHgQ1AqLLTgD6s2cg2CY8zxBztPG1EUsb+Cfu6ca8Zbe
bz/puQkwf2bMKbwposqmSJWJZKJK60e2MllHd+9WGb50345qP6vEHiITSk/UdHFP
B+ALLKQg8CeBxHGTThp5VAbQFoeoGDqKPFwgOMf9zegvBUYAbfkgl/8A1kTd+Wqb
i3scfzTVxjg2Tj/jb03MUg/R/K6MLEZWlXF4rvjcZi2Xq9vYnS7mVl1mXvmYc4Fc
C9JcCnjKBoWUuJ4YpTCDHD/P6mUHY32VmUf+RPJkvrJVWctCac8W0KgClz0RCCPQ
BNJ9/n9Gtg2ApULONwa0xMUIB4H4Gys3ScwmEFfZizf4hBOrzzqpEa3aiwWB5hMP
IhdKB5K2IuAX7Cj58rdfOctKhlet8A+M0aGeZg9nypFu0V4CVqnLoO3O2Ouk+v35
nn4gA8ya4G2EzFKr8XlqRK7GZGe8ZikiFHLgVeGoI2u8ZJOKPFRVFzhP/MmB4gEB
q99SWjqHtXIvFwbam2Zq9JeXQo1k59h5rpAWjHabDXBTXEt8AnJGY84RtGB3+BMG
yfIGM23CgcOlxe0Nb3GGAbvXxLtu2bW0NYrWHcLoiNr7rFT4dj2uiyRzVrCMEcCR
lRIydRFjLAWQPa5ryI5TWsaLc9yfw85LI12QjYTiHRoDtuGYHVpsZAzQk1kkz64t
mdatZ2NHYhHjkGQRtuVAKcPddVqmYzYk1MiQx7DuD/4rHsZsmwcRs1MPhLdl9Lh+
pobK5k078DfMdIl08DmB3f/Gs3rZ8yxLTD41zlRyB5GkRUXgewOw/Eb8I6ThI7Cn
7Xr+SxfoowY6bk7zzP9bmqnTx6fU9Zqbr3Evq5dMsK6dYtJ12p1BWIAofavOXeE+
7LNRWHuba1ODJPxvmIJDMHPsTwOx7x9mX736U+souFiNzoua1OuWNmhwVe2TSwXh
AzPIThPICiZKP8ug+hlkHtJRNH5SSTJ9eRN1FlJZkm3ggQ1cZ1agxH70UKl8K9cF
Iv6wL0n8dUllW1Plofw7Ij9yHUKqO4CNHxiagir39Je9j82uOuMzac42RY3VFmAJ
pqUHBCyjuql0Pynbo22pJwVpiVcTF1ya2Dvhu1ZtEHeSCNvXQ5XJEPoogegY2gEj
9Z8Pp4D0MKeZjBcTQjrDIJWjNMTS6YduwO87P2HxhJQzAMMhio7WQ0nMXz+eNyyw
tp0/6YFE5xHu7ChE7egPs7WLq6elY2azK2taRwOSsd9T9YUYIaEsW5H2qUf6h71d
HPTdPSKiuw+SmpsJRIyVB2RfL3LBk9vRGhtRjfc+ZXOxscqhkQLA+/c+AxGcweU/
75wnlehAgDFtl04DBf9LHRMbG0dNWer7hRLGprPI7ulvfPPBE9bF7XTKzr8adnPf
5Iikvx+3Cu2rBI4BMhDVJEz+EEoG7URePaMLQ3z6y90ToMweauiliMHnDKHs5ncq
sWSHWlSU5JMIo1xpkTOgyqX72aAVhElkIZbldP0K7RkyJoeoY2Ci0AIZZYOIWXlv
tD0qqkrJJA8dwDBgacmAqwaVnjV000PHqA2Ua3peeEvH3BaDHu1W++J9d8riEILV
l2l+NbF0ecqRCkY4C72szvW0qy0h7BH7o4KFuzdC4IQ6wICAWUUuEdjeFl4kSCI5
SPj5gMLyA1xAlfoWd31b1Cwb3I4iBdF0PvXgshX2GC79hxeRiL4H/DKRKKd2kzaI
JmaGz4oIjaSRJB7UggttrDF/gvehNKUSU7I2WuRn6SVgPE0tLJka4MEJynANM7la
CivMKjgouFG/gp1zhZrVGuWgngLYWlo+HJK9IRPrPZixps54DRNW2o3vcXCsQgmO
VgMCkN+iWIpf+P1E3whLZ5E5ErFEP5ZJhbx6Tb0Y5UmBugZOgfsYGbV2ro1ideZK
v647399Kq+3HoyRjNYGqka07/rJFdE1sIz6ZnyB/f1b8D+OLYE9f2B9ZRg3Regq1
YqmLdNGuqeIBEtlxD0Nzjhv4FP2M11swA0GDlnnrC5unNZfkLBkp8H7J31JCMzkm
H6b0VyFK9a3jEaDpYC1nJ1ZNuFc/8C01xoTb8LIPQ/XT30MMK1FNAbQaoKarn7Fv
oZ03rahMMwCnlcgTZIPFfn23zT4xd5uVdeKx7fdE1R7rldr5YHHJ3det5jYyRAC6
UOg3Sue9xHnVMgb97JEyUX81ybX554JJoWRcU2TY4fPOjvOob+Mbb1IS9fYgTIlg
HjaH8o5ZKzOD6+vS4kJTYV6zYtcPs5FAL5hv75V6yz/I3gxMON2F3CT9rh/lZ495
fCyhMBH5prrh+TsUzPj3W134vP99nQnQsYu1eCnMYT2RrruixV4aTWafUW0hPHMr
PiTZzSrjZ/KmZEOUebToprLL22q17aMZfAF55AQCbJCYpr+tK82HXmUJzeEPqI1+
/AI90idE04lMZJplXHwl/bvFOPeAQ1dVXBC1mnmvc31MTODEtW1Q0ZjLFtBjFzZd
mOXmpucLxX7QvcvI8CHFbZ2aE/1feVPYPpnr0T2LstFd8djc0XjJ67IOVfuzFkhf
cq7TYVumvxX+yN8MRU+DLbXTIunEZLDfcRNYuqStbMDWeiWh6Er12dJh1KV5w3+5
BbLaxk7gmAr4Uw85zzAgIHxzszLvcsj+C/de1UfI/U3JS6WgMbLXejFe431psbvC
dmmjUetd6nth/uycwuicBVk2xpydAUolFno0VGJnZFaDDpks1076jP14pX5KDYeo
GGEwSz1c5Ra5aaQQ4EwXZjnINsHHImw23q3EEgMlHoE+TT5nHtSkAuNrEKWNTVuh
CZ/7WHpipQYoMQr2IjZH91I3pMoPTIN7E/jIxO8B9VAS71US5t/3V93kLuIpLkY8
CM2kSgH16TOI6SjvQaGFUQwzA1anBAy6cG/UiXLZo4cf30A/EI0Q3U57fsOOU+cw
P0rLMReQPNa0ISS4em6djDdsaMdxL5fRVjpfQS7dCtBJF3HSnnd+qwJctX8OyG24
mKok8s5Q3ICXeqDU15HcRgPB9K+3Gh1Yq0O5OZMfkdUIq7IS9nEvAzKACnK+goRI
DlgTkbp64h0+etN2zrCSWJ9QbN5VcryYHq4bVd1bqdyrTuhjlsMvh2Bq45P5HCa2
KtaeDHSiJNbm1x5+PeXk4q68/piOdNA/+fiQYxj/f5KoD6Rm5v2bIa5PdUhes6oy
+tnBLz0VVc+S6zakKckSs+Q6Pn9ZFSgX25btsjErEQEnTnJxrFIw3bc9RRrR/DUf
DaMUyroMeptP3StzUDPDDYYP1+DXWLl+z9CyjWwURMMfPgNwPeBwWwR70wvuFh/L
lY1I0KVY/CTz8a9SM0YJdS1kcMCjnf970yfa/JqfJ+0sc6ygWIM1vUd2PC/ygdQo
i3QiILnKxGRsyOWpFYpeG0soGBHnq/HNrVa9V5Ne6sphCOa3exI4KEQXg1lzFa2q
lssA+swDvWSC7HnHpfIlmXSMulx/pxf3cY9P6LsQCt6jB6rmk3ftG00IYNCsW7YV
dlRzCr0hrEEWhVM0Ht6/Ku+xBoepMEdjepnxyE82kQa4gks3B93bLHgTvRkgnCaz
TRcBjHZeuOwrujfjX1zVUFrWvbj0ak0V3lSbMhbol+hc4EHlZ6PdpGh+PDfnVUiI
YKz2U4ZaEaGDhHjulykeLTle3fwBAwovDEOMMgs0ig32zBAUA1Eelwvj7ax1jONQ
SK3EgOUqKBqUIbAQxRnj0N7vaSP4VmWlpGEKOODY5z1A5k5IHzuF9HpIgMF9JCb6
YXyEDCSQo5bY+ssG7xNBF+oMvbE2HWAANvgB44Rk0Hp4Lwjuokc2FY/0r4D3uQHq
93qIn2M1T6Zo6ziehvroi+GYnWHyYRP4KyqAefvU2GcoxKWu/uJxxPR+6qtjzo66
lnwf7D/eIB7raOQbq5r33FssOAgahjmzd7EKvmrAo4/Erh+EXykEZlgRSOS07w2+
9oWyoUs/6fDaYToGaEVgcsMK5VfSE+sHboUShiSIwcBlZ2/hQ9/gU+S+z7qOFhdV
EUssildD3o7X5Sn/sCjdsYEAfiLndRYIeNOR6/c674oNN3aJGaUa7myx90/N/7RU
Rlm+DBKmiMLOy30yNmxOdeQg5XDfIJUfidWbMQMluFaibhtltdGUis8UDPIT2Swp
0wNxPiWF2vOBgVsZD/sscOf+NWPjANRXhyMLvmq8a/Vb4a1OeAgtb6Cm9K7If6yp
Dhq7WKxykvo8cNN7b21k904+DuUd6wbbaHjNZomeIve6+HwF4dKWS8hldp6GLCPt
cM0oC+1uOK7IMp3cv/ETo8VYeM1JCU5NrRo1z2eIEgTMM6QrPCvDWczhB2MdaQQj
iWVFQ/MFHS2DNCRqVsNzUiLZt6ABjCyDlRuVy3zE8KBgnn+eLr4VePx+W8NpHl4K
IdNugyP0ZsFKgMKnVLcl62+KJ6aq0t7Fe3PAeBe9b8IKWJPW/LeGsIml0Dw7+onj
84QPnNIeU4GD37LLwbx2dHoN+/LxkQfaV8RmEZAZEFjF4XJRYp72qSSST51i1DW+
HF1orh8T6X0V4ZYwOZ1L9E+nO2++Ah0fulVv26OVuLkjHmCfdTURf6OcVb2SNt/l
C1OOU+UnQ10K5I2nnFtyGnwH2vV9SBMeoezDOJS+lH5RIrsczumX1VtM37wIaTHX
JkaiYh72+Sk4wJ5FEcVCNXPjKKQ1U0KyEVL0WZ64mvwE/UmtN9UbJHUGMBuFjYa9
wzewg2wEIhf3Az2iRO7sHo3ZRNVSlsYq8lwjI2ZGNgorlziKqPFaXs5NoTPqMQVq
j8ga9g4ln0nBlAyS/DrNqrecucvcaKMTO66ydbMrZ5GaaZ1OFCDnUl6gjdW+bBpb
jaVKU7piwe1BtnL1y4T+2QhMEtB8/Q0tHAG5jM2h9Ill++9+dQonc/VD7a904ygy
O/jmOWVIcahLIrLhYWrSUUIcBg1q47CP7jxJuxh0D0EndkQgvNNacGYeN2L0imHJ
a2ZqJ8gElPSCgexAnO/754P5vTHsGH6DDpf4CnW1OrFmhmxSK/xFIGBM5Pwq+p8i
3qR3sNhjCsbZ2NH/GtNil7+e9sThtChS6IN19WnHgku9JzsBaEmF7s3X3L9yxr4B
xMLgOALX0hp5JjrOTiAcgQ3JXAMDKr4MewiGV6c/98i1i2A7eh3yK+WuDqAP01TB
e+drh7CYuSylBsC/Hum+8DzNgfQ5uVOTIWWEwqDOnKfGuwlVVl3Akklvikn9aXTE
l9LQdGc7YODvVPzGnh5HpNZTDxh/fzp7K5tHSuuUzzd9Mm9SG+crS2GqiqQjLI4c
tZCJNfe/d+XZG6nqFNpczemxv76nsFmdEGIUuTwTSIV3mRunNDyyvy8Y8kcbNBq4
Em/x9aChQFG2fMswNYbPIGQoBAM0P0k5wv6fbHsXewyDsgHhEiP40lDc48S5LJ/f
iaBP0nye6Yv+5YG47HGySjL9wykde9cswiQzIA4okHjc2qirVJfZtcoCJUDhf/CZ
+xbMnQptCcQSA0dA6/L91ageDx9C4Cuz0KpZpoxVUNJWJe1Y86+i+jVOpYDXQNvf
TeFyPXEDghso9a2QcUxlljZ4Nn7hO0dyoH9a3r9fSIcm60CcXHxsWEMXfRniXdvJ
RSFJZ6gf1e0BVnXe3lkBK/13m5Xp6DhFIjakowVrvnpKjhjdi44UsNmIM4N0qs3j
0gHrKLCopWq+qDYj2U8uBODAYlhyjEKukwP6I1zoSKUs7WmSREwbh7NcrwyGwENV
AaPpCyyRcpN+0As3Ahl098si1OtAGnP35jA9Jpb84oO2G7j7LFtlo8VOaI+rHXKs
OjO4QegpowzaxATWyAaA7c+sDaz2ZiirVwVuKUwJQCTtA1W0SS2+ggvjKUMZyfra
h+YdHAQgglUM+UU3mzcFZBncv5RHcEKZ1kmxvjVh4eotC/5CFXZlOhknHjPHhNQJ
OU7DwIEEhL/WsuerHP+MzAd1CVmX7dO/O8uUV+qQYyUWQ9yEpe7Pzx3JrN/ZQjMC
6FqEU/5i+puzdZjvwec+zVtDOAklXePCA7TIJho2XR/gU1vEVQnEkRfGuTKUVLqU
5OmE1l/JiD6qgnc3FkYeb0UNgejN4t44dNkxbV9ruFdDxOcvm1blqG+Op7AMwONM
aL5aKkBZurNmKBRoNOLHJdzk5Irbjv5/FQieht2OZNBxXy9iU3p5mdMPDp74A/9f
/YCQhJ8BfwrIuiFtRlybBmT5kgQSKzvagQa7RZRgRR+OcvWxdVvY2mxb0MlPPPyq
reHXOWgoxcoi6fSCgDz9Mq1pUmrB9fy8kdMgnmnrizdMC0H0Vjo7Fft9LIBC0Nr+
qHWUHOoQJZZjLoE4vGnjZGxifd57IbC65rybdg4KDA5x9YM4dsr7m1j5Z9U5e+hm
NQK923986sGJ8gCQemN55dYR/DBMZPeBFdYQHMLwW8YPsZaSVQ3WDLnF2Efd5fqE
JisUMqxqV2TGEu1sLbSk3JrXPgaRP2qbYiYDpiRFlWYT7TdPT6xhRhwCJmONJyuN
hZd+fRV0lvfTKDY75GjvlQC9a++j/mn9yBs0fBthOb8+CFu5sKUhjwOyaTe3Lpwj
8ym3XDuYmWpl8OP9DIwYBJpS1AfKLM3uhdRJNDtmERmRMFMWw9xc2uhfiFWMTxvB
235BjppjCHBKWkBC4YUoVzzWLJO9njq/0R6Hx4QLH4+3YBMDognpnF3lvIlLp6Qq
m/VZdmllQ4pUDuVF6aB+MtmUVxkifXPtFEow1JuNeRL2Q1oQqYarPE1T1KDrHY51
HAytFybiwKtuxjlvu5zyW/niX9p0/EQJ/dWtNTDDgRsVm9M4LH69tkT+c2SomG0Q
NDXLYFr9IDxG3NbKgX4NsZG76JYR9mKI7bV4DO5E+Szk73EWNdkkseshgcWNZJEz
VL7WqyF6+shMjf9BM46kdByGmSOSzgYRxTWUO1SeloKLMvJdn6CUv6FZ0z22kdem
tj++eoRKHEKy9eFOW9xq0D2NleolrH9GVl4owoT+Xo2MAlt8MJyqU01uaot+5z9G
vDu2Xh1IqkcNpKcikQV8NQPUb2T8gVdibukp1sH57CiTEMh8c3ykP2VFT0itC+76
/t/h2vyYULfoetJtaF5vOiDTuXAveLae619HNPpVZlgzA4rRz6N+TXX/bw9qR62O
LL3zoQFefn0+ULsB71FVNR9+PjUQ0vuigsKJkR9iIj2kxyIYIobOEdRXoFV0ue67
Ebjn+RF+22jHnJJ0dVV0+mSZSE7Hbrol/n12gnuTSrALCvnS+3c30LFVoPL72P9U
z17nyY+xXrRdzIp82VNhK/MUDwLwwmuwE/OkHwaTd3OL1sH5AAeT2FHaqW2VXlpd
WKkdci3h1ikbZrJDMlKSbaLKtu1UYEWqhe/qRsc1qt6eqKX/6Q02QEncIJL1E+uF
/aybO0xcU+YuWVcGTGuposdaJ1sSR1Ad9JByWHAH8gey6p/99kiq8WaLnXOe0qtK
AfORdKH7GvyTkf/dEIgUkyg2mF0UgwqU87f3GWtaDEvcCIyWA+MEGrW2mHWicQE+
RTX47oDBzjQ/ss8a0xGmwJaqOl3m0g0cm23TiY6UEs1BQPOmyfdQMGrB4yhpk1PH
420X5ddqUmQpuMAEqc3cV4iUcyLdx//bYQUNPX3IDZfePxRSfrnfHarBwYzUka69
DGAmgIZ3nYYrNuqtrJQ3zYW3+12IemidaPiHkqJ1Wh4DH1p4R7hba+EHJ9CK4i+s
RNLgUQeQqrIGu0CzICW/uIuGXyCVYZjPDwmAcHfxrpvg5MHEC9PO5f5TvC5+b1uh
/18GC+lrsfrXHBLxEc+zhlCr2QUxpeGp3KdC5VSrHSi/Zthw+/T0HAL8UcuYnwg7
xTOweL7FpQU4yqUzYZwLa3wvbm44AJ9yJ5JZArQV9dCvGRqr7J+pMcSdhz5OPRm6
kdiSFaazNzDt+5DJBqMiOP7gaK1XlkrqntdDoI/AVNnGJ4sOXA8b0TIkx8QIaCAO
FoRsyXUR7TQjrw0MZVG55dBGaOoqhPH1iQ7qvNnW3KbU0E6cPpXFALnUN08jBfG5
IstR+a+4AURQzBVJ0hJMtRXZgmDG1GQedjPwwnjlAzQczWhm3n1xewjUdhLbRIvU
Op3RrfdjMZtEtyXhSjDfUhOrOj2/LUWgIsj+trZsTyZx5RR4SnH4KAw4SAkfYC1F
ryLLvWF4ETO46fBb9XgRTG93Nng++TmQfI4joZ0Tdg4x9I3rncDdP4RlVbr/3unr
w1mAbgJVZtHUSlAQAluDyt3Brmxs7Xx1mjg0IGOWipnDAmUr4XQUNd35if2aKdKQ
tGRyZ0qN4F1coJpqgt2PCCBZzp2zBDx9QnrSVrlJy8Lgmo0xike2DSG0IXWj7tMV
uEAFzVGeq43emhWQ44vgXuYlmjtYrjbAYssITJye6nJIduVs7xt5BjTnzdsyaH7l
NJ/xGdV7G8LDipa51oSVw8mi3jz0KwSgzVC96PZ8Ggk6mqJiAQl7Lmklbs5hkcb3
uL2VKmZWJEKa16cxNTIxoZACP9wpmLc+vbRkYCIiOx1DAlxWrW9ugkPK6bMJpj4D
1gcSqDh3bRxSGTR/kV2nT47S3pUmT0YjWssz9EcjIHFaEiWVsGNA9yhwwEiho+1l
kmJzglwtv+yqEgERJLTGVo6Urk/Kgv8mHkSPzFWna0Q0TUZlro/U2jDpdZE6XY/z
8s7lIlXdQwJzOSfzAtBI69LpCvbiEFujkT1LHqOMTQDzgiEW9eZ9GHx8f+QmM6ql
egw5e437Qq80xD1J0ycNtXXWPNQbI6ISInNjEQwzphP4Shf/HBv2YN4+cl+eOa52
xvinEkooKGGI3gM2U5UR54Qc3yXG1y85bYyV5V7ujP2j6e7HyTIjg3XrUttXM2eY
juXz0W0Su9avn2qYF9E4+LDE2aMgmQs8EpUopjJ3W3642FhmS77xoRDTJmkeF/Bw
JUq2Z6N9Oocd7CvWznk3QodRnB0aIt8nT/7Actc3yMQUfXWzRjy96ti2RCytmDta
SfaKFCZvFEBBGaqp5eV+zvzs0XOBpSshW7uGccKQiThwli62AyXv1xyRr05e2arZ
iNpHwcXqJ431YhSh2U4V+nqIiznEYp/NGGLxn1J3esmGOC1mIk0U60I+qco7H5pw
5S0736l6H0X1ZW5uXhWG+l+1J//0oDJh8JFEKklWn4TkPySuyDUsWy6hqScWQp8W
4wL549fcRkyP8ylTDJWyF6FgOpdBpBIxWPUxDfK/2FHIyuQ/3WRNSvAsmuICuRxA
dFZ7TMXfv7L14JT6FjMIiWljD2Ta04j23rCd1vjOK7CW/5YqTWAVgO2XFiA1Ir4L
HsxYRfEmdp5o8GB5iIxA8uS2HHbcgsW7D7MzaLa0sS1uTgSfc1/F149HvF3yhswE
wlG9c5wrxavjnTUER4BAsZFH5XkO8ZnKaxjmaIrNXmVWjAQP+bTq0OePvJe4Obeq
RvqM836dgPOyH/pQ0PrxNta8CvhXVmWvSF0Bct4LZJhlxHq8JEOWu5aOlWUK2lqO
2TI9sCfoPYNIR9knJuAYUI05E12VCMA1tqXZKpuefwzSzYiH+ej9LuR2n+ePHshz
7Nv2niO/dzMOqRByOSdgTrHU3wHNx8uHlleNHYI0DshcLvByXhrZIk5FDuS16R9b
we1PKA+Rjpi/O6jfL/MFViLjbTq6zgqvfqCF6PxNkJtye/CS5J7Ion+rB5VF/K6t
1bXD0g4ruZn9GPUauE+DxIPCLMNYIfEYOhuWqUsUfCEqM3jsJ2OTo75FqUsShXA5
AzaMrfc4izIhJSnuvy5hCZgkRsLZNmM9hCndf43CivmpeVfk0BcCHf8r8f9jTgLG
PwiYIy0Gu+xCj4JlIJbhwve7Bwkgt2+w/+u7Qs7RzO21hL5760ZdBgwAUr0jlQZd
5WxH05FGJ37vRwBXMboPbQbbWjeGsJp9dpXKRB+NeDs7bBhxBIwR4dKLOQubG0aJ
vU3EdnEyDP1s2Dcr49edaZsfZecSxzIXC6tCqQeu5MHhUAy3BBgpBdWtLk+XSwty
KQkUWNYo8FGKVfy1MxqLzsXn1BVlvXJsPtoNy3jpGa/jwoIHUwi9uo/W7QFmDieh
IxVqRepW6x1m5HZJT7/xFtbBUq1jVBbtxl5y5LXWlX4JGHPjiozoUufnZOTqPEM6
gaHoyY17epePkZGj+Kl65G6QrrktppKFw6kF38RriHCZ2g7c+GKlTXpUXDAlyckw
mh0WW6AuVpWzjaE8U0JkEUvl5PzaLG7iYu9w6w95CUON+3pGvj69uGfzN9LZiAdK
hbwwu2DIeeZbKU23am9LtPpNY0V7nH2sCRTZsDQXLZBNEXbgWddQkoLUeZ4dOfIK
O6Tf++BNpcbRIllWWWni5UWHT2uAhzIJdK8ijUEsbXfb9iGl2y6EcfrlTUrneDxh
xIXsh/JNBvlxQXscI0f53iBrp0W8eRs2PIoVx1dOd3S8sc/OKLbbFNUQWTA+S4FH
D65QA1I234M06rgJ0GI+PaGnZxudckl/Qsv47bHIsi5viZ5WinU2L71FcyPEuXfg
20HWHvyBNjULli9g2G0UipwmQSbJLVu8VSBhwIGcoEpMZeAa6B5APppDpoD12h8A
oiSGmaufbugbBh5ykZdnDmU7hoOdWukEpZUwZQHhpYPWx4C8mlJNheHiM0344Egn
gWBC0V6n4HYJHoYWHFjSXGh9BEigKgU7Tezp3j1AIFev/UkcmgoiCQoYUC20jQ58
WwjYXb7UXtmaMaVshd0AoCVG0bKA+H20CfwO6O/c/5rno19QO5Jd/P8TJdLliasO
GivwBqk0LSvNebQIbSHFMmO/1T0OHEUea+Ad7fB5p3UYVzhvibbbY7lSHExXsXyx
/72yQd1CICWs5588h1lR7Qc9sfzcRxCZ+BLoq05WkcBEcDl+uGqXFuQjthRlSnqW
dn7Qy3PzrqD0boQyx9HTIKjM1VcNsIIa8V5Oreh1s6F6ModiIb7p5Kk9xgTq6Ob+
fUsQYLdzPxGqCNoOWVcdpVs6JzidiDbegNs4TRjcPvb9sNen/8XRofA017Qtd53u
uOcRLN/58oltpOEx/Nh2kFLgoiUDVXp5MQ35DyJ2vV203dt93bRG1cwomYrobdZ0
MK+ctyy5c+Zk3zrWDxsUY4JBXEFXE+WaQnK+0e4OTWfGm9zJziIKjkqprzoLRGQ2
Ohn9D+UloLbDQYz0vL7XBT2imzb/OZ8TCVNyRJRXVrk4gHd3QkJxaijhJAIOpCYH
0XiMxtZutpnjN29WwbVJmjB17teCkFHti/lSWqRmURNSWMnZKxDjlMN936eyq0k4
NM46v8SJMQR/3TmC1pfgt0KHzUzMe6UjBgdQ62cL4QBxGPD+dxunUtizSGLzk37a
ltwABhpeoZ6joae4TecSH4IBCG3MSK0YLjCWTlpqGR8hkb3m2jOQMohCXK2G15JK
ITcur5s6qaxtY9JyL6ECHQRMOhKvWhBI1pOIwkb7pXoaU+Ll75jXyr5ziwJG8QFx
LEHI4hoyq2DwpUQkbeO7LBfDApSyIqmoH/rTtMyHFwkv4UezabBnEFt/iQzdPL8k
xVdKOja8D5RBf9D3LTbhw2Zd7zoEQr5HGBwEK+/QI4e/95/e1tpPuDAFL2ha/7iO
ICWPfAlR2MHoA8sa1CuOznsTYj80WCYyjJUdegP6HYO+33qaMbnuARewJtQHCIcC
LTPl+MV7N39Q3mfsWLhQcWbT61UTT2RhLQRVu+L6eqZqHFxVS84DtkO90cmd6QEw
RXzyWQ188bfCDkovqthxcUflWgynjTXvEr1bxmmUhRSBQU+udv4dCld0MLG46OMp
erM1nelxi2zUe9cbMEwEpyAewpbiGPoX0zGcEGSkDy5Kf8n3h223tZKK7OK0R8cd
KMsa3HhAZH0LJAwSRpAQ3oBaTLYDHA/js7kSJiKJdPP9eJPZo+efmWl4f9GzeX/1
ubDn7UlVKvBJALhBZnvncfRrPVYYhCYzOwN3OixehhCHF7w8wNY5/DSY3Dl88t5c
KDmrA+85fiOV9TQfJqVYIyfywcFdUgEqwBPo4IWah9NAyRNTjy+Ei1HdWCoxlgwB
aUHHF4BGKPcsbhpwtt+6ovMSqDR/pbuLItNhWVhHYYwWcbu3aWd/UmmrXywJ82rj
BIC+rINtwSbGuywn/a4YWzd0LsjFtqzdyO8SAWCejlx3dZ052Ltp6XTx0b60ryWQ
LV6tJmijELl3/HWmbZJ0wdQlhF2eVHwvDPxs/7cRz4gnz+awSjXtXyG+f8WxFlFp
QcN3Kip9cM3j3aWFajwND2OpGz6a6dAGV6OCEgZFbkWdhqbjilbvf+1MKUKDb/mL
/mTybguuwmqV33BnZ92zFXGqKqK/eZXFTReH0FyVhoSkq29Y1Md5I5dtvUZ+BjCC
jJf/a/5zDGMQwMrtAOQV0PsqmHFzNYDpH26a0+Aosg1OMTx4tyQJP+V51bi8uzNc
VSSC/aVn8OZOaG2X58o/boPas8hmtEbi3Hq4YNQTeMoLFkOTWtUi3dcfkiWo489Y
+TMsiAqwjGwea8Z6iYYLf2lUWchPjf1PV2HP3xIrOAuWBWIrEFdhf2gUkPfjlaPa
Eq/657FQpJsxEyvTiclSz7dcslszIDOW2WfJjCRBzpKbQaUMLbi3BfxuCvbUhmcW
7Ds/0mC3nCoRerOEGPGhhTyf1m9xvhEzL/5JIOJx9kuSU8C1cMkPmU2zqyhdyYib
js7CWEZpefE9CkzoJKVkct+hf3l4ISRVBWX28BV+WqMaT6DwKQSK9x4+QePS7Pxz
7D64zRLd9qKWQ6GgxKcBs3gr+VqM0FD79onaB2wo05N9q+NhixWRljriZHPJuPeb
zFfGfGo/ffxvZFktn7nv1d3ibArBxTBjYsIGng3neHjJ5aWy09VOxWFxXa/V4bn/
YwAxsTUoReoxNa0mXWbDyRn2mGolR8xi1W+Mh+p91ui/kjGCaVzcnoBBQNnfHn1e
5N+e24rmQY/0Da539LiXNhxb/brkB4O0f9ilBqikgvivsak5j9kDN55wsaTEkbT7
kIt+MStZpU0aJthIioAbLxeguq/a910M+z8DmsLKkM7AoJY85WRbpENuh1hLIUbe
tM3Hl6CjQK7WgLLEk8LXILvxk3Xnx3z6CE9ZeB7UuM2J7QYU+Zamty/ep70ub3sL
9g81sLNPmBiWFJsqHUUN08t/26nEM9PU99b/JiPKf9WhcglPzXHD8g5gE0Y3A3uP
EnHNkPdOvmgY11RbH/rEgx46o/VIkfiFiD9+I9tx9Az0xyXN06XrOmtSHAibL8Am
FE0bH1VRh4WUOo94WImb6So22rt67aCId42TYbvII5+Xvach/lZGFcBjnqPhMlBf
76qXxdcxiQZt8IRQchJlu4tgAH0KlzdBcLfDV1NIHAWFSUTSy3HZ/cPUlV2PvDiL
b+INkr36vZBT1fSq9tZ1jw6zv5Ep1XT/Xe4mk08j5JxitB5LyJG/wHPZX+IHTHKE
P2vdUqSiv86Qnr/ge2i/P0JzgJIrW0qggpDfqMuXo+wJpeIUdHMRjwb2+KW4BRwo
/uWEIU8AplJ0Qw4MYVXOVhbtvZTz1HQridPWIO/JBImr3yKA+U4m+y1Bty2hPqHf
Es7nhhZsqduoD+Qua4dSwHnP3ljg70+o6zo6DyV2/AA0pw992ZC7XUfhvr+6Mm6H
GNKNcEBreDgkIRkhNX9PMkB3k4YV0UkV9AN3uViITNXo5ZQG5HC1di3Bs8Rileps
qhDO50uQimODYsk9JwBIgYtQ6RxdAnQd+EVjyKypeLbaLEZLq4Z2gISHDSok3ulW
oc2UuJ+3pbjFQJNQ+atUr+2C0s2wX6nDP3Y81qfWDCWNT9C7UahLv6pRkUNlbYLV
lMVXge4ry/gl01YvJTwS29dswfAcNDsjF0XbqqcKvDcOkJr5Med6EN+TjW7dvRij
jVwkOxX2K2SunyYTV/FqVoAT/03247UE8vFmHz5Udj2DNcsFe5SWoJaLDXj5qbeU
Cfor06VhR6cteGQrAZZDbRdAw2Ump1iK1lM9Xu2Hs2nCsOltG2iNeU9Q5h4Louon
9UZZT2xRVP1RgeGWt4MBpvi7gEXAdUTagCjO03VDCe5hTbEqZ9YlC3+XNwMGT/4k
nblVqtsZk5VDq/ESbifVi/fO+Bl02JLKt0z+FZLNEfL/DWLSbloB5Clzkokkursv
wXmCEjuQ9P72HjszvKIvKte/KZEFV/jL848xp7UwxMQswkK8rEPrPmfh0kT6goWv
URkocq3zUNxQA+YJedvWO1lyHkRw57foU1fsRmPTbh0xbpyqMmrR6+diLjmDIeD2
azWekXg9kkAyN1zF7XLhWBC3wzclfRvpMReJMepH9UeHAUrxVyBEOM8MBVTcKJx5
1REbZqB0DdzHCg6mHy7nPt000tbBeqo0U1LvNpsecqDYwOUAgEoibiix9afvY9bQ
J0IaqtwKeTHG2aoWxc8bsrzxo+OvKJiAd0ZSOcze5y4EvulGOHRkJJvHILY5xDuK
mRTPU/tdPghTLF1DqTN7EfSnkU/lNI6FRu4yHDqehspffj2c6ZPsMXex7GoRwAm5
0zjFJo6X1BMhuYkx3KoNsoYp/xygNXfMju5uyXCkofxRud/qU+sXEkWDkBrRn+BW
WM5lNtUMgs6pu/A/g24SB3aPB7IZzI1OqGoHbsbDKtvAwwGcb8YmnMwhcMauoR2r
qcoeSRFgUcDj2LyiN6oYeQvFlA+X/TGskyXgkZpA5SAC/JyJxeVL3Cmp4QH4t1IY
fKHtbXKHVOStYS8cYzLpEfJUMEkMaZ+6wkNuT6VMbEvWOJO39vr06uWeuD8PMa/p
WIuWLE1E3666pTFwXdIdiYQL1d6S3Oc9HxEcMdYEVsG37kBODVjwleIHWTUgIoIL
HEtU+QdAl80FPPbBp1GZI+990BDl8McAtl4ueNG3ytZf3Bk2EgZ26zqoGlZrid0q
zD3Qyy2FeKyCKm3heJhOOVIIIG45lPb9ZL2SxfQHO8YRsAZZGy8AKLahO23suu43
X0D2/OYvmjmOEwD1j4zNUSAgsGuMVmT7xzr7eI0SZ1/DMM8GR2ucY7tIGCUkAg5h
/DBqHkOqL2d6L0CjQkfGdCRY88b1IT2OS7XiZHiPGct2MrEN/8vKlrqV/5cN/cJe
MWGZn1hvqHD0WQE16Y8yUFWqMWcgWkjsFs1sclO9RviGUXMVjYu5tJNrzPmPhl2/
pT7QoxAotdKi15ei8ZmRUz0maNpvEPz0oyraXjYNTfn3QgWs391s6gzcyp/4gYkN
FQuW6qyVvCZZDhSUsaHZ5JOyyY2r75h0as8fVH9AZpVGzI6dhq9yX2tzaaewRfbR
C3uwcVHxOdb9dKpAGuQKV6GrsyMRbOMn4GUHPW4uvNCptY1cVD0tPlf70DPKn22b
AZHVlMssdjE52a+igDU9sIvNvzJRC58FqVD4L+uuo9SWp6WdZuLDxsqNDzIm/xye
lIGogh42SeaFd3Mqcr3puwCXpGtTaVhFXbipaCQQO25e5WUu1lxR4xtBfBJgV1HO
JAjD+YFy77dzFqLVqRAoVFZ/9nnK6oqgvhfHg5fLJ3Gtr1VFb0z54xwCzfDzIx1W
zPHowqWSSkF7d2WjEByl6+cyPcpZXPYQFspHUBkpK30izub+ge++9o79E1idMP6u
LPiIpCplOYg4P/b+CGwuKCFd+yKt4UghK7BRONAM8X3RGgvB2dMjiZOfMhwtUpEo
9VbkJcj3blYBydxvR1YHbia2wpNfTodMB7v7iRVTEJOusUSAnfTddqhC5qF23s2B
eBtNiqx8M3RQYdsHxytF3uY0RXGzCP6C5YXnOzj0V6gKapNeMYrKvp1ZChrbx6qo
ExshPIKQvhKkC5MyadjMNsa22+L0z57RShRDyTheld5E7FZjUwcJoWI/cTA381gq
no1Sx/01XRqmgW5w1BQiEmSSADG5ntClvswHQfHDa6TBhLanDlWVebdQHhGpEvwZ
7viNzexFlwd8Mem8Sw/W2Bz4ZB1euoBHJ9hGgPt0uWQuQyaAM1oFcseD/h3bEJ/s
iVfe1pNcU2rlIUYI301vplK0gE/3cXIYjN7PiXyB4u0EAuwVeMEbeGWnzYa9k08X
niSgB22FnpKrp7GYuLYU5VTqqqbDzqmsyYzzuz23cAlWYvuuUK32YF5xsvi1d/2+
t7kaYFU1UeyOFCtGkG6cCkNxIyI0+hYIwcEsTaVWXk8Vp1nMiY7uUwi8mASG/ycW
fZwSuq23LmEcYGJzvUvQ9PJenHfwnOLl1V+vVQaxtCRnWQxNPF1kgUK8yv2FMulk
mOLwh2UYShjr4KrrcpM25YNSQdkHj7ElK/9sijmTOqALz6AvTJ5HYnkjQeuczABy
jOlg3WhdDODo9q+AAiF52QvdNcvVViVOBvXAF9NqEpv1GXGXedrkyrDaWOa57mDV
kFeFRNXjwIlSPUas9y9LhGLuABpthNTTJNgIBQmvUx06kfZNXOGJkowN8yayU0Zm
9jIVKAr2Up9e5kBsqn2ft6Y6TKaS8lB/xn+NdNvGwJfhdvQDT0iiVapTxxStiRMx
MYF06R59gKt9+CUANRZ4VyBg6Z1mTlv/G3w5PRwccVd4SNKaN0aAk/l4YEkar6rO
w/XdHsU+b921ggYLkP0zqEHpUrnxWKKxUwGkTV5i2st88wQUawYIlrQu98ieYyWE
2eSKQ8dl2ndng80UOccOOx1wSiDEWhjE0bvNoWfXn08UK83992f4n+syuldp6Qrj
VeQimdAewMHbJsrux0XUOKLUbqq5+ezM8zZd22Hb1JSSDZd9rVF55wmuycFY8lIW
j92atsteUEMRT3EFdQgW5WrdpjQxASa5hyO4fZ6UAl81N54YyAZwDeIElRC+vEpX
9dgOnAsTi7BxOnsc7F7RcdeSF4G3uuvG9qWuZBvKZW21DdR5fncIzE6fo4HIZCxA
MG2RKJ8A8F+qbz6nt/k6RZtg53+uIUfqyle297qfrItCdEM7/lIO1uG8i5iif9tY
JF2HF1KFwlJVWiRuPfdQTnpvK1bDE8Xnr7AM41azSFVZPn3FlaUq1HJtDIhFuzWU
16mXTdmL5c/vXHaR9NedeLBW3HWwsV1kS1e+s/QD/lRVhOTZQk2mC+ttkx/LPkfZ
m6ImNYK3z3bCMKpNEaW8ofPOlXJHaiEqeEJz8AariZZXTzE6zym8HBUf5SuN/exl
UtE1yFJasnrbA9xQmjxhHzQ/HxXpFM5CDFnvyj6URhUqSxWoDI0pNsZb0YKjpS7b
882DkVWqnf6I/ZujSykVVcX7M/u+1aRV2HsSa2V83WFj2kyvLioL6odbk5N4gTQM
DcbjbTncm0IZb5yUtJ858owXNw390OVwR+zfnmjdO50vV5Nt1GCfMwRYV7UhfCgY
+ZNdaOg6Fpil/Qtlsv1gQsDMurv1yCqDcNZNY0m38M1y81cr6H6lzO52TSNz9Vog
s7TSlQuDJpnJ6TZN/k8Ec6pHJ440kZOD9dURsidmRjd4/8DzH/bzUjLLHyMuYnGN
7RYRgIQc4Zn4YK+ev3nDzeDD+gy/0QyFRP5S9GspGqU6GkVINqtIu1ogawt56Ble
Qk7swMtKTEWcygN6vSY325kEhffDQwF3RE4fD7I0OyuGDKieKvwM6BsFuM24yRRe
jpnoazRBy7DNNetJp7COQ3Ao2D3Grhn7sbtBxql74EOzX/H4Lv5XOMI7SwgjYHuC
XER9DwFPeiBUkikFC8l6glRqMSYkjb1TWQRCF0KB4uAla8OQezAAzofey9q5ZpDA
wqUiHKBr9x1NfOIcpe3UtNwRXbdjOSrq2i8PflhCngr1wfOL+1jDVkqZ3G9Mr7Ql
IoUl76yDATeixSopg13kBEQkQ1bj3OORZ1oXPWm7k6GEH5KOl84hAhRcXvvrv6kH
yHbweAwFe8D0DyDR8wMrs4ZKFev3tJ5rFIFQJ5fHm8TDKh3fXTRhXcwQXYz/YXps
fCP07MZ0VXt+uH9tSZqxUyfNj5rD1dv0a2MvoKFtHjIRNk6fn9zRlq33PyFr0pK0
r3GHDRNpGTycHbB9WopV+oyl0NnIhUWOwaBSNxuaPByGSZmVG+kG41R6/Ui45DEk
miI1Drwy9a6m7LFX/ViekLY2ElBGoS/Ju83uiRDo/Clg6kYvwn/dVavV2JT0Gn4V
K1WHpyu8zu7YLL20MvZygosrKtqd/d332khEH/iRT9/LyZMvFLEkH4bNUDSIwSam
62cKHrMRpvQugvQzM9iVQ6kfDPGDbxbfLeAKucNkn8ooADGnwMfm/wL7z8bC9SA6
z1b6CwE3xQhmFsrezZzqWz/FRB4whjBupmt4PpVSRqGSvXhmf8vSEAVz7Fk7rdTD
wyObR6Ob4GBi4cWmFWNtrgOkX0N63g7wVL/0sZS8QYOjjLp0wIRI584i1CsoXgJ5
ujiEua7J/3lPjVGiIpUuZQkv+F57puarHIV90UyPnDSuR97n6sgvgjX+0MVQPDdW
Pr9OrKS3ie4sAF73PJAMX+/6rQ+OmkxGbTcQ/+z+JDqx54kV4nVf0obAZiir+CW3
2eUQf3pH8CAlzjFYDy4cr8CyeI88yUuET7R7BV4BEa8A9Y28jDlu1vs/4Y53DQqj
vlYT4Ma1hrujfQpPfmZcbmfxJcF447L8arHmULf8ySfcUgU1SzUFkO5geWnVq0xy
0wzDxng3hauQXtYexdd0VoSbkz5VwX8Hxcaf2vLokhURLh+y5u+rdZHbz6J/yMWL
E0s/URsJdQ5hq0w4f/vD6LZeXWbp8JLqPCx9pjqZWIzrwsjDTYt4BR7ToCXQ6P5w
c6ya7YaJTKCiIE/oboz2TWDEX3iA5ALVOULtePODuQ8ahx96emJFOlUXJRI7JyKy
MZBxllqfU7yq9EV420CR8F9FtZicLPv/VDJwyrZcfY4JEkEB8ewBQIxnXPJvTK3q
mz1sziCk4r6pvs8fVJOsDrEo1kSpeQDDyMgBZqi1iCCaGuM1H9H+UhVZWQZJUsET
CLjAeAcgKpQPCza0EjYBNGprVkt36zrRSxCgCLHSwlj1PnfPAgNx+8mZnnipd3vB
kSRk7/5A5jCxbhXLkvuSMuUFPrkA89wwHRm+ZvdV8yBe1I1MfjPMrDjN9N6Vms4S
dA4uFwl+/1+OgH7gl9raK2gZUi1BaC1sV5MvBrE/uoFdOuIazOuw0PKczRmeGhNW
i1QhhI2tfati03algkHGCnH6brbNTTnEsJal4q/4lZsG6aCpS4o/ixDetuH+6XP4
DeJ5o7ayfvqI/tT+JMIp/pb2ryUnVXIWpdYx4eX1z6FGQqMS2NqRM62TxC9qXU+E
5NRgj0Jx2rG0vxiAjFB46ilj2PcxV7MEv5TJPaz8GF074G0W29y489hc4c/FxV82
7u9cuOPpvAwAhdLNN+nYnasxKinqxVPYt5uiTMblgi62zwNvceHdNj1jWH4VH4Lh
rsiB2svKoQRLpbLWVDY2AbV/W6Ol7JE8b7HM1lIBlDQZSmkxVdkMmgaA/af7QReV
JsDtmswVEwZw4E1vOH5doCucLio3vv6+6aLveqAN6s4Gp7YNHDFQEz3mljcJtGnU
Ygyc4HdnDaWGfk+vbdbWgVIHdVS89CZzgwdVmc4bmMdNg/q2YWX22tpguc4F1Ibz
1euQ4le30315oOraZwDDuYfKvk5nn7SCHg7lTGBB45P30nrwu7loaacJqsHhckdj
B+GC85ycZ9cxADDuK2pkMRbImwzVEawcbM/No11mf1oyDYH9i09A7kvXMbioV5u2
qmbGLi/LTq8EYC4sb0xYBEZLH1fe3U4WX/3zYi20R4ziOziDsnPeDaB/5qcPKG3Q
v6bKJCGkKuksCem5T+gAjoUCZ0NKQ8aN8Pl01av0+ple8Gkt/UkdxBnep2jQKmeM
uONwJcuqu6G/XA/fFLiNMSyJBZYTnVQDLXWAXJpP5eX5+MKkxWbnafUI/B+3r01B
WJsU0I9jiRes1v8SIGHBQGwHwkeqJ34WOn1pjD15ADcz7adW/Y1J8zi+y5AkXMCo
7fFgS12aH+jGUeOiFakigyjVykOhW9BfA8xAsLvv71o2UbSnHZV14t2rf6eyJ7VM
BY5DRPSAxw0LvXwOg7zN9Dxyo4nQg7JAxD1RQ7xvxT6unHVVG4KusbUMO74Oc0Ez
yJnK+M6BfdpsCFH67pJCygPgYPGi1G9bjFPeWnvlikkXQIRSGb3jgkxygXqhhj+g
fLeMtcdra2SlV/zoReCwD+fsGx5UxK3vnVAnoVAcx/nR5stklyJzyNWT0MwCxOKE
WoojlpjwIa5l7vItVA1ndNwoPwI0ysW6dzgPn+LAweCnKpAXKY+AK2R8GSJmeOkg
SCtFCjIvR3IghGe1LTCoTd+G8g1MBVz+TenSeTG0ZPyjKCgWQVsaLAHGFuMOm3aB
O6PawPYSg0kObV/qsDrowOLGkBrxyxSqH4TimxXox8jjwRq17TZKk3NJvIQLZVkN
PDR8ERTkIjoY6JqpSt+bXtlgY1hmiEAEdzskoe/aWVkMMLTm8O7xqUGW4dvBp9SM
sSabnGCfRhaAuD9D3GUJeF+OzAmXAIwzIrvugexTe0d2Qq+8Zrp6GOounnSVFl7g
ptDtcXOKSZMkEuug8Xtl3pmppJEyxMj0OZIpW044XNNy5QFSOCFIoCS421mVd/Jb
9oHg1rIZyhE7bavwTbY5EhkDQo/3yooi1UmGLMizRuLL7Se8exdsksKLtdyJxAhG
zd4ANzTGcYCQOvGqOVEX5yp0Ci1vLY2wTPSpOJUR189+wjVnDOY8XACbxK0aVcW1
zzMIoGRaMumw+qTnPNjSZLtzoMwG+sxgonyl10NVxUm8RsmIFz7R2WLtdpent+T9
yOhJkGqjyoWfBTfiEjXfQ0amu8y2EhtClq9VxcFmx2K9DhOrb4SvxUi93rEym5lc
vFVbVe3vQH14h0n6h8RjARaFQftwOqSsmuVgGxRyxyguJsaT2qk1onhP1p+7CeRj
efUm8+xVi1z3PkvzBI0H4UHaa/vwooBwL00/RUlOiuaGyAlTwzUDxux4cXz0oX+E
G6ZAVUX/GF3vxeiLMe91Ur3jeD7hOZe8BtOBwY4ZMes6A/csZwvJ9exR+90N5rHW
M78StG6erJu5LDuLq2J0w38gMTpZ++x8D+Vq4nWLiJtwFcgHcHmYmByx8ruUeTut
avsR5kfsLorueaKKeU/rS3HOc8z6mWZom3AOjIvmVqDmKGXYNX38RzTyFnthUT7s
fYQwmzLUelR9sKuQe2AygoQOEjxsd6JoJ9Qov8a0OtUOEFc59mxnOX1ezBlHonse
/s7lLVVA/MHzrmnUsDvBh30UNHkLRNzfWk8PF9/hrs4gz70iiDAOVAiIhswl6oc/
GtDITxJ5eCHcsjRr1A2k7dH3IgwvYilEvA02YA1kUEx3OqTK2rZe7q97Lqwnp1IU
WwkUJwxe5KphMq4vLh44a9KuY+MQA5GfpC2kwxSsSrHED3p7LVvzdQFRQqBwea3u
6VjBfxkRJAEd2rzHOgibfU6w3tetcpWtbDmrwFeBvAQeu+LUMDfAqezyWW1AoFHh
2+AWU0jWFYWbW10bFUGqdYxuRP61VRQON1WKuE0QtLu4R9sur57H8pp1ynVvh8u8
eeosbG4mIa/Jsxi4GLU17YZr/qi9ABbk4GN5dTooMivAnMX3Y4Garzz8FC2zsCwu
UrYkN8EB4+i2PW3tSLGdfLGlif6PWQyn8YS+94X6NxGZn57OYHR5ldI0WnILDbyL
AxH08DXqRubQ43tGzk/OxO9FbGUnnOfDIajwARPHWAnid0qRLdlxgnuN0TV3JpGL
iteC2XBKii0ZhW4uYaW/Cw85oxNAEKl7vu0unbwYbH+sIBO2kHOkC6N8eYLXqLvd
zAdlZG63aS6TwsxaMaK7e7HhlmYO9UHCpSkRRjv6QjZc5HOb8mKHHgFuF3+qWTyb
qQVZEghpfgjSHMwMd5eqO3QEQNvBvFDJ7TQFNMkZNEws9SE8r9x+ZIJIinRKCtp+
4zyWQpDU2YB8qABtzIYzsvTNELM7chQISFpJTah0QbCXJC8la1hC+LhKfRYrAfhQ
kMbSp7HjNidCyyvc9CUicbCGUFJ4uK9jxbsncWw69HNpK6R3kVDJ0acRx2uXhRsc
/TSeVsjPGnTk7QjQlnVvE/oBHI/m7zSLZp4kARTXN/KRUDZ52u5XkgqfAJU8fdlf
vwrbyQI4vyRIvkBNUJS5Y9If3Do8Jf3bXC3Td/ELhgjAPK9yuClzNbmM6LZNcMbi
z005k6OY/QP5WfceQaFuwVj/763z5bajbRzvu4HvwVJG5rK1ImFLsNUGsdm5z/ZN
EdmMIjYQzOVmnx4Rh9e/6AUOC0OKKLlWnmC5jj2O9B57Kfw4r7lEGJ7OlTLdXpvv
Zn0p3ndxujS0tG8skQ0M8juif0kjOgr2RxfBeGy8N4kSugroKEmeh+nPXrwFuH7X
uLrCwyEdhUKQcvU9IiWQUbK70CRh8tySn9dybe+Dm/s4Tq3hm1/fNqSq97V3ihVP
3L09xCzinqJBJYdD1GCN8RJUVZ1m1MffIHYSjtg8GnM6ZqxJAXs+ikbF55Bs1xe/
YRp9CbiRsDXpvpycBdvVp4ppArZIWmlX7sjrMuil99G/LdwfbWex8zlh83jTapLD
Z9Zqg1HlgVcvcACWaYOnxf7KbsB5yV64f8hUNd8fHli6uTfROK1wDFNKNAZgGFFI
Yf5osulWFjo99fXx+xKCLHkzXLe5e2xPQVa9bkmHlhe2XAKv9e1gQE9wV2UcVk0I
U2OysZul0uGtp09YBhH+Rg4G3vGfCN7iQu46AcpqAqZ7f21NX5/blysu0uH+Gqlt
yweMbw7Mww28Q2QNPffQwwZd05enl91+wQ3T0bkIoJB2GUnFlPmzvbBSWDBImvxL
ZmSUEluN96lX2myKjaxTYGuGULr7rLpFxwm0y1t1UIQRFiPbBMih/SdIpDt05OSh
BR/RGbJieExpofjQbYsQvoMfSrUFZSutyqWvgjkktnRQrQVWm24G6wIcPni74kaA
YFsxKTtnE/lX8ayKJIbrYhOnqL8y2Dun1IQjZkde8sAA5k+XLETdMQKN7FuUJBP0
P1yWKN3IP6Gmm48nlvGg9+fNtO5m3axJuf5AWss0ykCLVpWh18OEqsLB/4w+GYbj
HfOMSL+rWAIfrQYU01002fDTiGyCagyPaN3SS1OaNnzZZoN8V6fnZNewXgzEQ6O/
QXE9Tg95Dg63Ag7siQ6t4K0Ll/bp0RR9gmr8i/pNG+xdYTJgXVvX6K3pWQZ0xL3E
UPe/WAvlvqnX0RpB68pxbSFp+nD0I1RtXQtXrKjOse1FGCvBCBOVu5KGv00C0y8D
QHmqYw7Xf/0Hgpd8WUF4Xju4ZDomuO1qZsz+3T2aBl2mlNAYXOIYYC/rNUzR2721
vNsDEByyMf73OFwNgTyfSQDY+yhW9V+bhCHQciyPy8U09pROA/oRexkxSGbMGrNL
Dc65ObGfdneynCDphcAeBcwVSNCUAhOpmekNXCjw1O1XHzJ4tECHWsNfRbY+ZY/l
Pgwm8UIiTct3HrXVnNvhZltYoWj1ukv0W0rzNwp1r+apy8px4fT5ohP83Sq18CX+
k+IhhFS/abAFEnRVU/3sYSzI8al7W8kweLVLhxVatqPj90XantqOCwNOKyI/oeMT
EzDlPgA5WtZgOn8Wg6os3j7620cIq0ja4UkVT6sPMlP2RoX4TX/o4jkc7S8pTEtT
hpEpBJdImSI2oe6gEtm4DrMsg27U9i10Qo4ThSdqOilINFN6pEfBD56SuVWcDqad
ej2GNSne0iq3+dvF9sAR1YsNzmX8uFc1xHKsxtFM+JrSwRCEooKMj/VUsF/Iro6l
kFxaSJD0FBNoetLNK+w/UDvsI0NVwsONdu/ycuCaeuF32uv9c8X6hkAREG2CBDFI
tAli6sD9Qbbx8iSEHDw9Ruz1bJq2IL/KFgL6YsOBkHQMgKAT/4qVlUKsQ+SZXpeS
39ml4GB+6b03nGawmabcO64E8aoIK2Y+wLVZOfavEe9zFCYsWtgSxQWIOZnKAZZB
6P22UAlsXnnt+pFgiYlimeO5xdBJGlQfwAodNMUZXDmD8YVuJXJJ19y8WWVfXtu1
Huc6XiFE0I5cZceMw1YyK2MLUHcxyphI2WwJGNm5V1dsjGbz/kmf3xWOf/FwosIh
uAU7HSlky207v8AfoymqBKrBKFS36ezOCntwYb2YnlC270/0eza/jBNGtFRtZsR6
+4UkmbUNEHi0LCukPIjk7oYPmU4VtNfs/WRJV3jhNBpZpk0z+T/3jJ3YqZLDjvuW
aa18VBgIskMDocXRzzzkT7o2ok5Xcd3XVQ1CCmzXlhmb/+amTmVFuseDgWwsBFOk
fOl4+y7bGTokbXUbvQaaFeO8sEOaYFHBh4rFvi+485TpNwyqL30kGZzI8GHyqt40
CE29LDJZ9Hmys8FjdqShFeHL6LSpALQTU8mYgSr1B/PDwTp1XXNG6ZApz7zXDUDP
gGnRZY1tG7AkfBx2kiGkEdO7sHTNS32T86sGuyidfx3dNBKgaq2mx7qOuOhiugy3
wYxI6lpGen3T+07GnYQFiNZ+uzg7ytr+BiUDsnBM9jaZVqLJJUUk4JtR/YgGb9zK
8BxWCX8Ya0QQqNl3xpZJ/RBW6wU++rEvgFpxuSdEKDv8YW/pHf5FaWqgbH9JdzAS
HeCAG80XHnlEL9z1eHDQcwsNmoTW1RJNn7A4luutQ0dAS6wr+aqwWbojjvRbOEwH
k33MOAtbpkW5U4a2qqfjGsKpNfJPM9A4kUaKS2METHfOZJW1ftuUgkGoB712T3S/
lrUuuCrG+S+PsItUFmIL/Ca5+srzL96piefZ93r9sn2dhEgLYrl4yT8AsaFGiFQZ
u8ErcX6p71LlNhK5yjuWHVmiIUC3wk3TkAuRLa9+IQOkFB+VvqT4KQTSfSNMjyr4
UhsgUvlPe/0ML+70xf6/kVi6aXGtDHeKZawbjNWuglcwmbrVgHXvOPhWgB2yTBLS
RITfJQgy1lGzMbCcVWMtdYG2wZE+YoBF0czt2H9R5PLFVqUg8FRuMTmFEKG3oRWp
fI5efoLHWwEhkBYFwp+LY3oIckFf6ViKWewhrUsot1kYv2pEXIe2Q3ZCEpFrbqly
dW5ihzCEEYULfVV9/V993lLv1Hz11tQccO4tW99dqKqj9azLJ/EfsCEJxIFo5NH9
YvGWKWDPAtWUSUPiolcn8ZhV+bu9qI2OOTMf+eafETqsK2fBXr1W/3d3KpSRWqfP
Mm4XW4IJdT8QlzDKn69dolHz/gvLN7svrbWG3T7DK99u0OluCGOWDkgv7UNnttWe
PtX5WjWr9qBbQ6tE5OSxHatR/o/aMB5cH5lEl5x20ZVb3EkBrdCL3A/y53XhTKex
G0zX/+pmnCYDhV3WF67ElElfiKhYAE3NrGpkUlc71mgkRgKOrhwN2AQTPeVrOM0t
xWO9lQ5+UyUoITbKPDqNVNzXuXdycQ8rvFX7PNVcXWPGiNZ2XULFplyQH4GSIcrt
LPH/Ql6wFm8a08OvgRfTI3ykbrIPXA0fjffVW5Q1aNVx6T/2Dyb6DTi6Kl7IEIx9
uuxmKc6653/uhpy+2W/TgWrTm9MxYidttqsyhonBeKw9qVFY2gmvxWI3d7I5NyWb
P23S8EwEEfM4RsroYZU+I2tEbaWYtIE1vaei9mQkz7L28uoBcytuN+tMiFfFE1o3
QanVkV3/uDxFSRaPR/iFvRFbvkKqec3mbztjigUWjsnljHpwtXhuF6Xm3p33O3Lf
THV4tTVLzTbiiH4MpwHqegDahvfynCJUrJ3lB9/Fmor5tTlJgG0sFJ2pzxXg13n9
hoElwyNcha1oDyuiYrs/phz5u96tXuWWty0IlHgDtFvv8jHvMt5+zziGsb6nAcRN
Kc+C5lRiuLB2IX4uhOVcpZUWKYYbCUxMob3yYgVhsTcU1wZpxACrr3BeN2y9en9N
eBg3jg+XRSbAIaiGKF+MntydteHDVTXkEFPjwCWhWi+P1ju/2AFUZi+W1NjJUS6/
2yRZo+SB8IU62h5Lwn2OhQcKzARQTCCMIm1+LNNJjzDYj8lE9mLlprR1bayMonLJ
Y0F54RWHJIj/7f+V3G/IEkYsmxepfD5wwSGZtNE+ZSG52H6nbASSr1yuKZosIUpD
pq01TrVsdacIWwXemecR0VyUkFvMC/iltdqjjzOhA1FpyojGqjKOR9BtfdXAO3H5
sr2WC7ZyjDZJrJwFfwEoD1kecPeoCYlj0HQWNx01jM4k0yet+UnNLFM8cHmfOzuC
SOUMK3W8jluUbx90oUdTawX9RSFU9r8mUzrPBqUkW0czwamSKdzN6sR9ww/Ww+fZ
EVFzj1wqsfq1FoUO5qs/xKt3erVfs/IJQUdPjFosizsV1GNZbACbljGwhPLUPvtL
Ndw/MrGUhpXjOXfQbcU9qzi0yhT/uooXjs/7WRh1ITayb7hp4hLLjJktUxs6rlLv
1Fyr0qjB0+IKfwUbzfFkPRqFvT9islriBz318pKMHGgGKA+UdbuNizwvSnzGl1gg
0eM4jQDBrPy2vorzJvfCxkgbittDrYuIPomSXzUHyVajHDOoLsnlwpfCWbLF6knD
9jzzpRSXlIBndGMriWPC0RspunECNg6Zo6xXhr4bRLmVMljuZmDyAD9ZxYqKYSzw
RE3eX5WE31pZda7c8lAc9EPiPX9vgWoaczI9HVWmJwjA4zUTi6vheRXvqs5NLS47
8RPlhehV08ryqh2PqWikZrlft63ZWdyRU549LGfFky4YDsjboqBdFUBwmV38ZzM6
2uCTl/BWmnNjX4LWjZWaf65eKo37XO5hoYVAXdMqQB8NVq/7zfEZa31mNbn8wUhF
rMElb886heMw/moig0li8myKD6Q09F23l9ssCDHhJDUxtKEIroICMhGd3W000EZ6
eFaCBj3BLiFcHds0S24rwsHpelDE7/VgxMWAfsqAx8qEm7nK0LMSo/Hg7LHER3U5
7uyl73WOa++0luCcp3Q3KIkYURuYTZ+6ZkkoDxv6EdPvopht3Gctd4cXtL7mEp2d
WwClGWCM4zm3QMy1UnhE+qLe3Vx5n971qbg8UxzUhgH9/+sxjznqFXhWRctTQUmD
vuCwhN3vXgFxrPgUgxuHlpo0Lpx4ZX8GvHnNxsoXTWlQrLZ4VDDcps9kV7MYE8fz
yWsKLNdmyWeTpfxIn3ntsfdpyUqyLdcK3pYClQkOqOEZxxgIIt/n5LLG86k4VnlJ
hv6MBprY8zvgzwfAFC6Ut8ZDNIvfUxvicNRl1gozVrNWuudn7nakMuQK7Pm70HgR
ifvEJNdMyJrfgLsykgz0eEWzHgrrWoeUdz9n+H/GCgR7Oiqpd9RQPEEkYiYT5dSE
x6mNmedMoiTTjqQAArRLd1uIRNva7VxngviYiJfcUb/4XYqR6wPL+XTgb+7IZWfx
9bSddcGg4eORG6VYS4ZVnRHPxJooBaZMwQV2s/mGsN2xujSs+MdZO4Dub8kSIsAD
7EvHuXXg+5WDqvbBEVc3OdWlU0v1lNjAMoLtqMW4JxDToWG6vk4UnBLPdT8pnDrD
ud7S3+L6iSpyLBjKUctpG9OKJZ259KjBAry4V6N0dyh1bWIsa1EL68kiYSMgNl/e
P3Vr7veV3m3i0nsOwKsmVADucp/XSh+6675DuljHEidf485/qj0voug51LKXnczR
QXQgLCpZKVbV7SDdb5Q729HAAHE5h6irPsKsGodO6P2NqMTGhMZFPdSp4VZJtKS9
+r6ea/LLa5YQtI9B7JRMfZq2lEVICsNwWkNhTpED2L1iZjcRXJWWQ6guDVE7df1v
UpJummUMerrElvG3iX65DEc/eOoGO63sjVuDFK4nTcNwszD2I+7E8h/kMN99o3k9
JxOe9oawjmL89Pf4hvdwKMxZ3IQo/f7GKBmnbpw5VzpIaAHchOkkT1i3aowSAu2y
5wKdVbIp+RmteXQ4iIbR2nBlfyFaCgnvkrayeF3Xm/DO/93IfXWUw78fbgz5LCy+
ZmDUX/W9S1IVrODyVkcfOZeeYZgOzhQOPW7YJP9JiUxiucOSJCJuVT1mECrbTs14
ikmoYkznuxQlEZXm1kuDTTBpZzOg+3Of/lL3cyrXTidT0p4gcRFs2MSlvXv74ny9
vWBB0e8AEkP5vTauAZQMAZXzuqX3jtVC5H8E+wctzXP3PiLdlBI8uB+mulKub2dz
Nd/k7M39zRDKcOWqsK1eEDMGhSOXrIPhjxxkRoC0W/gmlhGr9T/T/cH49MPpwD/k
DqM7VsMhxN4VzQcMROzoE86DpkYAMb3/UVD7QoMAOXqM1gVOelaHDH19g0lo3rX/
lPMZarjL+jFfNb1TlvHQC/HE+IcYWVq88fOWTDCEUrH9uh8NrvC723aRjzhAk1hm
vCdmms0YjogbeakcJA0qEwMHZDJ7q0qIgJ39BUHo0rPl2wcSE+UScZf7R6AlcGYD
DXDzMYoppYUphw9azM5Mh/N6ro0vvN5O3XUBNAalsQqhfcyp4xhvNKNVTXfMM3Na
IM88xdqePSZxQ8ThmXQWXjEzPetdAIaW/VNWd4DrVZ3f21CargxI2eVrydv9O0qk
IJFnvhSwk/0eZ3TOmFyIwFZ8r1EVHNpznQ0hXhhgVL21xsDz2aYmsnvHZ8LRmv0V
r8XtY9vI2NckJpBARDfBHr08f/SdAQsBWKNmJD7IrTtGRWkg7vWp0Hfunl/8UT7u
BENKkwflyKNAmRqN/0VecH+8PB21+OUW4GHH47WWLOG5U4EtcsCaNbBL88u81Yjh
4rkq37LeTQl5LV7vxFDABnnqDZQEuDJm5rgm3kudi1brCykHAgXUc/Ri0LqarAMM
WJaVxXdSGSskPOy0c6AkHZh510n6/ugP1hvHxO3nJQ9HY1yw5KLureHyQQMYr7j/
+C2n/jkOgDmvwqJn+imGwuBBrJC1T91JlwsLBQmKZKUnwIh0DjxleifXnXwTsZOF
fQPUhEMq9E42R2teALIxT3oVMSwcxvdxSTcGqNng22/D3OFUqljXdggWEB2E7+Lp
lkeq039J222BTgdQiF5o7RBkIcccA8RljeFPfUt3MjwMYN05xCIcv+9n/+Hkulrz
mjsPWLH4pKcKfa5pCmJQJlkv46fpLalzy4aYmzsaMukhLkJJ4xTrLO2L7JrE573D
s4vqwuJuHGCebwyoW/Z4aDE2FwXUyFPCl7GSUzIvCJCA856IJmcoiJ+2fPlj5Km0
P379adDlsk1xoKR6iYISOe4FZ/0C94NIyUP9gx1ERm7IzGxuCjVkCmqSEG2la3Te
eX/IUqNbVWQSTBO3idJ50Q6yZCBM1Q/n5xuYnDsgbHHqTgXCPBOoS3+YQ2IrfUeh
Pc49qUUjsVEuXcBpZ8AmY9zQbf0baTg4IHCKRDa6ouNtjMJIKeQD/Mk+p2trxsvb
sZROii6p/qs/pM7N/uF+xof1sUYmtbgYATsKK6IxO5wQTD/46CxphcfCzHiPLRYN
rQlTddarLKTq/y2ory995kMGE+Ft6wy5AobIugdJBx11QodTqBewAOnCVSN2OXcH
OCqPK+FQ2fSsKj/8iljfbizTJ+nRQuLhYEkSKk9hUezoaHSujLrLkS6fPumaRXRj
QTjPOj3jSRzNGVjK/2EpsnQ+G7NtwjcHCPMyuhYGqWl5t0vfV/BJ4aFxlpHSKTBU
KTEOg8s+z0CLyDQinTITomsy6CVwFPy72COakQmbzCb+puCgJ+hVN1Z1Vaq+80vU
IgMINMSXMJ66aMHmYeCbQsriQ/nQodA8H8VtXZyoKo766Mw6nF9hm6Egt/xZxI8M
8SQTPAlbWGxnIY90GuS6ZgJrkpRDSxU/y/B4Dx9iaOWC6/knlxD5Lo1nO+865Q12
Oiul55HdgRtpPkFV4T75+EoTr4fj5Wm1YvJXxiR4XnmfnDnnP6MWR/xxEIYlwltn
Jba3ZooJcx231YP75MHsBfwCCkKg4GxTC5+EFYpUDqe8DR83+qCveqYQmkSEyeYV
WjOp8Y2jFvng6tld5W38wT9jx3torE/Y+ApBf8h5uV8WsUR3JVMb6bQyyLBzJEm9
ve7AgcXqD31L/Tay5xlSAoZjoAcIyI52g98s4FPX4YSJ5oC8xr9r+tQllYYXqiVO
drXdk8ZXlf0IwMxx58GCgSkVAzgs5JvIAaPojITgdMrEfKob92mX34KGmDU4edyk
JUm47Ukk1x9jkCKi6hyi90od5s/ur0JOh0J3KTxTaseGwyhM/T2Xy9GvKyrZO8sB
GEuda7H3ktETbqVeGJa293tx5PRQGXhp0czLQnxR+oNHTHKIXJhM/B3Tp7DvxOpv
9ummFZox0WB0SvWQsOrpGbjzw0QbFVpc3BHeOYI0bvWSwDA0fThedhPOYECbsCjd
FGaE0CkbK45Cc1vIlGnhJPGVOE6OqFl4zq1s3rQFWrBJyvdjy5DcApRZnRID7qa9
goIaWIJHeYW4ko+7Ak+8pgIc4FBzhZFykbmhWAjokv11pjfg19DJHhMpcRHNntW4
OhYGluPO1JFSlcasDCp9vvfyJCTepc1F9YBjBYRSGBhIQPGNGN4gz6cLX9Z90ReW
9F+SM1lJl9/43jkNMO3H9o9AX4CyL5WNhzK2mZNE6fI4GKjJ/gKfyJQSbKTPFm2g
jQEFajdTl8K/cAGdlIyUO1nr0gxQAjHdQWlofWGaltyGshy3ZRUdJm9P5QyEC82V
o7TXQyN6lKspFSgR4MFTccd2V1TWiGa8mtzSnya7pCSuc90vUtD8K2RRob93hwhZ
qFJ3VWTXyZgdj7YZ3rcJ63sB7J1/UscP5s+bVby38dCo//ZlHw5JAZA4VVqx9EAC
gORpWojewga0qPg6lvX+XsuqXSAChGSbXpBluA/4squAmG6/pbSv3SaSQPR7a51R
YRbaukjKrMFjk9PTNEJDMcSHR0FG5r9u3f/RFbYgkDE6l75TYaXzON7O8Cdm5css
QATNOQORr1/K8eDHwX+Oj76qNqoiM4Tsw6fbuzEV9ICRwkpchBafHQesLGQHclDH
MBWzfZGWYIABCWk60eRKIypkT9Sr6WkZ1ugcorMcSPLu+hKlGJwx3KDij/K8y+E6
26qQgLrz5cQmyIGiCy+RujiVO5TIc2ydB1t42/45cJg6fC1qNYl9PDel55HTJrgV
ZdWTSJ4DfT50Hl64hKtS/OUr83TXXs06Mk+2PXvtDww8LpQlj3LokBgqJNvlM9YZ
kYBhHY2Y5OBwHnPuGyKxR+Dp5vuizYAAIX9maPGvh22DjjWgdcdhuQ7QW0qQy6+f
nsFsyJVJaDZNetV8YPToUbkqEEpWRLfWnT2h2F2tnEWMjD+tYrxtBgGn9SRDA6wI
z2wZ9GEzLI89G6ofcFpKPGKlysBknsKDeIMRxgH7I5Edgve8xhFSFmTkzTCn5/LC
OGj3wn7FohQ/zRj4GyzwOX2vH5qCfIWRxSzwgyJ/zGph7Gh1kTOJsBRlX8pfr7gq
xzpyE3dXdjP7U9IHxdCBJJ32O6rzw8JGje679Y7Vi969rMiqCNjfRDbSSFCCAEAq
zefoRI+wZChs1VAT5i5u3mj9ZgxTQccTPeDuTSHVJfuGhPFu56th+ySeAQKXUxNz
3eMKKr33+nMo9JLQgWAHyjSWq/RoQ8RzQGpi8ee0D9WM3b8dMr/xUC3MG87eAXrR
C9LzIt/5QRhC0UXPQxmqj7mWM9r3WEoCLjfp87JOREAysaUyfsW46jZISRyXqJB3
AZ7ZZgV03ixbd9lVXuHW1kLH9aiNGLGedeL/YsXGfzKMI1BiZHPUs8ENDGaLqZg/
K2TUudTeIIbdKHkEa3s4u40nxedvhBQOz5Ak29qAkqufy0wjxsidanM/Z5NdePnc
AC+fmRS1QtpGgxwlckMA8W+AW6lhWBNa+LlSAnCEyN2NOF1FPLnTP2J12F1a7rsX
/VJ1ZfUu66H/pxoc8jyW5lSywW4x04XJBDievEvYIFB5QhrQx8K+PGDQKnNbVxIl
ntFBHGuzP2LjKwqQ9i2tTOoZk3/gST/d2C7avavOtojUWwnsIdQB2aBNWfrHjbV1
we181jqofhy/WmLujGREiGuTdsGEDClB1LizdZTkFSudXF6Y2LQtcGaPbv1q3a72
IoU0hHbRJ1RQy6qwzVpn1vcwVzOrHPS+EHbYatJ6E7U1araKdJLJRl1nQ6NaWZmD
a3pOOOPaA9MrY9f5+8qZ29d/wuzYTBcGqm0giTWxJX9YfgqZr4cfhMcZqNtAnUSd
U29XaLMcs5+ylMPFjZpifviPxyH5oONPPYWbNJVY+s4yXZlnyCjtptbUmYnpe4hY
Vo0MM0TN/4hbDk6Rk3oFiBSEsVwvLTJqe9y3busiHi7tTLbCf3eoS3s5rgRiidP2
ZNvewylmH7/1muJ63HMTD21SuTvWCqRAgtZyDCnLU46+B8FLKiifLYln1jD4Cj5V
PJ3Sx/z0ilRtegP6Jl/o4BkoEpCrto6w93p7u80bxzh9DnP5yqJiKL5ajZCYfZoK
dpVJt8gszfKcZM46h/GYocnbxGM5vJlI2B80nshXes+/3n+DUtpUkQQYA93f6Tif
wstENqHYqu050hyLid9fvL6Fyjcjk5zLlaDWlMJkmsm9XzO2x/b5j5ZXDAMmrxGF
Yb3ehCF0UKNRcm5rAqIyu4fUBonzSuwUAHkyyarm6nih6VmQCZcooXHQubMP1dxL
5bAlnKQc0/f85D1FowweTLfultn6DMtAeuUfWb6noyaiz8yKw1uZ6ZBONgxi9EEH
vUjgthJH8Rc5DPGcKW1Nh7ProOgWvm2Z5RZT8KnI+2wyLlaJap/ctKflGFMaij5m
EkGSWJ+v0ne7kNUWMYEQ/JkbEK7EULL9D1XwziJe6OeyOleprwEitiYZovnAGMyt
CBC2OEwvCjywyz4g7pTDJEPCD1ujkNa/jK9GVhJK07AyyGvHC9OfRXK7TiLLs8MK
cnVfG80ypqmKV6HmEKiLqrTXUsmUhZ0wavu1fXEKE1uDsWJibmOx82bv5Qi36SUU
6WQO78OrCO9F98wh02QNwc9/v6snd50m6cwoWqnwrfcZVt9VBDbnVMmgNX0trEuw
hrAct7AJg9e+bJQW1O1pViRsax0NeuFipGooWpH57A/v5oV/cyqZbptP9wBrmwPX
pFqlgnVsqWB0pMZIWShZO7ZPD1IBocBfi98BK5k5KpL3GVARV8xWNVLxglnTk1zU
VWh9SrbTIsjn37sLuFWMaJfoUPZ4qA2KyNza+I+bldV5ABPfWdmdt/ShsHR75sxG
n+z4JvZ2lHWF032/cBt/v7wdNnJPGjZ0soY00cjpf//pvNlWV77TrI4pkIgQ24LF
s/7QGL4k3pU1HWYf/cEqcSGoFrHvoAVKOwPoPWbx/JVv2WsO+eFn+j/5yP1lIebp
OFm10Fv3S96gXEtiItIbu+NLk0c4gca9qst1MsIj5HPLICi3d3+SF8VkgG+tgK0x
iYxwcxNt43B0Ty38SSsqThqiKd6DK498ygaw60OXBuS4fO2qXpoEkxheHBRKJd+6
1z0t9upArP12y5ZG2VMRB32Ctd37Vvg4Pkal2QJ9Sun3TPGiyO5vQ9lE/PKCtcn9
IkdrVSH8r9ypbjasx9zOTswv+S28C3DOM69VHvWf8E8ujHu1rnuPW4c3EF5/ZS7Y
NzjVRYPcXuMighda8P3H4uThUpuvlOBHdt8GKkUxhbz5Irq77nljaGgGyld7rFQE
5rXQR/+nGpugHA+zeuXIEFhi1DBgOWEgjs5A0M+rAYIn6xAE3RS+WhhLZVaNtpRl
lnMnT/MKX8eFS4I7grKyk7sbU+21ici8JdKDxe5L7hA8g7ycWeo300eX985+adFI
SJIqohygC0v7Q5DVVz5aAIg2Z++NyEK05wkpbNiLfKDzIIKwB81yqlum4zAMao9N
2TMXSM7JRkLCyJ1Vr3DwRXUGF8mroNFjDOf/8uBkW79RwIpb7oQrRU2IecsVnFja
XE6hAgvo3grgoDoXioEDxlAOHhFgLTwDv+RoVeXRm3Xhe4YBOzDYzgWV8tQAAJ7g
IvBr7tBue5eEQBP8saFBGFSdwxpryAz2yHb+zS3Ln2cUBlnWtW9vjkoT7IBKflqT
qVDqzEBMYXtnEGKTCDQi+chS+L+R1XTjCVI2bTVXQFdgO47ZphMvsaT+OD6fvujP
xrQ8M1JhU5yBG3R55twYx/VvHV87zzyCISxDz4klp1WUrBsVr6JtZaCEyIKAzi/m
juYfQV3J2FX9WXGbR6/d6DY2UkhDCb0AQI1uQIoEFMN3spldydxXC6c97lwb9fC3
R0R95kFsiRogDBgHxWMG9fpMaWnziF/UwqlXOhXWKTSQ17rK4t6y6hXIlYy3ctlj
KsmSsuGhlah1Vyn1+fD8zl7WOUSBLETLNkMHMYXgE/MK+OSuAfSa5BM5DV1mP9b6
rDfhK7dTSJ8CoHOYP4nWmsyzzqmc5z7+S7wuSVhg9g4Bdy8i3/WRBb4uEXK0/JXO
p5LWfAI+T1/bf23LFBMHu191rNKNqAUdhy6lSyGbZOZOGJ+AJ96o8PRin4nNqYjM
n5nNcKx+cxAeRjOXlxYhZ1icHs3h+EwIes8X55RH/6VAPg2Sit7cOxL8xk3tjK+6
zIp3nkFbdpQVExbh9Itbhd+PuC6bJSPu4mw0W15Ze06Q4YoA4RQmhddIeyIRrz07
591cdkFxpWLCqn579LqIpai7id4OguLOQMWXymjIBvghECE55jaRfSaRFilcJ+xZ
cgg0mbno1Q0Qedk6AfDYDgU16qRVFbchGv1qX/Vld/msgS/7y1Kux5e/CAB3NXwn
ArvzUbBi8ZtI401a3oJiNKkk0ujsWDqCZD6PcTQ3sgoA3S53fLu/nXG2xIuBALo1
uDauWram2zU+MTNL0otyPoSnaMH5iOde0BNs1fnYnz9X45w7Pg4nTFOONY9mFxPY
TxibXHvIPsGxIkUHYF6vVIXYiBOuh9aAYndLVFIx5cLgQyg7tRhDQ4lC4q6OcPHM
JTGqxM/odJYylby9v9/0LQznRTwgKYj5UOj/HESwsxuFKKExhsUbHBcal6hatl/G
krc50WH1TpT6zPNytLA4IEoVcLoGsUKRQq6O6+rE8oH37qDlbCCMkBDUGUQ102sZ
RWiseIdEToguu0SCwT1RZ1gHcNIosYw5iJQpX0TrY5o4PNPT3+rVr+6/gDUB844q
g9064Qa53yYx9V1YFe5tEnWPbIlp4N3C/0JqMcEM4EmEPxDQ8/ASTBKjPvq7Fhjl
OtZWhrK8LQy8Ioq9tPD5C+yxRcXoxx/kv1BXjJrQoptIgf4qAezeMRaC4NVCbet9
fSzDeUPsFPkSJ3kuTjGQv+eKHe9cF2dz06nGyLZtrhs9NbBStroLQZ+pHfeHe4Fe
TyZtC26/FsNNBD2KOaJ8VhefrlrzV8e2wcOKkLXd1o3szuk5ep8j8bxlv4UMDECn
SVSgtFvcciWCxNaJC9Fd2nE0W6BuZWNmlGiL7jHjhnTVAFPiZpq8ZwhC8BstXLzO
UT7ke/Bs4j5pd4vLuJVYv7ma/2zvcXUpVs1d3UzQjX6yLeA/b90Q5atXgojRnwSS
3CE9UkyDXdSX8DJbrQIvQPSklK8XiriTYh4TL6oRbTDRw8x4Q1S/dUjTX/QZNf6e
PnxRhPh8Bl/B8RPpK+DR6lJ8vP2Yn+kT64qyYTWsl24+0qlSRvboizDmPHy+xR4E
bpcRbr4DyQYvJQmCyAnFbbDsM1DdmxW/wrwYEAqDSViHEwpCdJiWadr8IJ93Bq4B
7f8ZQ2c0t2hEKpXwp01oVzTzLNpDTIjWyoDfqMGVjATf0r3oCbd/STwKXoCJt5M+
bzGUaaShZd5fCuKOOM66hwr12c1HXv3vhZbY1h8traqGu6bEa1udoI8UofrQzKWg
ghPHXPQhsfhHVF3DLyP1qmfoXvxaTLY+dYz/0In1t/Jou19AdNTnKTOvrKqhYATo
IjvrJH/1X9FVhQk5AMAMJS4l5f0Tpa7JZTr1lpprOSJVcI/GjwbDkgHpgYCqrS+Y
pelusMHIHy9wUsZOKsCGmhOnuGnJz+IVxvLOO9mzWK6a5YytswJPAmnCij9Httkf
2nCAY0J6VtH8qNp9IP1jUsawuK3Dt5sVH7FJTvx3fBsQEK/9hGgYG8SipUaEAQnm
rkq+wzMrwkRwrHbG/KOcmrq6ILj4RouCxjLPVHt1PeoTcHSffdTYXCSx2xXcdIuG
+00+JgCEZiTvPirOOSWUNX+24XA/Tc7Z8c8apxlaefE66IrFfKMbal16dMNfcTWV
jxkiUA8oo7mrC9367vcC6g3Dpbm4SuFk7xaPxKcg6MBrIRjSYFPvCKLxSnrkEqYr
Yws6hZS2NvPpR0GD+YnYI//bfakNUD67UNC41dkK1OXIuhd9QbpJvX49S7tJYNMk
gW1RgltvLrmpIs0PLSdv78oAREd8PnlCshmCbmqembN4aSBdAtRIpxaZviPpnhjI
T3fA/fi2krtBEz+0Qv1KlBfBAVq9Hg0q60zDk/JTPW3SCFqcJ7CPkGFejTQ0vZQ3
+UUVuIJibXN12tJVRhi7wrKCx4cGxwcmHrcsYaUUlb39u7xVy3qsy7qzyW3c/Z/v
EJYkQ7oSvn7vkcH/uWX/QPjyM9dlbC8YWhxbnXompv6C35gUSKuyNvs2Wxy0ScIr
Lg2vhQYk8ZAWpbV9xL+LZI2HGevhobkdeooi2/Xmo89ALC3A7ULfKrC34t/4HY9I
tNINZv4bWrqxjvChqsZ+3eNJwtSj08/N982Oud0g3o3Sytxw8/sXjH9Zj6yrgAh5
2GUedxhDQWSysF/mUCRaL7xIochDi57+fvnoUok/SW0Ysvc3YHUP6kMz6vV1dPE8
DO4ldsDVRcnDUKPv3erY5zTTmlOmqugm4E99UZvJzkjdD8gM5pgKGG4zQrQJIuK3
0+I5KISKK2NYuA2PKEGOfNi+FtuuCoOuZue57xexmTiCyuZFlZk4WLS9hy5FUIJs
3Q8m6G00gFvmObfh5wETDzqNFdrf4ETXzq7Pvn4VrIFPKAqaoO1Z1v/BrNWbqaDs
dW1h0k0mPjxACcC9ALa/m5eiZQYHi9H5jjxZY2II3appz14YE4vN70+HT7VK1VO1
he2JgJJnbdyW3hSGSTZvgOSASU4xPxSO8VJV6t+VcUSlkwwINofoWMSHxfs0zOu7
4Lu+K3KR8eUz/A+8/VZhQQFa+pVU3bMhv5lvZBxg8D91ZMW5/E19Fhnw4ucFl2Db
AV5mxiWDu+z1HnHGvFYb3PEfbK4D98+XdpLuT9LExLxmd0UpQzjwTVkuDXNIGpxb
kaOXV4WvhuMBQbxBa9VpSItvRyjGqBZ1Ey+nSMzIa1L+z+Bznsgkq0XnJpU+7JaM
D8ztg0o6ydbwv4JOcsZztFrQ2jk3RSZd7GNo7kB+QNffBPULtterIHpTr/aK9+Rl
NFQYyV/TohywF5szXgygq9Dvww+pzFzNPK3P5GCL+6EcVJ8hT7N8lq9Rv57JPMa/
AFahVYjkq56SLi+yeMN5UAxUA8E80YdS0A3g9pNrxq+JmFboJAo5tNfsKEYD4RJZ
UC3AQ5qnjhy1Og+5mAmd3uSyT94iQtsoXfcR56llFa888hFXsLWcoYOJ/nC22uye
gdO27vtWqVeYGbIV2jOk+mdYaH+WqAu4fNupmB0TkciSspuDB+MmgwGg/eEh/Dbu
6KrQX3E9ZwOyBjr4Jx3PCZw8bNGCnPm3O38WKY7rSPZj5r4bQ+0wyB5c2dO3wxUl
PpNvYpIybNMEXvuNoxtcHofIgJAy72Ajigd/PMmk9/1+O8v2MJkDLQhC53/zYb44
xp4BEN4dYglO/U5m+xofVTF4PS23R4MfPA2gcBIaLdOFwERigwfBuZEvFf/YiRlx
cm/lohry3mCk+oTAp1q3wXTFMLqpYpj0HHIJWvO4gjVJpoWq5JzUkEcYGx8ByJyi
zYQ8guITo9XY9/TnwAvJzuyIRPSGfSsaSiJsHz4apdneg612Fsvykq4uiDdusBSC
ld/F4JJlJfQLwmBTwQMRvZvJzdvZwsqy2p0fJXWRg/ux8VE+cA0CNJr0bm0LPTuq
6A9t8qPgBza+1JIgKrfjZkRPpy9dPITW4XCjxYCCn+wP67MT+vMxN6yQSTdAti4l
RlCwaCFHRLhtMpMaFnE0LZCOIfDNagFmcN577PdBKC1DcCYxji/0ekq0SmoOMztj
8xodsSt2GGK2V4HY5oJ9JzHehSwu5kAavF/Nw70Ke4GTMrnzkMhmo2Q1vf6u7pjo
8mi7Jhtag01xaxOOyPOfE6GYg2IoTcse7SGoAMNvJgiwXCfcHvNKEVHY48J3YDQR
A34w1s0Mmv5lBRBgqUQ2DGXfrsrvk6kysDYclPLClCMgxe6Y9r1RYl9ClHqqm+1A
vOlWE6sg8r2feTDv9g53KTvpftSCq5HmCAMdLLRiVmsoceLlW2j8p847pzXz80s9
rejKYXHB172c+WFuQo+tfqj9LyQ53porDkR8cr1Zj4SCZBe/dfn1VVqJfmkb48ol
VegIjGBHvqCkIest5QnL5kkbWqX+ItDbcw6XxVOHRITnjkSOyvri9L2strK1yMk7
YhuwMlah3fK5IdVv7lcnWkRwAT2MxWNqBnYaSukPxX3obMRRNSKedBmflCLwaA1Q
66pjGzD0LLo8WM4MTWyFklHGrtl6wpA8fQU/P6x0kL1j/oDKnet7w8aVMqA3ksR7
KdbM64P9E5r0mNlEH3jRph4/yHO0bCxtzbtwvwBY242UT45Af3WbrPBW0dQyORkh
hhZa8UynUdNAuYPTioTLgSy5thRTx2s1Pvl95aa/I3iLZhtRbrw1cMRJ1NUcK6w6
uWiKaUt9Es2M/qHrWaWSjbQaHhsZH2R9OHTIY1Sgi1XpVGJUbABs5/HAxSxLCuRe
v1QgRl6MYVFAGG+qF9Eva+10SiGg8Poq5wCR4B0hd7Ekzz7LL9Ld2BTQVa7wuY2k
0VU7bxkShdK0EaJXT1hlLYv+YLH7OhmBlJ82g8MtTqljxMU70HOCBrnPI96kegv2
YGW1MyX3l1khn+SvbqNJ4yrhYvyvt6DWFomp1qkUbKyTUzNT5jJ/CYktaIGVtuJf
Ze0cuW+wkiBh92xwzQe4eCtOF8YINWFoaCq903ZpaX46bdV0fwqXnmxsO7ZQUZDz
lbhbtxugL1NYcsfskdl1GxuSGPY+tUE8746PteRfU4OnKP32kuoyWHaxFdz+K9ST
qeMB+s2LSp2H8DLHWH/jXR14KUb9bZMkGUsQ3fLmBpCbItcoOXfNm5YsYPz1m+a2
iAUfB70Jp1BROQmGCO0Ts+mcjDiymWljCtOAN7i5kZDTbragHljP50naTwkLdrFH
YO9L0fHtvbrlRWNd2zq4frNX1ObSNAOna6Sjy/YSE9eyye7B4HGkmYfQAbH5ZQzd
um/O0HvpXbL1kfx8BT+1lu6KcvG+kLF8dy5VH+34DgePTPDIP+em8YRN39byw5QH
9DffFmVfFkqPaNb8OC9xskmDp0HjQu1z1E8Ylq6ExZHLEE1EOj+Amb/SpfJi0kgA
aSwL4wbO3kCFWMw2rI4IRghv41XKPLPCaKGE+FXGjoCOKVfLKk05HEEDDB9Nh+kK
BDMZXAZPIXGKA9WVv40aCdgx9JRlr1IzT5AR3q5R4jPRRlGAg+ALEvCZCXx499pO
LXLAFIdtQ6x0TtTxDVoPj4FhphFUIjYYm+8yV8luuAT0tNnaqv/xD1f1oPE7OmjH
WWz7x2u7CDlYyuVJVffjyOuO5ruQQS2y+MCErxMFhOE+C+oaVTiKQ6R4QycbmLfD
X/M58qg+G09AFNnWYFmXQXJaQGitGqOP3RLWR307rgkj1pgR03xZcfF718cFnMR8
zmpXeeLNvTzyc0S+udOK5IDjKG3zXLa581kE4DgZcN5e3AnPrwps1I4dAzQ3KoJz
lRsz/oyGcWg9wwBLaoZEbC7RdRLFzWnZnYYJnApRTUhNdFNnLhQuX3yD9esVOfQU
admLfv/8G2yjCtMty2TCu8L0NQuR0D4EJHOmntcFEYoviHmwzSgUL/btcCSbH8gX
cyDUUkGlx1MMT3rwFkY8ESvfMbhTT+DgviDmHO7mFLLkSxarrE14L++gPtwUa4CS
CnNeR+e9jWNg6yrpbJ0Rbn832fftthc9xE5hoZyq1ei151Cos8G8BIhUvKuDWYz+
V4AtSvh4c2dDewOkmuQHZiq5ljzGewq2l9yoN/R4HFaMEpgzdJYWUoSaRkhtuxvj
A3djf4hNGRt2aNAAqNTOKhVjsw61nF5tX9SwT+LW606u1jh0QCTMnswrHk2gHd6M
ryzJLB2sL/hhHkBfO7S1p0fuTd96/pXiEFkForrMELn5LCE5JZ68hN965pXGRqYm
oLFptDGWF3h7Mwhr40fuNW12D/ZwLFkJSWOgewRgX/2YzpgVwqDs5lCHRMay829D
S6XikkRLP835ltRddnfB1CDTegYqJx4l3lK6+vPtrTlc79FKqLUD3pVeXqUa+OVU
IGLDzEvI0r9224d9+Nm1zMndolIZz9wtyCaHu80nzsNsXB3XpHxih00yFh7EYzz9
1K2wuEEpfB+Jo0WYyOz089jAj2kvxJJtMJ+DUz6bhE4oTCXLtaF7yG/eJYms/pgg
zG1x6rIijye/vSL8WHpBI+uU+KiUEmzVTFH9LHfma5utAJspgQJacxSqCCSSpTKS
pFO/X/pbGD6tQaKojQONwtccmKNwnkeEVcymsmyOeE1rbj10Xuoj1vTrEU3+M35R
4piX+RCNfdyjYa/iVb41fXLqH/oiWOY6ZbjrLzWNh/LMoBf5uTKM7hIs/TUshX3V
EjBT7TJ4czJ0GAMY0+ReTvWN+c9vLgui0JP//8hwMrpT7hpnphHJkvoRnSgxR+Dc
8d5JtMe27Qo4RU84m9I2C/D1mQWZzX1KZWL9SS66XEMv9thQhvliJwnarjP1s+I9
jlIHhXHymFrydXndT4CRJ0nvok5sXBoRK8asPv+IXIIq6aQ5mOtIpsM+Adaiezox
3Yj7v1gy/ZhZpbr38NJ3UXvu3UdThSpYq/6L8C8KowrbUvGSl9uevYDREVOeBZ10
Z9V0sNFMSOCsaAM5SmNXaqUhcD0Mvc3SXLpVZFSb3Nsx3gvKamDVBIP0qMXOqNT8
JGXCHlUKln7zsxvSswCCs8qMLIL4WvXlHjlYRD340xs9p2ZBS1x/lgJO9wkblnjP
K0Qz0b7fbBwSmrA126Wxy/FjeK0R8njIA6gMtQbYQZggU9zFh8uxCGlN2IJeAVlb
ssUBrI+hL7+LQspyWUUd1CJy3EKDzafXljQr9chpjJO65DkTPUAB3kU445ZQcIhZ
PlfY4u6usYXEli5L0TgXtqGNBDOZ7it4ILMx7BzMbBnFIWj5qs0AvRkIPOlyRSRP
pKIbWdiuH6XkQBZubI+tJ8WvBv4MxGe8dfzqCqZJJI9912hkrWVBHxQ7fXtvZtBh
oOr1gC0dQA0/1TYiVQL54wtvSLMAONcKsM+ibzviNc8oMlz9gmFnhript2B6pUM/
Pci6y5hY/JwtPcee/ui1IFRawuV69G4IR898swEhy31xZfgYpNvrcjmVzFJbi/87
lO3GAMI3ljvIG3d5Jk00K5H/+ef0TfnRdtV3zSScTtk//WRahaj2UhqX/+mhtNuk
qijFuxGNtt+Tr7F1OMd8rleMyBuZNRWm+LHJLBHQU2a7Tdjrdg/lioOtGAkNpY75
OUF2T8KrWMKVKebymaSi87UqBv6aIctjOXoU7JevnsdL+HeY7xcX0CEOMLovsbCY
kc2NXVAcFOPd2n2/ij/Us6+7MQidvXGuEiHpY37R6ThBLQgf+Uus2kTKeuslG05A
ScTi1+sRFY5l3dfm/HtLIOCs98whdbV5l0kGccgL8EEp3LgRHlTjVDwNmi+4uvYV
7fp7jQjYmk7TJdbukpDF24Qh8k7mNSLX89vx6dCp/9hbzYYvYDjtapl6jPn0NE92
rnuoTRdI4J2gtytD+D5qu9HlXb1XwVVtVVeNm3AxsCOg6t/a9gHCQEYAJ63c5EOO
1VnoAezQbvsKQ5AjCf1xfw2AX+CZe4PE8Gqz0k2b2nE+pPvun6gEQMP9aJzqvpVm
1xsEt0Yoo1jmfRDyXLmsCKhqDvUaNdNZ8EAU+EAm2/oX3dhEU1oA+uWSRXGk1Kk6
ZXcsKKifHZ29DChpMfrC2nqMdBC3EPTyg0h/2Lgf9GpO9QpfGlwTC3DbjMareoam
buZdce5CmmadUhJz6IJEx+kpO+UdJ9xpp51M7xoJCc14je6XPtHfS7vZgm6e5KZ9
zkCPM6v4OuFRHuaoH7RAfhnaN8LWG+b2sLcz/dLmdoR4D+/NUXuw+Yg43UF6c+2t
53CW5HHxPkzH2JW1N06ySDzWKQDQ787qbGpoV6P+EM2ekXhOm1B/T64CT+LDtjcQ
FWHnDTo2kTdmZKeFhnyVEB4Sesqd8DK4bR7FB54wWo2zwClKfAUBAxfUFWkrN4e1
1EfnelXzLCZp+JBXv3Ff/zD2N9xUG02710//zMmP7eLDCFyaYXWztDhz22bDK7bC
6lwntk8Ts4v1NYm1CqnQKgJncmxRvONtKajsPHTeZO+BwktR9uum5pMEXSm0OCGD
V4J6GjmvW1q64o5shLz6Bvu25XhfqFEC+sXZqPtHN3lt1FqYxk28N1tH+3TV5yVH
hwJgxDZW4wp5SL5X3W/yOOTlvMoKAz934C4jYT4HmTodoJLNeKYzKDsoNaJaPwKI
2axZmrDzRw87DqdiuR1gfK4YHi3Z0kTRUXvmkIZu+AApXkbSHbG+86mMGDX1Bj0c
pvULyn+VQDoXhHvuIjtnNkLw0G15rDSNxEIn8wCjuT0h90TCrURkdJk61FUW4KgK
CcgJfXcXZi+ZjvZshhGnrvdnFMFpZh0Zp08OcYp5siONJvgQ0mAQiR2/a7tApNQ2
UmvnX+pGntpLzB2r1bf6jznBV7YTA74jxi0b79XCJKIQL1OjdbXS/xfgO1uXGZw9
XER9aDov8r+TFyngRgmLhbV5jXOEv0aOCDQIbmuZfMM2qqgDCb/F/UXTZwYpV0JJ
BkDKhGpSh1KYrVVuVwqXR86Q0li2flooyQ6Xjg6OA5Lnm6bSMTReYaHYsbA5oCoG
qyuopYysiIGA84mT4S2eGPzNEPN/uOPncxpIsLsKGHBB8Sd1NgtFtyEdBJr4/bv8
qalUbDYpCUvYFfrWSD9qrPEYQ07wZzTWeYVv+yuaexN2zLakw/StsfOE6R/16UfQ
bm31tqvVB1Cvk9PuWFr/HXtPwuOJB8tscoiJAmk1DioXKjtCR0iReRzP2NDEwPHe
AtezP6wAunfQs23K/BlVrVAH8LMtjCLasQiewWFT8uU1piSyIDoi1i0lY2rDToBr
mN9IUllLRLJgBHQUV2+VqU20z5a6afykeMT1WCyaEbrZIEukbn/uTZhdHSvQUBRT
1SZWhRsD9o5UwtLRE+BFj1on/UVt0l707LRbNsIG71I3NBNwmpxdh+8G4cB8OC5u
SSTHx61yPvpYvjYUg4bXs1LYy9vVNNIwayfcQWyqNS9GbLNQeh3Z1zIfUmwjdv0i
AlIrp19U8nmdw6n5JUQaQTirTo2DHemougPcBb1fKyX1urCmAKUvndZc0wuP8UUD
yehXwC8KF4iM+VN3Bv/lvsZ5YEsmRppVmTuklG08hQ5efa0Sy/F+FUAnaKavvTCk
peeS02lV1VR2BruyTh72Y8EEuNmV8sdIdAhzXZNHO7ilF4f620UoOlk9MSz+G4bZ
ZNwYTP0vAJlJUW0PEVJDm5ApNgn+drps1YG3SjpR4P/e7TrwDVHV9SZxzGgw3YOr
vF4MTRnegjqTr9uDB7vn69eaP6SGFqQdfKTj19aa0FqucLVyhyuJtL5vqmvaqm99
O2qQVJKzSPGpvXLrNg49QP5Kpf2/iWdDPkOo2J8iV1uSDjviT5q8ksGrAf4ABwCL
T1yZ3Luyc+ZVvm2CM9YGh0PZhQTgaMifFv7JPH1H6eucFl/0h7KpvPPToprdzraA
ZmvbcZ8+VtYZylQerD50Ac92PT9aJrG3wJBrbRseolqt21wFbYKtklRK/ibKx8NC
d9GUplL2nuluZnCvWLwsllY27eUCcjfvOAhntq6ChZymRt7qoIZpdp6HwbeOewXk
SldBNopdEL3SzJiXRBwiMQYTJhrucOvz8jzYZphY1EfkbbOA0IbKbklCYY/EVpJn
0nDKGGWNyBQRAyyj/qP41xeSrk1fi0dBUIOiccbwFRrSrQc/Jd3eceE6qUyKCtlX
wn9eyaFXQ/AgrYsr4rZA3BCJ/uQ8C3E5SS9s4XZmk8Onmkk4xbFTKw6AUHJJBfef
IHCPXqnChsiiEEdd2es6jTEAQt7//C+250JYYCt5FRypRyQYb+DAaj84yIzLp6Oo
G7PedK3AuI099F00Nyllv3YP1nm3l1gzQEkMX3t4i3RbzJfEQm/ngN0orrJL4yiM
Q8PCkyLdxIIuMrjfFQyy1ysXvDvgS98Qgb08dVd4OZ7CVZs5tsoWaCsSUXFQU67Y
6qliF5DFHtotrlUPO2IEHBCRCyGZPqiQ+so3CzXlr/0aYy31NJlIUuk+Ktd09kVM
NAZC/woGqVRZ5Z5O2r0D1iP9fbCfw+Ypp6JALNytWJFhmoT/XakVmwQTSs7Eqi9Z
Ei6+/C9HNlOxQxgMTmkWVoc4aRMEZlPlZsOzGkxL5kwSLI3NM7PiVzsUhR74+MbT
qbFvP6izhs9Fl9/PyhqsGsmXL/tlrZ5CxYn0AfuPVSZx2tg2v1kIkHK6QGFQbpTj
tpTT7vG0ep8qZKPIKvAFSxIvIOB+2zT1hzt0Gwa9R7bXlOp9b2yooaE2Y5Oo0WgC
JRDWIiV2lHF1VqnbJPK5haZwRO6cxWKk3xdab5qheq1D41wiXiLvxwfJlHgsaAdy
UurQzAImynmjz/VPEd4YHdfoKgW83yXMlBcn/3/JmDv/DUb03O0mnVlAI2WdCLSs
Y9AVE7NvaijiQLH0zicR1nj3/BXnyLTyu1vZuwevO45P9a3SQ0xegbx1ux/ChinO
PUYBT5D+qVCQib3Ej1RWW8mi0BbausMibjTsrreZHvmLx93kud6GVnyK6YrnrfhD
+tf2BTuL+4pxzA+tHbUrFjn6nCKFcownJv7VlAMeg+flv01YAXCKy8uY+EUGmlx+
oCXnYZZnwdBfJwZy/+kj6oLviCyHXihZ+aChkvacHu0zkJMPBhf/Ge98d5prM/iT
iBjZydTiY8wB1rg6cCB1c4dQAjOwNW1KAXXc9FfzCeo4zsi3ba7BOIT3c5jTEb1C
sHejj4csyc87Y+N/zvkAVnx1oE8BrmY9yQLZGx8jC//got0nPMuvuhlPFP8WjKB8
+erw47a0xW2UaXrOP9fhZJaOmpQcjsYj82Gk1BRo6GkmPtzpYIOMVqBhdHW1h1Sq
Jpzq8uEfPLK04aIk0N0btMdqFQapQwuC+osxPuvuHL/3q/RjG+l3R1sP6FKGtPHx
ztSDIpPhWvQ3LUod925w96eriNGRtFmBrbAR/iI089af7r00MSkF1bcACEdn2XbS
Zm0whYcX61qQ8jjm4A7X8HGC/cD402XagIahW3TvPTRcdJNS2i2FZhX3QCYacIRb
ylWEGI4S4ktYAUEEGel4Bvkk96Awd6aPglHtpuCBLd8DNoyn6y2jJ/bNK6e07UNS
Om6eh09Y+ln9GRDU3EB10TGgl0gkGtoRsgvFIHXE5fGwxXYKgShnotF1dUE8oRJz
EXkqMtzBDsJXlV+8rJC175cy9QdpiaG/vBlzKkDjZOnNgePlUu+mKcHl7JZmxzai
qH4Eip87/lSNA87alsKYO31aZBlWfYp1VrAvYHoPgT7ALlNmY3HWsPSp6Ny9ySlI
GzvWlH1K+euWZokDSRPmpE0lyd7P6tB74xJstsySyrsPDZrQJu1r8cVrceK5zej0
RpRdLUdgKxEJ/s4aLDzI/RVJugJ+FcQ82DEco6miRPghLZ/CH7kk8FVAlaLztSOe
7lpj5MyydSWv6VaGX1bSiCoJZJKIFBAkytCRbCvgvYNxYRcxvadoenpEK3hRcMWb
45fKJHpgmD1fxUiMzWL3bSefnPOTXgv5HMdUwNWURJBja7/EtxThfdS8zcEEUZJw
nP0W0/42Iknxs50AYsDXMx4fCw30l7CfSmD4SZ7OhOip6Fi8ecGn/jVKKUrkrbV0
sCUjsjgB5uTFyujUZmpqhTg2wMD7ZXoux9Lljf3N968QcToFNwY6XwQp2jMliCap
8w9lWwm9mGjpghilSL/TUS5vLm2Bqz1oPiO///J5sYjG6TvC1x/P5wEFTg2eVgck
Rfbnfq9UTzlRyiSnUkPIzrhW8zgppmNXspjTcVGgzNyAJASJbWne9Soxati5yef6
o4z2vMTOq8Wd6P5PiC+0aVkajsF+vdK+aMhhnd/P3zbmO4uFXUbjySqmHZhksqEc
k1XI+3RW42geYuePUviSPZQ+fg9ibpxQeb/xB7VaJATZq0bkqSEh5LqVC3FLz4R4
zx2sp3Ok9VZuOHe9M7eiFfi4yMebkFkbA7vwUcZePsx8msTvkJDl4a+NUoSnW9vH
ye2/VeB2hD+WUoQpFT8K10BEiLtj/0ie+jFO53CeK9AGoYP0TxrXep1rAJwj1BMM
oYsXS27k64xZINQ0ZKvC6C2tA4BbHuShm22sNVleldNK1S98n9UDk7FzsH6DKhYy
2SLFOYwXH/BcaFOJyNmP9be5iiKYC9hR31ROntACN+/K6ppVZ61PY8DIniz2B9jq
Jg2ZU0x0IIGPNSFp9cQ6QL05YYNSYlqiPJZpDf+RrcUTzmUs6RFy0dXXTf7dHGt9
Fvr/14bM7ymY/zwzHlSuI3sOGHaN1aNPhVaEje7WkJpl4p+qJFT109xX0Uj3y8Mu
OwLKG4f/aWzo2Iz5goc1t+PTfayYuW48G90BXcuZ2YDEHx6Aw0fe7xfTQ/uEtP+P
9Gkki1n4dKnzPZAjVNBioMHZiNcqwD/eaI7U0FhCllti4ZrHra+jPgWE+y+FuLQF
PeSGsRJMLm/Uvb+J+zAcPin2AUmPM4D+fYDFZEifIDjR+BUiKsiokaObnkxjxsyP
RBA2CMJNlPfCL2eZZ9FOz8e1RK0jo0L3P9FojQnUaPuJd/0lwNSOkmRS8KawTahr
NS6GWho9K9BIzB/CrROp16+7LS5pN0Dyv6kka5CJVxiQvMKq5T2DRK9FAuHpZBtb
KuF+87VOxG35kuwim9JoPybd1SvW7iRjFOk3HCH+4MMpoe+Cn5KGHrJCWAgiH1oQ
ViLoDK6eBocWXIdKy9ZSTHlz+K+MEzYcoCSLOCf7tJBBLMsaVSZpzSHX5YkzCvlw
8iPxoR3YbeQvQrdLcXnkjAp7Y7o8QkcwZNeqmmF8HvCZJYkhybJ+xb+GJ5NiGeuf
ozNPn7CmOYpS2kXelQgxUh/s1eE6pg1OcFcJ3cEdOCejy+yZyIwZE49sx9povwmu
yyyoPTvOE4DR2VJoEMGcFjot6XieVwjlipxbxjdMrZ1cMxkae/Zg6QGm9ZsbhTwv
8zNz69lw1Dw9Y5hrLFVBRH3x47Lm+2S/zTx6rUAJz4MtRLC0SuTgIK5ik7DC79IR
vkyLU0XkUz3t2xVNBaqO5mNfE6E3kZJTvXgbdp46+qF3Uf22Lg2W9UPU+9FUszCk
r5R/Dof7zJ8ofQoulaHDR4wIhEhrxCX2rLgfi5RkQgrG/BcWInRBfw+FwGe+BjEu
P+WPxL7aSjHtHaVFNfdItHfiPVBWs6YN8v9dUyxnz+gIqo7JwDyud7A7zgCidw2J
h812HPrM2zN4+PxFTzugc2ybgla8cfo3C1vupFaG0TMXri/3Nd77UKcI/DZSOQ7p
/GcBElLw5IAizUAleRPjjhBwrj7gjSDOsmt9a9ryWNUwiiMCi6IzfPNcU8l0j549
DZNAJoruCANpcedRe2l8shI+ihfHMtjN/AnXm8jygLhonkT4bOyqMBrp0Xy9IGYb
4zHpKddDaEAiq/7jfr5z/W1mXZNeZ7hpKpVXXsyCOqf2Bo25kKqbwN2cPTX1Jil8
d1ISR9DHi3KNgSltQuuQgX0FQomVufWJ+jFHeHIXMtNKbyrFbUPdY9pdiSZr057E
QiZHLm/9AnbfDuG+XFLJ21dMtwpqHmuqwDC8XL2qKB+Y3uEGJ+XxTqj2tg1n2LgC
uaeoE1ujFB7ybqDnDxCnv6XPAjHl6VTfPCgHotmH982ibW+WvOqTYInS3JtSG+2f
HkU/jWGU0bElpQsNKjpGMIlYelBKEChCY5S3nJxUi8MmyCUca6Gq6P+G7cpxePrK
8FnFoxl/VJeCbPDqUt1c/vxfHjm9qZE6PU/qpiSZZQuf8iJR7SSldcPt1R1IRVoO
rfNKMAnvXg6GuNwKi7CGsWx2wLxGFEYT1tUqGr9EAR7K+SHuwr8y2iJO/wsxCXfW
wntslqNUTZ7zd2Ti8z7vmhj0qVh83hqBw2m1g9i7NSXpbtcZtiHjY/ZO0z8H7XCi
O2+YuuEvMyP52/oBPLCmtwmtWPZ1fi30gHnNvZ9uzD3NHK/eEx2wCTfiNkDDqNaS
J6Z9KDtgpo7PiypeX2ANau5Kea0AeWNrlhcKfh6z/dZDvxaFonZb0NiqVBYdb/Hm
kzWNjk9pukYabyd7Ea6tsIQZqVGEifo75qhsnFj7YSxWBAzuTpHdU4Mgaz5qVQsz
amH49NOjLTTIl+kh1ayHWdEefNSFvQySP8qeu9gpLnEg99zdn9nzVPl/gM4/R0cR
rACn/5PQtJuubwCsS56UXozDWRyH4Kxf9zHlRKxivJll9bbpUc10/u0e2AGWDzcM
JzxheIVjzMTIDrQm1Cm0+Lhg/BZk1KipCM79OaCqFF6U5NlaQbspAL1ULmbuJs2Z
utCQF+XD0y+MbNlzmPNdTL70SRIBAiatFahzdrCpKJzqXq0D4LbaeQPWD+YCGJNs
H1J7gnn/CRGfJWqR85O/heqKOBVDHugEF20Xrldzq5yI2ettIFm5Uq4b+ZdwVKoG
7BVpvvFRreHSrp1mjnY8WnL5XVxzYoSMT+1FVvDOvtnGb2irL7ZOyu9I42Ds8fFC
3Ok9Sv8Up+k/49IitluY4DopVzwc8/eChpYBXiomkNi/YiT6oB4Pe5q7JHyCHgJ5
q7GIT+b0pUH69zWhqQ2WaXnX/iZgMTDOpS4ZTxpJnYrQaBs15o5soH8TjlzSDcWa
fuxbqgtOAM7BSAVYbfelFwCs6LO5dzuZ0cPjxaOgLP/d6ERsh+GvUt9yZERkyDWD
N0FR5PzoXAfB5JxUaPjgr8gyrrFoPZQVwLoc8R/3T/d6SXOQrhgWYxGznEeESeO7
GzdOX5iaSRObMqY1SRwwHxXwZDdtQ7MGAZQx49Kmd9yCjIX9MwUhdhXbmnH0L19H
1FRK7Qcz9gyOfieszNZUFgt80iRw7FE/zw80BV+3pSG7otpkvI8V3j57UqG9GY9w
ci7k4kcMWjER5ySyaOkl7JdbmEHQUSiVPPJG0iQJY/9EIZjJCiKP+NqLTeD2vRLr
8AqmLbMhXwnshzwUGn9oWZSLVZSkH2x7HKKuA0SYDSfgoCIEp6zEhvr+owNxofWt
Fgt7sL2lxb+9NX5Vj7Nm9UlCR/leGNk0Etp2KGbzOtJtWQOrZSxzdgWYVaaTxo3y
yTHSMpxIkp+KczO7YctvJ8URQvAzl247LkBPdEH6d6Iu49vMPtF9KTdZN/aw6NvG
u/3SV+JAcTf7OjHrPkDqYvQyevb4+jo6R1iO3e+4punY3BebtG+yAan1bEqPn9Ow
GZNLZCTjs9hNwn/iEJcv73e/hdUZdixgoAk88xirWOw4IpMweoiWrirXsxLUuMNL
AZD+DxNqHGcKm/R3+QtpkbLf6D4RqPl9gRLh3s7/p99yNrTagUS4H7XhyDKDGvlC
vALn6HG9umD1ojOykyu3o+Nc1Rf6U34lJ2HU1GpeejVySCz1RntwkS9L12lczkNc
MIK2XcUhqqfahFQVGUecn88dEnbHacOS4r1o4FpLEXVcZfuCYimBurY0c1B30NK8
nH58K1D13ZW4aFj8St+dpIm729Hk/HEYLtwXYr/iyAP3mBgbMQO2IgQ8vcovBXgN
D0M7rUU1f3iu+gXYlUawbeAJqQOCH5WPjKdhwePvUzAoEGkzmlssbnkGwBmEaY+2
BUc1Nq/ivQJ77i3SXXpb7aWMKkJLDV2iWch76xkLhRGbHhMx3oueqC/TRewi9Tga
7f/umdQvZOx2znXvqyfvTwyKB9SyqaO8I+1jQLHeg0g/Q6tdJMW2vUDDHaeyvgMX
AR5Zp6PZ9asA8EEJslqyZG/VmQxmSeAljlNDGEyWWaBVXKt+ttBrHuyhVSTGC9Xl
xpkxpsqaQmOBkQhpDas4+h+MJtAWZ1Jjqadbo6QblL2On8si1qvY1MZzLO/WaouB
q+LObKoyi4jYKDZwdGjRp4FvBUgS/yfP/+rC4bDDp7iqaFwQCuXDeKkQtg+7rmYX
KFHRGf+K6F/GA/GKKrN+KJVfZZiiEr+Ln30M0fpsdbYY7Vfq3FY/uzYZML1BFpQh
E2sdr/kXxmYD0oeuLoQ2lsHiRVx6KNdplMUFyQO71SNU+MsMDj4Y3+Lg5arzN6hl
4CiD7I8BjupNZ50lkt9rsFn3EYP5rox/Kf6qzohVlonsrbBy41O+lQIvsiTp/flL
aChk6LhU1gU4Xi1kBrYTT5Fr8s356k6w976fJPy9qwYgESXw0N0CpxfvVJ+/iTjk
z7KXQRKGy7Gj8UjFETzDQJjIzoyF/txk5uQ6GJn+oFRk/K0DECPXNiT7Sw0M1Hmp
ex8WHc3B6cR94FjBGXqSd1MsAB6QqZb2KDHfEEh2e5RgSYupo+16I23/TEVgzDPJ
Tq0j+c25l48nXnAycxCSzf9aTxUMT9UAlQozUIrdJm8kYrfiEUbgjcIVbVLcZRzS
zmx4tXarfABi1fjAfoFmhyCcJixcrcHmq/bTVBUkQ4QpDLFknWon1CCBRuHG1Mr0
6vhM3WI7ljJgIeQEfXgjtwjerCbCCgk3a1mXOJehsMJVq1gzNP1RlH2XuBaSZ1e8
felYYhDmlo4NZSDCcWHVVh6nhVF5hhjn/gh0IZumtBssLWPaXU9Y3tTeq9Bky/Ki
cmmxd37oLUEZQqoHrRBax2m6kYAfN9IJ8HZ9Wc2BJ7LzIadL0rsEUOoS8TXDVCQ0
4W2Um3Zzqa8RCOlywZiHtC1vG9raMTrcMsfn51Iw79p7+0u35x5TCU7wlMNwwWmo
eD9WkbF56AxkhwS2XPkmV8i0dm5XKjeEG3qnM6sWZwPvcvGlMzbhDAO3MlyJMnsE
bm9t2AQFVJkAtUi7lfbJmaaCXtGMoPz/1C2Yc0cQt6cGYVRuco+1fwJWcINccikT
PG3yks3lsehDyIyiBFakiziZH32zmzy3g5EXINKQcYj4wdn2GqO8T7Fi4M1/5HAO
1EcNP06JE6Wf6rMlrqynYtzzg4WKGUZ9yWAhzrbOzDrTY2yu4e3658uy5RGl+2m1
jdqiJgNbVuQg86eVLpc3cCnnQ3h+qFsafX1ygTtFB6lZSlxP6y9gl1IHEn4GGRJv
NssWIPgoyxNvfsSHe0VWPmJ4q+oM2MKacphwuHOM8nN1ryHGlSG0CdE9D9oyyeep
PrKmxy3gLwIV+1FmkjFoglRuHYG2XM33oaMQs88r63GcGuP88FZQxAVw0LrHTX/2
SoVlYKH8E2+q887QC5hIz0oxh1+65YgB/PoggLWRmGjQlUll455LOEnfGJripsQG
0wRvUBshkdsJZYksEWltmeQZLGuhhkJkTqLTnpiddUOiHS4Q0BeYrBtTucAfLWQb
CBF4uIJzA1qg+S48jnmgo5D0t2iQDv5cP4fcNkNHR4kXSTAnUXIkq1l1PfBhJ1RO
coYrRy+iniMpdlCDysH6uiG521SMIVWNc6QtvqSi/2yViVJdLLuCub4QTXJRM/cw
AP1M37Ec1d/y2oDrSA9emTR2Uee0wF2wVxPzIjn5sCn85DI9XH9T48ylClODO6TG
mmb3k/WKmmK5Z1GwLUgHOP1It0qf8O0ANAJPLrddQRqVJ2eysLfNZAhhaCesFydz
ZuZjac2O4F64jEUdBxnuoLF7ZLTgOcVkKnZDa90/eBZpLCLH5aPfBbiXMB62zTqa
9H1s7e3jGnEJy5fHQhpemjnzrbU10MS8GaWLAtaVSCq4fITgFrOzwGbaoLf82Z3n
p3mCuCvDHncbJv3NuaRXX0HvJaFFFYJrJS3dzOy61UCHRKbJBdJ4t+iHMxvMhizJ
dxBgmqKJjZf6kK6QG3oRKJnsud+yAL+9f5GFj1fGlF/asN9Bge8kP+xLwLoMlLrd
iE3+R4rV0sq7NtKer3D7TMPWWD7bjpTDWeg623geH9K0q2Fa08HO+JKY2bwN+wsx
UFMuw1alktnCKgW05i/47a7dtFUZlp1aUnTVqnqWRfw1/aAgdfzLp4nYf/JojQ83
GV7OCczoIsyMKX1KNTUDxSDA3i8lRL6K+qVL2BEitiXCfieH97mvyCD/QI5iYYA3
YNzdbBKIuvWMYeHGtIPF6hRnNdo7FYe9pZ6fTlXFaH3GNrWROW8MiuuLQDSYpuyN
jfDi+9S/hPmHnA5Ruafbo8uvR5Fx51weOz05mPPYcou5GeD6EnxA0+aufJO40hke
ZkBwc/LncNQeFPB4/K/z1lbJgBPznUKXV++xODSOje3e3HW/PFmcgLp2vBoKEEBb
XEsq7QVXUhp4oW7l4AKIyaAJD/DKEwZnAZgoUWYH0ZglV1x2PdgJvuzAku+NVImZ
slOU7ofhjV1qneQ5mx/CNoI6Yc0VE0zdnTv0Zt6F3BcSKbzdIIwagV1CvxP1t2ee
3DRwNIXbQsfUZNiBA+r1qfV3jGRLTORSNzZoPincLEB1d3h++amqMUcqB9NRMUXK
GMapnx4k1z1VqwFFccnxlQNXGajR9ttZOuYQtN84jGXOn/erFxGbPTqalcY37JAF
zsvzxlcMxD0ZcLtZncSGaCic6NOHMNY/WQzRg9Ed3rhVL3gRnE9FUWzi12ZhQs7v
kok00s4baeAw9SpmL4rMLsqO28XP0VniyUSwAvy+tisP4ItABYRD4rxA/oT8o1cA
1eHlndzHCthPXaeuc8/qK1JdIqfYos4DnR3UHnE4Yo8vEkWHSof3YKbZHz2wbTyV
ONI4hSXQQT+59juWUkQdOVst3iOmetj7s7Z6drAXFdNmIAxx12vsFyQUdAw7rPGg
/mZu3qpIIOfE4ku17OXOEbwHMhA6jZ8+lid73Q0qvjDQiDadFmOZyK8uO/UgB2n6
u5oHXlXk6agXtS0U4WcEIfm/SC1Y/trxOFdP39Q5JsCYcxK6zRg4pW8qVfYXfBwd
C3edg5qamlxA9tAFf5PkHOKBwWUsGjSVj/sDb/vmRII6bqR8X7WKgVenV7FoyWR3
BwM0kocsJV8ufNwixtDcnxL0SKru4eio2gjvinYWZ6HYn2zApERBLtg/Ni78JohF
gmfw2gs2ukYDbLZnn/yCmt5zsmTeNMRFNnON0yd1TQhryvUPHgeG17vVlyc8toJR
RP0r3rSeofzHmi0dFdWUTtpAdAIdJGT2ukE+d+n4g1/KWejrh//i6W8eYWAcLDIZ
SKX83DsguG96h68k9Vu0PtYu26oB6hxOx0hagdWLKQABOEqJFs95A9PJyGocOhAp
daQBNh16YafZRTZVEWwSRI/0v8HsDzz/bwJNt3Z0z+Qcdaun11IMmykAe2dJ0Fd1
HNwkE85ckDOsK//wQqB9rgWflDPHGb/XTGT2ECkZn9O1nL1beZYDYi8R/Ujrllad
9rjGkJ9blPTDBFheAe86A7G4x+mdx8wxzYG4e6O620zGz1cdvmfjrP9fTRK3uSE9
/xprkAM9ElF1MhMaMgnM5ua6VMcQHNvTLRAL4JLTV60o8gW6aOY94koroG0kIv57
MgmUInD9M/x8XwN8drHYF/ncgWMyq/9pvXzWaKcs5bTvnKSAaT43WQv4S4AZ4iMc
PwjpAQzu3WyJJmD9CZ7z2AtaoVtJblMN9EXlSxj2PXmSTZhTd6nhBs3LsEgRA1f0
FPZoHLms/QdU9LqtJRvUcKZGSRwCXX5knUlI8ajibXRZNdpORTBsaEKCAOI8OqGH
hUcaSTmV242HkxDlHlmrQg/Qdr2H3/snWlfE/8FJdiMslmNHcw6gP1VNQADYLwhR
cIf9+oqzARkdw2+DyHnNmPJU+Qjj1cRRbaEPX+iMQl9xGuI9IdevC4a6oDZqetPI
3f7R2oyLoa5XT7wzsvtyMdmvBsA374gv889Vx2I/lJ/BzOjmZuLWFZKL45Q7CbgX
Bo/HGn/GFfkungv1x0cDZkV+hQCYYPunlcmphbUiyv+mmul0la6mYtRFpxyVuU90
5kGzyvSAnr2FeuA5k5yQNA8Bh0u47BcV0hr7Eo6KFhrblKHN63HXdOyAJH3pQ/TJ
XSYp1qt+MRq7AUWaVFiwViFXeH3D043DwnZ7sgYkpZTaEzASIi+ng2CxPabsR+Qn
CnOvmgJcoRTeD9rX8Oj2P4HasEIsbIZUIwt9NvLxqVovUl0zi7O+wHP4yLZ0Ydw8
SJC3n6CHMpnZYqxNsxOkO4o+s7wPhbsZ1lPm8Hqn+7GQOSEzjjOIRVQKpp8e+7M4
VwpYJzl/vRy6MRZD0HlNZOryOvQ4QZB7YZRGbRp2z90gDVdCzCHH1TY1/U8ra6pz
qZfz2yXtf6iHMAX1p2hxplnMV7kdk5HzgIVdCSHxa0RIN41A7cE0QMgC/tPsi6vM
vLtJYayPUr39lwXXCGxXAVip1MOCiV3SAMJ9rrqXo9GkTvYQI9zgdd/GMUkruwe5
naNCmvwYxT2RvFTRoR68XifyCj6bL3SuGE7uqhPWBkuA8ZKwRTV8sAx5iF5sPr5D
ACQs8acg3wmZSulF4Xe/mo/OY6IPBUIzp+wy6X2+ukSwkbWvqNydjcZoocvMjwlq
USjkYNgSPzoxe6GS0cgLKutrDkfO1pQx/DxldCdx8cyA/XD4B6V94WKcPLSGxvR7
RSuD6KY8vaYEdG5OZ2mDnCVM4tAdLpuxrVmeRtudGnI0iO0s3AKimlfDlJSc3H6C
m7A5lKrpwkq54Fgu+EvIi48iATrJddKjHZGy49rb9DPDrPeiRuqWL5nd6sTYWLiw
Qys39SvBwLjBFeTzYF7CjCsXCMzhu4AkjRATIJLfdyLyWDlLNOutQzsck5MBiakI
8PYIE1OfYXNu6FfmZU27jG2qsFWVhb/tA4x7jTM5ro410BnjZrm1GRSQ2La95Lfk
ugnesim1ClqydHwwrqsW0tQSAkPdTNIFfQBhPGo3FydN3h3a4jsBWXuhqKVEYYhO
46OJWXjevdjoJejLTgpPA2mK0W66NNca1RSv0cTOVAJE3tmbrOibrEA1YA2RPzO9
QtGbviO/BV6Xu2Lowa2OqGsHLlARkGZufWb54iWN6s+n1XQQHFAwD87BiO8a8z2C
zsr7VaIreuqkGI8ubYYk3F/0KSxd664ugILyC4yhneZg/9+bubv4sszTpp6yuSvg
YRG9akP/oby+IlBYVmb0GKo+rnXRDN7TIe1pAgiDWCFTRuZvP/JdzwD1AXBWWdiw
LSD5/fNTm1J9UTuvEHfRmyhuH0crnXupsGneJk7diixh1D7xiJEgYq08vlLx5mox
FnyTy2xZBwYlR+y7MZarfslLL7eBDk2K+kcPK6/NVJWxE0BHRjgWCAtX7qMG+LkD
k8NbY/++eYMSoEIXDg38i6U89Z5+4In4gW3y9foILoAOoOVWKGUAgn3SqBLrSJj2
4rIfi/DCg7FMH/TOtwbHha3XBmhbYUykLgdc7Ax+MLl3SbdYpSIsxxw+SiJjlFyN
gnEeOZ7ENTZJ1gHBXAiqWx+kP9FlRZUZtX/N2rzspRQBiqzyuA8me+hwAJKXUvNr
aJJ95ZhyNcq229Qxtu+PoN/XjtB18aT2sHI9/IxgAVxlVqVMqAHv7eH1QjFGslBB
jQ2GpH8FgJUd+6UbUuSEKiCwVtCxp4qqQ7m5bRHiq7OV4mgazqfBtFEFoPuCQUbb
byKEtwmsp+yxCDxL0ITYd5ePzaXf6M1so1xJq8OcuIuLQac/l0YnWK3vGSrU0Jql
yQczSiciSpSS1hCLBRIDQy19u1bBMShWeKq0mhdpTYYFZL+gWVyQjMOc4XixtWDd
g5/VG+/kopEdVLAkWmNLQ9RgR0vgn4FF0vYTgAaojvoTXn0VLZK5hgMYw+ddjxNs
N1MSKOWU+p0chXeWgmZ8WVa2YQlobuFgqhFcNDiCBSLy5+o80tho8Qik9/WJV1rM
qoq1xTK5aiSl0qpy1kgYf2EJFFKSelkopFGdb5CWV+7PGCvJSGA8zHcUJbsnAQzH
97w8DW704AQc8VJhgtk+NeYXbo6mB5Xq2l4UcZUoEKjVPkzsiEgLaYipkRhkf+w/
RYMKCDon7D8Lj4tM2TsxkqHzX3TGfwo/VoiHBkllbG/VbPWokPiqSz+lUnJbS5i/
ijjQGdpWpHjZLu117R6DUtwmYyCn8jMEVGkv/jFp11uKghbEK7QIrlLxo89vsl9/
GFLe671lqJ+uZvNKLpcQXe0g6m8miKY3tctMS6nGtxlivVIobHVSpePklawMumk8
7PgMpmwFat8SiN7bvgRhNGqZUF8DLv//qao6ixeMM5skpFvaJjE63J9RlQvprZLE
xLAebtvBJ4T278dW1NNKKMAG0N5c0rtknJR406z6e9xTka2lU6GXCQcpMZeEZkaW
mdx9CJDo/E5qqZKBm1p5yES7r5l1st5qTCv+uw7Vk2Y9n22HGH3GvoXM9rliLJ4o
xlacFSxZ22/HvPIn3/06U7OdVP52WCFAjcoZvdE9Z9O5zfywFZe71YNn26rrTus/
LJzxNTzTaOCSFn4npBCz6vRwVwPtcsMizORPCjzccTFSsRdTVbUfPFsIdoKrib82
V9r4UlnJVsaTlzZZyFpizDgzuuQFCDOxIdAELgJZvRKVlBrrtuXPuUMWSlxyF+fg
GHXgv5wqgnWQU5cfNTeVSx1vwSFYJZ91kkic22Ocf3uusjc2jkol0uC2hVlJ//0P
GKK1Zx3W2i69r9QApLQHmY32c35zmuVTKQFZ+CEfQ9ot3ShaEebgA7fANS0G93v+
9+VrUWXyyPWeM/RD/g2dE8QbG7/P9C9kfKFyh6tk5QGpFGsTd4AZyZOSeyhKS8+n
MrPWFq+2vIF0vbnjWhngBsj/oRfKYycyadaS2t6R/aJzMSsn+Kggsb92lgpm1Ecj
iWPaw51j5pCaGLrKGlqZ2yRAxEWSPZck+K6vMBhh+eNB6pP6/gmW/rvOnSjemGgH
xHb+23tFPdAI0HZvuvgsS2AkqPA/TVQ8W+GmE8KNbanj0orW/H7i/Vvc9IenmzoK
ZVllfR0gOnWQ2/l9HvxvELJRvibvUmRUdXH/nCriBhpEeRJmeatS5rmYq/wWS88Z
fCNlw2RPAmx4mMTbOuSjtkZdTgJm2I19y/lyv4CflmRP0K5TJ33qxr49EIZLlEIm
Xn25YYy9lFqPjdXvhe7x613VUtcNLVsbeXipbl5CyahFs6T+44ym07DTyI68yTVX
xco7u0DiZ4HH1Y5OZktgd/2xcWkBAoHO0vW7Ua6GYuedDto5kQE8hQFPbI1fTz72
uW/6Kz0oxbRPYeKP/0BNNKqe+rtiZxNrrwLo9MYhnhRsfByFDDemdM49Xfccc+kn
RgQqgkXyMeD1GexAanwhHuf3XmGnecaBwQ598RwiTBSvmVBCfS20Zc6ubwfcbJZR
+aXjyUuxQahjtS+XujZ92Ac+Eo6bKVESOcNEL/qvNbtUVBJ9w/u1Ty5AMj85d+Au
2XGc5B6bizs7mslOB1vta0jfH43p/t144ot5Agk3ny7ESPMqq/bwWo6PQPnDhSKb
32ecGxpIQHefR1abI3wQyhl1kp0QZXPFfLJ01Frv8QDsEcCpX2gpFvQIHmg4Wap7
ZjQ4B/Xt+8PIerOW8b+koHl9iZkEEHAYHtbxmSgAqTxIcOoRQpbFgnarZZRUOEg8
wK8d5FHff32dhGEA0IomBvVpxUm+Kyk8Q/8BMYXfFRsfOPMvM9cJWrQEa9JWRpaY
OCZGARj7NeaBP72JDEybTYNqyeVUjxI5ASAvelWC8cKAppcgLpB9WeX/RFWQL08g
csVpBg62IZvyJ2YMefxqH/tsJbBPhjzRjQN41MfYO5TGM0xtv2VNrEjGi8PPb9Dt
IZDOZmTBYZ+NFMQQ51g93xg0S6lPWo3eB/+AlX1P/qtPFZd3bulLRDBUWIz5H68E
8rLG7DyTstzUfP7Gvozg+E9R6P3zp7cMG+8wXu6D54g7wiPiy4wdp5YD2Gjbo5bo
sZZbMshcHR+ldaipQabVYwzIr7vn2j/8DNhV5GlkaeVg1XjHdK81IvNPHyrg3RWn
W00Y1hCm2NPMQlrjceGtXprHA65Jzpk4O822KLmEVg9UMn99gvE91UhgH7gfpd6P
Q7RuT0YPelkVbZV5FVt3q3ZwHsT1e33W87Q8MFIxZXD1JqwVsonu/8h+xIHxAHz4
ZOsNxhcbWaggyQY4vcQWCt0jo6RpHBdXEALDQgBjkjAXOGg5dFCR4NfuWJpH1orD
Np81GW58NkAEnmpkoFeGM6fRHeRLjPbqGJA/vmWvAH9cTxpp8gFQhk1ReLV/Prqi
E1RJKnx2nZwxSPy2VSNCJ3D8a8HBdPULZ6/lWFez/C9Hvg0kma78X/+PtMrQSTvn
SSiUwkkQZrxhGYXKtqA96uFvFryUOnmU8pMvRq/sshyFOexsZlwa3vO6e/GG15pQ
ype9PvH+nspyVWZSLbvMe+SJjBpA2EgTGzdl+rUtWamfMMqqVrSpcbS/DtLBj8Jb
OS7rTD3/QOaShSK0075ipdmvtAT/uL1CEZVaRj8+wshZ+Zp3bz6nbT1qL+EH06vs
F81FCfeddNJea9vHmEC+hw1Ps/oK0SABK2rx6YB9QBG5P3tMZSgPZ6u9d6nQIO79
Xa8+LP8DJys4nmvW5SGmpPr3Aru33Xpvz68Z6s/CpkoqPbAdBgWRsJqyr0BhxJZv
Yeh1BTs7MSeSXZAE3uACN2LbWjIsGpR92PZOaJsC2RO28jUgP6PA0z8zwh1EH5Xd
QLGEvFPjO/Nt6dXWaxKpHhLBCaRTN88RtX9IHoBKwWW27HVO/YWwTXtwfjLfXEiG
b/x3qgtcpjdcButdBRWUrXoB68lEUQbVzvgxdAqKymKJs3M34sh5z0Xxg6El7Rlk
UTo6Rgb51l6ibOeL+8nIVh4I6rZdqr/LU/luoJx2qRP5JMepGnkr7bRhPECWs5w5
W4tBHKlKPCTr0vYaVyEIlpizaZtO06xTgKGa+CAoriUX1AC5Pr0YnqZSE/ccnuQW
20SuOkjzZRrVC59bwtLHR9R1w+V4TXOtWsrcvvZBmopU1NKsnQ7G6xG0zaDBe57Q
Hy+vOZd52eVsoQ2+gEavgmce2tbyTAwMQ1bkihkQauA5AtTtjXiqGs2awd+aiXLX
pC1WPq0po78JzOD+op2qGG8OVIjbZ3JV1cWjLVXjG95EYS6T37970z3pJd2MKw9+
f9jD41R/Gyo2XrTXxzKtAYxxEpwIsNKCAyN0TKhD+FlHwp6xGJ2vNXvtiJHUZjII
ZY0xHyVbkYeXqL3vYCo/lE6/7uP67s9Gl0xjdrbmI4qJxCEP6BdrspCqL839v4cB
LhIvUwFgavjQaeUYmLRp9PimWkLdG3N6Bbhxhftwe/E8kVB7Y3SLgU+37sHWjQqO
SpgwFC0ZJfpA3ycovmJkP7guWsrr5KDRbtbWqIQvUBgEHLYAI11ApVvYGU7y+JmK
YIbv2pi+6/0iq5VdeVfB9qE0941zf2GQNcMnvd50XDKOP44+JsrNPv0U95dzsutk
zwkbQDSE2AHbkBO9kFjItEXu6Kgj9hnQYzgh69mDx39rve4V8SMwLgmh5FrFuNru
tQzsG2BtfLSAwDsYI5aj3Ema4tIxEZVo2EymHGMB9kqJj953e8a4PijzeaQyaC/2
ZSVIxhYfNfGGRJCE0fTBN8WGeqEPLGe+SNdgleyJwhxhLhugG1WCF+d6mz0WFrG1
xCS26mExJ2cOeSNTMxFCHcK6nI1XedpDtMvzKKz/9WO3qWhdc7DYs+LG02hoIHK6
Su/Cz8IUE5SwVWKG7jDuv76Bl9lLhdRaNgu6g8p/RHnyeuYyAJPV7p2L0tUrZSLm
KJ5hD4u9tUthd/l1Orgg8xRUdkeyfnlhGMHjRmNFdChjQ95uyaoW4SiJj4eldzKy
4pFHhW1OIka6RqMVtSx3QPSpWYHIOY+t+dKQTF0P1aX+yXUL0gsBdH87q0VFPMYj
1oARHZFIGXnm2M1GIzpJTvypk+2+jLEbqsGp21rScIvvzAGZ0h/Y7RVvuRPzCj9J
8W7hQWQySvBYE62aVAAF6QBS2yhugSbWHvLwWqxOIh0WMpdHKQUYpLgJZlhMHoMa
TnZopehOf6xwl1FN8ci0OCh/C0Vz6og/OlUYghS9devBLuzwZRjSuIuYnwod7MCM
meZtrdAlxwilRjkvVXxEJ7tqJ0szB80GSuB7vLb5TtEEwM1OlYBXXDOOdAndsrS0
aHYjmIFmObVZEs6T+tp2tO+gO7aEdHmUryg9JQYGoG8UN3gcoTicjNtjfVD+4BEV
oZ4ng2HKzqgjxqFYglQt0ALFQixXcKwKmD4wVXzj+01H+iNlTnJoSYaV08hL74n1
eww2PF0nK9mCBYybG3BXAUUkC4/DpEtlB1df9apErQ22WZ7TNOKcKcJyd9LSoVBZ
MXP1ekcVv7vhvJXDS21qogB0r5y9JxGlYEJat6huUY3ldIMgal30tEbMfHtmgkIy
5wwnGE9EYYPdQcFA4WRFUYtsZSol92G+qJx1CHSbX92nLsCaVBRWpcT54zsdQN6f
0+gE7+yADc0GFi/jQf8eWaroD3NE+ZOE9YoYOjPNQv89GOqp/wE/c5g+1GKGL/rH
zX5Qc4iHDLmVY6js4NejtMMgYPofw982ujIEfCnZZv5WpxS7oaoRNe//6ZYHlNs7
ivyiADTe824blchGTi/K71gumpSYNLwNkwZDouBoRaDsr91Zqye5MuWKIApp12C3
5tbSu9CnC5h1yy4jToNA1xq4MHkx5IrX1hy26TvICaaPRvKET5LHbE/VLtgE5yUc
kscDh7Q9cH0R9QT9z5zXZGiecGt36RM8yQgRz0SHq9DyTwskEAIYCJBuG4sN8HH2
J7+KSEegoVZCm1eyCtNjzHSags+Hd5gWMnwi5xRWP1PRXjymZoFTQji9Xp2n2DoA
01QD3AI3gPo6/IeMPsqF/8f9MGY/T3KltEG3NL7BrAB76qeaGqLP0wpzGhuXxtwM
bI31PWuegj9Pl1Oq5ICO6DIWlYP9BcoEXwLG8HiMBeyKrCtMNppT11bRKThT4Eu0
br1ySxi8GJWdMqlvh9/0QHFBYr4tAKbjKp0KPlSvp3QxKlRZ54IhjNUBIbc2h/1/
7DcKds3R3bxYxtmr+kurBAtB9M6ZJPcwkPmpfGYGmwm5cAxBTuUzGLMPoLHKf3SD
PaPWfmTL011NuzYgMfCmyEQzH8xaqcJzHRpwDAsGPHYUyHD5z416vto9deQeRxvG
ygMxnXBc66ddu8TRNb3kR/nHw+QTYwA7a6NLodZfagdTxf9RkT8pT+tKPdyD6mTx
642jesBOOk4sDCNqOB6zlLd/Umy1vhlWVarFsLjOyGbAXVSyrbSqsiETRhUhCwQ1
MjthyiwoLppbBI4oGK34Z8Fm/ZXWp4bPoE37Ss2TRzoBH7kUrHIUlT6ztvKV5IIj
DeiiqvvxbQBGXXkwdBr1FowYr5tanOMAfxCHzK6IiOO+mB7uXe+nmjtnKqOrP2uJ
srppWXfspWC0bUZ//3j19MzYG6vg80ddHyQu9sSJF9LMbnOW4yo0FjYuGHtY5WkG
mb7lEOTQEarkebGynR2JCMAhEOyt9sN4g1x4CSAtO1c6z93jcZuY2sVP5SItaZ5V
2F+zBLrqJWHk5pGgmovc9uPHzq5OjGoOI4OgSlByZPO4Rkz0QlBkExTo+fIxC0rW
Uh4s4b1P7DA8pvov5zcLn5KdKQbyub72g1V2EZ/cjYpqc6w0yr4NLCNsyoHqTM3i
Gj3EQz9XrNZ0tqntvfrdV+3CSm1mJEUn1hb1LBH8GnCMIWfYuTAT0DHHzGeQLD2r
36Lz176zy1446UCbHkDNY7e72iRuBhxYX/dqeDa3OIK42q+1h+eQalIyYB2TuG1D
RFt3PX89rZN8xPctYj80s16xO8h486jWHj52NhpYfQWsH2zvd/SQHmcU4CIRzOrs
xmUo8vn5B3SdK57WtTwfSUExfUtFAfQdb3W7LpZYISgL3lqA3IO1fJ7GNHjC0UyR
zjbtfBI2PuPNkDWW5R+g6WqLfJVGpXpfju74W8o/LzBffVTBP1WoDor4EPD4En22
XFd40SS4tnP0GzhIbBi1i0xoRYQVL9T1L2l66Dx/A8gs6OmB1rnU3Tax6UYJjNIk
C02OuAb1xOlp4GZquhVy3wvBY1n+UBGcQKBMyHkyjzRAMaP/kAhYE9FS7jTaUtoN
DHuStKTB7o1dw0F14BaT4PoKsyPTLQOvoyM/tU3dpA53btqdKNsYwm/hGft/VSGU
M3Yl++qGB2zndLezBl+w0HZ+3iMEhEbaDj4E8yXvUL93c09PjDJx1daL+yuou8tA
06cz8eq6ThbxacDjIYy1zf9rIVTho3IBhmpeES9GOHtdwkBQECwQ+X/3TIQGOE0C
V4BPMdbU7iHBLhafUZadovfbk6I5wSg4DH+qPlde3PEbMZYC1a0u3zzPfvtz+CBW
KScdH8k4jbVQQ06LXBEQtmmFXJP+2ZjePv2DYY30lUfi99hhaTiK9TD83uQpj3MJ
hgclq779nlojcgSDfF58UcEYcXAEDdHTP3DhSfynKaYuZ9Ui+7Qp8FHd6cloqgE6
zx+KNV0Mm96MccvoYzjBRa91d9NBiKsA1y/mN7cOE4dB1VxmLYOzJobj4XWn6l/V
vVk7q1vq/cvptF9EwJFJWzapsn5VwfcJ69g6axiqrDKGwGIK6cEOK/8iWjv9Vomx
oH8FGSI8KjX36bBG6pWXJCg6aUOB0Bhektxcf3/yeCRg1vZJWDNaDs7RLdGJ/Ozc
uyXCFEXoRo4tA1klo23Snk85IiHxUjNY+TTT4HfqreAJSK7ZPf4DlCLOCtvgGtdQ
eTtkRm0hyW92GfzB8uzNWBAAsdkdmTBCW61JdEiaQCdpltUIhOElTWyzteLFMnyI
Rskw8fNdNZJ0PoHF3riKhCAtgRn040UESLOuYNV6CFlcXj6IJUiFbtTvBmxEvIg+
OymPMHz0jeT4ukJFm8OJnAMs6VJyiVbc2RcNKyAd6k/0nwubAjoU4asNH4zWosAk
fLNxLibRDeZf1EoqUdF8yNxB7srB17hMbOIx4mJLWBYlzbR1m0oRc264d8O20WC3
ewRUXqB7hB84QxfqyyY39DocalRTXmABlC2RnlTkB6fee3eyB7AWwBT1P80VYkX7
bgGX5DgJvbiOfisKbUmbRDagSigmDCSJ1hmmEizt1Vk1vMm6Mi8nhLQxO5/UFqEW
OLp6aFAKqhSG92ek4SQbOqd6lcI1VYqqNBYLMgCjZyt7UJ7eIn/Th5VO/HOzpuRp
G7BYWvlDM5123TF913iLiNnkDqZ0io0DcZUJSrE4Q/YdQrHRxIBvE+kLLVHZwef5
Bcx3mMULG5f59xENlh0BGA+YbqDO6MVn/jDNPNrfDaO8V+YwltrQgwWKY1JMGcaV
bIYIjEGSUYI2n4LVDG5Ksx3BmYxFMNJl32n26lYWocQ74ids8oPyLvR29kX333md
oOpNvglhbN+D+fhlm/qld3uRqSwg5/O0c+0gjUnmW0HBFJ2IFbXqlno7IcNPFa0P
ZuvPFA5AIPqi24ug7PhEoD6pjI41mqALEZgbcbM3y0yTYn8zAa86qW5fqVTidcGv
WxqBH9Isys74MoxD2PuV9Up5gJ01M2OmDrtztvUCZMuCVO75DQ3tDdXepgA6nFbz
4XSZpsi0zBYRAuuTdk0my7nk8UXVBmxPzbSho2pXYzw2AGRiU0jUUNeIxDGfqjXo
XWGOzJ9i9TMRSwrRanw5yGxxMgj6fxsTYELVCvHeJKmbGVIdPKj3tjEpXQPqhqVU
Z9XuKkyfuFyUACQ3AttqVq0aeG5rD4WwwaRTTttwqG0UjjWTRjZz396fNIrnchSn
ZLoORmU+oyDu3pRa8qDGXdY3cEtcY0v/QtvqmgjApq9H1YabjWkwQrjsrSrjd/Ml
NNf7p16m6qoNbeUgoVKLLgNF76LWqo8kujhU9A6Q/8SuEUOncnfFfWYTOb0so61v
bibHG7coUGI0hry6Q0IL/y42vpiAMr3eAuOdSEc6ixVwYDRUnMehb+NFXgK3p799
qkVFTePHWH5ZUC5sP7mHdZmiLRJ6BY/nDciX/+aap1bmG+Pu/mkBLh2rTBBv4aw8
ck9amPyYUlo6L/hqQ6WdMYcBAGLF5WsBpeC7JNEiBlfPX4aVWRSk0UTYMeQawACq
Ee8lQ1Spx/2MyP7qJS5OHDS7+xOKYfQdORY1GCtKVrTcoAeaYhEGXtrc2NbgFMqf
/bUeV9oi7S+xwIDCHlyF0ETVv21KFoAUcffWT6AyzCDaZgJZ+9GJc2f2INyejHPN
8sE+ZJ+cjCFcxCIA0hl1roNNe4QICMJenEGTeomFvf6CIGOjPsSC5SAaHo7ygMBQ
w5nYO/5SAH3VO87peOfDgT425oQxGUOWEGnCpEkMS3QKqxacjFNjSdku3Pg7J4es
lXBCe948SL9NIUiUsXvOfTMG/I0Lh+wn3bd5RbYJqLxwwejsv1YJ1liEXAOSJlv9
i7hwK5NsPwxmbMdOHCoiGJyNNX0+ZMyOCLHr+aGVHYbpvCvzs6JWPmSIvh6Jmag8
DsgG2z9FppKgxh8AVpcwJXdPp29BVbUFDHmLMTqVBU329Pik9rStBlfWh0btM0L+
AQnWyODpyb279MVaZmPSWeUWjcXHaLULbDAoTEtLVnswWnhLgjWlC3YaxYaW7TeK
mIVNsR6U/V1kEtxNT1qBw/Fvdmh+ydJxBfyfRNRIWTlrtqo1HB6+tXaAg+9NZlO4
Sjc5kd10wfRDsLlr17OmxQ3z7Yd+tF83NTSNUVWerhs3HS7hwvo1CnXuLqPaYmEU
EzB91DrxJb+lWEbzG/xyr2yXZuPCOK0vYnjmHc01ctX5i/5UUdDxto/Bqo+dhDyK
AGs/VZ4zQLekxNDifOIlRPC0/fH7iWhiss6mxbUWodtkTa0/35Y9KxHWhLHQuha4
Rd1qdlQxsJMIDuaP6HbYesuku/i7lpBufatlVhW4YX2NkmYBS0w8fiN0nMM0KQom
mcudhdNFAHr7hGiSRRZ6G4hEPKcuMjomtlWjezrxD1Dp/U8WvHuaCgWRFIgVnjgZ
BQqfMRcQhOG97ucsLyzUajMlHx5MI6faWFceDrHON/DvEzHFPQ3G0rcGB/UT0tj/
sno/hMuGrpSRiKuLpb8KzNzEoiRy8uN4nPfURByu3z9WUBTDouSX2HfsA1MuUVTW
oBPuv/xDo9K0X0NTswceCfbIdZG38igtJWlx0y4nO2SE0xzSHqgeepVixHdXwn5U
9vD6YlcYvesn4RpYlDE/gF/1x6le1TPSe0ozwTJ2ATSA2814AwNy81b3X5QdyCpC
kEggmnPsM0+thfgtzVVnckc+OTNEdcFshAoF77rA52AMoHlUC1jDpunQmVABtYr+
osUTh/LEhfosb74bxdDjJ3C9bmsug0/RWUsiM7pxd8mlKLVxX+bo5H8pDmU0P4Tq
SoRdO/cDfdTZHYY0JfQ2yCCnOhEM2nIgxHNB9p5iHF/cu69EiM41r9gDK600/DYl
/7I+LLDiRTGyxIvMdZTLnhIcPh3rVWVFTBvF9VDCMlK+uIx0w5JZqzEBNlr0tfrv
Ww6hXcmWvLA0W+VfqaHIMwjFK4pFUXw7EwenPliI+0+tOZuBTt/Bey1AQh8YIgwD
vKsz5m3eap26tvWhxQgJTEuxXHaPCy8L7Qxa9XmBWUiJL0JbZ8wmaTqovmWhsy1w
HuvIJOoQGbVyQoXLLCJwml0hrD1/drYoAoEFJuiZHJvcPc4hOnt5A1SKemqODnf2
5a6JxVmzV8ypT1/0w74IoyvTjNCj4VK9ZhQihSposDev8m9GmK7Utyy4UOnEryFV
N4+mD0zYxw3kbLZJHPCMihZqRqGazsaVrtlmTvThgCsOev3qnUyPYlB4eslcXDPb
Qwzg/wy2VTSpnKtPtlu8COASmAFcOXuT4cShMOT2gVBJUrcWDo85eMXmG+92Nc6N
LlqSh9XqGU7l05jJC9mh3lAlQRUnUpM/43gJMHoALbAfTieEH4nNCgjqeZ/wlEVR
Kigu5PjGbBYB4iBcYTMMifJK0FLnU2EEggtKjiGfEeZun9lbOlLPbRVMoo1KxrQl
hRpkofHXeRhLRjmTwpPTBv2PbT4pa00fptusvmcXmVReK0RwD35cMe18J4IIQX4I
ae/K8RWfbJ7HFVz7nbjZ9zqIjUy12cTVBxpkol1pIX9oBxyVmVXLmhjWfBk8tzce
KEdoTfr2huxORWdEmzDfjnr5nwVVH8lPY1vJhHtN2S+pX/O5EjqL3RzbWQi8bu/V
JMqLPOsqT/kDQndObaiK7NK5GdjUxl0Y+mg50K+xcenAZ2X8m9JJii7omC8PaQ93
5TBp48Z03BNvmFFgVAjHD9mrPp6A07DVYMygMl/7orx/90XVAjGhF6BWvlz3JPfo
RLX6y+1SKUWbfsrtqQil9sUicSLakZcGqe7lrOtvpXddL958bsGuDyfRXsse6NJp
gTfU+EYs+Gi1Hy1Ls0SY29Jcf7MfA4jIAbU878gBGhIpsI2cvS0BgCt3SYxBqc5j
7koyRJrIjCgd1cMA35KtHIiQNGCu3qKVt15OKdbpVKEVAQvki/NtME6Biy36q+nS
IEHrp9nmaSoJHsJTNo1x342gjHgrtGeALfnTSUM4duBT9FPFPqVTDLGgZoTV9uNC
98NtKYWHiS22NEPCdZ5wotzEB83CtyNRlXWBeUFiERSHbiHBm3b8aGJqWBMDZ+SO
cnjU11f+UDnGPsbbSeiaLAb58matnwZ3p9XYTUJTS1F5brJEkqRxhDl3x6keDOLT
bsSz2AAuJuiLzxVjTwO+g5VmnsY0WWBspaWOac7wGLsqQ5I1I0qHiW6sHFpqJFqf
4O10S8/IAo4w+zuHyW1rBOdQ1ONktJo9phSj0jkBspFm0W4RovvKwxm5wWXLLhvI
TeIxdYiRsZgQLuob0NCdRcdy4XfQjMJYisjMKMh0D/+Aiopgj4jSKQ3mRmfUnBxc
jVgRgJL+XuB+27LPOwsWqicoc4Np2Y9ZekOS1E1mb4u8q0g4m2WHGS/YjTD/w8pB
edJrnbNRxYwb0+oXAfKpi6Fn/yqJThIQlAXE4qudTajNQUeF0O/A2DpeFBM+p6pt
PJpsquMVh2rxIIbRu0xsyzD+3ysBz8AGJbvRCSufLWBqos0ko8IODoWxHIkGBBxu
DGT5r5ll4WvVB1E/rFpP7B0QVk18UWl9W2XfIMbnfhXJGhh9DLkUpreNzCRnPAGu
u3bedVOMGr4idOyh4c6ES6r/cS5VSucySWwRSswzGSUix+y4p4tg/aQQ1i6tY62Y
YHujKjgVsu4G7/xrieFt5xbNE+tAE6PXUR37cVbx0dUHk7sv8oodUTfTQFbtXgGS
yYZFzI4VhDFXC3UCY0DILNSO7FW3Z0oFIyxwgYcXYQdzS3bQJ/7FhUIfxCAYva9T
7QoTD7gU5oi72bNW97x0JNCiwtj5Lih6oLZnf6N925D0WHGIueptDUyV2zImwHqb
xs9iBSia9ft7Hu57CIKovq87yzS3VBLKoCcr7G/jLaVFk8QnM/7eHlqaENUpaXZq
pYEBRidR/Z458SDOUKW0jY0fCQLEonamwJBCR3r2L0vTqq3z9cj8VeAEoOpVSrVz
CJh00wYz6NERYC66BkIWib1ahLoPcpbopV3SdqrXt8Y+q78722mbxDLVcXFpZOkN
gBnuKQmUaFqAeaN1fsoqbvrf5qQXeOd7+A/NO6Quv/JFbWzePGEux7JsGZS+8ISI
P0FaofeSsZt5l+RxRC06qiOEPlFz0y8rwVLWVYMMUXY8p+/+npWGN1nLlVhBB4iR
h/47noqb5vYXBlJv/7cRKH7NvF9MVn5MZ0gtO21ALYJ8GtcwPGU4GmugQPkEWj3b
pAP2DnElvvuNGzoLh1BPdR0YUQiwaJafLcOf4VDjkrxs4djYHj8nk6TGUqPjT0jY
OZHsgfHUtkkXC8kG1NuPfcitw2mQGSwhdkr4K9XVaVhZECNfOTFClUhMyx8zMv1x
U8eW7c2RmFxNkeQ2LWfpPwifTSZWe1XC+VQ4kyehoeNbf8hkg0PyNL26QKcfrPCk
TvEUTLpBsbyS0JZDZVrpS0UVrQqeM1egJKUUAhy4/1nwG8+pzDPMrUCql4/hOup4
fALOhcnvkASaKGVcFJQ2KwmcrdMykmPoG6M9PpgaCD/dWHrOFEXiqd6ZipKzVwcA
4K3CxPvN6MNjqJn98kXcjsR5Wfxi6URFs2dowXO8tdMXyVEadiwKq11zI7t1HeS3
oHqAQS2T0dkrTZaVYKf4XHFzFQZphYRPlZYCNE29ikaWiTtGY0nOESVRECBGGkiV
/BEn613rrzv2n+rt7+QhguZnQp0RMadRkAMSC2bYHFadjCgQm4SwOvC6jKx2u4wA
l3CYLn1ZfYe7bPymWEDqkIShvFyY5hICXOTNWrrxavIpqGSQTFackOTJ8/YscEiN
z5iVsjEIeHHM0FJ4PIlj1VYt23t2Esr418/02LqL3x7OYosVPOK2AYXQCCoKJH69
o74zzm5BlNu46JgDzBBYRcmxYFy6HxpYOZRblVPPhI3LWHSX7Vb+i2xDosCZWm8U
tTOqFeNc+cUCzq+nourooWNUDvk9dVMNX6QbQlSO+eb06tuLZar9/uxmHGFeG13+
2UG9pTrXXr4sTthaVr6Hwy3jeuCHM/ar484k/UUGOjC/v0zhzqWpKA5sitYjNFB0
CCWVYHtbXHqK0s5/0VH59Z1amMQ49xBFq+lkngdeKDGeF8XAnGYQnF4/OCfVQvaY
1NnfpGD8+oyOdoOHNTotFL0SDsm2Lu/Z50kiIjtbDHdhabjnUmmuCcbjAPbvxjT8
In15Jj4wJduZSl0LvzPdA2MY59eHJNXPiB5HfnfcGqUS5pcf3byjsNdNx6HG11v2
7vRvY+hVRQ8yCXC7V94atOZiD5qP+TsB260qYGuP4R5it3FRANpllF4wbVcnk7fa
IWsYGCRL94W13OyOWhcIJtvupeiFbi4G4LOkfwgWf13D1WmPYQnp1c9pmT/YBGcR
VRyD7GGdMz8GJMnmX97079tFkCD+P9khoDCAVI1OazezJ+3dJhbCJgoN3zO7GTKG
6BMEIbVSmyUyAK1bxZBTYQdnnnsoDBYLXRuyVldB98+oJ9ybJvaI/F3JPuXHUTI5
78U5WnXnxp2ucjv8XDY1bSVQ72qLYExQqfAsr4FkFm9bCJy0FaV/VggsH8EJrbbL
Q4jKpcKeqPsNKeIdfzI0xcS4T3fk9edYFUI0kB8chbNz4k7Cb2eTOfz+K8zIMFVB
3o2VD7EndbZGcJXPKyHQUYVGusWoYGu1+LicveCBIuM2W1wQx9vVNFA+cIdYRDbm
tTzp7cOf1046+vNOASwN7x4fmYv8/0UphKvAVjx+SK/xVqkrzetwZrqFoswFH5j4
q96yW3cYckd7RGtEcBdFCucfoqz5zXKOSBjOfCSMTxs88zyFU83eFgVT6T4Y6Xa2
u4bWpZk9Mwr6uZ7fNWIIEKECmLulq3H1cx8XB1L7g7AvVpdvWmHfApkQ1LiUsLaS
/kzMLKGi38DINLpAUlpTj8ZssOlmPEdGcKTeILa2/sL0Dz39VuQoQdfCIRQt1p9+
KXYRSBfH/e+i6jXSsuGDIrpGFNGGnxSshY57YDCPEuyd0M/RPuCOJOC+U2cVwoqR
ImsQTLBGffBTvPcheOUDWVsZY4Xaqg5zwdiVRhukHQKiy3kuGY0CL9m9K/hYk3ly
b9zaOlLr8PbcAC+7s9q8FXGY193nSDRLgyxZuPvY0DiKp9sWahk2zvWDEdh74rO9
TLJQ2uzMGVcY750PVTH3ZapLOlpN7m2TBAb5/xIvMtMt8tEltimpe1c7lEpXgPZ1
wSlqg5huT+tJeqAyYhtXEyG7AAdggt0TK8SUVJPE1B5PO0VKC07gKjcmPZegh2Vp
aXcGc4aIri8pLsWdPFZOWoatmfFRQXsTWXmO0WPcKHJj6irO1NUWBhyRjoriOoYZ
csvGTwHebEoxzK3CmeVWbzgwBfHl+pyhTsIHrGiif9v6HeNj8paxoOoIezyEPh0e
4obE4pSyfijogibYXSuZBOSij9PbJj7a2zBvyIH08Y0ErIyVURKx3YpgT+wb8+Wn
TFsvl6pZrv5rY100L+AfPH289xhglnPtVuNWK46KTiEIzEGjvURytH/OVtklOq7V
bIz8+bn/UghtL5ZGYTDWC1g8bOJBDh3JoviiHZS8aLRzEjqnxmCcxK5jN8X+E7gF
IaE88LlcTabU+C3+ERqaNBRKc3cVHBdwrEid1b+daoof3yNaLVdLkPO1Fv05SRIS
3HDwJzthkiIBEKayazN2n1ogteIHV/wkR+SuZX4ualWziV1dRONzmVPVvsWISYg7
+NRdrOxtyqXO8FBxXf3+ejnoFoKfgtV7IqncpNGLTemWzpxYhdqsE1rm8Z8ZcyxW
zmiITqYpdrXF467TJjtDMns01noEpJfqq1Z1MBPyqCL6el0yzdWRmKBVyWJP4I2N
XIdXbi1t/5AOV5FDbfV0OBdSfuus8mb7TauWjq8rDkvfusDy+KLyt9U4+4sBT/jL
eM9vTXH++aFi9qLEWGpC9M/Y6UA3AAx7DfidtoLN2N6F97oq9YTZPRdK4wIREzgs
HvEvajhnS/OdQ38NNlkJf9FSkJWmW3cmzWqlNgNOOebwPZ2Y7IE9U5wpM3bIKZz1
rAvWMLBi81UYtLH/vAzLjZh+UqciD+qjZ+lEV7x1INoyYabvaCir2HJhuv7ijvV4
w2XdMb8fgHhFI9BORKsltq+1MY8X8VrfFGRgsMci5AynVcaI2M48ky7HP12BOVfH
PDV2KwqLUKSLJfKd8jptljHXXtQ+W15gi8OxKCcE8T715YdfMUSxRe6Iwsl8N9WH
eQynsqMH+bIORMSbFCdilPVtbhZEXvYOj3IA6Tgqt4236KIf6vaJ/J+VSiuJRo5K
qKyEdyAFsm4XRl8WFNDQngjV4C++bPJsUaNLTuUA2jdx8XUfS0If/uas/2eksFVM
las3MD6qIcXydEzDdp5QWxDJuvElOPC0BVDIochME6bDxcSNttj5Bw059RNCd1UE
Z9Kho2ejXnSrmfshLo/6smvl1mzkOMnFlhV2CQv84kQw05sVJQR0HBJpafL47bkS
oov8+oGqu6ph83J31toEkNFARiv2ZOG7GjkPg+slXtwKW1JT1+R+sScpgydZPnkx
9W1bmHCZ88XUZzT+kXooy1SIHmA2OJFgNxewpzUYDHfKkWeL77MlhO7qaDxahIf6
zlEph1zfqQ/asXf44GLt/sU7z35vas9vMQ0uvGTo5pWh6PJ2aGSZ/QZzh4IAWDQu
WkhwouS/jUP/bD63FdVFLXvX5rGmEcKuXJU5XrerwNbBpCTgj9hGjcVW3aCtZMbK
Xnuw0dik90Lg9I9rPd0YfOtDZfzMesw5aWbIQ5vf4/OLKwwNKQQtPUA7ZSCm0v5j
QQjJgeFN5qw4tVW+C0NgJ7QqF9RYYMeXi7e/yAeaE5kt/qCIJWJOdfJP3/9LdPU3
QDIKudJm35F43fVLysFugcTd3Cdjsi7kdgg+1KUFn48RrvCl5KBqi1SEXTFA6tmM
q9zfBlYwbcDGfDxcVzmuTJHK2hSHPK4x1T81znBhn5fK2tHSbp4r2fVf24RlhDbs
sLA9YqDDNQavHjnTfCjozDijRI6drsAzS1ngOeZ6Bm6I6DMA0jkxyueCQelI6GWW
V7v3YKeDYFdtZ4t1uB1W/DQw2h/GEGZFEmgHNeFHkYwlcraYc/2KpbggSwS1tUDy
XjcbsmdZfAMnka8hSsckLltwCG5GrT+W5n2zZzLcPWndSdyIetxliR7/03vO/y0b
Tp2lHte7vbFI32AVwVTMZdky6Do2MMtpQIKdqt/BeWrg7zji5T/CvyCsvuYFufal
u7+5nfT3siFy9Kc2wXnX7kmMbZoeO4x9jPl+pDX1kcoeREZ1XmIXEPjLgZPDeFnJ
cSJ9N+W41jVMyWsoJPzh1sQ2/W1DNWnVs9lQXrVd7zasEuaVNgYrS7O07pPQIgmK
l8IrvJ+BULRJnxnfkXWRh9bPo4MpAC/jRly9ZF9vM8LzUvzIWiGw9aNNta5CCc+L
BZTPdUrebIICxAh/4QeDKMqeUuhb/A5vQ3eoGzNnP1FIGhVMaCbWb87HA4/g80hY
kIiP2uDvuQW26ZVOTnPVabKWtAa/yLe3TQIxMyIHsPiVTWsFuxUBZGIAmH6n5SHT
9V3GyjGPYvXitlqSmnI7x5PN8hcik0JJcFAIwO2fTvMCVojv8yiEvlqHwXjtRWgq
sh/Y/Ks5A8S0m7lj7kYph1HN4OQi2vAygYTf0GmsO675iJ3pVmSgPF3B4NyfJMZ1
PTJcrF0QVINL+9/yxG65RSf6n7R8mocR/pPiZhoaHVSC/QW+JOaXrxhL8Ewd4kCO
FFJ/DMWk90qnf+O3d7imyUnee0j1/dKeSQKNHN+CFvg7xRy/AQAi5jIMO2XvxDRI
jl8r/KXqiEZoRIKYKevHKU1zZxF87qhOXVIzOJxyWU436pHH3hcEJatCnETJrjkK
rCGqrOjtvJSGnOniQ5CzrNpHtgAOPr8eBjaCTUb6nU4i5GgfK6ki5vV+fiEPUxzC
gsHoyzPKaU2HHXm33gw2Jbk8Rig5iKVKpha5c/PXvOPJk00Grjo8/Dld+cT0UW0l
chV8y7VMikJLTzj66sRp2qs5QopitaSsWXGixQTTLM67egq5+d09wE7Nkc71xlu8
IFCltG5fHrRlJGEJVZ7yd8q1dZ7aX8yDZCcpC8SYsw4CIg7WZG1LH0kA6QmN/Dqh
0iZb8//VR3CGAO0wKqu0IXBMYUfuthJ/3rmHsEIANyKQ5NZ9YKvimZ93wDsy/FE2
BhZAdo6qWwS+ZpO5UkvF4YM1GOwlurixJcFNjw0aGOmiOQUZjPwMLKNKipE1c2WK
9otTSPGSdPiOiGMWouq1CARGdnK1YXaQBBmizSw0qBWv8jSsWinvuqjYDiTMmJdK
13lQMuXqbKo/vGc+qtNx7TvT0RjoRkxiJJZ3wVpQpCEWIwZUZ7xM9e6+m/ncKnPy
wTYYMb1DKpF+LfUQPfOrAfGow+8/aTwjbxeU5I553j4zSvUIDwlNW6y9bOfQr5Fs
gM9y6fVpYsb/jDrkT44NNgacce5gT2RZ2/Z3EI5FI0fctFpfErQDR2+6IRrIiUab
bn8QN80M8xgPnU63Nha873lbejCm+Iw2RfBsF+M2gk4druoTbRm/w/Ag6NqGi7Vd
SyAv0hJA7SMzwIXG/7cFoeGj9HhZjJr4WpBUfqzkC+bX2seVzRvUo9zfd/zpv1bj
bYS/GiQ+2Fmc6Eb65cLZbxknzUQ7nu7OH4Ncq+Tf32fadMo8KkqMg1mwmE0jMPVs
2xOO/PECYKDsj/GxRGJyleU8CKndVJqgZwdAOakMI1aaOKfwQ62WiB0vonBB1hZr
/bdi4cX/wPcrKweexcQyvq3heg4QOo3nUJsc6+8WFvyWiXpd1k+JyPRTl93QwysW
nWTN/tjkRpGRFEFTYn38vU5dgfj5GXOJGdEERuP7j2acD+Nlo4tU/6CkNjRl/xPA
CUHE8uBcOkTF9MR97ST4IzB+sZM3VP5pqEargpMmY6zcb6RjuaYdEXZZfGl18Wb3
Tiu2cTlr/Gjtm71ujjn9rExJljHZUIDydGQUxLpFTPwP17ceNn/qQJzCtfLLL8Vr
TABDuMjOEmrYjFi1dhF99tiTHrXAqx4LQCRY9vCWZFs3/r7xojgQGi/PQekZJwDl
XFA2/QiE/rUcUpQwYgtM+64XqzJfhb6mOe+wg2uR5zsNMOaUic50iIFg99IeZgL/
KASGGilHAyHXMTemaqDQAfyPn0UuJDbNPPiu0Xzfu2eZ+gCORkxSBZwMyqsuQRGo
VnLWmUKMMxbV6viEbZs8tD+uC18y16i6zZV30SNAgBns6oFkNvQ1gYx/GsFdWbW9
FKI1G7mgyPvuKZ/Hu/pd75Ktbqk6BCuSyA06sOk5rmtUkQsHJDmE4fwinmKzJwNc
8C8uX2lH1FGBxF+zvOm6NE9j0EHqqizMipgmS/lyY5qRe6CLgbFU1w+wdzHqv03V
q32JacpBotTEO2VuIIzg8fcB7rgay5S/FR6yuAQaejIt41tHW9NTdoM2WYUWafyl
j/IQHIRik7VMbaAsb3uxmBjcsYQZgNkRYkCo9jgL8jbRYawIRj0zFaGPvAyOg83J
r59lOkPfFZP3bKdbsGlHO005TwAnai3SBWaDOGvteEIQfECujwfQ5kpAXL25fG0g
tGf427N49/0T5m9w19dpRJ0fmgVEKUc/ibnoCpO58rl7mwrqVFMyMuG2WUJ9CY0K
j0eFiLPsG2e4SUFqgVqZliOtmUXBh76yPtSEnoVLedJv88TiL9lNTNBRHkUM0v0F
xDw/Oa2MvUUrbmn6PiVD1e31ySucI9JW/dH2YIMfBHOrVnSdq2VtTJ7fTtw4npJ+
BGd5EkYQeRfWXMqIoikjMs9wWXAW4UI1MRsuoyw+MNhnIegYGR9mXNdXnuU5ZJb+
Gm4i48nex8anSqR29bjJjzYGVu5BYp+FkzPi1c1BDCS+EOo5jEO49AGW1BQB5ljk
X6R4nX3KdbFfo8Br9fqcu7TaFoizR9AQuPsEekTkgP52xLAlRisOLyA68gPd2oVY
j+qftttib72gNfKgXuy57uj8R6pNZDaPZW/4ZRhbZEUG9hwBolhGBBnAgXVMQQjf
glUsdzEJwj69u1gLhr3VqDCJPcLEPe6mA2fafgePBAHZo1JLDf7xIKKwdINncczL
HMXxV/WROksZcweB9IxSr0ybb1z5jIts/KIBOpwTeWYAAj2UEJsIJ35k06YQe/dg
ZVOXYCKNPfKJV1B+BXyfaxm/C237t+24V2LuE0eqPGQBLDNlpHjoofGB55+EmbPl
Y5T50jqxPYmgntcAkWP8OxK/l1UvUvxSCep6A+Q3tvF1oHXz0bLbp2HMSozhwsZz
QXvZ3Arvb7eeZmnchZr3QDnmUsUsN6QATMoKiCp+0NxR8Kr48QO8gCQrbUrqygF0
xa4kMT11JuDqEsHJz8p1G+XF++m4NMwr9e+0ys7Jk2PaEcUjG6sDXQ44MAC0OGRa
rRdJBX16c+stsnjM8qE46sxDbdssuZI6HmlgbTuS5Q4ny/An35q/C5phrJzOFM4A
SyfDQrxbnM1D27ryfQ3ZgMQiSRFDmyK8Urhpq052Fp5fZ9AJ5oGsKOek4eDMKv0a
ZTZj+slT1hTWccaJES27l7pVCbmjwhlXE233XyYiOKmCvA6GJKU0fGwjVLTa0oLf
EAGcKkdGJyo7jysaCd6+KBsRx++NFurDvwbf71iqP7OsqOmzMPrf0b618GScjh64
l12CtnuQZAQrzkFhqTGpsw2ikTpCa+MtG/bVekNl9hqUpUrWjwCLHSUkbch4LNY9
+Rqi/W/yB31AHbbwJfO9xhu47EEk0AkEs151GUfAsZas3Lx9bbNJUjaCIPj6QN/8
YDsDOc6UZwQPaG7wuHQg1EiwFX7tCbZp5GIt851NJJptWK2XEs2VsdzadKayZf55
Nf7PAcd/80PD+MnYOZb+Lz5uZEukNtvNNjDC2PTTevLzxEK6gUcGGwyxcZ3JCRu2
UlcNy0ZNrVaiu4Mbn14DihJaUUeuvFX9Hk6IJvn18iE8TZ9grb5eRFDCPdaNCQDH
7T6HxWwuQuuPkHL3imuF7SA2ZHNH9oseehK3aP/iWbys4fIB4qjcoanfoi40In4s
ZL3hwVvwDAkevniApt7UhPO2VLZfTA2ZGRjmfO29pk9As6k6+kNZ1YPhZtM9jg08
esW1J0f8oxfPUUKvvfdgSiBS7EZQRL70zcvEDv5AZ2exOAhklWlNQ1n+LF+XBpuv
oFgLd70zVxQ3F1HsgAgaCnOuor46sX6xs4dmniu1NPYvYYtsoM8cYDygqqpA4CU2
QYhW5yEqQAhkzSSMBdxItpB/3l3PiO9NGJU9muB5gr3g8wZqVALpcE2Zjy5pKvgf
aUaHdK6dkk4O95rv0++iYoxnZkvWBWNVUTTny9+0lWds1Y+Zs6NingtI6McMsEyn
Giz6gdIbn5kAS0dWkwvXlYLo6Yb64jbgd17eiJ0fIscJdu+s5fLOS9k45wdvwjRy
NtRuEqFC1OvRPUhaBB8kysdVQfWt3KxTia69sg9UV/ssBYYAPPLZ6DD4s+HeNmA6
WBxlEOnJ5nCsk/uojXiDPk+atMSnAo5sUJv/G9UqWXJ9fBXZNdCY5nhrCsRnNeNX
dAR+aRAWW0FkWkgdXmmypv9RM+Gb+irkWOc1K7vWjnS6zzVuFkFyXv79Up9igks2
BnOWw98gYl0KsZEx0/sg3cLRl+AHSKGQY0DS/zcOQ6z4dj1sK+wjm8pe/L4LOKWj
VkJ77aWbiqmxlJMayUryIWqgI3RRKR+yPArdjNWNwC+pqrVhtlE4MLR7UdjzumjB
XDEogLe45X3vtx8V+z2uNhlAaDc6NZZPXLYSIWL6LLDKbIxDUJWvOeZLoLdDOY7v
BSSf9Dj/u68TceQU3aLlzRT8r/c2h5BDPGVia68YG3v0X7i9X6NE4Y2czDhSWhnJ
aQb4eHusY+tur/k3q9PdklG5TEBqiJHRQjoxcZ2B69sJJCkOC9GDwVVPCt9Fnrrj
09pzmi+rIbdbBiTsaDSHOW4Chp3tk72JCXQvzuaaTSlSJgomqtyk9i2DdnPjugYV
cYiu5Ev/kjtYRHD3PNQTi3s4mRWhfeJHccdi549zTepiqwRyyPxu5r0/PpNDTpVf
ECDRJpym4eHLX8PC4SLIZugEYK+5XZUCEbeuRc8GcyMxE9VWJeuXbiX5/o3syCdg
v9HJdx69DbI0srRv4mhLCGidtFohSZuQ/ZwjRqwGgKj+gAEnMjJ7BT5WOcOjZX5q
K/VWtiuhPlastPPagG5HR9lLrY5q7aesDu49piaXX7GU8XP//nQhcp3Ukt4bJSE3
0Uyqk+QCj5D/KsWEo05Ke/yNMK5HRoDiVHB/GtO8rL8q0fK8NyN/tSp9nf3+ntkq
zuYMHR3ws7mIP6vviP+IFth6K+aUZAH7ji5dqbcbqjt9mzM3kDiw3LocmhSNwpKe
eLMmqMNdcFriQ1IJrtyH0RyprQg4arePHcMgKBDMyKfdnT+RbjnBikmoYkV1+ruU
ORlBqH8SokMJGbwCmn2BQdIOdVjXRiu6q5DFjrZqvUaX039muWrrl12nGtVPoN9n
WGCrJPObJCkr5h4BlCqnMCPjXl1pgsLg93843Biq3ypdAA0mlvRHbLbyj67gK8XA
WXRE8rvIGLoAq7IuFLb1gMYqkstfUcNhODyiJOOjnOIXyLyZopme5hs4dpNVy+3X
9gYxb/b46WEPxGaTScChiRlirtG0QKb5YGE+iVzUvyuNyWwXoJnR8X7GgPIVserT
VD38RGL9Sue2wV7AOQXMFlcHwq7NpWLH3i2WaEVzqDRfQh36T9S4VB7JNQ8lzsUm
jyjFN9kb4lDmnCFkbRSj+fkaHAmpgikC1zJy4kQ3ovDzqzi8VDfj1z4zN7xgvtby
MHruFtJ3MnQ6ldI/zCebqtMELGPPjolQryTdocP1eexuslIALViIx0l8zueEP6jo
zJXXi8wHf7dPNQlduJsGe15LJ6Hvt2e/Bu1QE35pbPxQan7fTLK9mC+afSWWBNxO
bqMzJAR38t0UWk6oDKnWUmZgHnU54eIvFlu6vs20uYK7o2qVrcGPIG/pfZvBNq4o
X2ifIqOsLYO+FXV5Lm1zlaZugJo9wrMalenkXI1F6xWSFK+npDY0rMgBU2R8AXrM
rrwSOIb6rojebarDAyvWdEvsX1bYA5ns4Y+ubp7VXVH8n6sMXY5hOHnXUFfLaG0N
/WLY1D+WjQS9t7h5GXFfAoG1YWxdPh1EAc/c002eqnqbn7WpkfxK7JXIge2Lrl+z
abDPplzO4itGIdVE317t1E9gaxd6IyQ2dlFxw67R0S/8JDcHbBWepsFQ2wAx9lTD
+YtfOioou470q08Y7lEwnIaziJPcuXnfx2XvADEubFvJXe5oqCG9cHuc4wBz21jH
Ikrs2dnJLwWk/mOwZVmVOFAt4LHyLtiep+0x2eKdpgoirGWyydvwl7/C2s/Tw9dc
S5xglBJQrDkcxCK03E9+VcUGqMVPFwJ9F6GXxGZmJ4omzGhEB5WYmHJPg5QUrZUb
T/GgnqbVQZvl52cQFZyPORxOSWkgHnW7GdeTc3MXRM/K691PhTLZxADspiDtM6jz
NoMAUrEMzgr6g+TJNwWjhc0OOS4Oqe7iVPf4gIJWX/jwEveXb3YAiGOJG7Tk5Eex
XddvBHPxXEhiRugeuagEHxOtFX9Itk09PcoPtl7A7RI2v8xvgVmZbVdUicx4KT6H
HvuvPB4jYuG4WSW8+dSSgMlaNBOa2Y8rhwSDoR2FYgBfL3kPcSl5GF+t7CBKiN86
w8ctX7Idyqtmjxa8u3loH0VILE8GL0sZiyEZXFEf4ohBAuIP6ZU+gFkvlkZals+e
B4W/cayXV4qiiy5SaHdunsZ0W1Z1uQXkxbJOUO/FOMo8yof5z6m/jgMCvFc+FxYj
HivOx/Y5aBaMB3wNR8OQPLPvEtsZUQmSu1vboKR6IhduqtJnEwZD0ZbsX60Xgzv8
aTp5kgjbWJoxhq02+l9+swdv83YlpBZRhqK1pQ2+D+/PDDghTIuT1noXIDolLTYo
eiTZWpCuxSGf+YsRO8pX5cW1Klhhl9aNH7I0tHrb2ONY8ik2wPV2WgoCLTsVpMmA
MPe/ktUyNogh1aunB22OZfBWxZjGNPUQ/BC3wojD8oECVsFEqGLUSyuB+PCWoAZi
71IvbvGTDQfZPJdZmsV3T9OFRvzIsQcatVzi5bKTb2f7WyC3YZFPjruVPB5P72Ez
SJZo6V9u5mBNNtF12JbbiegaBKR1Hskd/pyNhSBCIELu9ZdSiNEowt3NImwf3d/K
w0WOlVq85f0wVmKTqrOhAas9S8SWED9L/LohpI5ms+NCETrGNkljRPOD8JiEn78P
yhlfqllxpTbf/FvWJ+x3w2SHE5EC0cERp32NHCNfkRd/c8QsTe8U4BLMM0uBny90
LWy24C4Y+bKeQVtDbfzWaSi1plEd0jjCpbbAM9LFrtlyQiAWQytRuJVNi68LikPC
5STzexHV3rvVLF6IOJPWD6J9m0yw8DZHH2XX8as08AaLyAO7jgADnkPVc6uec2Kh
Qny33VY1W7k6XkntY0aECyHUzpmIjuO/UAaqOGfe1sCnx41ADNXsxqbIXRRek7Zn
qfSkp8/WGNGTv048ID/VT0syvjqyk0ewlb+m1Spq0rBNTmYmN+oX/fFGFj6OEMt1
QMXPjITcO1FhTyQYZs6se1+msOCBasQlBLSEyP1FpyhJ3gGvQBUzkEmmMY//smxh
SnmEFSVP6B1uvg9SRxPcb9+wojc2jMcn70cXby7rjNU6vX/u3hW1S0t6wEyYEZYg
nFoUbAvkt8z+I8KilFBp35G81968ErxnFr2kvPj+8ZmnnRSQ7tSlrbwMjyncxxW1
qV8pHPOsAJTtNX5bYVCpKmNytvqzEQ+yEiQ0t671lrq2XJKr5Y5oIHcUOiPGrqOp
o5wPbbb5JlDCkr99DoTbq85OH5LOrOD1weG+3sL5e5onk9+3lxTsc+QCGmZ1HAH4
cLn6fd00n5/TTB6oBX9FkK55JAcbeEZ6xms5HHcs//f1ErlgS1Rpdw8YEOj5XSPC
JwTWRna+ZPljGPWBdfufhNiwl7CYYVz+0eB7+g5Pv8cClPq/wZ8blCzwAgy8kFG2
ySy+g0LtHdqt6B3PlSfylkMPBxDSoW6VigE56H2UWrRq4rQ5ERRjejfnxzQHptlp
pb/RF3bXj3v0wbvSeGEI/Oqvqol4vF5XbzKd3nK0Zx/n+0Dk4iBqgIFkV/wDAz42
pOfHFAJ51oV2ogluyOHk2pmuarNLA4rHt2rS1o1WNN+UR1kqMstSqvEGcPL1FLFw
NSGlrNYzu3ITdkcZ95qwz26AA9MxVsAoRnaYosZxbf/M3OnYDtcSovaPMnM5m1cm
LyJj2fzX5QseJItm/o14imcqqMj8p3a/bwfQKOd2dH/yBRFZdZd2FLljdXjxywOE
N1TFThVUEfVGD86qB+b39YEipcujVhVcR1NjaANjBeLBHuXCkz7QUPtvfLgNHU75
eyDSyvVuRNGH/HI0P1HoYQcFXLpSj5hY6d/PfhDQrrvxq8AhMwyhO0441n5ANgA6
SvAZ2UoePPt56ncFPiyEY34pXN1P7BKwMbf5UrEsvzNj45wUcogn3oDVq22hUhDN
n0s+Ar29we3UjoFrTGvN1/Wzl8hwH9viBjI+bUuG+VQYFxT2WL+zdNTMQreJjzuN
WMma/Eopm34wFvxPDsQQoC/pJU3TbbP5tJX5UsQTENzpNGLUTXq3EzEK1uknUkOc
5GD+59+MoZMJGMnO0pIGvcIRIeCfuD2cLZQCd0alIuDzfQj/GvIg/lRPTotQ8F/W
ipwKGScx+YPVvPrp36Fu//nxli0CVMEqglBV7ja5gEAB5+ztJuUxrk+LRystbe3P
QFh50Am3Fb8hs/rBtbz1epWE9B7S/QtPClmKttXJWkFdk1KqD7DzPgM2er1DB1WG
IRu/WnitF8pkmi2qyhXHtKKIIRx4XcSx3qnen92GVb+iZ6PEfCtbjKWGTU7NhZ6Q
tPPbICTthjDVrjnNuwb531vazjheDw7wvK0RTHxV8IyyzPAP3Ej1laq9tbgUxeFL
rp4MHTPhyYKltCPpSHBuzBroG63MIcMjzbBdFIzFzZrnUi57YALPJFECW/sFqGzm
4VCn8NYM27lxKoHUFBF1iUQnPZuDnQucZX+N4IeosZAsu3midDVBB7VTLBtSoXvy
Y3DARF7lxMA8SUKiRsmecF/0PfyOdScVwI+C/au5fRHsYNdgRTwMICjC7slhLqhP
e/my2yveX3GE3wpT6DlQsE2fPnAPxK4Q+vtUkoTdWRn0cxQav+6ieuJ2mwKGpwFR
X5JsKCBQkHdjQyDsXN1lZRrPqRYzNMUbBQ7d8LC921tCJZj0zChUReImv89SYJ6H
wwML3ZXd5+rsF600TOW8vyyi41gHBevnorWOL1xr2EZNM0ruG+pQ8iFinPS0UcOt
i95iL0NixLt9AX5GhNAASwsmsAsD+r22/sxaSyknvn6yir/TwDMAxrFzJ5mBjoMS
g/I+sdyb4LUIbkUp/cGZlT00sOEfzULCedVx7y1yA8KGC15nAr7QzkBsVbaEPbL6
WlNH2qb2kkG0BqIdNEHif9/ORJcVU7rOgQtSjQTmW6xwYx37gXTDas9C1cytM9Nd
os5xh2pjJdUbyge12824rg8m9C2Rxc483BDC9k9wQftC+L3Ehzx42CXSrQmjwlEQ
3baoXhiiqgOZHbzZYRmlG0nnXxwM+GcDCBglxOJhYEXuiNJiczjhHYCKJ197pGkf
OHwOhYaFAAWg4jYKg279OqJrbc0fueZISQ4nLgSRXN2IDDpj7w2i63JqbuvCJcm3
2Ocobyf+MVOsRWeOTfelKnp/nS9u4+6D9qwILDBYl5urjdXzebD2BeY0q8qad4LK
+sUchBZMiiDTmAtu/NO1lbS1meGuqixYyyDkDJD/R3/0WlTh9J7LMalzL7irpgJK
/2BdEK7GwrF9Vplyv5knn2HG4Ur/WSMRMeCNMkviDZp7AtLsVI8vQr+ve4pn2ZeN
fRLa2FOqfFTlwxeZijBckBuQWL8YJJeZALcaUhNxhEtiBIs2l8KIAD4JIUw+bIWl
xP15hAOps7n1QdfKG5tM79YIqlsQNlLVxHopYqZj7rzLDlioduyZ3jnJYvaRGeC/
itjtbCMjKz4ndPljgCX+MccIPfEpje+l+WOxr0cbQPJ7V5lfmdn6EVJH3UB6LD35
+PR2j+Qs9Fq05mEKvlBHMi5k4SrCm4J8XOjqP+CrZSWTbKgulmw/SWEvJ5/8bmsP
lEF4vMdnxviRDyuDG4DSNq05U5qD5zM5Axp9MtEnJzAGX82wMtDmlJXC2i73igFM
QhsEdFrsIld77+2ySeTAgVt5AmF4pEU3dJEyXFhfBqAYQ6fGvuZ/XwZxRYnZcw3V
0IhG08U9+bYlXGCNm0iw5/ULjG1pLwk+2l8Z5FAQwGkfsKzru+POcvH3sZnwUH51
Zp6FkuVEvj38g0JAdqtK1Lt767YuqYofzQTnqJAhl2A4HDz83wit24vHrjP8s4mm
0AVbvr918o6La5I+7ek7NnL0sULvKRZ2omZPZKfb/FahILmnbxsxUDxrUH/60+Lo
J7bcSPLpQUGnWc9RQ5n7N5kaYbG3P5FA+GSKPAlvkQr4ZfDua2a01k1yc9358w/t
XfleAfcfvnpDZtYHDN3aCCC5A+XcI1aD4/KEfhZf0OahQ2EU21S1wGTPPJTfGERo
tJq7I8oCRg4FKe6jo+l/KXQlrobLmt2huxck8xee0SnrPOyWypmWPzox53OihHjb
IDQDr58CFYuzBm+ASE66GuDIcxfaxcLAdkD3L6F1mE/3IJLfNQGHxiSa1+utJE0r
lU4sA6YccXXMspAKacPpXFjqLhi9D2iEEJkj9qMxfuDSCmKf0tWpD1d+OZNZEQL0
bhLstCBBnEA05jfC33/ElC4sZ59EHIpMmVJinrdCyZe6KYM2h3fgFRbBZ2vZFRRh
DVDgzrRNm9Hv8TYYL4M9m5WY9PIxlxpGe5HOK6c1Jx9o2Wx/HHWDJMgDxZAVuJ5B
anubHEu518vAthQViQKDUyze5VZ3V4pHuSp9zN4ohcHL6g3fbTdKvqiRwp0h+Igo
pkM23g9stXGSnfGbmX5edqeVOY7rzqTVZf+rfO8o7+gBCHl4WDfD9gdqv/nAhVTR
Pi85/YmncnM0bs7od13vLB7sqDNIQRY8T2ZKopa2DBcO87/JSaBTd/JSgtkJEOdn
vs6Z/+uMRTIVD57YsDFIAfovbqZB4SHEuYXxGMJVT7VHARUMuwsuJ4gWzK0ruUQ5
xV6OLOikmsfEM83I8xXmocm1v24LbiCoWTLZDHoVeEn9X0sv+n7neTYF6/Q/zFjN
MPo7xoZEG6OXigmuVgDqydnyFsJxyA4CI9+DPo67yht/ylyO8BICdmU1Qy2ytyg2
7jQ/wCoLNkBu9g/Ay+tNmzF549MiZ28cWRE7I4sgWerMjJUbMDpI5vMgVSz9rfcA
n7bYwc1rlzF7Skq9C3Sfg4BNbgU7/omIow2CJPwfim57VLFAeyn2TpFkRmB0CGrN
y4ANfV/SbcPUNpyEf287UjWrBvTMaucoeYAD/B3vEFSp4jAYRylC4kGRjuBEpYiH
a93Bd/ofIhQ1BZKaJ5W3CRHFhFx2YL8cLDUhuVowPwK1pAUtwzs+wW4rs46mL/BN
4wwdaBNFeSXyNIn3YTUiALgeOJAR0cd8kRsD0cH5VFBkQzr19JIKnsTQgHM1kBVb
MK7c6Qht2UzxlCjnGJbRiH6WrToaueCv5CxxwldptOZY5gzphYe2PvA2wWWgBHlS
p9hdZGuBerpe1HJ3BiCsMAReR6PBgOAkrLmdO0u16QjsoCYO7CHBmHFYl9dCIcvW
OYHYtAlRFcEMk4LhVtMPAn6M4UN1w67FPKeoGfPtFyuN0XY8xynD+FWXokeDF/+5
yLjEspbFgPMEsSDm9FFfAMqKUagQfEEk0WfqHjJvu3/dnTkLXzIFRPdZiHD2woBK
MkJzZr6ewbAIUwpd/Z2sL41lwYvuamoW5KAkI55A5orJcNOJFQCt/i5WSLyQvCUS
bN+eWeeK19EGZQdNJ1FJrclQ0ZzER2eYbzTfVyp8ZXws8Lq24HwhUAeH3wAzIh+L
kSv56YR/GdIp+zH+nCuJJRnZBSAi4D2IcPgXnWZAUlR4IN6SDQEvdKF75G0YGhh8
yRM3mVCK2Xwg8yU8/bLkw6kINugSWdFaYSBM2jPX/mWDu7M3BCf4oeYXAD7vdFlH
9WqbA7LLkKgH9BEz1TSW6+hkAe2PXoV6Q6oKlnQ1Ty61KNABfLWrr+sskaLMjEPj
+ZtvvK7lWwfWi6Axi89fssu4b5OYrnNBbHPL8Z84dfj5DbDVnAUsKtlsQOzImgOG
fWjkXpZRvkgJN91SgwZFbxiN7BJNJrzt1BZ6TE75qoUqvUA+9GaM8bXUaDp5sHcU
Gf04qY2LNKc7Ps+Eqw8K3SNjcx5MxMLDE/4r7a7FuWsvy3YelyAlKFk8PE8pcLys
7cTLb2t3dYxs97R/qzngUwOJR2ixHN6rtDn4T5ZmKdQBuwH71YNVVtX7eOhH3GrQ
PFOKBWTqf8zOmiy9hkQp/L53IYqN8eQg5tRFuxV9AY98LOLD//OaejB3suoHAllo
d9ym0jU7cKEkJ319/RtW8MX9OrPF79y74CnbXXqO160ChVFfgHd0tNefLTqWmv1W
yLHeDRJ9+gw8QHiDvH36tB6udKDfOrcHqxN42fXuqmkNys4gUMIWdw5ZfGKcyyCN
uofvp4lQyTDs2cmzaAVieuSqRLd6fXkLiCpGmnt2fskBj6HTbH020WwjZJrJC1Pg
YXKWx9b0XjqdMqyYNvQiDmXUTAhRvc32gv3PqQNCiz3BdYkMM2Wf2HIeYtrOWls6
sfw4sd9e8OrU0h1TcXeeZch1gcxGr+5lzlnZ3FOCa/L5RxhDJdUZfkgk6rA1raox
BbUWUwzQnqmB/BtwLa0ubakmvYcxRmv2wZFQU+9i0Mvgeree0ACQ9bwV44hkjHal
4qqUUYWQTU0BvHuwh9ouTSygHZJf1r7Zj/sXX+T/AVonSe69zCkjHwd2z6BGh5x3
lYzdKI1Cag2ZDm4MXi50xnFyp0QKvpXiCfEMblIRKu5VR3QVWH3jEzqvQkZpxSYz
LdXL/RDA2iAa0NFnweZl0l4T3ebUlftukJRs8Du6vtJkMonBO0TVYhEO/+J7mdxz
FvjofFWpBLI4/jNTAiAYhxlf1SGkTVq+YKoo+Io7q6FjPV64jahRd7B6XPqyk+IN
mEYxtenzEgul8E0leO10D6VPe68U70gKRuku1+HBRzo33rfe1eSFy8Jp8nl8KS+6
plXX0PXjbwxfGNBxJPdl9nwiA2JhUOpI/NPitW6GTIUccbcmH/wbZFx5CSut/THJ
5E81GpLPYwXGevUAsxtv36PTzYt8SiAlAf7bFN5SVZ3K515hUxvGA4VL8KJ7UGt2
Eu8hef20TVDk6WoKN18GnKyBc1uAZPikQoRxw60hAp3nyd7IWsRYvT3/fHJM98ih
yVWXFL5feuxY8rDlR7yErVbCiZkLNrv2M1R+S4qh9ugPqNY0WjGfabr9Iq3sn4HC
kh5Xp+ytIkeJvCQQVtSkkrC3YOVgxJFkZbDBTqZcVdjaHHa3M+gcRtvHpi5EmhKW
wkyACe1Gs6G/VlwES11eUqGb6qazLBFbtQovqoBNvbCWYE2qlSqzJnGwh1YdZVPh
PhHvlQUGD8KabUGiBioQyoz6/ySMUvNRfJiPAHvas23ttWxY3FWfsa3P7twalhfA
KW5RuxZr5t384C1+HPoMbtvZoikQ+Y2e1JpIT00l7KTGnTFcRtYJcOiSgDii4/gB
VcjqHhjot6Z1UrhteVJRcEFv7xh846FetaCtA9ZKWlBW4B+sKL6pet79rU4PLe8+
hnYn1xldMPmdY66rDcBxkKsdhyvLsjH3o47FYJ6g6Nnw0SBQAMJbGPBA7tGJuXxV
E2hQobILqBiYNpIzHl/mg2CaT5BpIYxFXBkhQLEmZ49oegObFzqDTQw5/MscMo4G
hOaWyEotsGa71xuaeVCPfip/SlvQKtQYBLo8Wp11P2fJG2K8F3if7Dd6Qahf08Y1
LKrkexKljuDnoodbbBeZ1Z3Ngmsh86qF7hCLsfvSU0VyuSVxwSFX7c9znh3vzRxZ
K72kl9SpDQu6/Qj6jxpF/Q8EBDqMd4UEFhLCKUKSEFpuHH40YMLDPpUQlkKOfn9Q
Atc7fUb0ivXJHVKzfahOQatMYL9+MxBKl4g0ZusFw4qi+Gf+j/MzAOHGctvBQU7q
PwXphAIloik1zeaz0CCx8NOObuvjBaJ7JRnRVvqldupaMkBJJeTBfFWgZqhOD8qe
ERCBCBjT+YcTzZB+x38VeKx7+KQ6j8GmWiLcx0qMudnin1/4AISrXR4KXa5rwMJ/
oGpELR2DaN84bxW/2N0gEv3KFYoazcyHR2et/PpCx761E53ICZDx9h4F34+hUnZS
ZLocd3m2ZYzlZT8SctaYHMy+A53XLIvyV8Dmd2FmXeonaqMTpxxyICj/rvEgUTIj
ApNZ/REJe76BX9URycNR2A++4P8Ap+W2QKwc7D1KWVUpJE8exa+ONw49sYTbZUp8
WVy4+2n2GgkIKmXywjodVo/PsWPUMQYmd4nTRbQX9L2CC28Qngkjo0ep6KWgNSCS
/khdw3FhmOS+oYFTfJlxIYpTuE5wZQh0bzq1v7DrvQM2719uCt7idd7lp9EIDghH
s5HJLzhD5FTM/yNKRldSI27V5p+W3GGk7D2cJe5qwMChaM+Z62OYYRTzxfeI9zwa
jYI+2d3yYQxIx7KnaGGhKEll20C9zCM2BZw6tbK2SsYX4EFoR8rXVOKoYNeyeq/J
NFuOewGqPChI60nQx1DWVWfhDniaBDMnjoNwJ+qSb1RKLRTft7Ce5RXL1elKOCqC
d6d9y4ZBNVQ1DE96KWaeHHBG0LkOkru+bYI2NGq0Qsw95F1nUCbNaH9YOcfkDGx3
twOhngm10P7uj38IcbJiJAnij+ePpbrKSihLeX2iosDL16pvV3leg5y0+DxzxGZ7
6YjapiQlpe/NiJ+IIEKaxptMS1uPiTEe09546W7xglFU9oCw8zoB89anWDiXft8z
m2nd9G72wfHAjNyNEiTIQKcyf1rGH+ep2RwSuBKgtfPsPtjIzL3XUfne2yt6dvX1
0eF5VZu32iZwo0u+O6d+UP8pHCOGN+9Cl+H3P0De36GmnN3HkjqOhZgWeZDKKzMF
ZQMljc1Wx1WMIvQwLgdhdWca9+lWq2/pVAoputqWETe+kzYFXNE/10TwlUGmZDV8
2WWjfn8uYVJReUUuntuiSnLNgj4AjjehA7mgnepu/WZMEjAdsOSzlW6WkiobN2tu
s7M4Kt6DPs4HlvcPglz3KAQ3BOSeCCyzJbgEiLge6S4k/UfJ1R9kG5h6ITdoh6tx
N+dXfAf4U0ZHy7K+P5WT1OuAge+7Pmx8UJNNrpaxR4Z8KWtl1WEFywFzTObLga7/
7rY0LkQDDdM66XsN8dhpsm+z7AiCqp4TJrnHU4tfC/wmS3qfgGlTlP6tz/3DEw5A
4ilA4AamHPoZpngFMTpctzP3u2yaXHHrLEHpCNrrAw2XuNLXufhFJvRJYHWQ66HS
z7OLnDJQjKobKRdCe50ndtYPNfub+gyXOjMZKgmvI2b0KWq5HLgbf4ZyBfCGtvoj
rRvWj5kWvsXowtDBSn/68hWYOgZBU7bg2AJwJThM87o+pBgU3jluLXXi83WR4nFx
PaaHCiVpUuUMhIy3JLn5Bia2DeBU4yalNZ+7jthOAFWDAdk6753J9+LzubmwcAGP
d6q5/GhvqtZJY71j26ZLorDE0Fu/U1BVdVoJtqLHvivLLJx106UFfMGRhjoO0ZBe
2LJ1ToLMdTRIxiEl0AMBTAa0lsRn38KuvI49b8VwtTKzP/KnwsBTwRYsuVwXk8bI
PeVvrGFR0/QFuKeOm0wl1iK4ZEihx5d6tfEMH24fJxa868lOYVif+7BSBTOacreR
XAAFpxiu8ZoJqE+2qRlQNNRaH1Ata6OOwc/F4dZa0fcV4psSqIyW9xLcs9ysI635
gDqLufFbj14xNPmBkWjd5axPIoLACdEYBd/vNhyzsGSI+Wbu35Dtk9Ve4j4Iuhoa
5OsO6/SVEDYHV9Xa+W92A/vwG1wNYD9hfua3mhOCu1ykF+ECdpsi/Y2kodqoHKSG
wlMKqRIt/nFP7K278GCK9f3BPambKWiI8bMDOfJGh4cyZdmuC1kvskQYnqNFBe4a
z/m0t3d+xRdv84KkFm0j9EjB81vZF9OXCxvgyHVzKGCvNlUdtxKV+1BSOugXe4ev
CNDHwA0YLBklMV1ybEZEfth0o8ZRRz+oLmwH+Uesp2HzgavRzPgOgQaNOW9MkPnz
O3ijyPrLliFYoe2QhwxLGsbhUlgFFLHu9nt4LP6b+mziy19FhWnybOrldL2DEm9B
K+eVBtz7+37QhxsyXCLgFoJneJjjQ4nirdE6JeseLHteF3nzWgyQoj2CmhbGRk3G
kGMo1Yz/LuqHEl/4E+1EdOq53xMjCm5I2xhZFY7NL/jcvKQhUq6liwLup+/6dViD
Yd6OjP6pLQJDTWxuCfU6VfcGYRxjwNQctsN1ybSxBp/CkUza/zxq8dufJoWFta3H
HgoDY4z6LXMGpo+YRs2CJPtfzTB8HgLwna0IyvUr/kHbyF5vQUnNGvXCD6BwAVFF
iVYnRRqNdJUcJ67iBXWaoE6O9cxJPi4KPVB68k41omGb2o3fQ+klr6W6eoRqQrEd
48bUYQ1bDmLTsykyrJRsI+tZCvLUhd0FJykDGvsKXPEMBM5DhkTdVZquyoGAd65k
4hBGPPzT1aNiOaD+4zRZYC5+x1QaAHxgyKGL9ay+Kk5p9MT5G+tbMa2QMTlzDtsm
QcPdYD36xOyN7yeTMnUNgGEmm4qcIkhi8w9rtxLO2I8Banzx6xAZW0JKw6nLP7pG
XjeuZuo/na1cEWIugz92tiiUiS1VCdlAjlWS9Ijvoh5DB55UnySbTzlkwTBQ9umo
0M/OuUl3byiGmQKz7nbliw6x44JmzuEdyvLfqcoHON0lOuWDSPrwwU97NOXZsbuF
/GJgKusEluGX+nzKsT/xcxsFEzepIV/gggggRyfY8t9/OgyGTFs36Ziy1vLSFcVl
/4pGSVSUf5sWZ0fUW9AFSCVFJlBHOhOiR+SDpkM0fvsp3jpTDTfLRkLs6gAgjhBm
v3eDw9mDcczF234oTdc0OIJx9IkiDzlR5zhoo+hrHVbKtmp1Hpwmjhgh81jTqeE6
t9QpjRtLbNhqBMsUjsrqPrJdVHouRQO3b13sYqMQfBNSBwIO2htOIaHGJcZRpgmY
uhG31mOaSbZ3R0yDU8o+QuyG/TSgSwCJrfTL1V76kfQS3BQggNdbbD96ePr7GxpL
nJ8lkDsrkg5/t/nAFnlJTXy2oflsUWKl0L9CnyXALHvZ4EhpegBERWKYhNlI+LhC
Yhz1fgx65VXW7beG1WevZ83M0OPh5i30HjO4Hw2vKbB/i5F1zMDrNo1YVhfMZLFk
HbBnRFXbM4GSpR0xtYP65vAHLbTe78zWd52COBQrr3kwv9wSASBHVtBQmzDU6OgT
t+W4wDHXxaDWTyPfOf46YdTVw+SYl43UP1y+RP6eNqbS2oFMZwVG+L45oSdF3Nf6
1ISdYDAArtt/c4QjspQU5grB724b8pdrixhog7ixHzTf/307w3xNpSauOfgu5Npo
zhD3eK0A9qrJgyuhdtNV+pjIjadCNQtQY9TOTgjHR9Ncwq0phdGT5cpG+9PkULJX
kUrbpaAsuew0tsB90te4ZlUQ3EiLcRFhQEKwNoSum9CCDba314oDS1Vs9pxpIi8Q
BGTQem4zKnVm8U0fzom5ltOoNk1Y5oYF0UHUp/C+zsiR0489HkQ3ge3U+PKJaG5k
2zrRSio4pGGjcRJntErXqoaGBzuf4BqL0J9nU13qlrg4TP3MWT2QoaOX9hkMT3Xy
4akObs/vs+G18+1T2cY29n5LAzDtlbQvsumugSm9NHh1tC2p1Rrq3mbT20VW3e6D
fVvK1zgy0UJnEcScZDrN/DgjUEfZKiOMQHmDwgtQNBPrvEK9mLfxCn2ItSotSatl
B2bHKraQzTOjr0wTPVgvGZcBm4gQTU7pQc+J2sQikYvQaWNDl/CfsyxGdfYCRS2t
jT2L6mLMFO3wvVUkBZEW7FB/HnQL/jipNh4R6V5Lcz/Nirsr2aeH66/LZgV9v8WF
WEOSh9nBV+7ggv3gS+m1Shb7NBz4+70AcjEbHlSxmzpQ/AV+aWO3y8+I6x7lkUsK
D6IArXmNScOnlevstUurcdhgPF2zlOfzGRsBB3YBJxr6mPYLBIjHadwh28IkRhid
8fb6Zn3270OyY6F/EUo0P0LKJ2+Fh3Vtwd8EmE8nGdqQ7L/yHhSHgmURHs09UC3x
ypuCtgUXJwn9xbAVe+fyUgMHunt3TNbT4zuWxKQ/pPSt2rVYap/OzJDN4jljAcB3
iM1JiaxPee4DQdwtnM6bMZtZSAw+5/i3qCwO1Ag84GhL6f/MDfcSA7Z2szriWTp7
FuKPfrkImmBbcOjzso9rUd5CSxVY1uuf3PLRPeudBry64wJ4Zv7ZcH5xYEsAhFVG
74lbYWzyfUKxKsHdtjPgaGZxfuAhuZTd/3E01kKxuBgz+dY2w2g6KgPZMpcwE72I
HqbcrbFLRVYI/S9K/LztnDp4ArBVKeU6OOW19yAwf8ZE5hUlyZZ2HpDP5poYLfTL
IkDzIUj1NzC79yNWIe7dZdBseSCGavyZScEqwJvE2iSb/9whYIE80BVDQNKyfqmT
e6iWbFezIOzopVI0kVPENTLzsWPjaUlnu3rI7as8wYiAnGtC0dfyitne5lzd8oEH
DnH6ZOk1WYMT448syEddGLJeL6AnS0PlO6wTMGssPCuNgEg+Wv1ogDdvSiFouERA
vMZV5L4z3mhyekxeJWSsIGoPF+flyMxRfn/JvZWFmcBKSDY1WKNpYOlZ9it/YeUd
Cj9PV35rZWZ5Smdcu5maGikriKOh3ggRHndRNHRGzjY7qwA9o8FIEFsBiCjjt1EM
NIQyfv29CogugiCoOgjjUVyMkxIOnflyLclMIBhMEKnCk8hYZ8xPUFMVxwPDiA3L
sm+5+Njed7Auqt2YmllXlVowCoxsPV9NZOot58AYYjbiqLarLf4pZ64oKRb3H9GC
ME9lHAyDs/c83A0A7pTnKj5kRR3KJAiYnvXyYt/yqh6E6VBBRSnnllhh3UH8LHh4
ucYKF1qElHvK+Eb7dxhKlvYfVxEpsc+MbgOZkO8xMmwSTencxwWTR/icZjFF8iqJ
OogUqJqmK/tcq3Vntb8D0TtN31we7aT3MDQIy0wMdkFSpMRY8PTyEjElEiWbDi2v
XU+Pw7EM5Hd9VDk1jJik4RW1++O50D440M9tLLEUX20IU9Wf+xfs83Rk1aE6Nomb
o//tPrktF/Ik5acUhX0ASFBHih/3DBX4mcAU8+VzPL2NUiekrJVMTpzt18de78Y9
+wRyNq0VszUCKr8QKt9KihY75ip799iHXymUEmyVJ5woN2fziDNqN5e/zm/5NsHN
IN2s03zU0Pqq5nsektxzIO8Th1ko2mWBNLVjJuHcurPfNbN+Ffa1LEe3vr8LrD1U
1UinIIUWubG1PBOQ+elYKCzhI27FewIBZa0FsX2cOupINXRJWIw0y2KJ1X2ZJaVi
/VbaX2wr8Vd1BwDTD3SJ9B09NTBRWl0GYfSSNOaSLcLGGEkFk/zJPxL/LAAK+qvj
x52AnGyIO1YDkoJdD1H+QGWOq1BdSrbidrcNRznO76Rrmr52ROyq8yOEV0Vh3xOu
BZPDZ+T9ydwfY498dp2PjUloMzfJ0f3YoTciy1Uc+6Rm19pv9/g2BbEWpL5W/ltT
wr73K9TifxwnFTpQSWjwA52rTCTPI6ETib4Gn/sx4VfrYIqasWsZ4k3hKS8VSoKV
QuDQ70xLvMxygSJAamMhOa7VlvUTWjb33OBJG2V+WMiJOTzqGdJ7qcFwqRF/bx1c
sqydMHMyPFBTdgJOPZAP7bXRrc6ZfuuIxL6E9Okfz2Y5u9CrJR4y/FsC/0EQ/8i/
OCyXtCaRsRe10t3qmS9LN/MSrGgHejW8yCLlwxiwU5d6cdBv0qfFCn2/mmPrrvzu
oQfp5LXRCKI/jYrVcxhQlaWgfCUq5glKBaeLQMvudU4ojJUUdi4/jkXEmuAdmpQ7
+xwrHca8NST+v436+9jJ80lYU/9WoxLIk44UOzFeBeSMKWCivJO0T7e3stI25UgG
0N0rt+am6zYIRw9cG931WVK5GJNy2VnYCpsHMPOV3Cs0GyrqiYMC18zFRn0xF1Xq
BVfnmAqBgFKs23Or/9lzlxktDm4MrYqqU7Gxr/lJNLN1xkJMKj1pDqhjlswShxPl
DhrUlvm9xEVhA7EfsA2Lr7WuNfdlsHgnStBK3AxzV19pqN3eo7CvdIgHyno4JB/f
SVPRZE1bSCfRQeGLFjVOIsG75HqmIDW9w2IW6mVWJXJ09lwxTWQR3uBDbTZdHT9r
1T/TI1Fg+9Imo624xXxIIceCSmzFstfWOmswjGOkJNjmOb147HzZsAY33W57CUq9
THyOqCTzo5Von0l0/k8SUJ6hm9vSJQXTHx6+wmD9C2Cg5Uq+/bMUun8PENvkhWxD
nWDx3LKG+KSbcT3vAZI1fGu2GHAxJE0HxbKO50ppxzLWKm2xN8BLfLPYEyaya108
8QEFRVUpHoBGE4keqlDmDm6V3XOo+kWdABciFZR/3Jt/MWkZbsSQmTabp29ylXB4
lOsO2ibD2v1BH6oPQP5IS93Q+9Vc0FlrO03kIYl4QTX+L3Dh2yf6VnAw8hRUG4RS
OwHHx2p5w+8htUhZZxbijiwbU+BMSq0hIo2aJ1Lwwh82yHQXyqKOc7pE2qpxgefs
Lekf0TvtErmE2ws3ekvSRaEKqaadMVhXuuO09bBhvjTKr7oj1X0v47zuxLDoOglU
riyxbx79fO4HTM8aWyA2LhWQ7fezAsNQDCzmn8zjAx9uZPuLFKNJlGT0n/54Dmc7
Yl9PzDcy8uSRAqQ7jAcgO7a4uLFbbdAlOYJGXGoSxfyPO41wj4MtE/QN2CoYbs+O
bm7kt697cJFy+FkvaiNamxUw+HJlCwZKOGMlM1QDqLWkIZyLMTAh93BJ44UoOux8
f5V3v0Sw3KrktonVQ66zrROSuvxFGimK7DEfbe79ko2XP6E/l3Li/WeP3i9pAra+
iCjtphdRFYkn+0ebPz1toS7sKdHFbomsrZm9SyyBKwA2i9WzD8QB/wmvvFxBO6H/
Ccf3gsOcYVHsc0tQ8dNrsR4eBW210auTcA96vmvC9xoGiA0xThv5DUqYMRD7xhGU
4LkrbqJvs5AX/zZUXUox27xOC6AhhtSdlxh/gu+DycPdzMcqjt5CjW9/MEOs0t86
EsXyPSx22jB82LnYRwN6JNmMdeoeVRY8Uz1OkDqSZCuJ2+Uu8ah/Q2Ul3gsqEX6o
+IUVXdkyEQO4IXB3Zu4Q2AKZm6/FSNxeSbBF40o+8+iUavQOfP8q8WjIivFX906u
hxMKi/bG6vMUvUAbMTKS7QMnDrmEZOopvMYscuURmvofG11k3CBN9EfVoD9A9TM5
vRQI3n3zQZmeQbPHqjFMwhnDP8obw3ViKO2BuhHJe9Wz6WccXKrOxuexIbv6+Tff
Wav1uKwmoBNWiVlic5OYtiWR3vvOMmhh02OUkn+3UmopKrzHq4y9AlmRpS6EvFWA
4gTNxNw5MqHFC1qt+Bcre4n/jITB4xc5wJIs69+XZ2dqyHY0nXCH0yMGARll88TG
eIk9Rcw+xkEKVFltPgX8d7LT/FeJc0tkRrsMB9K+ph8BCaMfSiZpyYSgYkp42LzB
hCvFGR5Uyz3FaoTyP482Ixbd3T1BuVxOkPza9J1C0UNzZRaIwIf1xiMolsVxh1s3
7Z0pmWtsuqW/F1Ir3LuohKNE85B878cDrc8pySyLriQQdJ65FdALMkbyzugMyGHT
+/w4hhWmAetoeZav6OzusSzWdE+SMg/M6CdI6mivdUHkcJx9Z1A0ZxLhPfqfgYOj
7bBbI0yRRkThyOpx9HkzZ470UXCn4tU9l8Cf8GSbFx1svoKySMFbz9N8GJlnHPxW
CYiD0Vr6JcAsxFafrFjIngRCNSrnkLexBtoDtdbCCg54fAhXCE3V5SySs0POGaDX
XzIsN8CHFE2njGWzCGUVYLK7OzmRrM+UPOQITsy7/beX2LQk1yavofUqDAC6szwf
g/Utu40AaOyVJ1vYu0jSqENXcmvf3B3VG+mgbsYdwQTZQsQI6rLkgJSTTcvC+Qyy
kNkIlffA2uApTZH0x9FuoDVrG/pyPM4KxSt4Sh3nb10YmDgjdR0iIAgLWqmZHyZn
2j9L+lYsMWEBVf6KyBMkfVIy76Mzh5+dtsCZ2rhL2jcwwuIBwYEog8R7nEf75uGq
QDXUaE14smQ8e0e/n6Do2zVI9UfqTKBBNWx5xc6B5zCrNPEXrPKB/1oDTR1su3fe
qS/LQmie6G5yjqxUig4koZK5YCACylAICh1qKBwwSOheq4UB2IpKnj1RPN7P2ZwO
qPEsqubq+3Y8t1CcuctruxK9eroKL9U3R8r6IcGf2L9dxr1jiNj1Qh4fuDVEm4Uz
0cJuI+YGZa08XyoqDPD6ThPZiMdhrolQ70mGDolbgIsNYbX834raZHQ8eu0OdDC2
FBeD0JdKakcr2y3poOCVtBqM/MyXfWItykK7+Z3Jgb3RZ1KYSSDS/AT2C/rT4IbW
vbnw7l08mv51hYdYfASGxLl9saEyAtumyl36HLR3bs1TZ0yD0SATIyh9TUFqfZxM
4RUr+F3U5Q28pM1vFtWb73dIYAsfuyEWP6oTaQMjoADcDKFA6GGGLPHoQMZ+pTZC
CGhtoFuH3XWZN4I6wDZt/sa3tDc7qTGDfT9Tb9EWLr685w/bc+2V4599Ndeb5KVv
hG2ZM6fk0nPpDzRJpbe2YhydNoksBSEl1F5Rg+WcnsNdBulBrsP/dKXjcOCQsOqm
W7v08y5qDQkeQmap550IXqskZA6Xx/7pITOJml4zaYnPKuBzs2j3CF5tjMzl3nNM
oImDSGnQp8I6u2T9yFw5sT5U7t+/wRmGUn/8XJDP89dgT5wX6jcvZdNy5j7aDrCY
6osyLuIBku6XdRkk45ZzHLkp62VZmr7RtrCmIfMyzZy0IpArXP/KIHf3KSgcYQTl
3F/If1GXhXCpfPXqK8Qk/U4aJRzGMgwbI21D5DcvsCs0NMb2lvtmJWFha0TFjz+H
JrjuvvQeKYxd3Cpo1utsU2+N6tszqvdhzKoQk6FojzOW+s8oBkBrZ4758WhzB+2D
IW8emak9vv1VVVZpJNMty27X9loJTbizlK1ushNcaGF1q/Gx5o37I1J/7+39bnzA
sYL/P+kyhUiZQrDx9fy/aL41LUORYKTUWUYI3UnOED9TdHVgmkarnkULFxC9He4E
lBl1gl24+iJZn3vLUGBWVA9NHzujc2EPqnDiogqPcfih49xFBS6/cIfua8TSpg+E
fccIkILBDO4PIxyfqy0K0qAtc/s15fMmoFFd6d89hd211yglFn5W4hn4TtkTrpBP
PGqWX8TSBL+NgmIEj2Fe964F/TloQ45ItX9SM8IAuZsiyzmV7Pex+y/Urdx3Pdmb
Amfigdv5hLu9kIo+ZLBPYDX0KZYg5rceXSVtsJS392NUiw9K1X+Rj18Gj9R2UOw2
vQ1vrU2wcoTvrhtDJpiBXUGER+DOlwhYxSfORo2dP4ISaDziCGzP0XChWyk2w+1x
4eaLth5EfdcZq9WMzGNUwA5BPx7ZvJDIGcjlbqXHk9XjSd3xhlu8ubr29Dj9+G2F
WYESE3KWwlzZfgdxGgW7f2eXzbJZAg1bZ29rOLW3GH+lWTEPUmUOaMqbB3z/lwL8
f3xNdkuNhnAACn6Wc/CahQyBdI6bSKKhyHrpuSJZD2yiVrPEzfmQx8XJIcT3ab9E
S7L9CZSmNpFpSornLDoflDW/jY/M/3+Gvs4V5ps0tKl/o4ncf05GmgAIbS4xr0IZ
b7B+ple9VvGMHHiU4whUjwS7Gv8RedqNYDQPe9C9OghS9/8DBG/pYKi1ijcxKYGk
JPExr8svqCN+W/WUbkdv/m9nCxdmT4srj99RWoYjYIFEZuRNnVce8EWmj2KjzHkL
YETvdUB+Hnc33uFmQo607NeiyfeC2Mk6e7jaJSTXnjwr0o4UjwBlK2zZtD/RSY39
mq/d/50akpSjk2W/PJ6x9bRL3lbfyh9HwRMsAoDPS3mzfi9ohiKZ0QP6Kt4atDeD
gV0fuLpgAOttDYOVRRJd8BnyqwzD6dy+feVq7vVBq/3yHOI9a0txgdoWDOwIKgJO
5X+5S4zS0eR5nikWFO2K9/Mv38riiOYVJGAjQGZ2/mbBZRsi3UEyvmefOo1e/1KX
SKI1ukSgTkya2wLKNL3wea5HRXHhzUsjKjG+pHmNnAI7xqrtqILhZ7G/q7aZSMok
JuiDcKpjBOtzPtPSyNnPeXelHusbd7B1Q4gARWsbU93zd5qllnJX5qeBavlar/35
ZCwwIlGr60pkjmsHB4nmctTMaEYiJMFK4DjkJFHalxEX2tZu8CMWqcW0KEwAFfdX
LwrCO8JM1o5kIRZ1oQxRMJe6MrfmTXHs3Xiu6vMTMjrWXgn/kAD6iKIAU97Y4A4k
PY+iT8MUcMgmZI+3QWc3dIyolg3qLOf2u9vAcMRY1QampAstvwAZVLEx8RVHn2zz
UFlWSuRFPiKZFtNGXgSK3YuAwchrOQ6Sns91IsGG2Oljx7UIV6mG9YH27pQ30Ulw
TsuFRSUO/4xAFKSveDe9qsjPJExha9/f2WhY+gKLz+ajuziUennqhQdXHRpH2GZ6
cycms5Gg102MYQRdjFfpyreWybFie5yWhKw9gv9LU9WPbTIkvVft4tN9vorHoIvZ
PDC5xrS1M54ES+QE1/HY3TD1PK860HQVhHr+SA1I8NDAUZbaqF9L0ZNe0kpdEoPb
sr3dlo2R60UkHFfiiiHKHpEYHOivmXGrgnV9X7OYwCSMD0/OlUj5gCloaVC4Bcbq
GcaXpMp0yJLHfT0+DNsrAXqceDIa7dIiuT0HDt5Y1QPDVMQcRyK24NVzTx2fj1q1
OA6UFee1W32ZbMDaO9q3fBNjJFdtMJcdEoP1etbx4fRHo8Kyvcvqvao4EqeAyOxJ
khF5paCrhQwvm4Bj+0f4o7KCegr3gsU52f9WmBB6ZYkHcAwjnGlKLx7Q1WdEP4+h
bEhuoqtwL5KbbpZ4ig+9RzI7jPvOIlKa/KsEMLHd4B2L3wZz2zlC481mgzh3cY87
5kmzH9Md/13b9Q07wthY+B5LDKo8wj/Zz3iFJ/7PrGfFVa7qMMtAYygGYJwcWf1k
As3RF3UPSiNMfppnQt+JcgMmNZ9w7rz7Z+0EvCtBGLgKDykRouWO1oTJcMtfIHwY
77+/FIe3znjbCf1NXa4yVN49NjtR+WyskVF56aWu+ZSQxDbSWKtL2V8GaIA3lGDo
AMsvVUemS49s/AoRtkMApPT5BNZVWeh5jP8Ols72WHoNxxaSZIIHvG1AQMTgG4QB
2Qj9NJuzhnXJp8GywbKWd1eNAUOtRdVYxL1wVvvGnmf6fQiWAYkDx01qXRddq2UV
BeeIga0yC9M4gOw/z+j8wcbAKXsFyDqRP8kBJqZrpYNrlG93i9Jrl4+QlBeN9q7x
d+J7cX75JnoVyG4qzRpHdr/d1P0ZUtgwiSNEHWDQ413J3lJSsQBQaThSMS4ZcGck
oc6DyGPUq7cRaBwl6jFT71SuEbkTQKU+namUArsqRE1pH4TL+KyyHGNVc3ixJYlY
C0WF4/JRDKbc/aipopgyAhs8DhnVK7y2hkzsCl/Lt+iALZt1nmw2q2jnhrtSPK9b
VDbT/6DGXCZZab0iDN/W3Tkmj3G8yVVz4mo0BLlxUcZcHBmbqvKDWNB9x1udrMqd
jFJ7zvRPbEGyP6eq9RJlIOoMKWy62HDnaG3xUpXk7vls2YtUSuxAPfqZ2mHtfxWK
v7uLSQZgmbQ4ho4oJ7b7ppe0awNsOBdQ/wrI9R6A1EX0BiXM4nkbZslT6MbBADC7
oz4lwc60i3S9J0GmxrJxqHAb4m4D2n+X+WkOUrUfRhb11Y8p4I0A56+M2s1DwvDB
vWZtmalQ5DcKE+vpOUN6SvADxQSu8nYkEQOsZSFrGv7gVLGxnQ4GyL/8muO3Yw9S
nKdbBC+enVTW+LxIzDICJ7L7v5QJpAQ4sJ3WAprIzsA/5q/FUwufsgyi5v7IVFyG
f0RVi0/kwKHoN1OBgmBiWRQxhxb8JPYVH64O9dMF9omuwbsP3E/MH1j59+uXeakc
yX31enCoDQxIBLTyLxfH38BEtecNm0Y1IiUM1jzeVBEcRCTJEShu8f540ixBRdrV
xBXRUu1wPm7kDQTn4Mkprtl0XCVyjs+s0TIJzTHlx5/BMG3aCpdeDRBCy0MsiBoL
ftQCf06NFApbkEXdiBM6reU4MxvAuedG5TdmB9vivt6kMYugIe9WaMlAxDx0pj4p
gSgAkUUJKL88U4tN3tMlsCkLlQlCM5ZgzIlouadj2V9yM76a2EfZiEE4KT/y3SuR
SReZSETh2r33UatmVQOzHWjcQEXgi9eJq6r4xKdKbK8mGzq3jGiCJrSReZ2XZAlb
WvyatWPAk16uvvC6juuGNIt1piS1/U/BSgtRByiAPdCS9GVZm6tUvSPG6i10RbIq
2oUJ2Nita4j4MsBliySO5MJX03r4PuRieNZ+EqfKx1DRnsq2vToIeBJsTCdRpOif
xi7Db2Q2nhzf9QaCqv29UKXtLnuvFPpdQPMbHdNpTSxLe5ZdpvS2S8gvL6wdsCZk
cnYnpVn7UM8s/4nYwEbsp79AsnnPi44IcA8x2l3js4DmXeUiQqww9YR1iD4piaJ9
ilU5+1AfGjx3ZACnGamvw19D3ENUM8ryTC+wY6YFnxlaNAT9r9+SIhN2XUC+VUv7
7PLUP11gZO+x2q0j7Qi+dI+Lv9d0Kv9S82GP43VNTIF+Zy6KbcfpV7Kz0oxtxFOH
M74lFIGb6NJhTm77WM0rCQcopoHJnhPWcRArMkjmGoGiSszs/yXy9HjL9mHxCTi+
HXHMQIxcntdvjUmWJpy5/gfkDWmNw5gC3pse/mRqbw7v29GHGi2xssDtQjdYxUq1
LxzsmdU3TSSugUK8v9kemC4lAbfC8kU3lVqf4+oDjORum/O7dEsFOUw647bmWzIN
sXpRh1/F/xQEI8jPSMmXPhk8aPnpo1XQHorF0eiqxN3HQeUgLWbin3j3j4mWvRI5
qgf4V5DcSd+B76X3szTmmxXat8J+M3IZrPtyOzW+HAYwhI0c4zyK+mdN9WZxuF58
3Gr+B3vKKYUn/gXDX88SgcQ2XymQg0SZVnnKhVczjz/fN2WW7x+RYlAKpCn9JKoL
tR5Z73qe8CQXmbx8+2C1DdyW4+ThnFdJZvM/5Dw7gTbQ8VVFFtgA+jvVS/IYbeDn
V3hny/RGApk4moTkdW+Kv2fw5yp0KmEVHI4sV0xRJ1JhiZDnAGQ7gLwmacqM1dX9
XiCrvt0a45m2VGZ3o2fy09qosNs8nVWDIJtXQsdw8T8dy6PC/i0KJNCZlsQKZJlw
QSLvMvWa9Jr0k/Md/qJNO1bk4EqQGvPBEnhcMMJK31su7qpQZ4aUJ8PXqOuBcmse
xhgkM6eSyWTcYAIHdHi/mS/UQ1kFojtwZGs1IaY6UWlrOG7pxHkzHDGkvmgfifPp
CMM01C7iXzWYg9o8MLZeVK7Z7o56+qVRq7WExWFn4dYoKqxKAQFIi5UldkVuw63I
vy2BxUosjPdZCWglR68kA2bksV9RXSW4xD2V+sb59aXNc6QO7Pm2UwDJqqH2Kxp+
jq2qnuDtn+3dOTYzhJ637sgMLhsJ56acYmlXLzKCLftG/hk/aQA2ANEEbdnSjC5z
0SHbBGcOzMpavAjciNhWcnV55due1yLmmwCSQk6ni8fGHMQ4X1hcfN+PM35nRVYx
wS4ZePudMwp3dDF8sDvIGsGM/xHz1rGc4q6n5xHpmu0O1LtURiU59jb2GjLhQf5F
mZl1Txm81ihcwwioakaWvmmSPvXycveJIWdmZVTaX5I2/BapkmD39mtBjgrZF7Pc
rKmGlpXNKHlP5eIHi8zM/LkQ9VllbYf43iAo+qFuEk3lB/3CanFpcNBXCyH7Tymg
eWRQAYrKXOkBeiVUjbCTgkkMVC//AN4ISTivtQwNm448L4qi/egH3lCmN13E4tUq
hXqkwYXYF9xrdJ1WyFVaE1NCq6tbH1jvid/5mgBTtCopNhZqV6KKDuj3rgRNq8Ei
W9iFieIkJDDC+JGnKzyIuEG9wJlVyn2p1AVwdNwCkK64s0OhGUKru/HOX96dy7I4
aqFrk9cqyQAh0QOeJFj5udclKu9cOUZ8aYnR94KpObd6n/opu6k2H1eH7Wzf0eB8
KIYMESkh2EyJrHln/BXXdKLN38yyxlpEuLvbC8fVuHrDk0sCB7Uv/LnOfkIzFul3
AWhSKUdEF1QbcBBNN/Z6IDcN63mJhbJ8nqITAeDS2pM1E4jbL/8GpuwJI7DBFSfv
YvAq2oAJLCkSRPv4bTGlYRqCYAk3sCPgms7RybdJnUPPgNyCZPBlQx1ZjeY7jR2T
4HG+uHLZdaMxSi+y8e7nz4jSc1cL9fMfsdtBEmGsHoLPYE18xg5kZm5uixJLAsMZ
tql5ETfiesv3c02CIvb2TgyG/cm+A19rm5BW9OD1BVlTQy8Lq4Uk7LnVNT3MGeuj
praQQ2nQxe+3BU+Ailux3wHKonVWUe0C+Bong8xSCjc6yDUK9bENy5JHyCeqVuYN
2BQXolqoTXMo5KtmTpLKgNhLKpdZunD+WhNONLYdaz+lU52sdys7nYUM21R41v08
jnjNFuy8QeaU0+FF2x70WcqDQxxDV/mufFmf+tX4M9+97JLqAlWMMxSvRl2YTeIR
I6YaPDDoFXv9w4oRkGywEKMJEYGmJ/MzzwL/QQWE42QQp7jcQYzja6YEiUjOqit3
06cUlPWUgYndaq1XqZLwgs3ztrdxG8GJGzOJ92mK9IaemwRX4dkVsEcor+aHZJXn
3kWAK9YWWPyqUDDoLc4PLUfttEKvpEJ9V+hMXQ4lXiJaBWdEUyvcVIx9vrkC9Yjk
aeCbDA7ZcZIY1WOJ4K1lO4iSNSBlDCOsmovLV4Dn0OeUECzkEY6zDlLyzzmQcrgk
qvaApUsThhzF/IE3njANQznB8zK721tdTO17MqKjYBTTHMzIQsRs8RFGmB8lssRc
it8B5NWCyBagys/snxkOzsYB/qI6cnXyO/rb5zoD28DlSWzHL2WeqDTIce9ToHFZ
sbo2MGgqgx154rcQjWA2f6VNzhz6v2bdlhmTOY3H77wuT/yGjpBeVg5mCDQ01hUL
0pd9oQlN0tCba5hJPj+AficQffZl68+6tLF6M5hoRIO5tZ971Bu3eB8xkCaSoArQ
8cTlGjoz84VEzIgYHtSReDqBf79RMyp1rDAZ8o8jlyhqySkAyucRNQJkPBZJvlhN
MzMrH6DUnt8bKm+quoVroUx50NDlwxVVQjR0uoQYgIsOa+nkmc4UixWaqmWzGdtX
UfoYMk197roi3ZM1N+r0wwEmjMaEYaxnI7leBUmPVqDst33fHzYf1efKyxOSu1W5
F1oobwRqz/7/GA71qiGhKC9uF5FFMVnbt4gEeZjdMiav8AOxmzzO+vrGok17xZab
gQCc4pwfoAgFx0Df/Fpbtbp4kgX/iNIPYZJirj4i2gvGnzoK3QSBt1B/VGnphvdY
ADUS7XsuTU2v5m/Pe3CmT7CHcyZITasALceS0s8P5fkEZxzSoGn8okq8NE2bODlk
hPGrfI+VIrUU7vSpLy6mzYCikVZx7eg1RFcfUuvJzRFenOU2AZONPPBXAoLujJzl
yzI3+nIHYSfL87NqEMCRWB3aE5t6WpNEUXHHyq4m8kHAVNCrU7GfYiWffBof6A/s
V+qplUYZr6sWjBj2TNiX0uhIAPGkXYe3rcqFQ9vx8xTpZXFLfAilDdf1EJWtOSD3
s2YsNKftx7mqYNZnCezGwwDNtn3ymo95qcYCNr9RW7ceMupg690F5b0059bn5Z9+
HuVbKqaslL7hTMWsOedF232UDc0uK65thVxygxVBjqEoLFe25lB0lqow1fFGB/vD
EzTW84PQLFu5IHv5/GaHcTb+yQuIu+jY/3Dkw7MaoiPajjAoD0aUoVl8cjcXb7Ow
MiKcuufmEc5WHHzvOp0UVgSoA39VoIqp7pwEuQTKJ9gAFoZiZ6/+LGzlLnaNJ4vW
GLUq5tnR2gFWMvn5dzK99S+wxPGAd+OwAfbfOjFSRXh3WF/rdze8ITRSizsGBsVl
+tmtHBjVJ3OBMSz62B5Ufo4xtjDDk4+ecY7YLttX3Piu56zVYy7SMIBFkIhVppGK
TbLEAhrWzbBu95Ohu+RiDMBtEph81q+Dwx7AJrrrvRW1go5Wsup9ZMwQDyJr6pdc
FDcgvWs6/FZqAyH6QX07aM18J3puW+52cFoHYeWIUNKZ0LHAu+pYXUrUoIuuKwVP
C4vl2NkIO3WSwJ+IF+5yQykEAHv34Bdnixg8r5H6z8aE+Kwd3/1zVizVUtZVT6Y3
t5lNAzCbiCxfSapyWXBwj4Ijp0GrERuVZhHn/wNHSkx/FfEWiLsgTHnUuaZwv/X4
MYPKig3DXMTsKNweqaemJaldRu6IfSo0EcpgucrUrYiYsYAef0/u0BxgYiuOOe8i
dj4IFXKzkygEFKY2+zZ4Efh1kV5dP3hVbcK8aZI9vKaa21hZ3GCNttobQY64Lkd7
nh7r42ZyKTWhcyEZ7etKRjCdomFfJNCvV5z33s5vjohLpE2vIdo199zBFHk6Zxy4
WBSvH6+Kb0zbTBZAwDWp41N6T7pbVOcO5T+SU+7RYRaxcX8Lopnrv+gXQE6nZZKp
r/NfOylN9N7Mi/402qd2epAzTV6BozA+p44IaeY4beEFbYJCUkLaDVuVLk8IpOYQ
eLa1Q5Au4U/DV2/MBhTw8SVw0hsnbYs3XzvG0daJm3ew9JSW2++wpM9HXUONdPza
imAP+0rk0jGGhsnCh+yB+Ekg6JFR59ijwmMAIsssW9Eod56W5S31FXcTAXmtUX23
2szQnxqjWV3bw9JKTIf7pkNalEYfZYaePJ6QOCCG3NgIGWVZuCySu4IKxBMNj2uz
Y29QRqrpk20IfXWthR4jOZPzlF4MaiIIzQSqhrnh9Bn9E6jiNTM2o3Y7kcXcGRh2
NO71Umca7YoAPaWdQef3l2OOKaGwpBk0Ek9w70sVyE+aAxQYHlHOWoOuexhjWtbM
sVpMQT8Lm0/qL214PAqGgDw1CCXxEmvyP9aDZN6Agipd3slLTOYDFL2KE4PEGF6f
r1myE0Wrvk82FwLiFJakCRo+LJJ/HC2iGrVha084y1UMWue2c5auP8v1RDMs0E0W
EGtNO3DkWDnVGDaXr6vt7QWwXOF78f8ymGw6YDNNVBsGqKzK40DRjIEKuAHD941D
qWIkjfOjM/grGv0mktUSd5Hw5nU6VylyYnklc8pMkChRYrTB5Qk1r6Wo29HKTY9E
PMFM5kOsduSf1QlzC8W8luiP4YzNRzW6vKzn9MjYM7ixPjq+4GqWX2mQXG/UsOCc
l9Rh55FVeutzdiNTMtw/UHDEbpt5sOeLbrkKhlIbXxKd63RtH/QpMe86YmHGz3oz
mYX4NBNatFwPXav/czRrTsGNzlGyHfN2aApGqGXPQ0fbNC4w5DMK2BBs+Z3p5OcW
UYoVANqBYIGgGUxeBLKcutPCHiWgpkT3GcXs3gvyP79Evx0nxOm/33Tjv+JakOI9
YBHf9t2Thq1R1Hb3qxou1rIWQ+IHlbq2ZV5JH3BsnKwGaTgHxbV+WJwXskz4d83K
EdJN6K4fbTyiv93rog6S0chFB1sXP9pnNzUH6t2R/3WPmLRCZFSxwj+LXdzhY3kG
jEbQD1D2JBKb4uRev3e/XdDdoHOd1Is5uSHCz3yUdMQuygdFxI65apRWg/i5vQdK
rNiVTue83uEMJ22Ze+eqkSzJBvh8rtEHGhDAnNC20oqAVvkkQRYzRnId8jr28bSS
ChJ2lOdsywPW9DjYXZIqGuCXhCqi/k2GPAnm3VNZMmL6YRgQ8KeaooiAICZGpIMS
mjFNo7BgBQYR53A9MWHQ23R2LymDsiqi1pwOVTB1VE81Fg9j5EZPrz6Ty6aRWFW+
0wU/c8jFbFBv3GdMlxN742s4hPfuMbdzEnMXQqqErOFfYCZMGyV+eXHpYKNl2Prz
GBTBnTq9KKJYhFwuzLygroiVnRuCqW4h/Tziu/8cjz7WdggX/vQdVyvnjECIQRCN
geJqcYFaT3F5h50ES3kRQvucT8Erzp7qyqtEdy7OvYlM9YTrOrRa65KDUC+nTcki
X+8sPmeC+pE5QGuGBsP2SJ6qc54HkFrXHJzTVxK0esApvc6aJWTI9E6/blX6VoSJ
FBJwuSjMY1miF/GlqVx1Dg0q217TPgUsP8901iek2LO4i2sIJRQQJeQ+cncEdUk+
m/6Lw9anG5Rt6znAAvq65AmhkNq5Dj+XCEakOD5useXQRhDP4wWYEIU7GLIzaR0a
NQYsvwdn594vsGf2EsOAYmJO3hKB7qwDFAmLjgCQjHsisCM3UgMftwaGH0YV4DT2
OfP7IRbsmNbmhd4a80VoD6cowFcoDn+gcVKK63Pdy6judd2RvH7YD64xLgonI6o8
bIl1VQWedIXAqM/9nMR664Yd4pS9BKTrgZOgxJiWLsD9fLs64QfMh9iQ+MzSGmiW
h0johOgW3O9d56pjDc1klE1ihP6J+n1pFox7dhf7cfl95t23A4jVQuh6/8c6MVMd
0CL2Oinbw2m6ZpxYOtIb9jpIp1e6U7YXmpsjBjqNfjRRk6o33HE79wIM2j9l9QiX
2aZhlj0LxzAKLdMqdx6OkYIB0owEhSmtKx20OngmzOTYGctXUpKJO5OHeyGqfDiD
zOb83wWoL9pW9UiEE76WOvSYNAVmI+M1Eex+WYaQEeVXLGmO1E3nVNDQzy0CbSl1
MD8QAJClKZ1NHzroo54zPbuGHerdfAzcCIOp4IZ7eI6hokzKfsy6gIlbeT+xy1XO
rqEzdlXG/BKocFpLQ67Rcd9Qynmiwt3JB7c6zzz2PjK2tI1TVKz8hLBAxDEo3TQ2
37cVc5+ZsMrdXeLw5WE737T5jkrUYQ5SPFW5KhxBry4AFhGcE4q5deNhDF1t9UoL
rcaL1HPwH8C53X2LNiuvvINj6WlG3wfirL1gWd1O+DRq+lm7GQFSL17z1qZiONpr
JHJGjwxvGLTySkPRmb9wdd/t3Bq1V0NImPgGH1wvuxhfMOj53u630/CsMHqnEVuA
yjkMxeic3+XgaADXkuM3GKkCKXoyPl6+pwLUa1bizQP+9fNMLKsiCNnTCfLag0Fk
UAqo9LuIApnxYM7oS2Sc4dm+PFE/ycdj9O+1ljg30D//yop4gEqjDF3tEnT1viqj
xxkP6OwMSST12ym4K3c1JMiTw/PCMGp2fbDtcHfQIV8SMnmrB6EONWhlwkQ85Tlg
tizQ9w/91RgbX90dxq6EUkkwn3utxYxfTUuInwqjM1a0ochKRIN6irU4Zt60Dx5V
8iMsFFJwvqqpEDt+Y6Wa4HFVqKDkJ/ned5oZz/STi9/pctYdyHf0ivf/WM8+4e+s
dcwERGD9OjZKgg2E3QJ1c8rXEWEnZO/SP768JMf/clkLzOzes+uyv58zImytkvfO
ZIZLKXEDa1MJTr/S+XZH8k58TExo+pEfD+1d7yjeE6eGayD3HC8Cyjj07TmTOIeF
rNxn6UgvkQkdVEhcokZdXAPUVLFLCluhPvSuEJTMB/RKim+0WJdfv3/4wlxwiT8n
ZJpmQePOXVyaw2GVyWjQ4OKMCZ2YhBnqLnNPiwzoWHE0AW37LHsHl3W9VF73Qiki
Kr9pEmmikUkdlvKkWNeQIYM3powYwjYO4w+Gw/G09nPUUGWV0BDLGDSnxjjMu3NV
cP6V6RbDnv6fSpjcuDP66oShJ6ohzMir4Gp+L7ogyLeewDznHmzaHvUDRPC7VdGl
i2NMBI8NS2BEW7LTUZbmzW+BTiFpn8sRU+UBe9BRSZoqT+jXA0b3lOM5uG2YjP3A
92i+5caw2WvXgKcw2B9AJoZb9Hzq/NwkWIlhrtI9NCDAvjAGH16vT5qBEsjlxp2x
qKhoMDPcwm0wip6sXXTYzGTkrA9uCS0vx/oX1bhvj/5CepPq/WAJrSz6DdVXNi5U
rczdDQs+iqy8TmpBYDTsntbR/ltZrxnOY8Cm8N+Xr7nSHaLMXVGvOj0Hh4mVBjih
/39Jevbcda+pbWhx8AWUGTGNXKn7WrxCDuDGfjJ0j7nytgIFncNvudDHD5Ix6/LZ
WwJJKQGuYN7YlzW49194l2WdljsnDLCKLb1ydvx02OAv1WxMNzx3tJWEkRt8JK5N
k4c9lOli9GhxhmeXjnWCkHj3qvHzyDLSgiWntv87kxrCzC22o4zL7SCYKEFvTScI
j7A1Hr9xSKhEoJhl4ti0mPZB0ghPJBDbz24kluRLGJCcFIGQlxSZh/Sj1LvoGH/p
UA2SdzSXJfiovYkmKlD1yAyJ5vW93ug2/xTEouXHEUGr/v1Jc2PQHc49CIBi6HrN
Q2viDji2qkF6/RpDCrSvbPS9N1r33K683qmy9UCQvlY88hoXf5Q9ZW9v0JjnMg2v
MKh4ZW/4yGFmYlsw+sM0Q+bDmPbH2dS8vYf86XoLvgpreV1zSWbPi4VG6pFT8rxV
4a1Eh9rye9MfEUqg5AKoU/QbyDDACbtjyjeTQ18/RZn+PnoyJCF6hiW4vTdRm03F
mgNFJMIYrSXNKHqrc/8GyuzQlnxot37tDLeTsEFD4Ikqox1iKdgG/i4deuCeiSPm
c+7q3fIynW7Swez3N6vUOwANgg6/hLhcsR22lrwbuEZNG+v8fOuHMddV6ma/dac+
LhFkxImJNvMweNBCkrrFAvG54cwSq8ZiJ9mwxAcpj1Ar+mRNqZMtcZAsK0FNi/w0
ERW28h5Vxj0YOrmY4yrYK1G9Rw5Oh4Lq8Y7hQj00fLYDMUn+SHGickw54jjbr6Lc
T4VrnmKYlifzLCc3RbAjj7ADePQSCeN2bm4lXTbQfteO9sdLzb98B5y6Fg0td6Ar
Jm05wrjPoLpP0lV7u+uRcnMkp5jqfxmjerWIhHaMjG3eXJO7iPq+zDuCTeZ79WZ/
EQ458GSHuKlWx6+0R3czDdG+7ie+GZvKvKHnvqCDLj1lnBuUvz50roCRiyazeDHa
Ei+tKcKCj08tGTXqJb8JblnUVeWwFfsDWuo9a43xas/uO6Iw/t7Fl0CIDrt/p//C
pc76IOgjkJ1he51xBvCYfnJf/UdfF2OycJhFe33p4isYfUSXT7N+llJd6542y//y
zhqL60MUKHw9ngR0/6hqnSpmCF5ehTcQorKxjuug8HklANTw/o+U9+u7xBy7cPvO
Hnh4dbiAQK28urLCDWZy3kT6QBNQ8Xu5xi0fVqio/XJvX1F1HgWiUEK+hdOlnxHA
iMCGSGpbANLmh8cWuVns4nUHsxlq+K2Q/EFQlzjvvyzLKBpzQJZ0XnBvmozo6OtY
Dd2G59bWLNjMLPFLbV6QHulZ1hNXOzmHBzSpNdhNUhsoKQSiAE/muq8bduFqX+Qy
3LoTk6kha1512/XQDnZIVwforwNgDBOjhcMO/3jmLOoTqeBlczsmmdqr7b0eF8kG
tzrML5eUUVioYLMmYsKJpkh4xXfcxn2o1ndU2/tfqy03ICxsiVuvVcQqP8U7JR1a
hdmtPg5d+FWK09b7ONHv48646q0V8H5gDbOAySNp4myW7gAXAbSHE6LrDaH3ewYJ
lVKmuw6Hm0F/uw4TOZSN3njOOnv6H8jyPWq7fFTGBVi1hqFhKg38B84IP06aNTjN
7CuQO6uj7i0M/AY0xuH0sZSl9jgofQlcNc8GbnlaFL5+I0z22+KhakU1XgUx3ToS
MGPqEKrM2WaNuKYEPCCEpuGjRK2N+iwUjt5nZL8whXmzM3ice/Nprf/dnlAIBmMd
WzdJM4CQhmcuhD+97BLgyzony7DoSvQpyhNBDYeKFMFA/xbgpV8NBrzba3hobeuA
o7mpWBzJ+RFiy1z2gTglRSxf2QNXixSrC0lzVL0Qf9mhEPnwryKqH5im9dj7raQ4
WWrRFWET2ds3SjxvG11kv/O6f8CGfZX5mXQ+Q2Dq0AKUFRl4Ma9yr3hf+kLVMwUg
7xn7jOuvlhoK6vzV9RjPJWVBI53DSUfnJa7iH11e7XitQMW/ITJWLWX9fcYQYE7+
UKfyDt32xAKe8Q1iIP9nHBBKYFPULn9tY66rqdwQkodv2DcJhOjRUAQDkAbGMnlA
zJoC/IQ2RpjT8RVVwA7TBnsF0B1VV20BZRqyE20NOMGJPNRlmCAsyDLENbjqyWBx
H3bBdR5uLa6zCXdV3klhjzXyuPqa+ohy0LhESH8ZaSwOiFSS7eSpgyVZh3O00QrR
i2NchC/TS14jeUdnKwr6wcl8LEz3oegqeAeysyVriAcd71uJVS+q4ksgxxadgO5m
AFzbT5NmEBR5JmnmuYfMPQfplVk3E6iQmjpSTgPjwJ6OgbuLWSZfxfGRAekYOwLV
Qj2ECeTG9m6JpPYngoTz9xk6FyfZ7gbYe94ERipblhOuKK7H9wQv2Lbp8pm3Q0UL
VafrMQSOOBRPEiNvwX6p3KZOl6dNc1sVK4KU8qFbqzEckgwxSkGUm/yNkzf3gy78
PndojCZUjrzc8T5LCT25Zp3uGvvZyOIo/unwRlwz25jT85FwO+ty9RF/wVGx2APg
ODBZ+/arFwy8t4N+ORZsalmORB3bmUab6Zfj1UyO6q9ZLmC0ueFAvcixBA8NN1qP
iB2s1lhvwjxUUrAS/YJgIpb6AkRNl1y98ehs+kbMPakKpjLGwJ5dECGkam15uwwD
Kj1EOoWgwp/uV8rrLF4P+iucRTKAEVO3HfP8tGluUBfI8Q6KKkyBicH1PUyY5/ys
nh1y3pbwg3EcJXz512svCJ2eO2u5h3YFR9Btu6uMNkoekZB0DaHiP4BcZ/08GS+k
QI3gheRECwe7GjBqvQkktHXK6cyY14DPHSpaFBTKN8OL1keGrUkplY7hDYxv+oCU
ntp6q96wIcifRAlF3rEpMyuqXuSPCyKn8M7rM9BrgbA6p5LXa6XdERIWzhJIeGVq
auU3Vt/Mr4qoSHIUy1goG9FlJRmsgIUDHmPiolw3KTI3bIIcvG7hOoMRz3Ns4KLl
6rKyvXJhih5SMM50quqGkhClI90zR6ldFx5FPQkRcmpS/uO8PcGgCeiynpkVbnKa
mJeHEzhmNky5CJ2SjhkKkXPl+V1IWigxuf0crbk0e2rX9cHkXZnvgxbdFtEKxbC4
3zYpeT/BJjXc5UkidTw30Y94Pyn1I+e2WKn2mSWKbYbZAvI/BvKcuQwTVrBKuiUc
a+16fWkU8Is2bhAmvp/eYXzyDNaAI2LExu4+dMKNbr7WsopRq4Z5fwC1BIylyoJ7
vfJJ6KbPgrj6vf90l2IEZ3ddky+Ra7s3KZ+p44KLAbCQP9nb9Igxd80Xsj/4pMxl
wBYp64ROFjV9T61N5cSCnNbuBFdtiQHn65lFxt9BwJ2oJyHyXdpquM/CAB4I9FIJ
iEJVmJBlys2eeDmPMAVixB/DuqlmMwejg1WmErQJLTiIYNzmZH/aKJHBjHCC9zcE
vi2FDemzKGIYP+4CZztHJ5YhSqaVmxhwHngKapa41cA2MEZ83b6qhOZsVGcQDr1M
CpH9jD7ILM3pqpFoaSTcndZfsx6Of6FUy/v7ybyw4SNnItxywY1q15lMzBk+wFRd
wFj852z83aW//Q1z5lop76M4/LGejd0r9Z5dECDAcoGWnfZdEYm97zhCvnZR+LQ3
+NGlJdUyTCBd0B/s8ljoZ5GKlRTJOePJgdBCzAYxCOLzmNpA8LVN2Igp+ikP8iDv
v65Aqr15WI0iB0eezXA7/N3gLbkKa4aIkEsa6KG7/6GyBO+Gymc0fzljmXicv1B5
1AIisOaJze7FOXqH71bFTy7rU9IhG3wtsUQ91D+FLK9d5cFEf+TTlPI13linl+5r
SM4LxT0mrY2Xui4b/6UxMFpCYyH3bxfJYieAeKvi7bIJyeEq3IKABrTjAFmma/hD
/6/IM/8YCBnxBpKSj67wHu8xLwgItCqHFncpQjYJLfkpIHN4zEJlIPVhIYyI8s3J
UZfLNlXjbdyTDRLIu6uBO1c5/yfEom5LvvuTFZEht558io85zWNCSByDLwvJtfcL
fp847y1s4mvG+nVvs5ZH8m0mJNZcK4Qj7BTh2e7RUEUkRyrTje+i46fZYH2Ntkrp
Mfook/MWLwacsN+K4wgdXAXsXXlJVamZ6apQr4+K5Jmv/AF8ZkacLOTHzW8v8wGs
U3QG5bw9+BRwMnEcxFOuQ+EStSyaRcNumVPukXhki+Gifxef/8lYpGpZGFygyPwH
lhI5+T1E/j6jGp17OxfpWmOLHd0UrpqzFqCk+ApJ6gV1Pmj6pJvi1gxOvAb1vpkX
DTcqNBAj8JPT3G74utL8vydr5bD6cew6bHwwqEpnMcc+HInK0LEfC8oVSZv4stGb
lRcmo353EvKQIpvAhDfYx8T07pqEImtYj6ihYdRvz82nIhuxvOvN8Zdw2WdII61L
GKurqmCBsbng+Yy4hesZRJAj65B452IHtJUP1bBUfSziSpvmj/l6dM3ZEZz7TYVS
MdLSBoWoiZmJ2XmbErE+kRFD7PA3PqqKmJJkDyWgDUSIlJSGVZlsMI1Qc3bAJ5Wa
XhyRD1qLLmPeLnog3fjOVmmHnJ7MnNfvwL8iK1jK/cCDyBJs4tnmgbsTZw2KOf+L
Erqc0/ibMnvjoCHbdJpOzlTL32ISud+qjgyUN59/r9etuxqmgItZ/ws9bNHR4h5H
oPoCu2x/8DHYIR9fRp3ah8ThLUU8gn791zEWg0LQViU7JvaAWnogJKZ+TLcLu1sG
m7UKF2EDO9JfskPZ7k8cSMYiwJfNRLXiDiKJZkjtjzguHFjAH9Dz4Sm6O49Ed2ym
UjkI9TSvxjXuWqSOlDnf9fvbMeCDome2oUZD6zerJ7flf8/TzrXJYigD4pTS5N9W
WpnNTCJrDcoX0YTS3ZEo3YgEvTAp+tW/VBfPLQScdxGK06cuJKOWKdB2mQYmGg4x
YpqACYLQtHLQyvu3H02JCCQCMJDETHlOG6A2R268XPGauf2q1QwgM0+w/LlXs8q8
DJ9ACp1WsiMNSn4wPsKQg10eV8sQAOw/dWr148KZLU5derqltSHYKtZ3x1orVAXB
+8LyWligws2/xhk1uXRsiqh8tBaDpxMy2f+Z55S1dEu/g9MWO1u0yyvCIy7qZD/Y
6Qnlb+VytVawJ/S64ioZcOs2M4+d7TgYJuVugSGxq41aRsBqv/gvechPHbhcSRfy
EOg+beyLsKbKuP0CytWpDq68HmcsfgvM3wiaAqThwBRRPkAfw9vJ+5MH/KMOD0sb
g+u/zf1BMmX6Zk/mPqu/lyLX2YWevK8Pt2m4Xvnl2PAwnkMvl8mx+YCaaRTVreFB
BYtwzTVRtkSUEndcxE93qnfZOcKg2E3Y1PI4JtJXTToeTqtF2D3SmBDIhuZLpSeY
cVf7+d11TqN00d4TJKw7ZH4VgYqVqji1FqNSKRKGNvLPsaVE+/fnzIiz6si2WC1+
DQ1l7KLzCCepRefEITQvyLB3s2Y/sGZMAJuvm+9PjDpndhKY/V1ViggftuWg9/wO
6p7dsvrn+8r+Jc2wZhkWCL95SDyMZg4coElTjo2aBYqQ2ipwnq2FthuX0gLPWebX
EwxZvgMI2CcY0cjn9JJ/yGOfif39Km9lsb2UPi+/nx6hahSgz74wHFULd/svg4lw
EZbQATh5OvCtqO/sh+gdPnC/+qAM29fhf1SQa74aS8LjkVya7NrNd62KGh1OaOT+
Dn0ksM33O8LNpa4kwgxVrFyIUETdsiZI39Q0mKhizG7S7HuIUpBW7pyDSgTjErL7
jxn8BE9Jy6vq3sAXsRtLAwk++0XI4f7GdIgtMeU6G5DfTFim5vlTMNGXT6WpsYt8
Njk6aTKE6Plbjh+3+3Gy0NZrCnNpUB80XXQI9u9WGQwhDEThDOQEDyOnordoilqs
oXabHVXmYkhC2oAsjJGSjZiwibKVN2CML0fMLwn1seSORUmVNUPAPdw4kNPkqQDI
Tve2TJ9kVBohQTL451ji90pXM+KQooPskO+VYU5ARfHKu+fBWlyBiy2DYAT7JE0P
6MtD3L12q1xvLqmS14o4uRe+qroLmb4rtcY5y8OBQSfvNgy8nU0plvU4v48gIo+B
rEZOp/UrH/46QZelbliWl55cGUIKJJnrLfdWZWFliZQoS03Rlz7OucyiDYg9JnS1
nb1i30QDtrp4bANNc98ozGkgKtKBmvScln/wOY6UIfDgj8CwV/wnjwBWiEEFwTjM
4jzO87gdLmCqPhu0zIWmHZfcHyNTWrKZvffZeUXiDHkiG5EaAcWzuED2VqptvcLs
x9XCMTyJhuShWkEqnuZ6/HfZ5d/4ohCBOzKkYzWpIzzS5DsUofGHGmf2TCcC3wc1
t3AKxLqiGYUuCCBO4C55wgKFtPiGpbEhJnzXjb4TB9r7OI6nyC5KvoDTktSRzDRa
GX1V9vGIKWbKiZv/QS+l04OEZz3cGE70ImJ6Tn9PRg9D/c1Nze6emTNKlIX7PgDI
5eLVbZC+MLX0vHoWj1ua/suSvYkuzCdQ+f4jwnPUqM5jXtU3w626xRaIDcSQQQNW
dK4bQxnJ4pIF/Zi4/dDO67PDt9D9FsORB0Qj/N2qg/aeZw3E1G9jLgmxwT+LND7e
Gf+sc96wsTlDpXK/vPSvNhHXV44Ol+Up0865Je8z/pwFDxuW+/viMAz3TjtnxfO3
a+eS+s1tse3jdN7sWBONJXTmeHWNH2HDOEgCQ9MPSzorqeO5vWroSDes4YipH0xr
lX5TnL9jeqoYf/Ng4GYX/0Z4V+oWm8/5XBryIUHljHhmWLDqqkrfXrZ2POkFUyqZ
BNEQuS9fANTZVe7Vp166io3UoVZCFivrnCaEdzgCVRxzXmqvWgnO73DQfKwxFWqm
eStFg5pzgjMomceOT6X+0ZNd23C1amcHg/lNvuougOeV++PwMPIVGq2wLDYH845A
8JWbiIMGQWpPT1j+2ZxrJfy+pU7z1DyrfDMkdC15ggowSiIoOxypMg+CwbPNWnUE
a8fG+UVOEhQJwhL2poRcoh+OhSxIgBiff9xr20ISwKQntFE/zN9h9auA1A1Ma0HZ
Dvd0vf+qbRPlcbp3Q4WZm8MiabSvllf9G8STzz5IF5SRWXQinAlS0IYaagdfmutI
jBKlE2RLLMDMMg8WR2++003Qm2evT5bw1CwLhe/DHvT/vVebeq59bUP7z2NT8yoM
1qcvefiCqipNK46NrXzE4d1SXYL+buhoTUro7OukqosqEoB9fe4wImlgVX1wo5qb
mL8aIsQufAl0xa0PDx9sGwymmHiGNubk9npKFU7CY9/evV/XKrOjUU6NqC/KOL8c
pc10Oa7grZEOlAhLM3FxmyDhmtr/CK2WPkVf1DSSN9rgT8chG4M8GniX4pLUJnn/
/GzQSYoaXkNfWod7l14Btdp8aXU1A7WKKWx2zWVQvxdhbooUD0yQglOHd6i78wTs
C9T+yRg7rw286IwqmmkSOSZvneiQkvcGAv1Bl5bZPptXoIWyjGFP+4Gx/Ho/5Jfx
K/nDi02iZVOej19ekvYRw7QCG0BY7gv+mUucda6wnpoT98lYcJH6jUTxnSCDdpaZ
W/hLCWvXZrPdDbSeiNcmSGAW+Oq6v445F9J2z5gDdl3RmRtiFUBvNvY1uni4UTCZ
O612qG8NxVMOkx0mCsag8sC+5U99/a3d1RB0kY0WDwUwTv0n1wYazHR0aA8op8OO
B11zb8uVtDv/wEFgxpHvuXgH9DxNcz89BiPnFtNsEkK27UgnzOQ+DPuCwhbAeczv
7aQh9JkZYJvJCF9rY4QC4L5JK1qsoPeMvtfDjE3xVrp1beebBwj2EPlxFIiUUJE1
b1OoB42xWryPZ021j/kMCseoqZx4ZwXm+2WhUWnVdJd7D1rBO98nB3ik+DgXhoNq
qB/g10Fc9QTRwDnQP7OFWCMDsg2tj42Q/LGGi9Y4r/yHjp2YwToK3mLBMwFhkYLk
9eBfu5ibEcCVuoc1NoeNbXD7s3wgKfn47+/eUepfPKkFnMqzyMLBzQ0x5/RDeTuj
oCKTVxCmDvaTwRRmh3fc01t2Lwel/kKtcZLZT7VqDwiB+OXXPcCHq8j5oKiV0hr3
6cgdqhSm/NbNAqW+4xviHIH6Mi5GihBCEDDsjdV3CKJRmabON1v9PSSZ7VKbyjrw
eBmMGtSj5bzxGccXFtgXcbmbNRdCyP8SFl36s2mtRYv3nA5fGzLG5wI4GXPqoih8
rfiR6BbBkpmCT0e38l1zZ2krr27FhuTZxM9U5zOQopj9PPZrrwPVorbEd5IYrZ19
yW4Ras8O+vHVfgHtE2577N5dTrVZzOg7HxfDA8s/Ykm9kvjdFz2VMFBg5xpkorM2
FgdQ/yWvpybmHHttoZdiL+mcPilAQVveZvGfrnQR9oVBlFhqpcG2ZcrSADJuVObY
5JICGKHFS5ENPqoA5Uw+Y37ha124QNAR2yMpR+mBpWOE8A385Hb2ZWRAybojhCm0
C06bgbVFZRg2RD1S3Q/dm8T8KgaEKvOeXxoXH9cCXsGd7UsnjePFcdq4sfZuc77q
gaTG+IbwtpQu0WE3CA6Iut19e8YOoepeEJNg++HBf1DnXTuoG72Rh1RtrSoo6Du3
iD3VlkXlzsCcYm7jP4qK7+M7Hhvab4/BbUtgiiZ8j3c5mYZyeF0k91ayAtBZVH/Q
ARlM+XXlXz1OQwwEHhAP3stXgFwR4mXh/ZEw6nOi5slpGsYTlLHQQkRvo6Neyzk2
FHa5R7ksVuLN888bF9P2qvMbjXKf6I21eqh4ynYIv9oYxEdOSFsE10vSO9cZ7qFf
W0OekrKxqV8yssOl469PwEJh4eCR7js9/CTpAQUmdiryA2cXYLL+RmhI5Dmn5YxJ
zzYEy0uoMDQFcc8hLz6n7sWrRqnMiOvVdkMEbV9iBtjAjr632atrKHllqEMH2lAF
j/5osR8xYYgGN/2AmO103ORJe3YZef+C2ooPcif+w8yq4CKRxEr1B+L+H22foYLO
3Sh7B3vF5n9tO44cjm0/5yFu/f6XBC34XBFgChz8u4rA8Rtj73p0Y5XdF+IOkOBC
MHhJMksGaSX61hKPvDKTqRkzbOYfTE1ua2lHBfe8uR4PTJ8TmCVvv9mAdI5vSn6d
47Q8nol7hMFHDMYaT23PvA5ZJtaWA/MHBiFOWwtD5yECH1qVq8V559IShKfr4T1s
LmDGfPh1KPQCJ+efJBPwQE70luN2M9ObzoagMxJBbEA96A5QEICtgNzDnwIrckk3
Kd6FUMWHroOUYni2Jp3oXRbKw9WbYtKRGCq/DL3WiifDHowKFL/MLNTkuuvYSXIw
xb+ln88XNIfQoqVPljsHBaXPZP3TPrVvDwKHKvmuHVzdok6+tMAenQFqgr5O38SQ
kmmHI5tdTHe5uHVZ45FCYxt7ZvD8Jo9KmnbJESKPhH8DxWKr6Hgk4ups7ehwzrJ6
tYfj9x+iKwunbwz3kGUo/xNJ7yDyNxCUVVRCcs5r3veZs2VdleEhQ9sOLMiUzeDz
39aB0n3QZpSCgm2BNfQYjpnxnMJ3sfQ4Nr7b49tEqgBnykShkcEu4XhwxBPZuNKM
GGVOVpGMxZ1kxFzdP4zR5u+XbFuILyGXga+w5WvXOkn5Ij4iCboCE+lnkZVe5bdm
fVVdPIXhLsS5JIIdb0eEke2wAL3bp4oxdgbD1chzLuioBICVXEQs+cPtpLklAGfO
CeAqRtIoc0vCPM3RGfCrenKYpJv3w+hX3W1LtG/scKzV1nVnF9OhvwgI/OqN5MVu
yrKMny+yx93DQlS7E/MIn6scSY5EnN3RYmDH/AZiO2EgH4jujV7elwA8EmYxyyVT
lUF2GZ0oqoZhwvgfOl0tObapkGyyrkMmF3ISF98H3BOFnCv7xYF6fyNU+fgNL3Tv
8EBQa095Mhpm03HY0QzswoOTLwaFp+OCfvkrpQ5ccrSDByR24n8sLTHhYBb35RKp
XLVaC9Opx7aWvB6hHxj0NudVLMyQERe+gkJoVrrMwloDtDGlkME6NYKVUz9L6gb7
BjJT26znMW0+iUeY1/2gAKVZ+rH8/hAvbVzo6wC6J1fUWs8CPFrttIzK/IF9Q2tV
9vzUGwKm4Y1anRUC0QIcQEmo8aseV7W1tc77tBPXhVAnm3gImZjQJk+3lBdaK5iL
I/PYea/ybxVGJovq9Y+HjjVBW83Ualg/EkkgQcgrzKjImALi6IF8DEoZqkvPnkxH
SdaOUMpFjdFA28JP/06IPPB7IbHRDdLd87IYVB7nbRQxE4laHOTwPe8O/iQr1kxf
/Yy4NdWkTd6mb0KbfkU1CX0OO8dxeDLFXCB9uJDfVk8mAGyNXIQU2doIXHfjrMGE
uTX0HKcON1eC5aoFgTaRz6IG3TH/nItrR9XXhKKbj/BTvRXFlaRvXDLZfJPTrACH
JvYPJFBCmD5Y7lIZZGQX6rtLJBZH8CXdNVhq3epkRIPfBKI1lN339814oy7rKcvc
4rBJGAPK8tfKEm7h70D1rDuJxrOZ1IPBL9Vb9Su8Q+HM6VqzBj2YV+AbHTvpEHk5
qNSwGSWdYjcZmiLz+Y1ySNkOtJqgCl08bVJ/W3GYB1bCJfHPGKcfxnx5xeA61VXB
7hN3GrYIeit5muatAQsVQtTaIB6OCZhUDlmRmJDwhth2z8dIA7GCpQwZkTNef9QK
f1cuL8m3gc25AD68d6o/umexkc7lZ3OTixMfON8ippP7Wlwg5zkR6+ERcgJLK5g4
ZDXX2Pa9G2ohXmyCKUtJ/WWeufYMGQ8xTxK/PujXxepPY8C6suf5ibdA0wchGxDT
KNSfWKzWEuwNOCQGfz4v6WtTUQHQqfzfrbfe98rv3qsdpy72B8+p9DicMXs6VZmu
ynBpl7bKS+6Fz4rnbbk7obDWrbqFrC0bL5AzQo4T96fQDz1YGwUADvDBVTM7tuCD
Ns5ljNl08osM/qZWbw/eHguU83t5WSaB6eENqbrztGoUeGM8QsbzdAZVAXJEEaYi
Ek/uArxZB8uSLi3KSB8A4DhtmznohvlNafhgG4I1nr9MwyyKfqKd0vzPWbpXaizO
DmRqcmBtboj0ZZ75YAY8RyVvamMw9MHH9hySdZ/jm+KHdNgO5YAFdd0gMx7aJ/6T
0plyCDdaDyjiJdClQfzdJn4fNn8MeRM8Fgg+1HT1wWJONWD6hN+CJH1e02VQF9Uz
ZhmaN9rhrPAYcv+h+v3XlXJDMu7uTs/o6EIJ/EoXgpV/e5FjL0wore7mk4/dzNs2
hsoFX4ktSgKI2cO5BBXRNwq4wvNyP3Xtpm3ZujF1+LIzpGRJyR/HREjaqz1SjWH1
FC4ZNe/ONjMLneN+k0kiWSg/sAxrqBnbRC6sO3OC/rgskWNB7M0Y9wcLBAa5bVQE
tdbEXjv2JqGY1MMUtSKIH/aaGnFf0RK0Eu4GaOElZAoSsKhZe+nr0uxeS37XPjxr
b35PSfbfxC7JLc5QcAlZtY+apk9PsrOFvxYPb5VgTJaBka1Zm7ZrUpYcn/B5WaaS
ATQp37Q9AUT0Hhm7RiObBSBXVGTWXI21ei9afRm6LzMHVRrq4SzznIo53BAklPg8
hYU/Dtapl562h9S1AEfo6C+bbPpHhSLq1I/7quEETA39poT3W0PToBz271dOirDs
c3zN1+tncr1dMBg9fCa1a9HKcc4EYZ7NzmozdYXyhTMKw+ZD2KTobqr+aykrH6g4
vdf3Nz2ns6Bt6gR2YzdQ5pD7SLDA062BzKFKyszx8HRWqQ+PatAO/0uWxIlD/nx7
s8H2PXv/FSa5gTLYRDu2AWQoNpWmgbRe8b5i0CZ8503RC6SFom5d/HlaCpqYDu52
Ti2eiFNxnffIeBvgGXJ9gRQnjZfhRy8Me4MsmmFmhP1cZhAAKoRxRgLrbhfd3reC
7DXdm1AnwaYNVEggPS6sJ4UNy5gpkjoOxbbJl7umT6k4fVTzJ5os2z+infRW2hf8
ALq8jd/JY95aE7PhY0Er91NjqVpd+ZFtmAa9vKZ7LD7oVw64lwyZf+9YOak2YWGU
HxHQ9tyqVIKMuHKQDnPtFQ3HupRd3Oh9/nhiEN2lNNakL+igVKS0IWhiG+3Q9Rih
ed2HydP3eUSRNY0BS6KSdpajVOtdZ8CjqAj2t2NAzw0ILwmI47peTg16oRw/ijMj
XaVL0J4/BVuueE85JJCX9WExCFylx9pIIW+RplsVAcwGJLJt4XR94jBVYcI3k0wg
dJL+KshPcvPqUbTRKABOR/WU494x5kq+a087qP5hhb3lMcG/XxRIDYYf+14s3SRC
6cVUfVBqOvax/TJBzWphAa2ndI+rFFcf10I03d5Jrf3MD8JeIWrXle89yuksa5ow
1/lAa1Ob5qsKJ7ud8KKkqrmY+2E7GAsLjh7pYMc2K5mlThTqPjmxAr18dJyVJFvH
6XSj2fufWKO/UCR+aSOFTNPBga+0cvml9YavUGstkRMIV5oTGePPp2V2sU2AgA4A
T3uYrevxYl42cj7IXOCjun98qtpGAQrwN+U1a0uca9vK3IH0+nhFWED14E1ITrVU
r6Mq+1mMPN3uzOZ9mTbUEmgc01QeJ2EGDqlVvGa9qw7Vix6vAFOmKGuJFfjVln2d
QEVoczt6yhT367Qow3Lgi2wgHvzIR6btjs/5fKBZIVBeykBeamVH6FxCzi83oUNB
LTAsRYD56mJexfZTbxiNuZycBHiG2Ctr7iz9N/WtOAX/TdlAV2WeD6Cl/W+gTksn
UOmxZuo1eKP0Ku3MeLGBUOm6UTSSaEZ663R1uji27Mrv9CtLHO5RiJe3qOxUxgH2
OwFjOWj8JJ0g21n/RT3Rne8AOUKoxFfMByzEajqp0537WkrDvsTNXZqzg9O/JUUn
m8T4fsC8qzcjwl70HFaq+pGkPMsI+Ythud/b/T2kiAYrTD2rQ5agq4xMU5RnuZlt
pRERU4YK/s56ICKUTelb5vULhAGMnnaEzJ/GLucRDNLcjVtZXGyl33YKPbIMaYDr
k9GeVrSJjaJWdxATVVwrcxAUbJ7O6NkpFSi21ZBX/vWJdSpKVfW84xE51yyI3i1j
lNimLXpkEAICPXdqt4yWbpfkKPB769LPUQ26BuD6kxlDZ8qgRrQ6Qsu1Oi0OLCYo
dZkK0nUuBbgg/bKJ9JEb+rS0eKvTvdf7umRR51u1jxLeohfXUtGY5ztEeXTKL9n4
pz0KHjXCkQTjUyYP7iXpf9gut5S4s6LpQfXbbsc5bAnQPPXWh4Yf8isidxQgIls/
n1DbA7bUvehPpozXMNf+EJAC590Uwoqu+yqzo1e556Y/ou1AEBxTigNXcEUfbipc
X3p4NQDhI12nW0YcZAWzAuMkskNMwnfpsHdVqW6bhIEqRoRbHFrPAKsAN9uQg/kQ
CeR9123u6TJlG27jSz9N5mNQb+2Dlr6v9islqO8MMoyoqLbH3mHlMOpLHvGlTnFz
Af1aOy+dYfU0MnAgdEsxkpuMhG2ZZbELrQkVpD+m/PdBQPj+Q9KgnZCuJXJSzNr7
qLWAz+6PvVJqmXc/+rWPFHKv0YeHqGl8QtCwHTnfLg4eQQ4cJm3mZoODa7R6vG56
yi0V6zHT9Gn8T9J8kaNUVOUJAojPmF4XRZP4Jc/LM55Hk72yAtip9JvLIoV2ERFf
01I/13yq5YlZBxdgiBYVvLiP/CBVoRpaDMrU3jTc7YSaMYorzcUA1ZVdkmOBTu2i
8Xbeqp3FT6RVtRhssHkcl9uVOLdVO5VNCOkQ4HOQMa2vq+paQL/qlXVKaVpBg3se
XXrosDNe9+z5NBPiKwZRENHh0wG9UsB+GSnz5z56w1OFEZQWvGWIi2c+CRHW+Ie1
IsvlAGpYEYpEv4QyshXItbku0S0cZ/rqDn2X8s0u189OnipGdTI3G/gyvwk6GYgo
bndWDwAvxtp3IGpVBM6fO1zSSji66tAW87UCW9nrnQhztErvb9ldV9lS3E2MB5SP
a0NwCxR+CLcHgHcmR0h/iLESspxQ9qpBenf6cX35YUsKTZTkOqjkkfvLt0+dPIBX
pfmxDYWQNmdh2gqMARbn5FOzA311CzrCOIOOVPOkrr27qaIitp3o8PCVKXnt+xAa
kp1ZRDN2xsZL5ZX0zRMzOZpa1Sij5I8x6VHeIzIu0yrYpuPzjpnfUr8Z885scktY
iwE+PqxaETC5WIEVFl3ImuV/iPsa8lctx7auVT0Cr625s9SoJ5YsaTMB7FzQ7Qyy
3nO09c8GIBAVv1n1qjfCybONCZqhva1HZlKhnAyBxD4hq7UAHBc9cbmexYVxZJBP
UOhQZL5dXdC/nasVxRT6QndrCE06uDqJsVjIWfYmiHJMYIr4NjjkLbvaKQtC3ZC7
lOVYOUxyuNgl2q5rmgt+n/yWwuxhv0vBwne7ONlWE2cw5ywBpOUuJF86MLSBCSum
jsjr4usyK/DCjmHMX1siqBdnNGqE3lmcsnjnkyToudHtQ7T4Tc8J4FJ5UjWyC4ET
q+gYZxdaV8mZiOkOEPeclE1T01aSPSXWWxHduCFDbmY7HAee9QnzhbYV0F7gcbqD
3OQ15hJ5jv5I1M4d9WiqqWyYdy4ukFkr1jBkf1+OYPn+sjAv7OMAR+68tvPsrnTA
iar4JZEuNI6dzGKBosshhPUkuHhhESn8YfkftaNRtRNTWN4lQWeseeieitEaioVQ
QYw+9JR7dI/IkrCTnzkVvxqYOAh+vdW/gu70KarZg1kr2T+S+zajhfK/q5WUArRO
LzfJ5dG+0uO0kgHqBx2HxjcW6/drC/OLPXlMroLkLnPV1dGXndQGbmUN6tK5Apti
HDy9YP9wrl8s9IJHomW2t96DO6te83vTiaW6FgyR7/ckwzbL9hQrwgyj9boMHgLu
MBY8i3EwT5TtdTNNXxW3lQZWtx6QCcILTZSZFXTE7CcMy9rdkIz+9rjuOoZQH8Lj
PvDrz2H+sMQan4jae+FG1x3M+67XU4HcEnPIUSfxxPZ6YZqup8PnLu+ojElLfl7m
lfESdZM7n6Uv4xtVIkNm8/Sr2ztZQ9azu02BokoaywSax7yz2IS6+nVmLyKa9szn
KrmctPF6Zh1RmLlZkR+gTYxKyuuUWcj8PXEID44WM4APB4Nf7zxDU2eyWa9eJ/Sk
YFOp6HoKmkQh0J9XUcwZERQh0UbMyGpPJkpV7z/73C+oYxxEDZGVhLgsGGK4RQb6
vJCEq+olrhyx/xLra3DflLs7mIGrMjkfQu7eUgZV9k9Uo2hPucdAg/NI5bSEzps1
fAytwGbgoJMvkP15vHpDSVFE5wlRqSAaFsc5W8BUepq2Gb7N6Hg82aNrzgSwPqkQ
i0D0+83BjFkdjvzCvcevxJeH+2phWQZ5yQfyPv12gLjjBCB3Tz9E2RuRN0hLp7Cw
AQOgGkujGOoQdh11GVT/z34HrAbwYwalvJ0x8XIzU6BdLfaUFmEn3e9K1E2FFf5S
4vxfoz2ynZHWVcksO7CLozER0/q0O8ZqRjyqeRXp/EwryXLLZFoLkZPYTMwB0tkk
7oPjtgXRUYaojtuUmzaV+RISvhEzApUI2o38gn2Ewt3hFJ5f0WZJTWrHSzEC5AKt
3o5IIApUv3sxvKwSIj5sx4s3j03gOiUcqiM+7LoeMx2PqTlYGpWIhD422TznkHl/
/lQzRzmOMN0Vl4B8oiW4WfZf0nFXVoIirpYPW8s4NBP3JK7Hh+WTvndkcz5tQBRG
1cDFcqKfzGITR+sAeeCP8uS+bzB1V9YxvRcnmUgT+HYUDYKZOKJRC1QZQzOee4LQ
0055Ga7o0Sg3KPIe/De0hkBjbIyqTGhv79IWzQs5g/CDF5o2GofnL5vr0ynPd1BN
1en4iqymCtQ+bHIgJkGegonApdAuLCiKAudZNmGIPp34efdQU3LsEKBVHzPAXK6f
5eJpTzR0suG5fcHx1juMWyXo3DPYgTEHyN7khA+/oVn+VZT+wvsYeN2+kKQQUEaa
zZilBxz8G4Rl8NcFOYMgh83TbIHUU66kn+Gl+APfiDRhbQ6uahUvbMm+HlN/vqt0
zUavjMZdWvKnibmoKpUoWKRWGtGG7ztJScV0XAbCYX6mQ78Q8ih6v6E45/UzchB/
PImXu4FhitSkIqs9Bd/HV4RGT6oWXhPxW61fP4z+ex1RxO7RjGHf2Z/RBnOMCwS0
0yErTSfGM5gHxNFiOoq954bA9ad94/hB/JaUB+lzANGhQEq+oYVuDyvsxXegEXhz
6d85sJ5EsOydwCQwQ6UhDE606aKcoFq276uliWnMUNQUzdvQsH5wmHK6Gv9Rswh2
nycmnW5J84cYjfLatw9R7ckrzSK1KK31rDDo3fSr0liD6Z6j2qbbX5Xx5kbw/0im
xlbXK4FfYBL2dI5TK/TqhlVMyAR+XmkVfi7dSXdKoq/8dV0u/JWl2ryiY0U7ZYn6
26gKkynavVsefGlDu1A1zuvYagt2eY4j9D6ZM4xULHZyFZhJYG5Wc6M1Z4xvCP7V
u7vo+TS+i2gBFgTwkJQMjv0Yb0TCJdM9RSGbhuI81PSlMEZ9HZiPW4BS9flPhXtl
8BjJ704hI6HIUc7/ysqEWXUQ1YByMGQtCZHJamaR1rdbXbgcKpv+ndpJEfiSVCXv
rxhl9/lIp8xjSrT63xLH7crd9LrBDCVOJeuQ0Y/C/nklYVFHsx7sH6lgI8A1cOYS
BTgJohONrm0Pi+Wtk3qQbAYK7XSY04TpYna32Ypj76VT257jbP0FjaPd5FC7rp86
Ixt2jP+gGC7vj2D7Z1ATiqV6LkaluhnLvbaYvNjOfZfW+zWFXSUV4RsoNlXp2Bbv
lR4Jfxe3wHUsRNCA+YKnJ4j4anXnwPS05/FU/NNE2bNfQAm7XrVskXV62vT7ioKD
Roj66duNci/upzG9TL3mqeCFJCKysD7OOJu4Y2hmMWoWPmsO+yIiBi8++FP1SYbI
Wv0EYQiHf1GdjaavB97VeATBLBOHqbur9yzBhhT94UnMiyhQY+e0nLbs5wmYNCzN
JraldCxuUZ+qD4p8N0tTAoZSPmASDwt6I44yYka+f2LV/4WEs4JJfizLc7+7kWOq
7dGpKhJUx1iPbXzPkPPUOk1tyYJ1L6Byzm4pxNfaA+gcMVM0tzGp1hpQH+Wx5fvw
SYGa+YL2WCTim6vQ5/Z8oqqHZjYdyUZ/IoT/BwyQ5B1jQmWVjPbjn4QthArzBQOT
8xKTELoJDZT91ALTtBrtCqYJJGQjScnzKcWuUisLVdoS7aaelmQt/+fBfleeNwg/
YXXw06oBkfNN4tc6v1W7aQE9BAGG6gvDUeIdowtpkNdRbBuBP+qr9JzGArQoRysq
ZzeoSuHRSnWOMJ+2Z6oglK+O7eYcyQinecVh1lt8yT+V0WKGqo5g0vRV1ba3eG93
RN/nggfJYd4LNwJn4ftSy3pZwl/DfD6HrWq7T480uGqG/DTNjvGAQ7gmQWdMfKzL
+IEl4IEdRnMZe74jKuhcsf1vVZktM/2xoFR5UJC28pPxcvlFEjsrNETnRvSjeOKx
l6GH3HfsVidt/OAlFbnQx00gWM2zX/TxtW9sYXRyoyCxnrg1G/oxZlLRHCrtGNuC
80I31EqMeoRhgCtRlegsnJGOihTpWEv10F9WdDPcX8ipzAHw0j7YBJ7/n6MbVaVc
vW2q6eDBENsENXvUkho9XIOYonz/sk3TcT4HtYsITTEeJSl7uN1sucNS0hgZswKu
6OQsujV4PK3FajVw4q9Yf4MRBCbft6idUErrDrJgs+v6BRtPOFd8wNfUL9nw8Hpy
cNp+sOmitBQ/tfOu1K6R+8qDysYbo2wxVk9SEah/c49iTUOKfOWQsBpQ8RLpELOi
4IwpOTYy1qXkyXDWDDgnO1mdYu6ODhLBsoQJR7QPKRe8fT+xsu47IyQQyotybAl3
XpAHQvUFf6k6sOknvw20XYPk3CxdSdiS43cA48uvApwbEikxSHD8IU9fbhdgk3Pl
9zfUhB4/WZXWQ1TFVcj6wiJ5tVYqELmA88NJNgOPCPih+zDFfnIIUCyv2KuIuM/9
bkwFQ6v1DJ1G0C7tuevijUkZ4KEqHnnKWcVJDsKsYfDBMDtUJxjVYxrDZbINJVNr
sKZkhTZlDuEOZ51P2Niu1zepaTs14521KFHy9dZ3K/L92w5+5x0t+oRG/F8J2VGf
hOR8SLa6CrOES9hEti1UOyMvtGatgH/AY25Boi7jgVtI4Q719kVWsirXedfHOBWS
Y14jz6xtISAjnmcNQDkZPI2mKrw6UUZNuopizXhj+zEw9Wv3c8F+RI0ohdEYgVXz
EHKdTugtFuhHtCxDbPoiElvsJ/R0qNT9WYA/JnZO8R4WVXv0/yzezyg4VMRJvhUU
OnHrsw4EtSm+fTOT0ptmO98FBWb5koGSXo3HIiwjA2+OlsuNyqva7Ku0LaeZXo3K
Nn0fLiBYvvcIJKd/xyBQjxAoanX34igEd9NhkhRI3roxd2FyEDbu0woCEimDTsud
in6YGq7FIkGlWnwuOQ30qKl8H3X+zs6Mfi2eervQW6vhgeeDVnb4YvASFpOmSuca
j7satAUWPgECLtIiOrbW4rlHa1XQysZQBoTA3jcT/0NqkGeYdasRPRLPRPcAbp4k
Ew7ZNEC+RuTjOxbxAZM9ZLrVkAiW3xLuldx8cagkDFVLmgrri8j4hTW7kylWm8DT
UVxL7t6n43KzNqTy/6j41nKkTd8TSAjhHOA7m+inlh4NFMIZpZ6VGTMF74I/EXnl
eZDTbXyRXENxru0+dpsRuqL2oBV5B82VDo7N7qZcTvH+WGT9dVigLXKLg9NM8O7C
lk9/JeV9/VlWCzjDmBhpIHSx3PrDEqEA0dPvTwX2Xo4n/8d8m38RfC0mmU3tIbe/
MM3xOzvMa/zWNRzjjpqotT2Xa1r8mgYI/NsO/bClyo4j+Pame3ysz99kzlGpH6KP
q3+lIiXFySRPiKmYwIgrT02uHwNSjcKCYhLj9JuRmS4/hH1Gwk9CPkPmRlWZT3J1
Rf0yt1H5EanIpbfkGg9dVhzgzFfrcCkYeJgMtY+ieT0wQ9SbmvE5UE7YZ+AFf4Gi
WTYn8opLFgPstKMErgor0rfKtR59MWgdefGHgcXvI9fLtyR/eh1yV1cxbJyTl2VY
eHjwIGHY7jHUFHQyhXwZrl74mqCgqBOHGJwJ3WiIyT0XCbbfGsnUhvAU7WrCjwvW
4FjCwLt4re7IgxcqZMeg5Bv+JXkMQDNP6obgvfdFf2gLBLCEahfHeWW6VomdqQKh
CwESURpW1a8ZHHR3VQGIEpkos38po9yl1drrxaEPQwrG8MnuxxL8AQqw9nTi6M3X
YqzyZ476F6cchja51KaQa8W0KebNtZ0KNp7HRNAHgP1OjnjWei+RuWBvZlXz+KvB
JeEUHhakTkx7T3UaWEHD1BVKXumcEQcA9KgVAGX6j3mmxEIK0ErRRz6IrEDeD0TS
7tQ366D5iWvVi/3Gjv1IyW/gdQH2q34sKgvfnPAvV6xT29L5IIOkt0NiuRsGI4Oq
kOKaAxhqEQB1MMvW468LhIZnDj8rI6WJ3/ZV/Bia+yhNvBbe4XAfSKSaS8ftDBYs
WflSDJAws3w0kP76iiH18SIGmTh0bhMODDPvHdt35mzCxLngjm8MO/mJw0eyfC7T
IW9YXUlWooPwQcoUSzBTfupMpGRVPlTaUZvAT+TukcB5RrSBeobAQXA3b0v/tK7d
YuQxfAnM0gK9One14W2N4OlAFZK6MoGe+/0eQOCqhWBa6wlZuUEgGYhTthpkG2b3
mGlNoelVbDO2vYt/mP7KhFedX/gkKSxDHAeAYUEhkKRwGH5d2iRZa6AGGd4zq/D3
Hz4lAzo3e1A1ZZtR4GHGylR1n+8lXazBUwNwf2La9aZFxoo88gQR+pW0tCYf1LKo
1p6WAdPdXfQ0eQT6ngPIoUfHVDJdN3SLBqE0GaD11L6f4LoGGJTCBENezxMa/H2q
MdnVQUuYcGMxsfItvn07QpB7/vtnYAkoFYdGpDrsruWK3FqAHE+I6aGtiRM4tWAY
Ok7CNRv+VDtQY4N+GE0A/CfobtWBO4N03MyoW0idKmE+mgCSiaRtzur24D9LnBjS
2ZEH8i8inXf5MdyP3QtprXCSqUlDxGNfEu7QEX5cpXmrjROFTPW8zqw8AKSD7WCy
Z7qXWtLcVFbxQZ0fQwmvgx3mFFGPjcNPnjNbEKpXH+0y1WEOvYm2asQPsC1/YT6g
WBxhtOhQLVOr+l6C5hTjHqmYt9Li/EhPZjUTJ4Z0n3mM3LoI+Z6mAZ1rx2OsEsNB
gL+DpLctfqJvZJWgjV1EKB+vlZUjhqMQ6U0kAmHdLxYC6bIXw0KIPw7l7nIrjUGD
Sbguf240ZRc7ZfkYJkms5mu3IyBXYzy0yG58TtgaUkvo+J5B0MifiEKIkmsd9Qd4
GaBGYm0xiYVzkz/8JJMi+p1rNNtCa1pmnj1mtWb6PTz1rJYpmYMMkG+Iy00FvbGW
iPh2iPzA65MxWX4cMeZ/36WvwbJplKXLI+3r9ZBUwghA4EkO8v2YoBUDn3GbH91c
6YBAykA9eyiSBVbbmVGdXcnqmZO0dO31rkj9hGP2skvhXS3lDDY7G+jGT9ersyC0
QVmnDNnKYiGOqLFJS2Tbalwt6DXUz1lwIv4ee4WZFuCI7d85OY5OaKmnCE30aJn0
/FDLeqz8HgBFqoVm1PAY1V0cuJjbQZpmmbJ4k2a5itIwa9E1MZhory8/vmJOXRfF
8KoSlujCbqAjIXp4zGJI7DdMUadxqBjV6V1Slvf71488W2//QhKu7Ly9UUf6kcYE
CXUH57gPlARj4lcnZte+/ynIbzghewE+pRjgbhhI4vsmeB2C2Wu79E0HPckdIyyt
lMPv4l1ANIb7Yd7BUa98z8Vm6e8rLtIGZQNy1YEH34xcIG3imOdo6dOBCsRP+TNy
sQdOy7cWKixfgU8sEBfsLGZzAsHjapfDkzZpwj6q0Yb655Kg9fnXaSB5izHyg7YJ
HsWHsNGaAjt4sZRg6tcEHO5WoHBS1hhxcwJ8FgvU/sGZsP5uZwOu7L5uXJmRLw13
YNI98nYa3ka9haovNnwpWzhsQfNID39ns6Eav/wbbPmhziKika6hI9p3KxEW+b7t
5Uqr6pzEDZQtYcmXqINpOcNMEFrMn9q1YYhZsa/1f6qMa0RTIl/nYPkNQktQdLVK
jIHupdFpPrfC2qAuxxO0lB4BFc/goNR+LficZ6meu/8bvsarR8YddTVtfmxbJdUH
ULMkluZ7z5wqEuRHZOBR5qJbVjXkqrVr/aVHgRxjLQI9ldS8Lb8VIepCRrmw0KTA
LSLJgTHINqxrcNZS04uzVFcauwSbkrRPwIedgRXayxe4InaQLKVmMAX1MgHvyVaD
2M8mgViKxD43gdXYHms6wTXzspQga1ZZDR+8p1KTTbuOIWYmR2rjMbD3qfRCbx/s
N8JgwrrYB3lp8rH6TmPYLy5Nf8HSPRnxlK4d2I1j4k/kGHCTajyW6EfvjR1Xg5MW
KFpVhWqS80cMflWcRt7V8Oh3jlip5ZK9ol6hklEColGTFrKtvTitetDMYhfjDd/P
ufpZrqDWIEZavPInLGgNs7tYA69kAwgLBjRLIhrVyUFv5K6vP8sf8Slwpy4quuwj
tdyfOGB+4fDVQzFLN9PX2GgPwxXyr2DnpnvMKLkQws8yY8bkoDbg/TsF8uo635b1
w5RDIqhXx9JPmOlb8TN+GZ/pFnKZLlEDqH3Ix6xY4Gcg5tok4avdLpdHKAqpwwCu
2gydCwDSiRel6Id1eQGB23Kz0KX+zrAWfC0qrGFbMszNbh0ywO/2O1rYb5EJctCC
N7z5WtLAIiPzBtI9OqIL0VqUkmlpJbgttcrklMBOJVKoEU+bvHE6GoJKHJbgkcfX
bEmcCZzJwnmXsItnNqcSre7X1ufKl1LF0hW4B89LDjj4VXjBfIpMZ48yTDTd89mn
QxzeoIZ2wJ8wRSubv7JEOo+2BDtEkOSezqsGCtfCvdX+kdM/gcCZbWSAHWyb7aBn
K1wZeEbwA8MgKzKpVHuQO7/uGI/5F87VqXgjYZQPm+v35OyWoEoqL+cgc/3UXKY/
COfnV6+XwpskFZrnFMRMn4fBr5EyxWsq7jjnCJ1UHjMttt8bCl+QRXcsE/gb2B0U
p+PmJFevDjcy7MDsGqZeHJx/QRVW1VBn/MjlwMPo/R0WIgxxuY1KQViUX4h2a3au
OCOT2riJ7F0FBrYJvCPAijOzgSEy33+hKCDUNz3jEXpKZPe/Ux6KEv2h4OYRd5x4
5hcxLDE5x35pbVNjxwtsVs839n0Yk06Wbl3FAttYR/x5//8mOVMOcvVnfHZJ0Bpp
zlwMyu/vCh18gnLwSTigb2iizWv3NWeY3o/u9EitQVS1FnEllwGGga869lGO+S+D
nkF/98XMNO2NwD4EL28/IxOjByKABuMkkCgwnJZXKhqJgLbESiWLazdwIMSuJSMZ
dg2JeHEagSOtxaBQte3QgsdJjzWjrefUKOQfkHhRrU0xcaeYfpwdNBsAe0NSx0nF
0XB+GD6/qVR9RjGtpoOuN+fNm8lVlLOuemXtz2F+XCzokA20zP3Vo9KtoGgheU5D
Coqnzqj4qS8kgYAyL3V8Ik5tc3mfmjbGZ/qq8zqsrNbNpvdG81LQlKx+kXxbs78r
1vl73KSuX7gypNho1GVqi/WeAoGPvzzXQKmNkZ5e/QtpKEKZxUhkmbbPxmRjFKWJ
otjk90bNpNxNFRqmmtGTRXDgSQ0WUT5yRytXtzejAPJbYqGCWCrqHTMjFfptB2nR
uW3aY8rAJrJ7si1N/ZgCswFtMi3K/iESl8xIaRjJAu1tAFylCR6GnsiIkPagygqQ
HjArPCrKXkpnIi5Tvm2mM6gnFY+E6LsJsxxcH4RaMosF9sWdIjsPUl+5ajAsDCJ9
g/pzNxc9M0x/WXXntORjXeKaAipy99sFzsIPikddSz73XzhZxFORJS7dE/2g5A8w
7/gh84Gl7g0h/s1y6fXeEnTX7fmMSt22AMA0Y1ivwiWEFI7NbbEtNAa5Qi094ULY
ipjhiHYm+Qp83dhnFE/vYOe05L3nSBJCeBjCPuthIl+8dx6ncLvm4YvFDfYVRhB3
/x/k5zke2uZH6EskCZaYs5p0MJci/LSPX7vtwMihxHXKy62rnK/te7585aw+vORd
ZUGAIlWqGWYpKj1KiAIF3imyqBf/Sm4yzXQ+3xNLbdiVGyx3mSfQc65FMwmfRr9k
YRhHwqVsV1H6DJdAxKJeFMiqUTey+5z1Tign8m9iKlRMtsD/QapX8FpNT+Bc2Rj3
q8GUWFFsuHQHLXKOP/asxnmnbk709G9izsrIZp+k/OnNT08zvfTOO5P3utMcAS5c
4o/GzvW4MrcdAvIX9TacKKPm5aJLZwxIHxny/2W+YcKtux1THcBzka2gJyUC/lxx
oTnUkGJUt4eEv8lSnxQdihvApHs0QUahAzYYPntPbkUpqj4gGMTYIYY5VwxLvAvw
K8Jg4gavCcthOprYWul9I7FP190lVwQXcdC9xUFlYoAfcYVGaiWMK/0+rgDoXlR9
X7OXhayBs5e4+vwOvQE2znZ5cfWTAoRq0xv4wTFmNyPbj+50hdXTMzO698p8f4Wi
qM7ZyQ3LUYer+bN2CY+zhcQIYFUnFd5Ycsh6IuhFEiTKJ7mO8LRcrDBQgedShP+J
zW1rmB30lhRndvC2z4Tcv9r3bXyhIgt6yoEjDNVkELISPIWaoVV+ZKnPBK1BIHHV
k4Mw/z2vIydzS0jqhK+Vj2BEwklWLeP+cClKIdRwzPSAIxBw6es9/1tdTSjrSWsh
W/BpJNOJHFdKdjN6YlT6VQgK8gmUDG4LzMVvV6tlUeyJEMOD249/VwItcILSpFZO
P/tQjgq0JXOJWm0PCDa3gteVMSvwxaPYOWrIAH8fu7+82j4VlE1SewFvEiQX5/TP
m2b70ahI4NVSTp6ro/nOiG3u+vLMzkY8QQNQ2PZXGjYbBwdiv+ZY8LvbqmffQA1n
mkHDPPhdNkSDC8EWwFObl/seWgeefjjFR7L1QQWO6EUqogJN/gZCv1aUOgfr2m9l
XvB0vA59xcENNakIhk3v7YL+6IXEmbuRqBxKCAe3uaipWti+82OBFDsEhkCzWKJl
ncsSLhKhV2YEAMPsmUL4GMPfsiKfCHPDme5lPd8sk8Po3lSp0+xus7EeXi3PTZ8B
AOzpem1BrxF3ZxnHc7N4kXyjgFJqJ/nPUhVNqnnR9g0qDSyumGz5ZRKJUlbqk9ga
wQfcTtUBBFZxy7BwIMZCWHu3j1YyP4BPuokxetH5PZRzoidUNUbfhu8txaqpNsJc
n0cvZbKZuXiHdNaIYpB1Kr8KSWdPP9i4xoQ0R8LEuV4ecLf+umvYJidkoyntnn/0
gVhaTiyxEq5t+NpF1nAjm7d0DcdLLR7uZo3EBdnZJqRwWHZiiNNuOpG9W4CSyHjj
8H4rHXd/iCAjqz1HC+h8EZ1EGFhj7Xg/VRA26ddkYeRp/5qHRKtXNvpUx6zyI/uk
ao5BJyorN0wgHq3U+Yhtc8+hkXqxKctf+0iXGai1MwMP7hcgyhQpOtgz11DqOz3E
JExOZtV0SRgcTqkh5BsRrB3RSbr8opSZxW/KcDAitVDtH2FpfVwzIOiXC2PCwhOk
6Ryl/5sr/65nsB5KxABb7eVTs6yU7lRNTeYQ1HtFgGZDgJunAZbcqyBfQBOHS964
ak0CvTcSQqe+AZBolzaJsiqWWjvHbFhMtvZIZH6tpLtMNLlruvN023Bm8jI8A8ZE
iqW7CBEZRpVcueD9T/y2+sKt8wUbI3Z7s1BDzqw7k89Q5lGz6+NFq/Vs7bhqZpTc
ETVepm5948WibT84OeIovKIELZuwJ7D2LFvm17E5wOg7imdUWZ2YLZNz8vmFA9Us
Gh5ck2AvZ825pdO7YLUdkGKfqVliB4tVdrSlnYJyFADzCqvJneYVh1d6MLyOw/92
PR2c9FvxITGonh03w9s5lUXCfAJtuv+gpEv3diUDR4ehK73SqPYi22fDgLjIJenL
W6trKgV0K6Yv3CuL951dv8SmAWTRS6XBQQrLJg0hhBFsuA0t4kcrNdy1e/o8/TAY
YTdpu4sogWchf2pYzDez9u58t2DP+pUKn1XRPpjP40lgUEUYrJoFpk8FOfA8ViEA
FYrwFKbP/jPFJ+BVxrT+eA0IPNWTH/64nWo1+wUuCVvSprtJiA+mFxaAFK2RgOOI
nuEaWSMdk7nG88BcrUg3VSTqnLpPexoidPHuTGT52ImKrNM39jh5H4+Nm4NcuXOY
FhSiazUYS+8iKNLnIx1QZP7cK+nSvFO7T+M7EEDMZOOh3xyJ+euwNgtx3eYT4o1f
XVDlsL9t7Ojv8jv3K+xoC+JG4ebaJn3UMHEailbCRy+JiUQNwAvKZdGMyLs/cEiW
JMJm+SGO0bs+Q1nuVt60FzKS2/PVeAAW7QyDR83wweeR/8z/KeOFKQ2iFcMy8M5c
csNmS2c0daa+TdSLPipKgRYeAJrAHgO7vLVA/H3sHCI5mmqof4xZGxg+A3SkhNQp
OPAKv6vf8TIBhpoBf3EgI51ep7A6KgUYnHy8b/wzsU5+mZaKQufKRDfiRj8y/fGv
dNUww9RVuDr/BJnuXJsxbiQlrM97SZe2J392EGsX8Dzz0LhmFkY6x+Q4+u3eAFwo
3DQ/y66h5+Skoz0DLV4EUEMnBFVrqgo7ERrwqux1a+YRm5vICitUhD8uKdD41Sbh
8wSCpk3Jo72SxndpclWldUzUtuleYG/ApL5HyfwvMR/yus3u7DZgTn4O8A3FPgPZ
KIKEKcP0AZ260uDonz90cP4QXcMQ/TPQ6CEB1bFBPR37x+/7c0+eG7xxj/tEfplT
6nlmZ37xW+007890TJtipaCByB3KaZByJ+ZQ8j+WqZrto2ASdWd/oqG2kLn4Wjwj
yIHqNLBsO/BpQKe5qhIcaluPzjnj5eP05BkCyHB5445tJ5/c5DyB+op5JrHQ9SSf
2Eqp7Bszmjmt/eSs59QyVZY/6n7M7SDD4SqO3SysAxnGuxPpQQ3zTlv/Ma4gr1s+
1FDdwpXaxeEKtV4iDUqvuOChz80bvs1KJcauv4d+2wYW8dNI+6Cd9MyI1YtukqFY
E7VnHje3k8djPM3nzbPcsvBLnPz2ZYvO6vX6vh781cQ4J1Ao0haWo4e5YjvCfQei
lSqVfieGYBh8q5onOwGsQkSQoq5+eRpkVZ4tGcGjiF697vcuWXxJKiQzkYcP84tR
+7YqrP9RiGYLgcLsmeX6ZLcWgDakfTzljBFaLIRtm92D8E4zdRazoVbCaPlEKU5u
+07fNuml2zI4GmnzEVOow1GWClsD5aeGoOlm6s9HfjAeD+42f/PaWCRKSWuv2fnr
vcILGlzAWELW2dy+NlFxkNC8eR2g+KnqDqvz8lq5dsYxjY1tu6fmKUQYF4HgdIXU
a4cdkwaImaBHaQ4FkKhJ9x4KuMHKXm578mRwk+GwrtTAawC/vKifiseqU/BgWSpR
JHJ5oGxaQ2gNp2I30CHSE6ZoBf9IDkzn6fIaiB46BH6/+JsXdqgO36BWjPKva7Ox
9YhHZPgnXQunmawDkaXyBczcUs7Ghlyhi1ptD49wJzMDpt0hD9viMQom0q29rhp0
ML85xEV+/tvGta5DfU4nJRNm6TIIRjvOcxViQVpzQ7NSyR8sQjku++DIPsUOkP4a
YeLtQ23m76HRES13nYNsLV7nGT+Bu6j0TU0Kjo0wmMtVL0zlhDkJsWzk0x9cDe41
48mf+oCQ8DA4+X1xcENTS7KMTyIucB26uyYuQi8IxdF2DJAM+im8N/LUG+2hS5Jg
FMz7XYNSvdGCvyxAO4KoFLBeN0oFGSqKL/NMHr1+9eJp7LcekadZLZQJS8btLqEl
//dAlOTUDCtNQZiNLS7TRNCxZN3wwSGcP52Y86h6B13c7fGbk/8MYGdifs1lz+Xu
kflFshOyFjjehCCcrWM0kMvHOVvw6Ng/Gy/N6N1ynHr4B/K1f0V7ADW4TU4O1n9C
v4vu8CzO4ZqfbogWXkNxJ7rMusdpWvFYM/SwJItqUEZwjqYBZWqe9cc7QOVN/tlg
OGaVVtoZM2rxSJ056wtGAAy0JngSqbluBcP1/H13hkTXTfTtnRKuZ2SgiFIPPntu
/ycFrPjG+cV4MmIChFVtEjkNKu/iPin7UAp5gAlRt35Nwed3DAPLuxpRs9vUEk/I
/W34oW++MMbkCULtN/ExKNHUKFQtlDuMNr6BwQAfvyLguR4VAR8itdJiOIGLWgpa
uVuQ90jvx5btN88K8mbh2i8lTmAe8tEHijzeJCJfl1QZFV4+5qrvgXvk4dYQIQxE
mYRmHXXh0V5UpKKv64/YUMLS1qynKerDEOc076lgWip90THEU16inKuppZ3/9Qlb
xhoggapdj2aK7HkVyr3TWE7jKnwGzCzv7Xx+wuAwZCgFTIFhQ9iQ4EH2IhyaF7G5
NFxB+qsAy8JKx8xsz11O56QN0sg/tjy+qzPQgEFw6LfDn3javsjA++a5cAvdb1Se
XvK1/zTRhENlzK1t6Ceo0cHB/68P8OCgqCYDqaKTkNXfXSyq8iRUNV/+OkolerGD
/MZ2Ikm6ixlpZf+CNQ9sTnTkHuk+8u5CN0lrHve9fCz/5Q+0MX84uekZ8PVrc1kQ
hSjnpsh8WqwYAGPyg8qU1AtGxFhjLKOtfvRzllMwTNlGtVSumHovyY/MujD5f4ou
voGstZDnGqh9ztqn/I8zoNrXIMIoIiTTkzDMJx4QRmB0XVtgxuiPoMRv4qt5rozq
E+TiIs/NI4VgPmz/fA3a4lvY2cVp6bBwUwOxprP/HukJT0EtGr0wIUy+T5KFVvDb
s+0iyQqHwQG17Sk+K7AKx5+1Tyh2fhLMMRNCJTCwTFHEQqpK5CXfD+rIySLcblq9
1aX1I7YInEiDQ1Uq9GsVybMBDOb95TOEbG978bMK64iIa2bHGgO4CxuIKhQsmD0M
wSENg7jYOifmF1lfJM0Sd3pJtIz/Vw6JDHv6SZP+gFZpNMp/8cLU8wnoQ8Xc7Xa5
JHgoIv+Hvh806OhZ8VmYL680BrhAxWJAcrsfj9gOtlDfE145kpR9oWD/IFAKuE+4
+8j5cts2YTID8aMubwWsAUn9M/KiN9U/mVi63b42Q9hg/NxEEObeQhzMRt+4HrJn
OYfWMaVJ1bABXLqdQ5UbL1QHjPf1E6iBp0EfU22nItZGI9w34UQm9wzDLpa5JWr9
Z58Sz4J+l8am+2cBumGVd32Ip+pMqqnOPkKU9R49dtrsJpBCGIZWHi0ms5wnFgpF
mjQYtq5vkGKMJv/kPufPKWCpcV1iph1xSSkYmK0D2Nx6pqIRVvHWG28FHXVaLXKJ
+413BDNVCMeh2Pt/KP00WSVtjZJrMLBwgazwtHc760aEv04yCfg2WwUdyB8EkSZv
ktXSr8FLDsNFwa3m5OpWtdHaVPVEs79Qt+FiBhsgoj35amaJkFG5aKgOOfSb+yDw
4q0c2rxrgJbRWcxqi/sAy95Zc/4S2LXguvlpOa/GhsZOUYkjP59N0akA3Np9DOIH
JWQSOpYzdotb96ENt4egUJvaA64lDbzM/u1ITBbYCKtBBpAVXFL9vbQ0TA/xFT8l
dNwsjtudS8BRmJRFs0oFYl0S3AIXpR/iWjrPMqtfZVaZteWp7jkYaXxLTIPWQ+TX
NlgcrtLRAt9VjXVA2+zxu7EP9Hdvk3kwQ3nrTJAMNBR7PMsw3oTzG44/dSm3M2Qu
676zxpRuOvVOZOq7/n8q7SLMj80gAyEHWrBZe0MMTGpczVvttXwPiQxcYJQ62H16
mlUB98GdukTAb67X3q9GZHzC2QwchMl8owcIum4P05UdrM70xyGqDSny8Rlx/G63
R/hNJQjcy3Sb+3AfOh1WGLrseWlaomHBnEpL93ABFqwEbsC+WshX2/HAVVA3UG/9
mwLqaIzIZydyBrT7SHJGKE5bF34yQ1ZzBodC+b2J1d42PmhAbdSzq8RxxFNtS6TK
lCouVlijN8jmj7MKD6k5Pu9WnEQ74kq87OuQF0vAjCSASNoBkm71/JKarsgnyqky
SV9gp85RoGT5qI1lBTFy/moszXriVKOYs29ah3cQWzKqKXrPpBeG2ggxQdfZhRux
0O2J7Qv1L68A9oHBa2GW8b90yjxPcWyS9MKeCbnFnSxLuHnDQ33M0ahfx43JJ4/o
uQNGOobZdzQR3UxxpYAXd7AIUpgBdMs03FciauNpIcThwM9LjkT8xsaKfpnreo/5
7mNw1d10t8kEcYF1B0lAdnYfHQ2+egnKDDEQtcNxALfOgR4ThSBIx1W8bDhCoLRE
mkaC4laHLeskO1VdfihsyIIFpE6XIk9EPdE5v2xpGQP1uL3OKkmUd3lJpSSFRjHf
U95w838JWlskrVkuWt5MzQlwQ9wMY1xTtWk/kq9H3F3YB+9G8iocvKHyaMQwJ9Yv
OYIOpu3RwfQ+UEnBeubrqDcA/Be8PE4Niuh4NaRGrApdd7KVk4ogvyAukx6eQakE
PlT8K6aw+aHVfnwg1EvH5PsKw7u6M7m1Pem3txOSkEkqtAkBoarsw+Z23cQsUXwF
hdldydZMOkJtUzPJmntiFOWf0iLEa4INeK8xf5HnwycEG2aflKgqD279mhHjLce8
8urW7bcbHg0pTI/nBRK9+yWx5FX3anqkUf4qfhw7BgWn2tB7HioFo25+mBrxV/+2
/G3+22M6SXAbDteNKUbuAry6SiW53AGGh135yHl7UohB48nZxv1UC1QyD0BnbA8h
P3PS0RqRWZCtER8L87zpakxvEazlF72leI0mDWLUqm66qjQ5OlJVPV7hQhGmqPiT
+YKqUR/VXVI123wKNHpcx6+DOW9RUAX2j4s5qJbMBzRAlGkegr9eyq5DtmaYh6xb
FxhrZpkKftZxGTwu+7ySRSfw3XY4019xdjSb8uD8ChViW1lYwGkuHmC3BXj4cHNv
5D8TkltZAdVaoJMNdJlTCFamMYOhb559Qu27B9ijjREMlpm8VexhmNwu5j3Ztq6D
bYbOOmdw8ARGDJ1M6Mw2Ruwco/8ERdUOe3sk0/yx0uV01TIf5JuBp7Qex6/3PrEH
H7fSD/dxYWSw1By1fN8qV6CV774S773xyTc5YYfseg/VsErgX3XXEbHUDjy84ksw
fLgM5DCx1vvsaqzkIWW4AyDh2fgcLZjqoTic2LbPE/LTc6ytbPwm9WsyWs+2IwbJ
0OtjYFLG4PtS1YnINWguJs2301wjHX9X2NTMK6kgc7lhW/pBG+XhOuZR+nukWvEp
7/WLdDtLFRK4XwEL1VJrTtAVlqUuF7GJ8O+JwC8w6vsZnoVc86mHCAY6VZacAZe4
vF5d3uzwTVY3evsSV6Y87+1L4n/Nd778YUvMXO/uhhSzVHS5OtzgPPA13254Wsm8
+w9xL/GqZuX5aEHDrcPQcxBiwrAjX+NoOa0djTgze5evD5BIoLuVbUyZ+1l9IP3X
myRb3NZzKKbj8DnfvDicQSWISE0XeWIJaLEPx2KKS8K2MLWi1GQE3GRz2BDW21DH
o+qsKHBvRdirm09S0rJxCL3dKv2rW3GLVEnbuD9+fTZUxL+gQjStzlndFUy7j5jh
ZQK3qaJoaKkYVA2r8WQRhGq06HD2AVQUox9BSf6hMiBgagitOo0DD8b2EetLHFcv
j1yDNs0eW9Lcl7ztJdy5yUCcPV6/F3Jhj+gUOuHz0TZkptNd3mIpNp49ZH2kRwEZ
tX1yojqXHep7LWGrngQyZ+qUCB1tpYSA72bFOtXbGECVnr7eqemTu7A7PVWFSctN
uEz/dB+uXIxucIYk1WZrD3jLf2ZGKmAqsK2v1RYhkh4Ch1ABx9ZzNapdW05SP046
aBknD3GsuPwnHyEn8CYvCXtO7nex8lPpfwhmNEsFNqg7GPL8x4ZcKs34M7TdB+Y4
TVd83ljHAurTGZs48I91ZEeWercpXZ6lNKmKUUJ586GL6BMum3PThqFB4t9HRHZs
my2CBezrWBOrC5ZfcOhWJVlsMPfeIyjhRCyQhgk+1y28QDeDGp6gmuZTMOWDhfWY
HqYYktBqVxNvLJzjAqfZYXocigJIqUlooEpqkmT6qhKbFtMsEct1qNjzoJJG7qx9
a05OXD4oVCHDEnTVobNU/FiaAPiCQjsW3c77f3tz4TuUAFyY+SEeKRlO/GKvMhPk
vbDrDpz6SdCx6rL5IH18JrEZ3cVatAauPAudf/oTj6Zh0zwRgVB3eJZKDRtewncV
276bTJ0QXtYWCrErYFNz1uJq/dWKGSDTHjVqkQdKyhQ6Y2xqkJhhv00s4rUMDPDX
y44wTiXFKDIxRIzDBxt3RcCqxFV2LerrBqTugZtcTnmplNXBgF+pPyuoP35yYvGs
zMFZwF4y4ZT40Nu24DHHxOV1YHA/uB/h3IWkUeNwnrP0TeMfUHrao60xGmVL0qGU
rmNaUKHe9/887Xp3VWaXCG6gMyd0gO36gyAUSqri+CHDGnykQ9OSaZMNSxAmHXdp
/yMetK6n2D7OVHSsZFTCMuLWeWzloxz2or0TkGBcF4vbg/N2hD3ef4ewu0Z1lLUM
EDJqWA2HSKHqBBKyVXHuNIi5WAVnarG2/6zxLt67PKIqbtn/H756NgSBkMIYEAjH
iHkT21qxcN/WVX/ILGko6/Jez5MVc4sMjxFLOfNr5psxwTzCWZFySz8AOlztXSIZ
UISrJfX4N3BIln1D2Qod6eaTvACV954soHmjesF9F+p998j1HEaByElvydGrhTpC
VBIGj9M706Iaj6Xw03Li/PbWKSqIicogI14JVYDhLyMdXs9+hl9TA3ylKpvX8U0X
dYPjUfhDKTdxcp7q7f03c0W1OkjRiLoaiiBBfvMBSS63sFR3RFTF6s+XDV0sXnzA
hGBLC9uRqRNKy4nSzZeQPepRTfK2vU9M15iFcmTfBgWx241fXaaj/2uBLmPxkel7
ahkdWb3cwegPEabFq7y9ds0j3hm9sN2Kz0nad89Of55oagNyhb7DaNIHRzhH/nDC
KpYcONC0zx22tHBxg5OfSndDOV/kYaLVLCRbDmw7YkLUfKh5rSk/1OzxrHKurW3I
/AYrffNJit6OYq77YWNPOWGKtOm+Y5dSkjnuMqx2Fg/0kjtwJkH0QOqlbEUHBc0X
UtPxm9DDiS67YzxUepDXjE4YyBeTkSzekRA1piQ7iwb0lf8+iiyljxbm00jfpZcJ
/aDkeYIhKsvTZXBAVT+JuLO+zI+z1uIlPuxrn2YM4ANr0utuDtNBQEuh5mduizlE
Vw1LAxstWA0UAOmm86GAAUT5UIF9CshWuxDvN0vuezDMJgYdiPRyHf5fGH/jAzKP
byaHpGy1Tv6UUOudRb33Da2RhDztZAbPb8PaHlLOcHo4Bcs0BqAAbDg6bP/rGK4K
EPat1yTvw2mRbKCg8Eu70MmarN348Tsbs4Iw6QSOPcYgQSpoQ7BRlz1cT3JVqz9V
L630xA081/wzwW2GILMmJg358g8MdsNtSgJVvm/9OcSmED91R+chiLyzt0IrkKOF
0aRwVRmTshehWvZ1L3143b3pbXiYP+N4Vs14GDgxAl6yIIXeqVCZXv84eYgfR9DH
G2utK7we9qGlywVNuRTVzxYlO3niIspGHGju38+Hxoustkgrs4oodx+toeD7E2UV
yLNpC6VN3TkEgLA4+N33FPWb/+3oKDAr8/O1ETaz1UBs2JNznMNpVv7CaUxYf59k
WPCiSfUxPCwk3vDVo8iAoM5Gz5OCwisjiLUbiYF6cSqLoMkFZvXTt/w6sbQe70UA
wVfP7rYDKZ5oSBx5d0I56Xz2d3Wl7s/IRGD9o5aJkpEEFXPRRQ+jUl1k1aNqHZDT
k0yPe0FRbygRDnLQOdVI6NMD6aVuhrSc5sWFem1LTkc9nL8kjw0p/UwroHTgDI7q
G/8c7JvdFVuvqlrZ8KAD/YUox4NP1z8gQYNXSB38VM5ovURhzYB/S8JygF25o0Nn
WHDhXl7b6Xm2xPHSQCEAJ7DKtEDPVGD7tg2S9CJcy9u0HjkoUHn5gttfqwPbgQx8
M4hpLNpe2LOL3SRQxTAai9WhtPzog3MpgeYyZT7DpKBy5sgF7Kdlxh91aGHnWlnd
JbTEikEvH3veWW+XeZI0BDBnCI6zvUP7RjDbj0wz9oD5xWV5KpmfmeRxLEumQluY
qNYwS0EScEcnx1+uBSQ7b2ucz1g4epi2heowM5Oe6d18Hblxpi+IoS+qfCFqsxgw
1b8DlXqj0IbBQq7oC3U3cm4+DZmuo8XfJvhqDc4n0rGCs06H24/dpNPYs2fh52nY
NTD1sry4IpJI9MTaIGfkaIQtXnz17LXwgPairxlORUWmoUu5OWZNY7Fim1sWM302
xYH7cd5DtGX7qHxBid5yDuYam8lSqEDym7Pcrt8OuOztRrsU82iYs1FDgs5DDQoq
4DofmSH794KGqIOiVipR0dIpSteGuFg2Rr32+p7p7Pvl3/7Ts51xCZo/Ow0lYr3t
ACm/+BnUeYNP30VSQk/E4bQU8s7eCUhdxwDqcPTUCMNPJSevsjfqJ87Zj3mdZUZS
CcsrjD7nNR6h4pqQDmARSY1632RwvVxX7V++Dl12cdCL4ACPWkdqVmH9Q3AWgDe2
gALvzth27IdyW86t/Rvzpy8aJvPyqPERPBj9Jn44rYZ7b9xGmbAJnOoJ1V2OeOAg
94yUfC3rK+tXq7BYmhjXYMMA2FTjJiEFL5MKEzMWL2IWw0qECoCe2Mx9fS5xj0K9
8WZ2iiNiqmiWDzrXm1Xx0dqReIrRxMuUbZGHYLpJVzNRqO/49QL8OsEvXUqs/taY
U44W8I5mpKuiVCCmUfX1Mat105UytuikqjaM4X+UR3CCA08nTvBjYgPGxNrecJKZ
+OlJJztyoX5DBGYaYSJGSSULlr6xnixSVOY/VkXmVjEddKoEFCaKVRTGTYx453e3
44kfbbsln0ansbuxyLMowD6Y0A+198/vuUpSP9qts/9gobR+W5dUMQvp3jRTN6Y1
ItfJqhAvC53BGSJ8EBp6tdHlP1Lq7Dc3SXtFoORDMu8eYL6Rl1yN2Lf/z70MRUgl
6/tcWaMcPfRyxDcJAmZhKWfc7pq8gAi61K7oa22Wcup1NgPrq3sFyOZB05ce2tDn
tpTMT/ohC1J1DisSNNytfv5IgAj5yiwc0AMCqu5eKplLFH4EI9gSt3d9C0vEXyQo
jy0Kh8giHW5I07yXMmhO46kegayLYk0fMynUBUwJXESeDD4wD+IuZGXwKCsE49Z6
hiw3ILlzSXhmUu1gnrGf573qSnp0XwnmVWjQn7X77gSUXO+o6hNjndJMOLtDW8lZ
VJhHdeRXb5cSwXIGiZbT/9tVKPJqzHD82N4tKSLWY/zPfIwDunT+U2u9DXBqCZtM
99GMo5d0K1UljYiTNoPCQwwuH1Isv2o9oXbcsGQn3cdhETb6JPwvEW55rqMteQ7D
lSHpcUjgdIn/Mk6DzundIloFtxkg8KTcelIQHyJbJ5d6q8JU+3iya1FB/uGRi8NV
kQ33hoa+86sIIYrcOiTPBT6n98KHnba5jsK3+eIsvcWS8GTpqmk1FRWtyOF3xcdO
O/iQzlbmhzZiDHaexLIpfA+hlhLa8eyJv9fYD7uCP6Yz6e+UHMTDZr0TOa4vGyDg
3VoB71/CSgqGV7hW0/RT1FJbWPalIBH5i3E3YMFRFMRb32R45u7/l9KOediUqvom
wgfSuAuyQ+CsYWfigOyPBhKdGUmBYnUVtUqsGrHYhvHdzwuTm7kDhEkBYvSUgGaq
Nl1FaYpDgD4TPXG1v7HPcmK4JvLLklfCHKTp5sNOst6ZLirpbAgZ8cMfcCi+TpMz
7zs+uh6zLfVywcNTZiiHPitrRsiYYN8uqNzBljNKnzyF40plE0Pjx+aEs1hVpp2F
fzFM1bDaZS5O3aQ4cM84qG8ssUWbWlfWnFRc8qEb8k34lF9UaEmKGaUSEnBQNZiy
RK9tSBN5SSDht1mrLQUOZ8Bp63O3kXe7v8nQ6AsGEeVZj2UhLQx3sZMwD2ooWVUf
73saTpgKXLg88+2yC4Z8Dw+GnoLPkl6vdYQnUOGIg6JQz963mx3+bvguLoSCFCXc
USSJzexDUnT4DQcq0IoTd9JTzTggmF6lIG0kGNmxzsKxZENnkM1z+HVFGqU6tzCe
n1Yvo8cXPBVD/1Et1tTS+ZVXFjUpPOMbzZD8KCN5eH9evJEmV5MYljkqECJ/wweI
TFHuuLRzodmRTJu3AkGZmbAn5JrCMErwH5tddKChmVYibMqLa5cs8+Ds+ChyoGvg
CYLeo19oX7RjVEkHIc3/3csIS9xWLY5NxKMrcA9HJb9rQMu4rHH1v49ktB/PteHE
O43QeSlbNGSGSlEgJelwf5WE8ySvVv14fE/DMWdO/Q0wq8WzUuE/xWZfnolCObeR
rJPxkTPkUE1prUuVSZsJuKETDqivJCrRIQJpaa7Q3xLA6cAejDCsuluSJsOD3EXU
MX5JzG+fikKFPg6YQhBqonhPVNolCjMzA/w0lq49trRJ6l6eFxXHhimME5ie4BpR
J0FzKjKhiWwEcBJ6Rg9D62k+dJnimXviK7eElqJ3zglwgmt+kjS4zpmeo4l7Wnop
wgKnqQUNY48PknS08ynWyJBSVdWhlGmwTVEkW9HsCDMASpxCGLATKtEIS1CgfLPN
DnohfY/2bZgAkWDcyhhAoqFC/eVVdQ+yk4di0P+JeowGa0Pm1+1w4k7JumSPJc4m
IRP+z2iPA/L34g2FRXz82jrAEJG7AXSJYGOomxOsZ+/Jv8mQyFG2ot11B2u+ZNNP
ayDUVmgmI3Rg1foYX9hdDct2YcEDzjt9hNWUO6txNOiA/kWO0r5xzoVwZubM8aXR
Lsl4KnaP65QcnT5bFgCUp8FfCMK5isKYn47O5phlKHM8aADAWWjJdSxwzEReJkk8
uHWRGw06HoHv7QVuq82/NUZ7kyxzD2mmrWkP5NNNFqJ/DkRPx8LDq8iZoVZY3CiF
UfTl6RFktYXb9gfBlJ1mMvUHeExNzo2g4qP1l9Eu89QFh6vSI87t1Udj7on23rRp
vUiDKXenBNBvGrUshlZBucR0vkm5L7+zS6EI7GTFrZfaBZDk+1tNkkCySoSQlj7D
op3zpB5h0LYFRrgFTtHUhGc8FNk6o3lqdZR6c6hZVyaz2pXTCcvIzhvA6DWS2i5A
jLDCQD3qgY35bXlg0Jha9zS3/+802xRd6p/rmuGMw+NB35lznFX+T3x/UOmgOKYk
xguBzgSRLofn33JAkr6L1wWOg7W6hpmJbj8VIZoAhadPUQEU+BvEkUe/HAxyVmK9
67lbiSloY7foaVA5oy/8cDdY0NoB8kF1ddRf++l6vuQ18HiipAn9YN7qarJiiCpJ
Y+k3BXv+HpjRV2K4focLH9csNOIfg/l+wpo6l8NK3KaRc+wlqMvd9DC6icWALGqa
6EjlD8fhsgAOduaH48cs7du4UbQSJygTMnzaW1cegTLkpNqqtqnCXiJK7BtdF0iZ
iWvkjp18IFJ6MsjON6p0hP8wawus81UMnmzsYxBNE3WTUYcrWeNDo4eYk6np/vfW
MlmV86WLRcG8YxDKVZWHybPpCGjoxPzk/F7mMEWB2Difkcs3/Qru6V/QdX5/SoH6
DERUuIrxQrKlxDG1b8Z8AyoJwgJZyZ86m3xUOIgZbd6ob7UfDXoTzE4M+sMkGzDz
KkWZ6cr3qCnMzJJpg5AsiN95mH7m6eSAI+J/xPI4h2CF6iwYv3CwwUcj2M/TUNAs
mDVOtX1DGSGA1mrU3w7wbDeqUhcjasFG4nKA4jiOssHlTbwhbrXP1JM2i2iEO9Ce
nIPSPOMUI1VqjnRpREblaiKEDrWbgLOFpNwwpqWHXh/vzh1DiWRvOZcSeLVLcxFw
oneg/PhMCQSq/RI8XFzwtW+xxbsvL0Evxlzv3vvI5w29CvkrbiMn6cty/l6E7IWo
VbI4xk2dhQj4vC2noI8cgM0XNOWb4JKkIR4MuCCzP00D4XtlVdfw4EMJIpy5s03/
U0b4Fa4rmQ8ND1NPZDQYbJpPycCA/LUJX6BlUwMazQ8TJ1Jy2lJtIEFoHzzLC9SI
N6FPycH2xMszn97e4UVZ6Anruys+K30UuNURkybpNC5UUUjNfOgfyRwHk38yfEkK
WG9MXxjAhEKj/A0MgliiT7JBIsghmnQAbrtFwEIEfl+iZ/EHFYELLPKaa5yqFOZh
g2qIuipjrI9b36U0Y8sdhT2JdkYEp2p6Zlv3N2oW8+77zWLpARDSaMcx69L0z0h2
cDI5mhQCzCSclKH2po0KL90W3ThZEWgfA++XowzXsD+IKG29pBZRR/n7GPJc+vkk
l3KT5i53agRxB3JK062Ay0uEMymdg7Ru51/lFfvFiswRmgCS9/7qzs3preG3M8ff
gFo2OnV8Gakqo2M0zj++gvpeji/cL2gbsbwblXVpCbAxECOXHZ6O7ukzoiHc3a4N
fyD2ogDi62Tg7/IYRquIScYLwfpCtwHHVPRwXrvb8UZqzJkBm6vuAlteVlt4ctcn
tdRlMHoHTU/DnXRr9gNqKXHVKLzhTLCjQs+53mlamxdJKDBfGe9jxF1aLRMJ2tJc
fjoMy29XV0Ontr02S+UjOc7znRv6neVBEqXsvObwOFLRCv2+zVlpGg5H12fVy33f
3w/td8H3OIZ0J3dLhm73B+Ao5XGZmJccVqTjgdoW2fiR7dopybTkSUSEgPmPrx3D
PriZalbkvhc1777SUSfQ1PuyJiU+6jmVhcQJ3WmCAuNbAPVBh/NQI2ymfgpp1ixY
MQf3vlx4rcaH8+Um22cPAGfBASw31j3ec3ec3u0QfWs0LBpVmsg0D3ge4e7oad1W
+D3e/GRQVZs7RpW96J3SESbDDamHdNcl+3Kp6UBtUlFt9F6aPHhrgji1JiNlQO4w
aiCe0G3hvYf2NRl/pL8gZ2KjNbTwtIbGX1BLrIjmkLlRkZMeiWQezgTGOAbUEcnn
GKC3mkWJesuCFZXzVbmwiAaqgtxOu+OFTD6McKzgFDQbZGLJu9qOHcVOIJdVUqVg
IYN6E4/MglgMvs+lNEF1EbdVIGYeoVvs1AN/i77Fu7jz2DFZpekpry7YCbmHNjYe
GNbzN8TjT6RE2wtpCQPgZ7k/SG0vOZtclv322Xa5tqKOXIOHgL1He0DyOVKHv5FA
NOJuuvE/t9C2cdIbw9PKKXsmTTmKveCM0T0+PbwBQJaX7KM3nF6cKLoC6JbzKtqT
MsrKBtn6vY75t//NHvQ1YWOgqRubquryC7U3i9pHjCNbM5tUCXIOwYqrBAfcAEZt
bRNz2RLP5K3Et2uS6dvWFW8AIY7APkkCTb1h9YFXPz8AVMiMQLkkqxOg3Uu69kpK
MC674oKs71i3WAgHUcJr3H6pVIMrKdGVjjZEw2I3KTsPkJskAnjFL63IZYIFkICy
+UMz7LXQZ1g6Dux/ixvwz4sJRVxJPCz4BGv5SpACIapiacwOKjBzdDWyUWqAOUhe
h712w+FN7M8mb4fjniESgSLHZ9BOIX1bXP2A+St7xloHR3+XivmOv+r+V05cUSYb
EwLyMywNZbEIw0DNwUnrWyHi1dDOvHniJYfkotHbGbNCGq8dgPmNpDuZrx89cpCt
K/cE4rpPxRxetVbROLpQeG4ghwq4WjWPWaPRVRnbRFOftzhKFe+aTsrHG5yVFip+
wZDFeulsNgXDtq69NeY5rz4ILHjLnqmS1AAnYtZQ2idVc4kkRAgcEKYYjIYX+0qE
vZroEJgtfNEbR0n4cnsojb8xMobZxpchSARCrM3AWVd8zqHKg9vzawDPasvpl4XI
J8azcGrQ+kpOa+60F/aD9R3c5eUvVzfwdW+AMUT10kqQ/ZkJqd284HrP9fgAJ1fa
QAcFpeIZwSzNm7ZAmmy3xRsR5BxUNHSVCmGTtCKj0mT79Fw6TyUCwySeQ7xw1bL5
koyQRQ4B6pBj8n5w3CSw53LD3Swl4KGhvC97a5xadqFDehdwns+NzsmdqY6zKUYb
bnwo2eECbIVc5rACZ1bTO7x8VNZkVKv5RBPDr40LDuLGo4yj6Va2QJVptqSW+H+n
qIci0azSFc/ToHqm9Gki0p6uVHebYlN006Py0mmKU71HdjRdPlCV3cJ1/JOyBw+J
yhdrbbacH/w30StQ3YNY5pwaukXceMIuFaQYRwH5ICmb82pgaDS8XBPof/mml/Go
8Z70aVB8c8ehEyoO9fTq8k0AQNx9Kl4Q4Mv/6m9HOF/ucyU1vFATNSfcSxyr4OkM
rnwneHYVGfX1pAzIfUZzmz2Pb1ClGZURwDmyadzb07DXsccJqFxNtWcKeSpbxjSj
bwfxNEEEzCn+yHg5EzTFdf2XwZ4DiMKb/mxrvV53rwPQVV/OZk8FRu96jX0UH2HG
JpMVzvZkCc5nX3DEiZ98OJkD+Z6uw6AZgy+126cNAVhAsyk2lWgakXpU3muZO9qf
dJqDoz4eiH50ZbLq6Bcq9SKoUcexb99eUqpFwiHYdUvqAeB37vbHPVfR11rehLLe
RECBJd+6pG7XX84AGDsfonBxqjHegzAZRWC9Br5K10CGwXTwpRV8ZnS3FuXoT44S
CbrAs+rGcnS+xyP7lf+YjvVX66HGlKPZK62VTSnwDHvELAa87K4v9af7111ZuA0Y
gPgYECbkfnKsXB5o0DfK4eC4s+XglJDML7BL8jhrKOhjgS8UWUf5Ls0sKU73uDWX
T/jDV0c169KKMIFPnI/GdPqzZcmoqsTnxUYHmGYK00PWFr/O1VFJ1SIclM76XEm1
JCYUOXuQB+2VQ/PF1mJ1j3DIBu5v0U39NclJ27QhV7P8d9MMtAWR2J1ZljRMpHAy
rb4owS7RgefoDdlOwWRXqoyxwnTyhfySd9zbRXuvMs5FcLD3Fzkh0MaBspxdIInk
rGfbU3lu0nFbKzgX2PPHjLIWRCNrvwemcnFGv7JkObEyTZA43uH+bxnCnq2zchVd
JvDrBkXGzjsP2JP+ISxI9OEiXp85ksfU3oCYZpjVtU41APOeKM1lrgdD6rRaOw/C
fR25EpiEHeVDo5eNSNu7p2szrFDaBOz5UKp3UkZQqlstmrpiAUm4XH+E0Z8O0NhM
vyr/tkhqh7NePhcIiWqDtawkzB6XslGaznLSKkQTfA8wZPJAf0fVUc3qTi9CISxi
lL7TdlWjUU3vzNXc4paEHLL8semZp8GLuz4wQXvKc8mXUYzgEWxYuR3yL1Dbbpb7
FQ9mUcAdB908ZQI6ghUngU5c+U1nZ1U4GdySFpvRaFMfQCW8v5vy5N47fPxPnPqe
0+NQ9Kf9ORUmowMccCXaS5Ic9vgdUdSg2xkB+o+nXap593otKVp1MZmAXGac+4wo
NfcUWpdZEk8Wj1TceseU+lR+swZrE4MufkhhgMyx1hrVPtDKo34NMwA///NUNgWz
kZxZadB8KClv7ofCXrhzEinJruYNdBEafa1RyWDV7e7j6CeXtET1hLPJF2plJwPo
mA3vP15sSJGfdTHwfd42qmH75oQJNysfvPaC/CO0Pxcm583s6nt8ZUEBS4V+NQ51
h3IsPeDnVh9RYxTmqtPxTS2DPvA8mwCzXGm4WTdPxC+2ypumuucXkusctWwDoaKI
XgTIz4Ij4p8s9xJs3G0VujjHfvW7veZWq/Aix+mbhU4fEYsXO15fieabEfROnHEd
DBqAEDtQILWikjmTy68584VUCwsGOHVpa1NFrXONvt6+8pyaJ6+jxgMytP3SfHcd
29ACQ7uh/nBSM5lfvMImWddVhHVS575zhkm6/mOjjJU4ZfTcLUtBoIPxob7Zdd45
9nmoyNYr28ZUUknPnU1rdEZKKQ4IDCScvox6lZUkOp2qweZCfKg1J98IJtxG6jPT
AlsuoTQc611JCrmYf19/cYP035TBRj2D5axWF+thOHVdlV7+KlZLFdNnrpCFmwrN
i/DnO+FxfmOOChWSZhO2yqiVovHckf59LL1tjysLZWp/6rTqwETxA/F+2JqQ9rQ0
JQP7CUbNVzawO4n52sEUyATBxdUbgfdJkWFK1jhVKKw7hwkmBzpao141bm987QzO
GQHC2FOOf6PKyaYRMbFXryZgR1D8cd9hvvYH6PHRq+DVTsQkKT0797r3uUMzl/h/
kg5PKTwhnGrznQIVdW4nJMM8mWp3v9JcwEKsg2zG3KaIRBS8JyaY+jkQFbwBA+JW
3ccal/6MppobBW3LiCOhB8g30/0b8vI1ZZVfgGOJbHZ7s9Bu8q2UfVxAl+rhFUbi
FVrrZsoGdoiadepXOMvES2dzoAkXG7UlzXeLUOIUtR3kPbrxBI/gj5FV9Zmjp62P
l7J42UGravqbcfA70cPBsk9PrHVNjMXXtWCowNuC++EQ1GIoKpDvWVlqudR5zQCZ
muJ27NEtFyLoUbP30O0LhqUJSgLriMLqeTNKJrUSaU1is6ii5+T5GwY5QC7V/QQi
0cuSGi0uXwoGtLS7kcu3ABSXDFzKTmFzdGoqKYQ85Tl9455BwFD9KSs10vw2FgyB
p6RVM4IiL+GZtkz9ptDAlq17/UkeKz5Np8F7DfIfc4UeV0efNED78Uto+2qQiXmC
i1KqsExVu+yV5uQYOTKYOH/SKr7oU21ovsOgR908xFU28Bqw3OUY0WTeRhQ8neqk
q8GbhAutLxaaav39Vpw8JwklndCQ4Cd3Y5zocA41T0aMqwNXk34aj9r6KmoT8Zqc
4L3vOhVp6dd3kzXXltAo9U9GajwXGoD9XIKFTSmp3go3ITLCkI42mN4CnJ/XrDxv
k+Awn5s6XfCUf3wnWzS6yIqB9RSg90KH2e0liMbgrlY4siu/oOLiPgwxirVXAL3K
p3ZFOOFdvsyyhupEwO1Y08bTERGxgFuSfEUoYaJ5+BuozJZHqPmcUSu3XHtVBLMW
HY15hW/aaYBSCGeBedZEzuXmgW+IpiUC7jLoEPi6Q1GcT2sE1Klacb2FQsjtwWDt
5aGfy1rNskf7/DIr1boDGMfvBiYOYcB5YkOHyoFFKfKx8d9ddvKjVS6aE1Bma1IE
PJxx4FakKIbqpO30coU2DLaXBTmFal7MWxi+Rm1RONdgmK3qU6rR9RSzecu8GMxF
M3iQKgSJ6Nhfkt03FjmnQGDhech19ZwK9DWEuZbzV1AwvLxCvTmNhsdXVyq6KkNZ
bThsKsPY6Ky/x99i+hYIHihOmU2j92nTq9m+dZ9Kt1XArlPNHCD3zLdiXkV2B6d4
rvEO8S5bvk5ALJqDERPlnthPDTspZTNnls+DwbcCE6BkRrg4mUXuUExwpB50iV/V
L7xYtAMBWFKROtGGfBxuF82EZSVS6jUap5dZYm4gWLQHWKVnosYfkJifUHdmDqq0
c35ZXuTKqaU/nR2gBadRzYn5yIR84/UmQSNYU6INxzb/AweiExNc9o/WryDc4yM5
SVOwlTEZK+tZcc3I9WfMaMoG5EaNnQznD8VGohjicZSKU9NIiECclv3fDSOTE99X
MnVtw8V6I/m1XICWyquApoeUH74Nqs1/eIe1Mk4cNFc4h258gtuhFGBf7zISMgp0
s2hEH9HAT6EzGmsT/iUY/Z8hfoKF541bdK/Xjo/8Bdszgp9qSQJRfYW4Rt8DQVX8
At52YzZ83ni92ROzSJEBry1BA8nmNMS3CWuq0N5mqrXnHGeRONtguZiXXeNgb8U4
zOlAkDGizUfQc44YHbd7rGaQar8rP1nDgVk562Cn/d5LX4x7LKXDNLWuWUc2sJdh
jkzuEOPfep+DR+qMvJPaaoGDPGzardxCgYAGhYdi1DkmJh431ll2zm80XlEPR3PO
4fQWUP/84QwmyOeLwfmAl8Weaa8Vgv4XiNb3nATzS1w+04jr7Kr9loJN/oCyfiRJ
FtdY5aiVjVl2QOrwcr0cz6kLzcE+nAdd6tMcpXxhNtS3CUkzCf9hsFXiUoPy1l2w
CqRYpPeGlPQ2+Al/1o3PGcMLJla+/2TsGdn5QDVcYDh8TGMICdt6wEdtZcflwRQT
pczATJ9Nk7HY0lCmjJOkXZCPTtIs1/ijLFlmCdS+1WoiHYXcDHIcWGwE4fawP+8w
I8E6k1V86U9+1getXoQeY+LlnWq8oIFaRPT24zP1KKh10/kFwWcddmPvajvfkqIZ
HliA1+ZdmIlC2ueIpe+rhgivflrnEI3QiQcRmCzBSGsuU7xwD9XORqA+tVowD1Dd
XzjjGsKk7uzkAuzigvdHcbamdTKYjweUX/nwZWZaH0Ltfx8jFFq7Fk2XzUnVoAvH
mHJMnjT/4lnFzPIo1xiFF4s75q1ZUl5ZGNlLIYHqO9+7gdgWuH7z8UOWf98EKAyV
RTNb7FQ/S632Ji/U3tPtTi7isl4iXRSW3+2brXqF1MZBeBJhvp0I8kJpsYUWktyW
nvFq+iq26nXsmiUdbaaZaBzypxjY2WlUEcwLJVzqwy/2TuI/Y2ovjQ+UHsRxskEm
JF8TaRN6/A+TgA/S0U/8WdvjS3bwA8A7QYXQ8RNF6kynLCqq/6+fTU9LdVHI/kS8
22WVgbcZOaxLrPqJbQ/wmM5KMGopjLqajWwsWfSNOJ1NRyWA+ytRux6RGSfgwXLT
QdquwDJ/za1U3PKeLDrV26/fq5OxB5q+VtkX4ysRFgyjGZ4xWjApul2+95pCBnZZ
u/xBTy0qopVAvWJ+mhXZgW/jxwWINUARNsFwAwrPr8o3K6CJU6niCg72ks3KvwJ3
6P8qqvsMD1uDpG9nIn2gGYOuCZP71pp2wXx6UlKJmWFoOhSqyRWaPq7J5op8tNI2
7V0wrstfDUakDgwErzIVILTNd9S5YAD8qRAHFbijRl8LIR8I2d9Za/reG2WGLnS9
969KciYDUlXLbVOpwlPMY2sRGREcsUuUTeY9/gFdN0ckBdoLVDcOz3CQNYFF1PIV
Nfx2anqpokZ+hvXuqkrXzPW79VJ/CMoS0KbXaCHdY3vyKKdzdc55xXs0j1zCyydo
oh1VuCZr4OyVOCZeJZ/P5oU205Mu8Tt51CVVu8XoYt8Yg3X3Zi8dWutwu3KWSm27
IBdSuPuwWQJcPzFNv/H9lWV1PWM/8IQRrjsJ12XZz79nUFh6K97QWDPh7RfhqMGo
YpuK+ulQV+jkRDZjmiEi5rkKtrCkRwOjsjHhTulvhdqTID50tNPrcA1KE6t9z4bK
i7CPG2/0dRakyF1QED2Hi+CLSxT35yE9Ej9rwxF/nk+AYGm/AX4lAQJ6MSuXwML8
MatgHd6XHXmjQjkyvhgCRetiaT21QtwUPaQQ/9TvT1JUeik4Z4pPuoCdLDYnkkQW
y1UTdqch9fx6i72hkTs1Uq22JkGOyhEEPjBXBWlOo6ebYfiBNCGAvUpkXKD0YtnN
1dU0Oja6dwFmrIMrhnOpAYs9ypKkaGHnrWMHZ6iB+d2WfncER4QeufPIaDwel+Vg
0lMBQzC7NftyDcJcBe/9DF412b/Rji0HUxIMZAen/KQr1dFKHTCppZJ/ERzmv3aI
32x77GUT9Ss/AA+mx+y9pQzaetWOkVWSmpoGaSSPTeyMpX56ig9KvMSxThb+zHTU
l2ewkzEnTGTKBuh0ByGjs94NrzyH6wsI1LaXmmvqy6Jmxl00R58zZpUmJ6zEja9Q
phbadgggup8DdlEdJdZ8isL6sj6RVB9+x9hlvsv8e8NhOi0gsmOZOyWNSbzVwPsR
G6RkAvOkByV2cZcSs5j/ViVDTj8+dNL7xpRQgJy0L7HQxQA6uAUyLif/js9T+X6k
Gihp0Ue2QDaW/SJE/OmxoQAUXdVDBE3Q5IEff45W1bFGkH8uOwswkUfnR4TqK4in
0Y7etU+u3bi3XbH0ADuRnYbgzpLBWU7858XaXF14+qKTzNpb+cUi1IXCtJL1lpw7
DUKxa0YA7nhh4ZTnuME6qW8S4MfcSlgHamkJo9sQYKdYGqLtBBWeJbGNdVe15YRR
RzMdi0k8OzPLhDGjmH0gEOeWEnTyEFKARpVgL8Hssc6UcJu8ig+epEDCupWS9rKI
7Gjez6jTmM63CAbv6B4c0Y7ypMfujc857OHIb75ixG0VFll7HTKbWCSc1v4qjDHr
/uRESrpjdGuMShkcPaxc4lbKt7BPS3bBd+A6ii1GvWS7eK6+rADz9nLCuME+kn8d
yWZNFwUrcHgmyKfgrTXL2IVLp0vMHkFS8gb4kthXcTTvKA0Ba5IJ6uxQ86HBFxr7
Pu+IfEDZIQAYIHscHb6/Hxf3ZYxDst34SM5QvZbyujCEQ9zIsEidorotwCvglHEm
gkUw77Dq45dHoeI5aXqqLHRgbHSPugFBzSvgYKcbca7tcglXe99DLqqza0v/cynn
rmV+3bbTZmz05h5S3UbLUKznilAgAGkjRSIuLursgmUj2LifjZCOJ2bE3Rnjgpe4
73hIwXd5ooQaD3GjWk7wwhJehL1JAJpNWmqlBHTtmLvZNVoJ8dR09dyV0l68n7a1
Thif7++iGnYtvW2cbk2FyjxseebLX5KhWfagETghO8y1SvMqDfE4EIHc0PAG/Lml
nx6cGOTSOKlNTQDl4TPaRX/10gfLwzkRCsC85csDomf8ZAgHbO8AqFv0jMRRz1HC
2Aok2aoVD1SR5Fg9PmwUXYK9viJj6t2dMtPCeFHPo9s4667BcUjDZCeN9Y2g02TD
FzNw6agPrBXoVSYRtmgAuuzqgHKhj3onfjpEylBXiyeKt6+Elgcl6lxsXUr9fHDm
n/HcjrhIFf0qhSN04mtkg/imh3Y5dwgoUkl51W3Yl760qeMdvDLLnIOnejmIr57y
TD2vF6aw9bJGykomGIrC2WMxRJURZFNeOrFHjAriLLPVX0mlEvoshhPsgTfUZD2h
hZynmtAfVs5m+kURd+G469IqPq7C1JQgkVPwz8fU7bjrfnFLlYSFBQafaj8dC4UY
oGBu+YUX+ZHqDusLkXUAzfZJsVbGw2Yyri1JbyMAHb6KyeBBQLjMx494F9lWwQSG
fto5H7l83+r9JbtUtr+Ls96r4R/2BMBZ38NSlyucFeY223Jq12a7B/d50Cr0Br6x
HkSM60ZMW4zwCyn3ZB9Kb0y30gctF8vSZcfodUMP3MOVWCJbxj9pG3AdY2XECmy3
66pW/2vc8jMoJzfmTBq2TGjLyrNZ48p7cUKcBY89w/p2eCXBUzJfX8a+dI/K35o7
8GWZmUinx6DVpr84HoRq6Xsar8nRwvRohiwTsh20jIC2228MjCm0o05SJFoEmQAV
Y5HpNE1BAomUvN0JVzBBVnOR+aZHP2oP1KWxvAkLq0xGt/1HFpBfLGTk9Nv/o5fN
MJm1iJGfsIq0D/cnX80RdKzjheZ7tCI7MnQ8vdwq1MR11cz5+ezRnickhmfc9PGc
Nc7/iFvJFVQIjnqN4NURybxlWWrj6OrO3gsSCk0BH1WaU5wLlmXF5FFzG7i4G6iX
Ftqc9vO7nGOoAIF2ME1gem6zYuSuBa68v9Ifw++F8Pnb+WwpBB6UOR0ezR9xdBL8
9pQPDp031zFf26IYW+mJ5/sKDdGIB2OGrpkxOATYDG0FaDCKNCYSDZur+M0ezY6c
cu90PZpSsLgK4h9bxHCfzQvC0zBUJu34WGl2cM2rjfL4s0wXI8ESb/MjpBSNWJHx
tWmEesH+b0ORPHrKljkvo4ZTi5h4eUhFNeBKqLkeHDI2iXJgHRMqBsMG7vdF5cQm
nJqzVq4Eox6DjlQf3rzo3rLs/U/3B5mN9zOql1SpbqlH8YZS9pueW5DUFUFbJ7rx
TQSvA+dbxoXVjRmTgaySGTYScrV8+hvmqmepQzoM37hJWlGSnHeUi/CsJ4/KReCS
WojOrRZEPOTubCZbkoCX9O1uoCCdIr1ukmxxxDWjDUcQ8onom2Ve0AuFggLW611e
2dIFlP4angqbPxPHuiZ4jUHGXDQwYiJw7zF9g9NNjLv8eWHV8Z7nt9JL4v/KlvEV
hk0c9uLFXLNKupDtOJ64QqlaTmapTArKWv1GPb+gJ+/Yx5mWoQoMQ29t1S1zWNZ6
Q+bdJZ7ixSos6W4bJ2p2wbM1GYaAhjJzliprqHke7aCbIEirWv7BbDOOSGJq4bjM
tU+VTuB6iTqO6a1hptjuDPD0pLdObA7OtGyvUNBq/Spv45ZoRktEtAgg07KhZ0Mz
MA0x4l2/SlikBh5tPpfW0dFunXW3xXP/w772KkUsj9cm9jkf7pe4EevnbMGJseo6
3L2D8ON2V469BEw5PNYh82J9hBbeTLFFvGigaVkGRdNfFm8WjDA+Eo8Dyx4BXjTq
1P9EwHk68ysK096zf+RZLPxseSAQD+c03B7uTU7JOuqbzFKtVuMo+CkZdYwh0Qtc
/kxougsqIvmX2MHWH98SkZv+gB78OhPCwDCnyDV9Ge49t0r2yEOOTZRTzde49+Qv
PTYvcphDNP20bdf/K3avE9f3Ulg3EnR1h+JIarGh3pppVzrZs9X0P6j+Sny06c2K
ajLTezet372cnPmj90Y30KwyxvzGRfsSl9VZHZ+BAiv1HIyoDTObtF4E8LbXR6j2
lMGA34eVyw6egni/hwhlDhC1qPcG3iemsUpgtXunJa6HDnkBtqhN6aY7i6o0o/Fv
klBltrYyDBtHtRhCuqqD0pbNPWqK5BJH+r8LPrYx0XpPFJkpVAq9fsb8Mr8iaYwI
RpWneyAYRafy9oqbYIwMEbmQwp1n8RIiiAr8yqko23nElcfX071yd5uHB2gZktmT
E0Sw5RVucoZ8RrnzmsbvBWxmDb0SK4jSWMAoelcNU8df2/MwI57gv1tBjrB/ILFT
trGaP0HQKnl/AoE4ojTVZceLOyrrQxqqBHL5x8vJOesbbAfqlSHsEwOeljsedx0B
sTV9mEGsR/fcmdYTc9oc6uA56GfsiXKc9ml3vofES4lWsTZJKJxgQHtBCvWhaz3O
G0he2aTXCusrMQqRmXhbNwMnCQOsV3bT1DtBW0QVo/0qkMVyLJ+OWib9BV0lFA0j
kaOLTnNd58kfKyG0sjlcNRAkWfateTMt3qGczwlpU0dUaN2Jip9pgM5l3ZQx37yA
VIaYPaV8LvWDEzX75YU5nIgZLCc2lzjmImvPYcwrMpvF9rZI0nz7ebUdeCM8lZ+S
5OGF2ukQVpEoBzTt3MLsMF5RndAstt7rzwYRUcTQ8wwXubniRwPuYsgiN+10jyJL
PnbsddDVgkAugDTvsqjVEyrI1zIS0VUuQS+GQJjXp+bhXoSkgbKXDPTiJifwZdZy
pOcrTR0XJzVa51TXpQRRnmO9dFjabV51WeGXAV6t82C744IIwVC6spVebXX9/9CQ
2Wm7ZqfQOjacA5ym6CaDmp0aIM38crjDXl6EFR1TZ90X+Dhv7M/BQhy73ldilHCu
/ahhCVQ9ULJql7zSa9Qj/tMeVTYDlbasLkJOMVKchNpzWKgx3S4qVe+DNvbJT2kl
l/AMsUq9Ep5mwv0PIEA/SZOqYCcFp+z7a378K7wJ06c2p/iS/GMfzBq+IMpkwzrV
l9nYpluucPwshooTM3QFEfw0B/490TMlDMD2qQUbDMNAuOssG0v8oL/1CCIxMFY3
nlqApjlQk3qdti1+9hZkEbBCLgltTYuWzPlrDcgoD8yUdYWAsInGvajAxlSGaG7n
pIag+JAvPOp/mTNirBhN1hj+Q2RkBI0IH/wVODlos5C3NUcV+OpKhRLbNES3DpO/
CQbOOywiezQTAsTKn7WJ6qYM+Bct5V9HZSQico63Jdn5eSt7Q6Nocd3PzEpnflMs
9VXyGNmo21hUjy81OVSOOZBFUxoeNx0jIm4t6J2WY+KVw+Kjmc/MdYiz0ga+2Oo2
lj8OXvbU1W2p/g6w000e6/QiCMWjZwxEtemdjl5Vm1S1ehQVKTky1sRrlHPtmHWo
JO2NSX1Tu2R5Yakg71raS2/ybLRImWQCQ2ap6aVnU6YKPNwTQx/nzFmRRb3o/9g/
IUGaWsgI9plb/6cpkhBr56B/8yztHDvUP/Gt6/MwEp1U3En3ekUr8T6Il7O/jiUA
rjX5qCQ0jSzIg2UlVzddTeIkhRVEcX3XcPtM1IcCS7FbCfaY4cCCXD1/fcMkC869
OIhsRSd6UKZeCn7w7olYBGHIvwIghBBpN8HJFtYV6PTwsaHQGAHqz6joyF5DYLeW
d2Qz4cwgZV1gaRYy37f5T6n3Et/mF8Ue8oG9sv8WKJgDYafzT0tKIClcZkz1sdFD
yqyxMX8QxmQ/o1WgHIoaxwDCoKICXzdBv6OrZf5+gDPQ8DcYSSr4iOnHIGq8VYyC
NKLCIGRI25ERAQl0ASw/+MT7wgUDf499r/4J8C9PYcbPdlVjkRN69r9mDBaYtnIP
KGocYhARMHRTJbR5TKSjCakMXFsvidXwnCWHxgom47YTZ3TPFPPurDp5aXZVgPYn
23k7Tf7uZ+nfoQF1P3awuKwozFfXyXG3yf0khMyXZA2myL56S/WlHYddvrnGEipm
72O/yW26JhiWxA/oJvQ0MAoolUzcnrZfgCRbVXB0iAuII9Mu74UFWklwGK9Xob9J
wDc1ZIpgT2laeyljsFN2z/cAyNjJZuFph72/Lut7/DgAjMVZEBGag+7lmStf1Li7
8wb5ub1aSRD3BDLg3TJxEMW0xx7iAndHoZw8KqcN1l2AeCZi+PQvXdefqnTXynUu
zJMYZbzK6R6PIHVwghvsObYY5gmr1AUOlWdr5VuN2FTeagB5sdCjl0mCU5xhZYb5
0vmHCiXH1n3huPqe5rTvMTj8NGGI4Lc20tE5B73u1AcfcBcyYeQ523TT6sjxXwIi
ijAC/YEpAepoGfG7imo0LmjKQoWYQh584gtCwnKrCCu7y/hDZEZyL+Emepq6F1VQ
Vo2e3j19NDFJk5frc+55dq7OYqfvi/h1KvKLPYc9XXsnXfePi6jnyIXLw7YIMHhn
agD0FyppWwRXz3oEOVd4I0bvr591ZbTMdaTkluz3nH9xStsu+U0L5LCmK9OgBCB0
OWPXwgevBBlyn0AS81r07HuWGpWUuaJqvPvrEoAcICznDEDqoekhc3nQBhsjjQeN
LvFUJIG2p0cG6xnmlvvDEU+4jpdciTWihD4AVhU4315bunrOpDBDNBi+TZYNH0hH
ZpNnU9bRRdZrVnox2O97u03A3Z9XZpkhht7jzY9hn/CmHi6WGrCP+CGNX46Vqs6j
4zeKGH3c1OVyW3nHkJ6jiJdxjDoX9Rdr5ksbGqVImCHYmFa9zFLINeFHnI+ZARJl
Ff8e6LrxjByBT3WyyZO7nxWA+npO2CYSrajnGSx1IDThMc2mozLQfF5dnXYqz9Gr
sY1ZVmcRXAjAlR6IpF9YkFb9Hac6JM/gA2dpwE9Ak/b32pQsZqAkAHfpOB8RhX74
VFkAScIXTlefgwqxFuKpT20fGtCrdleWLShejup43uunZqoXFYdvgHtFyc5Bgbm4
axjh2lHdHBZxl/yBPH89yJ8Dg8bgvXeyIaz6TiZ2DvH1Jhw/dSrtb7B2Hjs0zfNq
Bo2HzM6Xul4odfcapDAcXMp4DOV/sdFxW3p9i6ZUh4NfdNSOCaw8mEuei9EJKqEH
b30ejjzE90KyihuVxGCYvRTRD/wy7wfrBw5HH2ThLYqCUWFTyRNuJrRhv1TZKFQx
Ps+0V7kTm9TXAzKjzkO5kfhJkzXaTwfrm9nWyU0WQH+UXpqdVAxYNSsQODdfluFK
HVLjmL8k8fHTJpI88TLvPQxYyMFGc2OAHaGYYC5y8QZFzqNpi92/8rAqKgji5avs
WyMfR3AYPqbBdZcGrxCYc5rT6teFFyodCXrb9xV7GXiOZ/JbalBCXPnpoy+Au5XZ
31BSp+Lr44LWkECSxLkX4BDQBlOdsg+rjkH7SvbaiuK8pnWFfjg9cD1u/wgPgsyX
58C2UuVTsERADPOJdr+0k4L1CtXEQcuE18ssLmKCbqP0py5rjZPJ/dOhpINLr3Qd
dIfQqS0y8oiiSrJogq2m6Cq7Y5EK8x2ARG5FszPqguR4lLkLpdpIIJLlmhrmnAEA
OcI54CKLnKShVtyyevbEhG7q2QSMHx1u5o6iIU6OANY8rUXr54yEEt5gpxJ4qHFy
UYghoD6Cdw5dpcD3/NNbsYPCgHKSN77WBYwcL+68LxodEM8RiMhY3hZKQAIdfFNA
Mab2Rd2/0xv9v32mW99r66+hsmbj89ZMivVP56ImjLPX/lIYPDTiBbfcSPxCLBHH
MEk+unnfgeSqztseCEw+LLUQXc9KgVZqZ15flw1GTFRVsTCBB4MlNnFhoWFff4Jw
3JcBXhdTH9R2n8WEmmeHghFawTwcLbx4plNZrE/fFmBIb65G0adltzSNZklw0gxu
x9a5ZjWERe5ErieWBeqzI4+xQTv3/xl6wD+4bfBW8R11H58f4TclwX7UlFWFBkXJ
8m4EQyn7oOuYRMdUL/7IOqPbvpvXzMdhInOcYp9WxFM3nU3fbc9DYdvsu4e2dnww
Wdhdg6D15DMRxIbqAUryqt+7ogAeHtZ1uxqN8FCzK4VbpenZgRbvF8N6mPKMXwnZ
0pNlQPe8rZX+q9nD/AGKFoJWGEFYHh80DOFAm6X6lkNoMCP9Aq3rhRTh7ABK/VjY
kka/PdqHqcb/Q4+MMVYj+N8Zxrj27M3ZEhPm5KE6bvbIOM+xiXc7F9cIN6tffUyi
UWQrDpXhpkET896xCex7hg9cL1lNtzOUvDj4KXNolphL+9TJclapOKixhX6ckGSE
wX0UcvKVnWf9iCXp4/A5WVHh9/ukisDpOOPtZtacDARR5/fln67GpV1yt1GlEvmJ
1sL50seFRYFmgMBIrmojHKjx2bd9G06oswb3qzi9kUrlYuNRzh43srzCNl1qLTSl
XtW3TPer9U/03YrvlEvWT1r4w1uNrgnS54tVgRUbW4Al1yhMv03vYMuA9Ba2WAPf
ZWFEqecTYqsS+G8zF9668JANqypCcHPTy0yrt8cFRrtyDtYoJITmNneplUWTFy4E
aTEPa9N48NbEhZHITwPz/sAG3NZLEfBJ7imhUWCqIZdk9MWlDNxjl24hX6i43mvp
Kd0TfzfBDGfMc+w8o+urQz3wFzrgXwW0HL2cEHW20Zj1o6xSPr5/P7opDG3V35zb
Y2/WhEZHd1fGRAtZUYwUYjuiTM5duKXvJTRRppmvtmlhI36QG/zofFLA/Q3w6V1f
Y3LHZ8aHaEBSExAr5Tsbrt64a7K1En4NAGCunMrRtt6A9oHY7iQ1XWaA36m3+uNw
Sl7/i6JNhaxZVLnpqlQtA/fMoZciBn0viDc9vnFoA0DAJz4xZ+urzDNU+CGUIMju
5GQNmoBvZvL6yu53sYiCbNd+VzqwAPbnSXKki3f9xNkKtXILOYPiDm3cvqfD0N/+
A+Ok/mIQFRZSft3CVCN76/BNNU6CHa+/Eydmssk8B3cDbTtyKksNUZB/7YgmMeIx
pRdABQsGsCPyfAObzJZ2cfMQb78VhazfUrrX5WXmiaWz4JIVMXpGmkSTV8i28riT
wIyfjk+MWoBwsAPBKMSSwERVOAKF3LsMgNSW8vNkbp2k5Zwr3KZTmN0PpDoOKran
RB7ZbdrlF7mCyih6YPXZEZMA3h0vwY3m5Ly7M+EwMJtLh+0zRANqPIGDEGSwi1il
aqTJxToMuBkKueLF3FQCGH1wrBvs1q4e4133e8+se5x2wT+aYhDEgYUldTUJ88EG
9ZsisIacK/BFL9xIOW7W8lg2wCzZnyrdczu+4mPAbIYLu9aAaTKGHnVhP2VE7HDI
a9O8wAQIhcRkoI4uQK1ieQ4680WHBKKMhRvskLr24x172B5VpAlJCvZKeUzLiNqi
z3T++aQp/JCC6aAh9W91OZD4CKt+NI+J3WJup4LpGiF4/oEvlKzSxyZWcjXVUEOs
ONE4fsv1zqDbPdt0DwtuQyqlaiejfWp4SNxgXfMCT7tzAXVOQQIilXQSl8N9rY+s
JmfQCeuddIz/OosB1IAShfWa6+tL16x+ethDAw2y/ToOlDTYD3dwx1YTjxglInz8
xEkWfXey+7mDJuHbRN1+PVsCkL9UWlFkeAMEZhw3OoL9UH4TEd2MWWLvVBakj7Sa
WYe7LC9C4NywKjfJxFAD1jvg0M7Hu+0quU0sj+d0yGnxnlZZgzolT8F93BnjTxFn
6nm1U00hnWPTCiN1x86kCEh4nusPzhgBmIUP64n6hVCSOZwIk50CkSn1X4XVyK/U
kQUHd9sBla5iMZjB9j9V9usmI9xPLWYt4YTsXyvlWU7s+Xr6ms+s/dkHTnjAdDKF
xVTu+CAivDqle8iVv15a0z/Ig3KyclxusRjwwCRSjOpOunwH5bN5RDP9RO56RMeJ
64VfX2K72//XwJi3U270jFc2BTa1rl5MsQeAGibaZsKrkvXitWBQbKvikJ3uv7bw
doLfhTmBdJkHnuHD+5bmcHRufSS93EuU1Hz0/qZgJdD5o4VzIkBfGkpPYdkQFhsf
yyId8dtkuqkAkWpyxfxpHjqVjHxoU5B18GMlJypymmA9FedHfRmTMIOZs4autEEF
3BU14jId7M6/0HcDbq/YufUOmsapNRIa3Fcqi+enBQFLqCviqXTgjecAPzaaMJ/Q
zBlCSdsPM0VBdkOXzItK9wxT5KULFQlkh5+P3xXc73aisoUi6yOEMZxaaIrMIcX8
ngE7DA9Zy8n2OpQ5nrq372D2otAafL9TgzpIrdNZMhIJ/RSsiT3Clk1TOOXpjh4s
80nVxBxlEDSjTmpNSkO1Cvjm8Yurmru86XjRknseZkqLG6hXfzfWkq55VJHmqxPw
4i/Q4rp3YU73bDtlokKSwboj9GK0eVTESVIeljSuUVgTK0izAQTSKcJHfqS31egQ
xdiNmo01ibEaWihHo3/bfBOHPTzqRHlLJ8DBX1lN27uF/iSsAV9BmGpgNMxaepwC
ZB2kyQ1SoZkqrI+9X1Qndg3hSFYfYcCMj/Ykb9K28QyyCc3YNz8KkFPgoXZsuJMw
3uQfFdZ3gCx1L7Jl765BB2KSl3VZGl89/yfegJQpVyH5ElXsKkQZO94m1j7LMJxX
Ptn9ZT0lVcSgCluQ7z78q2G6kB63KIQ72umXCxyJhxSsYqUANxIUlDiEdgMHsDyE
+J9drrzGAkJFnPG9nLESdgdUt/frI/YYfW6ugLPAA45+xhsQqwSKTXu6l2s4FKT8
a1jjqwyKAOV9dWaqxoBIOmpOkj/3qkhS8xjmdboPJsXvcbCKJGN6C6b1NllFynXI
1uLFR6+NbJrdv7VzAW1vbN/KNYm1r4gLPIpwKoLVUwXGrnnM2ZAOku8BJJAt2BpI
2xVbhD6IrnExBIt4rqW8/qtYO3wSMIMStbI1PVm4qDluBovD6uWSZ9y4o/CDcrke
LwFgjTIDCbwfZIqgul8PFu7uqu8QiL7K4/RM7+PbvjZz9xbUC5AarDQx2GO9d6Xd
ichnG8/RwfgyyBawPEOGMBIoE7OY+HFr53T++umoMc5DZy16b/kZNU1NUMPz4McA
36dsYwF9aj7ct0RiLAb62Rf2lHpwRn1i+dPBvGC1bPdtmW3khyca+h+gXcRK4PlR
hRDK0ozkslYqPfiuxjMrW0jD4LS8p5T4WBlknjZl/HxQJ9hUm3wGqnrLgeFYQEt5
PNijWi9/pWhOGaaOjABvMoY+mIKxndz9+KjUe0xB+7GY+UfHt+Yki6t/YubDMBLy
fNHJfUt4qAp/IACUhBmjOSiOb+xdwwVob2tAlnNG+b6J7DAMopbV7wdgJc82vHom
12w9Dt5wZgn6DTtVM6zdoXP1/ZhH32L+LCzGa4xLhtZkOSNqyJFCfaXQCJGxHreh
pIdmta8iWC+5OSiT1IJezZfG3GFvVeXKAoVB5sE6SuZOU6FDgAFTDc7TBAa1Azuu
8393No73gDQIE7nJOsrX/LrToK6VrdU1GThj/mA3w2WnUe5PG4IR1duDlT7MLl8g
tTPsZu4ahO/8t2W7ZQf1zQWJ+kJgli1yYSHCp0tR9kVIhWNNozDG10vxutpePTbh
BzWxBqHcViZESNOPThZi8+88FoDJdBu0DZjT3UU48/L0Zws2Lbv3wqmdWBJNDrNh
FJiPENy9Pz1jozFWKj/q+BZdRNzV8UxJhvAexiJfdmmPjGAT6r/8roTtlwWrPi4M
BLk5hCN2o2hmDc+o+T9Chc8UlS4VYJ+uqJwNFT67TIxoxCTFv98WCGlyWy6lc6fD
JLpb3olCK4YoiTKetpKIVUVbviZp/bRhJLB+3iwFtJpidYnnyGWwv7tdKdgtZ1pB
EdXbGsPztGCb0pkP1z/BMF6SqruHKKMPRKOcjCYG4oy9jtwiRZSnhVvLrPqHilld
iTBo8Euz+KeEuJ0PovWj9Mew65rLXI7ZMeyCqAwCRrxzJUZS2y9ELPdmetmQOHvN
5HuPKf3pRhjgjgnf7IQ9GadeLgQjeT9I21zDJNzfyGxXe+QKaRsiw96foSviMivL
k0o8htZSe0WVFgl2Kt+4Qk+CWBnaOZjwzCRrVUtX2ojD1ixEJkd6otSLNsgYY1gT
B2lflR/6wyHNjZJCcKeI3HDmpR89lgYhQuI3YCsJjFLzT+aMYjo5P7RchbJg9Gqz
2UvtJEOCEA+KsJbSTvfHclQHhCDLwMuDT3M9ewknO5BVKFb83yHrp4YILFwB6teE
H9XdWG0/X4R9LCySN7nAN+qjT6ZJWw9PglM6eyT/3k/9oXKo6iBYOFu+hOD0tgW5
Gli9kPS7NoNvR5GakP0Lnwwl7XyLoyvKDwbwT+KQ70oYW1yOhQ/Reas7eZLWgjyE
PinYhEIlzer+zCh/gGs2RUOBtuRKEvlQfD8nYy75lrkoKnVaTu8N9VO8Us9BZ6Ga
WBQip22P/nrbGt7siUU2XN57Np9yOpvA+Eo6VjV2y+qWB2o0fcvtdMpLOzVOwNs4
BATRLJzHksK6Ka0f5VB8YfrVGm5twpd7HPsfFM5+ZIgijBR6AJ8Gxq7wD9PbVqMV
wd8Hy0rEOoHX00TSohP/H4zbleU0w8renoQgi0fWodJFRlVv/S3EOKKPWK5CjmPf
iJgkDVazdYNzAutpGrjFQry6AxXowZIyKeC6c0ekEjqWR38D4iHdUKjx6wyZCTZ5
zmVCGRsbUEmv3NcFmed3TO2tG2+wAqAu4d5DV7sqr9aw4GvwBkF8cRZrZ3wKum/8
pd/BAziboyCGs93CEUL9jtuNYX7np+/h9OHXh9YYxV66k8D+XeOB+ZKxa1Jf6zxB
xkcfKjtGcwubBxGV+WQ3yTLmYVmjlJDZoElDkoU86wvn4CisxW2qCMquEXAZpF6w
qVfrFHcFdVJU58OIYdSGYnLdT0oerzG8Xk/QOwjILZP0tX/2/J8x19gv3VDz4R9T
AUl89nXD0IuiTY+iguYmdZ3sHTjANIQWuyGB4hYRPH5KfVvB+xp4Feke+eOgQ7W7
ITlcHoq1/I4/JTBwpPnE+dPOopgGNQgxYofbUzzWk4s3rJwucusAXs8kZGbC6GUC
sfXYQetzUOvIt82V/JW+I9gD73b/rPD9t6EwFVVpu2BvIT3F+nfr8/RE7WJX5Y+F
SP07ei2D7KeqWKI2PvXDKauux1x7IR9cN9vkOnpijlepnHQPtVciZAJN5+Fdwxa/
js71Ao7hFQpQjBp5TgrFWhrTsC4rbsgmzF50Fsrq9PbB4Hv9Kwl5QT5usQJAtf3b
bIEES5UV7G4rPyi+Y+hTc2ojezsxcNOV4vS1kr+zY21vOO43PI51w4uz7xvvwVmS
t37aKYYoTLZJ6m7sD78hspHuJXW1N+kpMTpUHr5yOL+4s/sOzbn2oR8sq3qir9PB
5BOSt5rot2wgBkgatorlJI2gqgGbWUB8icXaOEZiPDAG8sn8DOl4TvUy410J1ell
p0nBgd9h/SHYwkgMB2uOeQxOrt5MEAo9v5RNUnNZkropX8FN/5rcZsQQzF0X4m6B
MxT5dqzkoZpsx5F7GyMnTMDLza0OO11cJ9ne/KZjzp5aDtKfA5Y4zb6dzQjD8iTh
yp8TRvJaqHC/V2g/+oCgKNbGd+Xa7qqq1t0kNCyv4uCDci/Gv344b1vv60bdZNT3
BpU9Q+xo6UwiQ8zCNGU8MWmLYprSdQNlPbBHNlK+aMA7r2T4WcdP+YRD0v+szAWt
BbnnUloVlYh9UQB9ewviGLBCNylz+L0zdv0UICwMIrAdSOsb1S8PHcQgXHwZhW2m
Zxvkqe3fJ+NrlilMZkfMuLqhiZOcya2j5aOHPhs6FK1C/o/d5hBzN/NWmdWaTBJN
koNqr5pCwk7SSj+rDsyiragjRl0Ip1hvI9vW4n3+S0xrNja1hD3IwoNS2g4GosTO
/6CfN13Yw9OH5QDhTKcUdA99rorehaLp4jl9RFMUHPm2pTz7SyzC3D15gORSgHZw
gby1vJDxpg1GkTtXn4oW4hkoDlmW/ingI8dw8a0XrlU+E8yv0JWRIwQh3mRstdOA
Tt9FaPL4AoQkuvJiacgA7yjpEK93qmLKSBhmbwSwXiI5BeYsRApZ0wHcLA4vNaRt
dOvtMC+VAxwo2NKBa1Kr0qHLeq92nfk5Dg0J3ZUUh4rBIMnQm2lv9R589HdNpnlm
78JSWEET81rDffecrlr4rlHosZ2zck4phoko+0NurqgCixOZ52pMaMmo52fJtgmg
czUiR3fXd0mbAJm8Vjw8Kx7buGEsVY6IpY4CTDnBmH3wz3OIvKBsZbYRJRYKGx+v
erYo5ywXj7+EoMDE3BL0FnlGege2d/mMWxMZN/Uf9m+kPeZhzWJsQ0BELd8kmWfi
BIsZ7Y8Z/q+gnyrTyyxBibymkL7IBgnvLcmbBaDmys47DJ0uhyXgDxlSuGJHWUVs
S11a7aKeNlL6AIkPuXk2EQioeDQnG8GLG6GC4DY/EgfGWFPW+uCWI55S5CFg/wnk
8iZpKxJca2Oawx93V23hv+fWC7K9+RMI464n2RzA9Z4u3Osyk8uyzV4Dyy0pHWnb
XaNrUUTuOXcZq9oXxzvolWXZkUXpXoK+OlUIwHg8QZCrhf/Rhhu0UvM+GX0PeM00
8P6bDFg91uR6UJ8ZDDt1SuLAcdk4Q8/7/E73AkdaPX9/eUqtKJlV/e32Zx5DiKdb
H4l8Vo2xCSVbhTtvBIglADH8MwH2QEGDS+mLs4agiBWXKxVXJyuJ1NUV668DEp67
9pLj4H9LDtywD+rZCyIK5wkHS0epSG7jQibXmmEigzC/sHxyF0rECA63cgXI4Mpq
eXzUOCr8aWMkp3wwKdMFngxb4SpJ8BLDL+xmJjHNMXx2XpojzTJnoCt65BBa6FOy
xRGPuQ9pc/uefysmPWDmiUAfucCrhU5froqvXjXi2f7DPbPcJjjKGR7QVLHt7tgI
rUZQQUoYNW3WvTfUK1vhnqjO2l3b7BeNYGuHUfPeNKqzQJlVNqR27yvTezkZpq+3
YNeCktqsi2LkSM1KNElWD0Y6Hv/rj+SLQOZXB5YwZmNZfhPH2lEkPdpVxFAIO1Ew
tZ1ppPCzRKeWhRNQfwRJ4XYwEV4UloLNxUNbMN2slV7IqMO34BA7VGS5Lc2E0izW
oB9LZUcpjFxMJ16Kwkul9PF29jVoovDuGatPUJ/iXYlQZ+tdglHRq+chkPyMsRLO
vesXm0Bie94HUZM233pZdCfhaXI/AwwfYwFDlGGH4rBV8+LHNBzM7dnf4hj7ux8f
HtiG6PgT0o8pt2VP3NSyXVxbbeq/CehZT0Ucphk4Z1e/b7CcVfp3Z6t+c+3P65Sx
Qc6HMFUfiiVE37e36X8Gu7OZDhZp/ceiQNvBHujsahi/s/QOpnYOIrJTla8mjXEH
lU/fEbC36i+XRwCq6QLCaVtyBM2UmPNyQjLF/Yh47R2C8+McRD1kIk1u6MWGb97O
ed/g+G0+pakT5XSQdDjVTQfGPbPM8cHvdQ2WRjt/2ilrrrQMIb04qts6v8B5S/6q
Eg3OmlMlgHywKilGRb+NHS+Rwz8DlUQtpl4Y8hbk4JOVtbhjNn6IS0MpHfUKfRUQ
pce1702zNihfwm6II41ppOKc0EH1d124bPldJHQk0ctwbTdj13THnrOTI1NjcSHd
N5rK0iSdcar0pAB7PTEv32nH8WCJ7e7i+TdXaB6q/9xjdSg7kiHlwzvuIZUwQHJ2
syNydvXmvNnK68l8w6SPiGHPgVMYjGcf+XQ8INHyQr4hlTJXoP24p/qB9XwDja/K
UyV9YA/rwdvkh7BT1tZ70UIkeqSZhHAeTtC8IMLcH2feEsvS82SUvnKAz1nEqoex
5ZyHWVaGcHU/ZFRm4aCTOI4pAvc/wvipRYkbTrFWc01PaxDj+3HwFAZD1y897UWp
aEVlVWf+YNdZKLZzvR6biY2TmZR1YJK8RrJi6fZ753Fv4DbIAiK9bJ/26MeqO+ur
SgYmNAMWu1jqg73k/VzF1gAuRtoGZ1LgA4FGouHYWr8S155+niVg5Qtpy463gyS4
4CeWGgifpu8kbz4LbJW/WHe27eJwMYIEO80yiOcBsECY3OGuG+t9u6rFHRDnLiY1
CXtUid5JwWT87qajkNC668LX60pmJ9S15WhVtgpzlQ7tMJeRetrRbjFUTDzUxv7K
uH2ND/8q3BcQtdf+p+9bZv3ZR44Bzyq+rXgpCVX9jt2+P03Q5S4qZaRe77W0lhGy
WXW4TQ01UKuZ4K3Nc3pVTl0LxA8GkgKm5GHrzSWA/ZR2rNWAKV/6nQyD80VTBIpC
Qjypuw8SslBfoYTjGcusBtqXDmQWIyBYyjyEHpJHfI2RHTzMYvbD/DDSpUk1i/bL
GJ5KO1ANbbzYuG0PenF4KupgGcR0rtOr8NDt7o7TsiYCEtZl/zuzJPUmFpJ6caMC
JmsI3iR880fpoKPEWgHosIkMVTuW1TiN5xIp9Qs7Vyg9yPsyiVQG5ly3yu4a+00B
Otfa6uwKSpdgEAzDUG4AwMoxrlKLUncAELN7C5RXlKlNzcn9lT01ASon7NOA9mgs
jdVBpT5seLuOYuJYDIsNMu0Tx5Q3XpWzIskKDZqIEXQkp3CyS0dBCM7RouTluATw
KebyoPTiBly/DZ/aUszXJWn5bFiYMi9ZosCRtFhpehvnkdELakVaRaXJefdfeliA
82byR2KXh2AEZSht3xIy8vyw4Pi6V65ekbMm1HLd/ceRjgMdCay1jKyhSA0jnPiz
wJRatzBnozakRyk+gC4R5UlxNK41qA0VU0r0rwZXjQ4BZnxjrajSqFINM2j88wQz
rnfpPous/TwqtZh1Eax9rRGzC25C3MN7XfRyn1xe2ngGL4EtfRKWC+Ces465B2n8
fMhsnj48gX557PKQpoRKQ50nvavOEOV7YjD1e7QBmqEegnXlHUFljzs4Z0VJLaWV
vsQec/bYaXtVabDt/4TleKX1YGCadkdmhFuXfCzabwUrHp1YTP95zBmvkrDAFnPM
HPckWNrNK2WQeTAuyibf89TQyfwFq5lwq3SiMxnTrtkMc+g/Gf7DoKANByvUqNka
o6fklj8GcbirscWMXgB+Rsux5wCT2BCUFJLODLSZ8PSaERzweu1iRXLNCUz2kqTx
goiYwc5TEJKBd5Sxn2Wjmqnwt9l0y4fHRbfwsFY45dQeTmQDJj9GHZ98MJPoorfo
j2mnjpjokMMqspX90b19fpN4enQXrAzIsBCTgjxucEp6nRKS4ZLgC4/tDnoR6fmr
ZWzFwBMgPIF2nEMleGNEVdroqQHbyl9UO7n2s+4M7wVMrQIWorfVDpoMLwcW/7rI
hmqVLB0dpS8HjPmc6K3EclEvzV3Kbapluma+N00Hpcu/Nh5MOYuBZSBAFt29/3oc
Xmz8QfAPu0gGxUSNRNlMZty2bLVADDldfZAxIg8Q5p1Klfdn2td7B+dgtoPSsVGS
/nWViR6Cr9OgSWeMhM9yz1Tuuvxa8nQgrOup81VL4t+cRpIh/71kDCBck1kescz6
HGRf8JHHnou34BB6EmgRvluXDLYsvureWke1Zr1+Ly5roIiNodupJ5DrYtAfQw5r
hi0HaGB/gn4c1U9fkaIMR2WySrEBK4+KJ7C5DqLiNw88NxXtUbW1xgpgraiTJqzT
cJWXvxbj95AnMbci/CYanDRPo9Hdf1Jtdcc2br870tuYd9c0PmvLu9imw8B54Xvz
h4xRCECUFVcCQFbsFOOCtFQ7+0BE02kdH0xquDSKbdQsGEYqpMp7ZqO7G9xYo6Ko
k7ZNWYKEq+/gEpn7L2Uzjj8xjgVooWxyCrNw9wFjd9RYH4dgd2/VSt1tl0lPOQz/
AZ6GFU3Znl+PwoVV+v1/JwHuF4Fd7U45B6ocxPVPwlgQVKhGazAFsK+4fPZO9TLT
xrFnpwiWRX7jXyWsrAs5ibHHnl9zTa5EOvb94o8PAZYaO4KadpZtHaZZDUPVa1mG
dkVM8Z/YQawLWgq1DRx7b+XeqGxykgoYLsfg1lhJJpVIRkUdT20Z70Vb+eaGJVzi
tiefr+smIDw+FTLSxQtDimpBZ9Tb414QQFWUCfauRkxIEgxjfkoK5GYCEgK5lo/j
zyFBX+mgGD/yFPhLOslcGKXpAAlUhRzWi18UREjTvdttzOsdpnYH26yUr4lx6jFv
UxqKO2HEIH2vVwK3NSACyIr5/eFrpfMdNr9VoO8Fy9MDTD8h47dX8JGVA59DYFxC
9ef6XvHitOKmTbYHjX66d8M7CUBY1iUIfBfTzBkRylWoC9+XPOOvHPZJIWV8lNsB
hGIeSsis2NjGwEibqb0UFTgAipdstEokXHpDR0i7L00JB8we5ENmT8SXu1Vh4Dgq
S5rLT6HUGAYFS/BAX6IC4Y11rjWpnXB6ACENSnSY95kH1tkNXPMtoKjjptJc3O9K
dzOjwUAj2IB+PJu346+8HGcfCedvVJZ+M1tV3D1DcedNU6fkGbhMvxo+8aGRMH0T
PeyP4yYRmUEWups+3ix/voPkJbpS43ksL2mOozNoauN2Pui9GdcPr6cC7JiZNrnh
88WAVhhKvIIJp4eXY7kTrkiqQ48aR3CpJnoHjK5Q8hevKdx5XCiYLQCffb8MbzHx
PHEqBBRQvLBYuGyIQFl9CcdxOIhiFwZ4kYKi3PGzp0/vymxN9IpNDZ5WnO9VXraz
94TJfROS48avCzsF1kJ/ije4+qzsDlCMBrtAXOhG7VRZmdzFdcr5MsaxHr8AMe79
Px7MKAQiKu+oPIRAamOLjJLMhIRkx+fUshpBsikCtGb0QOgA5eBEPn87kJ38PoT8
N5CvZ1XJetsqIz6UR/oGchq+jQxOlUekRMKgEmW8HPnslB4BOKu3OHho//w7y611
ANFqRNMJVECS6B0XrW2utO0293Xr3Ri3s1nxbwdVeC0GZ5VCDr+Jh0CQzYocKNY+
6AigIZlf9DOW8EEldi7Uo1j6dWuylxnk2LzWq8H/cHPrwZbRLOZeDbE1vsxEQrSo
9ensrTgpEGY3lIyCDyNmUo5RaEAN1McTFg1ooanNnSNg/Zdr5FIbaviYpIjXftg8
6aZGVoONhOF5lxfP4t9Pnd4Tof9+YL7ZSF0rHrjO3Ek3aMuCMzND8jHX2lXD4BQ6
DF3F6C/a8iMZe9L5v4KEbEtGB3FpUWmr6GSwOemRJQ77oqaZgV9KIOecrmx6lfon
Rp8GwygDqfiqHE6x7prcGHVVEjwitolnoSAL2Z483vWgQtl4ShRUiEYilzyfxPUk
214YRjRzyG2Grh62KqPyxOHGQsTGVrtZ2KmrC7Zg1vX+re6prX9ruOeuLnqWBd/6
NR4PY1SuIK4bPb9OOfS1oni+5XhroqsIg9toEFQJFKmC2zOiBuRdny7loJpyPslc
h/JheQEHA48CEiMc6h/Fw+V+xFlRPB5DmZqZCzE7CC7Flluw7mHKgKVu2ymABiUZ
7rBvKaFyvCFITUA7Q7V8HDMssZgsxYi6xFJvAS9iDj28PSe5gvCXNr+zpt7r1kd1
1F76/N3ridRtdGzfM9lSSgS7jpAnBpXrRVCXnXqjjJQZjyVz0pKdFKQs0uNBFtUO
h/UwGyRP1vT1THWlpNs7bFje+s/Bl/pCj6qNjbGEqqWKfPFr9WlLsdaQGUpMPgnv
KkkCqBy8lQ5l6B/vM7C0/b8JEEizN4lX2+UclJhl7Rjhyvj5QkUj2Dj9PHQhUQRh
psFEmRQytidNXKyzhmo8pKDx2yGX8qYQIX0FZgLWYb54/IpoMifLa4BdyB9YDFZ+
WCQ4Dq8mfluzFDg0AKR6GzBRZQUmiPfxx3IZQZkT+vm+rJ4y7cUdmY4Dw89whCLX
5KCO9YuN7VrMyiswJDOrvZtpquwenQfSOpGNuTEdAS8s5KyArsUkD1asaQI82QvO
yCd3YjNYMLn8WcpsPDLs6dtd2H6jcNB84x42HKIXvBViRXFCtc/tn3Aa07D9DqDR
nA+BapsRkl9nGeiVIcZ/mNV3gLOt5/N+YvYkROykoKUIS6shilkhZQDVpPXpaxMV
z65DIsaf3iVFQTx9bS9PYmizdGe7JXUn544NHNMWl/nGXYCfcLO5bSZQn05dJPIg
1EUX+DiINqdiCEQLsCUUIB5TCwUA5vsMz3PDQQ8IlxtMRdne2lxLSzpEhWY3xY6f
Zcms1WXILrneoaoTWtq4Q+fOZVGp5lpKn9KwSBMtGHCGGBF9vuySBZQyARWAMg/V
+WXf1SpKbItubeorxcv+mwspXBmZRgrdod48P/Zari4XXRqt4jot1VmFdI4JSAN3
aZPYuSd70+kwH+oUoFk2bQV+XNFNETpZffCUivefN3ivpemDIp9PWsN3cgeYKgMv
9TZlF6NeLRnD879/N1ZPxkvVYc9uGHjhC6W3jKPcdiwB5hLsi9G/88+H4BLFPn+u
zgycWjWUfUSwsHy5vjxg3cgy+iC9BypfvmJUGjoSCzvJ/GeZT+Y4ZX9GUQubL4do
w+soI0XCBecQ8rfxF72Wo5h70JoFPPcZPHpNFl9KrwWEdl7jgh919SRbriDi9Ldc
IprE8bPbRdDm/FHIEAU1ifqdDLDErC4Jw9gLno3gRZuOQ20rUjM8ewuS+vHrXF5W
1JQPps8AyTJRfzLc7Zjtc8zs5Z7IUE7st4rCoEW1iSJAzQ88QNP3az/rosbSB3Hs
0fv+oadg7oxX2eSwUrWcezVSJPfpR+lRgzdg+H8qCzuKuNroaeM3qdUjk8fGjY74
pjjbH2jbMAxmaicDWg/gjRIdHYH5eYRyZOiooG7ofe/hnDQzvXZ7XxAKx8P/Psfe
wgZM+JNdB5dCWwLBl3fFiOh30bt0vaJfNMcyZeBR5xqdZNYsi7obA9C9tNtyGm6Q
GPoeMLNU9Jc6U0H7pDYBFQgTbrX9Oy8LaeqwXwJWz/JGzB/lcLOotDYfSgJjzKEZ
z4o7igAm344LYVTJgC8ZNg61Hv+xsvp8qkRcVETq2UovfzeUI6yfXAOcumjz1REA
TNJt34VEAU+dATvjDoEr03WLmvnqfVhKdalaJvSC2q237m9smn5PTm/hmn9ZUtMX
0qNmIiE1V9McfsnJcY82D+1Bcb4Xi02BH6ZVpY7Dv7icsbPckXaO5MzcdpaN5sRX
WeHVlz1fiF4b/b+zFi9ooPM/7yT0GE1+6O194Ljwg4A7Myy+hyu06kkKHvnjFwB6
y0JaDvtYr5Jajl9Lfha2/4dq0dtA3kgZMu48H3Y77NQ7bAhW/Cv66Czv/ZSFMJkG
gtuPdvNlJ1XPI3r1wNtfojETMEKIQMd6PSCJxWxwiA21Dibxhk7WbmSyiRxd2MaB
XVD1vJ77r5Iz1oUVeI879Kw5HBTXpBwSJlPOS6xPDGrPVf5+CPyq2TG78kRk0bKY
LxqS4gkbjTfifq5c5fXg288ICF8QjSL7Bn58pc2v6An+1L37gLJaNFbA/iBRYD3Y
Ylr5LqyoJL/6w+GWelV7XRBvxyn5IlFZphXb56x2U17m6JUNt31Ixyn9Bqup9vEl
L/6IR8d6EHmzUsiI+7raSmjpdrTeMCo8qJSi6u22yhs5f91Pjllety8EUlaPt+TJ
6qbGwjQLqhwrPtxaAnh6rqKsx6vUYHPuBXNLdla/h+2STu6tVOE+9TcUo9MbTR7F
QxyqC8YeKk95+rhoaurAK861Otza9/4XZVYJv8v1AC2lthm3fB2WLN6bQvPa1dte
Iuy6Wu8T7pXuLmx8uBFHvw1NIv2v0j4X9wnbgr/j+zG9BDjfFetFeYMQHjImjG//
q+ZZXcHcI7qhEDn2Wk9y6DuQLkWE29Vk7qpSafsuK8HjLKml6J1Sy6tsjzUG66jN
srzNkmQJYXwCAmfRHeQDdRjNgca7AY4/tEY/i+b+HcS2xpr6WoRL/csD50eXddA9
tnnJaSvPT9KBHW2mKVUZma0ghwE3MonLRVXhTEnk67r9AlqVm0bAyrF4nBHVKEKE
keqXuqOfR7p+HVfeLoHycnDtU8U2U+2Ba4Akgewv4QnslHnZNsfIh6y+GYYwXb7S
o64Fsow8nHd2Kzsl74KBHDGtHXbrUQwLbb/EObRGkjcXN7qeEeAhos/ecpxntwZB
rBJ23SmcxdVaCLG+cVdPDayNRMsh/qaYQWPA3czoNvkIa1Yk59rSipVQ2UNrJz1Q
i/AsXeyX/rqBDoq9p6WMc19hu8hjt00SqHGtHMDZaKF1dNjEt2GIR/ZWw4xBa91K
gBnadQOfUvjqLLGhs6j6rDl199d/8yftZqRE5ni3/dNRGV5mvn2axjXledJWzgUN
NKqdYheX8Ah+JGG7Pf3RA5TYiZOnPrBdR0N216HKFFhQV9kBqCPgjTB6lv7urSOm
Wgp2HJ/rrS2iBt9mXrtTVEr43C7f4jXA1Iz5RfjLNWTvi5OHYLL8PJfzg8T3bEMi
Zj9QG1KRBm6oc34w0Q3HCB9POgm4nrZthZRk5li3AwP9bqJKPeiq4keXV6roGBiD
P+Hp+o0oK+Rz1VO9RDrb8y42dNHEdRMD+6ThJwPMrJcGR3exE4cCHNutF6YGzqqC
naUBTklvrAs3DMD1wkJg3KZzUKBHYNiP/qjaELZ7sb5geoSSBfryrcxoMR67fsBr
N4JQ8yScCP7XdVUecYCTnUVZgXIfvU1qJhoVAKBTWAxASNR5pAkuwA7PQvB9+GSt
O9dfi93pzyLC3U0hCHo882cay6fgLElTt/2kcoW61cYiKim6SaAs4TATJFa0MsRR
hKcz2c6AQbr2asYCBOeYbTje6eW1vf3YLlJAOW8WPAHguYib9XKuLqtwxaljo8vx
itBIHIYO3a5JDMs35xB8YAhOgETeEB5Vg66VFmdUxZEEKeLlqSFVqEc+eKIWwq+S
fWBGc0/r7ChTFrra5EOiEq9/BKlymRXNXk8WsBQjlQnHQfodGet70h/W9qbDsUcd
79z30OZ2vYNkODfSiYE9qp/y0x3x/1/WWAkWi8cxUOSjQaiX9M4nu3k31LD0YCx5
1u0RToA/RHlTmabkh2t0lWi5Gkf8VX14RlLAIDHx6vevRfAMiruQH4CxPLIabh9v
jc0Zpzy5bXERdTx3rXq6fiFu1xOdzB5giHAB/LITs98KLQcv1DDqSscoPq1yvynC
pJlEiBo94b9waSuzuV5mUQnriFaG8Lza/l0wR/o2a2zxFLFXvabddWH5EG1X++g7
0/P7iBO+w8WO0bMuNKEAB5IE2+2Gg+tnOjTAqYzzv/WgovvnlPy9wh7PGS9FWuKl
gxXMzbyD4hpRfZl7u+DMubGntUtKST55suFQLK3KNCdSy4R068i6q+CWwXf90iKz
RZhUEk8pBfe+/PxXguSG0jeLnGz5UrgiPfk+swTYA+zKmJ6pcOU1uADFesSvFCbR
REWSKDs8T1gn1xcbzkKWIZqKnux7CSopywkjGUvMxSiPN0DMRlC/+ATvvrihw2hx
+ZjsYYyanwT0ziaPxSXX1uHbVFL+n0uDjXkFNWyVlhzYlni/8SBl+MNwWQnLPR4f
BtQEcsDYmS5pX81vdmrlKYTArwl/sqHP3kkKC6q7XBrD+0jVrAf0zQ2D7sRTjoyW
/xdybu2rwVWcnoTbFbmVPS6XL5EhIs6AA6G1vMw0Bl9y6wK0YBMINhonAJlB87Hr
A37wGnQzdJNGhQsHoadjW9nYR9g9xwBsukhBlMSFS3JdI3YhlPj3Dpnv/ME2o2tp
BY3guVob86/rnAU+/M8OvaywsTXyLnd6HlotqxT+ZBmak9EnfffKM1d9tScnUeda
Az5ZVOC7jI22bCG2mpIMi6IbECPhcRXylqDbVlxfPAQv7SgnCN2u4IEMLRZdIXTy
/XNmtjMb47K33FiByb5zwItvoNsnJNMk7OOPW3YL3SQgWoPxejPlJzWhL2zW5t2z
UqfN4aQNKAcICXhl5gV80wl4XAQfcxtx5t4cSQ0msqtqlNisGqbML8fUB4Y/3eLT
eCUv9iF+sR4XhmYEnc3uZaV2gUsQ6hsjbtVqc0Ab6h/+qt2wuL9G3Z+E5MpHazrR
q6rQoApgdsEIrfJrYAv9tWpTlao/iPb1mX4MEKyd/NR5OpXaUrW8xdH6cW68Pyf0
3dyLdNC3g0es5KYoypocU61YNaG1J++n9utEQIGf06cHV0a2Awp5CeOVumMJI8Rp
fh4rU8GdDciYrn779ZcB3XWGNry/J/nMvlC7vOWsNTexce0vPknKkSw7pMDmWjlI
BwaRUQnRb7b6EWtb3cwOdS0yYqouqLhPR9zmJc9B+kfNs2j7BDctKPKhxK5QzsDF
ToH0ThAHfkQCl5sWpr0H1mks6UZ81rw/Fod2Itw48crheS+v2zViSS450Y/DP5rr
YhsTfVBhDqloGTLlpAPYVWfz9tB5Brm/N2ArrQ5wH0OTH1kjVU4JrPvWKd9ZShjM
19T31Z0PRInWm50XsdSAFibW0hnNVnAleIqgwMHML5tiKnKNXrJOKJAFz3J75FTb
XgJdxloemqN8ev3f+w4VG46tCayC5gPEJFb39lc43l7CbonMDwJEMOv9YrscPvTO
T0Ke1EYGx4wzbvxz2HK2/G29rdwIN8nk3+tfJkY3SJ4Ex6PndTAcCriYGBkEf8vC
GF/F2CY5t4rgWkiwmoh5/N16DzvTK4rg4uxwEeesXcIHDC++SXe/76sdG2cBsUe3
5Qk8EZ9KfxzFaD7jtGdGys64cLCafAFa0IEJkFfofrjrFCE/u6kCTW9Q00eGig+/
ejPRylrxLagBRXa8wEWgw5RReNoZ0RhjqqPZIavnyyjYE9vmfMLsrkgBG5TbsEGv
/kqKpW+uw7XjnG1yiMdAC2XY16Z0XLrSMxPRaGjBJwepwN9vVR0CI0eziNQaBUhK
/hmUqbjdmU27hmOQ0VJr3Uxh3CIs5bTWK+L42A9tIWhLiV31klPv8la7jm1YPPvb
/XFZSnRxQrxFjvj4glSzRzjVuxK1o/5J4ihqUOLzGhe3KM/NoDil52pOzb1vgB5z
xEYILV/V3shTHwKW+uDBaFsSEboSf4Fq+hgI8LrPOUOvBpbMGgjvL7HMbomKZ+cR
Jg8K70v8eoH5cd+QxHuwHAWeOz2qAbfWghgUEdRnXXFGy95vPNAjl2eqUsjKqPEW
kB49R0iXa2nfS3vicRlZ16FZ/zmWAc2r51ZXVmba1qkFXn2K+KEbcOYdH/nCRNJ4
1ELxfHDRuljlIHyQPJrm829cHsWK7SlGzWPWWKY171zxVuIJsi7mHxw5TRhEBReH
/yVMsKM/OeoLgTGHfEKFIe47d83xhkfL/VhFe0CYLvFM5h+SI0XKXEnKasjgJ6Pq
J7Yml9QzKEeopaQzwk1tsk/QYHe8AAN8LEy8QySzr5b5Grat8LA4eFV0SSLFlDoY
GpOuvX1pJMajRShQWXtjcS8tmJLq34lqSygsf2yR0i7ALAYsI/iOOVBr5N7SM/7m
FEk8TM6dd2ab8WObHLhbnot4LDj7mh1mTp4JcWwNnkhQkgQTk7pg5GjPss35RD4z
agNJLtxE63fS8TcgtKIfqzX3mIwvl6DdyQ0ajztOYih0VR/+hHif5MmbzhSYjp/3
mQMXSAwmNy5EWW2IBiDGyA74KMGkPNck362cUNOeWTyr5c+/4K7WWiVV0JRyupBu
SMiVKXvyQSw2T/DbQ/aWFyfAkW3HzeUq0AQp7FtfixE4pxR3B7F9/nHebjSCuhbm
oDelDEWDE6QAjzFxHLzCFIUfUagAUtKE8C4BH9mQjNQynCeCjZyLnPzKTu3TYt7y
YymKA/kCgJeBn0z9hOOYJCMf+WUBWO58SJZ5iVkmQXdcNYjCosFeJY/QZss2zGuc
h9g839SvxsoFiPZyVf/kfwgsCLjh+f5lXy+wQrSOxsGHwt7aVdssP8ldJ6vzEOWR
rZ/9bBt3VhKUfSkhYO4ONz2DHQaOPu+Or9Df6PD+TH8F3w6ek9vRuI6TlGNtFNhH
5Nbgwcbsn+ZjAFM+1ugUR4bReKN7q25DWIlRNt7JC2tdRGYMHwuhp2XtQwXCfjyD
Cz9cm7NPr1moRchiAIg7/W+pCJJ6R2hCMsTyK3AgN5fUqYAssrvciIWkxWpPsg8x
50a0UFfYCds8Dab4Bvvs8DwSsWrOrTM3tN6Dtnf/wk6q4paEaetUJXT5N4RVIpiP
9Xpv/J4zT6PnwRjDNYDu6HM5J5hAs4ub+V2Zb1Sxadaht1zj1vT6YqOVFlCoTJl+
H31nnfllRP0u6aXKmHBGw+T0JUNjN9gQzkK6USD6DCNeeLknb3ryUiFz+1I3VO6r
2mMYJyDkNQmMJlWZqw+NxTVr9Le5Wku4UdGK9Co1IVzGQdfR0Cdw9cASLVvJjmUF
qeV3hKhHNwxv7/dUv8AP51t1H0Dfxc+bFpCEbsg6mqCVW/f7DJ248OXEa5h7oFda
n4Tg8vG/ymPJFRM7alIrkGgYUmrDBZFZ/qU4NWsKgADDZAX1kh3s3NCyUobQMTrj
GfFf9tKwqGz6amV+4OG8M5860JSduiYVG/DdUppoRrgcAzoITmPnIi/5HxrexvXe
Pe0kzArjs4iHLJwWeUlNEuHo1KcUYnOCrduhp0uiz+zDu0M4vwvmWPzeDav/OzUz
nXCasUGOKxXM7NBKroskwXf1z2rJNLaneMRs3UssH1x79DTbvmtanyka/1h/ZRWx
t6fbxnqkV9kkYgV65nM/t3Y90igqMPp+oG9mTNHj7d/lLwgPGAtOhCYiZ5YhFvAc
X97iFeISZ5rgfmbUmEL+pd0IOey7Hn7zV0F7V+nio3MgqOfbiMyhmkU0ugD9rvvb
4u6/PkGDLXy+71nwvdFn12KKnhssps3cl6TsrUiBvXucl2sK1zkjMqu0TubxF+jK
7eTohNuCloeJL5tweVtSmYvnDM5lW37oBppJoaJ5T088WFhrLkqmcW/XeMIzQeR2
dpTQgHkYP3S8MXCQv7H7tLEZSLK7n87x+W4/wN5ogJaCU8pkX4/Y7aP0oaN9E5qh
BVRx/dac200VJ3yi23atoSZ+rwEuHbiAfm3UX7aYwqgzQ5MHd37xOXZvS81sDO7x
6Oi25iR9XctRRUYviHAnYNF04i4msafAgDnCN6c7j9Ohnw2LJVZPiR9NHWrgaxyt
5CMBuWYfoaZO2ykZIS+ZtiNmDXJKiOLJHl2VjYTYPIe+rW6tSD+koRVNiGu5lJcj
00p1l6EfIABprEHtHSJefKlFMPdAbygM3WqDiu1QsLgL1vbZCwyeHFtTJkIc6uGO
kmSIYHAiSZXd1YYzxD7cc3H4Zm0rONsZe+T6jOx8Usa+F/U0jJGeqpK2xsPIiYT+
UEaHPJgLdoqpAkZx3T6cOSizOe3f8pkIRf5GzoR9gVwceq60yG0teQ2sjXhj5jUl
V1a8EM82V1A55ZUyu8r572L77e5lZYwKsyUPupVQaA2vSstlW58l1AtQCaM3y+l4
FKEqmsRlpNJYbkNh81ooF1HTJgPDzngWPTpdYpWdwfoDMGZVW1mpz98CteYlpC05
EYzxVHE0XDGkv+eycw+quc/PGxlS/5aWjB+aV2YffpRPiVm7csLgNZ8RNBtmcygQ
XiuKsO7VoT19pGucAI19uYy8kPVAy/7fijpvlse2ZuaJisx2vn42gQ4pzMErd1Ot
IW7eCVX8WuL6v8pRWObnmKXR0+5hkPsI0niGYMXfbApZ53IZe+570ijoYaTQ0irf
ae9oTMT5pf36zB/wXUK+aE4g1xnOMdo/JOWwOWbiifZgNnDSQpVxEOfBfcDrjJCN
kcmjRvPFhtyToR89k7PzQeKEI1Sx/22X4NkMnxHSxsurOMqBqJt1iWJ/202UHRbD
4aP0CHXeAwfBpA96kxS6K+uc8pS7OlNcCPqacDcppsNfYw8Nq9+ZhF7luMXmOeEz
Ap3av8guG0U4khmZFa1MjmBMGKKEx0oifNoMnqNRTbNZ9NJh3HjPAkUFmXaODP/A
J5LLQlML88FOL6C4GC0L/GSSEJrTft0Mu8N/eV7+YSfGA4IiU9NRKnps5UO3q+wF
FDvF17/oS3wkJcC0kHMcY7CAHlJCVejpUjEg752W7cCCrL9+Wd9L3rm82/F7iiql
3jN6nwPDuEJxJnzwNyINb5OghcZA6z8Yag5H2E5b3Bu5kJPE9jItu0Hz5FJPlNg6
H5Q7LOTvYTkudqMiBVcnC2KKlvBeKes9iJfXBzFktdt2ba6RZ2uuv5qpViVQSs+Q
u7KYzdVj/3vHHqXcD/3DNErn/2Kn9b/WfHkdBvz3M1ZAtonGWzKzOxOSySb2Zx3H
ZADruc7haXcCaZx1cmnE5PDojN847XYx1vCvnsViMiBIaO7fS38/PCng47VvRKkP
duABAPn0DEXB6mj0etq1k9D2gzveo6sMurtmKJ9jpHHxFF2BoXGuKxlGQpMu7L5i
B25PKC3LNgbeWHsa8+ED7ZhVHXfQ95oOlM37CQiJ/zUgWQS0DgTXx3lW1kGb+0np
7nvw+/d3MkfR2MghEDncy+kYq3+MUDBPybAmNVsSmqu7owlk/cudrsJW/5h0H+ox
hyyTKrQ87dywy5KBGYAirXqqcyUG34vt0WMZP5kzaZMEDwCVK9LC3nCZZ9BB+0sA
TLrJwnjGc/FOCCklwYuJIM4r4V+z1i7MnuaPBt2zb5WRlBK8Pq02iVTZd2/UqWkn
gxye50xJGGRINsVrOw6KkFIoinsQnZHljxUY6PV3QkwJgzOcmrwNySeXRhmSeuXC
uudlMw9DSBn+K9KF27oL0ifTY3EC74qVwitSEmSx2z5u+cFheUtPHjdcoZs0keAx
CU3sGN0IxMDEvzzTyY3TXqeUxwfQAPQl/bY8wGLiNv/ACsnaWkLW+qlxSQ6GrJKx
sXGmOcNOZh6K5VFYL/0q771AqUw/4gMbUwAalwRjFRbDnYLaiM73FwnMyfUuPPsx
fquQkW2nsTWrf8QP8HjVS3h2uVPyBfTUd+7crzt9wTKHGUtFuv6PaZiWuycal0V6
FyzX1tHSD3fIGToMjWKj6DLhxxeBI2nYZi/VMx+6dRCTMoYSxrEsLidRQujKayze
Tmn87jW1fGEO3hS7tlIZjuVyaSQWFER7uCMT73nMfsUQpf8+aS7f2aDmHO6gELya
ZUnO1jVCoL4WW4cinYm2rigwwZcKQgeoYeXJsXAcAYrhQH29LsxYh2hW2x4x1h29
0mSxzb24p92WakuLULl5DgJf34GHk+LssDVOdKjyMAdvOkutXYLG2AEJC85ag9p7
ZPEoCYMn2m+Qdlfg7Ec4twdbIyVMvZ2C0BatuQ5+bbuXPU9JhMOsNTcTCJwLqevH
zWXJ9yzrzHxWewEmkBJN/oRrLWAhr7saGEIs6JUXXz4e54jbturSR7LjpsC92q25
8KpfzOnV3GcUcjiF84dxtzk9o+njSdaUs2XpiuHkBdPTKhw1Ti3gi51sZ7IZE3mf
oOyimyqCMLfOQCGUutG58qbqYkg1yPckkLmxhnuFvEuo3Xy4Xu/Xz5wcofirLiqV
8JPGEusD/LICve0xh0km69fXuPFHVh74Kwy7e4HEmGnxQrko5O0KlhGfkVOZ3KZT
e5xFmBxPCTrmBZDWxKvayksTchRJZXF1aJ/N/q4kY8N/s1QdARW+TJXu4Lt3gJZN
rQNfo1ZBYb/R7WS6EPlqAh2ufw0TFiTK6jaXPHJSB5aIoWSQfHvN7TdLMQdhAgIb
t57f2ucu910j5gJ8dr12NqGEd4meIwKyY7y9RwpvfSmn+CpTbi7jAEnlPEbv19kT
ow9aK9AZLPYXQQGSClhHtWGts11Jjp3lEdQmCNoO/efg/8W1oOVn8S2DScHRetb1
eEm2j8naslMG10jWP/QmGpRoRxrTSG7KbqC1bkYC9a9jXQzQGzeAgBPJwv5YTkUc
Lz10NtXTP7LA545x8eB9hCO/omA6MIircH47RTA+dleh8scum8G1MkgpdsKfQGpk
Rx5lOjZaXnu1/zSwr2n5dvTqx3Su/JNyHg5SL1C5qJ7wRTVlVAhsQfZg+ZKU3r95
PFxciY+fJyfh6ZH+pLuOCPDbPmPqI1n7GZRy2+22Aq2NbXqsIB9oHSDhSiV6wREl
O22vfY5LPVeHFuN4EqjHtNvH8gp+R69IDTTiWHRjIhNlEYFtbJrwAoRjKvaty/WK
B7VjTL/3yqJKbhaHAxJm51ZNMAuqV3B/2f0eK6JxMf8EshfuQ2C7OpoDxWKFVcA6
ChhYMr5oIPb/469ZT57Umt1pQNBhKCM3fRsmODR8pIuv+E7vxhBJ9Fr5Cf6s6w6i
/R6cvI/ffuAZiR/cv0huMAt6f4NvgdeQt6SZC12eYL98FTVGayJKxn6ohF+p3NrM
XBjQrFDgT5iwp1PMcB/gP/SSyICLKMOcKCecUBN2RrppfSAF21hYs0yHLjJN+Qv2
oDAoN3sGLhK5YevxSQRFlDxoYEUIpGzgqBzE5XE0ytX0oAUkiPBem1iO0a0Q0Izn
5dp66Lxj6/Qu81aY4XTy1SV2e5z3fgEp2Z8yPYIM6Lc9seLPB033PHBGbfk622Lb
sVLGrzb8FoAAb2I+wX99j8WK71Iu6RFr4FD0xtX/KGhpA7Cw7HFF7bQB310RxfS6
0PiaSvS6CPpStQfvN2NYTM1vJ+BPFcIUIfJ5XyoyDDfFbE/+2OjaVLU1Kxrk7mr1
pnwHTopBn1LEqeL8hN+2W5MslZ6G5LWyTq/E7uyrxsUHSfuBeYSaCbRgRk5kprNP
T95Up9O7moFvHvsvvngJvT/NgHl8tW0FSV5NqIo5oOsJpckGxYmk8KCBr+dTjcKw
phH04YPJ5hMjbKO3xL8tlVpa3FjVqOs7KwpuaVTOKO5RP8TauIUm6AB1xPSFCytn
k8Jt/G+iec4TZOw+QLzIbejZYlo8OLJEO7UCl1gsTjui72qFCS6ASFwi2QdxB2cm
EaInXfhDtD2XUey+iFQc9hWX+FlS40DvoNlMwYRveemKScMXdHRgxxMdc4oyI87E
ryuzYxpQCcyD3k5BFuFxy32FUn1HpKc+/S1cFA7Mu8Bd8RAkiwo4Dg75/EK48le1
Hbm4Jp5JR5kh3TY/uiHG045wukTLEt0syHbdtMYpbkfF83j49pFyxgRHLwo9xD0k
JWS41PCWQXozoEeT+SCU9fclUqxhc7jpNDjlXM2BuB8x3qgifqedokfKGMcOsmkG
idpwQPbVKJXufQh4TzskUbtwC5AhYMhUUu1g4jAKYuBUwM2NCn3MLj9brWZcnWSh
dbuJtwEbPaRsGs4/r5J/9q49AgRqy9hi8QzftKtQIOBfacml6D3hvpwLWF2vrAYH
ouVGPuHY2Y7gj78rMdR5tfw+E3pj77oxfARBw167KrJe4R38wr51D+HgKzW8O1cY
Prw4me2uwwlAiAGxlQs+ASDgrna0Xlu7GtbpzET/39WsUEElYPJPWCAYyL9hN5K7
cwvJXFlJPzeIMvKlfzfvjO90NN8isCeru/pHlom+2VmRRgqJPdw1ukL6K8YXEMKU
fMAB2dkxbf7luvwQ3KB6Isgm/P58RUjjzaGRDUunagUXpfiWjthH1ODcowW0stKj
fKMyPrRrxP4WE/HpwfWOs3QAsB0gMbxwxsTq9JZ9HqXODIQMCgwog5ZeHgukE36o
xhLs5Pw0j2Y20ldFL3hNUZ80XTFlKHwRajtl3/OfY9ZkXpkQbNA+SS69NqLTlkk5
utKpG9EznWsOkvdlspayINg1Mc00DnR9VBwT/dC51CnRvHgC6KOAEFqOllg8woOM
GDHv8xZlBxfrro7A84XFIwFdLbQ10RwIkwks5tVltqKBXQhFO7aft7tNFTU2GOyv
DcFSjH0zRjwMscZviLkcit/nTXyzguISxDH5RJ01WDWsvXz1zvv7VBu6O7t2RVu2
S++Ew4t17fdNL7dXiLCy7AtN/O3JoRVh5kmUVOuiAfBBl+SZpJGzexz0rbHaWmYI
sYGoiOrMpNrH2owwxJcIgdyBjDfLZedjC+VolMvwADAoh/OYZtt6B1oMnnLdoR3L
p2+yFMgRWme4JIFVRc4n4HAq+5+JPnkb+Pv7xXmQlGbr83LeiIsCYEdEf8fwzu6o
xM6jX5beDs9WUCUoAmhqWgLNYZ6Pbri2wZF4O2YrYBTxVH0Otd/6qMmysJgiknV4
LMPGchoWVyl5oFR1MGOgfyg+XkDwqOd3t7y22DtLyZ5QaIWQzU/fsAammzJzt6qS
rdTcvLmzhxCjsYLfaD+HG7/Xm+jnoiEo0T4+uCSXrYmdz1WWshgH06Q5htJYF07g
oNGjHzWlT10R5EZAWbZIn9GBSejDsAizJotp8HV66h2bilFvvAZzWVW52ngLS4Wu
wyDOn2/1g+Zgw6DBSEteWQFEKi06il27gDnwmEi3vpPXh32rWQz0rD/eWejat2ne
5GzhoFbVIEJRAH6VsZPy97X0bXbn2/1B8QNhCRYff3jWogEiTnIp3mg0UwGL5QQT
Bdtja8SY//HsY6TtugoriHf4o6N3LzYXxkifn2HphmIfqqaWEdgyP5dH5+LP5Kat
61tZ1bRRwmuURxdUnjFU9LaMAXf2W6CqPgs6DGeTZvVjli+GtN/fTYnSjQEgUAtJ
iFw/mxIQSqIzOM92CP0VQ4JMlOQOy+ZWFLZeS1MR/25EEVOez1Mn/FK4/4JcFAHY
7EscHR0ja9H7sbiCIYy+x3NOoP/kNRj+g5ODYBIWiScr/o3zPfsBl4eiuLeFtkNQ
th6lMAVjpuOUZwaeCmlwJqi+5ol/YZLSB8xiGRzDpXMEBRMWZc/G38qSdIR27Mel
B2AP2lmvPWbJ8NieG3rsmUIHekW5ulCZ//UnxTYZI71MKzAtDbMGGLQlSL9SCa3L
SjhIcvBfJcs1IKT8TX5LPkXMvEpGCk0vCmk3C2VzhFZJs7zktBlDSSsNg7AoZoHJ
QjQ3SLVqmlHJ/82OIBchm6OcagNsPQYRO/ZImp2NmrKqzwgVLiDt4/UbeooTMNH6
dZHZTwTlEGK7zxXLEcoL1Mh61PN9EszCxYIw1w5k2lYTAxZhm2Y3BdMRz8TlTA9J
dwm5yUQfs/8WadpR2TzRQRi/eRT0cHbgfq9h0ZkZTxT0ENwhSw4MSWWj/ddWmWOT
NBwyK5ytQ7yVngrgz7mry77kQAStDK0Ivt8LsIQ6397j6JyIbxEwi/sk7xs5a8ay
HfAbMEPxk/rYRVwujeK7JDSL423slTI00oNfsF0zKTb8UjfulQROLDo13YEpqeVl
0Q1FVaRi/lELLs6RU9W6KDcyjkULQ4dBcvzjr5FjWEgZuJqpWHorcO8sRhI4q1td
5ZbxJNIYxEfAqlb4MNICeAODQVF3PzOYVGGCmkTSKhgG5A3PjZHd/dxiuqYt3etD
0CLRXnGtOvWtyX0MgVWjB1dbt87A+3py4K1VMigyhMmDk2pH7D1m1aswf8g2psQG
e7bDHCvROr8T/FPxnOE0Hcb7blwnDDxOl6FxLXLiSkNA/057h1+k3Ee+AlX7NlUL
d7h5lBeYyx/6p7W+R3sJW9Bh2hY8F1YM4RTjo1Jl9m/htvoouMGLwEOB6az5/MgD
i4vSQdmvj9WLgqkG9ZCtuFB6wIRyiVNLLvxKnHZuVwcxsQ+3qOaxnQewiag10Xfd
UN/srV0oH+bqsbw9QKqL6KQK6Pax8UrfVFvAB18DkxtMp9JYCD1jrGnec7ocxA3h
Fl6WfsMIQHvWlzIJK4AewZGsIRnAMa2f1zosJj8B+WHUNT/RZD3yCNJDp9/upeLz
LRDpgvtiyTrxX3VaLl6Idrtk9z6ASCVdsOBxkeGvCq3uIy9TM8XUkVZ4O6mOPoHA
AnHnhyzPV9PvxmEbQLuD0AQyVkMAI4TQ2VLCdRJoyfVBKXgIKU4uWiV0LCZFpPQ4
N8V0uBYXRD0X7UlW+0XtDdR9eV10O1ZppLsPZhortJpaUecdgidACRd2h1p4NW37
G+Fp2IIB6QwayeHvqTi5ND2rVdZWWUXZPsGbY5proZjKiHKfTjTwrQuBI0fGb7V/
lKAKQD0OKGrhXaZ+4d7IQTzjwswJHfP+6hBjmRejeAkwGx7bi8et9e2HUxihEhPD
vF7pTs6khSTm8eGtzie5GT8SJ2jV/gBh/Nq9iCmwfogbeRHFlxlILbI7E/IWyJpT
guoPXgXGb/NNDZZMTL/mnb4r82Xfe0pp6LBYm2O2XTRmC0JA7dLlaJbzZ1rAyGKJ
bua9u2KtCyu1orDmAASZR+QgmjFbmmW6JrNOvI/UB+tPkPS2mouAfUMdPPtHLmnl
LJcQNhonB1NUuhdFY0fV3yb+35bH6f2Cir7wxO29Qa9000M5AvcyWiuykvNitK6q
tMekEmBwSyOKes5apdo7VWG471Fr6DJ5GBEQt/SydbPDUnyD8tvybMwFAohHXTnO
CwOL9NSKJTGa7r56NOrHDt2xDSAH2su/cFZNR/snTNRw0obLU0veZU+dNZZTSEFK
kzsXsCzmVP6RG2mp45DRlJSNM8G0mcncZPouFKHsoEVA/tkLFcvXUvMtC0BKvMNo
8lE7MWKFfVALYVVf8Nw2tO+r3VFoT8eF3EN5jk6nmKLhvjJdBc+/meag9bOuS9zL
gXVUN1poELDmnQX2rgsyYd835iVx8OOBfyibBxKiOtyvmRAEYz3YghhchyEF1seg
+1PtvwPfq7B94spYqVX14ioeZECJnMjJSxTmTIkuuEbb47wOQrTAVWA6ncRnbW6e
klIA2HjpPrjLGS4BsqDoyLAwsABTIfMEhx+3iy9oMSFj1r5xhxBLuYJB7AyHoM35
8+LSo1IZV2zfhGkrcnW52KAz500+OC/jzkFVyBER9ihu0MD1HfOI5uADU0V7da+2
YGdECqatcsT82WPd+6Obj3TcDUAxV/V+MO5GGPvg+7vvaXLvRNZXBn3txXJhTCwI
GUacFpWHnVIWhi8vROm78OMmcrQyq0YBu6wcAQo8FMu74Jxx0QxwHJXuoTPTI9ni
JpCe9ZHgJ+WeHudfG5oGQg+TAzahdr0lDouOjAFoX2B8wxA4uBOznozgDwRZv6I3
ueJsenHEVe9hZgbqCuZvc23KcBJlAfaINH0BpNrloL1hM9LoKbXpXdeM1xFHfT2L
PCdRwMHna7+IXwOErzJKUJn+KrV+j2gRmc8wPXZTT0t+hFTnXOfO/J4iX7P7lOl4
pPI6QFC0kfDInLavzjoeYROq0VoYIUb6ETOFg0JXKu6y2yuZOsUOPGwiGhVssqdO
itdRoJ6Fp3LdebHmNL8Yn4JvPTBiF+Ip5d9i7fuUAqbyXJSspdWE9PDS5LqJY3h0
VVE6aGr5dyq7AAsKcVUpbKOfx1OWQjB49CRIaBlTt5m65pWnZGpd/FV6CYfNk0sI
xP8EkQHslV+6xVrw8OjEN8hik4RZlsTs7QgyqqVMPmbEIqj9s8Phy+Dxaipjh6OU
8AJt2eBW1LcsFYfTLPM2FM54SLAo57YmON5ceeMzFoEVFPOZ5L8hD0Ywbs8x1301
zbX0fXm6OsDUGeuKFnOJqN5Y6YaK1HGmK2X0QeVSyUCIOiRMgmZAggsa+GePvHWO
J9XXuSfBQH6O6TltfHDMQAbNYtI85o9iIa25cs/BvkAQDUqDqklxBO1/VikkTece
O/qA8wMmd+ec6yXYtVN3edxkRRxxv32AgAsbmd8g9HLC7FG0IThwqFJ6kjJDVb+B
pRMGA9m/G34Gu29u/tDhYa1haprKRffF9V5ujdPqKy0NZQhPfaOZE8ijSKd7KtZJ
LJnzaIkyVVtAtGyd91KVd3zN3jVdAS6BR4eCloy2MrKI6sphvrCR3bRMb+N9PPYj
8rraycKvRJ9kP9NUzpmsXu0s2uJH4wGoDSWmdbsQfwJIKMYTWYvsHV7WXSMyjKDJ
x68XRtsc1O8nNcibaHTyQtmJps4f3mzkCnFhinuEbNa61ZEPtN4Qw8XAbkCrOKCh
28SRz0wlwgDRBFDADsXl5FVXpV6aiUWGxr/nwwdedItiGH4O7e2x66u2UkpSd+QY
MjAuNfFcFkY3v38IEuKKl4Qe9TNnzsazcwHUGfkedKJH2wTUqGVJRmCb2n1Iy53E
IlsalzG7o9+2V4r7dJfh6P/zk3GHZgi9/Vsn9fvzJi2S20tSyZ34sOLIXnrWNrz2
JOdpXg+zF1Sv0Yml+xJw4DXDOQ4nhPdzX6DlGVcPjHWfV4tYOBRYHwZa83uIFyGT
A7d/ZsWlB5fxIM61TQJxG7CfryUjIEJl98aQkQvKTA8jcjH1jqvFr55Ubkk0uXTo
pRJhsSxK2D6whT8CItJD1QRjS06GXJNGdDANmcQdu+i3Amq5/b5gmiym7Tbl9e87
KIBKOGcyUV2C998nXzSG+vfXVCYaFmrAKX4Es+v6aoZS/W8iBphqd9aS66tn1uuR
7RsNOvBwtuYKPkFpjp82MZzlBvNSfg4AtDKFLgebz3jrHZtNTY06gApNwDC43sig
da4XJen6mj660ATinMGqAiIdHMrJT2mT7zEuM6nU3UXM9TX1dCroTJ5+2/NaSXuA
KhDG+C/dOrN+rU4f6EuvqRKOh0xQOlOEe18CP7A1ER5XnKQ8GedUoftxb0DonpvV
1NmKfBkKlbRGzyHvBkBhtRX8bDFKQqPN61kJHpwNL51qhpLnYZbVj4A2QvIzvZ9X
wLOQRdX9Z4rbo5b+LgPh/Oo8eR1Dv9EDUa5xRflxwQ+ozyNXfZQpxvJ0aIRJ26pP
nrG5jGaqfjIwTsfDldN56XsC5+1i0zXeUJ4CLjWlsobWfYaMYqah57d4Bqei7qjp
w73eIWoM5o8F/dGE2uNNJ6ef2v9ZiwavmI8J/bX45MjqP1ZPXTwB2+QGREz1FM6w
aNM1D9k7yQ+4RTj53DTMztuQKC7ONfpDstM8V70fQlckj1ooaW5W7zW5nnKAM3kI
3IdPZn99pxg5QsU4k8GCDi078vqiqHQqGHVEfeyhIjsOCkgEWbIKFV8z+CGlo9Jf
GUurqcUGeDK+bwIR6ImvuFPNBiI+uWuC+3RwtHIrRfH+AV48/i9Xl3vz9CZYbG6v
pjk6Y3UaABdZhqfI/8RBiPJX9YwCibD3qKn+mk8jBO8mOOaYFq/0b+hPr7sAmDl1
ERdE30A6GBAhkaifPEkLYl4netZ5PPSJ8DyFu0JYFXD2dOF5vq36Ae12LofFiOJv
NhDoZSq9WYOHTvhGWLRUqd8z1NWaEfNfmPY+1XgaZJnke4mwlLFnFVfAum7zDJcJ
lPBRRCtqOXXfN8xC24CD/PM3XuJCdeVsTvC28c3P1ryw0TiXfyyxrbK9xmBT/ko5
n17HcUVFxIBmYoOxMdMMK1JndPBGbXvGxKZErYwV2mcqSNpWl8+mZUsfLfwcSnqi
Y0n4LqOTi5GFKsRjl3I2KVcpjR7+Vqz1M7IJ5VrQCn+cCOpcuRT9U5qS3jzAOeCi
WO0tUvAkZEkSpjtfXSrvqAx+Rie8YEWO4yQGmhQAeyCVqH6rlR6sMSVEOLaKVSdV
pRjD7Ok6bghl00pp9BMrR5LIkml1bxI3wzUx5asM2mr38GTudDCtV84zdT5+g8de
jTJKV+QfI9j338uk/DhORB0xB6uuvzxTOjHQAdaZdm1SbJNr70U0QjDR8soyNSNJ
lOwUFpEKYBygfrtHMzQ08SC+f9xRfrXWfO0Vl3GMnx9gP1NGW4SC+yIUfLD6jhW4
KFEeg/b1OC68G2R8X94EJVxlD2gLEpibFJF/Ci+0z+EMeiruYTnictUyIERSIDCe
x5AWD8NC5luxBFNvwQKD0vl8gZQGadnd8bZbn7spoN6RLODeQkyttVnajmBx6dMg
y2zLgBy4+nFnQOXBupvXsp3kXqVXXgJi1ru9r/ZHjhELfR2KHv3+49tLcUV7h5Bb
2EWdzCMfzBpDmAgz2WKdHAKnSCqUK3C++ojJYIrMnMe2emfLgZUHZDg65pkzvc3l
viXCcHTNyhZfKBGhlVnTPQCyN6iN3/6JDnozZg2lJ1Y+5PYi141VBTuAWji3VQ7Z
VdlloPncchrfYGGOdf5nKGeTDeAssGGPWScY5I5p1KkAFzTlMXg8ixh2WiQ10Vgm
P4QuzczIlOChf2sccRbqhGIXKY/7OnepKsQjwnNysIeS6XhYYLF0i2LGNaJvrPy3
jXqoW5vIjdMwa1OGR+bcDPjgrKJLUCwMCDtBa5im3uv6PO4pL8boIeEk/OxBUcdW
Jg27vT/CVww9Usboy28Mh6/TrV+uZaKSuM3hBGYDxXwMJKIltbX2x0Q5Shwk11oe
xc7fhygUBpV8O2eKHmHJEB0+gjpOlMLV7YZ+G7W2nELsDD8DTKT/94dgnyYqkOO7
XB5Kvk4LUeEmeK3tBBbPM3MSv6WGfKvRKIV1eAQ9kqdkNdYOoNRFdwSwX/vjfCGX
OkDtcvGvmMLBptskfDtP6wSsFSlnlSet8xfY0/B2OkV4YiW5uJOI+GcdHaicR1Zf
hCJ7KjHKZu8X3IdihfgYV5tEVhJdRS8+zpF7dlb2b+0h9R6SSAnr0Qe4eLCH8gRt
kExH9JmQC4UDOZCUPYXODUdyBnoWOgj9Ze/A317v8FEfnEVtCIa4wYC9QURf34fO
ofJ+UYQjQ4Jf9nGG+ByKN5Jm2xdvbMZRy0260G5nYMxiJcwD9tSGvw2Gulieyioc
8JYbSfascn8ur3X3q8lxdH2+EwuOlIWBk1EGKOxlMV8/GRiZH8Q7UmCZyMsOP4tU
GSBE7Zugbf5jxg2couyMlTSv6d6/UFOd7X+83ZmsV2yQZkB32dwuuQwkKcSAncRm
BiIj3eVUASkRCEG93ZuIRkluJblJGnPaQhJKqIFSuQ4xHNu77tc2rntEHaZmqepF
IqyLYCXOIlaeBPuLAmxcT8+rgnLoziZTGoMojkw+EvIpfVkvHMX+a7eQyyaFwlCd
07LB8mHae2Iz9j6WphRc6OcsmV5iR+9BHeWon3dnJns1h7LisrepBahMacC3e+xg
D3nIzChr/Vu4HHTahhGf0tCVAa+u7c2MKdz9sV7lw6fqJHgQx3KXXJ7RIKAXzR8z
qVw1d4s5taIBPzSMOfIE6JpP9/MbO2tGidP+herTam1owY8R8o4cFncpreakMWy8
CZyF2G1D4FjtV1+58fBD+kkbJuR9UKFjFvMhoGFKKdaxEHvTV+GMtdP9DY5/2Ah/
sNk/r/pMobFEHrNsubqVSQoAYz+cPIUw40y4NvM/eGsuUQw6NjjPyzVlXJAM7hkh
sYIVRZaI2LwHNP6XqmTTpaxTKPETOexJmLyZLguIPwQ2SO+gXeVdweBmMM1V74Dz
5zB/BNI8RPHGQRp9gM2Rw0t20M20uoEYdzpR+qedEs7VJQ9MECO1JQ5drYStqreP
X+053uG8o+BgxLTOivsWKQjAF82171lUeilH6idSwq54kzghHU7PIM71eQEqKgG9
VIytxxkFuX3AlEG+9/Irtc3Kb4k3/3GAD2G+xmmm121zavd1gxxfK4FYQMkjjGcr
YdzkN5GMYuXcf5cccDWMAb3Pn+fzRma/PN61WECr2A5ppJd3gf3dw7GMhfVArOge
2ydEXea97iiWMocN2dxwyVkFzkCI72kefKdrWyc8VosYemJpuP9K8htIx+DjTCuH
KfL+LA59cMZ1owBFYcu3l88yVOZTlERxAK5qjYcctVXFoMz5T9bDD9qsD7CAdXsh
Mo5Pnm6NYTm47uGgp12EB9f56aHrXuevGZXdeWD1KOlsemuy6I0vM80clwG/NtaV
bgJLBKmCblyPyDlafh3mHQGRYbm/MRQlqH+IZwTkoXop5fGqupVT2zi74diAByBF
Lg6UxU2fqu9RTM1V8QF8VsmPnSEPoRxMDMZCd9A0uSkax/82fuflFCfn5IbdQ+Pz
yJ5FXYv0ANzDTIzNY3LHFSZ0Z7bsoAy0W62Ec0wKlOW9Lp8OWmaWsOdINNOB5dOr
BGs+ou3IfphrEgtKqLqJxQ0TaYR6T1Age8mToW0iFkE5zd04zgG6g84ORkKDoj28
3ZKetm9C1pL62b/kOcTtEMtptYP5UZoHGEON/34jomSOyLZTNTc03dzPZKAc8UKO
df9Q2LsojFyP0nAZGY67samVF7Xt75socDQC842AKiM19Dliv5W7BLBKP3MJclCI
M2U7KiuoNy7s6ECLi+lMVaXWH6AcbldKxOFVtRUsqnrLLILwhbp/lY7vitUhHXpQ
pMMnMVThedKAyB6CSF7dLNXvuZkBSMXcofYXx67y2BhSNWWx+hegreIjcn0NGJ7y
/EEq7XkhU58cmLLNTMZ4cOx0koJzm1ofgrv4kaGnYdHK0pI84Bm49Z5KrJmPYEhr
u5rGfSiqAUGQKESZb26/Saf7Z/XSzf389/WGh4xWfXuCvLM6jK9Zs1IoIQuhAicB
EuD9unTAbWkH84qmoXFlhVSF8RvK42udC9n+7a9YJUInzKMzEzHvlyJEm20AkExu
iWQhr4qit8v3u+GNUnDM2SrcrL1tAHAcw13ttymVo5ouMToUUOCEFTeQLXYDfGyj
Yza1KmDIvfPA4kdGwRnSBuTwjKqz2qgAUGQ4Rp27oH2iUNyZVo6XeqvF1HYtBeUN
seB5UQ/JkDjj88tc5rezmae4NG7Aza3TomEsqCmn5LZ8h3UQCfz2wkUpbrwTXqE1
E7oyLhlap6FE3sY62VLAwGSMienIU965c4tqsA4rQWOdsSUD4LweNJ3jRzrL5Ra4
guUKcOr4v3ohwCibcgntIThOADkpaUQ6fZwpnUzIq+TJlGEQjaqTi73YxjOVaWcH
rQIYz4AJB42kfegG5zaejXn972SREeSJ8ohVWzErAPbxCQiXhSLonVqqUoS48rHl
TV6Raw2eMg8H+dpHmhSjTeQk2x7NamhFo35gPOl9fNAxmO/KNdCK1wGh6D1unP5X
GpqbtMrD4HNzc2N+67HDHx9RDE5TW00Z0P92oJIHh4MBLHs35nLfrQEvNSuRcNkJ
hPO3dXM+ZLVFqtnL0P9XXx8B8kRFs2OROzTPE3dUooqZcBrFsJQ4UiFherSl/nr7
RzPrTFldhuR7dlwA2RbOzYXM72eLiITVoV7eCjRLKgfJuwB9EElLvBTFcOYlkkaV
5ZQMq79snDlYmDY/oOe+SR0d/K7mkNVFR86uczcsA7N+ssVBrX98H+GLi1N7Rx76
pV21k8JsGVnyfEFk1xg+xwaRbjqTptiScdhE0M2THvkZWyFQUyQHUV78W23ch6sy
c+qHVR7QPrveT/MqI2x5bmGFoMCn28UfJcnRNQ0Ea5OxZRjX/mBa6CjRz3BtzlN/
/p87NA/uC3gMnUzNJOvytJHEF2GtpjCkvHgQ5GhIol12RrFPfEcZjZJEy4eJyNmB
Ds4X6HfNH4ap1qWVKhpav1WvEGSz3XZeOL37XDeFt+XUM9Zz+/VdCfEE9b2AyWf6
tamg4pHxzTUGP2pczBT5lQfFCxtYdEvUYEoDyf8Z7vdmrltW29p3TW7JzRX8H1Wc
9HHq+Qm2POK/EgjhQTIwM433T1HvwuRpMM2aI2DznWmrTdjJYZhRtB8SeBsl1+qK
vMo3TPg3WbqVxFCH8G5RepbavRY4IVcy+w1O//U793DzGb0cI2+wP1rBCtmG7jvx
aUim7zIwK2Tg/rytA/P5Ko2uZgV1bJY94KrySStFLamcZWqeU4P3pho710xc9aLO
m4knGoXjMy5fPB4EYQh+cwJAyhEiSgM/ojrEzXiARK8D5p7+ZNTeHhUbIcKO8nCC
8o0Cu169pRqu41kfIkUYlyXz0xt34HGQnXLb70ttxU4YzGhZnajm8msitZj/yb43
WnJZsPxH2AJy4Gu7CFqy+1xbwjtkoGHeq4cVzN297ziX5bJqhD1KpFRtL0KGyAjk
1IIRqd6ipoDyt7JxWp6ysT2dC2olnVq0G/x4GKuydAZYQRyfHXPA5uY3aF7F3LC4
Uxusy8A3uI5PC7geKqp81qV2OV8a7UvrmyyWWv4Pht93bJ+btdREOBCzZtvb7zNr
Ii41uIxSUDGcB/yTulRFL3fpCSThSJnroGF3HcjvxuQysyNutq4QDkl2f73mvi5m
6o0AWtraPEWRS8qI6/Pi5YTodEIqnUwYMvQmrlN686jiCJNnex7tyi/+/i6yX/lz
BmmXElaVIxQU+J+BPj6S9nUR572UYbZLMI9cMCxSUJBL9UgDia9dS9MF1bKSccW6
EGSEsIIhoQ+HX4c+plKrHH+c/7Z2YAIrEQtlxdi05b8HdpqvAWJiJ/o5UMzNx0jX
zDRyRfB/71KJtU2L/v0cTFhitHlxi8dZat74x2O0meQAbUrvQiYs9box5w5G7SyM
HbG2kKaGtkwkf0YNkdFhKD7lcxpvR53hI++y5Lmeu41lUbcy64gWnx7N+tj3UHlJ
p+G+1I5xtAf6g4UR1ZF6amiJHCG5RX7qA15jKeldY9eNkS+Z5YZZWJLg747fnrMy
xCICwYtVFgdvt+bGHsZofsGaUyXjDzcyqMm5eaErs9p+J1RpSObalhe3Z7MNUrih
FHuTp+6OzujdTXgB3SVDIDxrIHhuOOmmgTCImtpxMWNzQpagM72hbM5AxfG04oPx
9mGcuHf7oZA0dD4MtLkhL3005CXVZpw+lv/1GjjUetq9WN721tN7cM0uFWtvKMa1
qqWRgi/LK03qdOPeZ++k7zbzzpuegbmzQVN3oMPIPgjQqpG6EvXAbbOnO5MppZDP
E0ibdk5ZTUxtvEuLB25gOcgnQg3HKQphrjjpknyQgA3ChdwkWC1SZYOZoI1McxC9
ejzAI5BOTjThkuKMTXbMMGNeeufABgaT15ANgBoxYCAETvcuOzI5vUBHNHh4RioZ
w1Qo1vvvXZSaVkvevTMM5CmaUTnwVPzf8Aeie5h92wl3OU27trA8yA2t9RZBqkSW
9LYjG9Y+KB4yBL0GX/lcYnuB1fsuOcrPWUIxrRXFbC/xoi1JZsoJUuRHN+73KFte
jk8QAd2cIrdb7+tzQu27yZSLx4LE3DNMPQUV7+7vWj0jG3sYKwq9HcYFb0+5e2v9
jz4Yeae+iXcJGaVuXE0c29r8naUua3fA/63GxvtVPCeZEDNm3esgfI8oTb+HNPGR
6RC1GvcuamPPabFZQMWclacvcUyNFhnwuitF6xKsAYVzki9NeCCAXKnwh2rvQtIH
C7ltX2kOLUj2BEHrhuwHir730V+z8Z0S3sXC6QRuJn5l4FEVb61Gu5rFct4rotZ4
1EA3/xXPsIrlvnkz+1czwPhKMALzFYcGxvGKJ1T4ag4WlZ4vfEzRdcRY10fXDAE0
M2X3flDRuwU+40gVpu2WGU6KDjDGNluMHsic/NXRqbi90/Vh+ECRh53SlrT+pT0R
yDEXJVLaOxtF76ycD9ajNH9v6TqpU2WVoWQ8p77Io8Yru4o7SYSCfKbmBdpw7Vyb
jzeK2Qnur/i6GPja2/oI17MggV+IMb2ZVOTDead2o2WYrT397JKmHBV51FtI0yLA
YQOxFcaHRF7ieJfHp0wwEeJDVJqx0UoDsHZF11Y7ypYwLA6rrTbQtEYuCNB/I6Jp
MtDdhOm8wZKN8Sx3vTLeEIdmKIUVrDLqK9t5rOuxLXCVBwMJhDmWNgLNBlcnXfaE
5BlduQih5Ngg1IUGM28IlPGDhzZj0lbsC1bKkNHM33hxgavFH4Vgul7EUZ/nF8+y
GqguN66LTRIGtOGfuZ5eGYci9gFBReoWkXERR21+t3w84uMHgpSz6/FVZSBwQZr5
lwg+lye8SvUTYKZKRf+wDlgaQZkrfmvV8jWIqO3rSxzllHwVwNtU/vxO9kTZ8dLJ
kN5h6r5WnKAt8mnVs6j5+0KHlVWNFtr+RK/5iZL1yamyzdzJvP2ccyehrzbpfhZz
ELtRkqIzEtGXkxZ5uMIWOh3J11urpCmmcMTMjUojFQE1qNtNFFPTEWfNsWMhc0/Y
WXiD1vMOZYAuF0jLqnI7PRmbW5uCaaI8b234VrAeXl4btuO8CnPzm9W3NgjFFwZ3
Iq1MGA/ARgArA7xCfcCB+j7eRdAMa49h+7EwPrABGcGuiopuE3IORgMy/XJbfInK
PLa1D6bFYpf5FT15hd3FNl43IUK9PA9CcCPZVYS2assnARIHntNjkIfLQeCE/6sU
JINVcD7I4cTo6K8MQIlji4TtUdozXaQpEpntLfmr1PLshomlIWAnNOVW3aUnebjD
fKumtbN4y3xLKC1ibLCpr2k6TVmC5VAIMNx7MiZrYzEXL5y8QFV0/fqnNk0byx5s
Pyc5MRB+C4aCXUlQZsfKa0S7ZRt9LN92kIzKHSs1Wu2ewqqZ5Jb6ilZNe8Qx1hK4
Y17GO1CiCVaKBBmzPwZ/ePEnTAXMkL3/WJ6697jBd+boVDUR2MA6mOKZzvmRhvLe
4pxrrb54SBK7Wv+FNZDHUvpIK4UG/IjyAmbjEFcRFHVWfBMkTB+uL4Db2KsQS/SW
0bJx68sayuQTfIwuojry9pt+L7R5+UEaq1D6VO3J8xDW/Oi65GuFzunYRYBB5OiV
n+c5DW30exEHX6FA8OnUZJKkitEVNkhsWaNNeWpJd7iUL8NcbFLgmAep7npTF1GO
RDEu2DM6WKk5vgJ9imkd379zEXXBg966w2jb4gArCg5DerKOKbENC4GZwnWAhD5l
9gKikM3A3oZK8vXJYPKhTfZczxhtffsgwk/qco7DLK6SQqRBtUeGcDGS6VZYktza
E8bNz9pEAgUkVDa/sC7OLLolFYHqAMaeFpmLxeYF89fZuEfsQSm8o6gqQpODe7X5
kzK892uq8pB709rQbWmIZKMChvrKo/XGi6Fj7dZ8TUttJscx8mefMFz/+pke4aPv
z3E9wGXuwEO+fIFYHqzdoew9q5cKhhcTSArRSZVELJ15mds3ypRnBFk6f7tcqAjG
3+yDWynKwLW0T2vBA9yjy2DTFHGrvj7WuOjqyf6TNuTyi5FTQdkl9PDC4XOulr6V
B5CGqNPYB/HW55WEL2w42NpB3FjM0rlvIw9fOaatLCa0yJHacpN18gYXKM2SJc11
tn1pXWy6UAIv04bc1t+bT2/Z99BvhXpmKvCis8l9pxjhoFPLP+CdsIqgtYZpfZFa
0gOLo9pxDrjgzKYI8JI3sAms0sI/sYwsoIr7GqDpl+Ypo8DItON46X5xbxsRebh+
vcfuClWaeeZlNqVi7SjhWg2glSR6R2kzL8L5boO1GBjqswf/8j6663ck9UdB13kV
MZChjlZaOtC92jKs56Fm4BJ7ehpQbGvR8oz997HEYGDw2Bj3EM0pFGk2xc42et9a
qv8riFNZ69kmA9HvnFTTScaTHjMYI3iywTMKZg+tG2LQL732x1wpfQR8dW082uZP
aDUQ3BzzfpemIFzCWnval/W9uk9poG2YuWG/PhnweIklHdrSG3v3qbolVw/qALpE
jm4ePX9JqiZxTPlNQh+QaOgjCklSzNIyW/9Dx8KJi9vnmqxwB5jLUDdembyU2YUz
JPJ7yatnFZqtAcV192ZoA9xhh7I+Kx9SXJegbbv/KQNhZyPS7sY8RS5Ic0edQ5Hz
rNLCla6MsR7zsvbtvi5fEYJSYakvUh1eT78YecmWwiP4td1KKAz9kCDbGOu1eOF9
4mGH3FufrJWpMBFJHcfxZb4WfcETdHHTTJmmt7k8cpvNnHSVVZ8YWoLHKcXaG1Xg
iMUDc8YLg2kjwQSmfsPDvElvBHrdnjcnWkdqo7jsLAdOttklWZd/Dko8PkIYIx4S
QbC3Cs5RvsG+BBBffrf4yIWZtZz1hS3Ym+8XzuFqgLs/V/HOM0E3srU60yHe9qCk
9ycS2ezgT7X8wBbMdaCcHXzyXlEeOmLxe0CoZKhHVAzTFFIFn96GsbLBmqDhvEst
ZWquDF2q3cw1WCzyzDjt0yjV1Mfm5xzmMH1Ri1xo6FUBXAT3MYnaai+4h579/zQh
stbAo5gl4RNE3QdLgxlSp8EyQvsXikXivc9uLvFYqcXCtDFXrnslWZkWvwT0xLHT
NeMGUM9nG4dr8mVKJpuXvK5/57UZmUwbSjB6oouA5AnP+uyQ/3HD9W7SPL+vUTFl
gpCpyL9qYCoOjVntraWOAd2dWJlBz9ID8oW2Tm+VXYVmi0ayIQ3fqjmbui/TqHMZ
3DSB4xRRthneBZZZkXe++wKIZtfBw+pRcgVX5JVYhSClJPTaGGifGi95beuTS+aR
LLKbn2ZJ+Rdj/2mqSXCaq+43DWGlB2jeADiTaTVM1FrnrFj5ypjOzSq6yuu8R9fA
NB34Mhn34xj+2jIjJxnSXfW744sXFTq4bumgp87D8SWEjEKXWEd27gQDHRE6X05F
ka1EaCAqyBVrRzB56dOhbHa1ZMFCB43SvozAplOQ7I6ECSVcgZalHFd0mBkRyjlB
S2joXewHBNwWtK1IX2Rbv/REHc2vZ+mPRy7SCjDc0ziL2RZQbfHYg5U0+FixH27i
TwwTiRytc90TAmVbn32PlTpiyICCLuHsX6dK3IOQzS7yiwRB21GLl2p8+wptuHDC
xY5Dtsj4gWoF5q4/wAc5rynt5s7MXUD7sfDXnMNIR/ZICqV3nT8lX6ye60lKoDIj
ODa8HODHS7semGYZ1Ncr0WoVYwwhnqdfzKte1YJ4XEXc2jdnDn1ChmtVJf+vsDH4
LCqitm84PYy3r/aI4H49YPBwE3PPFFmU22uIP3bOXRPPqhkhsOvBtPoPiyAPn53Y
8fxW1uo20BiZAGRPjcB/COo/3tXLFnav+t0miRV2KaQXQrytr8uUozclPZT91bdh
O+HYG8SL8IvrwyU6kcAmp09ZBEZoZKi8+Or7vOgdrFLkv4wDdGYCwYIh6xVPtg9d
qMMXAGWbk1WWFKKpwYDxj8kXJhl5w5Kpn2dWhDPUvJoFqOukS16wHRR/WCFgJJtY
DEUWpLMgwOJT9jXFwgOMan+kLRcaTQG/7SF5b5QMIQd1pjO320xYn54K3ViXr7xG
QRq5Hsii9WgG6aJOrX4p+VCGwjubdB+UAD9D8vA2R4rAkOlxe1Lfx7rgRquL1suP
DnSPbVQ66O8qAJHdje4RW1FM7VYzabcwPyrYuovX4l6dW7QPk2rzpjmqDmGBgS3Q
TqwjRwZZbedxlx/wE2Ryx0gDdjRCHENBMHziejtlCPOnTVlBsoIMXpW3eS070EHJ
muMM2QDiVCNgwHi7KQ3UvpHtKKzoLS7/3UzQ/EFRRHWcXD8VObGtjqCJLPzaCXbr
+1HebnFNvnSUeY7z0Pevq/FJpgEnyD3TyEffjr+OpiNtwItpwfARxsrVyQD80ty/
Mk4no3KQQ4Fx7LnPXQFwEhPSu1CenWU3HWwzBeQQEvYOYf0y3zYCWnPqt6E4JICG
w22sz8rxnFB/MGaUJT72XaOihLoNE/HVtsHLWp2+OZH+qclymICf1IceeO7B8r3F
pdRBVT0QXnqQ7fbqsodsJMRYn5/DAUl6moqUWrnq3EBV78YmgjDzH+w8KhpD/20O
QAbL+MqpUsnW/bzKMMF4Zhhi+8MjkAGiKeei9SxlwfjQx8RhiAQCuLPgtPFnTuw6
wiyk5u/asP7A7CqBYPitW7ZIC5GzzZIq9w+pAITHTLtuVp4oCucy7juMAHCJ3hZG
n6Zbc5RgWslQtIz2sBzbOHRa90nAfEOpoaWchXtPmB7Zmy29bIjkLc1CT9rRVBJR
9UJzvms5UmfFwer3GDqSaNkorpyCR5JNojTwalYwvoDED/kwIJtHlKVP3ZtmRFqv
WqSm5QoGHv6bvewlVmiWOFgFrUkfvxNxFqyT4dY0a0ZULSkRYw+Dx2E4SmNmPGzN
J/DRwczltPozfoP4aD5388dCYUgKNUUDF9bE8Jb5s4xiULjIGtETqqkO/goy4BSg
43v5894sU4XLJAhjxobR6VEzVbNgcayJH+dDFjHvql0J6sidVdIi3E+q1gOwtehR
uJM8+GHhAPqiKa5vYGiZ23ePS9+YgetzQMd4vT673bgJnZtUiUCYhpK9apMBQIy/
tiyyZiOsuzAa/PNBamXKmtYSz01QlaUhwyPR8tmB3qKfyvOV6Kwm5YZCXxIGSC+T
fOtpfPnJeyNJiN+VnWgpPr7+TNrgbv24TaoH1UNCumFw8BwumRylWa1f/RNPm7fq
aV3FyShJo//cN+UdMdhW12z+bqoIKR5PGKk0cFUGbp3PcMihqYqrXeQMyrYoQLSw
kagIqXMtQcB735dFVM1m1X1CVdnHcTGSmQE4gMSLfOEfw+zMgPQme03Lh7jCjej+
7UcDOsnTnugHn3Ra3KuWB0jCWQRfPsquWBOKSAv3PJ+iSyH4Hq4XdgJbx82K5bXN
3B7vg+oQbvxXXiqOsGxq9+baWbv1N6zrK8m9af0Ew7Kx2XzKgS09QvZxKgb7s2zq
FqjI/jcI0421cEr9ZhqKj6pjrSOyKNQi/qsomM2947s3oB2XFIlNbuaO5kSlaovm
eN6j6ynqgzPQzPbc+T0/snmwP2uEc24YlEpeW2nCLChlRmYe/zCdtwSaIlQE5HUy
V0hoBZCxsw7gmTTsmVwrdVQTBxFnJtFCrndcRnv2I9suEoweNWCuLXeuWLJD6SLb
0CHG2feaAlQqfLYYJK13TAm1rUUCXM8dg97T9cEX62PANgeSoFtfBWssuw09Eqgf
IAsNUKybTWIOOsQN4GJeAg7NzYqELuRzMyQ7nqbgG7v3EWKCNry/NHEHM7S5Mwua
DEMy8xqwrhMEB/RRWMcGlH1vas3rEZX/VREwQOnd2L8s6tg5QB7X+5+eAYp8t6Ra
dIFx119m4ztIxMNwNUs/79TnXrmWD0jAPxJjKygjf+ojwcTrxd6fUcKDuhpd7chj
SZK7Ig34OlFvkYfw0Vq0RPVHzBOaM+dJTEs1Pqe3vNAjcCmOL7pAJV+1+EE+y9KU
ATKE32OsTz8zancqoq4U8ELuguKQx3dFBH4MDif2NVYCquI50L3EKiGdnjtHvl6v
rxFHe1/abVt6wxFMZ73FHDiP8NWV6FmMF4aJmCiZdd8m2U2Bw/yM7ox0mT2E1s8I
gprt+UD/I7Mclix0q+Kk5YC0IWoli4y1A/qyyZrF0zdPI6cPpnGqDaUSz7B1/uiZ
6WROWpufqDZOrcq8NoEO36h/Oxzuys0plxaT4uUWa9DEzQ4MJB5aoWE2JLRLl2i0
BpMAEKkQ1uyQg1gBQKtsxVNSsJsR33xphHOjKcuOa2RYRA8CQEEMbW/ULSS2VupJ
yQA43B+yqKk0ZgDGBGPQ2nS9Jb543jYq8lyTHfR4dHvs2xy8bBE9UZD3Wf3oC39a
QFrygyIIERBgMHHtLsNS1TTNBXZ1BmbUFtmMOmK5zgR1vmohTl59TJYwq9M7hyCn
hTHcb0GFioKzmpE/jcpx9et4vLa14PlVVxrnUeRhJ1ysJoD1U34aVahkWu2pkO9v
I5BEIce0N2PkrlQHhG3bsMmQ+ABUWF+q5ILj3FIeeIQ4rD9wEtnT9qUS1d6BDedE
1KG9BeTxwzkU6ycHS5D1061y+NsrmqzRFlddGrpNZ7STgoyCgwDL4oW+OApAqUV/
u1taR+izYccxO/bhSREHVDx8PWJBmZ/Xkn0RDQSbbFsJtO0/ENql+X4fnnP5fMLF
mVsvC4pcMhIAShFQU4YWEulrmpUfs0AuTjAkI3Bowrj5wPEHt0H4jaOoUMpM8gqP
AslAbqiryh4/FPoM+mXpzEffY41IFs+34Fvef0SZP1wk8l7FXglqzo4NmrGSwqn8
NX91z3HutKbCGadxj8Kuujx/JGqj+1sW4YiXH00+ZsAtCBvW3FLT0u+yvqDBwIYo
4J0TLqpzA5n41HbsKM2FCb/jyXNPqxP5/7twrbcJl2uskB0XV+omhkDj+uPUfx0o
w3ltCMPsSXifLfR76mC2eMSDZkqU5DXHnoBsVfhbneaQx6ZLWFiyJqYVhsEtIzrD
+lAOxEaJvJ5qkfYsDNpiuxRhY2PEvxTHZkM0JXgUhGGG5ZOD9e4xKEHg6clyU1Aa
P8/0oZnF24vtYixRjfrBeAD9srXFK6wpsGgaG3iR0geBghRRI0ee5b3ls9m5w3Gm
YnWHFRoylu6YcE1XFzcgytbLNWhCdk5MD/srqB0BTehwzVy0nlHtPZLY905he+Y1
+V9D1W1JbJzvCx09ofQNAxGs7cJqzwnUfg1U4Lkk57Ik6dcqA7nt3gT3eIUTpGTE
dEZB1regFn+MKLK17f6mCrV7U6+V++gW6Z9lD49SeH8embhoYc+SBc2W8TVcBj+l
oTPCPYXalpp/HQ7YDOPZ8h/Jv2lGI1RdXD9YoXBq1I8S8DvNXMg0XWoOTnOhuuIB
L3V+ZFJ9Yknr04ewb5+9Ij1clpVkqjUtseaVKhmGguLvlcLx/u+aZR4AA9DiBcsH
WSmSO5btWJZmmwF3z80QN1KNfT00v71qY+3DMr04WyEcSnOHtFZm9j5GvTwA8Xzs
KOkd5ZZyjYc+cyIjcDBID3c80Z6duzhwOcpmrIsNVtAoPMSB6YkV++NbeAxQL1Os
FRF/vFGGXNofrZKIVnPwPjB5Szou7JVZQWtgB0tASTxVgoFV1FkR/WHJB27MLOoy
M3wWhbS13crlog0lytzgVBWpD8IG+tsz9I/AIwYkNE7BkAvdHthSlCa7jlHLj9zB
vUE3IHeOmnOxXONHJKvy2apzeHmty4kpu1uULTMF0VbuqkvNP0C2bfixV4ARU3te
GzChvWIPbI0TJTu4Impvaf80FUo7rN0C50qlZLZB5gbplvoftRSM2zQftyzD+sly
IWZY/DxqMuhY8Mc822iJaE58lVI5ipfOxpYPIXDKb9bypCjYKS5D/BuiQELzg4vh
J4a7UpIl7HH94mrb9pKhFtwcsFcp3Rp/TUmHK25UDCHUCXvo53okBh6hYG5+HYZd
pRMPLxoVVOKK5cDFD2TpIiYZWT/qRcjj7+DF9SyM4Kc8YVvNqjugkgFs0BPKuMBN
+xEjkF72EPTWNIHBpCMh4romGS7WTAXLrtWmhrEea4m+0rYvJQu44hZlNHJe5L3D
XlzNjP4SfgV3iwjwIi+M072uOSzMPwgMqGVwn2iYbUxO7+GCWXh81CA1fxEe6n6A
xK4gLtrOhB73xlRmKndTznApXfLiDOD/3kFpH15IOgYTL6YLeyo3sqkgEE1PcnSs
9J7hGTAwcaO54N4DH3pEErJae1D2xJlT+nuUYt5/WKMpKufRGbW2OQe+NP1phlRs
A/iV7srm356ecEwvUJnxts0O+CVKFBytU9LXJAmiOVtAD7Pm+ffwvD4H7nX/PHHR
G+1pYs/+/HBZboAJaH4ldyEVF5gjg+oUijgj5+iyTt30ABCiEET91bIn/RuCuYlw
FOjH6u5T97/EV9qa8LuWS5tgUIhrmdVCnxLfbTvKK1Qbp0p0+yrqtNPAW7XnNb9N
OMnqmMLewsFp68QYK2Nxh9SmK/uhqhDheQ+GcmR44lGdJrSWPkRBcs2kNV2j3ZWH
a0s+LYVDukTBJJaoGurtMlcsAeRJylJUUH66IT1BtscGMbjWSE4OxVvxzj/DH9QU
ahGBkzu3N+QoSp+QuOzsCD7wIGrimItL3ofO3W6N1WbDSpvSJnmaiuS/JJiercrW
9za7dIdo5ldHKJIgk+kZGkad/JQsfDIaVAl7A06vWOKA781jlGu8xew4YUkqdQqe
nVwviWkXA+WqQX/SU2L9CtCxPK8nXqpHppp3IA8o6Y4zN64RpwJvuKROxCuVzqRI
HcnM7vgy+Vdi9pDxBw5JCFpJX5ZO+W9JuyOkXMayCS2QFqtk9+gFLdp+Bf/xGom9
F9Mej1dH62fDgO7hbtNhbRhtwaSuLWVz7eHYyUEQxym5WomVJSOq0T6UOj77xRxa
jyxna2Y72HCI/IdfXz3uSVu0ZpQ/k+G1n1tGH8sLX0aXUZHU4ae3+9gL0LWbktYI
/+BXmBc84RwotTLO/7NCdJpmMXkj03c13y33kBSCF0+Pr6MENrrQOQ6IJrQk7xSn
Pmfgib/+eqQZcrTSF0VuVcdRsUSZKpbCVMBEjoF2UQjY3yNqikEPQEb1mq8XdE7N
DWcBDu/c9fVtXmrzicF0VoxTmgMNqj91up6Jismx7I7UB6TNeFFHmABmvn/UAd/i
MJdfuMwCwwy39lpENz78oCPz3oyQW/+i7nf1gRCjF446FuXRN7lRirbVDZMlVluT
zZEIUXgZr1jSuUB4gsBsD0ZYCXCyBGlS39C/RCCKNPQaPHIS5vfybhqT+PjYzbwl
YfkzlOFlN6BAUG0UCpfAas8DI+FVKgIToYBi1N+0XPZYB92OxQ58pWDbOFClTFxu
G9VpXCtqWEd1JnVLTcjZjSLQkVXay3KsXSCWTGaYwfRAVBN40mOhyUyy0NgSOSZC
y5BklJ9p90OHwR/skVPgjSnBTjlkbPl7fK+hqAjqr7Brx+80x4e0G/Czx0HMMTDt
9clWyunLPPilVsWsl0UEYlgHicvvlfL5SO103qZBPiamZnzt+awdCEnOxaGhywaY
JUcIsibu0D332XyguR6QOjIFSHegCXryKKaxTgrwjP1kQp/HQXzQ6Os+oWY9QSpx
IpHtwepey8bvmK+2Y4X8bNpyKsNbg8a+kwtNfbu5GXH9XSvNzcRSWDElqgvq9RnI
4G3bA+DepznYhXs6R2zyZusZZxw65dJUCcxfsy3nOT58U/m23y2BaLFOwE4wzFF0
qWXQiGnzEgu5Zhtd/f9ybI8EEMwE11iXSnZ3DEmDhLfAWlPAA7iePEI4h5zfqVEc
FS344HfOz5o9FEDT6nWjiSJoYV/yjV1fhE/DuvMWaWKtZ2LrDZtQxk5BYQ6dM6bY
WDQdRuFLllAg4+deYj1LaqH8mf3ZLvMtahDldZxnObNI7JD9TOZ8w/Qn7/oeHh/w
uiY7YnX8dgfr8iO6p6Ziehx+cFDTE9Arhke0EDlIsvpN5/AnATIefA2O3gYqNd8Z
LXRQwgNR5M/KvsB6YXK/Mc3U/xfXTheiqQFbJ8djRHaVK7w9AoT19V2lgl8nnn12
70cg1+L6xvKYECYTZI8Z3/FNw7UTg/iWSBU6F3UYAJcoQgbgT3efp7omAcTxpwNU
opB6Ofn8lsiFd7tVney4i5vA/+ZE3B4fIl5HFnDLNvqYGQd32ER3SZHCIqj7JGcQ
mbgi2Ddmu63n+Eh5K5shHb/qWG/b9Zd5mpF1Lkyx3m6XY5KY/tqjFmPULHvm2ucR
FfORs9fpHBhCOa8j9A05BLADxRLRrq0zHUPQMWAmwG6uFoZektL37f3S2Q/CKOo9
d3ZFoOsG5k12kIY3c/QlKLxEac3w3iLuZANy3tv2BUBm4vvi4GFOnnPuSgx9/U9R
RFqX5K9cCHxhFgMGH58M/EikbyI8ROYtBNRZy9LXhaHHsNc69GhvTsK8DRWq56tR
Do9PDH5vVXsxqColwaul4QvUGpw4YGKCBOmtaIuNygYajW2hYkyqU/fdquuO8kzQ
fgveGTymiLwqbm5MpRYjYwFCi7O+V1OUS5XhQhwlXzt1PDxHzvRbu80LJhLNpxBl
V1R5GXHsl4+2SYcU4LJJl8j02XOKqYxNu70PB8FTfZHIjfS2Lf2yNSPLZseImayn
aSo2rX57Uz/5C/qPXHHA3OlV9ZPMdzQA5Y94BIJ0UTPHdUYIcX3psQn9Ty1FsN2j
nF2mpxUhoQpqL2sWv3/ReD0Ide7pYOhANvE5O3ErZeOaQkfjxhtZeALPMcK/6o5G
XmC9xDOxa97p6Z38nE9GNU5LAMEIewOqOAwO6VtlMMtpGmdGwc+YEEwPAXI7OmYA
wcqjpKvhpytvsSo0C/DI745L+uuPKSkEb8sr74SavqtSOC96/6KbaXp1ti5xDUPB
UEvp2mgXbTbk243XdOr3XNpIOV6v+EBjX4tr8ePiuC3EIo87a5Yyu00387I01Izw
jLvjbPlSpeYZuYxDJkgWKbEWrgANJwBdEEB7d1xCINlidqHw7f/q1mk+xGxgWKqq
cq85M61UMqoc5++qxZkZJ1dNiTeWVl85dA2mVy8j9cb0dnYVaxGizsYsRscVjdcr
sYdv24MFeOXO3H4IAN00TQiws3oVmP4RGKH6DAvgz6Mr6EC0bZcwzOMLAG5JE34c
vvD2qg2Araq/qHtn4qpxAPaBfvH/34Mrw4sWJMhd/OndGGSCQiRH1Eu4mc64mS4S
yn21ovqEDVCJkwdSI589PgLhExtVSdh+rNQIDRJD9Zkr04WoFGMwhCEU9Rph0+TF
1q2BjZWl+zHq3Qk+wbmCT9X4DL0bKtzZXFQj2U6rOwYoeyWkv0GOg8S5SFURh6V/
brAiJZi6Knsk/SGHP2taDX+iwE5BhG9Gmb36mL+8zfEbKQWVTvrwVe+dq1bEnd96
7w3CVk8/w5dYIfwM3rW3htUa0ZtzoAkt5cH26YUiJD+Ppe3zvXwE6aWf2e/Tw/js
jKPk2vXpvhqY0wmzsT5aAP9J7FilJa6m0qkKYh+DjGpcTh0VsnOOuk7Ya1IQ7dxx
ID59FlQUomi5cdQKnNG2iL3jIX2MMGqSwwnv68UKdmiyvkO4z7rsifdXHGmJknZM
5wj/evSLBU2ZYZAc7GIvGhVmyyy06iEvydmOdznC7Q24fdCrjcR4IZWkkKRNRsE3
ljmYumlTA7lAte3XtfwViR2bhgRSuy+f0Y0e3JVp86PwOlOXyjeDE3jLNU8ut8Uu
YmiwVKaW8c9kOUYnO4JJnwsQCLRV7k5tWLvcxRhX0GSw+uumAFKFBWQaabppLpFC
lhxxA3hA4XrkC/73DS2RTJuC6Pn6+WDLstM2qQUsJTxVTP8Ri4gUpEQyXV+KQwmT
gGrd/7iwS1tL/M9D4gcmQzhOPkaf+qtZSFUZY7c1a638RYRKZRm6zeaYJ+UX+Ami
QUJwHYoUv8+emHHepOGaVT209HGznb2HtcTgU0NaogVm6dPQ4nBQW69nL4Vqo6lm
RVEmAKtSQDKEWnnIwoHVF0L1SAkLuVDwvPu/wxAzJx7ryeM4ZUmy0sGVHWD8YeB9
/dk0SBJfRXFSP1jTYOcvTqOBT8zgXdUuokuFgVPzP6/xzDXOKOxuqh3yVVUGZbc7
6GBdwkF7K78d+aD1fTKB8zoQy4/iSh45RHZr+oz/UH8OYlTVmGsgnFMH+cLzdnvh
6LagAGqBx+xjDQgAUhaJ1b0g/FvqzLt9FymineqX5IQ8mrnU6Bp8j5kNh4YXA5u0
UqIBS/04zkfErTWJsGOJUeTkl4nsChuPKjVawG/0Cn8Q3rQhNGUfkB6yKl40o2tV
exMKhReyePWHDg3UdF+26M/+YjahPOxKAZI0Ly5QBVZ4nqeHSDaVW6dxHHU0anDc
UfuOhV9vb1TVdOhU8Ty9e8iSECTUR3uwHp4VwZMCfedKuuAMQbC+RGE9cJ/963kN
opNreUYZyPKxJwNmv+AeUwX73xF1cUx9t6ur/bI6N+RbbnwUU9SFxRfhcnSz5fr/
+HF/9gEQidLhtt9MRYN78MAr8ZrJ49fBl2cRN/Mi9bHDZMAw2B4pOnPspZ2aL75H
dW2Ge6UGg0gsU77pOwPFvIDYplXjynuU4GZAn73bGmBQlP0cxc+2chYxJRv9j9G0
Tu+y15/xlYRWJu5TW51Pe8NZ+WOoWJ3hP4+clGWbrZEaCtKNehdNEvrDs5V6SyZO
OtROC/7zY5wmW0huxNr/3727+CD5utZmx5ZG7HN7504ecYEBlFMhNXb/e7wyqcI9
PX732RayUKEluGHqIPnJg/w7UjQ4JVQ8aliBVhTrFfSbnwm0ayrNw95I42Pr12lJ
PKZKvCFKnidA6wLVYUFMPGc/YN3Y9XOzF5sCtFQ9TzuauKGQ+gTLphKXPxz7Ygxb
lB4101Y+aRrhk6pU89pw74NTnLqPwigJgGEu1XkCJpp5fpEdt2ylShkxGKHe1AIa
A4CnsMTCpf+Cz6M9zYrTDC1pOWQ872ohI+Uo9le2lyIytVZVJumXes6u/wOn2TDj
uYdHa3jXfngwjGntG/ZRXcpfoRhS1/YuiZEbx6MVoFnUQ51E/ysTNYJupmEXYWlO
6trBSv3861agkJ4WAFQ/qia4pziPEi+4s8B1G5815rcOcRf5OnC4mhUsLuAsoOMW
pvJNfrWaMwXq8q+k5ACmHTgLOakFMzZy+i00m0Q6Oka+x3tD2OKnTcbTGLaLYEh0
MKsicYLSX57JyymPrAHBTgcDEgttdWts/qXzgOHKqYTNCp91Q4V6vJUol6NsEyU1
HLAey2XxME+xGleG3zl+NnPXKKAIWaPmhwa4qIeaIfPb1KK/6EdAOjoRards14He
itFcT8dxdnn0xHECYqpqU5nwXmrLd6NDHP99egyoEALBH8CVrzT9Oe56t8tdBsw1
BW9J0kQXO18dWprLXgfqAh5rr7obtPYBUee1/ApgmWgWG6NkCEN6vB2dtAQhezZE
+6hGz7MVMmD7HmKgPzCQLO9gb/BiuF0tVPX7TIqfzQ1aOmtqpIk53APw9tH8uF+P
cKnzD0iXrpHLL7wJ/ye8XUMQyg4Llv7YAsvdgNabEGqFZksKCoeIBIJiOB5bBAYc
RgqdjlVhh4N0NPqA+Ok2zazLu8Zn2sHCLdjRkJdEiXzV//PBWTqiv0gtyN5fQsAx
WtrVpqQphU+dvaC1rwh2ZF71kyATUZGC69Ku61t5uCyj6+IGDEkXrbVEeTgVlfPv
UnzTx7dZDOvjMR9VOCXAQZ1ggzMVfMH71PSb1sklXmvGduuJiLOqW32GGOi7XJDz
WxaBGgTjIhAbAz9zBqJ7a15MwYEzwaheP4EiFaVPMYL0yBy5flgYCqYZBXM3sUCj
pL/789R79dUm26Cn1+Jvqi0N9+C0DR3yVP6T/Z+hgI3zJaeLbSTw1+lwuR6GZpFY
0OUlFBq8fjBIORoPOxE7x0yZ83PFqO3rROOBMZSOSOZPfTwBGF4jVNr3oNJVR1zi
oaMX+eY8sA0wBjPeuKQv97IpXqaEeSgzXpbyKC9m4q7b+snXjwKLo4lon4LphaRW
UQNrZzTvTW/TyDYY2SqdFNyInwIO3ji0VsIKiUzDnzI+UjTWOQWHdIXqAfbsJgaC
Nk7uLbEDQ7Y4JHYWaX8jB0+X3Nrsc5eFMARshHtNmEnF9k5pB4+zDfch/AGdgKp/
cxyeiXkd9SNnNMOG6C7QHPw+bYPGJr9aBIufSXGP7umlZFPFEFI7Uuel3H/UR+PV
E849yTqXYDxvj8V0q8kzh7qz9zvozFQwIBuVS9a24S7ctL7WryZqg+yIS6uKGgIK
dyUEJVQ+1lWrN+70EmdXvpH1FKLZdl8uURXCeLAiE6X2Jpb1IKhwfKsznWzEVp8x
Q1FLiI15yRPa7TAS1jW7i2i5Lggjh5yQlasdM7qeDnTU8oM2eYRcM9QKICPSy4CK
TBLbTgJFEWZV4wLmB7WC52KICWBwPOAzRcVztzY81QNtR1yvLMcsYR/8ZUCDxsJm
sbBQiHMynZ51MWnUSDNQc0sx9gq70lpjo1C17xddGStueY6nSNIl19izqklsflAm
lRuguAg63+LmpCzvtg6idlFQWvIjW07NI7gE23ZGLnadSso8B7bkOrTW85cChVPw
1vqn/3jdw++HyHOC62lepyRya22qHFzdsxtnUgFB2CEzOL3q/5dFGOwHVsyVzG7p
CVCCW/Ae3OmKnX08JoNRTFAnZq9CicrZDvmPkIxsiMjdAVPOmd04A1Hu3YQCYTo7
c16k4oufFFt0In8HveOXlbEsj62LwJ9N4WqYyudg7J+BJBidrxnlmWAvMxkrEmzy
W19sDOrPohfft+nt1q3dAGTqRXoAl0SrXKoYfmntSogGepO8yIljWi5UBGawEZbt
4yCIOo684aAPjBrfof2Pp5zpoWH4SJBvAJU6d29d+RqRmss0cXDM4EzkIVUgiX5b
retXfgIszDAaJF5IIQVuQ0Sc8jAWMdPbYj6svsOXMipOTGyGJ1vG1KcE7FhKSMkW
kxU1r+fvIVfBTgY9qylarNR2S2S0rrRUjHE5met49xghnKNIjDkWFiISon3ce8Q8
yybXvjArM1TyZYX6NUFSLYXJIgiSm9UuWKsxx6m9sl3dMX2Rty8V5OKYz0YZmW1W
NyJdbCnLhR3ForZQrOjVrrlPyS0VBSzK495vE5w2LufPesyfE63nupnwaK1mMDC6
XHAlPm2PxMVlhrwWt6wcytP25lxY5A006abhXM0DtvcpCLf/wPUUgQX8C7R6b/si
QoYqC9mrokBhhTgLlDPKGP7s7HQ38wOXKBLgk8Q8d1nj/c0E+MGAKfXVj9OIxbQt
wP8dD+fcW7J9oh2jZ7cqnbaYselPDk77ds6UwoogU80Kc27wkzisD69HXUfz1OMV
RiTcAG9+GM/8160I7mqrE9FlvG0yhyz05EgEtPl1bsmzOYY9KqJQg9hRpz1PyacX
QqX1qLKW1Fq0gTRCyyTHvBr4aHhk4FaAW8tsEzGSmDSps5LCVP2MVLuTQJbGpebx
oqRfCWGpupA/ae7w3L96LbNzn4cnzftsoVKJpIiCniuKdVu9TN9s/RuqKn4f49c2
xsuQHMydfXxMlD3czesUniQL9ETWIGVl/evF6UtjypupaEVo6klXrrztj5IgjcC7
OTxQs+b/56LCMtuQ67VU36XY+xFuihoniOxN1Nv1QpF8FEhIIxwjlw1fBaZKvYaE
NDT/ctYztO85FBUyxPG1QspS891BBLwP/s92RcKU4psJdDPkvjY8VL4rwANak6HI
Y14w3aoplpFbT1MqVx6ub2DXy6MC2byCdeV/AcD8jq7yhXLTdH7a3JyTysw3oger
GUsE2rZ2q9kDz0XfPRCOmIB5dsQ5TA+xzpR1503qbfeQxg2YPlqHoA7PyKXm2uOl
keweYCJT5bzKP+FDoJ1s6/G/0kz81RevNHaniVMYHZOcL+VBb0g3HofjTzBhLJzy
7c1Z8A30jBIiCsMKvwD2XYWTctk9bBk/scWXOns/bhc6m0ldPjkYhJTelGtCj6et
ackMsaJZR1EI9aBlFgw97GHl8v3rU1QHv5nMehR9z6HIbRWVNHi0rmwojTokjtXQ
mSAyad0rvpESur9B5iMN+80SuqchtjASN8Q42hq2UHUDpeuEXdvkNjxsRLKhHUeT
Bt4RJ7JNYW/AoruapRxA6TCbJHcXBhvKzAECjY34mykkcCHcK6mufAaU52GW4odN
Ogr8ihuw4SrGkYY1vxJCvzXeADsHhKfghbbpxowCTZCPDOuA85F1SUO6ZYXAoh59
5BZwaxj3d74jRySoZDsoCYoDpDkmE8k5v7y0bu4cCBJIyXw1L7ClGQRjYraVl+qx
kB95Myq1Yz1PtK6PJzYtQSXjHSErW1HPal/1pL4TweMiKRnowAnh2jZZQOe6J6Cu
Q2ecyJRn32hu+DzbVVbIGVJtXi4vkr3JtiP9+e7cgsLN6X3Vunny8XAZkWZSfZ9d
a+P3IEx38kfSuerpak618ywJph2j4KFYn2mMofsdb3GwHA9p6vugO0tGqyQTPbD8
YeCQY/b4leo2C/ARc1c2eWtnRf6hSKBvWvErhNMMlUFlbIvAwDDF2kYGXL24HyZ3
qAu9msi6GEEe+ik06Ph5soOvY6uM4CrK1DG6HTPx3pWrxLTTvikQV83xemRDMfzL
gS+Vhib6sziqI6qnyUSYMxNjt44SGPRW3qk6E83JvGk4f0Sq+Bxq3tLFLhqbFu4+
gmlHMtkloA4sUZChqYXJWJ1aG4D048Dk7BboXarSOizDq9rheweNEuAXWGwOhItf
cd1KGDIA8+N/eIJMneYlnmCmr9WMXy18mLLsQ2REC/BN06bfruYAnMa2bceI/Kwb
pzG31uZgNiBhyi7E3UrjnR6DnuOhtshq5Nh6URjbJiAAumpJnSz4A6AHh1rvmuHZ
J8jAi5kMvAbpbUFjPMjPgTsYG/qwA6DbgAXDlKmMU2sJAtDPr+yjpQXPh/BPqjZa
jG7JVVTRkvy7uREwRxr7p0v6MIiWQ2L7wfcO8gczHKwnsgre0MLYirY7Ra9HDRt+
RwFAqISZZwI+1UyY4Qhay/wWIi75iT/vDFq6fYLvxv+G45glmJ/khW2HmYqmJbo3
WcwFs1E+RGENGkATGZWehOwZalaR7q0Jy/tGKYighx6en7ZYaT5losprZAlQ6TGe
rXemsOUcvs2mF1J6DxV3lYF/qRwsm496XAexdlv8QGpl/Ew491MV2ku4y9lS3tQc
e+vbz1BZzZJLy7W2nXKW25002JFDcJnwanr7xgZVxpWx2Wu0M0WwzMqRo+BW1So1
GidNe/S9UqfBA4tiFIoYb02azzYAjNEupJZfnV5r4ZFiImMCpjN4K4jylxorCa8F
YhRjQJC2mXiM7yLGj+xNBYm+2Q/5UcjeY1CEUn6dw26s2/waQfNDCuIqF14KFgu/
/s41EEkL6OlKNAgHEIHs/DV6WlHWw9iYPKGcEBQG6XVyIeDiIgiQ1C2ukKJMwzAn
Lu0ONHZK8TrrwbtajgqvkPbrtDtGehEHIBIlBbAM3c8vDOoCo7lgYQ543Jsc4UnH
o1RFA66c5M4idoavLDdt0wCIDI9ATqAzMlPG+UzxCgm16+aiuRjNM53hU9LY3FPD
LELJ+9By6r9sKqlkCTjFIEA+wcnELTRWIszQ6nFP3LkT3Ose5j/i0NPzy+GY6JRt
DwOHpSHC/r/1hy9huKRB3wqeKdyrIamEouhhkbQR52BZZUmEMb7ofeXI1irpbUJg
wSxjnjeWMV1VcgpJB3aWYa5rUyJ8xuTuO31dG2vBYYfIeTfJ+dTzuyTWBgiqQWpc
AWXPSlCK2+S21YYdSL5hxIzuGDERRazRw24ohybUhoZeQAvxn5Kgmvodo4c47lsH
n9hMAN/3P6PIzAYRJ3Mu22yHuirYTvCuq9FpeYXd3FEhlRhqKfulSrGyFFCFtxbi
CSztCU8DogR5wen4F18SFzcCSTKCc7pn17VnN06rnN+olUDnPCJ7AuljRuKYlM/H
spZxC6lNb6xMV5ecYZV9RN+b5Ps3RtTB8EUNkOhqHWueo9/+r1owiX/g7fbm8xcE
9R+yO2kzhr77IlXuGt5Zc6/LD7v8rJJJd5D3AU/fBURXKZDYxKRzd1Vdciy47eAE
8LwKmEKuCjL85BjkBkPHn8BVihZziLlm7tIvNjs0EK8suaHeDZFuCn3Glhup6jEW
3OKvJyFhxWFJaMwdbZL2fLLC9haXISGILzjRbA1AgllccmIdz4iFYVDMRxLDo08W
9dviE6WdVgWAPS7K3HTDKW87CNGKUiZNmulewKRVz5lZhZSgjs9qWix/Zefp90lN
p3itWAhgs5MrRORjeakLazGxxsEtAUq1+gnR+qU2SvFIxkdkoONuI5vyii0YCMIr
PCuCS1dVyKtGUcynPENEsT9IUDsSGjWBA3822to/d3t+QposGGwRNeTmWkLVdiJF
zSho/EfPrzsTCtxO32a+8cbTYKYv6mIKgmjjqAfx17+x/i5eSn03nT5x/yNXjiVv
X1tms35/svjyzqt5Doy4AeYsNTToudi8fk+YRWQ4Wq29zidrjoHGuyh3MgPTLlVV
XaTqPDlIdY1/U0DVakpSlnN7sNnzUunqrQSP82ByhWENU5Fsd6DW+8qZQnQO9Ppo
RMi0JbMNMMeBRy1ylmnK75B22p6S9L8oBEyxfFbw1gfF1UeEjTN7Xu7DQZOEY7mv
FHno43wUv15sLd9opMRo5BPnQV4AZm4PVyl2Q0NJi+LARAOgHr5Tj4yUbEfM9S6y
3Yg+YIX/9YwQxCUkmr9MsauFylz4Dgkeqm8uvs+oOHUxL3cDFRx70ZYhr7PLMVWe
B8gWe7F0Vk9s0HMNri+9I33pGyFnW8RwN+ax3GzXIsipA8bG94/R3kI47SBJnxv7
hIkMD+/wjL78r0K2UOPA81s2Bt/oPpGoBngMTtd6FfJsrXq1F2IVHLmhTNGZ6Tbv
a/tkvJPV5iAB6ejIR3tkUlNIGd9nSZfV+pODqfldoWsjOt/zpDWzVxH3uXbnCnwN
+GJ9QQI9kFMwuazZzC/Hr1dPEPRsmupFPFFaoWKjVC2ciha2h2CyuLMeLn80GPQ2
684+GVbrv9vh46DknPQ7BTQIq1+u0RhSPMjFSVuNkzY12MRVFhzg2SA0IH+q+7dC
LmEhn6j/qUhtW08WFlHWhJHXreHctbRt2KfJgasU8SquJc8qatyz15n7gquSGKXV
z6QPeC+aUPPzF9McQoKdk61TMBaeK6o6GzC51mhwk+LF1JKRXJvN4nAcB3dtQCvB
uwMMuwPQw8uXvPBVlNzIaRpmtXNNDsG8HxEmLw1NQj96Wi2jAvREpBjXizuQs65d
o6gzoJrP5NohRGoxHk/Ur8NiIKRGlu3MQuKUx72xWEOskY0xA91xg4I1yje/SAJ7
3qTi74ZkCyasvgZCjNnQqq3HykrqFmIuXl0GHTDVEZnz3XA1VZUo3f4PEFdbnYEO
5/UMJ4dH1JwSaSaXI9RAKxzTqalxq7oxz94C/T8enE0Wxojit5O/IMsg5Effl5kj
LFzOF2Bo3NyuLRVCqDOj/FSmVL9GxTRZvg1nJtMZq+JiFg1A4oaLtmRUnu1XWG3d
6xRm9N/eJn+je5GCY253mV7iwMhpBVIkzAHL/yQTYTyakihr4rGKheJltJMuUSQp
iod+C9cskHvnHeG4ZN/XKdG2XQDCfDOf6XLgYstl0KWHcckFqlvBq2dPsUe5/Xdk
0jNHQi8teHQuhSplwQFC3gYqAsWATZC3RAt6dykBOaEG7sne3oLhJIhNnzh5+QdM
nU5oTCp5mUfIwnq1PieIfcojSDRKuBqp9ZSRs2rXuPxYMIBAxosIw6pfSus1sxp4
Fk1NHT1hKe7vxc9twAvhpN4n5WCprLYZZF4ixnHP+kukImCIH8nbUdBciWiHnLqN
zhe3bIiddi6pxwytS/vPqOADEov4eZ2QkuC9rSPajQ3yZTKR+qXSwJUiPlNCE7MC
5xBgINIyvTVpD9EqfTzgy+TSanD15oqrl4qNaUmIETcEDFtFACShTc6bApLRYh6L
R6R9VrjVFZXq53I3AhEmyCKrP5uAIQnF1AJ75dzodLCbbT1JF0t8FYedMD01oYJ7
hOWH4eC47Eno777t1BE/7aBdv0MFQPaF2hEIqoYvGVfAGwcus94lx5rTNuNv4/AQ
zAJgfYCP9U+K2cBGFz7f7pniymnTXvlrqqd2Ca9NRZdyGitI6Bb5d1sHuxgiu9+t
DhOX/wIetWLV2I06GwkwMiI6jXBRXZ4pbqGdhPl0rRrIPDQbQVtFoy2+ahq0+BAC
OGaQLfq9HI/duB1QmcTEo/iSe9fUuhxDj7wb1SUKMmS3s0mN9oRw7j17lQ/a8/p7
LS85HrKrEO+c8NU2i6mKqCV3G8v8vzR1TyTDctRijPAwQllAdAgCw4ToNbEqZtws
dlNyEgCxmKVKEi9OjVE5jc8myXd4liUY6iBALQ/sRSvitthjl8sCvSB5tAB7wCEf
TOGsLYluxvGmeevIMEb3cUcfiQ959MxLmJL3r48AlSXEJLrq6XBs6z2F6j7W2BZg
w4cIgHWgs24138qWL3S5Kht6uGodP2KGN/Y4BaREEWptxyld/S4V7yQRW0O+PkOD
WavU5loKxKKFv9Wekm5plOd4FcAzzomb4Bd8r9X7QPtsSlAJMimMJ/2TQkmj6F6x
PRjyGIuzeI/F9LTdW2vHbPJh0nrdnFxywz4smGhf2vKKQooekPaJ7zIY8AAvm20i
r4PZUBga2xfsMa0HJMSGaEObfn7UUTMjaoUSxDdfJnq7XqIQNGhXztvunOawlR3s
8uBE5cuptALz3rM/ll8nDro9TBdUV4ly6Z8TP82swh2MPBVfVMqQsNz7CiHbG8t6
CzR+3gA1EIps139tB6tjG1ZAZHWZtJjLMMPNmlch3V7UDHFeo9hhDbheGRKmB8/3
Zz9ZseGfrFLJXovzJtTNMbVfx2eflrUEqbyGN44m07RKxcqmFmP/Gk0lyB2CTm5B
D+OwkOeXv5bZh1gkHM+EquTRRSrKk1jOeMPUyXwLVQiMPrPgAg+rJjZrPJSdpKkk
sc/Yiaaf4dFydgfqEpDZvgvlCkLMNJXFF3mbiX737pcQBB3/sEXgd2QO97K4V/48
S2FLhZPEBj1TowxTV49a/UllLcMIFnjDvNg8+jpS5zwVeVZkAQzZNIxgyeGcGVit
4eTgtrVUfMfU7Y+RI4CIch4z144mgQ0VpaCboIsYLNqsJoryZUlfZlHyYgh3EeBp
WbVd2+G2d3C7vDzhnicdJMsXJ/5L6UnentzqjVFfPha3rDqsPP4ASXW2ESJSDxIe
InN+/fzQ0hv9K8v/2EdA0un7F0u8GhJhPViOLfEbVD7mg+YJJYJoXT7efpZ2RCp9
OnoTAMCEEWHk1EXOrq+1ApJxlbagODD5Z29KhGnWZARNKFZSqNxvPnz1IqB5ivv/
nkvaNXEUuuftOpVZ3/58CLaXDQBn9XSD/v8HPXhSC2zgTTj2idvwWyLb+RfcuS5O
zt93W5enaZrO/mUQeq4GC8yYbUBdkjSEPmt96EA5JZxSmbY9onruCY6Rreo59ALo
2UY8VPZtThLL0ItlZL/GlNGx+DzoKltBKBTXRkPuVTmjj5wEN3eBvjpLIOYaizw3
3lMXTJ8gQ4eprgb9575Tg8O+6LTSnHVZWweDnmcxVvekK2/v13AoyWsRBga9rlP1
26cqkVQ2n+45CKFlq7u+f2RgSBBdbnZRB0x9AxuLR8xuNkzk57N7wwRLzwLZWbrg
yeH4x6O5iXtDD/Om3dMKq/CCp2aSV6pUAiRHlnGnmlWK2pc1hHD0zSYaHNpRVAvO
4XAeiQDwHSNFkq1HW+p88mqQ/+PMpDNc7FhnPOX1CgVmlZSbWsIsYdiHP2QBci2q
Kge5BHKukCr2bbLC7jakCuYmRnjTi2pVDSpY+yFe7NGVTakxOcdus/h9q3oxRY21
u9IifXW6dCPsbF+s4h5QtioZky/VkExW0VVMRi7eHtrZu7CRZzARBlOg8DqFh452
MnxAVtDekkJO5Yqn/k0oU4HehP3onb6IkysLSOLDjdZH7IFW9PIStHx0TwprBe9x
EkbkdVIvFNV+C4Zdhb3PH8lG+9u6PutjHaRDyZZ7oSjzH/RflyBocy11wkNgymHb
SEYM7itWDvwhTj4WZ3mLBAHzC1BI/ZRkL5COjVtyLuNF6YF/FCqKoG558Gi01myi
vGFsaxnX6al4tH41bRNLcRWUoW2koCeXabKPvyGIGmDYFKs+wcHh7z+kP1d1sHKw
3LxBnu/q+HFcrOLypxOY6SLjxZwQXkaNMEEOfRKX7bjgjDkuVx0Ha2NU36DIPU0e
7kbMkDdBY/JXT4HOx+JJbCPhbkUDUNCeQwzVDycuCmUqqr1vLhhFdkbM69hD9h74
5+hkaImqeFVj5zduPvj8iEPjrClfMeD0wZULfB2nkgwRZg3YxDmbnnhEWCz2PtvN
hJbhcfZhZYu7H3j4p0YyFS8TuMWLxr33D0/s0BPpc0gume2CHTYg9kfTE3k+0C2r
UE0CzqAcd9pbDlr+C+r3Ld/JiUOD7WAgcnPjk5ENgZk366trCxi8L+5CQiFc8OFm
U5np1HMyaKMhoa16DyGZTtIwfQEj0scVhfPPv5V3ID2BcXVhHNgRaSCO1JQot3JM
UWF+74/YHFtn3u0ThprAJnxMJbaIfMQUBWD5HmVe//5qVa4zB9J8lVwEmiiTmwmC
irxaQXEZhkX0karR69kHvROZfBlVQjIb84f4vlYDlOKgiV48SU3DaK7SEIralR0p
vPugfQdhtIzWZsQwP/qDN2RMuFdxWVtQHeAShbC6E0tr9Nj370Tn2CT+vdazRfmf
YF2z6eBMIU1L2/yiKrK26dewhBK963aKUwW/4ZO8GVUzrmukHODS8tQydVb+MHa1
JtB2M2RYt1yTvzNhMnr7CVYko7MXbp4gy3eDUcRZijl8X3iVENHdzMzyk6SNeU5n
UDsy2veiy1uiXJjE/1B8V+Su46/uoKeLe85Ei1bYGdgydH7QHALbjo5LozOu6uus
Ky7Mttn/NjfmA6n+XWcSsjAwxgpR5FS6RxBaeDVSkNZ5ruE3V9QBEnHx6dMl+KIx
/ZIxPfmIfdomWgklC2DLgkukidH52d08Mrhwietrb3hTtm+VSSezTp6DYJQK3maA
YM58CScuKWbaEfjWjayVYbBlvEsnARloS0u0fGiF1GFq7Z+/EfqH8GSXdMs0VFHI
cBFJQzLzryCm3CDibuJh+rykM32bfOmghfnXDXrc+VtGJ3i7GO1RHy1EtOJd+G7L
o0MZLfpPfwOAmVig810gBvG2bQOGql6vbdXbbkFVg99JfC1u9iuLUZlu3XA9YcNU
VG+wxxGxyUrMjxdkywwoCsFn/D8rsHOUNuFqvy6jRIVWp035KskSt832eFR2Kjxi
4/8JEl6fXZQ7zQJSMxYm9Viz8zQYWJLWWvOI9xoMboJGITI71x3Llk65zRD7bU2f
61DxBNEG5+eeMZQDUJNJXiC2UguMNp66SqZbIrTeAnaYtB4NoFDmKRXKZc0A5ZsR
ANpD1nWuFNNPJUwOiVg0exphYP3Sm80pmd3sj8oH5iwqj63ka1F9T+XcSbDmrBZV
V9B5GO1eJJMu06s0OWIZJuB0+F+fU2Fg72pr8kFR0cYFLN0EOnk9ZpkX81OpIBXz
1ZnTIp3oaXEbNqPQr+KUN+brgvsu4iPuCZ+TBpoSUbumbZmW88x4bacPFlfHhvvQ
OXK3rmucM8WaWyil6MxgpEpq0uhjnD1/3Z+VN8RF97q8ZiGkbPtIukjddIClKEPr
gDTubdKlG9jieq9KEyLmrjaH8I2J+YkccFJR4WGlLT9p/72KaWHuQi7OrUfmyBWj
/dx7gKizoVY95GE6c0NuLS19dgpai3utCldZSvNQjS+HP5NKocex7p/dLb8Jv5sQ
ZuuUfLyfbjG9apbqycjvqrPD4UHkDw+so5JL/D99Sgtn4l4Ka0odne5k8UpkWepF
OJcg2tnSdhA8XfwUsi13RP3v5N3xmWBR45qnwZR7XyaMvG9lNjZWpgZ6PjU9Mkr2
tmHeMan/RvzMRU00V2FpTKIooxAUAOaAcymrZapoe6F9gCBGFOYmm2CmfcWQGmRO
p9N2O2GIWFQBZhOdc27OFLQk2ikZm9DGJsvbhVq7Hy43UKwwkDKzyuVczzX5wT/Y
BpESJ9FnyvQzvmfZuppTx4/ZOPvqMYo7SUwzttkeY/OEZ9CZ9QEHyxvuIRg7TFRo
fjXwl+vLfD0VpsgP8MwpW8GaisDMrQ3BsA28WfNtW4b/9I7g4hgY0AR0Mtb8WJWM
u+9fV67j7O+bVnetWMdMKMSWybtUvKPhFcRQfLFCX+0mV/PvlLLJiY4FAQy6E1/U
qV9qIMFd4lBqcLUi2APaGdZOgEL7pe9at2Ign2FHE1OquozZ/leAwoc4vUKTslU+
FgVXe/JcnNilk+N+260eMS3JOcinMHa2Nj/ZgtObNMr7lwbHw9i8K4UD21WCy5vl
OMBgN82RbgylA7HwjxoOwbamDsjyOnn3TB7Vk3g+cuOYJZ8mqEdMpDCYkzyuqHYn
TFYGS6qHqGd1tGzDldINtMdDrHe62CYmEwOf6pTYdSZDAjxEWftrTyeKiKX7onac
ho/tDTD0QvnX63xE2JhBXWGc9rspAqaQIIu9v638vdksdK/saPfBTEFDvZvVf9E9
UQeD0cVhWR6YVg4+jxYiY7ZTgkajC7V6Cuw0rd6zWMICj+3yFiKpbs+lAbsJf7KY
6l8U2TtfnU4Tc+j8hUWat0tIIATt3E9h6tL66Tjzv9zrqgw8AkZZFKHo7Pl5BExC
DRkQAymX4/GP0jf1OaVi7TzPD2WuRMk9kLx08/Fnsg0mO/PFXYRiPScJ64vGwG7/
+UkdhbATS9RLe9/ItM59f9LnEo9B/P04LJ/9YIXf1O6quOyrTwWYlbnW7+6dasvz
aWJf/7w/NEfryTzYwSeXvnEn2PlTlT/Ktw/fcINp3tAXo67OvRrtB1krZOGu2ell
wGmVpO8mOj+6jPpPO7qh3pJpXtX/rIxBfW0SAhtawWG+Qv6AyLBsWhptIrIXMIJv
JRZnd2fqxh254NQZzp23cBk3fEebhWdHAm7b35jjcMCRHEKcuPe9iuRJzs7FVTaD
eS5fNrUfUtzzZuzUziFXS6wEN7ouFJ1NS9vCnWfvJOADUdW13+zhYnhU1Clpzhn9
3EyUTc/TqJvTXVQY/ryrjwi9KJ7S9Q82nYeaDvtoK5xMbQb7F2XKgcMcPEHp51VF
W/W6QQRH/ssLik8wWavke3kXCc+9BWIIQMl7Ggx9NFG5vk3YPtE9SO8jYBqNnIPI
H+UfG3TC34sVUPXuHXeqH0/YtovmQe8JDyXQGgU6PmbmOUMy8TBlQQszioJ1dOjK
/Rutx+Kc8qtUZd/uDEkl21Zb8m8S3Y4m+hyv+m4HtTfSxycS1PagyGGkAypKJ9WL
cJoMo1MM5kJcdyNvIdAdxeSUa5i2RNtAI1hU4JyQKYfyGgsDCjvAakCnHleN0iCp
kmwG47XF6BVa6y+c4wMig/IgN0IOHVP+M4pbnCJ0pnolmQ3Kz/JlufhIpONRLn8f
R/MZOXEAjwUCaNKgTXo5gxSvLRcPDBQsZc4GPpgV1qlFhLQCZA2Y0RqhublIfLFe
P9lttPbeFkje23KUjZcRFJYDk+oMJoqrIsopmBzEk60dUCQ19xcRisOh4PEpuUQs
iGB+KptHdDS1Cu8BgNZmMjdlt9sAL6J9M5OcxmgpKRG+/di8npgwzl+Dc6km4Yxi
JztwVROrfM5ErqmSQMAH0lAxp8O/dJcYDztPXEXQYyvkY0RvrRQ0Ilr/1mBm7Vwr
Nl4ZBEVJSaljIz7b+6CcNKOpfNKlDR915xl7aOukTcoXF+vteUBQx2gggBagldD4
FGQGIXoAlh96tMZ3W/so1RuF33zSsG2K8HMchN9ZJn4/NTB9jahO79PLrfH0poN3
WUlWI8THZK53HlUA6pO4DtiT7nK1Sj3Lt8vvdGNRB0avHec2dAmipGw1HP9MUxeM
cvJ58iRgNfjqNFDXcXSLzXo0Fq9sQLIhqEg6001FymEABStQADaUmMfOjQ9RyJlM
O0knVVyYd4N1AObP9YeIDXhfAJbxBVggJivpTQXoG/jGGz0foNux2ntfNpzwqJE7
ZqwaSpvlcyoOhIzSriar52GxAYmz0s5w8Iw9i+VNqprDWNnyNLVD2Ak60dVgCr3M
6nNhrB7aNB9sfCF3zm+ZgTCaqRr1L7idwe165EXzi/hm5zOPixzbwX82BnWVOgq3
UxtebbkufAabIILGWqTJpOpQXvOHU61x+xEs0lKZJJ65X9Y6Cb35vTJg0BVkW5PA
Es0upNBhesuFRKeV9Xy/eQ7MqyJ3zkXfoWR3pCipWrWCwetF0nqSaQmwuhORUwbi
DNrzgo/15SeK3R/RtNUOkcdFC7jjwm89ZMI0enPJzzVAbehFULJa2iCtUqS2bo4l
3prhOiWyTpwxf/wcuRJoWHWyGNms+18a6rcPnd2eRVr42IeCqLloTBniYlrtrTm8
JjQdokmoMJdT61WHU5bZve/jK1kO2uUaQuH4b/DyLvqv/Es+CJ6teUv36qa+ha6z
n/PaRRFqVDxUleRWgoQXmeD6IP25vJSepBGMTEZ8+ZHE5EJlSD/Z4OMCEGVwfpjb
EZgWg2DWMKxOxxGWTCOWv8QwArrEV6R8KCsPgI9a2En438yWprOUxZPvarzgeMvH
QrkbWMfAdp2FzAwE9tXt7AUSjymWyH0jU9zlYO0t1tnkSCihnAS2K//pxWfWUafk
VigVR/pYzi/ydk3NvyXxlvx1kvnptrAHhsydVSdBksZhtz2lYtOGrq5XNB67xBsj
mh1llfrhXLGSG3zLCLmqze792aW24HXkz15JfCybs8LiKWv+IEyuPE7hiLRQcdCG
WG8O7bDLSi25VJpH0LvXUT3WPLc0KBuc12kE20Tq6FNOdvz+mIZrA7gmQuJxoY29
FRHEq616vOgsK/80gZ/gFu5ZljjFUiG4/iEMGBMrV/vDVtfQUtlhmWnm+Avw5KQV
MMek4n5eqUwNhcDbgGG46uQKJzWKBPJ2DRbVyfV72vUuR5un/re1eKEFEQ2l6iyF
rbF0SVHPol2eyT3j/t+cWPW1IidK3NE4ICXt3khd00+EJe6RQnGscYenbS580S0D
SNK7v9Cn3GT/V59K79qjPAcIj/KGQyAVrwb0Z9al7NkhnH6lfx3iiH12PqN6PNe+
T2ImHk6SRad8wHVcyE1Bb3mWNpVqhQoYAILSd6RTidEMtpuUvruUdIMBN/MJdYIC
DOqBFyOzfmvo2i0SFtVp5PtU5n1MkIgSg1tWp3hk2w4EcrBv1RIfbIJuydD0U2Ly
R2sf1juMhXzI++vzUweSYrb/Dm2P9ou9Hz+ctmwLkPsXf1vhu9ONoWV05YenkrHj
zyL70Nt2Ovf0/c0X489wz94Oc0oRMAyFr2zpPpzopBl4JqG/NN3JTqR7VLwC67KO
OLKbryVvl447DZjsMXemuK9Z0iJA9Kv9whos/A9PTSMvV/PtpVPTK0LcQjNHfKnf
zzl/5qGcZkghD4emT6yba/kyKKZBmMM7p9iros/cH0GRFLG+DFy/hoImg3G79Beu
2uQz2Ju+1Tm+96tf+Zph5iO4qAqI5ySd+qxoYVhb6tLkNbHw+9zKC4ltgnC2foRN
fF27kceJjEDu5LvcJsbj8iDfOGkev4x2lY400XgKmX06WqWJdeutflLqrsLQpeaj
z8DYrtZmvUyMHzc/awHfydNYfdzyEHeoLlw8BsyRPHno7riWXbXEnz8gYUzrayQm
1/3Er8JDYQE+iXCA4+JIgT/9YQFQapQ5TzgUFrUiDYV0F0p7wnsDN8tj6ZuLyptg
gE40qS5kSdT611mURB4yPSKS3314A68SrZXLxXb0oByME/Q0nRk9mpjikg7EVCOi
8PAtl500mu/iV8ewvedFZy7oZd910kWzt1Lvfwi3Q2BYRMfNGCfz+4kU4wZrD06V
83BI6TQFRoHW8v6olJH1K8Xm4ub13D52fsSH9vzzRQmUGyQOlPu97UeFwhq5+0sm
SMIt5wsqTJn0h2vD1eaxIC5rKljYdZf9pm4O0uHPqbiSFsni/Fk+vJ+BNIVowueJ
vWRml0Ea3sXLXfaOe3/rGyne8d8yxN7I/hAh4C3EB45ivtn6Wi5LdXAChdoeTbn3
7dDBYqy0jBNGVT1LVSeE3Oil3pvzGgEDwuWWVRi9dDhf1QGKF5BEukPFKdL2NDpt
IS3Jq3D4vv7z+5pgme/SgjYxxFVzxa12umOk1k4/qRp+MmHe7lqcoPQhT68ok3OC
qnB1+q6FQL/3LMK9unPqbjoWsrBjh6yJodkr+9s4NISOBw2bLaM22fuUHxrr4HtG
zpt3u+jPRgrujt/eir091H/N0/NP1Owc0y8lQJyOTijzdot9F3n/YyXgA76txp2u
pijWlqyPf8UguFAKeH3dhnQ+N8sEeZwDDzFaRa3YBUzvnPZMS1zyl5lfUxZRNtXI
U8S/lPc5wW+G4XqTKDvF1IaHnO+r5+i7u6yo/iLF5a4uGaF/4VNYVPXREDi2GUHR
YS4GP6Z2NxUhDKi3i3qp4ZU/oKBxMqg+C8VYHg18cRxXfYk2IffUZ26Tj+SDARN9
bAMW3na+j3Ky3fBXnWMo64r3M59h2kjtKAgEP0az/7xbi+mW3vaMzYygViYQA5+X
peV34gnKCMw3jtGqr8VnyhL6Ra1q5FxevQuKcCjxH43+BVVmxbuTxfrrFAbE+6Hs
nkWo45CjP7LJit0drwa7ybGNkr8VEdwgMuEm7LLRrAp3uaNkzlxShT9yB4pxyu1c
pxwEp+qEePjL1fTLo+Q7zxjXwmYiQAWdih9TyRvpXR7hNjJDFGWqoYwa9UbCT86f
HR9TEgBTll4Ng/dI7GCYJAx40jusUq6otP6km4G5mpo46FxDRxNNR4ZmCBTZL6Jo
ncAu0++w76BIn4BRDL+kh2XC6DXgPeRgZhY8tTIegle9fS60jZcU7Z3wSAKT5htD
3qEdpY7KThFOv2SX6VLzPWdZ2fRIzAvNjibKbi1anJ2Aw9a7Qjg0RCYSmf1PxvFB
kIbKbc1mxlQeUT7iPEGVzRLW2XFxrfoNk8fFoCNMRch7ZUHQve6DMZIUmwVECt9x
Aqqj8ITr0DtGBjJ7phLsQyJvNIDqRs9iJmtjg+uHS+/s580cgVIt4wza04MVz3o1
8s0M6d25uwrPG+RLzVvBk1R4gSTfhpLrzlbh7Aj47/QrxH5iiRevBOqDqRxnWkWg
1/6zY0wnRCjmfE/a7A3w/fwzLWnbR8lDdnpWv6pXDFoL78kUURjgAIIxlpIduQPx
zQvIwgoG7mRmeY9v7Vqtf1gw+j3kU1/biz8z+2fTzjx5rY7+Po3qRvUeigNpKbNQ
SbbrCHd9jPv0tNgvBxnWTKJxHFM1BbSZT84fDhIv/udxh87E6oJ9Sral2l5Glkza
PdBj7UKjTqh1vWUo3AsD++Icj2eq6jO5EabD72vihfBDjo/IDtE5HaaYGnqmpVaA
i6roC09elwJutMdwmIBEttqGxO5QAkDCSG5+YDNUGdduPHZ01PICa5foZJd90dC7
H57k6RprrlRSpRL3CsRCEFpPwMGk9yF9MVHcQuG5jSJWcTzzIDVNyXDvh3DiIxMl
YbkVfSDjjbz2kkoGm6y66ceLu26ChBstM+knBwGCzfUJ3U6QsxhIzCrJjVkehILI
/SMjb93ntUCD3LuwU6EUKBUgHmvzNvhwC2xrwh2W1OYOAzaZ0P+k7JNYc+U8ZolS
6WIFB3jlitXwC0GFmim+AT94wf3dee8DafDFKOyJS3ZVdfqwhBHtN+JTCErxMW+z
FvRxWgW3emPcH54vzLmnbpxpvpV94Oe7TWQAiY4Amv8vL3XYO1Wyr6o7WpSiaR5r
7VTOvKRE+ftRyMXYQ4xg/YJ9Sbm9ETlauqNY+H2vLAMJtL7PAe2kww76+da1K3Os
FOf4sCy6X01djSE4BVYlK+3L3AAawBZ2osxDHotiXVVb5PzEB6S65SBiBQDtI4ho
v58RHX0JSqhuqoq82JppRHnTSBh8UdnavGg4J9Ip5CpL2pBoLBIObn8Z2UO1guBs
OePMNzdDnKRysoj1ZsX+zewb4+Zp721YUj8TJ1xRZMSIB1PZxIEhwSm+gRUBtZtn
p8IBdeDxwMfxADeihnzMZsuAddgEKzhnPnaYT9sMHen8e//iJH23eseHKYLSzgNz
tI71Av+LVzvOvRvkE+NAJrVBb0DJ9do9TcC+vUfNufxiaBYgbx7kLeJX7cuTR2Kp
nE47f8gsuFhCthav7DZrZD0uvqJPlo4RowFvJlyKEj3bDRymcmlD2ZiNxGDl6VOK
XZa2Syz9IqbV9+m53yFcfE7Xj7mgJ18t1O/yN9BhMoYYF4XUBUufappCAJfYOQ84
oK2q9YbHmFQx7X07F+m8NqOuTQlEdg0hSpePyjl+csDNGCYqn4WtTRnfYgORCZfC
FgRr8DScvdcAuEUJHfP2hwjXH0/0KYekrb2c5midUTsbn/W5Yhc/uh5ToLy/7tXH
jH/mu5hQrRozUwQPbDQCfTVKjUt4lN2CUPU5LOxpU1UBK+kRn4dHcYIXSCC2pnJq
kZ/hvcouebKRuTsG853boRD61vH9OI6KG84yioKLXOOXEsitmO6V36e5pA1+Od3M
M8hVxJJwHwiX2IvDw1mLtGaSmllDwynKybb+4H6CXhyFhGJlXBM6xK9L0bOrLI4z
4qkKgIep+GrGdcUlKflbOW1UqjfLeJXRwRWv7JwTeWnLo5KXqxCbgZpDdn7FRmJO
bBg00uX8XomoIkyYwel+YSH2bLuM5pk9zWy72JNlVT/Fm/AQ0xz0SJzXhNFFFPp3
YenBIu6ST6xXlD9JLzE3nowki86kFxJ4hpGws3Nsm35HAAERmPqfqrpWNXEnV6Sf
brhJU5rWcfFLrlgMq5bP3CxImIiBvPMf2kdNuiedlKWjTt2XREliBatvmTbfho1H
h6VR+wzBhoXdIN9k4oh8/o2YnWX63WdurCb8UStR13p3cfb6Ljwt/0a3saLgsL2t
3NqBL6J6OKiCEjIHOqRmLZQj9omw99+nDNdUQrXc82kEfSUySwGaiWA+7CkJ4jh8
2BomoIQ8e23XNLiuXiVKsrHQ6FMCmkE19PxSb7qy5ryU9B+YsHvE+G3ztVApxCyD
iIBgVt6z0c5IsYRhJZZAaNJylMm+tWRsYN5bnnhAtFqq52hjDxrjBrGB6EC+aLhq
UBIjLmywoBQacSKZXke6sn50nWiQCpxA+r+zQBkzXf19vxKL2KcGN+sEWwte6PMo
kBTCaMr6xnd47Mv11PGeTKrxM1DfkutVptIRGNoWVPAzcZwQgveFS/LGVp8c30+W
JEoNzMFqIVm9wAKKRJOiFwT37gwyoqLV1yl4JQllzXk44BnxmDXxQOZYyaqQmhVB
01ogr3mV5BrahZQPc/bi6wD7B8crgkMRpvHGEgSHaFhZnLyF8KcyQcFh3pcx6Wav
uR0S4vjmoyfedzz7lteNIQEGj1e+lXJzWQ9tFW25qwyby5xIP60KA+rx0yBdCldE
UJmJVy5CSIiKzQqSsmEz810ugyPf4MWe5ep8SA2TCx8o9VR2DKUwe5amU3X7eP3+
EYxvRORWVjbVGUqntnFScl0/+cAefkhEnmAV3V3UUFsdgNUseWSn0uZ3q7Nr6z6I
2AcQFbhL5prPGtTLYDjbaUZXRbe2lh+OwTjcDu7gRODPPacukvtW9gw1ZagWOdRH
2yeWaUmFSp5ETM19VGCmUKLihEmZXpBJqa/3irVQ6TsURHIioQxRSgN5FsCFYsL6
cQ9jTUN9X6xgSi1fDwkmCI96wr6b0C1wHqqxB7a2I0M6o6XgCbmP591chLq7wMAJ
bAfRRu4ZKDTk8Jc+zWc0rG8yLWQmrUt+m3AOo5YAuObwXElU+IUaU00EDgbuBbjl
HMLumRifwMcdAMf/a495kFmNHUyhMP74k8a+4GUU+kTODED7ghzwQR6Pm3Pdv8Xe
UYKg/5VNRo3i5EoommOCrSnLWlCs6hzxwKKwdfOANO23oPTraf7c4JoEF1GyP6Hx
ffmDwK0ddYVlmAh0ZPZUNKp8Rtwf37uuZGhv53DR+1Y3Z3KjQIPwU0qtz9AQB2GD
V8m0euhVSzhD/4cScmNTa09A1BOKtrJH+SY+VXbV7MYLBiLBWCxUdsv4FeRZkLLI
2LV2V8/jiSAAR/HSkpaFKWb+++c/M8qo9FpsOenkiDyX0Zn0V/lcELsEZ+oV5go+
ro+PGly9nWdhNMutNYbnbSdym31QEFps0QFnMx4c3AMpbVwai50moqxitZn5rUaV
gTg/oLIIbnhXHeHwCA8V1+Sk6GmWc+ICUI9kQiUYORLU0qoXoUwLQKLlSsWQqAS3
FW0pxlQv+TLCmiUr/ofApBecxaHRikpZyU/BE+DUcWtmhIbOhocRNvTJoLxF7KNo
R/vb0RPXdu3yeG47KoJ4WnCh4jZB3agIuwa+ZTulKp4TfhzC6NN1hfsPqMPBPZHe
RN0NOxiqRbazeG4DHLM+pnabJIxWj0DBJJya3toBf2CYn+Sw4SuiFAF3WKdviijX
P/D3EmPXN+9jCk3/UYze8xQmnjuPIy2B5nzHNaRaR0SB35jGgfHKQnKu9D6BSBT1
CkWM0hPV3Ym1cLk+QB7HjQaC6fprHS+rc/1z50oxBHcI5/1vnZh1GberfBsVkFVt
2iR6B76Axs9l2mzO/fPNpbAgUhtFi6z7eNlF7ozpSRcqNTrGXHRzH4yCzlU9v8iM
UXzi/BGg/UGwsZUCqP478/pg3QBSymxlnWI/UPxHUyap1tp7deAZs+Zz7nhMyu3P
QB+Gp+xMYp5Voq7Ip9ERzeh6UGZPuIeGF3t2xWPYY7RUDrQVGLYeLyUlM+T+/8C5
87aVtI2qwyosO6AG3sYBZ9vFrggkCfmN+CH4GtDXrGbEDvUOjLJ3jejM6cb9PDmN
WpWTFMlrA53jV5ldmIsdqvsCPLNjXTdb2Voa43J15sLI9JgIO/0CQxAHvMjgfWBQ
2/NaQEBFji/eXEF5FEHaOrDqvwzya8xz9DoLrd7Bm21ZE1hbhEe4PW9UktT7LfmU
zxjNAP9vNwYdk3tGLErn8bq1Q8Z6FqSzvSRkmD+JOoaDmltlzPVQuYil6nZZtwJg
go0hg+C4qbn5tI+WsFCHxTBHJh6Ws7FWFQyiQaBowLyLXIj4wbP1Dd5XJH94tVQ1
dwDxdD1aCc3R+0MaX5+JLxsa7helA7xfXPar+sHPrZXsEMGPrudz/WpRg2rMYAH5
v5NHHKsMWjX4B7qCaIB+TCIfcNftSpN0OEWjD3sWSrFfRVkIfVYiHVoRf2FMuk2l
hJffvzGEraS8Bl8xi4LuCC87A/oAO2d6qZE7key1+FVKkdEjRQtFTolgalPKVBrZ
ZflErI4ffahkGu3toegsg58qBfiJNGrcbKrB0+6xLFSA/t8D+8up48zwoCCOU1xa
6Nk1rZ7xGaNd+oYnudaepRKBUWHa7x0UShkqwFpmXTsOm3TtsvHzswWglX03/4v6
NF8D69tnt38XWeXRpl7R5BA12yI3wH9uRB0u8KDA/ID2GztcfoUzc3O3KQl+q4dh
cUJk3kRdGJ+UHCfTs0kY/1vlgAKFOVvUoEM8iqa+0az8HYmspEP3dKJWUGOmmNd8
TgrNBRDT5M+YReb4KQxPi+VLhz+B0/znc+2eRAIT8B0ew2y+c6fJfmAqQe/qPGWA
6PHZGlsJ0HF5kDM4XEYPCrxrsj5FvXodLj1ooxibVNfJsuhJ51CjzNr8KUSz85GO
fiS8jVlCLiacbjeLTvvhInWO6Zv/IUw0ixC8SZc12Z/tp+u8aTMI0mrghdQTFsyw
gZHMR4vWRi4ztVbPaKO6HInnmy121hYnVd2pEYTm8tAOawVTVcqHjwq6IFQ8MB3t
8p+nbnaYoGGG7zjgGqRbMsIzXchX90zpmEtm5/TryYcqVNNWh8RwkCX2nnfDN2xr
b69XAy79qbsML2vofT+YxFEEH1Hz+DxTSOq1e+49del6h92M+KzkR5hbT17iFuHz
Kvxi84EFL26473TUBDT9f/u+WzBrTKYe2aBGdWvGhWGTPuXUrPbKf/jFvADVVf+L
9dcxQVM26/cGWlIhhsAu3dzKM+C8xJk5GRUBbDARBG74UJ7iw18ki9acQBUktK82
IDLVti1+xwBnvzB4p0avNlBQscZGNrSX9XszlishKwCROyKREaDDUGs95v0mNGCf
PfPjRPGqx4xxkEK4sIdWtqU9fhRzi90juGmZwtFkgA5XUtLKjvp2rzFamRNeyb6K
CM+lAilva+gO4maw/jOjObZf6JgfAkX6W8hFrZZDD6eQGYLTiUFBPTp5ofDOqvIt
LsXXaHA3cMZf4h1XlElhk2MqGsiSLWf0Mtz/G2fuf5jZyhUFk1uhm2MUVwnf7CXS
cdXot715AbOwRAYxY7EsCy7h5dqCixkq/ngq5F155FoPG3WQd7s5fFuMaBVd597+
YXPT7tdSdob5lNF/PTqv8Pc7E20nwkJHW5J6DLKeCXS3/3wE/ttAHNrZrIyu5a0P
STPSeNoXXPaKUba3ZpFjU2KxJ+c79/Y2p4k3upC8v8enJ8TWtghiJqAontjmR9oS
17UOzz1JM3awALc0ScknQCIzaJP36sLCu84lseSbL2MwzVvTH7ZxikNTc7ncaWCX
em3ZOyUrmjGg3M6Y1YgzM5RCIF+QACqDmhp6XCkXUYNudsRKY8Aydgrz7WgtZNV0
SPcwUcFpOzdEZjLnCpMgwNpsHTZLarTwjL9kE1DPjjthRCeHifEydz08BkAnY2Tv
bXJRlEyh9eGtxGvhtvvFS826YWLBPcNkXEnX4AN/RuvjaCO7BJCb87O179+TsIi0
SMOemEbUqCTeQF7m/fm82y4Ea5zqQLl1TFQLe5GYH4zdvn47UAS1Rlm05nBfQhfl
Am5bH7L1g40rWpvRyiv7rPIQf6b8rag9a+Epw3JV9gLlYeh6LDPaFmxRQ8ONchu8
2n3ek0FfRVoY6QAdV1Hnm9gqKEySWGDbbCzXSNhZMVqX3T6x7/qDK8Vy7oCjnX8K
OkfLEnDi4wZtqYTNKszpURA/zxJIU90bUj7r8PEq9XWZldZuc5cU3AWpEhtI7buC
MEy61E5kofFzNCAlP4AcQZYCq8fzYfD/n09XRe35bpRLe7dIxw7qGLTsJu1LB3qF
g8mrvSX9Lk/grN2QD5we6JswMd4Fn3zWxBSKyyNqFQk9QMabfrWitoIzX0eCFA7a
7396tryp6gNvF5vh1aA3l5tDncyVZKyfTjeFuIUzsNHi3pKY1OMKyTATziaXAevN
2bQrs0b1MVz3T/gGpKjwuSD4SToy7Rjjxv1NpeG9xemFkl9pNLu/CiSt5MfbxrOj
2LdvyaDD7BWY4gib2xSQ+aiyP8ijn8mlncN/PV2wk0Y3lq4XYa+5Wmvih4YBRfAJ
XocoYrly70Shpm/nNwfFfF7EYwYnMqGmp4TYYsIJMU+Q5UGMVGcvaTMtFDlFAiSE
JKcuKxTBY407f0MRFJgncAeknpOAbUcHqbjlWdcZVNKRPRCGVZYGUEwBdIMZiH/B
rjzgIy6uW4NG2P16477ectAsdb8qn6ARfYFWff9EKNJ9B90GOHazRITx+bY63PXd
iGfxzVJ2rvdSJaXRaJwRdkXHpg4tcy2WHhfXCkbsavjD4vVgzGghHh3Yn/gZo8EH
ATRl/59VzByvULRsfotzfxos72lH7tjJOzTXgeQgmBO/Cq+qAe+bhqQuMZLS91JK
x7pRJu4VgL6WM5FSjrQVoP17uWKpifFWR4xd4rwHXs2skerEBlIlf/5QZzY+bL8A
cyeFpGhI/EHXgigK+nPPCaQG5mqYs/JsbkF782cKONJn/4ObCOM25Q4J2qz3I7zK
gz+n7xt+3rC9EdEGRNgIKbnkKwF4kldJ+UeLJV8rpXYyrWAD79AXSv+qcf6bbSV8
PIIxF56wY2Gp37jMVNJ9CxoHTCjMMmM3mZoBJq54Jkyt86kyXMkqyBVR7pCQodOX
ZzboIExMraYNZ0Z/2sZfXJ56VJVt3ZpCEQ/quWs0k3Gz9G3XlQ2X8o4xFdQpZ6z0
PbothVKiECGback9wuUCXzJ1NHkNFTuSd5HqlAXEZmPJJXDNQyqkcAkZtxIYkizl
0cMpcHtl3RjMtuJ7uc5nJ2RfUq/BTarvsoL0bq80YIaq+nZIuTF4GRVeDR0sKq8f
tBgHSKQsMbYQ4xMdAC9//fLc2Gu4AoqZGTvFK1jHDG7sJQpP52B1qhKOIDwxZ5Xn
qRZUo3vOsorOCduJQCBQpYOWnmDeN5PdHLbRn4v0/gnf/mvCa9nuxuV8oKYHCX5E
6dW8v2MVL3h/e+ZDLXkRrikEoURCcY+VwJSEbXB7CIzlnNBe8cTDXnSEbr3I5rpn
oYoz1vX267WXDKnJQf+JgQp0YiZhClTbtqoWUS/HikJOWcBP1y1Oq1WARZUcnFrA
GvHEIQPEkC7WLctGvcsetdto5nvqgUuQHilMXg0AurqNGYYvSmZQetqKXgMNU3oZ
Odg/F2cKXdlQ3N9OBcrrS2EGMgarDJUQbfTwLaM9Ybq57FkDC1VMGzlDFn6ffsyG
LCryko4BUj0E+S3BgOkoHnh0kebenp9S0GT1hjfkwQuD7W19fKHbXPFjO3jTbTRw
21zVHh4Ln2+t7VO06/kzqAEyba0PaxqCJmduMeYaTxmsohZK8lm0ik+v+xq/I57c
2ZcfpJcTjihX7Y/coqvU70ULCg0SW2t6U8icI9t4z+BADdEQlcN5fv0hafnHyBTF
d2eUocS3FjiYVS4puICexIkHuiRcXqsy9yi2yzOnNz8q+n7HKB7jN1AcDTNxLusi
lr8YSrIXNzMBR/F6aR5Fot1g29OhUXx9rNkjzU9aXSoz7aYvAau9hyAXkXZ1sKz5
61ZE7kRqvXcadRGNYe+t/PJrciOpI1xs++JI3xC7wzxVSZzuBKXiZ7d0DvOgnfQk
3ookii1h2Hy5AZXPmKCxOkUZAbjF8J069WZbvbkhS+46TR+sv6mIkuOp1a+x+9r8
Lp/bTj+U+6jjZ1FCOkR2AvQU8cFVHHEKOUYSLUmejsPTA+gbHOwNXeR1BDvnUxhg
5QDfdv4CBO1U4ckvYEzx4nzCesyb7zYOkkfeJMKEzT6lLtKsHUYv0A6ZGTd+HTXy
rlwm7rtrvRcHD6ZdLSg8UDYwfVe3YQ4JwFwV/puifM0KAGGkfufCBBmH5Sf/FD+l
16HTnoZCsxOW65/GB/+ktfmfK7XNqTYk+crua55t6O1YExL6iHxIxNccM6AOYv0c
uNBS9YbJMuKWCTEXMxsdOce43LQsNnOlzeHanY8IVWW5r9n40KzZG/Q2VxgcqDLe
GKVIHV7lw9tYeAzgc24PIkpIo1cRb8NPusEb09uo69LIVv1rfHTX1iyezosq69OG
mjHn13+eDX0hILDUWTesUIi4r4q7aOU7RXNDJZ5WETqG4U9A33H4Gh26tU2iSGXi
JynW9rUKIci803iJudnCDjPPItoDKhcAJ25Zb+tAPXPbnMz0BdyEDHUAh/JuGMdC
kXSflx+9EdVOrv1eOnFudyiGisnadQI0p30udVFbPynFFyCoFSVj9wJCfJOjy+/B
c9h673ycvuuZ6E4bVSx8cdIW82O+pgcsNCrfnc3sjYodyD5IKLsKtSkuAnc1Imva
AQPKChAuR6fUwV6rEODWtJW4EqotWCgyA/nZg1n78WJuMnUjno8vrYZVS4XNFT4o
KCVgTio3PmUuSYi1SnJPLWMXa+RFHp49n/GpEFaQigXhW2vAdX0tkAtovpb7mU2k
ZFemwwa1GPYVvbtM/ZOQKu75lpqXe3F888HKtffkqucWOP7KZ0byJCdYQx2PGH/4
40gO2GJCCEXAmVnWzrGHVVpiSwoMBIKnGz7PbYwn5/tM+j2ZUuoXqLxSVFJfqWez
iyneLwYLs+UxC+6O4+G735ow7Cc0PTJd/E+5OgkbPEAVOPzAt+C42dNNIMD/+//c
uIaO3GsSI/PRbilnm6htv3HER5uxU+FVTfPrJpOKhYH2kMUip8jGEyG6kxbsLjfs
1+w8w7O6p1T8nkwKbO60YP/TRCM5a3UAZ1EhETuqAF4jNCSHiOPIb8gKejNX/2SN
W3VE7oepPA59+qeOopb/cPzszW5bclXYZUwPzhMnYiHTwDd/JEKUV7eQXNH+oVU8
mP4dXtBamnrblEzcsVWc9Kt92Ffte8S+JuUr0uIgm8TaNAyr/1jGaBnZbLg+amli
ekz/kKdpTuQ2dOo2I94xYzKCMP+w8o0Sw2RpBWcZnO9vwQNhlO2DoTtLls227i6N
47v+BChz5uF7nQAuKaVtle61p2dF8rLFThLflLlv/AyMHs8/GMdWbc87TtY0BXGi
CC1cUqvJfnNx2s0oYxnTwMesY4/HOJeEY+kkFD6bR8ZdduftoYSkKI+KNMvAGDEp
1cZO562aeXm4NgDGml8N1P0L+EwvX6R74e0t234GgFnufOUXzBcZs8CHCDWlJFOk
cDtuiHL4ukvP4xl2TKRDFRZzIoi5EarUEk8ZsWq63blE9QpmpobXm9Mj5zQdIHWz
dAbiT7dBGGsvSlo1291kj050+gIOxj0Z3O0Uf9Y/h5crP7mM4vM7Az/w5UAqSXRv
sOpbSIW4rPOHQwJ5GuAG8onZXAhdiahv8/hxRJ8akJI3Zb89pQUUbWyZKa5CKsdE
koup+d+C2nsU+mRO7+6UpWW9lQZidzz4JrrFdLBRVDk427tqEH+pNEtxd6v+G5hZ
oCQMEi/bzg0ggWqGK2q7YtufNdFnLynfQIOBdP0LStN54mIOJJp3GMtcri41/ODT
if/poP75RviN2cBG73/Oc1+WjmCKpfp0xhJHwiRT5tmxPLLoXE54/wb6DXVnBR8a
IZpJP5knlwNvtKN8iDTOnIamANAipeO7ArP9c/X8lhSvT2tGQUeakqj5XmZXfWWn
4NXT1i/Hr0QCD8CJ2U7wBnBWDHoHCxOPXWjHQhYylN+grpLYdsav9T+cDcNSpVZ/
OVqqBN1EFwchMoKjvshMaZq8Rb5PSnz/aqSjf5HGTeSZjFQmQtp4XNe0gbnbILtE
GJ5W4qinl78grQVvRVQ/38A4YFz5ql9V5Vc6UDmPHA460OrC+ekTx2jZy3nKyodx
3xM/ng76QKv0cQeuV9jjDrJD5ZVsrSSNm9dvhTVRL2UKyrMxtXa7HEtazbT6gv0j
8dH73a/CDqZynR/PR3yb2TyO05laoC68ES7lL+opqWTLO1+X2AZVb45a+5Sli5Ey
HA/FOlCVmzGnclE3EAM4+fXCKfxsUV+vqfQ80Ioa2aS849cPdgFTy4QAvAXNeiec
R8sopXmB62DJZ7DUBxQlL6HHbcCZC9pmpIvvgk0cJAwBIDxk6NPr5CMKEQvMDnPC
aJ8CbIK469STEpYAkdvBW+TIFtaH0UaGU/uMXvKZfHH5WPYNLhX4HLKcdfIKRMne
5f1d7UxfpwwUjqSQ9MU/ZJSOvSPL8O2hmXJv++Y/ydXSae/gtdCecPeCjiZ6dyUg
WsJsqtZGE6KVaj0eehxbKvxYAfebzdfeRS4TqkhgZtXASh1aSAsW+v3mJXp1xRZ+
yMG1jRKkbsD+WYWFpalEhb46rdWD92VJ91JDNHuuyKy3DQt+fqX7X/t2yodtZE9T
5JvhTi6imkoUBLgMC7zA5RevM2q74jp32YKEpseZwH4UkPwqtdhNA+t5bgVlJkPy
KZeJ+amTo8SAMZKmqItTOhNZiSGxhqrpyH5IUarSoh/1Lm7k4PKqZOw/8otwfQyA
XK36kXnzLCGOEapcLlL7Vv6SAL5uuu7OEr2d6V27PwAOz2A6kVhqBjaEeDfF3e4w
NIroU/1/NWUM1yIY9MWfVG5Jd0ZUo7GV6z32mxcnrNAalb/MEq6iXUaQAQBxpabL
djQCY178uyvc1aLscPKPLlmAD4YCzshKdsTjuLVzRyMY5Av8BmU60dUzdlEfTmuX
9085PKuFID0gMSzpkHaFegovuY438xjCgoj01rQ1FMF9t5SdXqnulmNzm3wSbwxm
d0Ens3Ug5Hu7befuDxHdEZxVPJaLHw8OAHktvkeIiPQhI2rvHx+P3mod4ACx6qn1
YpKU4QU+Xqg89baj4SYMa7SskV2UWATazdkk+QWmeaxCB5T2L2XWqFadw0lxl2dg
S9YS+sktQVi8OZ0VJq3Cmz+/iC2/xD0gbIu6w2YLagtDS4Bi2xgzSHGslp1DYpQ4
i+PnIeZlxMZmxbmr5+LHe/NXiR5wvk+ZT9aRPGDiSyui3xfaYn/ik67nmXcvabDp
jNjOguSki7XxWDDFRTKVhDFiWdWHnV4GVtfB2rkWbEy7bsYM/xZaRBrN5L6ZPcv7
CVhVK8zIC0eMHHXJobZGu9Al6OEdoeRQsop1NcNzbR7QlxIu0rCHiUpLMSnyDN/s
0VRSskQIInwj3Mc8Bb+sjszt+vtEO1pw0P0WS5Mer7GieoGyLyJzd1T0xJomDH9T
KQk/H2s/O/imF82OmIMb1A9bJ5U6/B0O7MFI9Ir2JyPj6XRzZjPFnLWNoy2F1jgE
EawtvZJo2Fkse7VntqrQePeMl3GbTClcEkyiNZuBEr7C6dY3hm2LALGnCBf89eH6
er3QfEDnJA71RUi9/gq5kQDDdEnioDaO5SyEZPwvh4ox8RORG8vnvG8ATmM85r3F
s5oSTdI0738QggVFEBMdjBCnOFOfQ6kwX6B0HQMuZLEKxpWfLfXk5zHdFULSGimS
MGfkUH1xkPGgpbDD0ijQGhguWs+dRqn4BVpJb7F0dGmFrOMYXqUdd/GnNIeDrkrS
vMPTf3NszxedOEv9OHWu0l6YN8p95xMhQlHs5AfPQFpLDF//3DSN32SYyPI91kep
WfYkJdpXq9J9A/Y6NYiQzXLpe7wr1ZXiXzisbQEWqvIacbGSHFsa1e5+imCYuP3F
/+8ZyAxNzvnRIm9SpGRvNO6qm/WPbMJlwrvJ1noUPg+NNon22QlhsItu5uBEK1mb
z68wwh6zhQN6TgrukA6zk0KPivRCO8qajTgXnb/pxTsNjuhEoZCqVZVuWwG2i4Zh
NY3jddJCu85KBzXFb1FyXvQdlCX2x/u1ZqIbBIBIZJR2chGO+dZOcexrRceXFUMi
/EBMcgHdjsqS8Qhgm5paeB9lcD3RA1Pc9pK176V5bv/ki5oKoVO4kcSyNZrIV+6G
RVMl6FGJv+A7QVvmkdOYafDWzAG/P/GWN/L3tMwL7d+523VHK8SKhvWFrxnrUlvc
+e4QFwIz8YRjaa1++KcwNmstLL5N6mE6CGQMkGcmdBfnt++PlS10B51kNv6+hekl
BbPwLuajGHFkTsTWOxaU4zyUOfq89mLevjL0YvDfWLxRkLCSFSKRUQkWf7tcGhmh
ljNIAXQn+MRsx/Ks3BBhnBIgc/p4U53RKcegV0HbYE7B2Myvy1NUpVJ73T9v1htL
YlDlOWAti4qPLNAC3RPWaV2JNPe5tTSBH3XMAjlP3Ifss+VMf7pWbFHmpPRdK1UK
/tlMt/U4tujVfpsq+vT3nuT51VHK8y3cHjXsiuxysfvn8EGxzlkgEzUiBDawMHsX
DS40yr51oei47nDKKvt+IfIWPw+U3obrengaRCbageL51kayJo+2ubVL+75Gvjxr
uOn3q/cw+Z6WhiXCcOs4HTQy5VzpllHIzXAq5K+Ou9xK1ea71m5bl03TFMIQccgp
GgRcEsaJLxwAHyekAn0CqJ47F3b83mjkJs/jTfu15q/HzFAgiOiBM+NaKwrz+rWF
BVXuix950Lt41n/3QCGe75xYdgonrKEyFz94ZeRX9U93m9GNVjj1TaNPmxBhuBlQ
Micq85bb1cM8rv0uDPCZpRBqaaLlbNMbDB5F/+oI4BF6/1l1hoqVrU3JAKgKrO+F
8XXyr7NjKDa4254tyxKBRmwSS2Gtx6vrEDqu91wmoAny5uJTk5JcwnXF38fHtghb
OQ5GP/RmHSqL14g3N6Js8EQmY0TjqpgQpJu3mPF3LUdZGH/QlXcVUlGDawn85YEr
vFYfIveVIJaQXD64ObR59bUQiRkIk/08a5Ha/MGpGUfSWUFTw7u9Q5LFKfGxWAgi
DhT7zvaefehrvBjnwQjtu98D1BWRb/9TqsoZ2DM6rY8xgQYKTKR6lQXY4jOoSfzz
NeTQFypv+c+krKfro0qlutA86jNUdwU0wdXlQHZJManOwCsm3Mh91r2Q3578keg7
KLn5UWhrX+Rp/HKR73i5RCrQ6ymPOYMKiRrvdmPYZTERCma0SpqFHqBLJhEqtuqy
+bc1UN+cd64PqTSDX13osKF2zem20UDF2aOjmQUccAFLc2Af5GMUOKYm5erXtL/K
abCb3mjh2pPro0dt28aZLoCCTei4yBrJe+MmdSFtYUzoLXVWMFJW69NgUO0sqWEX
gnPL7WjAK0yYI0Mg4MoH9a6EfHLSeeA0p+0CgbpifTtRp/nQINF6Niecl9Aj+K2f
mRTK4zQNYR620hWo65UA3RX9v6Fa3eqh4Kf93jf6jXW9akODBDREFn+V0TU1w5ni
xwKB8p6Agqa8WlSya1eMPeUioF8yZ7cqywVIWv/4xOOR70FSjesk+BM3xR4SlCMn
e42ZwDbhh0OY/PYFPHJCHGkK39zQdVnAmIEGXJQm6guPueHAM+PomQ+avmfXbe0H
dbvO4byiXkZHaI/GfBvDrnDol8yFHMU36CaWd9fnspXKJkDQ6uyF8nqP6BbGobWj
bYnHPSlk9EasAOTN5Yom3bEf0MGu3mPXpk+2OP5ren/SU0WMR70vQSHJoBrSLrNV
X5ky1rYp/LI1guRSFBexvT9ClnBmjiRtDy04korq8LgEjZ3dH+yIzVHwVXUQhh2m
dlM+AwT83jPxbktKj0uNUjS/HZk4FAWBRShxfRNtJ1ArHvT7jnNhnZ9m7k2ndQiG
NPGnj6fgT5LWjT9sd2LOOc67EHcj4MC6wrXg8lDqvrr+5SISL3HaLxaCCbTzZBk1
xdbK7uf9sD9xX0TmCMa279u63CV3WHcMEeNrFQWnaewyCmhKGMErPh3e9BPotyI0
fdyhC6sfQ04GnbzlXJN1LUQcDhbh38b7H5O0ovLFFqWmVIepqUrEiBmWXcp4uxAg
RbLvUWTeJ/fcA3XgDqxplUwyQbDe6yNdcSYzKzy94737zk3gfIGrZrKICUYy9aRS
Sb2j01JzWWrfJ7M4l6fBTPVQIPu7f7vTpwVtXaaZgDj2Xi44mUAkOQ3NpAzhoN2j
nkmF1ST5D5vg3hxelyTW324Q5bi9IcX4liV3L/XInCXRAt1Kg3gAWm2F4892pj1k
HSKY1LjFgjkzsNbwqRU7LrRLq+EMyKBLDMj8GppRGLXCkKu02/pnEYS7cvpcWmZ9
UwRmfjZzRVjTPv/os21vTRmIVGXFqNwLPQW6G1qQWtXuXQ8YGP9DeEPGUzSSRMru
D2RphdU2CTJkNT2b2gzv/nr7gRW7xeVzZBM4GIxfyMjRm8+Muuj/vf//etmP8Muu
8pEMmIon7jn7zU9lup5cbBvOFRGER4WMafYFQ/Uj2Sc2octGTWPkLe0w0XwFQ1uz
+rMVmnODHyWcobSoIhW6mEXgctY/LR2TnEaRQXqSb7QyvWZm84XMTRhRPgx7Rhcx
Bg97FM1Do/ZN+PF2f0ZOGfWsXTxrsil4I6XZVCMZz04Pxifv1yNBNIQpdxVWaFFY
bapCasTU8yQTfwuLqVULwu6LfYFKaxUOdbclfFw6n2G/6Y7/i5RlB2CKljIea0ey
9dd16mU4VkDxtjfn5RQc7TvBuHWP1x7D6A0eTdRzwmHBxkaHBEYVliaM4WaL6xTM
0hVWYUshuwkal5e0lCxtUvLvdcwa6yBCKIMYMm9bJi96/Hw/F3rsojTdu8DClXa4
NesefrcaeQm+LH3l5t+yFfxxVwsqcEeWZ8wxtYZa6geQVGKvsV6D6uqhxpHUuesm
pGkMscENkU+wTbuLaULmdC1K3QrfRkSEkFJFpmHH1M8U4aYXg+h4N74/UT+oklY4
r4eeIBYnw7pkt59C+kMFy2dHh3gOorfeNn+ujPs9PVN392L9tKFBPWTNo8ysakVY
mtcgay+sDXCF5pa12iv3EOHLLwmm91L9hMmH4KM9tOt8Frn2QvSWaJ0F7zy9mBPX
ZQGEa7wlyGkUWrRPY791aMbzely9WVR4ICpYi0uSvHYS2EB8j0/sm6f2aA4TQYU/
ijmzYwESkq+rsPNLRlqb1Z46q1HYBAtXmx+i3lk7Kk0nlLuYfSvdyF8T+UCHjPgD
iHDXUddhUGq38YkjoSmLQq2ceaDRWaN/c0QOTX1uBQcXwdpmNdkHpGhH2NuNt+Xl
4Y+VxKtir+lT3z2nlY9X17xV1Z0OJHFgNu3kOm7pTCxHUf1aj2yIu8IHPxbkLR7k
6WdLKRHR2pIEvVYL7HftoxQPl/Vef1qCgrvNqbzXrJY+y62e8iZ2bQ3WkiNHiNTo
xiGbTowEOnSkVM0S1FWxdk10Q41kVV6t2X7zxfmi0vbmb6i1U9YSXDuuvzmylyuP
wfk54DNeivjs/xHHpnS8KcAcLtUMq4fUqop3O+Sdsj/JGIM+dqehf9T1E7JuxCPz
joBzo0rYoPH+8teSpXMSpkeeJaVGKrX6+4+86PT0CLJ1+w95z0g/I3mXfBp9Jcrs
4vhTivwW0qYdv3D2QvXqENz1d5iJwcxWA4RqRIfl2B9mWVfKvpc7ql+mexedKq+a
94lBNdXqR5M5zFjmiVjKf5ekFdFxWthzDJFe1VCkP2pPSGYFF7CcowDoCjys1rhT
5rhXGDoJzS0Mp3bRGzg2cXqlGRmDTNgHKRIJEolxdppZ3Ahqpc4wAw4TWsZFQfQC
k50ky1Ze9V9cdPUlRv437pujjFSZS4BOQ8rF1ZwQllHYIkLZWCI6rPXOCozhl5dM
WwTb9Uwrc5gA4tSuNsNmw7zDaNtyYL2j3/p3EgiJBHRmbN4X00tqPz63Kx1aFPaW
ly1SU1HL70qwAn517pi+7UfWAjSLQiZ+3WTtvcnVWSu92o+MHJeMuyTrz8LSAPsE
EXd/+klgDa4gcECrTuAHJESEaGe7Meqy0ahw+LehLoRvskWi7CLp5uKJRX25EbVz
LvrNCwyQndSRfiaN5QCW05sik2gC8oGcGU/951dMD8S3AcZj7xDwr9TZ28pFUSwu
g/hCmHHzcsuEVXIngL2Vie1TlqhbFMMJkhkPN0R9pci7KVE0WUKUIPanzQ0v0ILn
38y2DyJmzRjgHyCODPJ/AZ4PEBYevYfi/sUg+I0XfrgRMCC5rP04hH1XWuLAOpJM
yxdn2s4lppBGoWDVVsQjZU2Xmh0+8WVY9C9f6lf49e2fcf52YgVdaNYCL4Q/ILON
QLGFX3tKBcKFyPcn9BXujnraT89qU6G0Oe84M3xW7Xz2afQvTmRain1DbuMyRHC1
ie27+wFNNeP7CBABD4+7h0S/jKlVifR5QcbHZCxTjOnYeAaEuQAsVx3AoCzNpZfD
/aKyxah9IRMavR+1pRo/Vw9nCDmFgK3FBXV/BTN76QgK/5tPKGGhCEbmFtXblqPQ
xiZauLcZFRi9nvQc7CU3eB7jMvvbJPgD+7/YZgJYxHiNmvgphdSNi3ejetThIZZB
kJ4G23dP/oKwrl49sWw0UT4CwXpUQzymPPOXafkvKhyDBHc8+DN9j2MpaH8CKEog
5rN9oEH3n5Z8UlGUQHoGvfx/b4VoWwMkC9bpDGjocFRihmtT0OfwYYKpyBr5KM5V
ymYcwkIfCCRzA2jNtC4hvQjJeUv0Z0TVv0bRXicjbrGgklojhDc3/6O0ugDzCiWQ
aPIyxIk1LX9WV2ZTTIG+yKlVB02HozQtUtLJUhhbm9BH6A4b+KcEfS/ziVh2C72K
WEU0qDfpVpoO5be8empqzuX/CYVjxOEdJbAWIC+UCqMwenTvhfWPVKhFofXvUfqy
hsLSXYaAdsbqe0KwtBSew4UdZ5IRDGdqaecOPTeu2EQ/bYonVsSQB7b1ugN3JZ+Q
1FzR4Mnpihecw9j+mxjwK+GsGxE/uPlYfN6h80TxI/xST/tgKTMbxm1johac2SYQ
m0G44d3UMdZMeSTg/glh3GIx8Mcm8TVBdjlkRRbLPJ8bkIwXuYYDB/LcY2Az/RtO
jh86sQhDGt0VbtJ4zDbY5JgirnrF62HBcVJ6vp+qa9yxtrGr1azYbeOM4mfwHYfr
HlMFu6ERMb/CW7giN4IRqTwcPjBQ751DEPJlxY8wBbKeJHnNLAOmSqJDHr2fzZoz
ahCqpvsK00KCaN9nTEMjkZJtEKxQdoMmnYnh1bT9AohU8YBNoHGbDm/N9ys2p+Ib
zqLftYWUW1lMQCwe4BJaNTML5Q52CsFsMN9T9913EyAsqrNejZdp9QnoejPt9lZo
M+QNr0eV+deK5uIJgwm2h6KWq5C+rBwWJWeHVpYy6kDZuHRgHvR1BB5+OYQrsWzE
xNKix39KMj88mZjorXmCTeEn8F5ut4iq+4uxgrrPJnEU9azTH/KGrVT5ZO8jJwdO
vXsL0g50Dz1fAAbbOfNj8zMiayrSIlgMYDG36m0Lj269C4PA+ptMDsziZHK2fXz0
00fOGaUQlCbeWfnYH34wXOYnc3Uua1J1Xv/l+9g+mLoPprs/0DjIJ4bEGFK7OACW
n2iicpI3bMpxvhcCbCfXUfUzqDka6zr1RcWFpreZPW8z8mvKTLMypGp9wuQi270v
RYPFp5bTh+GmZZQk6SaQVTz7GIii9h1sdHG6A+vYs7FMUzMO4/GxbWs2fKd7y0Im
pkU256nV12jgwThenz3LQ83D0uWuXtbpbEIR1AlMSKuEfq1vp6fq/0xhOKln8h6f
lfE4m5qnEJn+5G1/mCGOeFleR5MEHfU2jVRFkISA4NSQyZXsrL2bZ0fl2UQFtju9
XXB/qlEYhfXZMfMeSl3c+SL63S99HW8X3hzNJqr5G5Levr4zjb2gnpXBrj/M8+oI
mHJA6Rm0X8qQOw8n60v1OY7YWITQEArOlzyTfxPoN7rS+kNoUL4sN0Qv6j0U4HoO
M2WClXOnNwZIDJ0WTzcHYAOFUlPVDEDoEqCWnHRf9hmTwE553816QLiXMLM5ac8E
q5LqCWOM3aPJaphuTxrFadocNKgvtQoqm5ubQ4hQB+WZK3H6xm0GdzzkOwmOSqI8
Rs6UjWubzYmbGj4Q8Qt8GGpAqCQY+MZR7wGDXHte+OawyjvHJ2uvNZAN+6FuatL5
LlSxjjtVGHaGqK6z8BG9YjWoWuG5d6vgsjB16EsrYqoHExvJCt8rX0AirR3cc1ec
2UAgI5U9l+7Y9pa45YvgF4+8TO1hDsYJk+ds8L/zsRprzvpdC2ojTRLAUgYxGywP
jDeRexb84FhTuIa9otP4LQMUVA1ffoVTHOeh4vgPzcIdJ+y2LNvkIfBM62Etyc/y
Xz/99nAZyT8qXVyyljuFYRZiuX1uY843nPm8bTz0te+2Vt0v68VdEdNrJ5JPrJLi
SfK5UFHvbz4m14KzRXmUOztoYb3CoCCcDy2lvwbKYwOjy5dw4VkytNhMIwVsOlJn
u2K8pxGaBRGJjMgMwwKsJCIPrhYQCiCTHibksH0fVHEtU/M5ap0TSUeRukRe4fEA
aoFzG0F0Bigo/6EYYGpFhOWwFnibb9fm1jBMEgubSAwIAk1nvCp4HweDEqfdJga6
4oIyC9aKCW8MC2HAUnkP3NcCo6S+FVNnGjuidI8Nj7coNkmiV+cilWFi/Srj0/S3
aY59z93yj20ZmKAktmz4GjEjDLWE5qruyCsDlG5pLDZbcu9qeJ8mBxL4UZHgHsh2
Af7l/3dgKa2fbXbsVCH7221krdlhBx/ONBNd+vuMdYmTxRWZFEc2hr3EKmzCJ1nI
mtfG1/NV5CQopko124lwhVo7RwGgp4/9fxDGfp3ZbHpZAuKuglEf210jzcmGbvCU
A9hv+4yOO0DLU6zpjLy8x9+8naIUaZY/Ozp3UBX3JyxA8UoDlZbM3UJY89Dxt2tW
8FBNlOfOEZ8qjc26IkqfQnXNNFvuXf2GywdjIaCQnE2xajOA0SiP82E6dj3i3lf3
18D/k9i1iuefesKNWDC6vLb3lbcN370IdSm/atof5bTNTGKqBFdAIReYDEvqBBoq
8qeDtO7PSneV++2E5zaZuQBDqAG/v9+s1nTl1j0nrOOLSH7ARBR+j2koFD3sxo+X
nt8UtCF3H7SMbrrH+XaKjWzaw0/wTafcZVaWsPTLfnVhXTSJDxunOSZXdjeXacJ9
4aBHZJM9/OUiXsUGY7bwXxhVpywpcZAu3wPL7H89eE0u0TXA892Dl9fcNGrdK1N6
xN/1X2dE5J3Dq9vpD33e2IqFOP05mF5oeneKb5VdRazr6qCl7k1AwdDNqGKGpcSe
wtfHYZu7bVhI3jbx82XUBTJ4UvQ7b7bzJU3/Ek6+3CqM/6nZ5gFK/zEJum+o0ybR
1d+uZ20a9veYGKE3nxYW+hYSSlnRXyerJqtSvpkA5YK/A04Th9/Drfmbp/sZHM5T
YcMnlOHfTsw/bF7/yByhekJKkJQsVBjlLpK3vc9H+l3vcngKzu4r/76Mkoo965m9
ZQPDC1f0WPxde8dhaSzkQAOChwbEs2OZGxe4uk9xfNrs4cjXcQ34aYW0zlr9sg8g
V7jirVXTlDx+LK1IamR7qoeButaag7TS7XniYWh2AeS7M1ZZaEVHBB2nphBa4eEA
lMRwWPlxNCerSJtbCyg2a2JFjlNt1JDMAOGSjx+RO/JLrKf7PfoowExvETt1ApR8
dWxwDDwXmA5Q8o5bywNGfeNcNn79NIXq4qqnhQtZlRlxGdEiWoCaqgwIs2OUB/Pb
qyrgw5dNZGrwUozv5Y2G4U/UGKSEwhcfEGmeqo6x34vw4+Z/gQ3bIeFuaVuI1q2M
2PDaRw6mQJy8Pzr/rHwxjNmgF0SPrMNksPSWYiwaxX7v1SeZDlrRPJEnAXu8nyuW
4S0hpAEAV7lfscM7Qp6DGYXT5i2S0qJwGia++3mKLf6gwmxbDJbR/3VHRruSHPA0
K6gWT2qmvmRF64eV2QSbVgm3ZxZgTP395TicF7bQ9vtC5/lrZJgcE9bC8jGqK0ds
PplO7eTlydidk8TTl7ZvU2u9GaZdG8Ohy5HJaTGISLKn83d9G+FQ/VzTnzZ5fndw
b6cLoy5cQlSd6gobqlau+T8pr21kjSK3K969O5kPgThluFIzR5W8+yC0xhKPKcVU
jnlmQtmxsWCP1QFEN2Wtwzq8ZknLKIw7xtqPiE8lNft83lnEmLiddpSOwlvqav2x
Fzzv0Uxq3vh224IBb16Mdl92rtwkyoh9NoiR5XE9sFGYJhDFLyMglkOobi8Dkkal
OGdkJp/Q3VSt0Jq0uVNujj32sIANUB9Cns+c2d3Q0a1ky5YMdJAxV25k+asoVSRS
AmPoT5vp6yJxNtI7ZyGw70u5M1y2qxdkHFvwRMStHNzrYp4juIx7/ebFVhB0Jczo
H1Lh3aqUGj+60C9o0huUAE7apzhGxi/nJ3+r+DsdCVdSzaqpmtl4R+ZNcFLKBfKZ
U5mAqprfEUm+57qUKLoCfyb0tFD0hij21Yi8MizHBrHagNFnsIt++KGqZIKfbywm
PL8QM53E967KSMflwOk/1O/Q+f5uEwSe4qX0dOwCq9A4aSjEpoNqd8Pkn/TJGPGi
iMCK1XcrLznbAgmflBntbN/YyyLXy20G0/0twNelUTBN1NKRRf87GkmcA2ihYxwR
BhdSzkPNSQ8R1PT9mxppyBkygCllGpRSPcSKHzXMWMLZFXutPU+em1Q8OhPWNeB+
fdIEPf0fY01Dg86LmXj8XGYMGzCQpNmyP0HVgjQKZnZzpxD4qf4jybLDa86uir4M
x/00Ifk7ajzEDO5hAnPWIffmXef+LPEygEHvI8rht7U7i2WF45vmssc6zYYQ3gtj
BLyBc1AcKMZ/JmGakexIWDROEaag8MSbZlUGSVQiOkVkl6eynnizoJdZMMpntNeU
8t/Lb8PoR+JdUGzaHDNjuxecrl1Kt7UGmjdKjhS9MlNpE1XYtfLG93MrBTrXGdHy
jaq3anCzjM58zbZ5/reT7SmnAK8S8yT7Z9y/GJ0YeymdYluVoZpS3Qe53nMMy3Og
vnfz9dJHsajw6/bLlzuCSQSHaFN7AzcnJe216lGTvAtYKY6h+jgxyhpqg5FnIYtm
7WTOfmImewLVzDt1KPDht3Rf9i3NsnN38K1voTkKs9fJdEL3o+CUAHKjisL2OhYB
EtKHMT2gwIWxYQwscGBqhj2xKajA8TLAw3CEKjkxYfRBcg+NjCrOZ9gdkHgtBmHK
Z6O930g2cPsOaaurlMEdGvd3UQWyJPlOhRvikiklJjFUzqVRgg707nyl+1lnulxf
KTbA/M7uCX0VpBx/t4/D/ApCjoUO3mzxPom/b3vIO2d08556Oh10OT8hlVLjs9NU
alAsFO5PLAiHExdw1jl0y1HEArLqD3raLU/cNCn7gDKLJwvpRRXtt5ecxTeWXbUh
PhOTx9fIIqOIwFTFoyuqW78YWMsommTOb2j0+F6vEJgK1219KBOhdD7W+1eNE6mf
sk2ySfa76/qRaoDeNU67G2IC+wKZREINszkiYX5Q2usP3Of48BePJloyYal8jtZA
tLT1uCY+Oi6uj5DZm8YlB8oGmI8XQFWpTbE5uW1CbFYcUEHkww97i1b8B+Oq1hox
dJi1UfkTzsrAKr1+fZE8qlWxyVFduPiaVGeFVYuyTJfEz0ZpUrgnMS7cyVNoy/5Q
3cZY1EZMFg8J86UN5RTUkyHm02oTC5aslFE4emz1ks/7ctPRyv89cEe7bWeCpRLt
ASnMKvW+hZL96x2GwYvPILfcwEHi0cbErXwjFkf4/mLntB+jnrh+GpPLZ27Ly88d
gy8EjaAu0mUx9EnFYUbXLyyktJVy92gO17I8n9sK/DTgwLlSEnZGnx1Ue59fJBFz
GqRADf8IP48APDFijJA4p5L3T79c3GYKxlsNf7dTQRaFwc07NV1H68jGIadRaaTW
CxWHwaCfHrULJFFXnRllEFvtiPxEAU+INvUDMkujV2ORk4N/eKYF9FJms6dZAG/7
z0+xQZJkFDL/muPiOcuoc5kYNH/AfYw9d8Tv3LVEbfSw+wbLbUujhKYjRElZK0bk
X4PsShAXKpurg+Pxn5fkgS+dlafb/PKhXNsJlJ7y/U3bRkiZJxy+jsOatGsYfc3M
2b+oIExo/MTrXNvj4IUdvTgzsAeiYsfdT1AdxORh8R7HpMdC6/4dy4fcJ1cy447m
jodxDxb0r67dvJSHJHLpIusFd9mysc90wmLMxNk43zGjaJbeLQZbbrOu8J19z7vE
P3JIEwWz8z5h3eK20Rj+QK4ytl2KwOqV7InCr5ox011BBSlddyTH5egK2ght/XdY
qcI7S7GivQmUceWorEyhXvGFvwPY7K2bE+l6jy/qSAuHioHptOATrYhvrxQs24e1
yYkUtWI8wKkibZSfMaaOHQ3Mm1MIyTng347dBa83LV0Q37QXxVn6IYLBvBMBfe5L
onf+AF/NqTweR701yZlmWp9gjfdqGi6QBA4rEMTARo/n2ZLJSKAjT8bgofRTKRkm
1JIMG2vhLal+IFS4WPQjQ3nLCXZZ1HNCQ2NvYFe2YS6gLGER0bierUxRVD2o4Cq3
lHovOT3vooxzlTF4WVOOubtyctpJkBZ4ifQ1GP2GU+s+eSVqOv+qAaN8yCQJPCNu
0D+OpykbVjbkQ69uYFJ9ZXRc3LL1KdZ6CSvM/1fOQAPlFI7uHGVzHeoOq6pWVsw5
k2c1NodSFE3v39dHAQIbtbneVHYzRNRCmdi2/FQSLuBAigGCEiOPvLbGYEL9SAjx
TLv9wvG0+6IuN4CdXf1ZPuCtx+iFgVIxBpMCtl8OZS5owHbGROzQiZrF6yz66EsN
k8hJh+uqwmmeNphfatd8WgHKgY+hNPyJakif+mAqrdnT9rmMfL19ACAgCs5sQkUU
TaTqVRpPZ0ijo4I5lpy6pafm/3ZZ1jGwWvDihPldnT3Ud4MtTW/bh8I3k05CSJgd
f4UZfV/uKiGbWVOjrldPEACczD4fSLzbHD/fWLPKlsBFpPXUvSBxZnWb8w1UxuyZ
JpyJu/BJ5DPMhs0d1z/bf07FTfOuImpjjG3vZZZ5GP2gxFxV8D+HytZSeWWoqn00
/qxC6rzNfxxZrOJWv6eTVtQQswQMO8NV5ZfB90DhF2bn7fL3u8GiSq+rdQy+PhT8
ugjzn4FXWiESsN+MFkQ/HArg/AA9tcxWKFMSKcPHorpRjMTVHnRjSQUV2cMQxjO5
r3CuYrZrygKJd/PBQjPvCtSJ2f8eJhZLptcNO4dSoNYi5nQsFmGb1ZOK+jMHSluc
PkdALGOJe5xOQr5IY1EYA1lu5RTt/RyMYFcq3P5JqfxdjgWw3elQgpzzmeOs8TSu
dIrbxnYhXBNDRS2Zyb9p48D+lEcmlFmS4tjjS4qGs7Aey1gvzox2BOwkDBCJK1X+
PVMfQ868SOHv6OXybs0Zvha0Qd+vYQhVtdEfksdvRFOFi85A82WVG2wVVu7qoxaF
Twhg3vC7L5vz6TP+hGzF27V7E037Ua1jdXWH+X323RyUsN7X6rzhKhuFkE6EAvzC
Rt69EGGLbiGQptPOuJqB7BCMAHwsvV4jl1z7iMakukuLo0stEQ9RTwhF2htYKAMU
pnyeiBkUoaS/QcNB4yirYojWxBdIwHDQUJRMIevfAvIOS7soMKe1tge0UnrTuDmf
JbOdmJ99rGCjs79W/2dS+tkoi0ihF9hBxiTMk3xip4PKfPe5QgXPJXu5WcUQHCho
LHwWZ/3hvQE+taYcfg0wVhP0hLHk/cCwBDwiBdMrcLjQ8gY6Ei3w4FN0l76jsLLO
LHuL14j09E49gXWklJmnhUlC8val5Tc+EALwI9STPUUPZC3JnE/5PSF3Wq/axk5E
/8yy9UaB//P300EtdLUHjrFSQl+NtmxOwwstYIQHhMcuRFCdG5THYzS6DIRR8ryK
Jr9RptgtwQqguMSY+YN+OyEmgOFIt1zKzVzWMYObYcJzEr/OdpbcKKXrvDyJd/HJ
aipn2fqyTkL0UJgzAofD/bzLNwyjExH6m5oK7RT3rbSpYuMriDDBDIDsi6gawGRQ
pr5TEjOeX2tVvICvu3aS0cPZ2yGODrJoiQa2BE+iKgDfxx/z8sYgn783f8fx9pZ0
RkRQdGx1AhEFoPAn80IN9qNRS6zwwIyT9UIFrd6oqGoAkVuQ7dBAznHTS48iN8tk
wtAAzNcoqpIL4FHCa47QlpOAXf66HiS7gFgHH9CzRLHbsoggn9rQmMIGI1vkeWPI
Vxvpi+4h1zMR5YUtROEw3cgt+Lc72Dqe/08yP0+0McMm2VhzvPy3pJAXPuiD61tH
bLT3Wsvw3dki6tDuRhkqzra2kWHdc40zBZ2Q9gDULCIvGi6BD70CXnsIkyEmlfxB
O1/7dmLshcs9XPBBr3rgw85aLwN2FuTgT9L8+4cpK0t7OxBcoIu/o5oqwEkEPvCc
c6tujWV19st3KlQh3064cwOXa9JvIAAZx6f1NJbTlahqjpVdF+6o3RFFL774Lyu3
8eDVJs3fsaT9YrWsmVMkUGM1gFj2JA5YmwCH7bvYrJ3mql5vnCK+xihdQpo8GlnP
BygJ5mXD6VdXUeTEit6pBLzeifsFDhS/RKUKizHReEuaQdPwOS8dU5DN0IFYUIA7
+DQXHmgbO64qMcYYUDBEKa9t9vKTG6PemU7SJ2bGJeBzMzMHihkTkpgvElFGUIC6
iajM3rJHsL4aSlTauupCnkqDBGbjc0YhhpCrbwk1H1qvURIfbcMt8RMUGZfB/Mjt
CO0g1qL/pjmsx5U5tl8PZoCQh2flYkVClixC5fyDTWuzPUsWXv7+Fez+zLh6zygv
pkjsq4nfgVnuJ1RpNewwoTmZ4gCTNazmVqMAPH+tdyhlZ5nwaDizUZ2DW0omtWfK
yWetfZcyxFo5f6VSpMIPCEZgL2qU9nq+vegOfMei9jS5S9jdk1BNrzbCzz6U2esn
6U0f69NSc5169nMpm0GXAKr+PnxMLyHG1LqmcGcBQkEwd1kmLM02scoC3EPt5uOl
pDyVPswSfie+fHai5xOrHnYfEUvN69VjmE4gqMBi1YCR/yiyTTXmD3YTN4WLX5Qs
iPWlMvMDokU5Xc5ZAoCvn9LX6Lz0auQjrBrGeW9amwO0EnLeK0oGIlHDSlSn1Hia
6B57b+WAvRaRlBTS430CT2zb0Rtj9QDkKasi04tqTNTguWtfVneWeFjUWw6emQCj
kKSDWM6n7jzsumsLy7jnRLraCQKibzUr1Fyh7RJc6wx/kSh//GY86EigDjnViSDE
yFBpbxY3aB4rrRMT/8kQeHnPR+CatHyOxloGA2c1THawwGy5TQuoUWxTY/a4JxIu
NMfHuBwM5FwKycSr60eSJPO4nQk5iZE7hsYQRSb/eSbdFjVKt7kLvf+MEVHRMnRj
vReoQPRfCI/mQpLg+K1txoONbX42Kl24TjmhTVHNl9x2s5ThqE3pKOZ2OTI/PsDF
rY9Hd84bxkdeP+XPntsnoRFizdNcUE90rMhzFQDEcjF9cJka1r5tpZyx60jzPUT1
uZyL0xvBxMZ8nUJjoJKK8HF8CaILanytgvSmlcwKGEWz8gLzIkn33Nql2cnzKm6J
kmzOt2N2Lark77RVVw10FwsuNoLI41CG2xdNHLVb6MZUwBAkm6Dht/G7gXps580t
OoCB1gjfpc4gWTfHfziHivVGl9E6IYBvYtywkPas2DPMCmC9OZWF80LzCoL+XQ/x
At0SxKwGFCtAi1PGQHfvovSAN0Z5G0WN8MatxoGkEh1shFTL+PNk8YlbbHm08Cmj
cjByD/wExRxc57nWUNqAVfl0ml9Yy6+oNTQuOI0/fxrXvBk2RBC6Ya8+DdhyoDRj
P5ihJG5uBut3SpxHxcvooFffPAQdLYebXUSB/uwfOTTY6xJmLI5WutYS826hedu7
X9rO+d94UI7GwKM1jhQaw6+WeTJ7hL5ETVtg6lSNf8e7G1/JLVkrbzxKbu4UVLFs
Mb5flPgPO0h/wRf9RcqS3mT89t1/aSV96kQy4yTWYOUUF0qmwLTZ4XBN5PdLFdqe
0cRgXuY5A3pwcMEHN7WvvhBiZz/gv0UbldsFTLjpu4lYnOokVYHfLEcaknJ9qUYW
vhCRYFbFnuIE+pwsD0n+U7VGmX+nAvMBrO0Ur6RlCi8lqp8BD6Y8Dh4izD91z/jh
AeB1YawL0egmNiY99Mu9Za0FoPidiL8qHGh+79lrqqq5Ip0MN5iejIRuzxYwv99z
xm1e1Lgo2m0rCXZ0bZQXYCSDHIiuTc2EwWL6cgHLzcRxAmKlOCmX5U02eh64AO4E
cf2xnhJlBmVo+IPBb1hnH6dGmi0V4FNFV63FtAvCrERHf3S3KVHLkAwmAgKbrKgO
SutIppeYQPXQN5/HdNyDq38+ZUgz2LyIa/VOtr5vuz/txO/PDJxtKPlvW4QDYBW6
L+vSef5Zs1AHnJjJnN9ByMdB1FBYe6Swe18gBrkBSJKQ0W0AhfzW0hcnsqhNOW+x
aBSb+2yxm/+a1Cu3S+I35CpwODsFbj3kbkjDUHxRQnn+bqlQLSQ4AU9UFEHwswib
m+qfFivIsTeWatY5k7s/G04T0tlVJ8WvBqQbPkm8YlVB3jsf73X5A2u0xvZNgkzd
NC07nE9TYX36czf0Rz56v0OMqxvUSeOk6MMwFHyUcFNTXZvkZSbbGVNr3skzh/s1
uYyZuegIgVOK1hCF9Qrt+tWDbpbwDa5u/UfvJnOatNl/lTEonlqFCDSggACt/qzf
678H4Q5CA+EW5qh/mASPFXxxE4uLGcRHWhEBW+vs5y+tgbtj5MgokiyMrmP0yRaN
1hXJ5227eoQIfKWueucD+z4kB6HncEByBgds/MaNPkZ1tCzzPY83srk32wYmv0M1
PzakDJ7D0UT68WY75V6cBqkEIJl2LzeSQp0pZbjfg6Ubd4NsLYWp8mANY64vmU4t
s+GKlnh0Kdmc6CnRISBBnq6JEgNIPS3TW3OR1FifPW7cX/qjXCNHWTz3xUKRPtP9
YdwiozKGuBXuxBD7usfoEcv/EyaU2jceUZvCAeOVDlp20FI42Fi3o7H8+B22h6eY
yuhTnHEMX2PZk11qHj9D36S626uYMG6NfVhJzCYarJJAJp7TXSQRrEcL5bzDHKYl
KrhMQ5YIIstK61vSeN5Nm1lBrYvjQ2pX6yhzcJNnqZXMWY7DVEtYm94VA/kRJUtK
h6Ul78WTc2fS4vahLw/psr864ED3cZ35MsW3wEW/Mc4JJ8hfx4dTFD+DX01ZGqSC
m95+dk27/CuBB4Q17HKEFcCNg3nUQi/PaQ06/Hlv6KFvS/dx+KGdlrxbNhTIoe5o
0XxxgeI6Tax32V515dAND3okZlmBr8k1dqMw09SxG82Kd4kv/StcJgAtUdEmc/Qj
rfDzvlyZoHuqBbeBT2sQglhH6kSxa8rCs9gQ2M6T5CB7uPkQjSqy4LItdg/8KZ4z
39/53rropZFWcemm/URzaDGuzTP+dDr3Vpyml0V6M5E4XCfGEt5rE7Ncn0w//ZP/
MiB0qGu3UpUZyhEq/thZ0SgCqmo+OQY9ViXQjNuV2RFKzDOn1SyoYsniePtLBy53
6CSNXj073dhEbAHu/kjwizhqsQk2LAiL6PwTyIWhZRw5HYW++kgHFVtGgsULr/OU
/vtGnEn6H5Y3IbYnRqAfXi6AMjo7paY5gzqdZy7LvZzWOXIOq2Ca2ABodFy09xNy
M2rlikLQ86HjvmxYwKIJnnZCDrm3rrRuiqJCgSBz121kBqxGH0q4G7z6/vlbg77b
2X9zECJ0AUWpKKAYcAGlGai79+DqmqVv7Jk8OwEmm9lPWcr+jzF2M8FVI1daNDBN
GbdxYLDDC3phwhQ905PKkybUrHG2z2HoBI2f2sZ6p+plarPoe5QSVwhA1x3xVh9g
BaI4sQdEwNoD6Kjl+evGhgmdutHuDoX4pRivSwoNSjGReD2T6UF9c+hzHLBChbb7
QeErYe2QYcpAiwk/s0dSSIACfFgM/JNqPWX6MERz7egT+UNnBs1INE/QCa7pXWCz
Fp9ZuJ3xEYVaDrgmGUxnRyR6dVQ71seZ/73i1yB0EKZ3qZwZRJcU4YWho2oYCsTR
Y7M1TvwzsIS8JGhKcfdq5Kc85Wc+00FKGA6VYhukeOGarvim+ZTj26iEISYix+R3
sdd/IhG234jWdJ4iFjQqTvayMjXrUi9HZ7Lm+HM2TWfCuVBPRjyXyhWfv18z4137
+eoM2ld+UnYU2pAJgeMvNRO+iio7RJtBYxVxmZOT3TDpq3OH6lSI3nB3ZiFNyX7z
8UoBYJMf7iNl0+Uq/Vouxh9w1N0AE2V5mu614QjrZ8MM4LVFZIb5q6CB9FS2tDFL
3sXWILCqN4Tkdg8vpN95bxx/lYbwkf7+VEKmRNUwSNw6MSKCPvdmdYo4L5+sGdZc
pmiQjFlwwRLTpFv884lsiA3OVCozmdLV4mv1TM118fbdGHippyGeAClXkxhAXdNY
eDLVAaMRq7TPosY5cD1D6XSNT8USmmlcsH/dUVfIWxDCQqbHRFlljbLjuNkwo2Ps
wCKAdq8FlYUelRGcYUWHLKO+iXQNXpwaoqwkIMH8qmZtt6Z5DkA/fBdGhwhtI9RV
qhZAsFmqgrRpBCTTqQikE1ZcBV8pKVcM99kWZxZYqFbYCdpgqQUNlvziP8f0FN1h
kzzYOTIzoedz9DMXkSGAIQw2Aycg9KA2bTnRhLLygX2JVA3tICOfma45e5O0MyF0
LVEqfLQrkefmdC9WXh0JP28R4YI6W3+ENMwbxAllEgiNKLWxcA850N2GkiwE/PYd
oTQcok7BcgmeTfWAbWVwivHHtTW9SvhsOnRe0zn8uOZ0E4AzXtA+flMCH4rDjGlX
R9smkATXTKu3cpKebBDE7hgaWHDLdx9tCxNfzI5rIgR4rlh1YyujE+grabKk14IK
QvfOaXO43603ga092ui88i/LXaaspTW5G4AybwH8VaSG8uKDIsJOKtHHb5pTPuoW
two8zHkaUVT87k+BCY/ZlLw0u9ghWSd3SyZiMEUFL17ibpQszd5RczpF4y6/Xuf1
d+PpI04EqNJbcuZ2Ee3czgKXrWsxH0Z1t8puuERxqktO24CoocPA20aUy/OGHNvr
Kfyohdour5Va+1NnWt7RK5VtjnURurbLiJdmMObyrEp2OzWqEbsUpWY5bKqxIy4W
Pfr1ekoPfNykpLMTokH5DFyCaIQdt9voC5e2MLp3cOoUd8stmwMnS1jmhtphdA5D
gfYHBWi8JHnKXrkftAZYczrqkLkkeLugF6bqN+28L3LXULV8I+9NshH5DxbgEo8D
Vwmwt8Bij+0U9lC9WeXpXBAVa11khqseaM3jpzWulehog1nxg/yer66Jc4KFDcpI
cqNiof50f2v6IX4U83bG2yh+a7enGlmVM/ZetI6E2TDEPoEFY1RquqsexIs4tCQe
EaTNA6odBi0pzBTulPJofvqdTD9SOuYv4wv0mTbpBS9JWivQtRwZRGPhlm4KAWiL
KbmhqhnAcdyotim4SxIeErr2KTdLV6alV68txsuysHj8gGPIODY3R5KSEH9/NmWw
2ba5Ruw2fnZWIK5rCWaEBaAWRTK2Sw2uthL4smKSHzgNPMY6V7yCxshGNeUppS77
IeEsjy4KA8eMStCgqJB5ICq7KPclEvj1aql3V4vX1ci3T8uJo5JMNcb1SwIrgKoE
bBt8LTWt9/71gsXoWBNxyTSP9SAU7GniXCdX5M758HJAaR8ehs09L18M5cDUkqyc
410YsxmB8Scgpa2xl56C2ko3M51k3TxaXbR4rLTgoBRm5/UkAujAmhohqg02njbH
uPMYsuMtu3J7iZOC0jBjDrofiDFL5qOczA8SmZ/YBm8lB2gywL+JbYsDn3Y3Fb5Y
vFRFbiU9AYFTa4t29goRvz15BvDCw83AImfiy+9XBSjmO29fKiUBq5f9AL8Jay5C
oW2k5/QlVk0HrKvog6705HQSIHms/9ujIE25rBXoCjfOcz5Vy3U7epqvp+hJ0l70
KL9/3t5JMgEWJVohHPEQlbnJhOUscGIKr0/bH0g+lKBkZ+XIsxosJh+Ai1cPNr3X
ChxI3EK94/N+gnZ18PQnDYtBLitjbmSFnlvrf8z7bVkHycqpD92nytx0wDTGaAbI
NOB9gZHEj3TR/mirrcfX2hlviJB4fA3ks7H6+Xzc8NlrYrEMmLFKI2b14jMPo9l0
Z0KF/FS82jVE2OJsgsHrNN8dRrODFT8XfDIUtsDJQujJMpp6FwodWI5rewzshUUo
8eHSykUFO+O/E3Nl+ifHf/EBGz6qiN/38mAqMNdMcT5y4arSEmNv4YujViVDv7A5
/UjC/DjJOzmUk86h2gRMtBOyzgejjBW49XVx5+X8DpX22pAMpn7h4qHT55TVcnp3
Lkg5ubiYqlMMM3xkl5qXLAbXd8Sp9oAeRRm4MGqYV8FRC1DC19FDZuPrmKUkI1SS
N/48PauzIOjXFZgae+d5yXfEzTfr6rMcNRs+tPbXg8WZZtVfw2D2w23sWCdqsSgw
Uz4H9JTwj2eORYgH8BxAzKEfAZrAgkKgXNAJLG4qSVhUd4n/ZVIjvRI8JqzSSEP+
9Ka3HdxwxcrsjBZLGDNZpQ3euGgWyZVhWlFwZ5NswBMrdboGsTNoWDmC2I219Ce6
iiBMYRNs84wO3zqy1bMEZfmnOpnZYZtrMTp4tPsB79KCBksc/0wQ+nTRyi14F5ZZ
Yo+uZuoi0FQ1UnbgGD+MJuD17UwuHlknE9zzN701hLLiJ03xCdLsjSFhWzRWqcsL
GukdLL7EWghLaM6qoly6ZRYaBrearQgr6DYPJKHANCDUks7qi6VJm6cyltuesD8R
lZC8s/aXr4B/k3uigfJfFS5YNfsElnaMx3V/8OyY/7CAtk9QeGyBScs56ZzJ7okw
OBPwRU4VzdYd5A40YtGvwEGc4OaSRqk11vzrJIxxiKswpCFDFJj2BirRkORBUkIv
PBUR1Q26OwVURm+7g81Wyz5/jkPvkVgHgaMRFt36gIY7bd5X14AXYq+5glXeOiuF
XBromHfV/tJtWjbgEVLGvKgEv/rk4cLbVumvQWk5W2HIsfgMgOceH6asO1pi14wI
eoKm0quwex3v7NcGK+eLjzb4iP7iCWA6sPnzcbwq9FVcp+i4h3oknUbpqPmkbWDq
bfPOtc1Vn08XWPTQgS7G77GJIslLw/Btk9g224DUMvaFK264539uR8zzhzG1HMj/
8b92Ubc+Jeq601prexI3SFB1ZvvrX/WWKqe6r0z/ClWlGwINT6GvLbbQl7rxYkIP
0hD04F9xDCLl+5a9hGkU4PRzrTBrBHEIy1p1sKZAy950P9fq7ODhj5yxHylezSmg
KcSsJCchHqAvBEYo8ZlPf363TEv9XcOdIEgt+/1/YJSdJ2MDNOP9vfe2hSnUGkTU
FuA3PGsP2pMOjWNw1V+/cMUiOL0uyp6VInR8CFw2N6lNfAOe2TWa3zBmxg+XL7GC
yk66Y70+Qjf+m/mLf2zSAU6vjrVwfMNi73uzBcu64YF1LcmkRKIkppEor8s5itLy
rV3HB8juBQm1Ut4SVtEF1qRUoZn9vm7vopwbbEljhSElCo0tnrCq3FWgFdje5Nl9
VXDkuqQwCdtwlY3DEWb+M7z66l9wt6tuSZiaMMVbE9vfqZzRUWXebXcVcuuP5NYN
Y6GJm1zBf1QyWQQswe+KINb9seAjB1hg0rZbTmLT6KhwlUsIb4SWwxlyBVAQJ8i4
NPVM9Bqa8ZErnxmhBXhp0lAgKVpokLDe1iWITpmMyv/lWKtxj1azd6u6wqJCkMHs
uADzB9aacAu8b6VygYwZpDCQaBfKtAEmduDtELTDyPcGzK00MuIFm5yBBwn4Ke/P
Z9BIh4Q0aEA0Vo4eXACOQGXDsxyNweQYamF0+HxcUqRF4QUEXIZOmlmTFvYTW+wh
bLhZnSlps2gM8AJ7OfNG3fy5d+6HY0MOcAuRw2p1sfOuZXPrR+hIlpQm/LBg3qnI
lAPYKCJztNW8drg+8/qagY1+DIcdYVvsFw/G42n1nXxo5NsmnreGtq7Avk75SsTN
Qq61j+Sg0HEInUv7DJN5zjnG0PFX5fGqtXnctq4X+mjk7IfN1xzA+j/GSSUqFqsj
5L7tcE3qugOqIqtthWz+L10XH9+ahafrwN7pnlWIwKljwBI75XvnrYa8mPCxDDEH
y4ETNcvnRuqs/tYvSDI/230/LUINLhFgxRPdnj03WTAYCW2aeQ2pWbQylCQSFAJM
9duag5U1MyZ3eNWkuQXl8fjFA7gV6jqZDkxensMa1zdAr0i5GEy/LHS/GepQDzG6
bF++lGp66392yShQoLBijIHS+xgZXdza2ssqCwLtXIJqa2GWDrp2UkdV5LReYLUt
oR9ireWsRhwwzMyBP3bQ3Vn0zMEa/zWp9BcTwbU7kgTnyLmTvNeSC80HXmcPkRCB
j5n1LqnDvQ5sLHgMUt6vk/fT6JShYlp0jibyY0i53rP/TeZY9yUdZ6i0T77AFZOI
2weKl9dXpoBptha+7CWLPb+PPYiEGY40DHcLqdC8ZiC6Yz6qrWvKOrHVKsM3SNob
IwkTsPGPN4tsHtFaEepe5LAushuwB5AnhPba6+jwSukfQ59uudcwT10PY1Rge4Ep
ARSdwfMHUGZgJ6AxqdisII+UkQzJF5IwJxWva9yYh4pO7Kp+jefcAYYOfYhouh/a
NKB8CXrgz4RkaBmUrsPN1bnf5bcvbbY7o0+XSRuQ34OSsgeLZ1sSkjpIe3y0PFFt
W294MLt21YOcFmIOBKXbPLbYKfySI8nM1hydUPB548Fy68mjvETct426XJlc31/V
1AXTpdZZXCidkQZZ3pDQEslZDlBJdnjybsGgpeZszAAtHKYp8WbDLmX7T1J4AKBP
sKZ+NWwUpgyq88Ek4guLYXHMtx7P2hztZ/irweB3hPGHT8qRm5wF4wBQVwQ+wOX8
7tHWh7MFl35iam3P4RBNqKskzLAuBkU7vrsFlN6WkaNEXwmLjAf1NQX3RiAzhzuQ
6Vi+F+oZrhPGADCGYYnsREqZhRS3FiK0D/IaAXySKNTIBuWE2FTcGze6Rxe5jFcY
ttd0DLgcPjyATWq6ehXmpB+1YeBwrIZvyrxnAsJvvDTUSFgzGMZULZffERNWvbAk
v9dz8REAzgT68POSMA1QT2iGgofQTN78T5QmfqPPQQwNAg1MA1SRbIPAldNWp4ZU
3ka9OOa86RbPqLaBokTnAoakSDZBmgdR0dB7BwK1tl7TFNN6UNOsMKH7TmCAhFVz
SlYwO3CKEet/7oeN9O/OSWCAvJK817S5GbbB3YZN7+93YFpw1M2ZLuP0BdtSsm70
7owIm57rGExoKb4oGcKUbXH2KTsE5AD7BZgXYuJVnysADcD9nUB6Kxk+8GRu1gUJ
MTHCxurpxJn5FfQy4rqAHwn4OcBF75affvEiznVKCem4miSgIhrmTtspv7/e7Zqz
oXU1Sw5PMz44RZfeUIyiPjdwCrCM2tIHUgQM2ORCM73Z/xEkHUcV1eCrN0ZEnlV4
fAPn0oxZcD7Ympp0ouJpJ1mYddfoWpljS2x1OZaDglmnAguSv0sYFIsEnPFFAsxS
DZzUY+QKqD8rPpS//7saZ5MyM4y3ElAcGEmqHCcftw3LpXVYiESvvwxT9DP8FZ3t
FfrXSFKr5rctpk1Jf9LgPK/WQ0mFtqK+NEzRG0UrUIBiRBz3SGQRYM0OfxYrlHJY
plWFQp2YnfzqHE1vDIv7b09g07a8lFii1RH/pYqwlmv9rLYe1MkQsWvoNC23Vhsm
w80SMdA+qfh4Bvalwa1aUwEBdNN3xDc47GwW0muWW0ryIhZZz6PR2wFB398O2utn
Sco0VSgVmwm4TPP/w4tK0lze3zvD17mv1P5uHw5kQmW3PgSWCeCjp/SJ/4JQ6DQU
dMrKvbh+4HWx9i9b/KWCXsfvzR2qoRrwYmFncHnlrmKrPoOWR8vO4X5WH4+oBVDk
rtdryHHq+seJb9m+RvwH0pn6+4EwJR+PVw5Va23Ow5Xff5dbd670Riii2NK6ZnXh
8I837dw22h3CWkk+qkXi3zUQsQbxooD4w+zMCMnb+kFSlMBWgPSuCFmiEhGmmfRZ
KpJZUfhS+TE3zcsVvp1Jhp52Q0zNLS46N+ffFA6Cf1AZCUqPqycuvffb2iXZDEqr
k+sDlsZW6R85KK3E++2BY4DycElukfSnY37sYiTmLuc2SMiRHrdEn3+6/qqtkrN2
e6UXyL2ND7c0XI/xaCml2sw731BhDn3OSwcR1SBNoEOdP6HGlZsW7O8JbEgD2Po4
lsFYb/X12osqabCyif9lRGDWsmg7OdniGA/e2Mn8xuUuSVr704KYS7FvmJytlPiw
pjnX0HzHrxYYdHjrK4znx7yssbu8wiFNY/4lsTNtrb6blj+M8pC0/s+XH0eIWwFH
We8/WWSXQOhnftOn5P1NELJcN8pFKV0COOpwgR4fZgTKTKD1UDIOvR1RxAT13ofl
ZzO/cMV5jgGAiFBPU05Ecrhs64f8f7E+nGSH1ZjVwwnUc1PkfHBebC+nY2yOsNxG
KaVF09R4uKZjVwlp1zUry1u/1EJe2ykrn5OI8cCsUEDkvVa/ZmllCyB+FU2rUYzG
GWRmVEDDmgS8r5LfRI9mEOITjM9lDyzMTTk+W6GiHujmXKjdntEsVP5OKzTdYwRD
3l48ZbcrAkc/ZdzzmT1+k2/kdXhWCWQOv4nWerrk2PHocvxdeTRBJ+bavS1DExC5
elsqtJOjc6EnYeNk8wdAxz9ye6BxyxRjshin4HCZMr7n364T5qaxDuMh2k4kDrYt
3yJPvex5Oaih41V6/0gh2I9Zb1Zq8mvHn+9S2HYsx0HHY4tgwr7hd4B/hbV9Dlzv
InMQFHeCrVg83RQs0fcz+hBii2nnMcRitKl6YUFe/aV5GSbKyW50npaIelAJ0DfD
4AGsJbRgPFHPWjd2kGCJ3T/zlMH45DDdpajWblNEvbdjorqBWLZ3ig4Na1WC52MQ
lriJZOZG5rkZzQ80TbAhYWkHhmZrrFmTlpLYzir1uDaJ+8JHc3a5vKX9suAmLw3f
3Ef8oGcu8qd6jd0pBwV2w+l6rq1sBtugpeuBBhx/HS6dBu+0QgL8GL3/Ikk50WLt
V9mWAXKnypM0CyipsHgSR37f3345Dz7Xh/juiqJsmVdYOsolDWIvSYkwBYm4Sbue
IyMQJ9Cwc3l2OdxugibO8PhCSBBnnHhC+/aIYb7mzY8vSNzm4avK2uRXg7JZolQ1
JdRXOvIinU9NTo8pbXd5O+y8t/HJQCJH6O3sNajHKgziHV+8V+QylowATUgBZchq
mzTUzTjK4HfbBt6gqF2uVgsaafaEADJWBbZzw/hEOOGIGXObw0fHQVPow/MCc71R
qh9KAaHdQ361AQaf4lr+hUWnH4Mc6giLQtjqtuFDoKa9oHOV3uq7JCPmH34LM8Rp
cjH18g45qrxOzKIryc/I2g4EbmPD3CSXimMRO5sxpYAbbiixOx1wO6O3mrM0wzXo
cuSpeAvG3uWnTxb0+xw5ztuCtE21FTQHAJ1tvCg4moUGPgIoNFgI9psh5JtsRN4s
7hCDNGQresZErw27+oUx46kPCRNiizVqo55siCK61TcjWV9HjwFAT0MCrjzeyjos
zfcPN7IPo1D7bNFAKH87tXonBgvzV66sdFwKLU6j9MA35OXU3AdUhSXRkjTm4ctg
Y3rEM7xZoC12/DqiLJkRwaQCDgmSMmnRkBEwgbBzzGPEIueSgAcm7zkIB6Tup4Ml
u0FzDwDYNl1fakhdbZKM6lDzyfCoXxWPVHA6ghQK+KcxSeNs9/H0tublObznytoq
72ecwbO0q67w3UaivfMQbcjrKmySlSFfLu+SrpXCcAsPi0R+eCnzXUx2DOCfYiQ+
GnldilxoIdGqZgrgbtErNURzb3x2gavNPQags/SI1dAcK6oerEzlokyDir6RwnlK
nJpVQj5eL0olq9/3f3cIXQeDXuZNN14HXv4FUD40vFE468rXcsnZl7Gl4LBTTfqx
CXNKHlCOJYOUJvEyHY/hPybj0QbKgKWJVBNrNyehQ4UZur724SOsvA1zEXEzcjff
qFvJFPWPTaYMz4bfp1X3SQv9QWxcjFA+FyzkUqDYpGcuYFeBgoqYdyHMyKZ0AXCu
3u0zLhJA3UB0I6KjCAHVwD5iT5ZumtUwcVjuSFLHmuycemjbRMObLvVriqC1zGV8
9Y316wjzaq1rmW+cKtotuuBmFyV/jvqy7r2vQ1ywg6VsMMz4M4vY4wgxZmlam0VH
5m1WOCQz3FdEK+g26XttanNYBXIKpIpzrkJEW1Sc+Tj0TQjYeFHb/oju/5JPRNgJ
Hft1Ga5dkIpM/m+2AKQySPtn/BG9sQjdj+6vSvAP+R46a0idyU0HWqS/wioCRiuq
ch/0/xZAZ/3uKhppW6tjY5i+c9i5GFjqWHiNOcB2XxxanyGR05EWmx9iKqfGL8s3
26M1PS7gMzBwgbi8cnkwjDK/S7beD/vk7vxghKOh+bGZvZht+h1uU5KrrYdJvVcE
yWnS61G3dICM8Z8Ef11F2XNgYVNBBMXSJ9CpaI8cS3d27FXpnL4LwyCteYh0Mjw0
RcI2GNtOO+IPWyXzSsaLZslppbGICO/dv6ObEEtDjrem0tyET4gId3GofyD9gLI/
PHNRWdTbDYkXrNcSUv2LHPV9bIFhs1yIdiSgWBFEuTnLep/hza//leLLPpKWLThM
0mYjksW4z1wbg84GVjTG1GgHWG3ugdG/XkdRhHAGShFsIpOqWKHTxam4dLP3LWR5
FFoYEqHKmHMdktC18IW8/D/b6HjHto5BOiBeW+rPzFYzU4kMAJhH+ESfcoez+H24
McGV16bWfIxtdIZgK1Q29xLHAjOHIEQXajli7lukJTu6IMLOyX5Z5qyYN23z6dEo
VdHxhifbmmmaaUp1a6+7PtuUAv7hteFFJzsfgCWEQYDYg+q7w8MTjZWr8QrGZnsx
5izWT9s14OJzJTxnQdGYYNLtr43nM2JJPWWfQ76C+lxzFNoTQFV6UAnegI+QT31i
S1bscrZx/bY8uYIQhSvelDdnZEsqdJH87dL6936IdkYv1vqZFBWunxNRAgg9QV+S
JNugGBz4EFWEqHNIJRGvY1eXf//e7WP3mQSLpJPXdzfcFSwd45iEDpKMT+mbXQr2
mmJ2g25BVdHH5vNWaHBD9Yv2XPHmqsZpM1pEd1d26Ulmtx4lodNXgabsEcQgTg8s
ZK3cWV/abDCqptidCupomyHl4ooVWTb1QhG8tB/YHPb2e+eteEBwp589TtD6qFfu
C6THkEagrevaoYwOpPaPDjzGqIF56EN00EVy08PcHJ8vgaM6LFKjKeTcnKTwOqqs
Cc5xrmaN37GJMXu5FS5VqUUsxUklRGj87nAicLed0A143yybCHUkYiZ2+OmcoqXK
rMDnnYftzvsJbRc9m7+UI/nN+V6i2fU+oT7Y/aIbMVvXXrCn+3LN/dOg6HRJh3A7
pqtpsvk0cs2Q85KTKcnnBfYsub8hbObAhc+KF1PNuVPDai+CKN6/WBXmjFf251/c
DvKpZLaTQpvY7vAyEbQ4UUR7wgJtaWh1lG6Z5VP7HrN+/WfZynA6khgFwv9BkwzX
eBHf2KHhYr9uKpWSF2ikwaLB45QTabHGvT63WblsRB9SOqmfI+JHN9dbO+excgPM
+65/gATbNPkAHUKHK0y9wfzK0NGLzjftI827OhAZFgjOIoNpXB3/2tV17N6ScRVw
vQ/wT+tdabOnk2yKdOZi6V8YEUeMAUObW++uLNGmYSdLShIJhrMMFBlrf/khYm09
yn5vTMZT1TRxpoTnaIa745x7iPbROoXx7hNvwPi1Gn9Ky67vj6J1aMFqIDUNT+5a
4Yi05BgSqn4k9bn9T70lMV08Y8cnF+0ItUSKlHx9rvScsfNO+cx+e3mqXj1FRe5D
bdU+kuyx2CKABBC5fFs4XxYYCqyI9PZAeZ+Fv9VA8TZaro0Tcl0rej+Ne7R1RVpx
x5Fhce25PwGcqhzpATmvrawqHCvG2GY7wRE9HRqrqVECniaTa1e44T3debJNIEtZ
2Dlkh5vCpL+FHDUfSBOxK1f9LS+DMFgs33bfj+caGTwupEc686dGqMX5rsRXxUJE
L7w1kRWKQm5PBL/LJZTS5UclDp6/bJZeXkLLdQXFhyJCXNDzhtC4b2vzf/jlo55U
lFjpFLptToBzSQXkglWKyfa5L1rUquD5OYh0AyLMa+fjWch8UEqWK9PIuH5TeM7W
UiyOcRHeP2poEMjSgdKzz8kJ/cZ+fpag82mW9LIHv2cN+Nru+4G6bii6QvpXshyl
O6ApFjzFIqxy3JGMOq1r3k1EysRFdRC99WPPBHGvOcX7Q4/PxnxzYYQGHestq4Ek
wy1aHYHDFTXsU3Mvaf8s8RHr5VXHTwccQ2Y4LlvwLut5g0ck2wHJnJxFOVTuGsry
RbSozTTl+ZPMDBDkdER2q1jFfePiOG0UAnXXmujeEW22VfrrOmYr89ydWC1P5tmO
g9ekgM0FWJ3FlEYUP2j5+Bit46JdRaN/UlE+MkSP0BzqeG3jWglaRSpmB++7Vu/A
9dxcwwXW5B81op5ZBBhKbiTLVQpRc7q3X1UNndqvgcTV65koGwW9IMwVKMdTQgDJ
gyBkXJ4QnBdvFoBooNglY8aESQO+qED/wl6TzggTyhNF9LVbaAgtzL6gQpjHK/ph
Yb/7luQgiOzq+Ugn8DWijGWib2WTZLQEQEJddw8tFhB8zMACzNoRuLLy36JxMfh8
IdE39Oh3w+DkeLgfvnabOlWU5XhEFAzswgMBRdDxCiXFMRAXlICbj7OKBZD+FGk4
ICx3UGHS8xkEaqXwNvYSsGAIRWW62x5HNUNv2H6m8KddjdzgJIyms/PK6OcLw3gX
m9f48acARXjwji4ck2asTBEeyYw3r1yqnbO5aQWzbOamDSFZYf6xc/IeIPJkS69p
z2+jVVkSq0fdoBj68tTt46OLPph40HhJbIkgmGUX+nGvhJPGPopMLnNXDwEXKVjd
uku1f0H1z4DzhMOrCJU4svnm+Rh8WYS2e+b7BRzw5y8K/RF1d8vsUT770ueLUjkl
xG2CItiUBEqqlcxhSSF+NRqWQQZ6+/EJ3bP8i/Zjefu4gWGSJRO1+iHnK0pp+AzK
lSA4DZ0K3atFYVJnZjVi0NQTLqcpeBggLaOBXpoNqDfcceNtxPkO5nkMv45TEnQL
UXvczGCpXg0xVAZRGZl48I8cq1fCwDIu5vBNY5DYH6/Dc1KmctGZwHSpzE9XvqpC
pyrkujFo4CsXWtNHMrlr4+iJrvCKQnHIYP4hVCrp+k6MOrCEg/Ym1vY4cHbWYd1Z
gUowRsd3941KMDe4WfYB8Hwjj3JCmnVaXEzAUHBzsZConT/TKWfk8fW0kX2ZwLP/
pMDXuEfzkFFPfigxe3fMKT/99lHzlDh86PxJ4I1FurAPEU0+h1pxGzznVTdVHsHn
Qxn+/gZ5IYS25fxdp6ewKSXw5QcOZ3KdeaBIaeSYMzkFz7gxednr1AbbrDNPJEOO
yLK7WXac5RmZqxjXmQV7ZuLytTYgB7WPkGOUdGb3sxg5TOc4vPr/Q0u1h/VK6/zR
SH371XK0edMHh9TLX+iI3v5Z3WHQU3rsq2ktdlE/IOwvJZvUGtotS0d1zRLrwWF4
++WBMEWU2DsMp0ovBm7JKNwUF/+NSUhfF4P3HBUHilGMOgvMzU/R6UDzhxR+Aj0p
ppwIPDbfmGrBPFnTnVBQjGXPzsD6njpVpCHhvHN7IyaSuedKbIZPNQTQccElrXQd
MD7LjA1Qyd/A40t9cqJc6iUl1oapm4Q0dI1zBHWT1CNVQTCrABwgEP78Xj/TZeVT
CAt54mgCyIkzHQEVD4rSeWzZVw5BKSzskATIaYJRMvbL5xCB4/75r7chPLMa+WuR
SLKGbQGbH6eUXv9SSJKvB6QaVx3MaHmFh3wlDJsPLdBBROcCcJPx7t576kOqDE0B
QCIvA9Lj9FtfX0dcRUSwugZKPsXfBhM+57ROFgdk9qkFuFPC5hbAEfcZ2rGd8RgW
LvU3o40cHjGtz+VUoMTiqW6H59Qw6jiEHC4SHELnsXp6c4XcWbIYf2Lsf7M26n+p
WSPKisWQt6bslwbHReXGPE2lJ8bU3cbHtOOZf9sJy0Qpe1vi/v2h5DDoLarQJu8Y
1x0/pTNYLKi7SMiwcqABntlBGlrYuok4/+nlot77zlNbF9juhmlGaVHJaMSeeLAr
9gPean0CpNa+E9qd2QSgJ+I2p1hhXAKW06qsiUNH3qVz5eSYYotX8Mf/dr1utcBV
becrdc/ILEuDJv+dJBnzus30zk9wzs9Ei9t17yF6Jf10XbB1StjZt0L66a4dMsw8
NBhd9YUrjfQMajZ2G0EtQ466p/++E2r55NdJrM2KLRKndUOSbMJbc8XSF+ZP6xug
dBExU9JS1hE1qy/CoC/k497JSlq/o32c1tYEtmFzco38P6JR4MwnBQxWq1ZAiW90
elRxRjv28E6uHLZuKpPjWdqOVj0mHgvTQpxQe7dPGNv22ntonDnJl6ghGAfv0ROn
kZ/aDJJSBa2MJYt2tjOSCFLl1IqGXC0tv8szVdZZWf12U/udAWHSTxXieUJVlZdT
5OYqLTYxZtwMKCS12WKlkIodxr19EMa/NdzplpOg/cmDovJ1n9R2MrHHv68+lqqS
9IlT6w9pmR/Iy+vme1saKtBH+Tz8KWA7DuoKHli/+TKszs3b1DTqc5+GS7lcpXJx
aBOSMH5NoQhjvaYiXrZYXFQM2HvzhDs9cX3Yfmw0Q/meHK0e8vlnSdZH3v60vcNI
2YPBav4s53LSvmHm3tC/HvTmX5X1WlIPIeftdV6kJNdtEUNZVuzpUlmcSeNk22Gn
S1svUmlvnCfLAmTP026lXfVVm39hVk6oiJPMSoshz05bfRN6kaplcDSGwrWmeqRa
Oo+93/c4GOSKUzs0tC82ozSBX9Rt0odYxo1o9O2ECIytu4vYMdm7xKYc4AGgy5tU
cZSI9UlZJi3QSgoXt5wO2tXUgwt/bQqg9ENz4Go+GGcMjpLiDy5Sqt6AzujNa6Db
t1p4SjQgKJAjuKiVHrvdnmRcmwTJZdNmm8QO/HrGGkmE4cgIbnXN43GqCWwK/j7b
aKavwLv3h3h/CmGBzhh26HZ3di13a+e3d6UsUUgX1x8tmbXv9G2b4GqcHPA5HXFA
MhZqW0aRl7EGjGYwupqtdI7uiDGhgLW45g7vv/8DO1PT4O6tGfIhXO2BCtV06DMr
BWqCZrr9IPbqs/FBlPTZNRR1XooBwIaTbir0SrxanNuB3UumTHbULB9UF3QuEQkG
379/Fs77HEzlaOmc4i+gKX2bFBM8SBwUoZZQELlhphewkX2qC/1g76yX+V8euNJw
7VMx6HAd29vByjnXY9ZOy3Qr290LjAmMIBnXHUbCCZyrcSym5elmpKEVna0tfzPQ
365tIHmgyamRa+h4MkKr2EFcCKxSLdit+ljDHapkM1UAdiy29WufGHOOdh1Qfz1Z
97A63DfpxvpJQyZUYmvbakZEcdtlTXJd7PmOHOtRy+gmoHD8DndC4Oew1nJh/R0/
1HhJNIwMlFU9j2xWAHrYR19K3DNJcX6Xs1SGxGR4fBrYvh4NbJ2bOadXl8BhlALJ
8BEnax5zlzWlFbFMlu6QWpCD+Rcv67iF4hS6/HNFsQu+wH4ToA8RMpt3FTv2+sBu
soUGbV2vdc51Fu/uRdjxnKgYoYncW4BnTmdm4XWcOjt/dQoszTzrFuQydCk7yKxy
QW09zIqTsl2YB3b/bYKgKiA10FPENjqGqBV0bi8SH82Bn7n1WlWD6bwj352X6pLD
OB9I1Xj+TED3q+JSNriJ0At76DbunKfndVK4PE9LJ9M6BHP4zVB1ZDfv5uhlxJA/
DANIJcwlzFC6Ts1nzby+rPXRGuVcPriFV9bzkJtQhaRIG76mlrYNt+brhG93kYXe
oO0hdI8ujgnj44bKatU+PHBhXKyIr6W08899H1w4tmiGOaCQIyMXSMB3UyGEVEJI
l30wCQzVszhWvBTSBTbtS+t9abS90X+rFtq1K1Bqzq9Ecf/4WrLg5ap9hJXrMIDr
lH4XT9/8IeexkLr0UyClMPcM1hp1pFpjtNk7QGlw6j4ekOJ86NH3745iG/OU8GUm
JcfQVkvsrc566tZ9KRdriKgvI1FAOkrKfxrFD63gHuVGQCpqOBXU56J5Kbw188wi
NO7wPoqJlKA/OBtBcg244lKSRU1lbz9DGBYNkD1HI3P8z9/Fdhc2OJc6Tqrb/UW6
zksiPUQt4lwIOcEObSTT49hYpxKLhGLaTjSgcz7XNx8Vu4fVKi6Cks96+GRdU1e/
DzOfZKL4qnBq2CE0k2JrTmJUnI8NIUuJaaHrFiNm3suUwg4Z+T3f/o55PZLdYHN8
2YDIXpQvMQfZhcnUEmdfGIYEyE+6umH3GeqfG4NOZvzKz+dnFHXovU2uwEoob4Yy
nOmHmYsZT4FRBddAP06kCDKd6uBoR6LNhb2umPGfy6FuEN0yBJcogXLJ6LcQV3eX
ZHG7EBzLpFAX7VnBNxx077TiZQJCsGATpIB1UREWARM1zoAqlp+ITgWlotc+5Z6+
Bg+0cdW3Yf4Do8nwBEVU8Uua0zouhDQRPVO8Ei+gAqWcvbibGaOvqtMty064Em7z
e/FWgxgQWoWWBq/0lKMSfcXdFxvTUYR+vkYaDF9VJtACRwjQbADqk2dzRcrk1E4K
qUscdEYXwGuJzRQ2zaxYm7FujLP5NgPA6F3ssl5AMlGHnrAh7EmHhpuLqV6YPQ3p
8ijSP5iOmyjPDej7dXTM8weuQVMpU5s7hIjkNEj4D9LF2WnouDOmw2ZIz3BJ/vPA
LpdWuLf2Ko6SG0igLPVL1y1XgZf9HN/9buSCiLNwpIRpxJi9ZkJwR4d1J45yPcn5
4JQBOFl3yQbfxHvLdjU73FLYhUa2f1VUhLRCuDH6mtldjrO8iwvbHJU2kcSfxuQE
neIxRhTtCrDYd9T8GXIuEGif5CFFwGq5jcwbg925Sw5xT2m1yPCMLZbaLbTAATHK
P0XSNMi8A0bY3Ux/mqSpRJ6TY7xINoYF2gmMNb9LuIvntAs1L2uJXaG/7q/T6yFg
NGQTfuymenNTU++PM0/PpEmOOBRwMGOl8ftCAo0SmrJHHF0zs9YQhiXzboxJnhMD
HbE+5yInFJFtBepLUl6P4BJCkWq2lUyXNoVZmMQxA5a+97Kx6aJSGhGxjHTB+kob
0gYi1cgBOBqtpQnZBD0SReHIlHyacxxOdRtjFh2eES3tdG0aTp/SpD14NOEP6hpY
LL4CvnNT/x9hTNczz1B2Cr/Vnfl9U2GwWc/SzuueLvZ7uXCPr3QhZ+Bahf/tcOet
wQ0ttF+sBIB1PAOsfgGdhRqSIEDiufyBGBB5A24Vl60GxzoOenNhnU0lBBeVbSu7
G/mumSQTmmmyxpVmm0taAVPZxMZM/hr90WmNN/YjJkeL3lxg+JO1lvtlCLL8psZn
slkDTX3m9KDhym/EFdqeMQs+uAUzX4Y7n0J6EL6LaUyxZt/VzurEqK7f2/Z026ln
X93Oekbq7SCkcQ4DSHYw2sPVl52isrK2RMkz8PpkbZvEYEcSYwQCej7Gi16r8vl6
Emrfb5J3c2wR0kblsupqY+IS/8PkzkLBp9uZmc1S8s0K/9RmkCIC2ysJz8kop2ou
9h9N14afA3W5FfIaOun4pirh13XwLeJzlllgevcxr+x1LxTQLVsQq5t04xX7Vupz
ZBLDsPn98wN+c87zDIGL7RqbgltZEsyBVPUPA2fNeo1H130Jh4aWJk95ah/MoXyP
ZnKyGYqlnjnyptk+wHuuMJoMYYTk3GleyDdDRFSaVmzBUUu69eoPElc9Te2Yjv/g
ApQPY+nvR4TsrRg+SwbyF2nggTVFrRamX5WNisMWdn7eOvTMWAKejA8VeeC5wj1G
YpeqaLvaDJ9sNZ/WUXYRbBFKk7ThgO2Y0SfXHshQtyfVxjB61Vo/UH9tE5T5mSOT
LXrWpN248o3owePdW3ct+L3H092br9wD2xJr3MuVKONlkTTET3uUiVItrz11YN2F
tBp8g8Pd8TmJd5Ne5+mEzau/wLe05sfrVV1XKIX9XqRNyEnF3XeNYEwXHPwSjtUb
LqWz4Imla3VltbVTJcCyuUFT89ep4TWA+8/wbyKLRADkNa7FcRXTbs+U84CiozJr
eYTaOt6f8k81nTCkde0JWA7ydynzXMKWQSghBzF75cV2VmuOJDKnuUDgjOharUFY
3O2dGYgwB3nFZIttSrX+BzYjy6oZ1md1j+OBG2gyh4/+RrsOFJ4bRL4Ya0i78Vjy
mmwWiQCi3wY9w4Nuj0S3JtBBcmXkXjqi1dB3KJ2k+wejvD0peThZF7Y4zm6Aq89/
rOLIOlK7khE1FqXg56BwMqrTV0xi3pp57zvyBCJZTNQHJqJHDbucVooJ/AcY3N4N
mK2cgn/pxO7NLs3qq7K83fq+NuXxOI1MLLOUO8b9fdprvDBCsSxm7vGHQf4RWZ3s
BPOMfTeGFh3NMf1QYsqLR3MhHAiGIPSXg9/JVQpuo74sP1nPT0tYcI9ZRjN5HxJo
y9FtUJVJypnTiO1rbU50TUhKH7Ydt7QPCDPBpC9nKxaldN0S/ziiEJuFTVupK2oL
bPwbUMsgsXZvSSVh8rFoRnQ4Pq87NeNF6ewCSfEAIJF75YfIBAxrLfrp3Czo7VJ6
nni92n3NBXlZ/Pp6/qbuCv0F1tVNDWWt1oF6aXgFy5iXZfag/nZP+VhI2f8Gt4Sa
6nVyv76ENh0UMYCrRJg9i9BIyjg/Wv0Y3fTD+jXvkeEIFXUY75qIGMSzQb0MdooM
Rb5o5e1oZFQpwuuCaIRApTGT2mMAAuUXY2y321UHTuX1ENCGoJlULkDAq8elyL3w
ZsBz89U9oGKSNOjWNMfrqLbiPuaUJcQifuNios/wYbPZOSq+HVAYTxZGgOiibXVP
RHw8qP+6gw4ujwBULs3n0ra4kqPeXQ8VPL6txA4t6CZLsM9z0CjEJRn8freDQbwX
aYypQa8WPkyS4yeKmA5SIvqGiCkGZCvAuIqYAiiO+JCMfOz/T2dn///kDEyiASll
4YYFsI8kWRUx6nudKFy6HhFB5gHK3n7Wx0AZT1CCbt3Qp6a3fSdFuE1cktyU6CSS
v9zHM2RqnhWppTFZH77aapkcPJcVODVTAnUtxyu5EoWc0vyXtx4DTyXHVdAndoLF
NgonwkqFHzlaaqTQOFBdTvi2dIhedLxBz2IxW9JdxYCwlj7xY2GiHuQmrlwQvU2I
mFeD8KMBo62vn35IOPmSRjkK3wbOL/hoTqEBob+1ePdVvtNy/UthGh2hLRX51nrS
fXVQeubCzI1kn5gA0+pd1t6617z5m8kAe7HYUMk9liczV4TqCfEwYkLn4IxZB9GY
WDwREKWQSQMJavKNYa/4OyXq4a77wIfyPeBQns9aPtGPRx60sxJaDVh2nn1s6aEA
ju3ZEuZUapb2+nYR8HuW25Ju1DgZGLbYxFxhEXglMcIqG3lwP+iKq8cgMoFhjkWk
iJ+uIpXq6Xq8aOh9C/C9s6sEwRqR1cWmtvzO4YCEIplFxFZYo70qeBK//9dh+oi4
b6GLXUpDMtlNJkcJzPaR7usdx5OgEhJMcq4Ns0ucZNsLhv7wkAXTHa6Tj5mk5ByW
naqGcOrUPjfp13LZEa44l8Xuo7feU6WqAFc58ch3SDXSu6y8wg3hCmwJ9zbbq7vn
bmsPJRU8qqh4cGhuyfk+JS9tBBPy/nHLgIsYx1b3acD/O5THVr8vrsmprbNUfKV5
GlPlZsmolgTWtrTH/0Vm+ZnNSzMkzrdbNim7gH14Do6f/ndYsVABDen3uxzZHLQu
xJGVIB1PE5sq6RhGBZ46sXqPi80KmR6nJflMa6lhyo045Hl1y+KI4W48LHAMNAmR
X/mH/vyhLTSdS3LEde9nB1lcUo5gx5BHUV0bxxfB2C2J6cSaAZkE8Q9xtxPnhOl1
gRVa5T0Ab8sGOoCGWmBcmpTnipMjGXIYPfkVeaImC1zBC7w/rw2p6uoKkuYxbvqS
bQXaljaRU3GMobUSl9GHBzQdDFNmrZmtwfDmxi/SsMuUIgWQonHmWSkoCu2grVQu
yY95wKEu6dl2VoUfVeDk6zZS5XEvCZK4gMH4ypLHFn8UaUs5Bra9btPGC7m1wMqL
WofcqNI28stRpcMd2FL/u7/HgJ2bjFbB2aFjX+u16NE3zsPVqJ90lTQWo5h6OMrV
TbVfHZB/T080Lv54sNYifK5Gx/1ns5nekSHLsDh3iL48AQ8x56ZoKGBTwaH/26h4
N2YPdEIQ2366Gz5n9V2DvPfW7bLGJ4rCm5gWT+cvLw+9H9QVpUSX3Xg79GmYin2L
jHFvz3xV3fcFeS0u+T9TfL94HmJVBvdsPxA0d5f03fIhX7FZ/CQbECTE0AyiUDfz
pXRIH0+QpL+kAGBHfraEmfJFvBwoeAnZXA8n207iLs/SDxUpQRkDnsw74+QBxiV+
clHN2neiisXGBSl28Z2LQWLsGkYsjFc9jv6SREnXgr5cM20ecCCg40Cp0afF07Oa
KPbm11psfi7V2lMzHaOwwBlGKU5j2iROXlbhHSGEzCvyC2qgAT22LtZ2nlIfK324
Lij4nUFAhvuBKeyJroxVr7FRYLtFXa7ISKYu4593kVfHohf/KqwPOVlbSirWA2yS
ukQ5feG1x4ekWfeZHn1u9pX9bmZr95HWSVDKmrS8XjcZncBmJTT6plhDRyGSYKrg
3U9xqhnMxmQoVL+7JmjnKmbaSDkY5pADk93YFn+uYP+jLVRoP2RqgstTnBxffD8V
yH+ZimTU7Wf6ueAsYhmoN+41Sh0w1NBoDaBGlduCJwQYNEn8z0nHm4AJcbqTArTb
LWeFlQgyQINKjL82BTyQ1SyF1CxKgd6KdY+Y2LV0ZE6XIh5VzRpeLvfRF9YU3H4+
aoEJ4/pe50Gu58oRTkgb2w35p/M0rLhM/JanBD3QnhrXUSfBUGGEcHi5dpCc8UJc
oPemkfEl6/dzM7BcLpae3dhuSLMFh7uar9UUYTuE+5g4OOivjyAhc3XJ6GFqYv1C
agl/AMH/2oM069F8k3DH9o4AeJRyc6yyV/TMbfJrRLyur0bzJcaJ9uGFH6WQJiwL
ALI0SqQtuNFUc7k7NCUQ0EhAArR5CxFNl6yfAGlGDoV41MRAmbtDWkXMlyIsn0Fy
PaqqBdVyRYDbyuxr9ngN6NkLFP8/dsN6P7lShhc5ApRpXDTGYoHasH3xcQcfVvLh
YYDAVegvrfxoBTlXZhR5ALY38vGzQx9/KTDa8q3V9Uhil8vXIxZ3AIYAMxOmis1m
DRtLkLoQyEJBIvnIk9hRCW5CFAT4NI9uftL1ka8ykm80qV+73NFyRtg6TphC2LY7
1ftiqc2KVkY16obGDBNOKJUJ6aoM2WaVthm6l1uPdrPCgN16M3xSbLtZxbasMJj1
tFJN0dZP+ORQNfC7HD02vSdk9H7AbVjcj4Vy2U+Tna47TocfN0ZzYozTPWe+EzUO
55evXLTc7FzBC/XTrZ7mD4c7LiymzIhgQSzxa3oPU5kWHrrwqnsGrumx31+CKSPE
SDWJuh6YqjnbrhvXCi/H6U5Ajfg8VVltlKsGlLNm2MtmCTR8v1wFvDJBsWaiga/n
HCV09kLKn/6Q9iOyVgas+TZjZFAE60g91/FbMNeT6EjYKcdHLfusfrOnf2+f0i0O
P5Nmql9eAgGhUEj0X2kfCD7s+S6sbNhjUaFWFIrjb0URsZOA+HuuF/CteW4R7UQL
gkrhBThBx613R9nPJ3LeRtPRbUj8p1E1o1218Y3OrmLdZPeZu8RouNsuibUW7Wkn
Tv/BTOvbGiRUClCqsOr/77wg9IHt3JfNSrlepe6tsKKv/QRNigRKZkjGzJoWb1uA
JA20jqdsSVMj1FDVMTEezrH0uf8nuPZHoUoW7o8QlWeywpgk5Hr7YNI1Hmsao8N3
VRK02rSgE7oaBnzbi+kzsiKhIL0RQepCoaGEzYHZdWC1/W2ZMPgrGx6QUcohyCc4
yRynBRkIMBOwx54UVWapDSpBPvq2tstDfJWFQdQ9F6E1qcLWXY+A3Sqat9QTDsQy
QbHilgC2kU2bQVlFDsSlYkcUjE1jLnxEk/rZf4tha4mJpbDYe8OhiqlVvIxhyv3d
2FPSdB/aFdPnWYX4KfQkfFU43Jb3MEP5Z3cEw/IJwDmL1VL5B3Xkwufbu5BNiNXK
fOVjSQwK3KpRUzl4f1wWAqJmBjD/hlkxgxKpR3lqHEJL2hLYRHag4FYTkxKxgJtL
oK3TYyzGCexTBkAslhGcfhVgN77L4VyruV3+tkG95kSaRcmdaZT1t0QiUcPNwOWm
jVf6hQz7Q8e4oYLqEIg1iDzG0nteBdJvMqlcEArkY5+Ap/NzLVpBZudfKO6VPHYt
NjqLyZUsgUl0R1ZZou1vR36tGyNGu0oqlSMMyo10jAi4k1PL5mVxQa4YV68NNTsv
Zl5fiPBuqmS/iUL29+Bk3/auTtPsgJbuJvg6MsbPRx/ZVN4DJd0Qi+e0OYGKEm1w
jsxpIWI7kJUlJjGht5nCp35RfcUu5o+u2Kz9tEKG1DDAgNTOBVLWgBzA6TYtol8Y
QlTqa/cmYeK4doQlUX3fRiBgKcXdXcRJ1kkJQxtZfzeqyYIi9pv9AwPrLIbFelMH
TG+5DaXvUEVh/pYK8yAdxRw3jcEBrJiXc8Xw9C/gQzCJN4HnyoXKhhhFrUYp5uAc
FPGU5FCmPy4LjcdWwHC/+S8XPo8t1qjOm+wjSZbM1HQk/XK263XjyOhSvcVPR+30
4I1T6GZEC5oa/CFALN3SengdXMOnq2ln70q7gE0usrWursUMi2fnfF8LK25/n5VX
0Jn6Ifx93safCsGZ0R5FhLTsXx0XJ5fa8/GXxWsjfVxbO3IMCfTrsyuHmTymo6Nq
mo+PWfx0fazCu4fploHw5crnsMERjjLWVEq1SKj/7kD/gnBjF2rrWDGid7DhFMk1
SVyBWkcM6RcB/AviO3GWCuO59XiqnBkEFOPARJnMNbxf3TFiz0pS+ei6c7kdn6nw
zlzbToZKrMSIsVh/a8l1kqiQrFu+HTr1zeLYaiw/p2tdVWHP+dSX8GCnngpqRyYc
An96a8PvP4RGZnhX6q7LdiyLDGZp1SywWpEsoofN/Gj2wClmyhw71ZewnGj2MSWo
4CHdxmtYspK/43Fi7npxGEh/pM4tvtVSL3lK/4m9r7d1ctgd6aRS5KADQ5V2xEWh
wRxUxoLjKTQc2XU/VEKVjXicxNgfu8dLrEQ5wlwSvPYbwWo+6OVNqdT77cZIO9mS
ZxfVWLdteeIEezxX5HqqYubWAc5JNX7NQaJSOeZJuCO72mkJdlmZDhpSYOCOV9dX
Cmvgogdqbh6piwzjh638RHPHys4hi/k1ruIG/f+HeLGnEjEoXaMymGWfm0zz19OC
Ak8IrGJMkuCJJg9WekewQdJF2J2GBdCVenVHCPJvaAjtSaLS/BF34M9pwCUrUbtJ
2FYSZusZQ0LJt7GhRKTMmCkOmnWYWmUaoA2E1BBkL4H2K8xsBbI0wqSDnDmevBqd
VyAriwO2yfMmpdvc4kvA9ibXNWMwUD+ZVogs/od73du/k7wjggNyW1zlMBxoRllN
4Sb+iLuh17XgvNUGD+WfvUlqW0uyJ7Sj1LRvdwivbtASNnXSvSgBmBpFQ7OXweaU
Twq52oUu52Ah5hMq/r7OlF6Nai3ijxuLo+vsodFWmbs8mO0LfyHzmtjeb7hxEGA/
bgQf2OP8cxh0E4J9DKcGQeZDN6HPG0n2/7w8fvgh0RY+oyjAy2jQvad14WALN1+N
6S6Bw7nlnNFIYAqQ9FKBRj6NoyNSZ/GvWX2P6mVzJWbwkXMMmd1xVw7ssja1ygkp
plLRX+iSQgJOVg28qedmz1p+FdtVaRRz/t4vbsHWGO4TDeL66qXEhl6K6P6pi25a
Y0CIBZQwlr8R/8zs8HzquWBNcXWZi4jYF+Ids5Rb+3RVyaUW2v5Xi/ROmnJK+Q1E
JHEabZJ33qzNJEDOerwTjZVoT+/s1QUBaXlk4Z57jqL/V+TxsHThiRUgWF7j0GQy
6fr2gekajGwf9qoZNTPGXq5yesjcz2ydG+SIl1JLQjcy/7fjt4LqjFa7Ey/cO2qe
BTJzOpF+zTok18WMME6IwwlkEkki6m5cpB1IA3YbEBmvrZj5vVunG7a/ph3mLEae
K6NuGn01x6voT1LCeGelMn3qpI71u8ur6HaJ0tIVh6z61GqJlf4uS7keMZcQwTyF
SsuUIRKEykKDnuQXAbkuAidS5+y4MPmBw1BiPLphH24eYqagFSobtBANxrpR5iq0
aWIJMpZEHilYtg88pKRqNQgoRY3bT7IbfD4mYwlRW/Y1OQCaLjgXO0u1lcAsk6Wp
JCNxkL8fK6SNT1D3doeLThEKEG0CRudecWh9rp39PHWLCrjyr/i8DcKfdxuwx6IJ
fOsdHsrlxeM4zrY3zpIoFnOJlnMwS+Osc82jrpowscb6NItp2tegoIDTmeuLJqFH
mKGmcGjWSrldt+7TzVvRSxrJl2s5YdR1zhNXfBFWjEmLCVemhhoNcHR1DTLuc1c7
MPmq4NDDCmBMZqmJ7wJBn0358DPlfPeqp3FVVagPL+rsTJUfePqkqASSYvXEKA7R
Fh5D+jATkzu57qMIl7GEsCiV0hAJdQWQCicVZMMRYmLJZsXctGK3ajbefT5YbPW5
71OOCrXZkzGPM0R/wk0btjZsj14YsxC7GzCtWfVa3xRkr1SNaE5T63Sy/1PrYX61
y9iwtWekog05fke7uHciew0dr9SGlY5b85dQjLtQrFfy2Vdk/+vB5m7Hpli6/WnE
CHygOxrq6XSgajI+nJkACHQL0r9f8qa23Bh9fpozzNm6gGZjXY0Jgm0VTLZOwiQn
yxNyvcKbstQzro1oWesoBb/vPTOH/WCEJ54Ovm98gFBG4klqHhr2r853Ead5sEQC
YbOFdyb/RlUONDgRpdt1HgJZ0xR5St6pqPQxXDI/6V2PJjpzydzFkI44Dp6+JP/h
Snft5GjntKx7C8UIJfN3KSPwuPLhS+mMVURgjowL4B4jQleqfI/ZfbK32eTJkrZr
1XbY1f4caUZjZfBhI8nnr0UJuPBpWJ+a+s9VRCIlKhiLmjf7lA6dvIM+e1x0fBCj
mr8BJ0nKAr+n0YowZkBo9SQEqENxt9prMeTG6ALw4KqOiEMinn4VXVs/uGZN10rx
dY3+t5DsKkxRqRqjBL5Wrj9esz6SXFKlLd9A26BIv1v4btYTfeCQQ08zkcjwn/1h
l7f0sOvBElXOEWyHZ5klgHIDwQzXR2zdNjc3ngjHB67/VDZ0B+MHNIUUzDmYYG/S
qhAlbznXaM4A4w4K8VEZ56gNtKATh+v7s2HhhTN2peQQQqbty7vOqXkQYQpivNi4
691rY6158H/qO+em22aPDZC8mHNxvpvIZ+dPzqzjl0B9BAKcs460i+xH5QixywmY
jwdWYQ1WXUjoH0tsazybGR5jBbgWfJhKPFeC+a9WWXqs2Ww43dd+bfxN4xq9Woqj
bOyoCVsZcD1z+zdMfksZwANjKDZIFSIqq273NyvD0c+rDpU/0SZO0S19hYgufAmF
4jLa71xsnU16AALleCbMlg0KhvCt0wK+HK08VGpOnzCJp+yyUeI/qkWC+OF/Qfu7
ERLlG1hFGgzl34x/IR0n3C/tuD9cnLccR8/gWrgrmJMlbTnKO48ODTmOyA7y8tk9
jk7Idw/Jq5JTjv2ptqMoxhy0nX1KrHMTEm1Hz1KCNDbjuft+cpJSiGuosJUGWZNi
T1vvVF8KrT+7agwwi2gPorKbXcDIC4GqCG/nkqQR7CP+6IL9nchT9vBiGgDIND23
qEXPnxQ3qAWPKVQiLH67GD6jPwiJvQly5xhPhjVuwowYA5LeUw2/ac9Onr6YkGBb
KxRAHkVEkdI3d6PXaHV+rBJNRzS9MM6CEvhsPlBnzUnLhb3BuCd6b81BKcSwW0bn
PYX+GGH9en9KTPS1xvULi4XFUf+ymHj+HK5RB4SrnPnl7qYDgU2qOs8O76g6ZPS9
ofPYK9uyyQ7uAX1hY0A3uMEUiA/qfA8F3aSJt1fuNJdIYVxLntez9wBRk11KK0M4
ZrxRfq4hrHJWlU/O2v7c7EPdpz9UPvWXZCG/98MTafGu5aaN4i4H2Zu453/rS7rU
bdiV5RyyObwECqrGah5qelwbMA1NUGQFuh8CXJsqdrjan0J4CAiAgsM/Mv7bnHEu
WV7JVB9/hAdZvDBl8FuZxt+tcrYf/JRjEYlhmqNo0CfZOlVkL/aFAfjV6ZATDu8D
MzZoDIzFM7cGlwiqYN4eHOgFIH7hdEimHFyjGXf/zvYb9WQBIXDGRrpwoQKVpGH3
HiBEFbWN4G1f/lFGKFKA91dwgMKZ2D1azXAflmhZ4WF+xuE1Zc7OtX1QZ2wvvxMh
dNyh5KCyJmNLdmGf2rdhIQIzArRhLZbpo/+wSeiTvu8EKke52KayEYQ2G2d4nwEy
5VQCTTucIRtvA9GYj9ULmTG1ViXs+m6erR/GQwDabye+zkUMk5V1K5bwUnKhtm9L
sUqmJTsNOq/FmfYgclfq5Xr4vBtm3QXFVNOq0cHaSTTSsSsB8I7Fd6nDXPGIWmR1
JeHqbLgYTwepTa7efa6R2OL+wl7fwzAbS5MwgJaw0Gj+fTobSYcJjYFNum+Jx6Cf
221r2vPHEUNIj4V2d9HaPf6muDRvq8skGCfB71kQKxd1lrJ9M9xTUBUuGXCeHcff
xtoXK4gAAS1qbFeyWCSUQ/qt8XH1t3KKvmLClE4ztuGEc6BiCtaJcnAsAwsuqjTl
bNt2NV8zCEqEcx6KISyBSxEf6u6hqG+j7TrCEgkv8F1lF7HhjDL3Uj1YXOT4VYKY
rtegNJCFuG5rFcUXm2+TaI2XUarGhZpTm/ZHqQ16nYfSo+5TPcydWtGgQpJC/h0P
Cl09x8YGNILSnU0rPqa9iNMEZcvQkUcp6fml4CsQ8OqgiuL5bbRBBXKD+Hvg0qsa
tnOcUlUZAqw/iMXB5gZuypIMzC7/VxqfmlDF10HwyT/9QOIPZOGLJQLjvNi1FmtY
9rPhcgkiS/bfi7pinW8tWqyPpl888GQqCe7l5zwOPgOvPkvQo6En0Kxe2SkbtKld
qLRLcq3KlNuitbzOANe8rWe0dZQyy8bgGYm6JzR+ZFYPls/a7bAy7huCqEgiDjON
EAiGXp6UesDjzGY609RK0xS9mFkxf4UEKRGo/+EmFRDqzYqbCvtKzAITLiXHLOXz
hzrrS+mbbi6FjVcncm6X0DHtOYRUHvcGS9bXfq1CJKdioYDAUr8OaqfSlwmqkiyV
DKgYPd+pbOQWv6ajbUMb47rU7RRBEbTmu9eefdz7Nj5C1CG58SZWV2Kx9dE1Pc7l
QFXAz2pq5VccvrmeyLVi/HsTv72cCTTMINcxP1Rxx6QemliIETmjACmsqLFzPrF4
V4b84sRayoq7FlFgN5V28bWu040d1FUAYUw3DBxNTlGenlJftODlAMAcm9uquC+H
yz/owK3K6x+jRe6UhaX/kRl1f6NLsAiFYAAE8n59lLxeaAgjDh/qsklNbJI6+xnb
6Z0WBsYXJCqjv2NPMABx4H0rb37KwIoNO+Zy+5N9gTAUfUJ3mHdJ339lITDeX7yS
u4DFv5aMzZjKnjGYvYKpxLfjcCIFdNEI23M/yLncYGnMIeNBkofFH1r3xqQL/8IK
CweGPT2h0lvYl2omRqt+AgyKwIKx0wLHTfETLCfSbmhpDOE5RlN5ykJoKs2Evia0
FiA3nBwH66X2thPXfoHA4+r/36wWSElMbBEJHui3M5zmI2Qx9jWCPXZmSFCxminy
VHae2NB2Hs3BLCNpqWH96vdhzOVcU3ZWTq7uPdKK4i2cr88pJch+89W5+m4lWB4B
CSfevKN+jABGW46nXC2+sXkStlaB+1ch5cv/Y16jMZ8GWuXC7ZOispCAJfLFhtAn
wGR7xyen/DTkMHl3pED6LrLC3GqcPMlH/PHum5ljZPUEs/v7rKHAyOYcUFx+siHM
3wbLmskC4Fp74zJ93yLluQb1dCItpGR6X3iTWPjDA5yIz7Qu5sVEFLmnKiNl/uNg
5FLffsM+5pPayduLwU+Tx3asBkV9wpImw1Vo+TYS6Kr/WcdGrRa7WS68sGOAPcyx
i+ZJgebGvRqrAIUmCBEmYBJKc3BGsaduviAAQ/+EntX1FPr7LHZIHGK3grm870k6
PXG3Pw+0/nIoOYDPsBvCmcs9v+9cOKB/zbdVpAM61Y7LvC1cZGkK4R27VhPyRc6x
tKOIwf+YySoju/t0+F0PIAplFYGgDLxhODjU7U7Dvmed6jAjuriTSNv5ZFuEW1np
lSHkDzxSp7xHthQClulL3v2xYRKzBp2ZVxqGuXcNngrUTwKcLYDq+vcW9aP65Lsv
/ncs697Hqln5MfImDj5BjJPIZfIfuU9BbDeOSbs3rEJnk+zDRRhKB2qEhRgjiAlI
gEort1HQhb9qNYtJyGaU1zvFK2LzJxJH656L7Z4M+tlkF4+RbaNypD6cc15sqUTE
yFShwGfKBr5Abc3EgG7G3hXRtBmUuZMZnfYwRHpIa7eiM7i1IV2glaG0TVmVYKc/
3L9KaozzM6vsvAFmuGnQ00BmwJJW5O8tNk0AJ2eIeZsgnv+ea0cEhCdc6TxnQmVF
3n3g0l1BdAaknuy88+5/8yd5ahTI00yV1fwlw7fira6D5LkL8fwMCqWRA00CYvDr
9jfoz8rwLxi88HKmmz5a2CNZ+bfqL1R4eeXIJiPMPPecdAmRQGpELMWWlCNxx+fn
AdE+a0lM47C3MhzmTzbpR3Ilkf7+jvf9nu9YJvLeZO/Z43TTM8pl31sBDHrqV1nd
bhPDLx43aIFSnmpUrCLPWAdBYp44w5pmMo/1kIYLWRm724bJ0QsOPnsYa5F1kz0c
o+fVWb0PnXiP5dMOzt3oOPvN7+3S2tjlM5rlX0KOIHuatgjj8P4/HiWDmk8WNCpw
jQblAe0QgvFmX9BFsWmvwsBwGpIx/T0rKLfw+LgyWzcXHl2WLGUijlEV3IGTdnYB
nSsV0u6B2iE7UOtyuRpldMd5CUOse0eL6JAbhMSAPesBsYTXVTSAwLEbzvOvx7dJ
EipNJ6GY5lSRYfJq7OBTObgW1Ync9VhTSJ9ibyKXOpLopiVhNHOXLbqZlKpsH7F2
BJeBrl2MLgbWdwuacCrO1r9p+2QCt7ijKLyxArTEEtv+AbM46f5gk+KaSPuHBUyR
ZyaIPzqGIPBq1HNL+WgnFEgZj6fx1fKy39x07ais+OQQv/EFhR52ve//hyfRIED3
elqYpItpnITwzkqy6Gj18l+0n6bUqcAJ7rLXfqiRHa36aSzp6Ih2WkhaGUGdlYRF
hP8VvnHpv6ecOuzdYUkk3ZFTeVRe5h5aogVZc8mYb90pR9pLg2IwBZY/DbF6fq9s
3OttyoEZn1gYlbExwoNd3ywTWLB41+WqVjxQ/3l5PXmQ/4wbPboLjm6lPTGq4fOO
upBAk8YDB5CYmiJDkUXzOC/HZg+zioU2s28md9c8vCaB6fWxCgtkeM+H4CJtuhme
SEoJPttZG5XFFqPNJaZcuvL/sdEdvFe3jCMY+ggZDwfdqyQIunDSm6qgfHmL/gFa
cvUE3EdJ1fy9sQ/a9pbdKxuub0ZAbfsb59mS8sN0bXAHQR2zhVTKS7crCCvIxtS/
epENKTlg84bTg1V8YMIvhZ4al248yHxromOU1SyRmOLoH61fotL/QutQO2yaWHH5
QL0K++ff2XJeKW4F25pJ9F/lmuToRmR9YF8Ycq3+tWKflEWsc2XYKLXO5ugCo2h9
IMA2HFzMOo7jBn4lJjY2VOmKiu7dPnUfBkXOlYtTO9zAYl3dhSM871F2o/Eopyh8
PZ0iBuSPoOc3NRYT+rcK/JqCr9HoeJdEzJo6SdzTyBE0lS//fRsAyjuDjeGqNtqR
gvTc8Kr756hpY+NEn0qng9WKyAQhsBBbdOvy3E4a6jXnlrQUX9DphcLw80k416IQ
LZnu8qAToFXv8kiRh+guAkX4jEvPnZN+vCfV6Wdfkp/EDcwadH/MsZqEp2G0trzh
wtyL079Y95AutPsXWYf+9QAde1v6USNJLJO1xEVQH57SgGa3uOFlcwjT9n/5v8gM
vpcfMsYwOO8q1/JhBQPIa69+8PGqpTZo4tVod4nWcLjw3ChZDVvwGdnXyTvtF5zv
VW9x3n9nLakhCaHBD/ZXTl6Kp5wo4VKWJKderFstKCvU4WckQ29Jnor5yAiWWOTR
tYSH3QlzYHlTOPl+W9sK/Hd9Ea+KGHjwBvbICmD+biJGCselBjQqGvSZTZrXYCNf
e0J3Kiil2qkfJbxMrEUkPrq6AFtLd61gYi7PxMv8sIXv5JI1mrlDMyXOXnz/ipuZ
Thb2TNSLELn04NAITk3+hAAKQCeWKY+9ylcWA9o8BGOLnNS0iBivpP9O+1AAMCuo
VRfYk2l1PrjfVCopABziezApLfCa5atHWmAY/uLI0xAn5znPSbzEWZ+SnNLBUc4C
LlmsTRZZZb0hSn8VycuhrqjaSqQqN0+9h04I/Fje+F4EGBpEvl5yRQ5iAg7TXT+g
4wjL5g0Y4W1ARdT7bnWAiS/bSjiduxZQ5T7JHETopLc9BrlSU6uZJQd8Ejy8bq1Y
+ONTVaVxjdK/v4hsKtTOI54t9FhzIKDGDgdZpCb8+X7ajlxkFeedUIFFQPuDlSyO
BfqVUeSEgtlYcKoaz52f6lB3ORSqOlHEM8kAuySI5Iu0nFh64vEHmhQqcZbQaEB5
90Af/gjaibzqQRXD0KA63Jm7CTtumSWJaa0Ah80WWOZKq8j8KJw4yRzlOMAYVyAu
uTqGsllGxbP7bgBxqrOENfZ18uRrUZkCUxtsXUeKgB/WpXxvm0sx+G9sNAnjG4u6
GhV0BuA0xmC1QiYeg0T0zm++D+bnh9cIpG+HX9VHm8LjrBJnPMU/H7RgwrNSFuex
dH+YyLEPi7W3LBw3l6Pvs+uoeDuA9j/KLYf/rBLkrJBIGsvz8F9rGfGSCDR3aF5q
Xeffrtf9qPkWipkJk4cz1ekZnnt6WF7Y8ljxx+HFvqWMyZ6Hnb2KqVXLhh/4aePg
LLKNtLzG/UQ95vj9cyixFuJLL4cxoA7KXJvwtUX4tF+d/89yePGlI61QrpbFwhKX
MKCBC6AmxykhNJctQVF2SBfNfzmPSHk7dJFqHc1Bvma8K389PRHHQo43lVb2w1Nw
iu+ddU4POMDZDKkT+7BtOdoTe1oy9qiSPp9QVUCQqOujgAcjt0iM1NWIRNTRJHbd
dgRi1rsCxVP7EhKhNlYesehxKU9HduyuwCEIU2RMzXU4SKPGb89JqwOzN5WrNrw0
C2Lis/jjggP9UBeXgpEBk6ELWuSPC289rZeXyazww8MkjWG7zyWBxqZI0Vhca+Z/
8QcTg4YRpsdF/X62L7UzV38TaU1zz/N6P6/H0Xt3wGcm9StjnncdxZNXu2wOBwJp
qsp0G2F6pH2+5CYfrWLnEkYZdx6LXF/bjH2OoMZUDGcf+rZFJMF0uXQuLLXDjld3
m4cerni0J8NuvOyZwhe+zJ9K/SEJGYh/2G+O3a4BwKYLdPb7LCSukJJ+JrRNuOe/
yymKElJGu9BGiYuWlmS8kFTxEA0USDysA+GjcXCoDVkzVs9axdGpCnqsUH0MgNjD
vffE7LlbycxLAQ76125GAU5lwFu3xArBeaEB5tya6dDEW1VJpTv+KWCpZAjgctcR
PFPCXJgaSQWgW22F6my6IrKi/lHyjlgVV94p+Fk5G4tR2ZR23qM/8nx1JNAQD2Kh
P5AGSWeRJ0W21w1STuaiTxmsE6khsPCu+bhgh31JQ01OChVfkGMuOgg9Ivmnqgrs
5//oimlXzmS1mPdQ9bGS5wtoy9N94z7XAxCYl3i0cO2y3x3GJF3+Yg2ar4yRDKY5
u21Iox+KFT3t5NaQ8uhGXBLGNZtQh+NOUFagdlDNf+Nm/W8AHBprfQr9R1rlLt5A
wmRYzvpScgafvcRfGG6rbXUvQIN+vshIsicogqxjjUmvpnpmDe3Xlm898E2/pGYK
VsiPKZTLlxWGEKmdK8NOK+OO37SvWOKPfQKTLBmtbXATRNwAqnG2l2yHpEL/7kN4
MUmkl1yTJDcey076sxMsG6BfatHc1KvL6+NYK0QW6J3EKOaXa08uTf3VdLcq5ghk
tyi7c7DlHB6wmvvn2O4DV9Zte2d8muBnd/zDIrcYAT9h2KD9HUka15AZ9rgBbIYy
rT+y51Ij2ZKk3omQaml51eYpaM5Gzz01ute2wwBnLjZly3AJSfdMunNz+aUxI7ln
31QY9OcAhlQjiBLHt8UKPd4PVeV7saX7TEsm5CGaYEW7Jdkk3kJ5aFuoYxxSkHOT
fwXxBNbvGNVdvuwARMoKprELgnhReDzGbqVQAeJgldtbcDVatytER7ATDmm34spn
Rnuz7fQ7sagDlkoFPJYcH1QZ/IfQAPlJSywfCRME4R9CEJrjAeI4OIMX2+q8zXaZ
FwBsmeyMRIGcvx9gZpQiKK1lYT/cwU9qelJeCYDqzbHWf0w3hJjww/QtvZYfPwvu
OGuMTq5MnehoFNbwnC+2yhf/bEYc2XouIihLbOLcX/Rc3FiQ7SoSAfysgjPN1XCL
jySjDuTRxByAzy40CJF8w9qEWVEAkmauVLh9+/mv0N0GNYocCXMkwt1m0h3W7po4
sPP2MEmrIwIKQgNiqL41HyZKsjlxJB59i0mwfKUkxB2NJDmTEWbKXNUa+VkOiy+q
5oi525NslIjmLWjuo0VxafHOYPPVyOZf6shmuu+vZfxayQyo74SXNQiJ8P7/YJu7
paWGe9EpsQvUYkUj2yFFLS540YJkRnA3Gr5grKUtFE0q7ciEeJD9cIDUkB3aBcUh
xsTiYmBpy8/Yyzn6ujuKV82Piq69Imf2KJ1UKmB87qNgbsF+Wa+B8+5XBa3ptQNw
XnYtYxa4CC+7npE9eoovF7GqS8E/ZaLMs0KJw7Vr7Uui4drHUHyair1Tw8bfWFq2
WOOYtXzSPRnHRWboSa1tY0FEgasBZ5gsdiOJ5OK4L10Q+YdmmvdpLiowwiHDvx9a
TZNucWclGEcnfUScCUOY1CB9qUAjjTvJfntv0ZDrMkkZC0NxXvr4LuLGhx0kpRjE
aw6e8+ka1XknjBm0lSyNC06ZRwcixm4Ed2EpyroLu+SDDBIYxf7Q1AN0L6LTN4Ml
U6Zl9wc4/h2LOgOLUnMIe8no6+VXk6NUYnpLqXkQ2nJnE3rkQInyiYtvqouDRN0Z
Mk0Vf55Pa61sMNFVJUByfZgcuUyi4MbUy2IGo/qJkYpDOpY9c7ipBODZ8yEUOKQu
OZaa3fkr/FfaHuY2UX0wpN4PncfNpXn6fbMttuWnakgbhxgQnseX4zFdlfjw5KEd
fOtjkwDFKBUXR6ODQhK+2QhfWEovOHJBdMIRr2DYB1RkYfCdq38R6q7mKFTdGduw
g+rG/ZDe1NkQQKC//Q3nsgVjRu0+AKz7r1sc9GycfIHRzABQy9Jo7PyQvQFTTygn
bO2DUaFv9BGhMb0puCxZsbkFOy+Lb+efUtQQAK5B6uEhSGqOmDTIa2g21p37w2+m
/UenNPcv/Ss2Vixj0lBmQyV2J4B4CUPhjrjx6Hd1HTwcuRQA/o0YeETBo4ZSYgFW
S1sxTGGpzT017uPuHiNwirBHEEj2/nv/uRa7eU0LoBe8k0cwq64DOsdxzt0Zl2oz
n6B3UhM2zoNUX7GT140g6U4ta02gYO+/JawTiTnP/QdCTRSqnOW2nL5zu3w1VjIl
eDsXGvgJ3TUb9Ie3tyk+cJR3ZHOu+a5AfOewv4GkunJ7j2RsNt/EmbADEeKOZ/w7
a+iIVDaOiCKmIxCM2ZdvXDpBZCQWflcG+e8rbzq0WT3+5cvapDp3zyIvTQfeBpcI
5DT7lBAktkjdT/NkPP3ZA3G4NI+kqgarmimsQF5Nl3Yake3Sx2JgXNJz04V4oo3Q
JGxsACbRuMLSkMLr07dchPtk+ddtHMh8J3WXPs3dEOVHNg8qFUNeKzrtO1hlxd8P
Di9RAPGAVh1UzLTFiAF2iTqX+7BBUmH8G4qscwHcLucYhgj3ZMk16JTpD3auS9+c
hOxdBFlnFw24IrvhZJC0wdtqgUq+cJHL96k8MuPr5gGf27Svjt4dRbLHGr5J2zc/
cQdV7hHsw6/kewzL2ghmPTr1nEtCh7xW+2ZJiere8T4sCtlY7MZtOthuESrYze2r
ZEvc4isohFtyb9B7dlIkx55EVpgUhl8ME6vVXfMYIUrWuIhUZC5lKQE0csR3S4AH
1JhL0Gy0HYN4R863eMH4M3czFUnS+3LMmqJciL0UEmWSww/PTmNXWCIMcpJ8QdYg
r9y9hNkNk5GrJXRbEc+izz+UVBBE2YAnOA5545EMfc8w/MUTF40CW5jWTm5T47Z/
STnOINtomDSdR33kgrW1G9doFEz4Fxkpxb04IDKkc1VmgOYandCzGMPTFcWLv4ev
gbzgEnyQtD/UzTllhsBI/QQlDkVpFS5Arx6qZm6l+21OhW6PHkGI4TlFj8TjCTAI
EB8YvVpdzbGE4GB3Ucx8azFyhcQDXrJ/WXK+GYlFWgqaEdCpF+kE5bchc+bg/ken
RYs8vDqXqMAzJi7puMocHUmKLDU0PZvkuS8v0S25o4d/Z/8nKYw9iu82QRfGfuwC
+VuhG72vBCX/nAFb++lir/Lu4RYcJt2EGRnbB8ECeh0Ob+HrShNZ2waq+D0Po0Ym
Lk+lzHqczQtWJGRyAFToQmKau9VcodSgT7YGWw4YEqdkOwY8kmjLiEvxC/vH4apQ
HrHn96Ojsoi26M6HQOteokdd1e6UL6PGg8iILTZ5KV1KcKVU0i7afUb4V+JVuWKC
SLO0yGgrdu8S34kk/4bcJAGLxswG16wUPLocWWBRJfmfDKrgKty2rqvU/V/FrS7J
O/Sx4Zqe5ZN0skrZ0DbFn3imr3gd2J1LVT9ibO6nhC9Qv6SydnnhHybJJG9okkaq
VStQF2ow7AlbNtA5x1I3rY2xnlfB0tMymwHzHmkekazSsEiBd51xABqvu8g4zygd
QwOWpP1aSjZEBeS4c10wJeArUmgt2ex9rI8YJ4YPzuHZrhuUDQ5iYIHR016z4ENl
6gvu+/Zhv7kSVKuI4sEjPD/t1VTMg1IFG4FEIsN72zVUgvS3oDHN1BWAEzsWHT4L
xkdW5foNo9aeMY3nuveeHaVTOZvjMrVvpUn1pF52KUCc5rlNxIB7Kp8ZwTsSG0Vd
TPjszGj5SkyAFCM8vw4mWHkIMxr6eXyfEDZSAZ2NDNWVLxlTZhjTum9XmICwyT8n
NqekDoC1GKDYvESJ3CuYNo96slpfx4DG5KCBOKfnk/WdowKUrRq/788JGydsXO6Q
F7gW1hjfcJocDesvYxownu8N+t/R5JLGOii3WjmoHeMWqKYE+pl4nN7Kp/4FPeIV
eVBnFo+hf8+N30spm4ZJaK4vMtNGq6rJgJBhncntlFVkEWJ1mQsEVNGKHQmHSGEl
6V4VUBqKbEmEB2qglBKwdnnbV1Tlw2VyQ0ak38qgzKCWOlobUXiODN3tqoVX4eIy
pwIxyzC/PpoojH4rQIZZU5+RXtHgc/bq+7L9lvrUaeoZkwsDEEzFxe0J4Ff9hg8d
wCHxnLZww8xCCI0eZR4V91WJf8yFsZVt4mtgaL3PDIugz5iBAcgv97VVGksXXJ/C
r11EU53aXnABNaktwvraZ92pn8FT71ZPHyXW0GcHqdx8XzKoQAoVAZg1ymNbkxrI
TEPXWvJYq5ukbA6ET81TU2zYL7V5IlYhnSFcZQYYbtUItUF+Tpoyw7zqW0GiRD8s
znlvwxFk2V4K8zW7ZYYhVCaXEFQpXLTBvtT5bNfUUCTAh/1tTwkhUUq4MFaLBMkX
pPkhJjVJh0uKW0rRFC7Qqkw90jRjAznk4s2QJM7zlrNG9QYshE4l4XX0zKYqlKzN
CBv8SILO72c4vKxAXIyOy1eEmLvJeTxGpaZekUFLPIPvQmw2GQkIDJAAqFnTfaUh
M2/ZAUS3nF9OymO3nQiT63YMWW9zUqu827y2TUMl6mFU8nXcoFCbggMpcVy9RfiY
bfKtt2ddrwZMZCzQO0oWZMvx5eiTZcsBVP8d6UYwdmcVnP+y2kEkCBBCg6Yw/Jeg
6XXdp+TJ+X8DUbV0ECoi+a8sUsgg0MquSPFGvdKHZYhwnGUqIr5pF7Xti4l12nB0
OB57tYxFhvIIXd+aerd3QVXhJ7IYM+0TZoq0wvpXjGMfcqzUWtsq+KXgcIcVnNu2
jkpEtUvz5uNQAyAqzNV+p5coZKWHaxbi3pKeL8t7kOlFY4CWx/JHKfUsM8DBt7lN
kfnuUpIvWVvNztd6tslABCDSg1ru605FcdPHbS419pl5AFwZiDzpB3+UHtGZSiTy
8fgFc3AK7A043vFg5nLAI7P7bZGRsim3yEMZO6pF4YrOq1/9yf5jJ8iA6y/e1WKn
w9tI0h/6/ubFcazkjZvIW0eUheM7/W0Pmk3CLhffUZvf24llpXNLs5/AsZ8xpduT
ar5koA6KCVqlojI2J4LE5z9guAemkLtYSYaiRRK45g8Atg+fRw45Q/3ZV3NVANtG
TXbKR3BUP/snYM6JwsU8WmAPTK4JMDWpvGbEAZQQURl5NEXeqIYeJuWkwLMQwddo
ancRcpbC6jrD+tV3IDGqza3OznQezW/gwdGKtchFaZ1q+M46PAZjIcngaQR2hGkD
hgZxaDmrJlIg2yn/QBB85wQMaMbkE/joh/axTsEDl24o5dTRKUGrjlbN8we4Te/0
Bv6QjqG/dy014SSsCfBvM/qp28NR7yg+LrsejZkSGkCj0A/WjdDsZC95GDVfGtlg
s+3PUuU9E11eygBMV5JharrFwLIkCDFbs/11vhYy+HAqEEajaKIyBPA8ucMK26Dm
Bx9FCA9CEZOkpUjFO74F7PZ4192DXSiDyawDEjiHyBYzRBrFpze480ZS+mJ+itX2
U629YFgnCJ+gA/mNi17bb9jYyRyO6+0M1nozNmjLZ9NjnI5Pso+WO1E2CgJI2wj1
1VxOQIEjkPbbHaIXRiQKBwbE/PVB3Z1Wr8mPkEykrRVxVh1uMNOkYhwZ8Mxfy11f
EXsdITPqktkDnt0RMDUm6/hI6FBBiHxjaXFU3imgOZ5GuFhsmxMPjb1W+zeK92JA
xESKiblO6644aJ6fkMSy5dG68f7Ldk8S37PCQDg4A96sefA1CRQxb1pW+KCrNtJA
cdTIg0tQCy9nrat6RJ3DECcrLiKI4IPlE9wLTOmEgbZF/9AGfY5b/sQahFqnQ86/
WIOAlco3fXrxzE5RCrk4KgIveBQ1VsYRP7FMuCDzT5aRaQC6m9yc39Xm303r2cME
8c3Vcvky/xVlWJpUr3Q2bqK50U+XtvkvMqe0S31/7+lmbYZics5vf6Y8ctgS2dmn
G3H4eRWc76Qdgb+IfaDaIHxa3ns4R9sJSqXpnTDBMeS/r37n/Szggc3zpFaixXj+
oUVyQwEuFtqItcNkKXRR7wxXsw+lf1wxO+YHCgxitnHzEYbCoQQF2aXg8EPv9sCd
t3IyTi3PUUDbFWJI9MDEWSqUeKHpkeVZPbMtquYP7n0ZkHz+1tObs/oDuXAXeO5u
ryPKxZcCh/V5dTqM539T6qNYQEKk+Or6NTsbtr9BjGShCHc6hBcvH08KSrg72Bbj
eqUm+Um86Q0lFbFnJyeqqYyr1OSHAllNW+pVcF6jrjX+5/vf1xHtc0BHhbiSOuyN
Jx9BsMj9dKumdZhaIod2iB4YX8YXx+cmrK/Np/bbz+KqNrOqrU9OYcexQBvNePuV
+VbTrPQ0TQKbFYy6iX4j/7v0UhZk61nyHWhqmjJUrsQOBv6lfZf2I7FJ2oE8i4EN
4a4B/dcaF+W+XPdJN6UsLiYxaz+7e3lqO43lCDSMkie1BZdnO2XuOHh2A6izSGQn
xOrvnOkb4ZIXSIMZ7OVqpoxeR7SaMsQy0tV0YLZ/qWsjer9Nz5LilZ+iHim0swWw
uvZ7bCnZX7NujTTeMQxLpMmfnY3DVoZ6jLcf5oLn0srkLmDPHPLtqF1dhyJ8k8c0
8sYflk/PmE/dJa7qo5hwDDJhFTvepPJ4P+WA0fiRTH7NM3lpuTLwieEgfx7jVxBS
ZDz1YIdVhQWuLyRWhLtJttaZ3+HXmacniY4zBtPGupOHeeDt4csOAQHPIFZbALGw
4IFoKdFv0lIkpFk6FJHj3FDc7WOaM8H8mfeik2oJg5avLipetFsUS+mFyL9inUKT
El3iGvzzmbO/12dZsCaJHBvQhdxAbhcvUtoOcjJCh61i5w0qQhmU7PaZCcIXqoOn
RUR3Gusmn+LY5Hh3m3TwV6gz+yTOfRytufg2AUzkyZFqrx8/0P+AVcVBp6CiyTkM
DTvXZDFASrljDy1FuVNHplVuu4jf1A0D6/xhbP5+/gijZRiCyBu/usGcO8s/23eR
0uoLilnK8QRaIQcGMBd2PqSoaX034IVxN2qHk4Naem3QhxTy6mlr0zgfijfhCAzi
a1O3z5vsvkqDTNIxmFDVJueuVCpZojelCFQm5u/HFw2MZAk25I4zyi2dpqf3LCyH
QRO42PT7HbnrYRB8FqwoQ2td9wKQmrdA9q0X1xgjrp+b0shUN7MVs0nqRjtdyjL2
w6SPQ7IPjZBVjlU6SIUP7p/BpaPiwkgUC1WDWYmXZqnR0Jeh3skO/RJ7TF2++OLI
7de5q7MqJ6Q46yjqpr0iE1zxmzj0JhlF8EAVgrgqWAHubnSjSV2uTZLSzBSfVGpy
iKiqSwdZwBenzripUMVkR1GPcUCXjkWkSasKrYR6765QLWYrpQuPSmUMr/gQ+jpw
oMaSybdvHKsGRSLok8I2f3GqNb7ZtJAnDqxWn9hzq6c5jRqpc2ZKb5qBbksvLw6u
4quWH6GCQXWFvfcSiV/gFcmgl7D44Slxo1f2fEZA8bQQCkV5Ex62hyB/TXvtIN5k
2W+aI1XvluVXF1OxJCjthAg6Bl/YWFOGi6jHxMAcZfv26zw6fmhnf9VUiaQKtxsP
YZRIyKyUsmYW+qatD/CaRmDune5CFwb+CDchxRsfPu6sQrB8H5E6P05+DtHqnW63
BwNpctCbD37EUJS432unaI7niU4g9qr4foaNuNLrf7VBQKk66bwDWNXC/VaD0i8a
qUy26AGml9kBnCt+mEa3FLsenVZ8KoWQZis0X+Vn0KPU0+L2NIIlfN9gACdnBTTl
OZMr2tTbL6AKPrpoJu7TuvexNEIr2yo+eAtp0Z5VZFrvxNBR712eNYVFB2TPs33R
SLf+PcCdlpsjPP+di4aF9KgHLl28ZAcIhx7CBDw9WvenEoNnilPziBtIrqyKiK5R
WrrrWwnvMjoAEMmbzOGZwgNsLsFPTnIaSoHf96NXrmpEOEI/c2wZNGVN1ioDaVWr
5F14VAo9QLDa9K5U6jlqGihmiNVc8ZX9u8IDc5qdbWtuPlwav7AWoKgjRwc/JU0c
OQLg1UPThAZT+cI7t88/h8NPqBLZy4dw6SJYLQrlpwQXYuFxO1VfQteKAz6puGtE
HSY5D8j+Rgp47eWeo3QWx3GHF5ieVYMm8wBJqAp/wxeF0SoQgsGKzZmHxNlCsL+e
FcdkCi0DzS6efiqaxr6jwQ9XANp47fQ68GzT98alMhp+MHhvIAD5CuBW0VxTLsig
yT3QoSxzZvxCzh0R5aqKanU5lRRmdBKvdrsn9V/zeWw10XsGPhEqSV3eU3Jwoo7s
h363woDZvoRLrBo1qf3bh/M2O4jgwtozu5Oi9LcqWs5braf5T9jpdhq1cR/5tyCw
K1dFxTqbVKF/nPm8OH0eqfP3Kxo2F4krRGys0ofpHtpt2eBLk5hKpX7A9tLqSk+N
Me9lvv3MwvhYg08LTABCVXbHmZMH0tdF7Iaxm5a7pvc1BF7C1IC+NQq0LXqsHdQR
MxEZ0oGHoUeCsg8A/hmwKYKIeLfgkIPj81X3jSBEmwWk8ZBrmd+M7UBoTa+0XkOX
EX7fJLWAkgWZ6quMXtLx1Q/x+4ntV+Ck8o9huX1iZM1faCXEpuMm4pH+3h3d33Ct
+WlSmpK+Vz93JWMdtMIxaL4NSXLB2PkX/rM56HjpXM876PBXW3bfTeBSqE0WcCz6
ePCuUXmOgl6xmk9MLFy1c63VXaTDZ4AQymCJeeVX78ek8iyrxSBCj+a2TcvR2mss
+2ge2ZAA/v0hkAw9Ppkb/NvVJrKvMBNAqI0oKBoW7INyzAO8xSRo2G2bqp8DconQ
c1zm/seQy37EVNKQMdl2PLbkJ/NJyVe1+d3TkJHj0Ap/q1i2dFRqhc7QxJK6LcZt
qGh2zGcky8PgRXwPgAOwFXUpIhmZbsVvkKCZqJhEoN5j4+TMLX7ajQ+/jyWqijAp
9JhNKQXDUOkdQjbpf3N6wgVyQkZkxtQcvtW8VvYmAyY6lrt+tMps/UrXoL6Tdald
5npqly3C2m2b+NNtDq6dzh5f9JuAyYRwLvnlYoMDOdT8XvFKEHg6EuvSKZIJW2pG
GONo0kKAX5EGU7vDxAQcCYoEbM5ER8sfBtMka0hyx0Xozwpx/aiCX7Fw8WODAe4P
y2hD9fuQIxRWJnckEuc+ZrGhQsClQoG6Fy8vX6GQWSxEVF/uA0GV392n6W87zm5m
fz8hTqj5kzOcHkLAwqtmGdqyppf62AivrT3gxFH8prgptVOhhbR2ansz6eZM98em
DosP234nePoJW4WH71F4PKfLCTC85Z5qkkaz1eWBSY8CBBix2Nlvc07sq+nYSfW7
oz2jxyIxc7R3VO1/fCc/estuyABqtNYeGS4sSy8KE6ZBje5w0dJ+gb2vBuEuLK7D
vQJlm6h/6ldTj22VQxCz1w0Iz2RXJF+bPdn7I/qRH7ZHf4peHKt3x2K8DOiov/n2
pYbw3nYLS25E9VIWsjo+n6d8k7IvUtjHD9VdoeUb7mvPi+KB7viKqCDXtAs5HtMb
p8xGpVoFFR8IdQFsDTG/zgS42MILwhz+ckwhHvIeIWpNw8s6sdzwIa+jX1kTnTE9
pcKIeOsP0yjhOjUPEMOwd1lMTx4NxvJqqEMA+wG6lhYOCXc0ZLXXFmI3si4OUaxb
zTQosUJjcP5ZAnpvJYEU2UFiwrTJrMJzwpiHbIqmXG2S7AXseY0aPqxr2Q8Hgil8
tHqflHN875nUwAZTwrW8C1XRqSYmieQIJEBUQKopj2Up6fhXz5oBNVSLP+yPg7yX
W0wiYA9ZlhcEsLWmWxXg7QBm5TCZFl7p5I0neff/AXNlPIaPvc9uIc2vGQjWJsAh
dT37uLDT5UQODMOMrHtxLzfz2uofjravZNWz39SE9yjdizRLc/88sOUssfsYkmJw
Eyz1/8djl9ye9ucn78u191bflSFPvD34p8KrnCZRoZoxGi7g+ndx3FfApWgMUuSL
POAtjBpdTpRLb3k/42Ycngrv/XDtdpDCD32oGs+Sh/8Wd5qR7qviUCjWknXTE/Bj
IDqDgUp1fBxVMc9I8RMrTfG2egzcf68A0ybsExVCUFrggVmILUknQz4DQDIUp6mz
HpV50XTbhWM4xE/U6YhuvTKRm3tmUuAsUhBwemQFbXnTP7ciCNH6le2BeEHItWIV
xpDkeFzbMcn9QRlUaDOemTzAFDL6ZeDvNqLzB1EfKQ3OQ3lE0GFtJna7QOAx6ahr
Bi7WwA/DZOVZ+1w/6Ei79sDY9RSQUrfHKNKqrjZ3xCKPIA4TOAIcQikuh1lsDzCL
wRf5tntM03NJ96EeOLMU93uJtAlGqPSltCHYcivn0C2OQlNrZmupgk/xmvDN3Dlv
eAuhFvMtrYTrHmfp7N03P3pDZvYQdWoTKx+5ApcIEMBGR749oNc0hVZS7UEii81o
k3ERuDvs/fyBai5bRe+r8Gv1S/ScaPjBmOyCSrf53bEWW3Tk16xL0vi8UFrz1zOE
uKAdWYTtTytAiuhgoquRV5KNw3zqTj7sBlrgJ+uqgBCUbtxTasXuOHqdUEIPePUS
s4+uHujMB3rli/D4AaA0oxJOEbHPsRgll2qT8UOEmD/973vwv8Ci86b7EGEV2mre
kJRziA5kSMIBTJDOZPHdiWxGgOe7KzLY6Wm7RSRO+mcaodLtcwkPkACk5aKXMR8l
QsEYfrpRv5z0CPB/BmcgbVB0AE2ZvGUvMbC+jU3xt90pEy37QP8bewHDn2LK4yHF
eleyUGnQyt4hLzlWhDc1SlNUXosK9o4LZ7DqN5rkD3JZoPy7PdruJP+rd5Un8fAA
dqKn6xNIt6ND7e9y68jqVzce95DcFh1KNJ6Hvh3D8aKRo5vO4/BWHvsgdbutBpOA
KszrS3AEYoEjKuejDUhndRdXikcSE+chNQ6qjuNcbZ3ywnnkI0Q8aOjjv6sQigeq
7uxlIx4tHwI2Al4/9XVV9D+NtQ7+T1kV6WnU2cqS+e0rJH0q5qABRAEyZLfixATX
J7K2OL2zZrwhYkoTYT1YvCc5V0epBTCfhfUh0A9VV9Tgzdy0d9z5EMZfhVa0xSha
2lbvNbvZNT4IOmoJaYQMgeAxfc81bIAvtt+uLN0Xh1Qce9zWoHbLbN+DJ3W0jR8+
LBwl4ENg3gHdzd+sl1KnhbAl6CMMydSGz2XDhCY5QLiXGExhOLkLtnPsFtxCbiCg
ce2dLKXA+GbRSqKgcvzVDyBmDrfuz+Rz4/+ibX8AoGE13HS/Xi5egWSndMCFjseM
IGRWqYiTv/USGMZHB0EcrQUXg8X2qCWwueJXRS9SDs9XMhbNbmWi1TTfLPWtGA40
8ztOBwi5gDhZ7Rj0S+AD40vFtxPAWGN7PmlsaZfTQIfe3OwzG5eQ0S6zgpXdRe1B
NDUB6Qr6uW3CwD5hJ23tQxxoHBP5beikl7p9Xwrzv7ud3u8eh3+4uNMjFzOSnpGu
o4v76r34sdswYkznKiTWpICfWj7Sn0iQhX54agcAk1CCG3sDv3QoYgpxZEQGpYXm
z9bZ5tmylZQ6FVWsoW8sF4Y/kNk8kWTHbiooRfrhtYzp0KhSNRS+YK+S2MDjc7Tn
wMBq1u0Fc/AMwLWP9H/3g4YyQvjae0vyAvzqYUi4AoN1JKggjOkIM+HtR4Qp2ipx
Z2jT52zjPmoUUTgsdUlvJ3lIFNhFP3mBhJo0jkVq0YkSvVfyEzsp+cwRc1KYhJ2h
VUNSmJSOgEnskPZAmPoLPzasMefm7iYBBofIvXiwPy85dG9aLTLQQF6Bha4ivTUb
GXn28zt3cbp5usHNsoxl78jJR4fAmQwgfjypznyYK6aifp8d8MBpSUZACj1sEJl8
7yik9yV4hmvqXfHjXjXP/uFQH+Ejft9Fc2A6qJKw002QZvHR2KVjG40/Mj1of5v2
kXGfVIo68CKDpayg7EqYbg4ZzSawJNa0aEVJXI+B/t8LgjRqWrkJZCSKVTq95IZ4
C8f8hBITWPKcv3LQUe/d3LbIDls8RVwr3CckjjHCZDs12UeJITSduB/nHY8w7upF
+Pn6Ke3/P5UcH+byQX4F0WbitNMzA9PtPBzZG1GZhJ44bgDkzGG8YZ8A0NEYIZod
iKZZ7IEK0pnEOpNLJUNIXOHUDJXgFTN5IosXWmy80iNJGDzR2yiVBgKXs9wpVpXR
SFoEiEU00XRjToo/JF6OOUeajTyMGkvhNbWZsx9f6fEsf90wPUr7UDwfqsrLxVgb
ENiW2seaja3dLoAF0+watTlmhx6LEZ4n3AfkJPRDEwijmG5uEm0xix5BA8nM9PWD
ZbAwgyDBZX9givIcHFSMqwYUbdO39883SpA7gNkz696k7x+tPyF0tNvJmW3mGbIR
AoETD3TYGErzq21msAtHNRYBI1PraAFVTgRluDlpNg1Xabth17DMVYSEy23gzDNV
+ZIbPINRBsneqec15AxGzEcclNvztas6+CW+0d3I28nrdpPd8/qH9lNE3mV9Z5of
gFQq4TP4lJY/7ENLMQlK+a8C8/Ssc/gsiLoSTOII7xMvXHaYUdo5g+5DSQmrMAOj
GYYMeaSO3WnYz5+X5T9kHnIGgbeoQs2qnTAcQerXwoR9ML22MlMpZWgpEUxVqH4q
/0mSnpPE2P5p39kmk2j4sGqBaC9SlPDfFMr3fnBcOOtGDb2Ryvr1qOv95h4Kv+Xg
CEa30ZwQxLSlgnjQflUmA/HBf0/ZGt3kWz51ws6VxWrRyaKn1I8dcE8poagIJhMZ
H5xkUaWZ3jEBxfhAhGjzBrc88aYAoczSnIy4I8orJX8On5xs2qqwm9VHC2nEahUz
FFB3EfU/pKDWoJM5m480lHAaLuhBhHT75VJ6dqZd4YJdfxZ+kBVo+ls/UHCChQU4
VMzaWpyZK5P3LADokrOzHSs3fhxJ7PEHCFR+EEIFcrkfXGe82ZKQ1ntmj1N0y1Lj
EhZePZQezCd0Y8aw3D+es6OOnd7lRKn+pbPAQp2NsS33GmaKDEvja4wssXuQqep4
P0cGJVIh2HxMBO2IHTwmWY+cfuzQ48nld/udtSlTVKfsUXBVFE/VfIKpQz0ZamPv
u5Nap5xLv7AcmXOp1Ta9MicDgl9oOCPLPBoX/EFcCV/L865MuwUcd6zvoJu2M5di
4aFW2I4pejPV8CjbFAXZfMxCmjn0ueA6Xk6b4hL34q++PaaXddCDqnGEsba8BPEo
kCJvtphW9BhHZVrOzVIYf4lq863KIU7dBaznoWTBo6UFaJGCwDiIMkL0EnfSGgaV
bdy7MOoM0hpVcucq6UO1wW2LlcIuC8zKnQDdESj/lhMfReTwSYTGJtdzahI91GnA
OtVFXJMRkSmdU4PsIKissXueHo/ZSTBarrJSRTdG5cYg9VXp2fsi9ysoPyNL+DST
SxenWEM3ZimLqUVp8+4P1LLkr+6vLhjyDm+/yAm/l6XkwQWaA5OcY/bDyN7Gckg9
VP27WqpqQoDutHk1Se2IiBobpr5KHcf8ezMTbUOS9Cnyh+btYuLBspAca2r9m15x
L/t8tppywnjtGeA+Ee6J7FtEIYrc99CJmSd5NQxCfHvHo8UaqHZj0VjYmf8WO91L
fmbUEuy9+pqOOgOnTr3rn+r9iRYtogkcm6vjG1o3YSsuKzsPooY0xm7ulZb5sye0
J1g0txjc2dLRcGeOhnq8SluHEr/k5EQ8jQdSiGlDS2d0SegeEVodYXW/C3MlZfDy
f7Z/vbpENWMSzIOV5oJhYonTHiZkES9o9eHh+pNFGXnAOuSt56X/pAE0Oplv/zgl
+XpDMdEJL3jDgbe++6zrT/XKZZmSjvivzQ7ExxMqzOgw/3V2xktlFUkUw2zrzbOi
7up18tlST9XS/ZdXu5KXCrPJgbVRsc/n+Fa4a7Z19KndX+jlV5Div3ap01M+R5ci
VZwtdbz+5/8PWmgrBD65ICBZEULI9LY7kFLTAjsn7TEAQTJmVYG6lOfUjmQ6U4R7
+KY7VvjquIZBIWU0VzWH8HSILoj9h01Pd12tJpKTtgq3YKRvjmwYtlEjodt/AGAZ
Mh+xYkeYeeQNqSkbskL1SDfJF+jmW7qFR4zz5eIruRmTFF5qYD72zdeSmnm2XS+C
Irz3oh786tMsgk/C6EDcD/OdXrkEEB3XIeuO8Sq2Qpu9EZZ5PTxQYQ6MWbFyWg72
hiBzbfffyKckPqSNYuI0t2T3TohjpkePLyCliKNWRBwZS9p/7XI3XYj72c6Hs/0/
FRR+Gso9yQxzrCd0uqvF6FOV0Hrp82VzR1dOo3NILDEosYTzEDn5GkwhZDRx+KaX
COvYwr/a3uWj/Us08oTGRibooF2EJer7oq5yRXRuyQChNJO/Y4Z6jHhdJ5zoW8Sj
fSzXYcp52n/72tfAoIxTZvJQ2HckcS0jd2BY+F18IkAJBYRBKPme9KINuP/ptkiE
Thchz3fIX5rmf9zdYbc4ti5HoJgZJUqBoHbD6rPTla3lGGxq/jhJhxDfZvooXbhm
7StRTM/AU5fEvuIrgq08yzwVN65mlbJc6JJkdIhc7JUlc/J8b/Thq28VVcHQ1C9w
B9SjCOb59LAtsUwDp66uha7V1sAcpR97BgnvpfDU8hoKMlBfB8h4peh9wC7WTgqq
g/9RihufWgyVxhSBMMTF3cRrtzY5eCK1J4E0o7m5lJeGc1Yeuq55+iwklYM7UWxY
5vf42is/mwjKeHKuJV4BLih79nthyPgoPi+PUO4gQUAomGlIfdhYPi+IJTuImFg+
2gi5BvrJ267qkW+d3VkpY5qgAZv+NktHxV4TYaDkP1G92mW6Kp95i3FedjrwBKW2
1zTkiLPArHPB2q9qiTvqfMWl1taxWhuJpadyZ1bRLdwJY/75GANf8onUIK1MndYA
U7d8ENvZS0Lerp17f9CvkRpb1DKO+k40EBpZ9prT4H37i7dwO3S/qzYwyqh/OwkP
93IQgRqxB3v77slSOVbcT3ZaZvRBdtomBcNcO9DxALvGGTzmFHSU5KEyIGfMe4oW
OMLjymM3lF+1LXfO3f9tJ4xBAAm83T8MVzfFe9fkV3lesASNTQbqsPyShcjZB3BM
epnWhEmKX3WJuDWZcIkKxbjTPNCdWFI6d96l4TcIamMJQ5YPPpjJ+c7fIfV59PFr
JeY5LfJ7U0CWek7VhSqjvf0l1VsS9IRhWcaNimWakJlpTOVB9k0RhSyKy9vds3ym
/mhDm2SVVe4pP5XKU95e3XgKbSmPHBE9Nq2X3u5S1h82KBUvGLBREw84eZLt2kdi
et7Lb1yfmkNC3SsehLN/O/Cdql8lGzg/qvCq5w74GIg5DW+O6s5cHry4QOis3TYd
Nz1Mm+5EKF9tFBh8VPvZszZ6WG1bK7EVEaqxNDFdspO8Ka1Dj1dIkr6a/ba1zuQp
KJnK6mJ+Nm/yPl9LjQASU+yxKfiuSw/RjrwGJH3b6Hb2h7+Vzvz0jBjoHHAHRYGK
F477GiywtYVAbClT0Ym7+k06Wo11IUWoZTAnZq3mw7jXn6OlnRbjk/lcl5ca6lqT
gJmxy9Y/Wf7oBfq7IgtLtlxU4Ilb+A/Q0kVaOpCOrYWrFoJq/O8y+CuBZWS40bs1
gUlHvQ99NkiCdNt1piCcW5tPTcrY7bN83YhzzigNoHSye/LJ0AnDmYO/A7RjUS+j
Y5WXtbNGMw1dw+yd4sjgVw7hM6dUr7X2d91Hv+7X0P85lWZ2jiXuZqhEMBVSAMQQ
RaL5aN4XsTgfrnUcdSQxLSOr7CHy5CAg8dBPF1XUrk5D5g+hR6jRQjt/K4ITKecQ
ighzlRkz+lfQzIsklPHJAEvfeBGfzWjqoXJlwyIln4y05ccYiuxlLTZ2YAr2Oxev
/2ZtaIHCUZ3/DTszFDUMyUW/vZOUKypiUy6d9ECOjvypAUK7OniRtIOAVSts8O8w
y3DZ4nov3XzT3REQqu6VnnpGoaMFlIPTuJEKI+2VBbF3OjwGf9InQ/CJZHrUxkNI
IXVh6Ke4YXwDkDTdC4jWwx+XRjvUlKynM2ELbjymXX5yS/yvNtJrYU8ubpU1lyKa
XOD0pSzhBxzEgcLGd4Utf9pRSfU/zmwPmSaP2x4RfHUPSwE6j34uCM7nheWUP/jy
z4o0YSLZOmgqnSR6sx7Zcbx8XbTi2JIS+ScOaRwVaHvfCwADHxk9vRgenk9ffzer
QtgWYqDJCn0ZJUfnpiLwSfOhaQ9ikz8bcyy2+rCmei1wewZR1vmg407xMfnnS7VO
Xye4b2hhkmTDBAubRM54HO/4zNBl0y2s2adx2JNKPWQn7qtXysnrY9YU8ZwD+yks
3s7geBOzPEKLZ5o/f1CzKrohhI50xFoYElVmLyzfQhfsLHIu6runMCwogrveLlrX
hcB8pG6c80fw6O2kzniWg5mzSlimvf3L6totVIdrHu45SMTa0SRWWdYiXqqHKI0I
Dlk5SVE2O81Y2FiymBWbB+FoPUslARwpy01m/ecu5RCpEflUcU1Kl+DJ+Zf0MYCP
g+XcjfrR4jfimA55VnJYceYiOaaQhNXSYZY5uic0CdVivnuPKxbMexLCsUyfM3Rj
Twz228X9iHckSUQxedLdDNgwwx1jNLccV4iNndlh28kQYizc7ASm5S4gxZPJJr2r
0TplprYbLom4l0IXnBk2FrsODeLzR/OZp38zryRce9H4aSq8e3Ks7kQDwAyOZ7Ds
gfR4KZL1hhiKNx6KEO8Gel27DRvLX3ytJUsBpAyTQByFYjjdBix9OYV2oQ4axTeE
nGEbP5lmGAUfW2lQdH2e+f4J78S0pycsFz13Wpfkp9HwzItCTIJKlkkyc/rqlxDk
TwVCQZxvuagwOu221M1U2e202g9FhFh35R2PqsliBDj+yl+IjAD2vN89W70ujL0y
2+HjjP0vrxhelK0+mnxS8KRSM/C+/mPnbc6nn3vk6klt8Se4mQyvpB+dXJL7iRVm
lA4Tri/b4KODUPscHBtqydrFY65+pgdpk2MQSb++6qOuKKC/fTC3YE3AsLmDubmz
2JU8b08Mas80Tojql0oobyBthHFfW5XdSHz60CV/aPHWuAfB2oOSciXnNkPnAnbt
w5bqiX2EDWoGBeBq2Bap/E+qffKhR8/1aKZmSNoqx8E3lIpQa9JyFJkAuGKXpfgV
N6N/grjWa2RYoi3pXcuHXZhFdbBGe2Tr1EbGYOESXxnKGLCHun+Q5MF3KTuxI8F1
jenKptTtZJwq2Rl5n3DB5i293y5EK6QALYFkaqjHA3k9eBnhBK7bY0cCVcIJqO5C
g5FZzcHEpq1lEO20qZ6DPSr+mPpcoNgtxpz+WF9eLsr6E0u/CqV+DwuMrgBJJwc/
R3wi4oS4ZYpOZokLsLTJi9psJkbCBeTZcfeOlMmZ1DXYq/s1hze8DnaeEe2B3OOT
n5rXzPbS1AOgm9NXuqqSqqLRgxOJ66nragIWU4Z8qGtKzmolokQyhvB9hnf93vHd
cmIE4VMK8CigDhFbL+qQxwlv1cQepaUboMAYq/QDqlPNbIyQ/Aycvsb69JUsZabM
NvHys+nuePyajSZ9GbU3MH5DEB/ex3RCp3Rh0MxFYs31OX+Pk4PZiKT/P70tTp53
3om6wEgV/YaJA3vZBFn0Nl3oDQ0HQQxiSdias8gVeUEEJWtXTBrMS/VIcPhlBDeh
ZNTZbCyH4sC2jflMJIc2gc/SzEfZ/riKBhcHwEUIlaCsBK06xi1kw1GrnxkGXlfX
zOwRfx/NTnOP0WOOEAxFpdH9saKG9aJm9LLsYQfRJDi9LIuoxZLGq2zVHac4xJov
c7EfvHknYbyuf1yea+L1W5YlCgVNHxalRvOdFsv5u0470Q78eRaz4WeLTo5crYjd
ZS+9l4GxfXeER5LHly+wgpvROqftqvEjpim6HlP5pz0KWADCYox7IKfC1ncS99+o
m7XiiMOKy/bNE+xNw6sqAVTMxMiiN4aHeBTI9A+0d4MRvIU4qB0pi+KjkK3LZLYJ
6rVTCl2uft507tuO7KcCtuPi/QOFbhZGsQGTOjBwtO6Uu4FQiXZ6cP1c00TV/W4o
Qowkj7Jog6uWoxhPeLcwDhv8BAueBDnwWnk4g7u7sLF4Eq/vy6jpesDw6EqpOIyL
rgg+6KRFbVAqzK6qNaD7x/9IIk7B0RkTGhiniLw3hkRZoPAg+e/3XSQTU6RL+7L3
WZ8LSEP7Kq5fK9qRxOjU9AMl3dAkQql/lYnJ/Slx5Gx2VV13+h7wfIt1dA0GRG4q
oABLbaCzxI9D2O23k7EWjj8FsaGXh8mtLm7HnAJLIVI6RjiGz9T3jIv4cJExUTW5
s1avhiv9u67JEUQKDlOs8Nh7siVOqM6bz02T6rrFkGLHGRokiPb5ULKMizU9FNVf
k2DblLbkM7f0M9UO7IT96O5qllMrUTYAOTHUCNGBH2AF0qwyQnWqxi39vlflp+KV
icEVuvXYdu6GrijX+IEQY1i9n+7aTA9f0fI4c2egfuu44p7qpNhUM2r75TSsbBjc
LOEZlGJu7syE7JSp3xWs9eFPoW+Cx1RfY4WIdgsFU5VDHrQsBCYBhKQY/QjyxI3c
k4Ji4SerW4b9NJDLPWvGxh9Mqwng9kKergYNKvQlxkRxHL5Jksvn6AknllqWAxrl
AYNdrxSLHM84Qk2hqfCRXkYuvNpHiSdKQ39f7Uc7087tFyAfQ9nYTCmZqSqLVbnU
HrRNCeXHemT9kodlVAJpOfiPvnmApaTw803Urt+oGdV+ThIj5Q6erWty9NvKjROS
gdn/qAWYgO22WY6LlxRkZ9wQpuZZsCunMVS+jHAb8qPZ7gGPDoE/CWA3XMHYiSIX
4SIdUXssWmE05OQ82SvxgH46iAqcOvUgqF8Wo8V9OIPFv1aZOgOu+0YYiiTLq+Mq
uvyHV2p3vFaYtTho2pmc0XND+KfH2Rc35q8gy54RBL4iEqF25+9YvskLL7n7Z6kO
h85LyCMswd3W8M73TSzJwxOYqnZwk0FFqFl86DhioGe1RTleuHM8aV8pCaoMuZ4W
OjM95IBC6IbTs30f1Y835//RfTa3M1t+DZBZlhllMGsBpsRAyMl4lMecP1VsIeIP
icyE3qkclAI3K7PgeJoRk6gxoePttmJFBx5ZVnBWRm/AqN2zj3nENDSoWFFT2F7P
RZ2l/w0P4F3DMpAaTEZRK6hurfU1FTSo9+/uJuOH9n1PU+wvS8Wr3wEfXWZRtwM8
h+VvA1vry2I2OsYvoUztsvr09UTAsyXFjRxYvzv9LbF+KLPQC/baarv+EKhFvx6z
pxVNduFvOkt+mwZ7ioHKBoxaBUm/acDdyTxhUrqnvBZnV3Sst1IbDXiZ9Ag17I1D
JmFGN17yY2QwSWSENcIoK1HUFTWv46SMuDZlBkWtv6rrKpMoAamAS9ed8FeBZ7x2
Do/5iFJBcxauVhj82qYEnnD6RedvbnXV5a2BI4vwGyoVRUN3OL9P8am5C2b1Z9de
5CC1sdjuwe4tgko9PgTUJyhLUYgy/l+ir1kZ1BiRnnojY/ZMxB6o4uQHy7JE5slv
C8kUU/FrNfwaXtLGQzPllvY2ikdpIRpB+d401tnbL51cRj40G3Pl3gWxSQ6TPc1J
U0d0nUyje6LMBTmsDVdmYl9d93AApFKGVWjZq1icm8ffI6DHRSrLgedqxwjYR2C4
IgBr5cNLwdejN2KhY085ISGqFPgd+HCi7xyuyFfZoCDZ+GWDaiY6XuJl05lhYqj0
VVkG+zw/UxNnh06QlxYWGKxqaDH74DjjmG7EQUPHMu5t4cIODkGMwq4FRqdJ4z+f
njVYOIMQciXp30J0t7s2h665vz1V/wQ63AU0ok61PUfpipQ71cpii8GN2uc02vs3
bI9lsd1l3Gcvf6iZmbzYA0h/JmvKQhO+3LIXqLFrpap9BFcnwHYP4LP74scKhm9B
4pbxN0AycB4/fSXkh4UuVgnFNvPRMrzWlrZG6qc6cm/s797ie1lRtjQlhl1zmI3R
73G+5Nxdps2ZCBjSHlsQ3FduH+68y9m/Hfb+tOKcPZ5bQuzTulanqwGve59ZT/lO
MB0MP5pJOQ1dGz7FUJY0xO/4xpDIs8tZ374c0AwJMKEbnTNsOPGtAwQUzEjNw7zv
mpz/fA3hyabqq4NCeWXdjq+DNKAmnVIRHSY3Oa2HjI3z534TcE9jl7nD6AfK3A/e
uODwUjW0zpU2L9ZS3zhC4+7LyNJ5mN2gw++wUsG2dDiT9Y9nqN9UQqUit1NQnV7i
bCSgJVRgsihFGFxSb7sJXGgbvzHwx7dPoiyRVdW7lRPuVhMj4NPb+a94lo9V40ds
x6Q2XdUB3yGU99wcfFEH+pWFhcEmSnLt7l7WkFQSh7gm3iHn5ndxW8BdO0mz49+K
kIJvWphTK0ltBO0T9DMgwBuBuExudDdmqDwS2x9IwG91MwjhYduYFtyTITz0cElj
kkSRIOndoWEMsg4GuV18K/vlVXds9zZEOIh27d37DdLCWa3omGxwjbWX30OfQ8Ax
a7eYofwPfdiBZ416gn4cYI7R37c9GD+JU7taPX2rmrK80igobKyFf9vSXSveNb2K
TfLQgTTWaUVqmVa7qJdap0O5320tAMxNcGu0A0tsgHp8U1cvTzZ01gUHj8DaDgol
xPBASwoCWPsFc7wuSKwGSiQlE9Nd2rVsxx7kYYQCfKPED7sN8U4ilc8OmG6pUWZH
gHRCzA0wZhvFzhAPfUZW7prh8GM9LBYYynmuXMIxHD6zaqICL19ZvysJXI4RlfIG
QCKPdIVOMiOzunSTjre5panCmy34ZT/osIwM2F9O33xP3cgiRKXdajB5kN4od456
S10MlE7g3C3LP4ADmIsfwhpJRXgWEMGfNdZIMni0CcgJBtWolxyM/2doC353XCtA
c6MdMMjLRPR69C2LPmacrKgkQe3pw4Ug5LFnDZveHORBOiopkrG1m8gjj9Q4W+fg
ZJxCEnLSDnIZsVbjpNod7FCSPFDbCmilRuJvUDO4gP0nUpif66KYM+Aa30Fhe7RI
2Y/ub+lUXr0s/LgHr/JBXv5eAiq4tjCs08pS07f2QTt+iaNOGFextRg3n7uohPMZ
23XW/4J78Qgj1i5lFwJ8hJiCVi3QU8nMq+YhRAfzTOOvIT1II1gWJh5wfFbxlnWB
thsbniBsIY9o/fFGkr5Jq7/6uDkRuOzc78aM30xGF1KB5GSxdgzydulZbBOEhsKm
n6//I9ozb1zn5lp63GntZdOOx5bHnE0Zw9NE0UneRN0JM/KTfZ3bwFDUZUV04Kc8
lfGIOAhD1hRMPDQHjrrvAgM5dXwn0bXyMiTw6MEquQa/nBp+2Wop1wImVd9NtzaP
B6xpU57uiuBn0nuanuo6Zszmo731P/82Pl8H0XqXNsz36RuGKvAjup9PocChybfJ
eOdHC9IqW11fJu7PrTxi3h7GZzaAUUKbZX0z71ytsRelXuK0j9Burhq+aAIMfzou
aqgWSBHwSO+v4GVbPoY2fcJ+4nGEONNpoM7dpScxMtFwbg5UdrsAvzKepKK32EYS
7cbl3jHuu+JMdoC4/hwS/yC2A8vh2tdNNnx4DL8iYBox9U9F1h/dtb3qof3ug0Xm
XD77UfoWPF+8teaeXXH4gSQPMiGKNpe8IfIzz4VWvVl9BO0ZjwB8fiwRgZiM3mur
BSuUAyvaAVmuSHsAWUnqngrK9rYutbTXfLLh8ID5byuGIgACcaceZ9fqDVLcxZlZ
8hzGD4zPmjr6UP5WxBqZl9nf2WEe+2FeW0pMFnxCciZv4juVgYYntwv2qGRMDANu
h/wYkru1m2bQsF4ZoANs3/LTruNqQv07opmiPe7ADk2Nl1o+Tw8h0MtMpvlSfCFQ
DffOdDOihbmVuGSzLB1Qln/QzQTdqjuYEQfiKrin1Wk1BJ9Bm49wJmVy22Nufdm8
fMtnzLVGhs4x/jPmguO/0Zfp1ljzHSlV4Z+azUUJqxXIDSVSGgLHDBkaGzgKamqX
4M4ewyjGlbi0cTLlXoN8qEljAFds87dLXx4lhZcQpxr/OkwBs8nMij4Ryh6mol7G
jgm1Q6Jsc4SB98hOABwqtzjM2u08mClaC203O+cb1n1AKiiWmsCfBLvySL0VVILl
YQtmAS9nPVngT1BM/tKMQw7MWUKakhugHJ1Bf0Vw65sYcQRXS7kLPGp3eYcOE1DS
jIuoul9uPzugQcexRDGJY93zVkQcIWmUbAB4+l1SwipxQ/rolqg/NFRCRSa/z+X3
kZl/FffKq5pfbbWtMSS4AVNDwUyfZUYNQgdISDU+JcNz1PjxcMw488HluzhCTEe1
fj598XrqI4EXd64yRPi57mWJdFvoAEYk1M2dsKnk5qvon+aNuHHglDggnmnkXBS2
Pm/QjOHIOe+dJywE/T/Dw0J1U/nReKbWWOPfVuHGeaVyDfH+bLxNbdxnGAmKF9NN
2w/t79p9WVGmcIKVSDxOzcVAsgu6ytI4xHfnO/1jCpk2eX+GOMtFtOaAVzy1dWNS
IYw05T6wxpMbZw3GVj2uoqKn+8OHrOF1hEgY5FqTbKylkkqvHfWDrv0VrgjbdYDl
PHuxV6fMX4+i0pv5e11I0oSrTHLar4OeNxLR5j1vk6wnZcDS97fAPmwOnEHnE9u5
C95HhMp5DIzxSHzjqjCRvdbclOmS8znU7Ca5OaMHKbKoaoOJAEpCdMqLbRK1AShZ
7U13x1HgJlwNlyLNwkHBMq2Lc7iWwKfwk3iYpZvI0o/fatoT7atXgKm16FcK5pTF
btqaRxzIRE2Tl3Ymouvt37vVB2fEB2nyPGBhm/1Ieqb/M6Qw05Hworupf9jtfpq9
wd/GZlCG1ExwatQBiEk9phZlbFBS+yG9hw+FUAGOayjMXIiBhsskRUz1jkcj4lFc
Ln+oxNr7wbbP/bdlHFbpr1hdzdrb/varwCWzGjIzbdVA3CXZ5Dnc/QYOSygH3EDF
xQHv9CX5Mgwrux+zmAAoV3yFixj6bSJUs14ctDWzRvyU2fPteEZ5FEmL4EJmHXkw
U43M/gmo0vA/fr92fGOlMpZGeGrmGyOYkjj3PAhrIQRvu/SBSrXkIFFN9hHANGj5
AmoSpQc4iCzpffsMXRVnoY8vMBqP3aef4vKXyssctlyG3ReQKZAL1oNn0ltK5YG3
qy2FRSZuNPAyJ9F9oE1PF2VJHBLjrPI+rGMIPOhUQv/yE4+tckw2JBYxVBUbsFxI
+106htHedMHjXYH1muwE3/DXTquS4IzQUv8RKPn5PBXjFEE51mljRGiRqZVFppiS
1uOwaxfjR2ALTckWp6u7sD6ksw39AeSLgNOSTkaig7GgL71tn+PtrBjRkkM3JCiC
7MRf8H74oX9xoWhlzQTa/FWMbQWWkSNInYUET/YO5HhhTEnY8XmkC4n4NjFt8lew
P1dkI/gFQc/BQLHxBxtaPY70sHRLSf/NBGPRD5W32a27j0f6TElzFEGEoZCCU+S2
W1e20RXsoC5NKwAs2DYcfAxRZz7nk5H4kd0itvWyS/hiO38WAxWL5xxX9ir3UvhB
yiIDfdVWQnI8T6thZXbJwvlFG4SciV4D9XL+6JajdgHPd1utKEsVo6l4upFS0EUU
DHNrLVuWUN1yVUyRuCOhvf3bSApS0zr+6mDNU/XwX9DT0izWPBVy3rp0zGxl6lLg
nhocgEwXT3XBJVjDbGPIl3xJqeCNuNXiKkvgzwFYbe5OpH83YJeJUjOIhpZNL+4R
EwLrLPeVZIw5vIEIS3biGOq4NORbvttokkS69jlxS8koQp9AcTtvxK4Ixc7qwNlR
jBWE/MU2Q+k/A3gxDcSn9W6zfWQ/s4YSTbxgwcEzomdpN+nL80ogCQFCUBIB7nwH
nInBw/yOBH6vESoCov4VNAgWoc8voLjABI33POeMzMCKvQQeQ0I33yoNOECoehKW
t92hakLSwyOGtxrQqIn8ArAsXPBaG6Q7g6E5BHcN6esIBWKoEtkLY56Xq0Q94gz9
9NJUAUgZl/CBroCZXSvZEgG6w1gTGR7BEeilrApp4gBk6J6Z0LMuIppbRBFlzgoS
M2lQdk8qh7AaGgJkCZ+dtixCJvrAJ0pNhzle+bLxZ1o0Afp7k6fOByHwWeHPIvsL
wd0TyFOXyMAs1fnZFZ8Bm4A2+hsa86vdH9WWJ9ea27Jzg6tIM66xlPXORBg1+8R7
KgSzVUCjnMjHJATqevKrn/ZEmnisRm2b9J/5/cE1IrBIJyomYi9Qiq/g7J5tr2Qs
Oa92WUBsTOWE3vdovh2rsffetP63vfx4WImX03PAdNMoryDj3uiInfjjoJxJhMv7
XSLDdeIRr/zusELkEeKhhAL+pPVWG2GoEMUFNYaD04tNAZIXukA5w+MwpKIR61SK
LG8MElsODC7FmEnrQ5ec2LQ1TjjYdCIQGvZqK2hrg23mW6cMXqxJjZ1Z1fICKS1N
xoqdr8hllMTZFeNxw8iUdmffOHu6BNCOFaZ53WjSJ9OQtpG3XtXJ5JwDj5E7MJEJ
I4J3x6Hs/TXJxtC3fTrc9144KeClVghTfw6T2WjN3v4v37NPKJF8mtJqslyLM2hL
4DILrDq5r5OKObZ6Yjkn5kUupohmkFY45vwE6pHthmUrSIKaLuxJctgnQ2LEJRva
JJKd8aDaNkMxiKSA3oua48V3MnaWSiCqWioZD02FltuV4hbg68ZhXX75hFkbABQB
yr8L3bonnNbQfS6LRtyDCkeVg03sBmn8Bq5or1qaJLs2rJSyEjYzNM2UwWzOUnIZ
RjHzsCWxFQIHHTtCKQEaImFAEy4ksCOpr8SIKiTiuR7dV07kv8IX+xZJ0GvEgcjm
++de9zYIaX0SNQZeRSXE8xBhILdX4rFRzQztjUkq96Jagn1wE5140FVOf1F2Q2zB
DPHQF/B1m1AbLpdzeEVlTtsPwu5nQ3mWwks/ZkpXiqMv56fn4RBLbuwkQYn/1uzz
2VHvQP8ymyDmi/LolUuxiWTnpk6WnSMQfOIdhpTsogZL9tpHez3hajT0YqoXI+Mk
PI2wBPk39pMADc67VjHG5L5VLju6k6n+b7pUhatv2obDYaTsly5w9TsUWOM5EhB8
SATjjetcbYDapFi8r9Apz6EvMNdg4bicNh9co2Ls2cKshJrBrDXbmIP7gmGbX4eW
PCSf4NevQ/sh3skdQTe/glDOFbc5DAIPMawl8ByfYxKEbRZylBHxQ/9M+SmARJeF
4shOVLYk1FHq3RR1im4OjQg4NzAux72YSGvDE1JQzg6LvcPyqBHdz0pZyR0frQ9O
ZmCH+WeAcWbOQ9w+i3mhDjZFQPVzqjWBOaFntkS+zjFvMFdEN0f0fZnhh+dXo0oM
zRbHtj8i3N6i2xkdizFmDclRgkcNxC/s1gL8i7vkvADYzqAqbrxT1Brx+kCgRHjH
YYjWx3Y6KUgd4iWp92hE5ujJXniDC5pA2PyZHlW7KxoMrcu8Ri50Q+8PtCBMNrTf
MRPRbFY6ZoQ8Kr/MPfVc28bibaeBUyb4kDYFYksWdojBYky6UCL4IeBmmwZBw6Wa
rWbHzYDNZif4QgLaOoxAbVezW3GPgCYlIAcojoEoPWeLXUuXrlwR0KXmm417m1bV
e5NHeuMUmWCwFUM+zRUQkqdkyDlMJ6o5vW8n7QsOW0hPksSFnAq4E9+ZmFRR/Ogy
+e5ZkSmKwdhcwYI7DXUMMCGn2nJYXEM6EZEeXmAOKeQmlM56XHAIh7xKrDbTriOF
vABSfnHLNrZUOWrzI9YNsQZUdgk1+uuAG7IyzjMNJ6ZPZcHYRbC9RmdJuqzq3Uj/
ab2yUpMtAEpzZf7jCoUuQMmTwUB7bZxEAQ1cPpBcG3dZM1tx0mhZ9vdTZJRCFVvc
Qi43gWOkdfHnEOOWk5XPfMKzg0STZrLmSvGMV+urVT7D3d93spfp6ykIKZcT4W6Q
+TSs5DcsjQmkmT20L9/UfwfHIZYXqYLtsC8+3VbB1W9hTnXfeY4lJY9FZdFNEaK5
TSXitCfNVTT3QvpE70aHmbEVewlTBsZ5m/L6woFb1sqyr7X+1pvFOuZsJlbAvECB
yh1PpyXa3bTBQwZ3n42FlV9fU8c/aWfYSeXoLbGuRH/APg8TshPaeRaXMFuXKVeA
5rkXqLnAAqdczY+gva3PtztKYMlycEu/NceBYgFYB9zJo0VNu7GJe/Z5T6MPdkFb
zIkX7haahezem3tnRkvXdLW+rjWNazxQUZNBtK9wd2SHXbib2SO3l8kRpYA9jkh1
QxFObSyYUYXqVm6kYNptBVmES+6xgNPbEi2tXuor2jODzUG2hAoLiUI0zsQwmYQz
krUMH/vntzhucXGzL5vhj9KVDIPzvYmUpt7F1R3iDSwFd2fpYZJojgB0Lioxeu3F
whAawfRICpbgmEQX4fXR2iBOF+E8UEk9MxtMgx/w2N1klmLSQynKeVAghpD1F3lm
phNGCqPb2j8HWhf+D6dwovHUUO7Wfxh38pVasAWh8SJdCBMkx/IOdIV3oGJfbNSA
aqzjO8wsWBue65352TagDHEnDbFw6V2OXUx7NHurh/JGMPNiTiBUYInMSTq6pmlr
CgUpWDBqauClq2VBbwFn4vcm1y10/HTmLllWiW2XkxnDgzVvEqs7WH/8+PKuU3F0
JTxLCev2tVVNc7HiISlqH1JYEhUoeHqQwoP3OQzXrMWLYaM5W9mOzuDE1HpDtZOH
FZtt2V+bc+xnV1jDBAzuOsq35IrtajiGjcuuq266UKH0EH7meXu73mQlxwCTc6qM
cgkD4Ub3N/SpQNZVnbdtXH/yetolvDl05ig3Me0fv4vADBYqkr8bdQe+dzq0+abR
Bjg0TY3wiJjoT/rGFEga9XAsxHhSG+InVNugEAK+dOWuwOXqsr/m5bb7aj3TJSnG
cOJ2OGrHCuMf6IIHNPBqKSE5hl/OqFii4R6WeepVo6wrCGmWlJs65viqkHGj2h1k
Fh/pl803OsiQRhzH61D9/aywlYyvTPsGwaxuAcF15iDm1uWUa5Z3Qlj3LW+uA2xU
NvceC9ZJIIypcz7tk3GZ/6z9rUbMnndIDVjbGaz0Gr6/HpF6/HtBbloiy2qp7jj6
9FD5L/MswabOYWNzK8s6qOCvs76AQzfytkp0aAVlTEUhw7LIYAcslLguHk1S7j+y
g/pR6OUYyBVxxnk4Rh7v3Wj8VFn72u8Dd3I4f44wMQrKE0fRdRwW+dbPnZ9N8cuj
Z5GeOHo+06EYqPrFAEAy7AoljpbwDhRYL6IfNIpexC9HiuishU4Q8U3ksEySMO9P
smvxU2inQFeQ1JE+aGZEcSvROXPwjKrgW1qjTNYDp9KM/DZB2q45uziYvvTWvYvG
01VTJO+x4/jO2jg2Mekcm39iwMPI185whYnyiou9v4rIe7Ronsb9AMZWvLCtl73p
EQjsFIrC6fB9L2i5ISrasmmyslBsWaDBvHpt4ioKNXgOSa+glxK0nrxb7rD+wKy2
IwwfG+kA4GlJ44UzPtsuOYvrk82wyMJDZZK906YN495KtEBBK4EGBwtj3rarDvvt
BRWfvsL5K9vviPoLjkll6HyiVa7qLkjMwF8lSZ2bUu51khDOsSFvhkZ6EPO6wj+J
Tgn1dFLt3SpUMDBJwrBDxV+73us7tYHQbAEC4loLBMvxHVSAaQAr+g2wxN1G2PSK
OhRX0D8fAX3r2/CyV6m5K5ztyBg0vr4RM99kYtiHEglBZ/VhECovPJ5fZ4s241gB
yeM2Fv8XdDgGsUeXDJiTVo+Y+QQ2SyUuffhB150bjdlWrC4ttme1AeyHRgFkB+5z
fv0DEhwItTNu0xBYIendYB+Hu0wRcHojPOSXC/ecwFeHAJvR0RB/jZBepLSGaskh
AXn6+7/xm2rTW8I3mMhEN8bM78nJ4motpP5B2asKPCXRzANHPNsEwWTNNjuOa4wW
lyUBATjsCV3xKOa6diYH1OXTvnusMY4HejwyO1cgA2CEdi58YHG3vP5dHtvggvqn
+EBkQJbtYFEScpUFwt+RUjAinGfBa8C91yBQkRtFRUP3Yw3cCYLICJ+y9gNSwWT2
/sBLRWLuhKuqqEBYwYh25T0lLJ1pkeVKIyfM0uXpJanevMu1CwLaI47DsYIR5VED
YpyylVY7/IndtOM9ps4Ez7r720/8b0VeWNgBiXLGgtQRBd4qBNYacOOv9Gt6EVxC
0GcAaIENcUwArnIFG/gYwKsEviTPZ6z9yAubahhaze8Fvxr3GCGceMVWZyuW+kBv
cdYO6Afw3B1RH7v28R4xma4jEbWhNyXxwKqj0oqCYTUM5vMX0aDYphS4yhiYmTMk
wr9qVCeqbaAFMoImqGawFBfjWdZqwPcAeM0fRwAO+jjONx13VoBNXqOFu7dBOlNZ
ztChk08aJZ7trUOIIx8bC32UYcRyTeD9t56GibeciKoY+L4mo0fwqUNALYEBzx0f
jvb+m1NhZaZ/dHnmG8mUcIAayNSsgwcZgZ/1PE99sfdCIJnx4XdNInf+mUG/AmRt
yQWqOU91UkeSurDcRKjR7rPydz2lef6myleGoaLTYVlI394HvVsi6wfb7Wkl9h5S
X1s+LaopOGOIwFIFaxN8pOZq1y5YLAtAE8+dB9ikFVUInOyE8maZ9TjfJe9K+1kL
bGuT7XdPvTHCZ32IKug+guPpi29CpGO2734Hjk/EWynuX1B7+Qb+xlqGErfvwFvD
W9Cf+D2rt2XEQq76RRd35LEHEyUQpsCpXM8NlTYj6kUTqEMuv+Czx90rgITx/QuX
q4DMLSj3BnpQricQvz1AMA70hv3JR5LKxBEPBJgYFdQ73QaDjA6F913n8JxKWHQG
w6r5HUnA2rHckEHW1IV4Y6CVgfum50hbC6Lq6QFCRFrL9h9HTvqNlXmkwYjKa0Ll
7yxEfTLhKezvouu8zIyL5oSVZ7Wtth13JX21jYk/D0uVJEnVqpuwhsTD+WLv8e/4
MoIxuxKwqVCEQGg6jzLXrGSzrP+AOStlWs8t1B55p6mfYFOuKM8l4d3JCNzjaXS5
asaeu2zxqqX//hi6x4yFTPUtUUYyqcFkAiWj8z0r6CADwI5KK+OcXz0/4aR8CLA2
yOSERjCcGE3Xr1h9Nx97e16Ev6KDQEo/9ktIXT6KFqeKJiGo9B+z8vB/n6wdcOuN
Ee/Lo58dU6IFgWz5EguFRer7e31VRxaHIZaMHkV6qchQSuxQJTQby2MDALwe4wWk
K6DNY0t7m0/1hTPvaFV7OqoVpdd0yeC1DjWXt3HNzpK8b5cJBc5zm/GdN3hJIlUj
GeDkIPRM7rc1bLcJgCuj5B7keQjojd3AeBx9SWA0IKP2tD17Hxv8hFweoT8tXZP9
4lbSZVXoZ1L4bEihTA45+YdWCPGbq3Jc/WjGC83C+rAB3JhntppN15ScwJeE8dFW
wWyZAWLm2TmUS6ThwYEkr0L5yRBDk5UjaeKxHtf0b7/lsmF6VyzoOJfOKPGElehD
r+/Tc4FmKxDrsICugs5c5iqsLQqWKXAOltIwrEfPK8UI0JrXpQvrsktabpzbcjbS
LIJ1cSTd449EAkuq+r3L0mGvF6dfxwDGBkxbYSFT1+JjJDpzkHX6S/RDDSLkCOpP
dUahU0a0CiclL76ckxYq++GgDUmdlL9AR/lQ3BklFessGQfxhA+npxZX81cEzVyR
MuuK75lW9c3JxN9q/AsZgBjZJDiYVH7oP59IOLr4wWRm3XdTFLFKIPF08O2VPb2J
j/gcCAWP5L8fKKD/dzd03biYPmf5fL8uDPS4oIketMK965PVT1JtAxT9NjBG10Sc
FtYu56UjlU1AX+Im1kgePUeeK6HcSLkKf5fWr9A66sF0V9+tyGP9R4dbIHI0HZB2
ZYm3snjnIOSGQDq/q3+9mjhrCxmj8YtnDAqFluoYOD6M3rkw0VGzOHGVyH68TPHB
3MyTgFWiXMJlQXByYxM/qWJq/26h8xIZePjyrcdsB/vwyPpavvhWaqoHjPzqo1jW
HcIz3VyekPYaud99wLTCmv3ZkFoVSkhRR2Q4oJ/3dvxHmNXYCleaDxAQsVNZp7to
2Cao+jct+tCaofbpKs9FUM8rYrX4SceAXcIRJSvnSsm9oMB0ZS46bANSfNd+9BFN
4bQAAzBXMoZa7A5QChPjbMd9MorWCx3y5OdzU3ZWLFcsOkXnWzpXIzkmzcdB0VJH
FwnnOrzwJpAGCzyFxBbKsUEuIKMm6CkQP1ncXnZ636LNdzJsjAEGFrKGSRbw/Q6b
QKSqe6B7T0OS85DvjSJPlVc9/tpiucIg1j664yP/TIsIRNnPyv/BKdxyl+5VKByE
AcOSZVaOOxLYqiYQz7lLa31g1XZrm9kZ64NVfxMETzckGpIDvI8P0sWYWRWbiSL0
Hl2xONb2jobiGx2gNUGO3toka0+ihmFdXcHdwpb71Z9yjjUyxDhHYH/8wK2iWA7p
3CKXzQSAF9MJ5Fwth4+Mi3RHkfEBKDz6xGHEIm6uOUH2oiuTVpqlmi8xNA8yVsW9
wHS3Hj/6Xrc0onXAfmFzTlf3ZmZxOVKQD5nmVP4kERlm7lmnvNLSuF9LFxb78StC
YoizJQK7W4qK5ETTvoOr3uEssMKJuCrlfzW/nW/h2/pMET8jk1kBKbmd1nqgbEM7
3EIl8PgH3WjaFFcPe/hBmbzrO17b9qBDn8RID2jusonqaDfkLEdQrHUzeSQvyCYO
2ssd9TpcGgGduSUZE4GpvdQFn2dBinQyfIURydBw9kc/MUj7KomvcLV6/5Il5u7K
t3f4rGP4az6eZB0AW7oXvzh+c1xMjeUFURGTeGPSlRy03zf9gC2hi84qryxppylG
B9fPeniHLMWJsW4I0yEtkDxaRRAf73MAvBDgwDjY42X/WgIP269iMICUNmdWHHr/
49AIwmII6WH20dq26xc/RqZJfScXhEA+M8L2u2x/TUwuuZSWUA3J0x8PGjWCBDZU
UzP3Is1WWAnu0VV8IkKdqPcPe9pMi3Cae9VctEN4OnkY7+QA2qrpvZCUF1C7xw24
JxbDEC5gy2U5sBpYfskgKBFmFIcSGy4vmrBN3WtnVqo++8zBWxJxpumDywDDAfZJ
ix1oMQ99dQk89CbhPSLU2J7O/HoLuuOAeqi8A1oS1kWnoQ7NqyR+2wxEwJ7Bvq+t
NtNYOLN8NRa0IRDDQMKpLlTjeUVsX9QxzEjSBxtyrCOIBadu4NnAecFN2yK1GP8i
c0+Ht/3LsealrAg2GDgs6GWOp/z1PLUPqVi5C+QkM/6P2m1YpuO3Uc2uQU+D3ahk
GFPUsl90qHIt5ddGCrwyIjSkCVGIkHWCKvOuhW0xZT7Sn3NlimAx+ddq5vS2RgLK
zC/xMgjeLhINA9QJyg7IBHB3Jbdo+lGp39spvbiWemoFURZTqsGpjo0vdbwwNRgj
jKdmWsaLJJH5ex6lfeCO1V7nQji24hsk2YhtqKHXT3Hac5Mp/QR5AnFN/DunTqhE
vCAbZK3/66CUq8+kjB743Rg484zGZqzfZ/P3v7tcAVExp6NvIJiX+dvsjMVPBv/J
IqCdyjo8FTiZslAAk7hIqWed5p5ggUMsERBTzy2D47fGaSFFxaRy5I6nhOhr7dvx
x7kADWVjV+5qN2/JiYTRokdwHNkvHW6YAlqHjJ7S2gOEniBNAfhOEFw/tAbsWwU+
6aaDdTI0sP0SlaJWT2krZHe2Hn7I3K3f0/dJY6yLzXZZQEdT5XoJoeCldxcPFtX3
2Fw2odddbViWmICA//yrORWURMDL8l/OkLNjSciyKd1eMm5NoBPOuVRZ0Dw6kEoO
3+HjnN323vojavlSBTKUpOV+WyXvsxYA3cEc9d0Cqk6DeDykaEgZJmQo9QosjCmY
vAprMUCYhgRXQ4WrkR0dGP9vmbRgqXAv/EmpL1kgXu4E94sYesVggIbAM0BHv3MR
bjTJWO5iWE2UN/5j427W5R9isZlwhl7Dx8uPv6nBfihmFBhkZ02fg31JE88yySM3
2+llL7DxigtSRAuX9qOQRUpiZEaPfo8EKrlhbCQ0yp7lFqp9cNrnTYCgw8IeVjEO
2gOC0AU9I57seUmA/R9FyW/KaLFOGeaIsj4D1P8VpuYvDssv5SwOBxmi9gxBH2fs
VMlZCh87PWDbO4htTJiU/OzSfeJVOpaXzGiXyrAfTRqyIhQxoRlsRTO0cCUgGPzF
8H0aF5rQs3k07F0SIA9eq0v+oj9vHeFmQTxQDIs1rgJcvINhFwLGtlx5N6B+07KS
oOwaZdTZByut1ag4GqHdqHZP9ce6DnDVUusPWhvLfhyCN5tYS2kxYJvm1jaeu1+M
rIm1zBt5wtMUCIS668w4x+KKI9Hy43Z25RG5o0ett2aJzUY7QPZn/2PxrCAzieXL
54u66rcSbretYywCZfNHc+YOKqDzJQcrhaE4GyG2YIuZEaaS1OFj2gBCwmEWKtLD
0tA8mnIjfDoPpAc7koCuMyn8cHAfRzhkMTp7yCRRktCg874/57qd70xtZnohCkJP
spTjLm7NidQPFBsHXh2LTN8Qms86VfrO6bibmAgVBUx2bkwW0c3UVdpSFIcuTtsC
YIa1ypoesk0slwy1zBBhQBRttXpPzuWDXWratJg2oaMfGrfRKbE16NgZ4RWtmWSU
DdRxz1CYlr31lrbGFkqOfenownF8sfFk5QAY44+EK8Ui18oXb/IunIT5RbkHm+4n
4xCsI2yRWI2tXJx7M3nIVpgHlAii7sb96Pjawe1FlZscqyC0FB+0QZKS918bMZ3G
JrHqo+ia6qoTGAucJYE8dr3AFGbuLEgchkImr/N56b4uilsFn7LEM6JwZP9iKsM6
KRdUYAKFEqMnaUjWn+DVqOHv2ToW5NAiD85yfD5SaUcN1hX/MDq45bPqcfvwrZ33
g6WBuXbwnv8uNHh1z2yrWR3G3L6uOYIc7k9DfV0dyg10Myz5zQA9TGZVaShbBCzu
EIpXfgxBc45j98ihEE5wY48Dt86YLL+xpTQ9S8uHQwEsPxPrXBWslKc3R32vsqOD
WgrRfn1ssIFFqjhxUB8hgAH8ewqZ31+uQFeDRxy0bm/mFakgycDMrBB4TBUDecXs
shoRRDC0rOfPeK2Dab+2omaq9aQV60ab0XCLZVD7/5ckncnWBcPLzGMOt4WVDTxh
lp1ssjnUElsbNRvIcyjPJErFqoeO7jUdZngWlNprVJ4M6SWAE1v6DW2+ZN3au8lJ
3QE/f/pwQfl8OlvDisio4DQOe26HPp55Wv6QYXX8PYxiWLqSWIvNYUZRoHUZTNSZ
GGbOTcloQ8bs6ojk9KWGpq5l0qU69HDda3/yYvR7RVQliyMdzzt+ypj3pyybTzO8
WpeB6PBPuXBT+1En4eFQAohrUIFWLRwrmazINeNvGQdsda65tMxNw/0R3KNYGVb9
gVcJjUVcfWteT/wTwL6V6vSW/6N+zo3HvFhMeNERsQPyD0pZyv7JJAldTnR+4SkP
c3m+XPHISt7bqHAJWbmLe7GeFlvYjYXOcOgHx3VQUo29mfZXSJrZsVg938K0nnNv
9MyKnay3IuacL02c5RNxqLiTzpyAWd+soRCdaa188SQNy+9W203RK3Q3AK9IIF4W
OkC+8SuL+a0OoON4PIVywUwbMBgn2sEF3ZSAObvHkmDDaiQxzzL+x+IOy66CUqYR
s1jzggqoCXrOp+1khmMziSHXIUP+Z8DuIQysoxZ/J1JdLLnP87m+zgUor1+MaFf2
WCOcoiHmCOzQi0LtRAJ9mIwN/QW1ZJGN/0TkBG3n6GB9F20C/lmGZcp0j/RaYd39
jHhZ89AfAx1Vtftff9XxvUbsIwjKmPdMtm2yADZUXXAEN7eWDoqGHgE5BrCR82qh
qGXnCf9XSllE/CKmFyvQ4WOkmBbkEt7WRwl5UdI5B+igvqOb7FnZ96AM+gxtvdVu
b16H7lY73Po6hvqVNNe74cvAoIXJ+opypSan+eGJKz8i8V4d6CPDydwUBni1YUnR
j0C9sfv10l1X9E10SSqdshaZo56JJIsh5NGWIeP08ABfp0Ma5hHIL2SmHUiEQ0g6
FYgRXqe3l97ZXkFaDhftc49StAhdICiX0E5xVcg9oZqX/38ohaYu0cKpTkuzjski
NaoXRDPIiaYTZ6JZpxeEEmJU9I2Zocr8LVVgodhbyL7k2mtS2wCa5g/+aHP6GFQR
A4QghjAwJPBukpn4guZjHbtQwE6/02ECNRaAo9PnRfLZn8cYd0pyq+5ldC2LCmxH
ccUhTCYnOAq/AoUesTFQJDdh6Jl0Faq/PpzWkFwCFnErTriChcUHSQ3YxfDv+j0f
ovqEUC6tb41dnZuIMCWbTIhhEU260zP/2We0LV58SWvAawHmcK85PLEQQEryj+pG
o40bTug2+KlOqcAFw6/Ov5RDpOlu2GTj1YcJgrfnHldKqQtC92uLjXkLw4kGXehp
pzweEdbaQSD8fO4uSqqTCKJzBApf8V5ENHVManEeuumbW7ZHMMpMOkHaDE582CRL
8xgG0fx+g1VIyBU7cxg9FoNwO1BZwB+qAKTQywRmJO1ddJWbwIjJ+CES5/joryny
Tdtulnf37XFxXZY3gUyZWbg0aakAd9HU4QxgD/U61nXVGh+D6v/PgvF1AWzEEGnr
wcoqkeGQMj9syOvWv3xUljxihMjThp6bIEenQQKaTq/11PQg/sE9NLBJJc1JldKy
L+gvT19wvgS5aFr3W9TdKEi2eUUWY+dMXLC+oDwcLkYifph51FY0GfS1oyDiaxK7
OD72vXeCsRni71x6Q5xh/Gh8aDFJGOGVRTU1EWieZtIGhkiG5cSvWMQv0qS+TJiW
wkT0RWQQ8fzEK2z0zY2EpFWihoC6tUmz3TvzqCj5PfM/YbIc4BxK9ZVpPh4ZkIlI
KfUaqtP7hws1khZixhxHo5AYxEmgWUMEpoDl8amNU4s+Zv4SFKk76U73rz/o++vH
CsmyvxbD0mL3pFUwrmQ3e2xefk367y5DQ5Rwg4VJVxouWvlMdyCCx/EKvQJXT2/T
T+c5fZMar7L223nzmJT9uT/HKsk5YNFvB7bqxJUi1lOk4udth403cBK6YWWRyOn5
kbGwlCpAj5IyOO7NFRYdRN9bfeudSpZbGWgrZjc3Fowrmj6b1cNsPISUb8ZVu/2L
0P+CWNdH/JBPqtpszTWAKD8XBCN4AnJHwNVjAFJwkOuR7SmiDusDIIgTiMWFDhP6
vlt8RnMZIaQWRTZHY1Jgf9jRsRUTg9XGmY+HY7gV0zXoKpG+8MQhTre7GxTs5kb2
KwM4DAI9Czcg9HZIluM90kWzhks5qHXk01OEwlwTePYIoRGpoXRdPfWEOuaFwdvN
InOlWELlfdACHAe2f9rxtEwt/JMLJ8OZ3xeXq59sc1qMWml//nuHQsw8jnBAi9DH
aAFSGiLnfJlPiR1qrP5lYpkyv2dr6UXnm+I9vwEZcEX+Gvh0W4z6K/6VSnxZevDe
9wd++rkKUWYO9o7c1jdQOO3/hnqFckWnfqsi5y5hDM97dwWF94prqskKzClWrZms
XaJKArZmj76W3vJRJR2vLY3gzwvtlZD27vvilRx+M751MXvMsfgtlWq4l3o3sweJ
qOgW35bD4eQEaz0oHfrkF1nzQg6WesGRbzM61VUPjGvXyHeUCNEE2WxMk8GHVCa2
KXV7wz0cUVJz/VkQkIobxg30+N/5GvxoCyyYYomOAefXc/LbjC/FIdQIT1dKu4Dg
S6MZX4jubvYg+LnM/KUXFb1hyUkB90EiqZveui9IFeSoyZ+zuruRxZH82KCYYvBx
VS03gemgHpYYvOi8xYSASWsNz012FPx9St/GB6B9grZEfPxJPtBqj4YT+7926WLJ
n7iKlSo/kemDkAca6fmS5LgkLrLoJ8xmpR9FoEAhiCeXTpbAOWlGCT1YPToQaj/+
MrIgwpwTAqKdazT6L88P5L+gU/fm+w3LzS7iINr0dbMcLSYz+5Av3lbvF+6fjVLW
AlTrpbXiZHSk1C1RlZiZ4vvXtP8LzVMKkj1L0ECs0sZ6/MMDMMYHKnxwFwLRs54g
xtw1PcEHvBR78UvX6d5k5kB0/Pxx6MCbbV2CRyjv9TdCIzyYJF0hcXAl4dSRsXiU
HD1bUhWbf/Zzo4ZSRRj0eXFi9SzYGMJheT+YYSad7VmKW3v7MYLUctF/eTGt9SQk
1WQQ1go1GqgoUNf0AflHQA+S94ae8o7X/axfSYzaKpw1XWDeU5j1Eeo/ObvDXRqH
jdislzv09egprR8IvB8QeH4IZ4MdvcTiAp/N7RSnG/LYL26FH7OYLxPUSP2EZZu3
Z66fSuxQLy1lH/0+Mhbcup4piCQKHGHBHD01JUDibY80laLNBbPtVhVDVPa3EXUs
0pyM0KmptWSu3INybexFGiEtPZHT+CKQxDy/VfpHiQ0/1dX4gqk5cl9bcySyMQqO
9cKWbWazRgZxPwtFij0QunXkCwxceed71Bq5bdD6YpQmANJTlsYQn9BYHI/kvzmF
7K52XirJdq/boR/KDD8PdMw6KJZiZYh8OAXrAyvBgOyYZXo+C3fxwEA2EfKrfkcz
eVrt/f4isN7DVe33DhwTPR98nZfiYFWoM1K1oHfvYNZtYWYrnWZ74lbVgwVbXNTI
uoMji0J199t96D1w18iMctIkv73ffgOmOa8ypABvRGUV0ru7+ozdfVWDUOLXChgc
u2VxUa/DDNpv0gmRcUObenPSTjYGOkKMbQInT4FgErHpRp8JLSM6XINBPv+izO86
bttT+z0SnGYnCzj/48MOApFR8fJuQeBzM+l1FlRVUqySyRYwun3JifgygFa28JXN
28sdPQATJGD5syqhD95n+OdIgKoBjUSc8EUq5L48XFwAbrGuIbwWCMWQEF7dlJXK
BDTGDHNBoQRChybUpcNPH3K0l33o0Uhy0FHjNd8tXaSeNdM2sMYPXAB1spuVBFGQ
4wiVgmkaA2J9+KYIC757AFPCB4UUaH1H7VitpODuJ/v+A8ANOKOQqMDGr6br5hJN
y0GymOaEuyKlsrzmJwA55eWUgZhkg3woVJpP0pazDbYonXgISbvNwAZfF7lv3yrA
DsB4jalo97ONrwjyZp1+35FbDhvXKM7uqgc3U2H9FLBABuUlYUouXDeXW98/dTuA
AkmoEjzZAmZ6Ujo1Awye7di7g5shJISbUm5oHK4mr/Gz2demvB1QPL6D+jOZROsZ
VXLOSeeL1om3WA/6zbbQtSDqlUReNYP9+mLovvFyxph5Q9zTW9Uu/D0EXLPHhFuu
LBbK/zTJgHmYQraHM3ocPH3PTQyIDeKY/Nu6rgFWsqYJgB1onMJTGGcLjcENOV1R
i8tbI7cIkAusnRNbH/NNfgcW8giSyEW3k4B7+71Sknh5lbya5G1CYrNMx14yFZ1b
Aq4SV1Jf/LTGtZp23iAiqk83wcuC/OWkL/3s6TdEvrP/2+/PWFUNjim4eEq5X4wC
lYNJvupANd3t2dd82HS7++pqpVxMOpkz0n9eMeT3XRgyS6JOwydZotyAi1fJbpn4
SySZuqY8P37lWWdKuBxl5nDeemBotuFCWOt9xK1FnZqs2lzgmOPlFP8UwoIwKHwL
9m0KifdIuMD0zjzd4RFNE+egTfUkD7FXGQugQM7A09jZTNBcQsE7K7LPyMnzOfmt
2bsZfFYgiIZvzWM4YL7fGmTwkN9lf8eJdvB11QKBi9Sd2c8N82Xk6CgiexU98q5s
NlUr/h/aaWXhwgwwDJ/Kvb/EcNfn/wS324XmETQpGgt7ydEsMjFWhFBG7okThT8+
pRaEQxQg30RmDyXe8FpcVfBiCWLCIdv4FyvpS1JiP75Lxa7rWsH6JgeVByCWO+5z
tVmUlX4itX/Vnm6VC2JYL7obryUE7CexURSWUH1suas2SMhKU3A7K3+HTgBZOi30
EXktdtli0ClByR33we2crSCkbPmJGu0MZq/Dwr4MIMpqkWsqfE5SONTsOI98+PSI
Xgoz2/4baBfT8EtPZaca+PQpnP5EpRtBQhuVRgmQGWAy2ExEkJJke9sYrFwc7vE2
nbOcK5pCYJ7oxbPJgN4e+9AyzGkSwf5RFQvI/Kbbt8dbubyxyC7n94aF24oznw4U
H3unTn3jLcvgLO5rDUQBFbSAghVudwZxTEby3LCoCdfNP6DXXw5jmOSQFRxv24xX
+c6Ub0pjGTH0EkOfJ1nvjJpmDeAUzGBLPzdHUHcGdKd1T1XuUO5tvQ/IzUg2G3j9
6AVui2dM6kGCLBEDH/n0KRZ8BevvcZI7XoAcswkmDwgJ59wdN2iqlKN3E2tIgY5R
jdKkdgZFKWhXqn8yaMHzLk010J4j9Ty7LgXWR8sfTvtu8OJbQWfCdlfHmiibDLXW
WLYWJZjEI7bkxCBgZGDALxDyNagZHLXE5sTYPiT4Q5wngiIwKExolgP9pGhYtXn1
C+p55jg2JQyhQZFRiN3JQsAZXpe0l1fwn4L8zen1IfusbZRQLdekgsiqIfl09WVq
Js37CAmgtJeeziSAI7ApdmoVyzjCWnGX7k5/z8Djc7YbKc3zY8h3DjVfGWUQJN/X
xL7qkfHUKyrEJYQytvVIIE2zzxREK0khIMQRXL5pqAt+3P7avVAewtLj3Zauh43e
E7kNYzS6KqJEOPJhmnZ1fRAjvRiMjikWaAxNWBNrIxKak9hyjYmJNdQCpFWxB6/l
wguNZ+nPHgBu7gLi9FYHNWvT8aa7/omcFLjHwGx3zuQfcTXkm2SV3dbhNfRhq4l5
4YD4JCnZ3QJ0mTeblusLtYsT/MMHvGv6klIViBPjlz5up2PpvOJzqoW1uNzPufu8
bmIbtLKjOOu8lW8VVfjwlKpfUy2psSeFzgXeHhn6EVUwvlsTKaqvGKnsyrMcyqe0
jf/tQqukB4H99Hwu6Q9bsOjshG5g/5rOLYuyPwmqtlviDv32OtCjRaboBE22oMtJ
EskrA3RxIyW+zyHheKxQkfclAcFJJZgtCzt5BjK7joX45UJpEE8E2eBUTsfa+XIl
TYCwAWBfhM2dqu3PJBJLYRIOHHD65WoXgmSZwbGIS3Ic8SjOtw2RNsOtAm1sk5un
rIXYLtjPm/ahaWogn6yy3U7YmWI+FRX5hR0g7vQq5bBB0eQ7oMCXyKaC2GuFULvF
LrcoBFuIPqzoNg0xeTCfWvyodM4Wl7qR1opaxLOtsMlFN3yYCRCnDNyW5bbbA87A
MqGbtXtxY7JyK/dNZbNGxUbdelQjwKkr+VN5fQI4CX5iFyaoPizz3BIhbvVcw4mj
SHtlPfuHNpJzouiAlxKHWpPM4WunZZIfCjuM52viMCG17qILNXCLj3M8y7su+QHG
XV7QAD2FAL8I30q7yl1z4cRpsEAGeevNYU3HFWOoZq5cDrLHgMAR74EotSIV4BQW
MnxDwF/LakPhZ0rpEz78aI/kucYhCJQYxaGJB6qjYucdyR32OUTeAgncYEv4vZxL
JEMoB74pQE7BfDrzHKpq/kcw0LPtgT5GzBDZiFYqQEs4NbatLVjy0jXT0uycPjiY
g4UV66rhsLoXqEgV4dbx+48l8S7YfMZEbjjUmaeUrJNpmLJWXdhXjgRatG9IOcNJ
vGRGRPR5lOv5yI/QBKmiV8v3bG30sJp50fkw24CY8ARGAdn9OT+1NhRPqo9B/kg6
WFOF4sCThicLn+TTZ+l1KgDogbrex9A5cbl5F7ji0I64xtn0Ty744rmXQGJkMcC1
Fbc+1F9v+CwPkIstwSVaEqThs8h57HtcAW5wWuROChImBpNot/3yucEVKsgWkU0u
nYzBmCJDHneX71dMLAF4gRPeCsZRDHvVSPx7p9nwQdJYqtGGEIUtXimHAz8Vs6dW
cfpOl8Y5G0hg72UYneIpV7D/N6p5/0rI08LJH6rZVvvfZC9yhLf2+ORsX0/5JMjc
RLmxOBBTmqFnUy/EId6xWV0YSiVGDirSOHAn68VKhjsdqoSBHJwCys+/xY/iIRwh
xv6VXXAyqI/4rcJ8ZPVr68sRwoFxy2LbtGxMFeRQDbcsOrkj9Afx6qKnrLzNdnyZ
raWhrcabjXfVyNU6syVW9vFKMlpCEcI3vMoytItklQCG7AHhdYAO4Grfdm7Q8D8M
bIgaU94XucTHzX5CrGdcrxCLJLFLnwM/u0T7KqUb9d9r6gpV1hVT0N+5OzE91WMX
S+VW9FqQ6iBXpO7xU0ac4WE7bcXWrAXFHljuhrTDt6XAVKwgvVcYkfRho1OFjT+Q
/n0fH1w0qR6hZ8sOdcjQjfWCFNWdHg0C3nSdFV17QtqBEuboI3eIxzvgDWTNzDF8
WKKXhHPII0oT0CluwqqPN5izjqZ3HfhW0rzfzVYuhqi8nMdBQ3+YyRrdqX15Qa1h
HI4qc54r+7upB0yiYO/Dor1DGOPOlX1AhIfL7WIY+qJIZhdQlJyXfJKk6vAolm51
K9yryf0PgltezSplewaWnrNcvrKtnGefO/O2EPrYG/Gw9SsiazherWONeNxeRuqW
tRHpe6p8okUOmLzh0OJB3h+WhhFlugAUYRirLKYp0ST2QW2A59LYB3T0FFHEmLDX
mgx+CK/qPL4GpztmabixAt98eAiGsxeRPfYpIFn6lVYnYx741VYagL7bRKvfr728
mic7scghqxZ2n8ESqvrc1pw9Yrn5YuuZFfpJZ/p3JSei0tzJvI4FzszoGbXslM+B
HShVpW6FA6Iidu3j8LuyqZqhctrTXN7dsFsJB6aRb0kjoGppIs71fpFDdpLxMSPj
w35wxS8pJEWm71+AOk+rSt/8pNDJJiyNrWzPCXDKLPC1ntpYdoR9klpkYCE5IyPC
UTmmtfy9u98z7GtDuAWgoX7wdGuMYSrLw2SepXvjHqFX25E0+gjd2WLYXHP0bXY5
YFXficBxzW9oAI3Xy8eN3Zg+ehVYrBYyyQL+2yp+6g9NelZm4zDoWp2WzXj6FnqO
vq136kt371FCArWyqA81SKeqZCXQxYhpUnJXb/i50h8LsV04OlfGRME72/l6GP65
SLsVapr6CXtuI1Accf8tKAAX0ltjjzHNRBHI/cMUScSbS0b69iX8FjKPoGQx/p9q
X+xEt6Twful7+WJt5Cj2/TkKxa/2U2Wpp3TwrF5cLMTFgWjkRhiWyk/ort4/+gWZ
lNS1GvYgsCMwC+FGORV0QM7PqugizRYLQou79D6rkxe92UdU4KCi8owrxLM3VcqP
4GSv5IEvguRA8uty2ALBXeVIeM1kN4yzfQMuq75elf7dhX41oTlrHYvKoOKerY4S
YrVtsEYFUc+baZbhRyInfLyQaAhyPFYLaJfJc6feivmeMWtuFQZKZkDsy+P8CRFp
7KxPboxc3ACWULM1sjKNoWqWMbhmU69wkozvAGC6LyikDZ/xph6nPj4s/eQoKnJS
o7MMxo3X5RYZBeHhSK36s8o7wNTPG4poTNlWLRG6ZVwkFSl2O7ZQmOgaYnghRgJb
UoisE4/6Ht6uusSWPjarUtYs8Eo+hikXamFXzvDYmmIqRv7L6Wp2Bbx9wwA4d/NQ
ZUZ/YdLJkqayNuxjw187E0GPKGm6p2JkVsN80HnDYVxAjo7eL3BXmplm7ai7Zwxx
M1lOtpsHkIx+j1eB56wYHzoLT6i5EH0mSupQabaLR8n3tqVnlsc42LiGzf6R3LKh
YUXDGik/0cesocRENFpZZGEv/WAhYRbOevM4MLX793hq6FZCFRZ55oJmX30WvFwW
HoKcw3eX8QVfPpG+ddrkXYYVp/mk6EfDw9k89pQTaIieDqFnTpo45YaIUK6BWYfv
krpJrhMfim7ih1XcaDrnEdUlEQ78tqSMtm3rdDgoWmoZWs3jrBef+1yCeBUhh244
3z164qLZeWo82VzuPOvnrVyoLzyAB/nbXiDBj6x07XbN3KLaLxerrMg1cXFyBFNy
XKumnHDxmdCOv8OP2oCrZ26PYhCWuGs53o9C6yMUf4uAuVODxRW5N9ZEoPRK+TIH
ssYcfoq0QJGZvusKi2YJ8PZ7NgSrh9bfglbXqrCazcWNuJWGrXT5Yenrmasr2Ono
79DzMbxEXSRzdcthOsUoj1aAUHOlgfbNgRnEHIL9GBN2TDTl/p7lGhId9wb+bXJZ
+BeEc5ELuHnLbFL+G5/OuLs8eSm3DzQ+vSkE++qvyIhJNdEXJ+y6od2S1Ttjqu7z
83sDel/Jtv7A9T+uA7U/r6LcIFOqR/5FU3Ya4zz/7kKM7nr7MbQiYHqOeMlj8Au6
BnewNTFcF2mAwDXj1BdR9fMUaZqJH4pDyVzPFxsw93npV7XIvRWHpQWT9kYp/xeY
k8o1r6a8f/PpJNyFxchiA1om4WogRP1UvwcImQ+z4CpNIKiRf7C8jO2yzdZX/W8n
wk6+zoi8wVfH3Iyz88qvqblsvFOwCvn2rs4I5mRukCCkO1qhxP+JoZcZ9NhtYy/S
7uMFNC6QmcUUm2Uh6aivPQFFNqGZrLpT1XHRnZLaTYgoX/mIiB1AzDpOFHRkJxSU
CArKFIgKhpl+zaYOHhB0ZXbmNF1ywXGnxjQLipv/rtHwoZ22FXUwWOKl/LcjrGyc
8zOIg+ck5sX7vCzWYamKPaT34fgAWzydr2OGEWyXQ++AxOp9kimwbGp+92tv7JW4
Pa06WmwjrgQOEshJe8mAyV2+OFoFtEo//+ZjhWmsRkAxHuZD+ck74dw2b8ak9P+C
JavhPNoho6IupRPRbW5WzsLzC8mV7yWOdkujUW4Gu12kcevBv/EUFpFe8BI/5Mc1
4eAgBbWul9piVdcHLax3HrJf1fNbEzmkGfATQZL4lMyVeDP1qjX33f+afi2NusHL
tVoLqoGkhe6HE4X+yNT74VbqTdXJjTQww8ptWNA1PDEuNZhq55OOycgjliwvk4UM
8JM1/EiJlwIBfaHvfX0zKN6vderoTkhkxHPE+C2TSmC9JqOWvSCJ1XMZwWIaOjM7
602vlwT2DYVbwkWBH4OUhyo+5EIC9YL0LZ4k71jhzQaTzvtG4iCg5TPTB/DJeist
Kc7YqZzLP5YWxYkuEouj0tWtaUxDJwqMPeEJzQLvdbtt4TjB55fF1+ZkY9NsyoE5
YvHPHruCpsKp8R0X5nkGrgkJHKFjnp88Ockgci2F4OxJNVawBx6JIzOkv599J+y1
EaO/R2cHg2x60TKW60ytrASRHrVxF2VZa55lBASOhnDu+VcOWfrqYbMrtAbpxhaE
dhIYwGtrLIl2cP+ICMYrysN0floOjPKYbktWjfKf91cxQw3wRgevBZuKSFp3tut7
JKZbZfXgFjt+pGuqZYvCw6fHto0+NPigfDPnk4ScmZAZeaSDPEhcCSf8Sd5OXyzW
avjWp7qtQhXOoLodiFDu32U2G1X7R2Ljwg3vHilOokMGOClkEVbRlt40WBq3hn5l
fdYcmTZDu4fjAuwRsNcDwObPEpG6vdzmGuxAeaWSKHM7r+tQ2uuwN+LqmQJqXrpi
eMic8/MCeeY6iwyMRnIYGe/rFVNXTWicP0wdpQTF88CNk6hvEAJu+Hv+h38cTway
j9VH+LaoZiNH/kSw0WxS4/mATFW8G1IsXkCLieZRHiM1sEtIZZi4naRwD0dRTTnD
od43rSVVkfh767cUpaBbhQc96RoIAzyCVfxgN297xPMn/V5g6MXeMRr8a0VitEys
bLtsm6CuspsaTZg36wo2Ck+ezcXDdbNRkqhiOHX+h9AEdr1laBMMv7rZRSbozdma
A4ksbX9KWgVdpxvu5HSUSzaM+B/boldFSwSMadhqRFK4iOEGTxK8aUK8z9my21cQ
s+cOjQzobgWHGeVAssEEF6Jnd2kMBaqptbFMGtxiWJrB4yiMd/eeu5t/wfpfcnZY
K2Plqn07+4b/wm/joB9zGQ60+zF/49lhhJYqgHxdpjRH3+g0S/PqguQVJCFWwmr/
wUxK9s9fZnR1fRUeAJMa+QXY4R0SEoHA7Q8RCJR1zeqw/FPR46zd1XTeLAZxe8DQ
WouEIhKn1K3YtDRvxx9Xa66Y+cZlLJ4B/MxmJ+/0VyeMguxEeTta755vZB2ATyB5
A8vO7mgVfZWbRtfPgi3ZAfGC7gwc2UTYfJG2r640uGZUbFnlnLo2C6MYmsDZM8FN
kYO6wUrhIrKGVjXLyMqFVmEWv78z6xEb5nNxHf174I/o2Wu7JZigQFaF64QkZlvU
2zR/aLSbiG1qrMN9OMu/lK1eQ6jG9IFyv3svF77rehU8H7noZiAYXmCAN+UQjKbh
emmVOFeuMCB4aDWR6rvWaUmYsSADqt1uiMYCNPaHARu+nGVnmp0kYSLzQ1ujVYdw
VIm6sGxKtB5FWmJo/YeUKU8NLECJ9VfWRa/9+Sa9ek+RlvZcXRmsob1NlpjdPiZF
E7FxKA+75l9M507hLGpiobQx6kpkuCIE46rc0Dy/9S7isvlF48h85YQHLA7Im3OU
jr8G4J3xCOWS8a6hnIbt4j4YHJVNeXvEbuW0cmxtQnK3OGWe2VBzXamWsAksnWQA
MYyy+tH0l/eFG9OqPm3kWgg309Er1xhwq695UKujrITXRAv3L10HGJ+uIxdthdOX
Ej5Ad+9XzonLfG/rqUHZT5IwUGhn6EOpDjiyE1lr58O4UK1RO1+nRfwBU3vrg4is
Gj1cbiIvxIDH/j/Pj/IQQQx02yPBA+rywQ02Gt0U2sMMRzIkEbkA73BdwM/pCpG/
/Schd8sayFrzNUsgQahVBbrhMZoPUBc7+MPKq/oCr6WaTj7URzdmH5EYhoVOea7g
4tstnv8D4xOWwnKjvEuavGe6AkFsjc95ae/PIRLPLz3DIPEsrVWJ26kd2RM9tmWF
tihHEYOgDodsUS6sPCK+HG2vrH/YlJmtRUtI/0u7rwTm7aERqVr6g94mSF0Rqi+3
/wk+2FBOr1/5mAsEijearZJbiY9ik6K/o3xg/KUGpYLAa1s/GTFtkHO+RXlNLJuJ
hc8xUEeZyLv4QabIap+ywL1biJG/2YmppyhULnVgCetp4l2lnzh0oldO2bdjf1Im
xKdyi9tWAbnkZWk9aOxHRgTeKd6ZBnUsOZcE0Fr6OQPjqCc3lPWvf9fke3o76EdL
H0AgOgen3WopKvqzvs2YKH4JHyHmWJPQjHtZbLtPUiGT4+WbCeZfKMhlkLiPd7vs
hqoY2lpDmXYaBBz9kWKjMUKqIGnx9zMGF0yxrYsjaSqgXMA9ZlfR/iHSXL0cRuPJ
ZW0hZiMx8e2YCUolZqBsSl1cTgG1GDx7AO1wq9tTLnNEwqna6epkIza1OHBxux9/
5Wq+2hCh/1kSL8qnfjEwrRMuc4IuLI/72+T1/eUPIsGHOnmZ115HKPoZMq+gfb5v
2ZlkG4PaEHgy0NnrD7RP+nZFu2PwgrVmwMjsrEcME9ewFwTJiR/otj9oA3OsavAx
7Iv4ac971lpvjGRk9N+gods12fsX4FNkaw3xmZdhCnJPEbsYaw9imCHVNWvz7e/q
5rZs90YhAgDTFnaoaTSdNsmhsz3I84N4nIOpmejBmmRoRAJk18UPTLeMWwzkqZkt
rJZ3NbKoeKdjp1ddBa26pjXefMNwu8/i+Z6X/aT0CAmfXuzlwcjidsh7PlnzcZTM
7SWNFyMuY9lGvKOUxgUo9HQuKOzeMp7s/tR7qp2HN7vcBODXyurbZWsmO5vOn3r+
noJGRV0tam1PEQflIVPljvo7Sg7p2ab1j4U0/pL45i8+d1dv5dKJ8WE1M6cj77Dl
F22D5mRBirfFSzSNIHUXbCq+GejburrUlukZjdxF8+ODonZCS2WXHF+MWt3L8e4N
YHdzhZgc4t1jrRgZPOaAORCOWDi/LdW6zyankWHg4AmXVDFkur+cx5FjtiATGx5O
X00hqgOMGY33qqn8skW/CRO5MoWi5TsygfdZjxNsgpadtkQSu/O2leAOmR/AKcIx
3j32KVnmV3oSfaZtBOdhQEfbVVIHdnovn6568ZGxnJdale/ztTwQTmkcf21ssJbo
ts71+oooUpTACYE3jvtQsvALWDEi9dBJX63GBsjE0FWV1Vl0H9TEACun7ghoR365
aD8+cGM2fcRNpfZHJxKQXvLC4kR8By/SaMV4EWXQSmt5FdolkF4sWug5kLo4wFtu
Z58/2TetoA/UVhLaU/5X6o7YWjGu3LcvCa10HVgipexCbHNm2afwsip2yu+tM7ID
9QfSwpvUyE8mNFFCOflapmESwiCJ/IQH4m+CTZ7pJCRkCuXRnU2cZ36I0groUIP1
GDpd+pN70iMWf8hc2BBuGehRf3AtnLVbOIjysGTQPl1vDu9SFyY4YQiDCHOtgxNj
X9xsBjf9txaptAcIBKtqJKkfH85V49vyyHkvEapbpPOWFtJ59yjVT1DZmhDWkCv4
P27ptfkvtRBFV6p3JHyrH4EPOP0d+8uWkNx8NNnyS3uiFo1ZG/3md6mHml9yDCrb
iw/FY/vPfwwgIZMl/li8UzuiLM5lkGsZ+3N1vugCVE0gF2qzpgugz3L+p2lkE7A/
E/n50hveoXxzOpHwauCc6nRN4cSeNPFrgtesqAQ/K1f/6wyT6IYHwTYXnyWV2AcU
nZmHQIMHKxtSkFQ9pa+ipGiQ6I1okQE4/rLSpsIIKVbL13IGSt0VSdXybzmJjrj1
w/8Rur63iNqSFh3CL46XOfUghALF9XRPr9zgtkPGtn/Pakf0PZq0Xr2Tys/9fczI
Upa3eR6ZHlVFEmSWECuTD6Czpgwq5w9jFiEJ5IctWtd+HrJq9VWi6jEqByXsiZ7w
ytph5bd+ixnkMhbesaqNJgBXBwLyLPp5cddeXAwv+KJqK1raxNxMBRdctCnXywov
IUAlCsbo7QJ26j3nECMj97pQY3CaU54nbgpGqE9iul8CUYHkpO2j8BWGthg+HLo1
xeqL/StlIxOiuWE0poPqNtp3ncC9rfF4zIQYdoiTIomUkgqz19A9XUlWzC25+ojx
EBe0El4qne95anFl3TMeZJDTA0JJ0ykSe1u04tbn3O28S3AXMr8998VcLr815teT
3eqVQTqmMa5LH2MX5vsvilcWqbAMFiXToaf4mR54rczyl2kjXJ+gv0fgCVtQFbEa
pjsmRV4WwHl1cMGuf2TlR9JjwG3DZHPCie2h47hkTc7LgQIQSeMyTc6oJKdL0qMY
JnjAkzhHdzJL2zIAqrFY/olDn6C6jxuk7QJHVDW6OV9be9IzArRHpFPkE7SIsFC9
VHRDqv5vs3AYmMCGO3fwFkwwJFDFUtMxk3Y9xjCwC0y+CCjdT/Uae+247f6GlWra
T1P6dTIR/Zjoo9Ke0Qn6U/ea+LcEuy1+HuShhe9TjL4RZNtL9MJ/mlCZw/VFrnp1
UjpaKvYe2J9kBtig8x4xrs7VHBo5cM46ubsND9HxDpm+oT1h9S5HTa2lvTB+9pq6
Fyyqyade24PyAIrBzF4SHFz/cNrB3G32Oig/zgtmZgrdMGv7FKhgvc5oCBxV7NeX
c1B6nTa8kAWkwqMDPJIqXQwHWcwodv/PlBNls9Yq0SWH1PlPbgpYuqNEfknAXlgz
V0f96wf9A637Ww8mHdMVfOdGhh5TgkAnQEhru2SsldYLU56uL/xD82oD6wnoaJY2
orLs4IIngXR1zmMgZXaR1N3mLAdCkWOBLV9HysolxutJYyIgVqud1dmllYLoQjpG
Yx4cB9aevDaob1/f7P9vax57E99NdXpTx0l17qRu7yUPEU4u8BR8InLAAnLOmbNh
VBplF7SPULEpnvV0p4jhv1f0460EGcM122wdXx/Nj5m3lu5UfWsWVakM1OeHu3G/
1hBDAKxv1rkJgayZnVLhwuwvgRNUTDSFyd7n+CJKI5VZkxY8dWUAZLien1VrrsSe
GVpfmDkViVrgUOBw4L5RBjKBICBH893DV0rpSmB7V2h0L5H9EjYM0YnBQt4njaby
Re8wgQg2maXDk5uCEP6VYIJYHcT+UTiQFxTkp1IuLpc7nAOuSaI2q5P4FtMD0RE1
PEOo3z6hUXB7mlDBoVCBNNp6aBEKZ3MmynoeAyY1rePwC0oZXVhdTD/6nUwQF90P
ZcP+NRr8curE8Nhl7HQ4cRYaEsKJ87msQwg9j0/VZZ0WouNmzYK9my4vsgiLulpO
yhJ+clvInR4E1JY76i9PnWdA9ozJi/fWXdGTZHDZie2He4856nMA6OZufa5qveyy
xqd3WiAGdj2HYpYjvz9HJDX8Gd3dqL3gWW3vWUUb9Tkv8q71ThyRIYjpG6QdO95d
H7YVjeQm0sbKGja2vGolU0PXjolHZpIZXP+D8Odo62nD+YPkuS+h34yoTr57FBfz
KTA5Kf7x4SyCJAJtC8SGtIgyXuJRMzwduSnWgWXNAqQp6nhFu6NSV7/0oWMYJniB
XOXbxh56/V2T9+M5rIKZ+JI1qtMnRyjwhBrKItcjxDYmcb6vh5mTjALkgi8vd65t
CSrdRLhDBThl2EtSEjhVvdDtl5a9P0NSvV9CxZaoWrz0rZLWZ/Y4XdL0s5yxJPC8
oV6jXmPICsZRHuz+Fb9xIi1clnBpUVD1rZaCdQCJcLIzJDUn5tfNHzr0TOur6dhb
yJMT6OIwbsPFSu17HOK+gwhYYmo3gjHEBi5r2T3lkfC1e4JvXN9g9+J+4yhf5yfb
C9o0DqBexLmMhynrbs4rlAKIAX96YLXDfaEc0h13qLoPnKwIascyH1PRWLGZhKQc
LEuKY3ZXUQrzH9T0bgOGNqAVhpeAiLStZUvP89Rqzdrt9FRVHOhxXwN7E/hwyQe3
w21HgDGRALNwWVA/n58YK1Bg1kLj4YgCCjWoNPRl22yYIZA7fgi9NEPeRYefUsz9
pT5H4a8f/oV0HiozH8wfonXuPeoXieHO22twD1VgzettB/LdJ/mWUV+e5wctKvng
2Y74Bn3X3n8PSlIXEZRlT0qfk5vAjXjlgYFb+uXPL8tIG0RvxW/uxkNzLb4omP6H
XW7cvelul7zGkepCZjIwewqeWNT9U29aRkwuIxga7DFfGGT37KEGcjyDlCV3sWKR
oPAEzH++ld/RdsKXIM6le3rbs0CwMOktBBQDkOWLcHsElKHkrkoDYVxfQV/EudJ9
Iufmj4/Z7K4lQziuvc7dDpLO+y+xcW0GjHz3bB32kIF+kNdEy7DTz+NNywWerc9M
3NVdcaSQ3JxRPE9fvKOeuea1FxPcEGP3glHe1iG+3/XTZyhFYCus1xULxkTwkqw1
yPAaqt3moSD7bSXWaFcgwwoMrZ648Gvz9QXpMQNal3oQooE5bUueaeQPycG6ECvd
ya4j45B+zDl81q+IVPUuRmOpAjDi0M/aEuiEpOMdEsvQvxrhUy4LnyvsPnUs6CMj
WsffSeSPf5cu5rLbtsR54a+8gkZo/qbJ9MDDUil+7sAp06Satc2LEknPcMrv7K/8
24H8QuIBg6DV+aXyfYeZqtAh9I+Rq+6z3aUUbS703D8bL0bSiAhbHBb1es8DKNRH
/FZ0qM5CxYDvEWfAbXm0RfOm9tK0YQzPTUXgV2Rb6xZkmZefzJAjN6CAv+cdeKNQ
rfOK0lhEyN/mVkNb1HzSKssnh6+FGLJ9yuNybtmStrL0gm4VUkXE2GDESQcZsZrr
iZH8KUEB7Jertaml0X7n2PUledzmhe3mfM3VKL211/9CwmiOxFjF5uBvUn0/Aup6
un4R+Pl2dMzkAL+7QZB1B+3vuOELaqt9Hy9r9BSKL9XenfQTCFyWfPve1ZFdxOSS
24RIGRgUWvRmMnyLHk4R6aQR7AKM/8ilbII390IjqoyMpwgalPI3a6s/YjX+fIm3
uz1ESvxz1JdQ4wyTW4gNe9Ida4LFS034h4CC7jwoj+a4BRv7RUVEwryx9HPIEFYg
LNtO+Z2ST++sp3rRDie8poQQnQLzmKAzbLYMWRIJnpwfYuI4auixjJJSa3msqodO
g09YQThRTzhfxaUMrJ3d0AN3DHtpKrUF5DCIDQ829UffAanMXieNKLSS951xzbpZ
tyUZRqRAIsLqIVFgOHMKrpw/Xp5HSpb1eJi8FfC63FwW5KAdMJ7tYcVMkdHflA8H
tOlSG7KQ/DJ2Y6ldL8xgzGQd3BR6gTecHMj9W+/od2+APBL6WJHJHEUuhN9WHH4y
/5gEqcIKXwpH3hFS4JMISZtxnhuDFFEDasrlKH+qMnLWoBsE/1z9HGdEipHgxltA
tRyVLwEr5X/fi4iWKWNl6cIVQq2Lg31kLY0+HWwxduMdC3kZdl2YbDjNgf5nxaBi
FAHIoBWJouBPb/XH9y1cxbAu37C3CUpQYtOm2lwKAiu2zXV9OCiV9qn7vAUAjlxe
YvrOsm8+vzs5F+fRjvhGKft6nVyTHYoTb6LUCd6G3epMeTczJbGM8q8K86QiuNY/
O7uMK0uLPf4ZkTNvSeWpMV9OG7OI00K3yy9UkoyFMS6gY0ClUB3Xq4qpkbcTCy2c
y1a5Pd4o+iBkt21x4AP9lubag39Vx0grERRDpARjbsLekGqQGPeuHRvHxdGkHap6
oqJ1s2zJgIidGAAPSxj0MFmvqG35Z5iA0aLKO2PBemAnShHA/wUuD9aYHfjaU2eA
S8xBujlexTBN1DQf3cF5ISg/WlXliWqgnyWTXRFHmjjBEAUztwCUbIG+ibJVoOE3
3fm9NXz9AHX0l5RO+FG6CvONVueRpoljQIFY9VEwyEoyXdj4jBeg+Vs8LZW+yuRq
VpRl5uvUKC2Q/DORvM3RE8vlz1Udg5f7UCwgLBWXi1+SL+wlLqFrSfCK9gfF/n9k
L5spS7CfC0ecqXm8roBLp1U1VLCwNg8w7v4NefqBHUm8c3XRRJSstP15zEy3bjDQ
Lz/GPfEovrg49ATs/+mJAK7QREOzkW3vydXimTROJpc9bEZGKpPD+Y0xrd2ATHn7
sIAkyFYJjyCSOFblITPkfOuOHnZ4lemtnIX9j4vo1Ct2BKNVT83hVUpKMGe7MvKU
nyid4jQmDGFxyQ6ucNgt2HyfiCrdZlBD3bhjoHkHk7yoqmu92QHMeRdk3IEMAuP2
+mOnBMYbjMBxIeApEgJGDf1N8ZiDwYYjdnB/0KNv/IYypry6255GQpZR2Miix/Cd
xmPhA/rHMfvKqrlGlRbEphv0zde7D5xpW6Cn5l36pbBYgV+B4gRW6ag8jENiqYSF
Rm9UOdbfTm4YCecboumI5Iq+6ukG/CAHcEolugjOJ70XznHZjrALbeLfLMlPzgV1
P2Ft4y3Nu52Hvu7rxXVTLP3SwKHJfbqFo+uxfZUyzvA6oiaVd5pPwwLgesByHlnr
/pYz+uqFDwM/yp7lEX5UTXsfB6m2BqNUnV6pCOfuwewO2B/fl9LH9i2IHI1Di/CT
8thrH3rJIomxs3TuflwSggtFrEeqhQxCESverTG2MLuDAHj5JpmZefUnsAb/tYvH
so64eWxvTBK+itZ+WRbUisCkOXTMwUj/bI5rHqplHHn8XsU28BKp/UeGspLyQh+A
i0T6pGX2bprnExtLiByjKkS50E931T7IQ1hEcVca2VBsxBDIsBai9VH1CKsZRCLb
FjeUVgkfzFS58nCSzHao/jy7vQl4xE1cbpLmtsNhAKQ9kP/Y+coFysQQBNyBzkkw
wgF5b39Qdhbubg0ftfKigU0IphkoxsOwRhaVuoE5yK9iV2ng30ZlwLiHMfs6i+lp
SUgYhLGp8/jsdqfrXx0Uhaho73YBQvY+HanPGZkNF1FG6X/816rj4EbnC87oPzU3
rdhMJ0TfkUhZu1cD7rJoF2U0ZoPcIScwT5s9HxJuwUScFtevPXmh3z47CwAadlIL
FcdpNEHvzmnWRtpKl9ctO0M+wpPUWoTuhBtNDdpi/QigvyPjwaua4BZHxA+Bj1jq
2ESp/7a6TBvGro1+yRN8lqj0ph4Y0WGR5tLsw/Dj80vLcTxwriEQtRsiPv2vwnfG
aMl/FzBedn2q+Ow7pvgh+C0bE4ywcvKA1lJZKb/TRbn8UXAY7Z9qkw/HXk0Hx8kq
QBnbkIue2in9JovN0vwl8fUPkvDgafPrgnS/7vUTKK9sxGaElIdyVRVosBzi9N8z
8iQw+/Jy3IRuZ1Ha+8EofwFJ+/bJKTwNi8IdaXlG/524AsgylZGAs3eeoNEZTu3s
1u6r0SdTXBzmfr8kaa6N2z8lJ/htvtLOO1TZ1GeJPaM1OhieBIbn+yd+AYRyfkIe
B6NeJ/+3o0HyykWFs5OJT2UCfrnT4MUHGzUq+LzfQ8iQGW3MTV6nIgrnlbkhIBFj
M7mF+Z2fC8i0oUjiMKABEeKIu19hOl0m+oVioBX7QynNGcWYoyqG188ugQXF16g5
jItDMN06vYtGB6pPnw24h9I0ziXzdhFG2/gMMQl3bU61acG3Fzw5BsiDxDYl0FP9
M8bvuWMCgtFDrFmVFafOUB23VM20k2pDcelVU78O27BNlJJ2tp8N+kEEjCsTIUhu
EypWs0W9u/FwuSxAzkuLf1k/mU1xbQf7PCp2REbpB5W9wFjCh+t2ITn8+aHOlRhn
s0WGaNimnmKOKH5d0pqMHWyqXcbB7HkBSXO9zcT2UfsfZVBRxF5eRRmD8QX7Y4YN
PJdZ4dtdLAKQ7KFEqGdQ+ufMh4OMpM24zTPo0KmBy2NEXUvxRM6XYlW21ZYJDta/
IUYlFpPAa4TT94o7LF2VEQrzGcABX1bvbwrKkUt+zSRdllZtjIQ8gOq0I/gFWRa8
D5X4SwJcOp1UiZUgdXwvyEZ1zxVzBwCJ5L92XDzqyCH2LxX2xS/5uqX3jUam35Iq
yUV0u5GSxky82I8JIXdEbMxdxGhxdcbelUA4KKlzAWUBp6wxHogeGStC5aHHD6J4
2ensgJjpCmC+GaDG3Y6TSUfpdvi37taucPgf7As495B9NjvSwSyvZO78iVECtF9Y
PFD1DUfTjOmPcpD11w/DAWuWUZrncMbdinykKuybkHIkC2v3ausPZ/MOVTE8SO3u
PngZ0zZRHQdBR3XssVx1lxqOCV3MqbwIKPneCaPTFzgn6dDKOeSlrpEYWMOhXj9f
RY+eE+WgGjsT4RzmiigyP/cfM/+UyU88mWq3whqEqFKn+sL7FYUglSuZ6wtgOgEj
wmz2F7piyNb+k5YOwI8XU/+zmSY6phJ4r80eeyNQY8PCFdHjhIEuxsKZOOikTb/p
qNWva+OEx6dAPdsAATXG19qIcdxNbgZbJrHHRwzMDm5NkC2ABft+fc+Cwb8n43yi
MeOXT9Sc8i9E0nmyoO51ISYMC5sqvnY+1TzHqytV724pYZDJazLge5IueZdcIFhc
HwmD93ES4WYbHPYBscEsJiqstFwzLNi2AlSG1NrzQvQuMUhUOeNsChB+oFI7MxQh
aXZW0M3aZsCvypoiFpZGjCv58Josb2m4DQr9YSwvfeIXJFmnGy2T9G6Kn1p/pfYs
u9yoIrcqJW4PFwDH4RCSIorp1UbLSHkFdrSDacg0mR/GRVBlBOuB9TrKNns2CLYi
sOjsbbr2UUTEbCdzJaVBanyGaiADAXtIO7jO6nlB3cHdbUq11vFLnSHiAM3T0r96
UDo4e8f9rmjnFCKnumwYdgTxaMwNa7+lzMXKZ0ZoqCBR/48CT3vkYlIyAcaCvHoc
mcAgjTGo6kKN+uBYVCQKYtKz+tbdZ4RxEf3TbzFsssvOO+Ee2nAArsr3jhPwC5tR
ZBbU5Osv8ii/R1g4QHYGUnHS3WTmJA3D6frInipCOrRs9Yr2J9LbEVoD+qbWZfAv
IZ5kgRZeVge9BHLUqzHMVCJpoQsoHc+qpkQL+05zcTsGMuV6hf6dl8vujgQljGDk
BAYbCfXnfheZsXNZ+U2jQl7fZIDLjkSM5Np9MN11Ewi4jvdRiG6DJgWL90rpktOi
sXgq9e/pfYjwTd36/v7vcQTFbUk/aOOMbArh+8HnqSY54G7nHhPxRZKrGK6KVkrY
dPH+hi4r5aemRZJrySjg0JBB6sg9uYqfM5FTEXZ/gX8H0SogaBC0fGrttQDHRCOd
sEqkAP1U3HAP1zn9q+FdTT15JCFl9oMS6jtFZiXFv0duxsGGdxCGm+77NR+VjyNo
j7BFcTnJFYRRFLXEyaNXD7+A0bJhPsTpaiRA1A+Q4FQFvzU2Gx1dWJ6mq7/9V3Qq
BcxgqrucBZ3nx9K4pYw2WfIdeMWVJAttqANJZHhHVSgXUBq+JRwz6jhwQVBv0E+P
QV3fMiFScQjlwHYqLlx1nvpkC3Eche0i94Ynb/hQ6iQSCvt6g9Vb/RIcNPWqwt9i
O5VS4eRza4jP8xZeSP54qLUDPyUz0X1E68Xwz1wqQ+5zif9NGCA1POkKT0Jktrf6
+uFDAWlh9W2DwMrGuZlyYMOi0wGfp6JOrv4qEvRE8hlfTjyDwks85lTVFZSGuiB0
gPjf1zmyYf4BVAhDINj8RbeYm+N9Mx+DnInhP976zI71bVlcdLYKlc9x9HLM2tEp
3d2PHaarwFKkZPEFkbksaJXg1jpYOlUmhUwuNAj71o7gN0bgr8vBLgKvAwRCLcpe
utCgiVK3tGuXFRmQ/uUmN1S6aokVrq/Q2VO7k5U7U0yQKd8dFshqd/6f9QEOYdn5
mb+HGJLdWH7nE7YpPk5AL83DcDQLaQAsr+EwAIHEpNZVF04MgKhrq5brCzC/sme2
hEQrIDt4iV25FmAP16EhCrOlhSKuLF2P4cpuZPIAQ+wRyA1w6nCctQ+CvtnezOgv
nF/W1wDmNoBpZdz0n8/KEEGBfryBsKDP6rsP8yZX05Qg94GkVBi4m9NywEQauxgK
WzBlG8dIzAGqDar1PDHBgK1/SI10QbtYEsk62BCLoqA3icalusWmU4FN6jGKdT1X
vM40eIt0alqb4D2uBYQeBCuAD+EuKHp6CaGqmrX2zmuAXmA4F4rjkuVwpwF3Ghoc
8dtxOVwe8m/PCz+jl1dg9ymTOZgDTvJz6D2Va+ERhjG0LECFUj0mh82m4Tszz9KR
H/duUykBhaKlMeocLWx7tnI+edQYH8cK53vHHJSfOmhhOITlHWqkc4MCrxhnRpVv
VGstG41A7P2PMn4SGiKhUMycoyS7W9ZqMsygughLy91bDn1tgtmlFa5YpngQ7C1s
oVQnwSN2k6xAhonq5IIv1skaPwnKKZZ8C0blDiP0UojPYLvajc0vSpq1RbRFgAoi
PXa4gAHL611T4U5TkTCQ+3aHtiCgd9iLzDaj7Qgfiq6ax/5tD1YapcY7xGKEuind
5Khec7FrtlZWpvzS7mH9YMAF2h9aL7pK5Xexv8PtAtR4I9Au2xTFe9a+KNu1x3HP
wBsstT9KP+yt6kA9JjjYRVGvpZvXesD8/MPzT9Z8U+7oQRb/kMNVt7kCIVS+f9Hw
c+FCIVitnGguga+QCr4jVqiJdipn58lw5i3L9qxNnEpmW/VbYFXD3Bx3rTjo6Dio
VyAO8Qgs8SmNajbSPVMNIq4TSma0RYfS/LN1qnwZ+UzU+m4DPOP5twe+Bh5k6KtZ
2ubBDYSymuBFWDBNqy8l3i6txcot9t4qVHIyM7XDAjoKM1oXIaOI7ChgPtSCXS18
PiL6VoaY2K8uTF+Zrbf6CrYp4ZXsfKUhWGVcGUsmrHUPuXX+RQO3skBmvmTkqpOm
Fk42jaWr2WGSDpYjymBk0Ck7clBRuJrF56xR1O98DiiMaey9ODVuQv9hxjTk5RDp
c12XuAg0XCNVc/XUu45cHzPoOkCZAAck+IgqXvp7W6eh4CT5BecyfeEdO8u8ztsl
HNB3e8HyZa6jqCQa98jDW7qFdofMoAXXC55I2hHVosPlfhX6NEGAYaq4RWU9r219
Ek1J6HOtlLiFkPP6vGimr54ebvOfO1/AsFn3ZddJ55ULoX5LslIPX5feeq45Kl+W
jAaiqZner6EWn6FbMF32ahRkX43d1B4NIwAT/VPJBJ7XXb522MKxCxNZTSuqMo3V
mBv9oLlyIwT/0tZg9FA9/QgPJQxgMxiQ/2zkYc39CbjaLZZEaHm6m0y/CaZNA9I8
Jpkjln5nhlCTPjLYKRJbPd1QtzziN2zFnePFQmfuEZNVY8aajkE2kt/M8VDuezmA
eVgLlzroyo1a6Nc7S9FuURj4qR/3oMLPUWNdz3xcy230+F7xHjoqiv2L+OquSdad
9Nrfsa+bg9YOR95wbJZ5EjdAiuKRx7WqLO2Zod/MDV9tx2GOF788yer9C7PUWmhp
3cwUruBNwMNAdSOeFKEOsCuYGTHGI7lupR9ZyqLBXeVqPUdY2T6lwioiTu8UM4oy
ECX1aHK5Ic4SSA/mFtoc3qo10O943Fp6vy69ogL6ETwKWLW45/JDn5WWQWgDmYql
DRdWIDuosKG79p7pjFCt4a73DzLsc94Jm2mGx6QNXtc25gcrk31pabV8lLCcAOlg
Cihdx9nOkfn9MXpAUSY7JzRbM4n1js06mgRMUHOPTCqzIiVLXJ2NCdTYDtjnZMnR
ZsjKiZ41M2T18O577toySQDP5unvy9wVu8RJ8l9QYX/+ngBmN1s37MBzoOnsFD+W
0JcJwnCKCVqIpDuq0dZG4gh19vXx3zBiNKGr1xBzBwtMaBZrjqhDWwGbYJSU2egN
LIb4XUoABigvu+c3NWUS0we0iSmyieElUOzShztcQSkbiULahZMbfD2/ujIenseW
ACXIYIx5ZF3PjgH2yJ9vop35qWTU0U/eHvsNbknmx/A6qsPXfH1rEZkq80m729EX
EJaBHCSb1FtmJ6xvxmyswvqsZsoPIBsa6XO1do8a5qHMZeq59bDJX/1nLT79hHzd
QcyszyqlfUQATdIvXrGGY/1ITh6T755VdVPfjERmyVVVhyLTnozBZKlccYhxpCwI
SxQaKp5gR49+rTp6tDuusZsS+vMQ9owWnXU77DCx5C+Y0X7vxp0SGhstNVO+d0Pu
/yPPF8o96GqZz7GPX5RgalIQNyauZwsRsDgOvS1INBjpW9LUg0ApIwdQlaymLrpI
xaeVHPCgaKdCIvjfi9NGXGqg7OCdgbAycrrYK7dQnIklDcMOSPKvmTJFGa14YjJc
oqhu9+JaypgDzr4IlrLw6NdSBT5p7e6eG6yoRTKOSdQnMKDDDu4uk+13pgD0v4qE
EZoB5vR9w3YfCM3Ji2DPPwgpVFCusrvyNRkJg7M6lwffIR6DagRcoBSTLJvqqU5O
LBFE6mb/Ao1fWoXPoztI8qHdxlCEbY7HzvMlhp4SeUWToC/b5laJaadoQaT2x7em
/Vztryyqdo6MRzTz0l1q+K7TrcqonyQYNoiVd4qYCY+gYB1N7yoPmA/D9PmjtYPq
Rgg9tub7sSJptW4YBqvbHjXQzfoXDD+4j/imZeMnVi9xoV96rYgPxzW+x35+JwNJ
J23GijXFQIy/PHaJ2Yvkajyn4dh0RGurI3pDbzDnbcEkLzbUmev3GpfK6s6GrNuk
SJyLHgmIrnrVgXoG2phMHm+Y04lv6ZoLeqi+LkPjfOPwz+6sDhu+MUs0KcbauzJ4
B0lRNQxPbE72Q75bZkTynEYUEDIzpNdF5yPk8zdz+2sUiJjclTVROSDPoqzPYC+8
20FputsDGzK0Y8Ba2pjutvzIGsNtoyUa0Er+kJ4cddLFO+o2+AVSsd2S1TBt355T
0L8f11oDxIVGrBQKFNkyOishGSTfsHP3NuMC8ZTdU1teSbTyjxvuQidEkwFO/NOb
mPrZsdOUsLet1c25Ch4CPzE/qjWQM9b3+pFilssAjMBfyCwhhzjdI2k0cS5926mS
TO8CS0RNMdMCXGU/XS69WwQfyVDBmGyUK0ymdwbGAN/jOvEIWxVqBqwki5yQm8bN
E9IPzQJCjYJanzh8hegndFvSjlMOXmzxcPUNFnZn+cm3weWSLR1noIHHLtci6tex
H1zjYojfElCO+8Rpcm2uGCiiPdp+awhhNFTOdXv9/94/tLG8aCC0Arw6ZgXEdXXi
HxJmfBpei78TSmj5nqN4yXvug0PThIpBkw9lQzXq3wuVzme8cF7AvVijNlKpKZX2
8Xu1zo+xSZ3s1lBaPJ0XTIn6yj9aeckHLxYHqTHFzuBwRIfXZVb9gkQYuIlBBugv
kFG7JJxRjYTlmdkZ3tluV8VyE14y4iWg2ie0RphRG92+aeWqWZ0hQ9NHrTLJ6SYp
g8V3/hjvhgJCopC/r/M3IWGMcAvdtDMdW47zbmJ0h72xhvcvFtpkN9rzXi8gIg36
AqDsmDzZ1tcInLIa4Cw9fESiZwrX2b1Xy6YYR/2gtDYV+HZj2/qD0/QOlhh1rJ52
oIegcZvkGbPEiClJXnGcO6DCL7by69B4bc2QuIO7z9jFn7Usd7DejGZHa/5Q8wOz
J1xVdHj/LvCGbqhV4u6CmUhOk7AUdwQkvesyVJizb6x3H8n3NnlwQAUmTJ+sojIb
BiKqIAEYCcRNWVQL+GGa2oWQBnir3Ra3LBhOYPNfQkTOuVaHsKNq4k6nxbJdCLVF
Jiir+aZ8svYbGTfjYoeebeHgRwXlKJe03xGtbKc01UNsDVIxc6LFXO3u+/y1Ky3U
jy8sdQcS/kVdjxaKPjrI/xofj8BEx2ZGMjHXXwghMFM0NdAXGea/sczyrRk0PsEM
b2YOt0gaLe+lTN6KidBSZl/84pvbAgnebP5hzyA8duFjLhHyWoVp9YsILGDs2K7j
awJlImFgD/dFHjY9XpbKxLVDnQQZXtJWGGSRDQhudigEICt9nPUn/F1IoTSIrpur
r7xwmq5op4/dGoLuV6L2UMrb56aZSUZJuIEA7enKr2LgN5SJmBGAHeBPNuJSlYqn
/swzKfBHJEVUIrQkbn1dgvVm19hsZh8YHuvQtCdktWlfxzrZkjpiPzVb+vS3Xh7R
yhqw+PU73df4p4KwPAl4BAHpTkHGBnrB1eqwl0Z56D3G8nhM7mO+oFui2UDAISWY
NsjZ2oMwFLozyQDqzoyWUS0mz5mzXkhiXOqO3S0oIc1t3Egid84elcaKDBBU1eVF
O3om7pRMdeQFFyDfHkjG0LxPWTPAWC0RIWl4PZnZUItUthOoVGuGr9ZxETisT8Di
6DAVCNQLdFa97CcJ13YRlNqKxw7ZnBcsFzh6BvKbwsGd1/Aw2tOCnSMz/6Woq3Ng
/SYXx9RQf9urBAQRYO+LLTRV94nNoHnHeV5TuWgfYlj08nOWcnyuZkCU5Jijsakp
HWnYIR2dg9pImXDJgOxSnqnvf+0qM763/k28kWn0F7ILxV/2qIJ12WMLRnf57Dxw
ZqQr3dATRQLYVAp4asVahrKZjycQz3JdHx7heF0aRnGnar3AFMs1KWYqQVNhfKM7
29gxndUYFv+WXY5YWoIm82x0akbVLOJobuTHAPYoreHZlGb2eWC+uy6o3923iQmu
DZbY+fSTAPqp8mTnbk6bGM2VN+lO1vg495yvUmAauEb5TYg9+ler3LdiCpltOTYY
hT0T4DlBwH6OGO37+9TKxgw4Mqv2j9LolMjIQjvvgJIAKuc0Fg/q21fwW/0wOxVR
7omjK0n2DR2UeyhB3PHYqecCqYzmdWqfPro2ctpKIIsYvSVStD+AW8kHLK1wxkjo
jpB4/S0WLDnvnyNozAsKJMU5mpaMVfUueY8jUUHLukDk5aeXPeyWWuHvIYEzq67n
s22hJuepGzKCbbLns7N68a/tonll6ChU4yTlfBKFLVLlhpRK9Y3Zd9n6O08JNppY
aMuSC4gHxJwxxrsmi98eWbH58s7E8M3brPuDqgUygERw8c5RPRmJTkMvUB6/Y6KD
vP7BJT+4gWZiSs3rL+UKsB9ommx2wW9FpIVdiNB2T46PUz00iaSmMgXF7Keoag1e
BZ2ImyMua+brDPqCW4SERnjqiu8/E70I4aL1lg1hH9tbI2rNE/neWdCQyZJTbNpk
uHe73h/nWT/+LDt8/pyDLjktE5ecYxwLspLVlv8tFi+LzUuoGrtMArD0u851Rmlr
BKjNnvaBsl28hN22Kei1vWcDqrWl4Vrvh4+EikXmzzkfCnZF0fJO9tdkqxaBDkrS
8Q8zyOJ9eu4epqmxUT57eABazqsjGLPw7ZOjto9jWWo/gwd/5XX3IS0E1g6GfyXQ
2g4UwpxM6pG+anCjmdblzh/LW5TD75g9UB1Qw+SIxX8RvQgqO87kbHk4/O8LWdI7
s/HaTHKLWZQ22h4+Ypq3wHnV+Ol7n5uc9wDO2k54oUtnU9vFSGqEljLh9hL9Nnhy
+VxwydVtqSAOPwLiPGJ55rWKllXfKODmsc6ZbGcUamJ58KET/Us6tyv/8rA1Y+ya
IVinm7NnqnVd4Dy4VE8jBuQVvi2bLaJvAzbCOwAec7vjFKJCdfYWhyj3fnAVlmWb
obnDJUyZ9aBPujxfbkWhjfFBqloAFqqLLTzMdSb91lIzO/SinohH0QJhD1PN8aWt
BPpAv/nuYHqAzNTAR8cEuuN1jIeokpwi29qrQDQ2wpXPJ8iFUq46xllz9PBhGRJU
c9IQKatZeKzJIMus75WpuOggA+ZI1bJHQQrlhna9IXls+sbHq96c+jTRiZuCLvrh
4rwzyMqZxS7UZ0nLbVQ4bj0zJUXpA3tEAm2n3Bq9MXj04e6xeaMRlJDMNoj+hGyy
m2lcIB85MybQb+jy2Fb7c0odXMnpV7tTeobztaqoyGstuRz9HH/r99rM0ptpHDvJ
OkO1wKJhTzGTpThhI2Lj3iTPZaVBZw2Xub0Qga5PYWNs4NkxK0/MCyk0n+I6k6cj
z3G7QaM/YdcIrtR+cSVhtwcP67RlQFxR22iKOtFzBOh20qWEOviFeMi/8nOaYyuT
yYF5Yg5J88c7sAPoaUkkC9EUd8wwei/y1fT82hOn7yDKsT6GneDS5xz0e7trgUQq
A3MF1UBt4FHWfxDqPPPT5eKtSmfyHK2lbm7thgOy0NFtR26Ttxb084GTrxY8IwQ1
EzsdhHsUIPHFEZc6AKIN0WoBJIQSDr5F62UKFLTtJhQ03gpmH5wLFj+LNqmPm34B
bAFmM+wNRZAdLOpX84bet3LyOOM9p0PiZdFZ+vY9YkTQiCGE7HUR4HICTLxJa6TJ
RAxCp/CVQlq2KoxBS6eXMvBnIx+tt5SpaA8lGHm4TwWA6zOfPlpKi94UbM0NUxEM
UQUFsQbbT3e5qDtKXZm2fpq0looWQFt8iR6q2cB51JQMpc2ks1mYXQ2+EwiQjw62
CPvG6AAZRxSz3y1Mg6SwdTS5eOBAXNctn1LDQVLWXSWZ53dyrf7vkS7W4W2KSl7g
RnQAOp06M/FFCLmC0V2u/x9aDNl/86yuqaYMj/o4bs27vxE0m3jERNiJd5zKO4RG
6L+3HGozEw93QUOxTW0/JPAAJE1rYGxYPmvAl8+h9PaowZ+Zmj4AkkBMC1xMF9RO
zerB9xvARxpZnTLRMq4XgTaPUj21XFsghZocPnnFQ71903NzfhuBTM44L3V6XPlM
bMlSbG/l8l2sVYU8fh7l5z5E3tCoRyyuNgg5AkDOIPf6+3RAgDMDhER/z7IgJIB2
27RNdU4+jcAQjqV/zlerKUJ+QLMb3J30XkRRDTz+4IiDn2ZTEJCRxDC0zzTf5UPz
DnEo3jEwk5cfNv2NMqih7z7c0tYOTqvUvJ1zZp86nIxCwVHPfNxzrUiaZ8/Dp+Yi
cqan3+n/tr3ARuuIAGoWWPd5kSuF/mIl/02rm/j/g2rIYk3w7dOV4Awtwl33z78X
bABy3s7rUkQz6HNTzUFKbvId3VTU7pIDAT4x4BIgcISqLilWGlyKSKeIgbNDMFml
1ac/clYundNDvuV8g2aG3ORRemPMK1hUNplGvJWTaoi3xIjwWCA0PSfMpU809Ehh
IlQJgaCJfv20B2xJD6VM9AEO6P4qgKtUy/JGs0zHlh9vYN6H9NBF2/ew1ikDSAl5
TByECCsrzRWCWy2d2QYTsbiHSIiJYjxFOex2e+2lQBtYWoxTLnxgiFOOf/zrz22H
LqO1ACVa930yuOn53SW4YxIHeb2itFJDkBHQH2mcLACgehSbDSmiPWrP1aDL9Q2+
aR6pGWZWx/3IQrS1z2CZNJcV0nZfHa+KG9LohNUs8WSJQrtTpymiYPDP52aVnMUp
H36w8x9iXPxNF+HVFQEh83PaqDmG3xp7svvH0UpSBsbHEn/8NKBsK1+YR0EEW6bA
OiQEW2YQrRATqXIxu61gF0VyN5xK/8jPnIxOx5woFDuv0kHXjz81+kM7tBY/To6G
d+rr862v+Ynb0s2QRsEsHHYv7VwWCxTI+nwGMS/uek1hRaV4ZHP+thNKBwAv5KTp
rwIYKlTzWxUKgnMhJBoyij9xGD8PZnUxmAtUrAwGi6tpS/uqL7vUiRRwlqDtgIo2
EydqA53/04AMDUAhcKrCk14EMd77eTxfH7rguSNlOKW2r7rk1hmnlIBi51Yn1bao
lm2oVADRReVA6MNSddcPhMWLqzaYfin3FDu0ayUg/fbkkBAQYU2m7wBvIiijpMX7
UHu8t5jiaeAq8WpAog7L1KQ/tnCOm/KsMpdKIMcK5UmaoyL1nnpC9bxHkB+8/eUW
ZRVY/NEGAJPPBrriHS0hs20pBjefZj1ddshSbwThWywZ16So3D5M5qYjSktofV6l
cIYUxeJgamrdqIfqGINZWDXKRokwujfiCm6V2s3MlDOcCV0cffJX/1LntI+xMsaX
6CvafXluoT/MuwAzFoSaAWn9jZ9spu2789ZKrcRDctgGrfVriDKen4XQaOzHtLLB
mGJuPXnUbbxX/vRWgMBQG+hkCoW4jHkWmQvQ7D3yAnfPOCaJu3gMNA4da2aTKmMu
B6XTA8d/7QTlLoqycYJEWOa+zAdE/UMiAYaVCCYUnS2T6QsvEvYV3ck653CC4JFB
+DdobX1EuWy9JDJIt0a6Po6FXulMYNgm7vNVRphbVyH8xv/snJi12+19yCEU4ey8
6QdXktykOleMzHvmyrTxOtEmmsv5aDcNXqirWNV3asKBnXU3D751QOYX7/uDJ/nN
S1nKvIFSg3BHH+6HJnbhn3mydQOqPolagJRuAVgjoYGUaAJmz+YQghL36NtBUojD
VFXd6ZrdSZFNG4BhGUI55siRYf9VOjNJRxzFOz9JREDSxaoKMp32+JZAxn20S6f0
YGmAJs/5Fzla6CxmGjem8WfyMAF6yg4vkDNTynTyWvpINH04LH+Yy7GK5APoKj8x
zaZD0q55GzbQqgmOw/A8gBsmfVrJPEc4Yfx79STlwdRGRM1n0OB1QKektRLC3OYz
cmg+U71nAVnEc+B3Q1tDFjx0ptXJ6LAQj3ULaYk+hAjw6i5t1jPUrZX6VuLl6Qpz
eh4ZY0DjnHcEnKTWatYRuvENvVwaUZqdXG8WWi5i7i31CkDth1fQ0Cjz0bTTyp43
MJT11W8pIb9D35fYI/fMnKgwm61pBIysVj/BEXULj/Qo0SOhbY/SbXl5q1Gzc4AB
d10ToFWvKxKqw1Zs/LKfju+FFB9X2Mo4sgxPCrq+AL/S4JWPRtmkEgn2QHBwhG3i
vlrcOIsqnJpqbEhdiSSzmSvwsCZK/IHytbXhgbhXzovJDW8xro/HEjNyHJnr+i46
39LY72mVK3wM6SxRlwxuy5Vc8f+82I0f6Du54xXpb+j5Ac2NoSqa0Ofr81A6/Xzj
qNWdgiPnOHWzEe5BfU4rb9SUaZe/J5z5qUDtZdn1H0MTbTTjZ6s5tBZaiDQR4eOt
kTrF73z0E29xvtqM4O5LbGBQLPFiPoq+3ZYT7sboii3SuC84iI89iaOmR1BH+dYI
HtnCtbVCF62kLm5YG0ee5iydpSkAq/DDB6SnNmom4Tgw6Mqw3FFJk40rEIm21cec
5skcgBASES7UB2DBJ8SgraVwklNlZxLNFZpnzXpn2ht8jEQCiT13wdUJdyeyQBA2
hTkZ+yPhWcLzMEGahZ1RyymRwwPEWTK3fno43611GhA5inkuvc3U23CV2cFsCG3B
ONcf3VCBk3BS9SJpGukM4AHB7zaLqAshqZFOcFKbo0cvB3+/mErBe8uxgBoc5/V9
33QYuUbqO4xQJaSn35hcgFpMIRj0gWm99uDK6AOL5WBhlSWMzAZ/eEJE+M6imRTf
yUpx32nsKYmQ/Z60+WeoBnDfzRdvVJD7z+lvVH1dVP7ygFKrYjxeCCQ1d/iFylPE
8PSZva875EQEk7r+4ND4wB2cAozAW6BEpOsur9k7nSLLyFSKGUQ5owPUsKOa2559
Sl0cJUUjsSm8Hyht/rdVyjrDaDJ0Us8DmysKx+sqgC++SPozYmGXN1PMompZM+wN
KCQeyPu5u3Icgw8aryMQr3MHDpqE101N4VhgqwxCTZTvjZKwmJEMGQc9Ts+1q//L
J1ahV4BSe+neIXVaPprNkQawie26wMCAbFB67qO9TxA8caSUnEcIdZCePxHqFvHH
VsxD5rQsGM6mxXvAHo1gQ0izziFy8wtz5bTzxXEWEphtbVcFMMOqFe8P3RjV04kZ
9/yiquRn6ZNt8mjn0HSI04jiGiaTqtK7n3MrzT40kFMCnry65IzBvUEg10olx58G
YrYNzRQgcLRkaQsz8NwWgZI9L3syxZnS0ehVIJ0W3YUhAMApndbcXH3E8JeACPKR
1xosy/GN1KjaSaDDdTIRTfjS6/oPmzwSF8EgQ9tJ+Qlu85blvtkKZYwmqmbpjC1b
0gePtFYkEbgpkub+6xbMYpRjm9Iy7OeLnl3vNRQOe0E8VrIqYkP07uGv3zbaRBud
HcY0U4iU3V4CdtsGSq9XROOJaJ7etmvqte9xI6tD8DKO8n4UFZOGmbisbHeTCd8K
bcC1607qi4q/xpD7XqzoVTwDSFelG8i4rXD015+wbznM2rkOTwGA0t1XnL5DfxRf
H4fkUymtOYR+dzhJaQW4nO3t71N09iYyIRbCN9PVKkE/yYpwQ/KKYAWeXudh2VZU
1vDdxmO9TNfoHuiUYzTQhSHJ2KXr5goCQgz30CIYh1qW7MNf01oUKkftPjTWjWLh
GQJ+dNBsNVzK0WZgwwdvP5Tt8rdX+Jn2a9ApByx2NJj63xanabpgjo/VbP7cZsV7
MQ/qW+4W7x5W8UTfjI7HJ0Q8YXMOynXaNKv/tu9p1XCdvSo88WdiYU/VTGo//ReH
VYXwt54mr7RU8bhDIv/k2VTnPEhJHk7XGc2p2055aW8V6iryXEfYr7QGdSYDK7iB
DIyxK/a3fEIT9bxG9HJlCl9PbEwFef6pBrAAy1gJqN3Vyb7wJbyAHL3BWZp066Gz
6T5Me4XUbaK4ewOxqjNVYC9+ewWPwhLMCUmmH8/5hOcZ9EkCIt5wrnfdkZdMV3Vy
wiZQMUAJRV/R/nmEjIvKuiI/j0eJFNJ8I+wUgLbcmssdKYI3i86nX1vn46/lmLBs
CK3XrFYMaYFp7vnIgJ0yJgvVH/ez/Yr+cCyricx9VgUREFcBgwFkO5+tGZFgb4C1
dpfYpwMopJ8mTCIkpx+jZguqoAP1kunqxI3O7Sf8RV89jKa3529WZXNteqd1MX57
bpLjFldRp1p1kzClgEWKpAbFVCzGMWf77DLMTAjkoQYB4FsPb1sZOC++m9pPFCd9
LB86gBoiLyL0Y04CX6apk23exaOGpk6yIquK3fNd+U5pEv2w97xzQdS7iWpVqc0d
XEiJ+TusmyVzqTcHj71XMXWYEAB3fDE+gu+6eqg/0ZerLRcVyXT18Sa4okvHnCxl
LJbeA5kwqk+VjBIFQ5DJUnTaXxa2ZMIQ+aS695U1eMFXvVT5UrR4+cQ3heOZRXeq
bClxzQbTHI5ORfQNQzmDqMShc8YrEcbeOWkG+X098u+a6We5R6Irh1qSzjP6lVHC
C7+IPcdv4VRGCj2Bh4sWRI4YMnmylwCecvFe3MMweNk0LKR0Lh97mTglTMKS7zDZ
+t423sxTPQm+9DTu3xf9N94oClcPVHjWtDO2y/nf3zePrIroYozM/dtRzkr085DE
Y0PvRVx1pzxBnM4plFMfUjVkmMtP2lUKE6qKk+BkvBsdPsraY4+hwiUTNj5BuFT2
ws6bT3SY3bBYkw7TtgI4/2GwRgQc2yTJYXtfK25NkjSHv9GXIGs9ggkOgZpc5CLP
CgdEOX1wryhjcumJrLXPaZ+HK0V/m/aLZsj6ths2Oe2qsKAc2kjfi+HT+g4E5ri6
jvfrZOUUB3wJ7bz495ohaTMg9e4oIRalVEPQGupQkduld650OArJlKbsZK8lI8nK
fJx0vMofD2dzxRCHRY7LhNQfMfu6TMAYmMHY6pIHDaOimsczYKv+Mxko15JmlINN
r0PIGGInD1tbAokFtCXsxaemoI3dRzsL51SVwoaTzOzynjEfCSK4wNJut3osCdQc
eiPDqhB1kiOqrf8PfwOap1kAdKgxqWMYfpxbAkpdzemR5/bJ/BZ5So0Wfn/tWZcG
Rb06OoH0csbQekQXS9YFZOVwBk3HzfQSHKXGKPKAbKaYa3xZspc11mHgKcGITouQ
p/iBcLgc5jo6WYgcT/iV/p1d+KX5BLLn2dYcSZi1gws7jztvSYXGKND3jWdXipXs
iaSwKFlg7coapopS9hzI/uHLlDBncLF0z190/Ei/Nq0anPjLRzZb1U4BigqLRZ3I
jNaOIyVZlrN0RzSo8Iq4Iik3zMp0UpJJt0XtTo1jT5KuPoFlut32XSPgAnRyjI5C
ZXd+ywRBHKRHsgAeyvs4+gcQHWG8BOV39eRV5dizZwX3YZrnljAE2SmMkOb5zFb6
7MSa15j6B5nlvNnVOpJKMfWP21B3h9gtdGRlQNwMJ7pOgeeqKznrJ+YPqnssAVwx
AvHEFWy7eMkiZVUEkOiVowmyzvf+4HOb2WXTUpj3qOp1zz4ve0a8J3TfeDVXAnea
7uijicFj+S0PU69OLjjJo0OFHnS4OWHOi+whxoh76+sr5Fdyascbb4P2FYb4Je+a
uWML0I5p91XH2bnYyb8/L1YGjKI3sXDe/EGDInypYtUQ21NEnhFTpelHHsUdQ/V6
CmKc0RTccbuQw/ggl8ckKphszTJfu6cm5YtfZt+mW4o2fDGqSS4cewKFn8rKpknX
sU6IQn8XKS3jzvPIwzbcVUNio/eMrj1pjeOCb8gf8wDfb5n/tz0gevfRTQLdg4yW
/vrZ7NKJTwKz0X4Ev8zXgpWuwwUfy0KFgV2maWiMkqfnrXR7whKmRtZO7Y+OcnUq
HrjZDqHm8PaBulPlj2UhEy61+UNe2Zt9k4lU+cB4jYcHqCJLc+/54BpbZ6OzEzko
wyx8nCgmcR6IC4L8oaLCX7xR5DDiRzcStT6oNLOkae5Rfnw9Fd+iDyQ1B219ZR/h
tJRHPRN5XCnYA38NkpC1s7nrXR2DfuxlOEv8kJfsXaSbadFL+jt7+Q7TUXTaWz8L
LSNGykYzR130gW+MtCTl28fC+p4SSdGXty/OR71i4paRPl93OEaCLUkyzFacLJnv
DHQooYjIUuppEBhhJde9kcgjNbdAZ88X3cDKamaXAJ1L3Ac80yhiDiNQK06j15ZC
d6VdgQrjOk3N2pkvTZPrkoRHsutlKsB2Hy8WqNbl1tzw/yHmEUMFXHdINjAWMQX/
ksZpoYm6o4T7Hk1dCegkQQyKo8hU/l+R89H9ha8fc9VMzO9UNbrMEdzlnHIiej2f
cS13jqfHvluWrz3/a/lv1bQ8oX5S+NCUf84lfakgzKRaIml4THW6PDVf/FJn+JL4
mq0GG2cuyHCoNuzMhGBKoJL6D5iuPd2ab+v7HoBbohPWcPNmT9fMoVvJaG5e7fCb
qQEbptfm352iEOuV8/hHaKPOgVjRh1lO7VAY/qTojbPH1e7v4a3MIUgiao2O8BU2
ti4X8pQ+V4x4lnnwfdw16CuYo4Ccx+BK35Oyd2rIlm1zakIlUWmwFi5S3wJE+h+Z
LujBdsY86yEPRT+wtYBoj2V5hs8qY/iljz8t7n2WWTM7HZttV1hSwbBR50ZlRop3
WyTxp/lLT1bhOSupswih0bIT5OhNDqaXGUojOEOR4jeWBFEiC1DLooUkIXoyJg/o
ekhzDTkNXCnxAIhf87cRoCO1NYYcPgTWNv2AXuR6mXXkPn7BRIWncvIV0RulR+1o
p77pKWBg27PvZ6VmanYMLPmX8cIuIQTtAlNQi4WRLSk9suWPPGR3I7FU4zkDM7jE
c6XndNnVCGIZTEzjInSHRXyO4lENfDNbbx1v2Xy+U+UDpakDyrTdpey8oKkKHQtm
3IzS5z6/gGaOi5mUAGhEhpvt+k7GmZiyy7kFp6wy14JBUQq+m6es0VI81i/w+egg
02thxAZNOVm5kz8qb/RbADeTCledVvFI9bB4SfMufCkoGFjuQPKMEwzfy2bGN+oB
9YTeRV/JBI5RetVUK3uSdd74hFlvZS+JfFDkBizLy8YX43fMMRKpCuEQMfXG2NkE
XkMQT9/e6lMWvaXUJup5Zq3b3/6tmtCvwwV7kgCwbxV8k0d+Or15AnleG1cA0RRH
tdgAtggUrBOatpOfTWE+Uh51Pwaq5trWdDE9+0sxRBqnAWiZDNDQP0nQzevJZbOH
8BsZWs1Q2Kt8CmQNIrBsfbXf4uoROugxAwNDQREiUwBE45DTNfA6zmRWhNEY7D+z
y/6u030Qpio/F+EjulU/gIhJbZNZz8GE2F/AboT85Ea7Q1W94PzVJdEejiySz3T5
nR88+sPj6VARNJ1T4/Fx7wXFKhAmDgRXlKwp0Vd1TKZIzbhJ6Gvq1m4y5+3VwNt/
F0kue0gzyFIAw03595ZDJ3CY+8xHRhfifx92gyPnNfyNnJH7bshED0OirCdEgrPa
dMJPu8JVKs0c9bdktva1Tw5AUjrIs44ZBU09xVz6f8lXzDQHVqKqQHfBTEx0yM6V
+v0+hbnfafKE4MVQ9ntWr11wGuoJszum0tAFG4N1MPYGm3xx/kB2bynARx1fYdKJ
k63Yk5oFXWPXblxrJQFfYRn3bC6nezwQSqoyCbmm5vxjK9MF52xvUVoAjwrz5UJ8
2XvXsTxYrAAurKn3nWrVLc8Vbp8fX8B1C3AB7Pj7XveCSeE1I9LsVY/Em3cUJkkO
Xvd9CDXAG2a8fsNQMOt9SHY1YV9ThUS7LRKY61MwchDwwZ2Ea5ssUFkQAMCzZnkG
T6XARHJM3sQ659kw9+x6mW1ytqFyCmsx9IskrJ9zwq/uUZdXhYnrwwX0eDLhEBkZ
txJMv78yjse4LAmwtQQ/tSNWxNSJbOv9+Y1UpCygTAjY2mJzAL6ay61WdKlZByU2
/Gealo4lF6L08pPK91/KghJs5GrFuy2s10cNNgwPfUIOMdC2NmkzE1wjnQXzhs1J
UrA1EIO5UWbomJSatSXGKEqgwWFqQYSnzwczLnJRQY2b99gJse+tC28E9zWWEjZF
48x8vycwifisFsmSyEhmvurO/4+RZLtL+XCfV7Qeq0wifn8RwLtj8ZmDN/1lZs7q
U4wTbudrrowlZPjA+bJBUibFnbm1c4C+n8wm8qA6/0v8zBRvIcOWHLXlg7IFcDWN
esRUiXDr/DZikCKS/l3BZ2OC4k7zpifUnPlPtniPjmccRWBX877IW8pmpBMhNOHs
J1O0ICSUgl+yQh4XKwq8uQsd62S6H2V125WaHgBY/nilBWeL2sDBrRyvn5ilTKtG
vnrLSd29tUjzyUAuDpavXbkBLcOfE6pc1dTOv2CCiG2IKa6+joCM43kwcTlkBOgR
JwvdEKZfOQDXt/h/bL00QMIj5MgEpjnNq+MRrv9xqZfimZk6lr69crH7oAoIGuRA
SrM3ipbT/eUfLUiWJak1bsnTbvlP6fvrrmbFjtmqrCATnMLnHKbpRaSz2PiEqap/
saO7xxNbOWkFcXPjelbHLZfYH2BvHvjXooIGkLzDtsrtmT8PWR2fDHYnRTtXAZfr
TBhKet/5N1X29llm1Xzngt7z3Ud9fR8rgsXz+4RIcba9vp8OaWicGTVNmJWSj6JV
nVcswH+8EzuI6GtbbaVQ22AmxXdvoVYj4pRDaHrGA8Fpm0uncLTSnaZzPrrDyO8P
1SrgAvIiGJQzJDliyN3Zln6k4KYodPkJZKO6LseKROuOGNMPXsOeXVaCbxAF7FxN
wxZpVR/ToOMiXzj6vQJ6NEep9XmtSsYYLpr4OBwqmn0cRqlwBJKRqQM1JuDZlCtL
lOz/mnBH3lL+QhFPBeM9xjjl4mapBAecnBWQ9HKtGJe3PBGtSjy9V2q94yMagOc7
f8fTiZfRtm4RPtYTzMDgH/PUkoe+dbGZjWegktEQwyHcKn3q5PVbhRLHPjrpk0dn
BtPnZUCXwLhi2IIvemA3oTuBwXEwex6HkhnKZkQK2jPc7ODDmRi0/q7rJYasL+1/
h7Db3sHveg25vdq8i91v3tbu86p8lTQHlRTsaEb1Yzh/OcImqFo6lu9p31jblJPl
xWveShM1/fuqGYHbOfdPI+JLqfc7ATeLDU5xY5OireB/yAOAkc/cktrPi8S9LW4I
/eo/jsMSWPmng3GxdNqF3bmK+cjc1myBOtRUUn86PWzgELATB5rEBC4YsclkKBz+
TPVd4rfXJ3659QdTCmyfZ5850497AAZxWgm3ozg/uJazUppUOcNb3f02qwmTtD7B
6HYHewMKzyfaoC/E4h6fY+YduwMsOX2tiSypLrVLiLAQQFJBkqMfGWARwJqnjF3s
CPAlGxkFL2Er0475TLz5sH04GFRSqgvwgicIIBZ1/1JLzsgdcrOC9ZWkMJ1q79mA
jh+c5Ibi0p9mX82eiLrdIjwh92Vg9OPYv3G2CBdD4dEGZEdVDfYUfjZf6j5ao1fo
3saI8D+LNXG8WhGWPYxauyn8qt5S3qovZnoDQmjUCAqVa6HmyjVoKpydTJ6Ck7Mx
2herFwx/n2pNH1MB6ykTzvDtzKkD2Gn5WOiCwlm0kVD7XXxVGqgBrupT137e7i08
qoPcXcsVKjrWwyOhYUVEcfA0+p3TUq0Vv38LPauvIQq2LR17eYvTe7EMxpsKvp9l
6VzFhKDE6NeVv9muBaOnp4or/KgQPla83M29TflnQVtRPsABO0sLOtV6n2xWrt59
ApufRHVDOcRrptUXMM0aBYMUrRwuqZHfyvr0qruyvFRZOaplzNMrd8vkZlU7MsZi
hoJLWrG2yP6mcIYBzoETCNs8M/QvLlbSiSpheUMlkP1ItI4t77yQkWL0eqfrCkgT
X/xzDezcqPVrHt51ipqMWIeA1pma5X74kN+W0lQS3OSpKP4rMuQCnF3WpMuM9Ey0
k82z7jYqw5YCe76FhdS7fC73Y8d4pcLzU0Gkc251P5joJa9XZD7fluBkL4JqMP5m
eegtrqfgsxj1PJWPF6Kyw70ReOjq96sv+LgObArGxL/tFB7hM9DYaWHeMt8Jb2ob
twfO7LEoRt+cMqpXj4ltTWN6vI9Newd4UKZcUvC9yg+VDF2P88fF1V/aq/T4UTU4
G3NrE+TCoxU1c2HbmMmXFmYCDFx3n0kaDI5PxcHEDun0MR46pWYhzQ+H4wBCUiDz
6myi14bVkO2QpwzSaI4f5Eonh9o+VWEDa6D8npeITWoah0LIGjNx/we4xBPB+kqp
veRyp7MHtIwZTp8X9EFKg5XXh8NU+oE8uxkUK3WCoErRs1wyS+wBvtygKjkR4pQP
B7UORXuDEUgWen3HgXF0ss8L3jQmADgKH9jsQ/6njX7SSCNH1a4t07ZoFO/tyn0T
La/h+QJixh+VkOqQgRRomdbq0gJP2LR/LHKzY4ref84YWkbFxZuBKohsnhctvI/X
QfKjitGuChvYHWSycIsi5UFQ8nAQFMTeQvTsUxHLhsYKEB7LgAf0IJwgheffHbQC
PzZEOT7MyRUA8oPHuKOnaPe2rUieOt11Euuhn5o0QMU3IqzVWBzgYF7gxh9znf0D
PFktfrx4a73BFyfD273KM+MzKd+Eb7AwV9rPPzzf4qOLmu1F5Os1R93Z0N8zPRAR
tbq4blsLWgv0zcZlg9cC16RI+u7tRZ1lusa/PYxoiMoJLOxfY/7RRm9e5ZNQ+vUz
uBjNUkShwV8sSI3DRQRW1I7+HwsJWlMHAgVvzHCukpx3JelC0GD6cSWZlw1+lii3
FEvwg/8O2IPpXTjgKWdbJI1pjA3Nen4jMlExHw5ZURWN4saC/lP4RvlhsgoZO7U7
qQVxWyvA8byC/3xmUxTVw3xIctDC4pjX/0gY4tAq7pw+KaovpUumwHPWIZI9v0Bk
sH1QYQ3cU3lC3Elh2RZ+8FpZ3xfuhlnCBFxi9KRIh/86rfSyfzvPggOYRr2adTeU
2TzdwpkMH/b2WyzSvrJgevyn+u9pKLrkBUXQRNo1b1jT1+LQfh5vwR+SgXuzCtqr
7P5LY90DsEwTbociTSca2TnVk7MSCSZhnFS5Kn8ev1wnD3QY8r+yvDstWG2/eTIe
oBYPWCzGVYbGxjJeB+yknqhUFepAPKo8Or9CbQV/rk5Zmsj8xIGgELMAGFxDSRBA
D851dTv4OJieEL7xSi+Ph/dZzZ9GuUHfAgxOzLAxtL9i170K1qVWhhmPX8hfwH4P
Hmlq0swiDYjQNOnyhh4KHEv6/Bq19IvDETq/wlSGcF7dNMHrvICTzwCa15R4HQTm
+YetpiNM7RHhYeJK+P2zxd9wPFCMx3Myjm7BARSjeaMAFGaH1WsqPXVOzMjKwDEq
briBCOFVH4pX3h4pfBm9PFvw/QV0DbAPFA1+eaauaUyW4eQmkYSzYyMmgQqK1+4G
7XUfeQuNqlSAVUjo/p/aUsYryQOq2EXyHj1Y1aWJFOM/dbjLbHrRQ3j0SvYxuVB0
QzfYvzqt+jtLvVzoqg6YwCU8mV8p7reVbD7DMyfpYU60btyOGXPBuRJDvLDdLY/C
JPAKfKrAb3AN0t/iLLuJEPBH9XCq+HXMNUvqsr7CRgitxknMKAfx/zgfXpSG8oG8
F+4rcKuKcQle48RendPTtJ5GMBfse64BBvAKxOJhP1j2WSNP1rE1e5PmkL/+X/PM
sx19734uy52dwMy27lsKBXdbXdWC+ZmkrVkrLiW7J3MkvOyD1p8JfeLPCfHAjKJS
op7xUpF56j98J1D82sbd+aJK28ZrC2OIu/dgBxjjGdCYgT34lndwGm1O0WxDUrNi
dxLo9Zb7Nw6T9mxjDHgvD7zjxHTmGe4ZWK5/HiFY+B6AEWBExPCPnm36Ab6am1df
XPIJdS5jgNZFpPHP3Bufx2Rp9+uKrgM925L6tcFFe44kVxd7RVSVzkCgZ4YwF/t6
zK7kKMHt7ZD+dVI7GxT67AFHD3+TByW9Kz0DgQZh2cj9+kQtnfy6tFRKtEtR4SYJ
eY7dI1yNJaB83RDMyLfRyVHfPBcJC0BTqFY7med1M0ZBTfbedZ0J9QGj6Cx17Qw4
osv7sapO7A1EbJNVMtIcg41WX8yKVH4UQYarJleHj9v6hrMFRO8ZyND6WFPtjbeY
n1gtLmEg7FEVk5595mk8F8UpGCmG+GjjoyIBoiTzgIWOArlQWXloakpeWJWjSzor
ho6/pzWnU40qk0FnAIAyIGMG4sQDImIZRGIpK6lHE6+G8uv+TJynrH2cxRTvkNby
0TYDKRyKqnC6AjlAACH7ptIExG1Dk76Qa7DwFLg6tvfMZQlrhZucfHCC9bOIHI+9
rFWj2pfBiLDJVDK6l6JeecUAj4QMBHd/YnHLNDp289KMTY/d+3KYxo04/g/jxVPG
JG97VJhS7QzYxyT0OjaPoLtgCC1x51IF16hIrDMKztkfcFpIou/LrFhgptQ3krfd
IRXfzAHu8GOcN92IK+hyot8Lc4DKjAkzOFv31Y+7cPkcLwup56B0iFsJojSg4EUy
G2C0g8dEgVCvB0zuNeF+AS3mGG+5EBN3aHm6yukD8OniZ++9RIybN8MvwRyEGCEV
yOwy3BDnz/sJeXEY1K8rC2xCm6F0Cg0lMw1oQsT+6ZupDSjxka6iUxOxzf0iTKvs
JwlLWMnp6SVRo9cQPntZVnkbiXxiK++vDPuK7wKkyqc/f0CH6MFdASLQ+7W6Wmro
FcjpRrTOQkonatQI+kCPmJsu/FnBF9f39/2lmpZpxbxI8IkVLX8fIgVJgzG+bq9Q
XWu47nqIMSzL5OC7szLQhXMM+pXeISwGSv6ndEioOZyOz6updmc5+KRGykHSAta9
aYbkcTKTAlLn2lcg5KZKsVW/z6f9FBknbnAdT22lB1I9dhxkWk8aQWkMxp1p5zYx
/OGHelF+ZmyoXzmm8+2zE9YrFUX2dNlML1o6J5iR/yypFTHBhV8WtwVxrKOftwrd
StPXN09QOP5qO8huTnlBTfykfvWLzq3aJXBpoLXteRMfZoIozvbWCpGT2Vucr8dX
0qFx+Sf8xJmGrcMik2q8nRMC7E/CCfU3+WjdHb5SckFTCTAriTqdJxQ5uzNqyKVg
PuA+H+9rdm7a5esG+41D2X/F6FZHWoIHkDv03gGwoglpieSGhiRD+VD5szhcL1GT
8fAo9F10ZWEWbh7VHXFM75Sy+uu/QFpUknLmvXBQTZqLiGiGEQIjmS+5/MzaaaV8
KWPYJaioq45g0Divbm7PcwHZnqnv2lZHcnTEc3HQcC5X7Oec7TKMCKo+Rkt9Z9dv
tQj9LoAcQMJrhpIWGGFnqY9k3I1U0G+0JU4PYQlsKewan5Plg5A/6phTgN7rx6Xr
ZEr5fpB4a58Ff6a1uZ4pY5NsFWyMiqyYvRlQZEGklVTdwqRKnu6/kT6LuTBZpVvn
ORiMrdiHHYrvQFkrURYYkdfzQlrgVFYf0bsgzQ+0wdOfT1HySIYgIsHPhwFw+6AG
g1UVdHLpxTlIl4A5uqMBu3aLnbj3loxQbXENvqFx2cdcsOi8jeYS/+l88jRnhqhN
vj+GhIj78EOJBCX/ORhsZdK+g67URJKhFWBesycrSF4uJ/6l1jO4EhFQ5xrRB/wx
qwvB0jwDUGHGTQ5zQDWluayQYb8nAnZmdTn4OMnkgRKk2qO0UT1dNUoXG6F1tI8P
x1RDtKhorMo4OUma3Ys01lBW/t+zRg3qShdGZU3Kpg+HrcUW6nT74oGBpJznIFrF
LypsxuKx61UHlUvhJvzm9bFBlQj4IYblhMX0wgMh9/CKb4eszQxY3lmeMFLXDWTY
/aEcBkje+ktiLDeIRDnPd22xmv5kIMOuoripaX5x7tqA4HVJt4wNCCzomQ0esv69
3tOUZC7iR1x8CF2hWUXXZgaxkVQ9lWEwhE0KjRVoM5e7Xu3jBFTLySEXzPqPQVd7
N1rk6vMYhZBEIz+45AXui6WMqXTHkuK8xRDHItRBkwis1179YZes4iKtJG8V8H5a
pPH2Bd+JXcK7oUgEbjXLbO6D64cp7OX8jggbegQ9nGaeZmoRAhmMTzyubRRL/5i7
AW9yJI3CA4Ome/mWPzvOLiVmyKebjy0WT1JbawVbL3DloN6cWMSloIsovndgUsIP
S7OIEwz1tabP9RbeFzzMV97K3YBUUWfjdU+g+oKWe5XKw3gf7rsmiRnUoLshkQUk
3hPqWYo7Q8DDrQBMl9B6uXH7ZRjisEef6nJp830uCVVHL+afQlO96NDPLWdFs5u9
o/YnFOhH6izBMbvaANxxQuQ3LQ9c1SnTZe/DOWYzAa43qMJTDgRZLaM87XGDCfBi
ftutLnQrOMCgIdNeXXDKjRFgZAl+CjaIrVMGEw25QcqwZIVdv1d9c6rrnuG+x+Tj
5g5UofVs+D5nKRf2C4yHGhYv5zc4IDFTTWsECpJJRnvN3e2wYjlwT8yruE85PGDm
QOGobjkrfCWtPi3dw66lwhpwy90sc7m/l0X32JThWtB0TnQVBEoxcMTfSBXjNstW
sl6WuyA5iZYyi0T7f2jtIFtfXfeodCTIhw+8UYwmUtGwSSLyxMk/P6z2DPaGDBcZ
XMIdYzsOLzKUmEKNrcsNsdEB4NrcPqs2aKUYGyNaeaiK8JOg7E+lHLzKSUPIOxId
C0bdAku7jLFtzDLutX8gaoQWZvNd/rrCISM376sgpgkKSlDf/8h9o7L4rEyArDQz
fz+AIYxvQK1m4oRGNK+5NfEz7PgXFJGeCm6OwCneNtEkgJA6LdbNSzA8cHjjz7Cb
7HO74Ky7RDbgeJT0uUujMjlB2rWy2NIgurYHmi5sp5ggMM239f4HC5iuB4ND6Kh3
4cC2UBxLFgFJVn47sryAhDfKjJypH25IFzNdqGjqyQEacLHZY4N7/Z/q3FFI8aK2
iezN74GlrUrJzOfpM67YC6vrRLJrBdi3W2rC8l/mnJ8rTjN0qdMvzhlaaWTE6qRU
CyNZJUk23+zfkHvcKE8EvW22AE7gHQaWzNcOkc15WBT+MA2Vkhgge2zwd+IBVVsZ
wSwPnJivUpl2rR9EQoEeA7hDg/xwH4CfdcSrxenouOvq8Gutke4Vxj/dHVJAg/Oq
/cA+IsfeQaiUP4SLQR38OIsK3pAX2zpmQlicLFGKsZhCS61/xrWf4rf61zdKbkyq
LUZLFhX1tm2rbVmuefZJiKl4C8qK6/uR/chjStxWtZCGGc4un8kNLqBzaM1M24hW
05GaBCOD1+Xg6oGFQPrCZsRW+tTBUyMgaEFwsGp5mv1I5g68nrjRWv/UfQsEtOf7
+uZKDYQYDUuL3C9GnAxbgEgdp1AJ58OLSBdnO8fAcN+pa0VP4Yuy3dfK6PK+rc8k
6kAfA59GvTB3+mbefbbUef5Z5PiRNSrAiGishaiyWwDc9oVSo7TJaMHLZLl/QMbb
C5c6M/FyTrFvMdyLyp6optOXhb1gE4vqhyImaXhH53/tKhEQ1cOGteLuKiiySvSM
YkAFKjxV1mXXGF06hZXoTo6ogf6Asy2jya81Ej1hnguxyF+re+6pf3kw+iaZrDsc
mJIBqkng8Mjq9UXnlliKuHjRJgO18tGs/pTHr1KYTzm/YrysN8aAzV3Hw6cbiFRF
1prnlXcltbwhTGb1L3wC0+bkQ7ftTLKDeMeF1G9lQkNFMyhMvPpcDeP69JXNLW4P
ITi5hqHf+uwTpVHy5qFER+KsgaLOw5+TD7pEGmcGFtDxpxDfRIN/sQR8KA3gr9eP
Ai7XbRv8z2ihLBwrKB8yKH234yrlQhLj1Z5n9IsVUAtsxwSWCiV7VWhlYsNNLvaj
vHODJk8Bi2cnUhQLuNly3sACakloN5tnB8GzMY35iowMDo7CFYhrtzZmMRSo56TA
cPQvNGjGJ4u/wU+lTjPc106hTJeT2PuHU+T4VfEBPaYEx0r7Jhpwqpl+wEOQyDQv
p40TSwl+TvzR/7KOd5sYLKL2AHyFNLqAEOkO6U+02Z2xPpnnC5qx7hZMdHLEgxyH
3f+93mFgjJYF7TRvaVtslyrAxKMaVXngMbJ8KjVL3lIMvd6PT2Y7ooMZeog8GbWb
VsAoBzjGrlgtx/Yz9nLoWwaRYZboujt9TaN/TPd2JVlFGZDKWYR8YX5NUTQyXFtK
FM/ie8Z+Ivs3lW/kjgVA/Uj/L6lIXHuJ1cM7a4GLlL+vLAj1TJT//txDX9ou5kxU
HEHNQxyCRmLFhLoOHke04ng6STeuRQJx2+gEtQU6HHaviN8mNgQ92cIjYcZ1YPhO
zXtyJHh9skfbPgBBCStvp/NTb/VC0k315UTWQMOr0/jn9YZH2qHu5J9sxNym3hBm
ivoCi9TMOFUjwwPm9NgNRYJhgBBIwPGEBhqmCBbZF1faz1I7QvIKzIPgooOPk4qR
WNtvK+J7l2DGHn4XOuEA8ucMMy1IRY/M7wbTspA6v5415DsoKDoVIZ4P+FJawmve
padH+dZ3l+TpBJc3H0yJB48xnDDaA9bjOk3Rms8ZLFSSlrXZNMSoW11bgZLJFubx
Oc5moM0qstvIfZgDdvgNXY3NWGZsu2Xg9zxmuf/DBDkShF8xB7J06VOdGACbP0ri
ahNOCetd4cZdvNQDBg/lKAozdEJpAwuA04R/hHnvonbj9ol+h3APpOahVuLh3sNs
Ev/mHq1ZsTs8XA3orwCmoZKmxECnltbfebRJDCn1J96Tkw22nlWtKmc7D1ygPPOo
yprkdq3cVksyU/6Otq6V8bcjwC0U9086V+GXIJpbXBSYy+ZrEfr8KqUkkbAOXVsL
Cmm9BaetyBAEkmYcMNULUEJ3QydQ072yFLjS1xRHELZz7wYQH2ziY5uaXX0k50kI
0uKeBUEnebfZb8sEegyPG3oE69+7rpCAOSg11yBA0kUrhypqqLS4w4bqj0I1iJKP
lOkl9W5meE60IdlTLtFc1guHg+jk3FYI7hb8sM1hw70FokS00Ta/FCh0VdQ5yN/s
yH+VsFJtF5JXnERIl5MGGbxUjZ7FSe/hrswWpTcRBDwzHpLDgLlziTx2/v2RCReY
aObqiGuxl8YUcyT/aelcWaMM1NHND70VrRHBSg3W6WFzMnzfRo+3XipC3DU6RSx2
diMVR2Ebj/7rUMVAkljKMe8TDXYncwwoGsGXI/UbLSFfIglkhUCN8maQIwLnOXDz
W6ze/YayZffhP4sPTMEEs0hbNlZKeqZj/8Pe6GFfbtGXOveJ5odUUo5nicOv2WEs
D7wV3/aylC5YBBygKuYJqMaxVUbtbA7QuS3qdXJYDQ6+S0FxoBsCrhmwevMKsDU4
S0u9bLJ65WwyF6u4aFbt2aabaRTkrC0mqaC0JEt8LUoPaCSV+Rruo8VEPrM/2Ui0
GVtZd7Jkg9oiJHyrOEDVDPQ7+xsKrSb5CqWScaXpEqceKpKTY8Dn6GNAkc6BkP47
dLhKDZfmFaPdWd4KKOFL37LU3z9ORazMYpGpyjVAjSFLZQ+DjiKj8bl2L4qJsOYc
YjeXOFKIPu/FicZte59CO2B6gqbA++Ng641Wovl7hGNT9alNi7URjuww08w79ZCE
ndPwxjbeJuH2uQ58h9Y1UB5KLLbkn1A9AuYxgWLYOukbBJ5NaS6tB1vh5igslzrA
ddRn4B1aeZoSLdtbGvHHCYWoGvcq6dKEuFGt2xyEQ7RddG5z+lmMD6fPqOFa3sKj
T1ZO19eQM9YD0xr/YT7BCLsQx3OVCkoziXO3z0Z5/C5rzCWFzYEMp6j2swTVVbGt
wUNTcOCe52Xkw9YF95AoICZgDX8h3Y1XbvzHURMIbb61PaU59KR+uYAPQvbOTYw/
mcNdTnRkaPknLK5wLX9QdmZfiRuzaOMJFFu3+2dne22jaj7xXeVEvlHS+CMtXNOg
Jzhrl/0zWw9H/abQe+aJO9cc6WQVHtL8nMmSh/3OXiw8JWkVC2QVE6lk5kBMlMsr
2bmTUXn7u2YhG6n5GXhRoMtTiGQB5ryuGPIAuu+i8/UtUTWOg5AjFvl7imnOeHDH
SSox5CffsERmdR78ZpVSH9dGQ3WgxLxqyZymhvbxHvdU90qWTuyoI5Fctty7I8hO
Beuk18M620/ydYzzHpLQfmATD+DHLluDm7gZyTjT4LV1gNpF335z76N7GKdlOj9S
aAxUNCbN0qoTYWDGFZ1oLAsNnqpWgVNpnAwfGunVvZwjzivxLj0H6VRj3HE+p3hJ
PDCvkGJdrgYI/5WxAEhWiXy41Rg8eHfTbNqN1KdiP6q7zyo377xgNJPkMB/zkuHC
zGKLUxJUrEGOnejB89OH2lS9wWnXQx6MhsD4sHa9OXpEkLs2GmLMoB6Op/fHOOgS
xinrshW+I7aN+cQcmbdZzvjkpaj6/B4N6ZLXw7Fyim+JFh9y4MtGlwfG4vMJXlNe
yfahtN4VUkHBY6wZj6CNZgIvsVxA8boBn3tWFGEIaxP7l8pk2sRl392Zndk9Uwtl
XsewKwhABW+Zg2GYOX6dhVtloB3WybJsU5YEg3iBHP5xDlLFF21hiVryMbrU6E+q
IxShyVFnLyJCf1yb09uBfqUsicOQfLGaFCxR76AH9oTLQjVdPA8YWBrla2TftHV1
GFGxM2vtmjZUO0J4W9wz3pByu9rK6Hp6CXQn6IIUWvvvKAPpkAuFnbvtMgRUoXjg
ryino58Yhuwm+990TBU3pxv1MNXKiEx4zLyf0t7pwCHu9URA+qgLN3oREHc2DhK1
Wb4YT13EKsuAx4LWQokeKycPiWL/z3tQxR95fKzBEEO+r420emM5cBRGXzbNKbyw
XKlTZBu5FVEBCiCUN5wmhD08vEIbTdaDtYlwJ0IDA1UP/xJTVZwEf+DfNsQbyR5k
o7qnlqq8eqJbQPYT2jt6QCiGeJ0TuYYWC6IR1A57kyyaWPjTYMJCPrvpmsS4tn8+
aeSPjokFPJNTUu1H5zMeGsgEzIrTl5P1x/O8eFqvmmeULCfv3LJe5FJNXvc6FwWT
R/y7/OhyAb47GC2XpdZnzoYaUgygH0CJvxusSpaYlD9cUPhGwaM4vUjXNLhrARXL
GyYmMqtXkZrfyKJD41pEVUgq2jerdioGs+gaMTYO8ixNTuq++9dqdMKNpR9In/Es
G17fWDWM1RpieJchqL/jgP6lBdMQUEg/FTnjA2gClWkCZvrDRBLxDGr0eCBSDQPD
OnD183XgT0qUl95ST9haDLwjeHSjKuPD6AfAYYyMfT4p7UeE1q4z4K8P87TSaQzJ
qcGv23CuZufVw3nOoMJEhvCs9nlqb0PmXVCS/gY3JWuvQ81C3ON9Pqid+Vw1dTrc
+afOlABwa0p6JpivfEDIn3Qvoz1qB8wHfjhvoFHcrU42gq2oKdmF+wbM8XyF8oYq
b4XQp1mD+ap++S5UT1NMFuwhWAEy7RQNqlXHs191c8z1qxdrpQJK+9I7KEPOLhy/
utRvT6iEShDeXbHTNhfqJvi5l79o8vFmeQroaPs/eQHZbo4WaywyIIthi94cA6Ia
q0Ku5HKdvt8RJySqnF715ALReFZB/2DIcs9RY2tfNL04yRoIgAQQg3jqPi5/Q7vc
eTS/1nuU96ySgkF/J1IQxWuY5twsOOnj406xpoFkFxdwL8V6P2HzOkRKxtIJjPXB
Eb6Q4KsWGFVRpUaQ4br0oOAZHpcJjD4VTD/wHrMQST5IY/+9QAKCKtrtFQdIbbTn
5zCZqqKVUvZ29Gt9c0iqdYpm9MXBTY7xbziCSlEH14NLlm+QznZBrXPUaA65nCVt
KNmDphwDmQCHHfKuDvVLnNYg84JtZcSG1CCUHdXBElX4Fkmex7EKwgPx3ZoWZ/a5
NNt7xG9j50A8fUO9kI4QAoAdd/+w/28jM5Dn1PfQSdtLrUHfRrQCoMyLrv6nH6OO
EZAsU9WRMpoOkpOIGapvEJKGdmWKj0Ln5nQ9QlGfzFKUC6IifrXvuI/PEyueqjRn
osp9IIUG63v4IaDRAmMJarNKilMhhzH68486EFA+Kq8Isp7CL8SnDD13enKj2VRr
5iOdLUtQFRVJFMrTkzIzi9yyA+BnHdvZZ1yeDPSOOzTCie8G3Mv27tx6WVY9zTc+
wCbFVsF0tYiEn1BaTJTncBB3+w4nIXGVQBuqFuceBaTtLpxkSX49aThhrioo+IoG
qsF+Wu6JZkUJPDWdoFNF9XkrGXBy3n/ysGI/dQPUMMNMKT+4SYvFrsH914ctbOWb
EIutZMUHXoodb+Ir8sf/EhR2BjMYKHk0lpmEREGiWoosSfYhQammfeBNHu7pWHJU
S6XO0RxV+IO0PnGnKm6LH9o4HrH8hs9vx4SdCaqQtZRPY7eTek3lbUwm2DPvsS19
hkYH9K4ChFp/taJeJHMm0btDJ5lrrr5tugu3q5u1TQZ9b84P5Ym6Fg8j15aMWA70
Ai2UTgPKg5EEBKw30sSH2fQ4SYS1TTLk6Eoid7r28n6NLPW4LxjXXVgfx++I3+S3
pYS/p7vBXOhKUK2jT166eg5VlJOz+zdt8/MwtUWy1wiR1Xmm8iLJhyssnuCHW4TS
NxNXQLKgS/OcNnZ2IiK6C0Bus7K7YVZ7AYE7GF8/xp4sJd3yLGl9tWFXNunvi9RA
Evol2SuNC835O3akBi/WsgnouJ26cH2WJ8spxobBWWABK88ypAG881bvN+y2Xp6H
nTFXQSffWo/uhHXjVLj+Cbb1yY95u6ZWJzzH+5ijuKoGCD5G2fjWzWGPWuZNiJfR
QwDFMqleSAucVU89EmDWtGcf7E/xBagLKA2TFM/dZ4bmS8NedvNNbn4J3rjhO2fT
7JYPQEdHVYS+N29PA+Ap7bYMTSJYNEcT7yrPPYZPvokv2bl8ioPj2xV3GVfk7X0U
LE897u2hD22PBTsG5hvsrrU/98btYAVbXk/4MP6W9TwyEH1gY4kvzGenznj2LJvY
GGsyLBi/DlXYKVwEobTFfTT2mq5zxxpLRfW7k1I6ZuRXdxmyuF0Z/RU5PSuRCwJ9
mVGrNR6yRFcZoKw64IkH0wpUgSWuRLQI7ufDZbqOwp1a1G5AYgkKVDsEGIT8zlAn
gxe9dHitZc2jURRKrgLYaJiRrjiiRaNhQkXGQ6yhrEo/DdnEqJulcI+Pyee9c3nf
osvsTGQHoADfu8ZiG76cK8lBV8hBUTPxwjeZzx9jPIN38uqgenhfs2dpHDppyEPz
gMpNHq6/KFUbiA3hDHKgXYEZi4s4bqn7HD/MQV7dcx+oQmzsN9lPm/0/ojJpS4XD
CUWZvLVKM9MiKjExFOeoq+1jpG7SaKRNKtIE4eLVM2dgh0LRG+O/VqC482JJoGuU
0AxqreyczHO7S+yes2b/lvuarKM1w7IZzb+TBU/TvaHEh0/+v4ZpqulrENJBd8Dm
WWS3IK2rYfndUL0KVsOchJugnAgqD2v29LrIEOQnMPYMC5FqtSujUG179p8qhYKJ
53TYt9NxJREUJhU8b8Za+uPBS8CuQl+5iaz+sj3+8KO273tcfU5aRIvKkEIsvK04
Dsc4ZeUVI3cd8TQuTdXHlvgt9seBuxrJ624Az2qCx9CmvH8RiO3WYSpjD//6MvaB
QvcoIFNaxkulDcXKjcjLuvmc2LeX+PtEY48WQtAfFsjZqsuvaTHEvzDxblwpSofp
ONTsasQMAiGsiMEzKCv6+4N945QyT2Omvee+iBVxOlql1k1bhyRykIRfYPh0SxF/
8ROhVSsWrq/CCNvxltYOn7Bc6GjAExhuD/53yZmP+tqZC/zTJTiYES3PNe3tYev+
WPDHC3R6idbjoqnjLxFr/ESDh5BI2yR4TUBKqJAEzkaZvSGp7xRbiLAlsDPB/FjO
F2FFcfeNT9/8EfweUCw2u9mjG/EPYTHqbrRukM2CQGrCRmTPdg3iBqKzUdxC291g
N+xsuKnne7mju5+WHGp1A9/WIK31dCqotptP8bv/l3CCbGRTiZC/6Dk5D72A7PuF
K8DHgH//bFBrowqQQ9bV+BWsJsd3s6WhfPJaLGGcsCZGPScAGM3su5/BM6YLqS1J
Gh1FfJ76+rpxpD/rdTsR+gKbEotNgU6i+evQgkcsnvN0UVtpZiBMTPaLQUkhxEoo
q18BbHgVoQ2VqFFkL83YmP5v09UxbxN519WYVvTHK4Zth7Sma4mEOQRRxljUu8X1
dwXTyUM6GR6G+/9KCDapR0+yRbZULuPFI+b+FUPyc1fPK/iIX8VWmKp/phwo31os
4+2vJ6hcM245YixCOspHRjkGB7MetixxfQmKSeUBeLrMr2kN3v3VGULTJNJZc15T
ue9xkoWk0gea1FsoNrCdd1EYrvC+olcXgr6BHE6tTa0ZcjPmqwSbJAycwMtFzrK1
5JPlyblCEHiiDx91gbCeHuVbdvCbMImBkG1DusrUiowMighu+zszy7QmFIlX3rua
XwGllXWJ9I8AGj+OWZ46gzdGnaKtw0iia4rYVq46Ld5Ln1evBQwW34pg1ox/5Geq
bWYxmvhm9810wvgTZ+o73+7FW1Zp09er2Z8UT9pa3u8J4L6idpv1X03uS98Krk7r
WfMOqw1HE70IAemBUbwPp/V6OWs2hC8TKICEAboeQH7npkOTnYDJ+oPehJXDdUJk
hG+Z5wjNSaRqOqE87d1PAOiiTP6wntYZCA02UjWqZfol8EJkutuOmj8kfiBUOosU
hLXK7qC3BPJb6kdgvKjNjn5Hnj3BFAdqSjz0Er/haB5eMPT9lPpJ6mlucHqiRNSD
Kenjb7lCpuPB0OykyyOhEnkATgDYcaDLDOmtJnVMIjt2evHnugJAGIbRkNmnKZjS
7ItVzOdRN6AG6u+98rfkm27u430P+pwbMKByyCkxclDY1VTrAz3qQxuA3M2hAqxk
2c9rza4/rZC0QMpzUVAuDxABHa0NTgOZKYQq9O2wDMrckJqYTQqoqKxWwZn9fo1R
xjLLN3Z7pPQmgIwAUjGVFKnyvrFfldnhiT+6K5lXJsU1vBLXiXs7x8GRIMLP8mIG
Tp9aHR6DRODEmafgmQ7iTzRTDMk77jlSFxhx1LYSFy2j6O4eBXO060DnqA67dPL8
DUTHHwClNOjG9jPO+n5HdRM44P1e5MQtKF48JxuRyOlBoUbcDMJC/tQyw8i/sy7L
pXKnDXeSKnFMXaSDhzbapGSF6qFKWV1PpCRy2VR+RSxfWVoIxGF6vM6r0IyEcdZ0
CxmUxBtaqoOI0iTqFzLgNhgVGobhnEHAnkEPKHoCJjgnR8ZLUbP1Lx/zyCHy5y0F
3XU6kA0UevlVYwqgIRiboGWSN7ihztne9/gw5BMhcSfpIZFowwnWcJLRemmxUMAn
wb33Gisgg8RGdjovin8sjS47hWtHrr86Nf/RXkFkQ86Oo5Hu3fN+GHN+mIyAXOPy
FP2DrrgV5F/aAyrsG9ZaMYWDfDdCXpYPd0x2OVCJhFncGnkFUJySQzYWX4r6RoZy
Vi+AMHn3/oEOwQ1Tt1+ZvmnVwhltR0tYijceno7thyzdXXUb4p24rkRCcvgicveO
kJ9meaAVcktY7JCR/t+MJqRd3rFTfFMvz06otQsM+ERzqTnLgKRroXperkNFz6AL
eyM4FQ4rKoVK/W2fqocTgvyJqYhgEIxYo1ZUrlDmIqQCjBn6LLM8WHvvpnkwZJP9
9KbFalQW5CPCLpa583vXeiT+WO37wqcx1jOgGzRZ6Dq/qwFvjAoUEZJxV/mCpfN6
XIIMWRx41+CMeZ48b82l76jAIqbBC9RbKuBth1moPC2Avg9etpOlMqF1X6pc5FM6
oZO/FmNMJJfAm4D1SW1KeqzhJT++E/oKmlp80rxoTpjKfghrn+OeD2LGJzMZFD4x
8aK4wHs8Obr0ueInOu+ucivae3cpcc4hxuWtlOrsOl0A1sAL3v8Sib9L1LezdFBE
RYtDxAIrvEcr0N3bSFr6wnmealmNb2zkd1hoQmOcCnJSm2MzK46sRPqI9nbAs5Vy
y6sAgdlOehNhlsmYMZb7jB/Nfgye2Nz4nhM6AWPry7zUJ4uBmonOaoXlipczQWjg
kJ/tFmQ3P2dnJkM3d8pq2Oq+kgvzHJTFdfv9WyQObyZHppV1OQFUa6/km4X18CXN
uq7UG1x/IDUWn8rYxrAs/AN1i6nkEMiV0KyW6TK4nhI9NGDyws9K6BT9daNvIE50
gsldDPOWsFz5ASu10no5AvBRz8YkJa9jQ0hhx3r9eK3gP91Igy1/MseS60d6X1Y8
bpR3bYN/i7iEEi9kCA+vCX3T4Q/O0oU/epy7K+b59Ro3lEXHXfNwQGY/lmH+VR/A
n3Xc6UXYr9zrm/lVxCmO6GxImKin2KHPMcuGKEINBvFPYKoiRfdgposCIXphyA7R
Ud0hvqemLzN5AnwD+mcwXZYWt9os5OY9Kn3ykf+VaM9+/SL1eAoAdKIc8qKIrTyX
UqfaoL7HEMCSQNMe8+zaGcu/NVFm81lXrjNy2/q1BN41Kt1XRhc28JGvmqZ5Nm4a
vezMRlbuseRsMKA81j9s26ZVrWCVdnpVXdQJjkCva1QFJgIPFtXuVdMoMRvLYHMk
KsuddbRhdxD5qo/hgFF/WRXH6rVPp4IauNxL6gVvmhBuYuNbcutRgluJ0REAH+IC
tAWn/HaCZhvL9C/ceZgRy1IaqCYu9eDF1jOqYL+2oBe2gxyETtU2Y3fOKI5jgEGF
MztFRCAIM5ssBP7DZ+2Q4pgBodE81safuwXqz9NJupearLW+pX5WHsxWNI+CF3gf
0ZlyXwqlYSEt9xC+GeFIcSW63XIoVBIwn7/51veI23nxhpf/EvOHiKj/Ka69GLCw
BoYLMku/kqye0mc5bjqeabaeRX21Vg2cgR9qJQEERgDbJAdHYRxMNWbYbpPduSl6
MZoDR7eNyvhXNFc+Ej/2paft3V1mS6k5MXqM17ioWfpwxOy1rQ+pFpEhaOplWbSn
fPJAtOFh3PJRrnVclJOFcOkYIYc3FFwBdgRy214+arpgVZZ976wZ8OrcmcQ+HPGn
xbe87P15eic4UEtEqYHvuprVThkZf26dqsBsgZ9d3r4alxlOF6vO2ij/ahDFjHuh
17G+sf4p7t95rsS5byI5z5pscXLj2Qd1dcXErxXp/BVLecTFEteUWVxzlXMkd39w
Nsm1tYl9ZQG0OC/waKmbexuzgMENWCvCuuHJjQ/G166xjnsodxZUpjJOWBpUVBSX
hzjDEn/pUqJzRzDFC9do0L/taoV0EFYoV9+aMxDjjy3Vu8B5V0EepLUQx4xJXtMQ
mwjeShKY5efe4gJVowH4ziXm9mRssRl8qksRDIT3c3CyR4x/RISgk5wnOJeh3rb1
nfWGH7rQ0dH5adMalF9MqYyY7csf6UR7rs0fRJwUoJTbH698Mj/03f2sFal84pnw
tUiin2jfKQXKKy4IQsDFItnPFgRak6NBlvQIrTJ96xozMSLmF4Df0bfEM6JewEVM
DpaJeoyn5sZbGOo2zakugIiJu9qCww9vZSvC7dQ2jrFs1YTbnKZIW+CbyOQZUu74
4XUS6xmwFvQ3jIuZaAQfB3CQNzi3u/PGMXUJwjKvLSzwa/nnH4RL1CvTchSqZrdS
qns1dD62agcMVuemlsVbauuj5Bg2XIDLGIpqtLItgZrN1Ra3MAPjWAYuuCFe6rci
25r+FixoDx51Mna21UynsBHx9JvbceYyiCw0FSKrNAJoN6OJQyObJehXC8qlcDmz
yqZna2lg7ju7iQk9neTdsakZtHvxVOEh8C7rkf9UO45exliSoYE7wp345HHsv48X
5gvXqRv2mLcC48XobA7T7iGrqe0dCu1YxFEAQ0YgBNe6Xa1Za9+qcvActkZEj0hA
hee7IZYnkV/Mc0mUyOEVrFtK9HI3wiBkqzF/GkS4dquWlvAK7sXRrxqrNSHulCoc
IKwRxZusow5e6EG6kkVUxPRd3Ej7PFqFlayd7+l92jk0rkiG1iSKf0pfl3NePqSn
vVL/IpFFyJu0zqwdrndrVBNZG3fqcQ4Haw25IsChX0nd0GVWDpTEFoTbMHsDpYtq
Firi+/a6Nc/t61MD4JT8+MUCndzPKHBDat5jN1WsTVqLsNPPvaOOZiXwtrYyQr/8
Q/inKByl2R0ut/+58I6D2FHccpNIwoxGnGPCDoVo5WG0P+a29i98vSprTriQFyqi
Cp50H42KEw1ecTLKMPzmu7qSiUPF4Pmv1Uq0NvheN/3LgKTRwP1sdSD9ys6lykR7
C8yZK6czxGeqaaksXXtjh5/u6iNuwBcpzDOV2lzvFE7Of4LEV7TbsCa7rnTaUvzf
faPOoRQ7DsL34H6A16VqxmG1ywikkSy1QzpXuN+aEThLMdO1FGjbQnXnqv6yFoGy
mjegrqqSEEHKpMnwEqoK4MTi0mqwSYG+5FBFj73dNGrQwni1ev4y1ak/4SHXPlWZ
fZLgWSqZWJiCxO2FnvHkeS7WuHsTYFvGXYnIo0ivE7OTZ5T45jS+F2xSN0zL+19v
J/kho+w6f3HeZJ9uYxzN6GsAGo9jBejhiJjB66gZwav9ozjNn32Y8TJ+2T5Zn24t
NRkWxK6IboOGzRshtyMZhNk09/W3ogbDX4MnDqDz20HSkw96LSs0L03Z48Un2EDB
8vgVm3dqdqB5YuWLlPIiOxGkmy7SHe98GIyWwbaElcG6YM5127EB6mZaNC0fCspf
/iHa+x9nS9uvWNfGpnqeRbsdvl6jRlthbpkQOJoQkqwIcUoXhJNEFndtyHQ8URCm
AsKKsZ0WrHuWeY5RYiQlrJ6IfT5m7w0f502gVr3ZuzSOZKm7FsSMeZZBajnbHUiJ
u0TYT/E1uq2ljo7JrIunSqv9NaydkVBuiMtTIzjjS8qN70v2OuPIvWEvdlVZJ0LJ
xjdHCzERG+dmXzmpgDqXJm54+bl4G7KL/BsoN4+70Cb5MXBF08JSuOhrRwYxHx2p
6VLz0JeAuPn8td9O1qKSIOV4auUvpANACmAmnMczBNQJHU/HD//UlkWX/fbM6EBA
x+l86wo2gHbU5zRTpiLDQ7lk5xCaY8zd9v7w6N3Cb9BudIMARo54PspkgABp0hD3
hek6+Xx8xcQccQKwmSnyxTXnhZbgN6iV9iPgXQVsrbAJiE+QXrKfRJnIXQwv5ebX
Su5LdXThNv2l62lT7U0KXKQRWrd1m+XMjvGYERDzUY4bNDOCbOYKPg2Wyy2ufkeJ
PIpCQ99XXep4VTzNv4rCt6+kU4WIYROdn4bHiXSpcQS7jTRgrDN6pRtjFNoxbexy
Rjh2XrmIueIM5QUzlY54F/dgXMI5S/IibAkGlsFXUNS/E5QdqgjGncK+9wTi0cFq
Yz5JPKGD1TgXmgdCpVfoGVrRk3qJs5+PJB3oyEpHMOYvcJnyMpQa1kW/fRQgnf1s
pVLAAzb/5Mtmh7+muVtXfxU3SKsm1rGD6uOIAqut8c/+7M7VCFLaCsfKzz1aQ281
amgzQZOydPvgs2jxRB6LNqNX1XDHPk6G7HVLpb65T+KFr4r6usFlJzinVJigYsbP
rORhj5UeIAX9jULMWsW+/88TyRf+e2i19tQa0CelTFW9dKCVxlaaBEv8xZYlxQgF
vVfBInk0xMOLaDMgbag0+ilKRMZoKrWGcrVah9XhojHKBnRGEJkyXUIt2x+3tOHm
b6vWVI1PRz9xa339LTgWLpf1CXfjhRcFRFT3wFuQN4Rqb28E2NXhnNw1sHrRrMg6
oOyZFcvF7BkBbiyygmntyebKLZXB+STTPQAzYUbDYKwjtcJnecznGlUv3GsDd4JF
V1or1Bn2EKcfZtgAH21CzkqG56QFhs57i2YPCok7/kFSa8CXEWzTQAHjepgqhPno
gYOWU+IHd2cd2+nn2vMvOFy57Q296V4b/EzUwg9STrfDkjb8uhQavLmj42jjQFHy
X6gCD9rZUUfJlRy9FkSI/Q82BPY7VRZiB0EUMRmCX6dcp264sCEx+h5S3FpgWbzR
r3lER12l+0r+0+wpfElgLZH5Z9JX04ovpDj9QZBKX9ew27tL2itMu0PV6ZqmakIs
Lim7UKoPMYJ8mE+kD0napUHWiiUahGmRl9DuPGoOabBHTSh3sX0J7uVlf73t5+yF
Vayjj+z/wjUOQXW9rHRcZHgfEE7Rr3p50KAVE8T53OZIqOIw4jAaVmb3yccu/Ot9
eE7vvuaNPcT7qt+Mx+UR38mptSTB7daTV8PmF+bVT64pkm7JwEHOhnpOF7cEzade
eOwhDEdgHMsnnqPa0Hz94si4D2yeDclYTSo9Mal5Hhs6PgFXWVeedZNj0DM0swnF
V/6jzSvDIjbmCHfS0DrFHM2lVv3ZFMW2mEK1RTM0osjbUuYnYhnX//r+gvmnC8rA
1jYpWkgDFK/zmQoaWQEzPpzm2cOE/qnjydKNu+t/7++L6UwjMSn4Kv3TWp8Yh8cf
9yoR05dPb7+OoZhIzE0ipurPk9sA3BG+5USLyVCWowb8P/imyor1tQb/LKoL+fPU
R2Da6P5hxMNKlWsfB/WwZGFSYYtHy1eBEstBWBOD0cbzuoptRPJNBNpJqw53RoKu
EBuudKmNFHMqsHUwbGGyZQ4JZKCssMc+6q0cSZmaLYl/mQi0KJTOe15L2IY7+XzU
294c9SPqV+vCkP2b9UmufYAA6nedQiVsBR+2EQ/2NTbDq4GqQB5xqis2cL8+NnfG
WkNt4AMWaH6w3ieojmMAZPQnmaPjRK5kR0sy4d0eQKdUoR8qah00+pR7KAxuIVxK
9V0quIE+jlz7sD74tmk158r6lZkwk53cL+ffwyMS1/SIkBKj+SDsxQaeg1Aoj7q9
/q/B7IJhCgsL0Nw1jhJ8megw264xX/5q5G3HYZgzhVKdECbh8dcU1tYLKYYvvTLe
gw343YWZYSArscDCwit3xU4gAZ/rgJ2yWBBknYtbFCxuXmvmYQo+7PHRa0ltFt+1
ovB7A5z9zIIdhZbESD+Wv/78fSTNP1O0PaOJShxgBfbFc29TSaEWeMj/xyXlpfMe
Uu9HTJQCDi9jmjh3YAAiZIlbaGSy3yLvSOcDto/B86ooibMKG2nOnql9fj6Gbm/A
L41BGH+cg1x8p8SAQRPg1uDlSHPrsE+MbQsKMywsG96qrPzWvBn4VeTjN4fFh78w
S1SZaB4ozmI/GS7WKXK2F/WKuliCmfEZgEZ506DInhGzU5A9I7Eut/cIKfQGzYn8
1V9B8ensmTuMvFhQDEO4CffsOowDiaFt6X77aNezRcOYBzmJ6mh6zjJRz9EpXRff
0SoOXIn9uriQyWjZZ3nMmaaP007k20xvpXf+A+SpCxq98Lk5bCOXjsDS4BLOKcff
oa7snDoioAXvK7CSf/2d4GSOT4R5ak20YbM2fBlDASBaOlcvHlfZcIqmxXjgsmUE
Rocv+u9T08CIUgSIRPs0nzQ9oTTH2wilH6BmeFpjfRv76LA26566HZ00PPWUNnXh
aL0/Y5Q21W+S10PIC9xdWDiUzQ8KiC4xyN2/JzO52FpuvU5WSI17qbzvv+vM8rd8
x8RPzcsV4s2FAhxkFUZOiHKLTBy23dZQJN+UQcwf2WPthUZ8/oju/ZZnR+uUCZU+
YPVXCPfQNTlLvYaT1bULy6wtvsiaAerbT7n+eNoIw/3JrEQC45sBN+vdijOKNHwj
svzL5ZEOcCa3JMQBDgnjY4Zv0FmtC5Hyyc0KXkvdUZ3C8OCR3hczOXxpaELXsE8T
xS/yBvAOHcqdNoPzVltMoaz7W7amYsAxjOXswGKWu6WHiCO0tJ9MrcDHmojLiWP4
9dmRne3F/B5IQcg6K2Q45ylhQCu1D0NXuLx5ZQ2AkTryf4Lsee7dBOsEzZC2xtkS
ALHu9Q4ngrL6AwhuRtn80AL2Vh+l6Q8+C55hiG6QI0pmYibCdP4H5uEAXlN/qQ6y
vAzXZagTnQ9VrggEWIu3YCuYcQ6gQ2MMXDWX0iNm0Cpd3tvLBURJjCatM/pDT8R9
4wt85MvJFWz9/Oh2fkm2iDcuFDjGCIzI9zqgrehaMlxkKvGqd3dFLIHpOqLhTCsG
qu+8mm7M90EfqwBPYYY7aAFBTPYeS0rnZ/GOXEiSXdPrKBh36I6jzo19cJTCrjR7
wKwRLzwTq6tNJI1A1s8vjO1ZsygRD7jQ9/hqh5IJr0mtlFXXfWe9RuCOIOnurmjM
BS0cCIRoQJbBTuhcFfsdsNjrSfh2viKeyAIgVxTvXOgz6/X7PrV0Nuabl0WNY4GQ
lD4aDi2zL9JQWjI+jS1DEBNer3alyvsSFMT56wz9Tr0QNHmqIOEzhi4vBWqwnRb2
53Bm7Oefia1Zi9a6Sw/fzn6BI2iNOqAC7sy/zRNKbli/kp/88kJ0AkKnmZHzndfA
J7Lp+ygyQ/BRc2jJRrfOfoQ3nGdiphUNMYTExqBKzOfxkRj0RbcenjYFq3f+lZuB
3rtTehbQSODS6fIAK9jGtXK4T6haTaRG2gYlvm4CVlb0BlBA/N7ZW6wFVFdhsZCc
ZqXPJOB7qrU33COEfitU9yywceEjxPf9Pyr597WSOxVLAdKML+rMDe6RjUb4jha+
QIFeP3xlRDykNrrZF2Rg97Dx4sBBq/dMc64Og9sGKAXUsfEhZpexoRfdtNcwfapz
64oOLwonOor0MZrc6fCfKutSqz37u8H2SBiR6VlOLNxpQLceDN1YazX6IlhOcaK5
/HKo0/NHloi6wUwuaLENZbmVLQKss5PXh2EjYaqTWUKjmKrdtwnKh2UyVGFDDsDw
s8TFzhp5emzPALMYHHpKdoawJWD184fRJr9s8R/3nvnZpwpo2AzsFGjNMKI28Vwn
C2NdARo++aJbnFKgz3XZhwqW9yZT35Do/gs0P0M8zO3Eq4Fp0xx4AyLkqewTHT8Y
vnyG1SSVkrf7VjjiAyzcn1sP7gX6nxn9qkIghcSAMufOsptx1XpJUcKXp78xI2AS
znfLDf/DLbnoAFvB+6XSeppziRCCDrFG/Z9oh9IScYY6cW9zwJlwvmolqyOTsYrx
p0svd1ishRCDCXcX16uWLSmv1KzbPQTDzNVOV22Rx3A1e8VzBeIsrXz381kLhiHI
ZK3Wp0GHuWYcoF1o58nKhl8vTshJeHCrRiiqNsqxiYdzMqTd1NrQUcW3wXpgx29K
RkI7xTpmrGP3E9psE3GkEn03B3o0jvgsCu8SEpNXUYFqWzzaD2aK7OfR69bZs+pl
basCK9eviUAx2ShIunNC5FFEZBF1tIAxRhiWPVx7JCcT954vwpss6Xm9TaajMknw
Bxbgo2qlO/ONFqSsgG8D/RXPBRt+yQcrfXCbURh8YUAF/u121KrL4ynoNkEXksBe
vCMKnbksVups7RvbZto5sorUuQUpIacYQ5Qe8rX4yvJ3Q3jLQDqbenhCzJjCnZoi
Iyvzi/zDpRIAF12j4WaSpaBBbe9phDvoi55QfO4JeQvAR7Os8DslXBFjVJBLk8ue
deXIpw9AnZafnV/WJkyYueuy8Bczu0lVAm0DCiYxREVLru9JYY8Jatj5RzCgAs2K
BzXIR0jm5OWg6nVefpjaow3G6lB4h0utxuxh7Ukfc0Z5cuoqs2CbzY92M60KCvvp
XsCeknyzVXMO/Ih6Pr0e0L6Zxn1O4zokyyHwkhDijxlg8JbvNvj/iKnnkfroPTiL
S89mWP9fTVdYf27QWYu1sh0QoaZqj4jiS2Ntb9wwO+qHh2xNHTk2ZxWwbazaXnfR
KsfDhrtwMFPAHbPsnLueotDlHlHEACKwG5P2HQYW4yMrr5ia6H6GmVMyCjHvHGwG
0tvy/U3VBrycuYAF36o6mBk3nQm2YLFvFua3I/t9tf3icFMzi0GnB1DKXvs2Y9iH
D4kVAlNdT2W9JiTeDHFhheYlbpx9HMy3IS4RW1r9i+tLNRXabNvSnLSYKZXWiVqe
aL8Cw/3ucrw7I0VdQqGDHIXYcl++lIs1k9qxv385wHWNL+Wiyyujyx2f2rvKs6tZ
Z4i2PygfNVlhdSHOy9h0qll4xWkH9vYN9oyiK9/QAtcpF0jL+gzjX/d44A984XcR
WBxXNKTDiY7QdHLFF8laq+4InTfE8lUL54/dCMrXJAWl+Mp4XoauWxvteoPfPldA
wNKfrlq2y7fSD2orA8x75C7mB8l7vPMkSh3tI/3TDUUDrws7vxG3U24u6t+Wlxta
YIb6zr/pi/vDl4a+1G6O5cbEBCjc01g7d6Ygf00XUHdUJ29SvLRHrNQEqU3WXc+R
Egl2ICh6lSlzakHfesjMve5+7SDGgZ1Af/7EaWJsPKVUY4NFhv2/oClORYXd5vdM
2xxmRt1gfZOCx6tJoQ/ErZivnDnMigOizD3aXRQgtRT/eePpUPYrnUi+k7FvS3/t
bzsyEmrPu9m/Q3NMihjYG6FU5OhLtmnWgLjg6BTKcbSEpUkdRSE02D71rplO+RIJ
AtVIpXMJe3M7yhBskaIx2pmGYsa8CntZUvS6VZPPv5obwvBJzVRGs7iasiJ7OhQk
v3xwJjzXv7m5C4kZSsuOyj7BWUxkWIEmteNlQf/L70JMuVvU48oLMo62BHMdkteq
g3/L2tUh0qiFU+rewdhLB5dv9p9SrXEqCC3ytU7EXP+SS2FpvpF6F9ju+FiY48Tp
JvAng/t8hS9f61AUOB03mHYv2o8Jy8wA8vkhCm//vwmK1TEl3lhf+yLvUvE1+4uu
Qois2diiVNPpaqy+U6OkL6HM9K7JteUM9eJ4xX1Bjyyifu4o2vEqr9ijQCZoQpqL
4rFgSGWwYaZtFuqR7UZZPYLj9wKN6So6nLRgM+ZuXY2OyoQfcMI/zuLKuPDO7XDK
QhI3CjXeRXG6spqpYFdeJ5vy2fNQFnXaY4oNhgZqmFZPCutIMYA3VZ+dsf4Vd27G
Nu7aMJODM5GRMpw20dcP9PXsiY9jVgXn65G6woBRFZw1oATUWofcs+2NrH8EusQX
AM9DO7exPLgbfbzB1FQrECv2/fgzO2aQVKHAATjmZYsFB5glw3isZ1ZthqJ6t4TI
dzaK5tKuJQfBz8dr8Du80b6LVQMqETQfr4UIdDkOloBaOwfVIqvVDtqUxxgLUKJY
hanCKM2IJaSWUbB3G4gS9/JiGU69nEpgytSPKdZXy7QV+kqiYJ1j0vA10E6XHz5o
vWgN1aEI/kap/zjGBzeaaH3WMPydyOxowQ4M5pPuDLXFga2njS9ILpCoNnfhSOf9
anWD4O6tQEtdnbBFj/feTGZwPd4NCpkRZZ3hzs2mrjpz1RpB1BziA58Yop0WdSTG
/BxIVBd0nCtVJYFF38MkF+VHBbadsfQXjjw9wsZGyeQtbWBtIA56YKAr+o7Bbbda
22SpVS1kk2JG1jD0SaWVW1+19PvH/Z6aQOyODU5UVL07OoskCnDQfJxFOvfQr22l
eGFHE75LioR8EYUqO5tIpDQq0xPUy9OaF7S3pAVQuCNKgoSMMEP5eMzLblWSa8FJ
8zMDrmLf9HTR1h1xAcrGTP7rOwb/q7ZbBgRTqnDJ7NbiaB0ZZc1OjbbrjZQfUVSJ
J7sjbvMPN0l8dqkWTukIXaMrWXPOz/20aVm9e8El2UUt7AtiOlJB8xXlnttrdO9L
MUnGX5HcxnaRbSSZW/BH1eKkmv8auRbxzhyWMhf51HWxKG0c/9d4h62RLXpberhR
+e9CM3ONCeIOpMorKbuvcX/X+j1PdEwnQlU8tzd7QHLCiYQ1gCIFdWUlRI0agLje
0tkwc4lFzuD05KMrmG4lVH3AhBtsnlYZLDF9h7bcUjiII7tWgY08gkZsHwHS+otj
pI/W9MAGQfEkefNqReZnQoc+Vtti1tsCftJS8uvRDljpTDjdAyUO/ecrl52Z9OnF
YTRrLv8h8OyBrQfMKNRaelkRJKDG4cOq6E3h9aTFNcYvQZ8WOgbOj4KxvtRNWO+E
RthFuw3xMLlXZ0ve9X39QsupmrAU5f4EN8Rk9DbsZZo+GqCeTk/jzvmAhEjshF00
4RAG+sw2ebxvlMCHk8r+r7o/eMiu4jHa1XsI6570oa2yyu3Mze8m1bKQFQlhUJRG
Y21SAeP7LUhuT3HzJaHGTqxBmbmps0Shu684XwC1q0t29xQTWYEfdlo0o8PFAlaP
X2HohMtfLCjJTihJtRiUtsAiUzzzO+wiRFzuyR1mRH8A0wRaA8lTfF4xnGM9Oidv
2ewVLPqdcI1B3J5OyhhWxiSUkhrpDgU38dksetnVnQjdjGHMdYf8GWR9WxTsl7T1
/Do9JOfz3ZPwuV8YjJvdCuKMEZo3KlK25Z77pTFHpHVlYDo1DueezZSkM2surFtn
a9PT0u4X+258qAdGb2RrHDhsj8Iu9uJAzJLONALp0SLktKAgi63JEE8nbe7Y2qIt
zdqbrUDG6Pjd9J1VGHzn7tZZdcDQFRgO/66JsNZGAGXAdHvkjDSAEO4SMR4+EqTc
Kr54G6bJF06IW1mkkoFtPCzMfaWrLMv8fS4pRtCyu3pvz/GK3d7BghxS0ZC/eaSx
rve4biwOhvADkmDIfhsXMrnjkcfNL6uId0tEr22JivZytpgdqKKtbKIO5fethkLr
gSOnbc6HBawQCiQOiEnCS6YVi5xW8hxBe4+PnM88en2HH6u+pJbC98kPa3jnCrKT
yX/5s4qYk8rli6Q2QAlNlN6jaOFFx2Thmg5IC4NAKWUSnUKjGJjXvAxYCgW7Joyn
H+pU3TTIiw6C2zQNeoadqBQAIU1i5zfY/XM17Ah32NT9OeF2UVmNmvGpHAbpFf4/
8oN8PE/B63NZhTs6IuOYcu9nkTAiCitYuEbM2yAvyto+Dnac40dWw0BEooAYSpMw
TjZOpFy8Ojf5ObsziTksgzbcfgeVhezNSXo5htnOOnaFkTJyr8X4bpz/pscKzLdR
xH20Plmqj3J/c0Y0x1q4aWF1PEYYrH2GTVbt1dw648KvG5HWhZkIMyYrqD96Qc88
0riL2XcsdZKzKtW7kIUrDh+3bi5qbZUF/RcT24Ql+dGDhkrd5mes4CI+yZhC671h
keHxdmSVMGzCcHvIGR+7+jD9liXkweN+zfBGGq35cTo1clslMt3uzhXWg64vhqww
eZe+07xbPVTxoYPku/xNljUYV+wVzwzDESmGBO7AcvbPqqQG/ooB23jcXLCSEEZw
PTQNvM3oAEScqd0XRywbTYjseMw4KJNAQ2qyXb7U3iUKnJJTvz/uKFxHZkNF+VpG
ROhiaJmPnzCTczbtDaczmLuorbMFrnBiOdtxb1P2668wEWFEJ/axrWeCEMwTO9l8
hzwy+iYoYFXMJ7LRrR6lrePGJfSQhbXV6suwNY0+FJR8tI9HuMORFqMuMdaMapKQ
CpiKmZIFg9RcJ4ktetn6Z7XIvGJP07vY7ffvvnfSFC3WewN9galazVYhJDvjf7k5
YNeNwaB34fgNY+wph59AYWas9M9ev1B1O7jAdrZofw/S0+wbVQIvvTw5mJtyqLFg
fCCgNKdNEXz3/aw/uj9V/3+oebsfrMr507rWIfHK+xe+5MjijMqNKljuDA9PGEoy
OSeo5aIPyex3vmTqkWM70oKxRBuORpo+qzt8VE7Y6YUEBreIl1+79DN5vCxOkxlA
OwVKtJIrdQJmq871oHMG+os+RMXpZzvG6rgt8NNxYxNTv0KKubR7cmCAtvIu2kwL
awA7qv0nNVi3aU8zA9IoiHUEvhvmlYPpsqszV3H4DNC1j0giMzL1wk6p9Um0fy5G
zSzuC7EX4TihYwSXMCrEIbrAQwNSkC5+ds2BO0WSXDkI96eODPvW4TXrkS9QR/rH
FhqzfG2KY/v8+9zc7zN/pEUsm2lNIrqx+Ezy14CuWnLgX2JNC0bMEC2fOMutiWo/
oRrXZvNRWwWHYkSuWQwOX36y58lSIe7C58f9pll23ADBgjyV29de3g5qy9SIIcr6
WC0t1zUUArPiK6uxcdb6zKfDbYQ9mDY6obKRL7Qt7cl8t6+/VqVhctGpqvCLvZRb
oHN9l/ZsxbwPUdk7r3vrpSJ51KQlsrDWeKHzsfyMW6cUOSL0SRma7Cm3vynJGUHS
K11xcIXiKBKCFsJrGVJFNMOCfo0GfJkcfe/MNZhA3zayIE25a5ttxBzhfn8Lbw4o
Y+es+jEOwCXPq6QePLRSW9Noyi+32Hbe52VBkJfjmts+GHPeerVPXioc3zt2S9CS
QA7d6ZJBSOO+5MZHOpo3GY6WftSBEAs9XLFp5KnZnXfPqhIUMBnkFhbGrTirjerZ
O3awYVDBsLsd4NJgXuvGxrvMetlj16eOLQDP5Iy5XZfD1wD+vxO25Ru7f9tZYAH4
6Wiy8YMuT1vEwK55yXlvP23zHlCgQfNDdUzy8GG/SJcURDinu1Ym4MWWO+r2ASn+
i4yqZdNz1D7cS1I7lwErEbrOfqaRC/NJGuUyYJEdVup2bzKMMcfnBVGngahf6WLh
9nsxaE2bHOtNx8r73tOw5IfO5bb62Hrvd+W4G8SrF6QOOjiNp5x0l63Zj4V+BG3c
3JDXd71zzHgHRiqBbpvV3V7C87Z7zoZ7ZOQvCenDYK1mIVn7nzxFVqkIWD6mrqOw
lVQreAQA912zBy7s2ixVvNjlGcHCxBzqZHGI9rlnrjRVPak3AM89DeDhqwlF8S6u
Q4sPcsirFsKlmh95c7C5Qzt3bCC4Z7Nehs4XeFvFEazJM0y8ruPLfK7Wk8u0Z1sn
hQ9bfbPZOD4c/85nsQYmnkmhnjcgauLvaEEOUnDHvUkzZ0eJ0/pOUuhnc5R6Gv25
9rCh4ddSc2DewG0TmiZsonxzJSrmTJwIDxbi3Ly77+PZGD7ZqOCXrhr78mhjldn+
KOaCZb+0PqFmgFPQORG4vPVSmniSTxzUPjrzRQtfDd2aDIcMiwj7m6xlMWKCTyd5
gWykgXToVPu/lQSTYHMlEZG7efWPxiRZhG1WXz6gcmbAtqhyGBQbP+En4IYk3t8o
PBQu/aWRW1iZLf15zzdmS//SWNnU2vegU4Kqvhzc8pE3viXPptOpjdTBGqad0UB1
hjK1Vy+5PPQOzjCZ7sLgur1p345DF2w6FaykZn5OhnTZQVEdIiiNwAtQ3ssh/J+T
CRgaYQ4aN2nKx1MuUvbINoHxQj6xi4JWcOQ8zBApy/Xt0mL2Qa/gKVoSkMoAik/Y
cYqCt0gnEU6m699VuXOQfYH++3KQnWlBOuUYiw70YaZU4K4ByyMpn9MqDhRhM3Bj
NAixsxEM4HLyvD/iLnHttO71AJTl/Cc4//COLzSbiu7KS7PZbt/7oMi+v+SfdQdM
x1VZOjvyU2njLhg4kAshtPseIBmLSEL7ZU27lddLGJZVam5xrOXg/9XohWNeip1O
SjQbLMefgvgu6+hV6miKkyiSdMP0secqGQI/tj/sgTx92OAvsUZKh/g0MXbb7YEy
z3t0YMip86XJcW3C8HyumoG7AtDD9wJYGdygaJrWXorNey1snm/l3Hx+h6/ostzN
ISuZ71tMcGvNryM/U3IpAm+H1UBsCn3kKpRZgjec3ZHjZqXFlX9gqWRFufhOqOKj
xn/8HvFBGWHF3HiFEllOP9q3uBsfKxeSPqIVClbD0Zo8vPEwy80W8uP9qBpEueBk
V8CeIhFpVYtAw1BXLamvDD9SXExDJ7L4AK58oZVPLjcL744Vfx+LZjIqkkTWxC0h
L700TmBbSueZ66avuUkz3azdcS4oZxsO37tgDUon70S2nBXnMhYoJoeAeUCXnGrD
iUL7yDVOJnIobZBoq87zItnpyNzlWyyu0z7hD6XgD2N/fXASX/CDoSXiig06XfzD
2EQ5RoUwUiRPs1VzZo5H6Lvses2qpOvRcNQygZ7jcaEThuuberkTpK2iwtYAgT4P
BioW+dIAW7kEg0MccV1ExD/qzzc6N+t5ntbHAAvgJ6g97jyTlszT4LSUSbmIurEa
IceQWyK1dx7KdZ4QmwWbqR9exLe2AeTJSHZql173vmhp4eb2e7pPHCWRwreLP4mU
z8tbY65T9df0HchsvSNE/fbi52JyEsAduff478bZHQy3A/Uv/gDZQN39ClcFRrzu
BQTyHI8WY3WasrkzFe+EKVfxqTf/bmmM6QK3s8V9wO/AVLtvP8HUQuHquISmuzIO
U7YdO5R6befHThPM3sNzMUDR7T2N0kddeNQi3+sPli8oX5iBoOHrWlOolRBtht/E
wtWWDeBQ1BHTbWAAazcqtxX4kgg9C587s6RmpcVURhR0r4LpWoG308J3QOQAFruF
/+t3NT71k78+YRuZLJte8dVFjIx6exwuSUzP49rhr7KBdPF3eS781cNsFM3R3Azf
/w3SHoVW+SPspQ9yTwCRzXE7gfh7sfDqZEoHZ0z/7vh7ov6MTJTel7E/2ladyi7y
VCtLap4Hrrs3OY0MWAm9KOZO8qiDdCZFfeNmYInuFbX2EdD/O7TLjZyDhevjH5+O
kegpt56V+JcV0Ade+MLKtO8ijlPBtf7PwsdpMUQ2479Wp6XbNDv9r3ka5D2PHC1+
FgnSoy6SmpkVbAaZYyyZSdQx++yzk79eaxi9f8Uq0tgbs8wP3ORk/gxxY3cx4MBB
BHCr9ULL6n74mE4u0KjsAnx9NKltYfMrNv//sT6C6GAE0QyZtnfc2h0yJKp9CEGf
lJgJhb2Bq+RMWZRVc4JbMUiqIIW96YvzbI0jUTFV8ZKMo2fmMdHI6upcCRhiruTd
dEj11fvLe5kvHTol7MI111cf0lF7oLJFc8E4imaluLU2knspOhaRaEFNESaRvYnD
UkXFVwr+gqcV7UArfcuraRSDf4yJ5XNTwcCCYwUfmF5Snt6+sweBK2UtwV1LhlaX
ZO+utHCqFILHEpV8TUzOH8le1gQ+h2agh2O2slh3ND+ZhAhk/tXIdCHRrbx/wHjM
4D2fdbGXgLh1cj536KJr7lsEOZmLUNAqyqkuHxBZQ/XR/1l47SnUc0JdyBp8hcDc
mcGhPxM8QoHBQ3Wyf544fWfwp+AxxWRemWTGYNmOhgVXtcHQ/QrCd6pniLwr6Kk2
LHfjArT0gpDqrOWEpQMxkRl29+AVD/QbBoG4QUrotemppF7JsCVE+7yCK4nk9sH0
f2WsuT8MpADojXh2GBm+mmgeTx+NmmQCjHvlfgmbjU5s9XLzdn/aUPEDn1Wb0GkB
goB4Ykc13P0NN3jFsPnIt50EoCGb6E5rtlF0j6Dy5k1CRZvH7W/ervTit2FkQSHT
OzJyvruCBCAepHMRTyzNG0EIyifPpQKGK2OwwACv7V7z3YAlSpZS6/Rx6aOtsSbX
L6Gm8ee+RI8U4nrWjSeqiuNzDvI+CYugQapYZW6MRFR1AWQ9ILj3rEkBx4TFm2Dg
BDUQBFGnKOOkkmZutpczZ/UVN02HYJs0APr0jQuszcDxv2pJKVkFqLRDxaqTzqzo
EyTM5DT7qTXW5FRt0V0MUbO9gYHIe+8VhHBWKYoSN+nLHM2qHHqQNG2cSCuGLy1b
LEoC+H+XecOzXzdWFPDACz6dhwqxbhul6TGqZ6HcJHVclxJAdIVPKkbEXv63nIz7
F0EdF6BOYUviP93g+KFR+CC7cAnieeTwOl7B5n4nWTBu4Pj4UDEXeF1kcrXmRsDp
eEddxjCwzJP3K6dNA/mBz+QaIQm8hqSd7VUxIZITljbX0CuJtYObW/jcJKRVGkEv
8+cbK78vaSzW9YiuWb4qxn3G4sMZ2Ff29awlKLLQspmhjT6OzyqM/ezSZh+99hNp
xZ9jKYsi9FfjhQM201vBR9Yr2Gy6YQPsWA422eXLZ14yhTLlspcgQhd6uYYD6vWp
wDQGJbHA58+4e1uG1XBNThLGtSOoww4JpNORl6WjMVuAfCjfla3OAjfL7gnEojDk
AlkHzJYMRmdeBSKWvzIB600EtyLa1KraBLUXWchMC13V2hDeyJURJP+cHjLdV7CO
5UDc+Eidw+adSo5c9b0Ne28Pls8n0cbNbTafst94Jw0XghVd/zMezKXNOD+ussTD
dqHYW4K5g2eBIymLz3ravfQ7FlhN2mGKxgHhnDWOys2vf4Xml7WIV54NkWeVZcmK
hVSMFHwDSo8w+8CWM4+1GtRW9TvlbCoWnGhum416T71Et9ACGrauP5tM3b/ehrv9
28XGl+lz+5w5KWnB86QqwGUnT2wHmjptK/+Gluei042xrxR1F66APhorURFnbtPe
avymDyKFGH8nTf2DUqPzUc+DtFX62XFCZfs8MrmaU3dTjHfZhpxznOIrBGHEBXeq
tqfFXeVkPWBJytcIfUtLg+/LvAd3URQ/9cdC+sClx7MysARkyn9mHUo+XOb9kLKT
KLH/1XzrFlSkdI46d419ccwa2k8LK4vC4F6dDQRKkcDBW76C6ZbvcuA308ti/arN
mLRYwS+tw9WMPolRu3qqtV5pMTruVLx8Qnla1QuHeg+ToZMF9HJ5MBx12MDMEuCU
JnQBouSMz++FA3ItaKsGZy3qgwFKrnEYoguG4xN6OcQ6fDh765HdVIW1ix9hsYOD
o1+zxSbe0yrSVJLN/eiOlDmMVuDtBZy5NGUI/qNegzXcEWQtU33bcouTzRZgDD6N
1icyO+Et33I/+8TRp6Hc1Kymg9v4Av7QEJPMeXAua+rQE3skCrPJYmrJnsQBYIUJ
YllzXsN3eXYR8A19TAn4VpL1alY0mNH5B/mSYtaOnpJbkN6sC3xeaf2MKVATVMEe
32j0YESIwPn/KGmzMQ3g5XdjI3s9zFdhIMllGxrmqYLfP6/fiOrWerwb7xRcDANF
mD3Y8dYzVUcQSuRM3BO4lbopvr5U+BAEogISFfbJvTEXIwNUmNSS9X+ojHaNEN+I
yGFgjlk0GWosjPG1vpX545/GePuXAZ7G9d1tSRd6ja1Q0DzQQ3CKVCClkq0lYBmb
898ueeh0t8F0KfYB+486NM6DrQ9zXIHfNuFJyj2R/A76kLQyuvxsUhBoI8q5upBo
0PDfI4l9NIvCcfPyC7DlmVChlbx+VyVvrjKjCiXO8Jg1CQpsVmGMTChgBseRuhjH
6Ct30+1oML6QYNLlczKKR7SZXdqWcjHGJY30//t0hIUXhWMbg7eJAYlZt7XZGAoF
CtFYA8peFxf9op/Gss/Gai0qrwoiQ31TUtsIgh3MYK8j7kPjhy7ByIe0o4SeTY4R
EHpDWU2hGJEEb1Y/6xlnmyOcTwZjeQuwgUniSnBlDOOFKIbV49QSi72iJfUFdGMY
7uxsvUQ11dPj5BBDcAV3tV0ISo0JOh93cV8lpG7v5SCmvc2xTWJxnDgX4ZUdoanD
b2KPzYApzwiTCjiYYUhgtJth9uVRd7jfyiDLkkBesd3dKDHI63W+xwE/z3yxhdBD
ZpQzZ22GnRavm0FCZQ8+5e0up9tikZ5z0p3Q9jkkRAo5D7i50NfxFmJTAsfYQSZY
F8X+bTBsDz8FUD2PW5eLdA+YaOhaZ3pfqbLuKK+MMNazgl+nVBeEvNR11SqDn3MI
ISge9YvmPkgxiBjtJD3VzV9dw/IeBcXgFI4WntMWZRsagtxb6d+C8zg1+K8iy5Ta
l0eEKQIpKwUuvFkseeZESMlePTnp3undfIxZVErrNRsEEHfLmhLVGJoTsNVilEsD
Cy5PIPgpfbCs1Mc6Zf7UYk8gnbxkjdGKkTNAJGIdr4B3IOPbiea8IxaGmjtrkrgC
lXpc8S3cMFE6WL3+dmtRbbftKqYOeAC5iiXxDubY27pFniPwViP3E7baTg41hnn2
bClKcxkBIe52WDb4k3/FWUlJx9u5dTJhySHwtxi8dhbnVJ3cwHBQOqGv/wxg+tJ4
6oJxt3E6B89uio4RbEYWZ9/UiTtWf2pMdU0P1Xj25Wl4AUzxRA1H6ToBmyvCTtl5
tCKC4nzV4hDbMKsMon+dcwjFRlWs6bs6vta1HxQ3gNQsC0677HTL6sDOG5RtYTvk
0MC9WFhGQ8R5Oc12JLCg1p/6C5JxP4VygCouVIPw+P+AAnuOxnv4PrEVpm15+rU5
SAQSItjvsVq2V1YzZKhbM1UXuiYJmTvb7enLPcjDnzxvVZwO83NguCKL0S4c241S
u8xt588qZVL/bOf2+wY8HwEwxhIRuJmvf1psbvDeAnzeNkw6bdW8ogT27HzeHYU7
2gKj00Bsiw7uag8CR/R290a99npFPXYlePC6kzPSkmjm8JPPIHntpajdNbYtoRTP
Psp8iYB8vtquJCooV+0dYi4g7gfP9+W3sRzfBBukDBYH5sn47zJcBs0fXEBtVKNV
/92Ax5sujTyZvY7QL55w5fYVkg+1NY2jGRW87j9LjbW3MNwGE5oV6NAE54PjOw4+
cSYH+CnC0aYuAmhRho/xSyd3jeltCFcINu1CATYO8xlNoW5blyAHMcngdj9J/jJG
8mK2sVRA5BIJLF9UoE2WM5A3Elir0ojaBqVmj79yBTzPyz0r45OkZVo/weF2FUTo
uaeHMxCK1Lu7eIOHHK6brtHN3npbXrjvmCHjWZuT1vp8xs6/n2DnqSoDaNF6JefO
h1IQPgktUGoQHFy0wsUO+vGM3FgdTwYPQccMQ1KxY+BJasBx4CThfoitefUNLhg1
iTOzbHmcs5Kc3WJFU+PLfTOjmAo8ljLe9evnSU16l70O4myQOoHdbYS8t5vzIAPz
azgv1edSbobEuEtbF3ZTSF2NSL8hQFQLHIdUkTzpgPE/7hsBXwFXTSyGwk5Ghfpp
2bTdfVPISbi1JQayDyoQ/+zm8mRML1xwOxsDIJ34hUrDBNlLUwSXbNOBgyhotlLx
9+z0QAj/6tQt5PuAwUFTMo+1ISYcXMvyjyG79Zu7AWrmjDbmpUKuokyzbkZI4QpI
la7Uo0GN1F5y/WbWA8qbE/7ys47cAs7mZw1rg+Ttxq7HQzl+6XwMudzutIAQJU3t
/e+OS9u0fIehNSyJIyoKI5PXh0N8QpAUBjiU5Jb5FkpePALmxRJY5hMLC2uqTKHf
MzRmTY+iSBhYnD4vgF0TgQCmMqk4vDjMMAMRB0h7Ws/bz08WwCuBiNX4a42TABct
lH4f/RXL6PX8AoL31lCbVL98XkOjEJ9jJUaW2QXu4FO5pYr+ghrSJ5jAurL/DEKJ
BUhxeIiSxVtgtG7rc7NlgSg9crMiJkQo64/ZqHk2eSViITQLaU6rsK0QGV2mer9g
vJhLos/zJdOx6MDnGlhvcoBNPFYOWNkeJlWe6Vek2KLpGqsR1zD6PHw0z79ur2Kj
/TBU90fsvUIxj+jFDM1QVduevtratcUvQXrcPFMlOUC9pBC5mtfQuVzNgk2fjmJp
gUjeXIn5DEXC84EYfxbU5hGwWTDbFzF6WrKlQJjZXFQtU51qzrsKG8DamdBFYEnj
U2Tku8tLOnCU5AXnMAbx8FBrDmhmb+W/bAx70iGcQXll4Jx9tglYAUDpWbUlHmSA
/zNZJ1E5+nJ6P0HttIMNGOJCGTqjZ/aLbmrxXEQbVb4Qr5xrxGBqnFEz7wnzwzZf
sBCiDoJgzA8PjiV/7zjQByQZOr51Pp37aouz/uzfpntsagwthv2WCEQ5v9nig6J8
nxTUCwktXcg635rn/QAE6/BqafNvMM0V7L5ORG28Q2jGF6iMISxGpaV8MTon5XUh
jrUgrmYcLkgnhR5p7pa0Auao1DcDun22RLT5qX2JloUbUFl3kxCJUtnnEy8FF6sX
L9mn6WIlxq2tCaCtxE2M1sjK9LnzXOS2H/lz/QSKpA69UUSRWlSJQYlyD6HZcM4S
vKZqLSWLwJthabl4H3rL/YtYu8eQzi5Uwxcsg96gKUuMQuZ3iL4BnhTQFKIgZets
wp08BmC23ohQNjF7NeuSnIIIzVYJj9wmeu/BgdkWACHG/K3dE/mmzcUYqXZq/tKt
VRvDKVhv2KrAcD4G/jl8GiF7IHLmew9uITJwwo2hHJHccm+hCNDrN4eKMKS/+xLW
PqW2v7WaLSmjPlL7eCdmrgsqsx7aRqQ7O1hdkxW/Ku0oi4+eYUyWkOKt3gCxku69
pOqwxwGvdnFRNv7lwolAnXzFOqKuhmH9j3d/kaDOKu8XRcynFBfeq/ZfjXHnta/o
O/vX32bCSqaiK5Grs2aaC55685vxxvac9Trt7AR0C6QkQMt+niXVqQIs18MwhSZl
W6BOkwgEF53JfLpzg4lJ8rXXtqxr8qvMC4E42X/wXv4JMicCuELDMvE70azBLs2P
EegHLxnivldmqmID0Pc6pZWncJhNs6+H5kOCYQos1Zk740dxukeVd6VZjmzPYK5s
LVhNUG4JGHJRxy/vcdYLZ4V+2YM0HlAAXgL/NHVHRhNCMPz+/UOWTuU7s5yrpbna
+UfuXi5ACTmdFo1g8aRVYvvHntR4B2TqCc5BJNeu7GT+z1+Wd7wNcihO+eb99/TM
tSK3WEfPpRngYdfVeE66DLMnI9Sa96RhtPW5UC3SwXQzzyUgTdvfa0AvmvNoFYvB
7cBTDR7V2UENIMs23uIy4aynoV8k1qfH8684T3HL+C314azipd8vOw4rOD2CJrER
abaNI0poLW6IJzh+KsHjazQUHsm/ZSuwwDnxq7MaAjw78ztl5VAeNPj5VuJ4CPRg
S5YAt4N3hKNCmYt9JktyQIUF40H06cX8r7CGXancJDRpkHqFDtrnYYdRsAWooyBX
kzyVjTp9ji7cX8bii2ixOe1bQfIaQ/1IsYYyJLQ35i4ZyOzL5otAox64I6+JQbIW
KgK+pAhexd+oeB6lxOMtR6NnrA15f/q7MyhcAiOl1p6rwGFgoQ03Hor+qV2sXq6N
VCHckTP9Qse5qWI7geUo3Eu1Kl47eDJ6sK7JxQ5IXDpTFKH++6wb3yNlI3VwA26R
fd0iubxUkB2JySxvb5sG8btFkko9y/EaKjtZt+mb363tjZpy8bb2ru0SJnB86zsx
Vu48TKJ1S8ItT11mg19mcCTKwfqOV/4wiSCUVV4R1Cj8l3yCivHGaASOQuJItbdl
83BZRZJABnWQKJrlDGWrndPBqmpxwZEqpjfKU8oYyePjWo2iv6odZOgrYNEOP/Rd
ev3UvQ8t6SA6RjicudfbjCApSxia4u0IsN+jl0XbgIoW7CGQXDxZwob2fNlGR7OP
27nipw2nC72JQmoHBmG2uf+FS9Z3O9U3KEzIoFV4PBiu687W0f/kFJWMJYfE6Rm8
lxDk4npp3L+fXeU7AQKriOnm9vfyOA88xcWH2U1wcfSTe3G8xVS+MoNKQwqjUHqK
B2Ojp3Z3EeI2FZLg1hIvo7zG8PrfhgXNY0gJXGOa17CDZuS6t5L/tcKnjbXLz7nV
/orWsqDhJIM9LBCdzrZGQYgrQe4oYthfw+Hzubw3WC3CnJetBgbA/88otoG/lrxR
C5CydSQLKwSMTFjYH5KBG5cOUNSppddCtQhHpVUEqQ+nZd7pJesV8XC/SlyOcAZA
FbXBT+W8EjmzXtd6V/WQ4X1CupG+HlmMIht/3rxOvQLT1lWZX66SPVOXSm7TFq3i
+WvKnPhNhdMYZ9dBz9T7ZN1m4OQTnH2RzietF/lRTyDQ1wKMumADLcIodSsoQmSH
hvBXRJLMh6PbOzywLAOxHWIYjcIITkEr94/zSWpEgCkrXH9XBuUjzfhmlxcT57zY
dfsrgIPcylbWpgh7gAAblklBAxFIIrQTqJ0jNvBpSY0OlCBXVVgGIgLIoD9wmAVh
kT6cNP9c62vlYwBBa126D8Oc0UKTI5SqYibNiduQfs7X70flsm7oIBFGe8jlTYp/
m6T3OtWecJ5sEd4bVJo3oYTMOF5B7b4WmbLduSCZCHF4bTE+/c3zHA/3+KBDeLOi
h0Mvz4dM+UJHxUJ488Vtdw/p0+WbITv3917UaN8x1AYUpyIXfoOnx1BtpPJXJaPF
QEDwXLBQR9/7zqTJV8Rhsz0E59UjMwyc1pEUNMFmbflzKq8BbIsch9hKb7j9PZNb
409GpGqjQ7i36Gbpm5uX5UjskT47A5dO5Lpv+vI+fTONE2RqPcZo1QSLe2jatNR/
xWTD7OCUkz8T7Fj+RNf1xeaw6YsCs4cDbwgNnhiVdIRtpIj8ArzS2Xx9eoM7ORFp
EsOl/Qx0sfhqUBpQiDw8iLRcIQS3R+jp3wEpN8xDQvrdaYNwAxKcLMER4rGQfloy
f4hWlzzoQdfyEIOPFDfHAXhgCqsud7QYGIuqdszOctS5JlwDPgrqjFiQnYMRLME8
/vtqU1jdrigGCwOnhKrDsHBbrVxtAg/9lickC6MA8TfIvqID+ptBYY+sLnzqasrN
jy5HfG2sTlmfPoBZ1BaNoNxOl1jImQj8PTPFsfE3b4XRMKJvMHYts7qknZ6sQouZ
dQGqulas9A9sqDHb3Bx3NPyXwD075RihJAGxG1i+gN1EjoCsmGNb3CU6our8WdZU
7AO5qeiIQruqUMTfRyCgleTQvFnCmRmT7j0wIfftOu2ZsS3SXYTBlOkYx05Z0Uao
N0kkAMz5FewsgykX6MyE6MrOfn7lrS3788dzQ9ulWP9zt2xn6hR3YIE5j63cBhDO
74FVhVo/eBCXlO1p29c7TPeTC0/mPDWwzPqihwzYhRSpjS06WVp3K8Hke0x2KSVi
Y1tWZcpUnS7YKBKXDYKRYaJO+DMg75R2/NSX3bS2weJtXWhoeBKWs7X75JuMxVdV
3ESHjXEl/S3/Txn0NezsupxHHsVVRpPYHBzf8zvhIFi98LBH/eVyEhphX/WUcTpD
6+xUnIu9g0Qc7D8L7MuaPVuJ+4kZITSyTe7GjzB2fT6STl0tsXf2aSc+BN5TC6ir
pUNqtapvIbb8kNQJNMSVetau93Uo7RiZldKFeCeHSbUH9s3E8EDO9nUwsEBwvRwd
BG5KEF3ARw9Kaz0fikHH4yMcymSocJNUd3WuQgN6qlAMmqjhsOifgJmldi2LHKhQ
WPDjirjVOYtiLfEE+loZVMEoi0LL7h4B/l5OJQ3lWIQzFG/3Gj0B3x67zwGUiFxz
eOUXFxfsfqkVQvSP7v76uju6zFK+9qQlv3KIdgvZGSjYgSiXlLlicoCN+zX9XeqT
i2Z8lOLEURc5z68/Qd2LFzqqK47C0JegAU4glDkCh+HxSvYwJwB2AXydYxN2LBKx
pVhh2E0K2t0CiSpR0do8TI9r8jczzqLWkJZoaJw1s2B9jeI9+1bRwVgrbAiA5kcP
m5RNS33cX8A6k6GtaQKt97yrtuZXX7XTs8AGSnVCpNReb1Hc3Lzg+BUWwjLLoQQ2
ILXni/leDHMvJRlqhVBPHkqJ5ty5OlTYpt2wEMIMnAUIc4Np/wEUei65yH08CLYP
kVd6rbMwfT/vkF4okithDHCVm7Eq40xAkpuU9dIS2GDJb7jIxAOziYc4lh/iDswJ
grH2OccLm7iv+n1tt/R8geT1A9eKsfBBeKrRUJNk8cyh/KiH8X7oTm68SIfJKZ22
Df8O0FPQrAIyIqlXlcoko0cTfJID9Tg3cnr2Rn9sNKyglUeyBIwJ9qZm4unhqSDp
boh0iDn1YH0tm0+0dsWrLn7g1k8XSTMKANp5vvH94n36ysiJQ9Q/jzJAg/h79pOk
yMW3ePg0CceFloletkU3RYa4IbWlgAkJXMwD5xDu1DZedMv9w79QxRgY0szznqdO
QC2Z8eMbJnoFYLJRLp/juMvgRh+YXCIEmdgwm3iYYyWanFcGH9h9vwpYVZGwZw2u
D02/J1JWnrWLwcpbSuv6OKLCT7fPub+P6WX/FKn8iee5Yx/83g8XwFvPbBzOjy7f
T2fu3Fqt+f52DJzZl2b13oYpvNIVgfjnuRm6viAXUPmI2zCTgZFhF6fEiQm9kV4v
mdUsIe8arLTn8VipRs/HeJBpWpzw9IO543rcOuu6RZQ+PXakPZK2NidrDrlV7Z49
zTiJStJ0KTUvUQivjyhbSxynV90WkqXHILwGm5hBATTo6+F7l0yYVtSV3iRJbtba
YeB4z4Qyl+/GOc/WWJtFbq0Qmwv0Ws/KCLgEY70bRFoFLndLU9O5NDaJT35XODjD
5yd4xGQILT6rvrZtJnClU2ua/4jbOFhOiczVQwwqj9rir+IbRlaw0APX8J3G2WhG
XFpZSme59OQMAxU8Ux6PYjLX0py/3EJQVuxRIEnoY1uh78pA429NIlT8jlqIK3rq
ZUnu36SpKEjAhxqSO/NEW9jCf1N2F+LuOZ3Kj/ndp+adZ8/Z6M+lu/Nk1h/Dp83y
QKZYQQ5I4gRrJwn5R16met3DVVs7+vf3e7Pdn2TG1dnS+2o964L3DdfxN+RcyuT3
Q++dDHZYgMe/4+RQq3hoob8ClYHTWmpcgxdsXAWoKq2HSjEVWVmTu+WNwpcWqP2O
/2T4pg9uXzLPohGOkjagCsCR/9YRTR34k1rj2C4z88Y4KFbGf4Ct4NsVwL8hjFpE
Mw/ysvpF1PaqLiHacmYIhz8jPTmmgP3/DUGjC6ktsHTAf1Wc++LcuZqnr8teCMqb
Qam1X64nPBzThnsP2dYEUdZ/iwdn55iKAbB7SVMm7ON35ldIssvZg3KSsc9so7ZN
z2jbGjIUO17pwSQ7wsZ3WtfMMlH9cJEo7WdjnqjRzkW5Pa4Wbxq8xYHYKVd37Igr
74/z5+sxHCyulguYLs7QBE0JJmcAK1mgl0o+h/2FPTYfH35zqpFA5zfxgsfaRQiL
f4L6o6iZ4fXQbCQnAXztA8d3TlQRUqyG32ZGRshtFpORS0cnkjjTWyn4v7ZJ510B
sAhn9FaM0ldDJxy9stZlL59DIT8KiE6/+NLjWWxg3MYA4TrtJjEYrxeEtvgF9d1L
U5IfShP33ECEEu9L6C9lKUof965f+aqkDxZtVkmULg5k186XLhU8e63GxyCdvEl7
MjLCEdO7iFZeYD8M4moSerCU3Jd7tzRpzUp4i3+j0vZyXwemFNIJ2EHsHsRrsZEU
Gn0jh1evEin183Pr6OYG0rFu31zbfWAn3zDqshujB72tmaR32LUEWfsauNE4rF+A
PZflGXqz/usrllAD3QNSz53+0AxPTwYQ/kY8iG+X3Qiu0XBT/Mbd/4sdm1hD0Nl8
Yy+dmSflS0D1GGT3HMArYauLJDGGvgjG+nPdBXHhUaSDUKriVDATTjhzTqWTXqUM
lPrzvnEgyeTOF0vRsXSSKAdnWsVqR6nFrIXcYikuv0R/M/mHJdDOjrUiYJxfzmnL
yXMCeUTETjPI9HL/MbNvf2IttH5TIAKLmvWgntPOJ2cYPgkRUT0itjnJ3B10tFVa
6drmteAHET2zZYRk539y9+c8wU/s+XzF8zduuL3xm+4ayMq4Pw24kj+/n5WWS6IG
6YPKaknn7Dc4ZRNZtH+nE/mTidIqQViHbiT4WLfdeWF1iy2+6e2dJZSfjtU76nwl
SHHUCCfba6AkXRD4XP6X/ntuU1kftuh1Qb9uPgEy3cCxiYl2tLdB3thWYQ5E7gEi
3lTUiXOzNhMRf+NQjaFbk8aGT4vtDmoZl+eCiGyymJrkzGayrcBZUaajl2173/Na
uLtF8gWFMC+bqGLCDUQZ17jPHf2uvwVangwgjppThZW90uCU87RQ6l8tDxqp4aTK
HQyYVR0xcbbabpwdDqkKMt4Zxa5lWdt/8rlkVshZl40X8Z8HUKl/IHvLwrZbKC0O
Gfwzol4VU5Lh9Ob3ll0GjznxChS0jJYlFbblQs6/AaMfahuMHIewUykKi8oRHYCe
dAi7MSHfFlhYNqZAm7olVrVfTK3e5V15xIeAcQjWOdLq75r5QUfi5e8SFHWCZflW
xjXVMesR/DudHA3UFs9HT9qF9uRNhAQk4LMS1DVWovdktHpDeVsXLoCfol7BqLb1
g5thaU1BMGAkISAW1Buj5+uukDCg5cDLrV0x++f+YnXG+pHLs4DVSffti5mewgMr
+fvGqg0Bye9z3mPg50W6i3QLMyGDSjRwEv+mBrqY9s+/Cus71vdEFCfD+OyDwHzV
Khy0kScshiQqvWylmBr9gr/WQ1ydcB0LJKPBKfquPDll9/M6/Iy7aDeXisx99V89
wXNxDVAeKjH3M/jb5KJxo3aahF3aXXJZBYS3it5AL7NwcovBqjQeeaJxGuW0dMnZ
vcW2nemBQEdaW2yTa9z5wQuj0OyDKFG8zUzzCaeoRlku5bpO782TsR4FKl4dI/hU
Qhcji22MsJHzoeGeA8pLb2UxT2oUutJuyBYKXylrs6gq3ZXhvHrpJdM6U5AxZKxx
FCF8RN4KbPt6CygIRgbYtFLMbXsHbPALsCMevdSZpQucTKOXgMrTxSypiaAX/6oJ
01jGOMazB3X3+WtynEHC4zwTqCPJLQz81kIcIPHqtFtNQxKZ1V5ck1F2gaB/27BW
kmpEvk2/LYeD6NWinZabYulptSE6LCN3oXXyHRTc2x2PNd7cB+rrL0OBESr5h/t7
r8cVa7QsiQV4TZXzscut5utuHJ4v8L4lNcQOaS29H0iT1LDeGLf8TMjFYLW+EMR/
ygR1CcM6QBq7+cFKuAht5a5R4azpMwGz00RJS5bmvpHy2307Uny5ItmHH1/v1/9g
I+rYCNY7863S4GnL/JOxyRFsarUjkFs4IGt69Ajgj5+RglcRJDg8KsIFUIG22sMH
Ik04ITGKQ7JKMujgSgKVUfyf7A7o2Jlqo4AIwrFOF78jSwkhT2zvEzjqSounEKN7
xRUadocigaspNWg3+J9bWr+0ERowQ8Veafeu8kVypbbGA6DdD2AtN4B8dCjT/cZi
h4OY7TaXdPC9flzQ+XuX6wvRPJ8SeeOxx4qdPoZPWqNdnFdL8tLhXAzXD/YM6Iq3
sy+OEQORgEs0L+QQXfHXMydjacv68hgCVR8QFqKm+BpA+ARX5b+kLNSDFc9k5pyF
DkuiZN9TlrPLNYqwYwRs6NJ6J21I0Fp5d8SbrtG0SJOO3ZhcRSkEzqxuyy1v8kRg
srvw2uWprjRzZ31TPB/6jGktpJhV/mRNJvY2xE1793PbGIs8QfSPcjDISBB2mwHH
gTPOxiw0PVnBs5BcGEYerUG5MQ5HLOUVtVT0kYWsHuGvMu8o8uFNNDsiO8Olrnpa
UqoVKJvjPfxOYX8tKDAb4zGIlxWWJ0QBav1DkBdqJxzLU2rUfZVq194FgOOpvuy7
5dqNFXBxshQnwrpA8aHSS7sDq9tBRGN/7cwbcOc1Ma5tZy/uuIyEtppzWFGMlo1G
s9oN1JtPnpXq1jdbeokuW6JYy3SxF6cFloPobGhaTixllzSS4WLwCFLXpus/JFYB
13aVxoRGJWyYUoRikIC/LJ8W1ZL1U7OREigPmIBYDdYKqOYcUrmxCpstJpsHQ/Au
Q2DmxVTcQWCJXTiW3h4LvWsj/Q7WoAZanL3hxtqr7tDtQn607Y5N88RIlgnNtHwr
hZ3+C8AJRs6IQaB/QOEL6nT+YaDgRImr9UIQep4ym9YGjQXdfkSwrCWWPkkSisO3
4Cpi5n9y1OZH2248z6DKZxl7Pcp+HJoQQ3ZS9fjcDLqJ9sRIGcpfAJEH1NSQQ37A
K5GcYdqgcFMUdo+b15XF0su+b48HAite9FoI47WyI/BFt9wxIBxKW2IqALHm63QT
rpjMWw9eL1L7I+5qQBFhzleXi0YpfUQJWaOzAYvtC4cr/NAcukV0wV/qU6noMVOf
sN4/HEMSO7CHJBvhCp0aSrQTxwAG3U0nQw0DXrFPn+doGQIZVHGXfIRnx9zOulgT
a+djsvsFj1djUH1tS20oW2dO//h78JS77iXmFqRFCiNCSoScdhXs3stFPUNSCA3D
esNmPc5SrPsmSyTQdIdcAttw3F4lrcOMuyBCxxbxvQNx6h4ai9qNtMXeJvlQVBoD
e95J0I/LeLED+PaoQcTUNyjcGWASLTddAawoL07wE8f+VbTPs/Pz7/xo3pVOOH9A
3DnYCgJc2PtSH3Gys4VIO0uOiV4MhVKxv43taCBKdUs9OPaDIxGpt8eMkmuBPKi6
oGouSAvfnngsIcCFOuQfN3YPcKaG6A0WO18O4msK7KmYzWUAyZmZk8/AC8oF6Fgp
rSAqtOxqZ0Oml6HVeveMWxf5SdawnDkLBkSicwZqMkV60hJgRfxfqmYja8UgQO1k
0UJM5hJdliMr82sypfv56XRDZMMAQkq/QRDjq02Aiq8PN5qRjUmVjhD4sEVyL/5P
4W5rCRuydr5zXRaw1BHprWyXM3dcnQ+3UU9ke3VrANEn0Eyzz+Xlv/UDU4KpXQFB
5UQkoD1WAUfr8vIinPAtiyX8Z2kADcHujNGlRe/OZmHyW/gBYDxw2UJwUSlpd6i1
X48aCF6QjGxh9CjaaSUeGpkc5g51ybqLT4bMAdW8YYXNlcoaeZ6p2mLTPO1zKmaK
ztN9AuJCLOgCE7ATU6eJyyJQHWx4JEa8Cj4HB4G4mvxkihVYBPTmDy8YEtc4sjUp
P1PM2TBvv1c2vM/f+YxG6nstW6kvqfR0X+ME31yHS1Q39WmmPjr9vsC3ryqaMFe5
kTwMPpRfh0FHaMbCB/tIz70rsemRY2JgAfxflPMqlra7mSllOchMoEoRljjAE4kz
2reC9mage0AqhTzkDXp1K5aniubLCHLhcPESpzEDrsZao/MsRWRyPtC2UFDn+NCt
cq3k9bsaMSAhBxXeNnOA6xDOlIsCQkanB5qb9DdoMPcwVxNOas0xoUDatlMLXEO6
BjqvHf3JoNODqYKsXqepoaj94cE/qH4rramxnXdedE+MdL4dzGwQeEGenAjkKGSS
dJHinF4ns7r/nIz3GeKAZK8M0EVZ5lRuDEUw7b376ol/HfwKNiT8fAl9yhjamWbt
gMLCwkGO2JGuyT/Rm5vV0VwmRaXB3kHN7cbg2AQqTxGKRvWLRuDNA/yaNsBQ71st
C+x4tWqYrvZ++EE0A89vKaobxdUWFGOpRNf74nRedPV0yL97T+W/OefhxUx/AKuN
2VaVzBkce0S/Vh2NY57BwfyElTB6f170zZi8i2a+fM/2MK1/sCsOCBPOFsFNs0Gz
XrN8LeNXpJu2DPDekjnBR7iB4/geFFDgsJtRoO8xdosjds1ipS8Tk2MfP7TGvt1u
jWNIGjiGs3KBAuFZwR4Q5L0mh9T7BXtYz8GylSdslz2tT/LPZEDYe/p+wGBH9ulM
6/lFFMSr5MxDRrbKEQPKy+eMm8Efbn8SY1rH6nNqs4EZ6SBF4ZU/i8q6wXhr84Qc
fDiHJlliioAJZHxc0nFVVLhwQ0iLecnMfwo5PFlPZPN8hXLm750vahVRdBdsaXC2
AhoVH5kVZAxpvB8dpIvW05aISKsl1LfzeXkgFs8tdwma8dU12TNXIA+Ya8Wb9PVm
aEtBL8HfIksDrX/faR8Fq8ZBrCeYUK2DMyM1OmLtGB6ZqFu5YqmGrjgRIPmxFtmF
gE0vKONIgmWP70TUentD1W0WBEEl7cc0vmLqtUmS0So2GfRiFRZHK8M0td+1fo/O
4g9RWNfGtwCFCSwx1yjWmD6dzTzhexZ9CCNYmC7sExFVU3g4gy0ZrhiCdBKbNHPs
tisFf0TmDngbEdBzAODkM3dzCnHmou46Zp/Gptg2oTNkfSRB3lwmc99sFVnUSkMZ
mKHrvJP9nkja4iHeNY5xJpdvB5/GhNT/BsfzSZrfJKrVbeKnzZL4X3cHeaMVpAQZ
XRUmBLIBaXMh7frwbfWPUwWrlwdtqSbEHeX8uD8F270+BF2GBjYF2fnempCVFAuF
SHE2RCJYWPRYTSoL8qW12R23a2EqgxXLuqrwpj9KMXEn8TuNpGl8+WlRKw2AInEM
D4He7/3N2KpYk4mOjZYpHLroY4ZkL3t+UflUR+WCLMp84msuxVpiqG0Lbvpjhc3v
fqtz7ANUrNA/O7FhZdYQr905Lvj5LgVcuPoxHOh7qp/9ZK9D1cW36bqbGe3FE7/G
Eqyktx/lySfHOhwAXOdH2AUMJSV5OyBXZuFpD6PqllyeVDhZX6TM9Q0S29wFBVHr
DTxDLkRJGo43Q+nyVnSJRHQ9PcdWhhACiHltFCbSWQKOblpaE7eXWs9i3dVhXwXW
dUdUoX00tRKhq2hsiOD2g7Uo6+G3QqiYGX5PlUM86PLMUA2bFjQMn4TbdN1XCaE/
8eC3yeAp2r2y5wUUjlEklvf2CGi4BenZ+dokit1SWyQRVBgb+5MWuNn5fkGLjfgg
B4JqWQoeEsTvq+6RAXEutlGotya55kRecYe6N//HdobRE+OY6ulEbmYrNTKIaSX1
jxt93fI0WZ5PZ0bwsSVpKcIrq0QqJNpjgO4PJfYwUvvkSaKGuWP+7YYicWBLcUdQ
hUdpxwV8chOvg7bRP3NJ7etPEkCtpLvhazx4r5WiOw4XC9H9dDNxELUgmnEECJon
AYE57TAB+K317yhHvmOPX0peBikb96/tDRACw0sTlUGROd8QApH1s7b9Yb0LfF8Y
u/csTA4IIAkIKuhUU9u7BJwZ1Z4MFBbUoBOFGoNr2h1p4KlhJrY+gp1sjdQBn+bA
TbpsnX3WRVrWpwz8NaDojiYFWWmpJPbkY2poGhzv86ryRBV/TPsIhUjM7uqg7jt4
uhylE0l8lZtLnW7qKMuN5n7IehNEIxh7B3VlLZzE5Q0Kt1dBfsyD7yrhzUz4XQ5Q
wVAPlD9+NJbXx4OHjHnOsl8mEZ3w5ha9028lp7WuxPtRELoXBMPBW1/w28kQHQ0E
b+qllQ5V5l8+aHeJMQI98LETWyOj8RnlkQLe2pAIcSDfpDtZ4jQ4nBBtT+dXYQgG
u8FwcDtYvi7oPi+b5iRPoqQOriT2gxLoU/7pFNaGJJIREAlfTsYMw3KIw7YNrfMy
1d18SPDJ2I/DixwEzaxAgITHyiRux4dVZ00t9eb4KQykYPhi79XnXNbJqMYvPmm0
6hAtdq3E8R40oQ6jn/kX6ug3Utc3iDnw5xPmzK31Q83FMGQA8qTgohNgRKlOPncB
ARS2TsAveX0QSNpTDwpX7ZClr3PqZ4w4gZLF5Ox3FFbNlPdBZ44cgZsCVEWUZmM4
eVgu7xKLl56B4DrzV2jJMm2elkCtjjz3mzKLvuCO2OGeHAJcpdjUdcrYIWXL65zG
QcDca+fEX78XuwgpBEs7pvCYEFJ7M0sTKk3loBiMK3kxqayOc9vZwOdRyK2pI+rC
n0ZfAZCvYW6j2PljKe6M5MyclGXFqndhHFl1aoIVFxw1LIpv8hxNZzwuKe4HAlBn
oZb6wIBHpsSao2iqJf1B/0haahPV0sc5ZHzZMF43XB45AbABaxL6Dqv8aWy7Wa/9
0rO3myDhJgIY3KArd6FvLddMZ+4/PKoiX5I1du/8fTT8I1hNxctH10DF55Bv3UcR
WzoKdUUmdRD2ok3Eeouteg66TZ2na4VSydMiJs93NpnrVjxd+FE7onEXuDwIJgKL
lGmbHZ+VWlEaukNOJrWnaH4uFnqxczIooYTzgPsjGUDFlw4w5Z7Ql+rFIeJnWwPS
Sk7fHcbV3vm1IRSEtsx+JeLCD6MflGB+pmTAoC7+RgrlgMBMKhHnbRmtBYT1aNXO
qQgT8W/U/yt8Zd9/oBIBdTRoUEcQFuisao968JFIucCkLsEdViKjL0427yYePLAy
qBsuF3Jvw8BvkLpWz/BkAv5GqYXgOlSOgP95YMk92zZa3uYyjK9cba1moncE/jsU
HxO9yAsemlHdVgwVQ5VdqVtzpdrPBLREEOn89HscoF0vBgu7pM4A4cUV9PXajwQm
WWX0LPPJi6CF32r2a5X63Ts+y2OgIfMGGQkDwswVskHHrF+qeQnKpZmw9LPGMNF1
Wlnl/sJDoOy+iV4GA+VsrMKVOR45nP5RoeCE8wnVLIfBE0MuUcwyRvobg6mwqpsY
nj8TFqzsQga2CyOIaVzQXXfQ4CpsEi/yToNcLUrfCA4stoknp74dVQpoyrfJLy5A
K71gwuespMCyvlR0VcyOm9nMzbRLhDh/4GH3p+4mm6ySHLv6kTibdh/vA3iSIxf/
OR1x2xyfomJpJ8j186teFtuZbzZ86BLjdDxunYWRPMjvW8WltcQDlASsUum5oR0z
+RnOA/NUts1jII2TEixVuspANgy+oB13QUShobbCTe/HNK0cuCUZGu9OWe6BloPU
0OaRnmQufonkn39jUdacOz1QtQ1KS/yr4OaDbytya9092t54w8krUEbiMlZF41/r
2znfBNFfGmdH1x5c5wIPrmAhiXtLktOhznWSWwfkgkt4fzfJiRzMQcLWYrRNiOJF
lGmen7/Q6KZDpeWTqhY4LStq0FY3LyiTOZz1TOO8PakqjZ11NBDIWks13vvg9214
dY1V9bu+EdKARmjFF6NvPSbj5xwxI2L9xER/lkEDL1wmmKla4K1v4+sbgXW5xtXT
FmrVFZbiKIUaq8Q1ltaIGdg4c7vpnI4mluCDk1eTjslRod2gUCcb+e6Fsci7ayJH
1vVeWmfXvwUwC42KBJKAJipQvEVTXXqGKvzPENuwzUhEqj0KFm50Hw/8wy/Ognh6
v/I6j/jMG3AOU9vvAR4M3bNWVr8VMo1gVvcx3IoU6nOTtdKzdkfSHdBh+ikpsZQN
/6uUPwCOMENhEjeMi134JHvc0eRKhGzUI6f3+VB/+2ca/eIzCTmKuowASyho/P06
KUtuXoW2Ww+BtOpiN5ca8LKc2naG+b0uuSwPqGJxPPI7qBtb2DUgdeNPZvWy3Gz9
J/7mqTTJofR2ya3+7jRXORccUJE7JjP8TM/ruAORY/p0VB2lskj+Gs2SgSfPKJkh
u24RtUQarxcvFbg+zevNID7sxLeCKosvbyiJ6wJd5QQfTlrtmlFIR/WKOqkV2BgG
HC3//8aFJesilz0bZqrCXKU5o58doMlLmKfR7Lk8tgZteRha4qNVR2pL2dVkl2Ol
tPm7mI/37s9VA0mWS25poDmzIDd7Xfz88+bWCWxCiC2U20JOzWBek5ODqvOz/AMs
nTUaLRS/ntmON6K5iiwhVS4GwH4JOyunNzqfPv1GV12RTcH/3oVV0OkOwh8Ee1Sv
2R+k6QFYdA8omC80XveZI7cC+Iew8JM8Evbz4aTbee1HP1fSewKoN4W9uPpnCBTM
d8hzUOHpBBHCxCyaPtJDW/78HXLvyLETGj381Swy+sq4j43hvi+JbqEhjC7NdEXd
BTgwGybGNQyqMev8Hvse6dlQiqYUWvwbP7W28Kcg4QUAwZVLUe3x+FcanV9AlEJ3
sfJbsuXP7If1H9tVQfvyERC0v1nSFmVrTYIxJnGlVpis9fsMLpL03xFdSOrfB3FX
xbDZ5LpuddeCuwJQgC6hdKZhrGjmS55YVFgANteFULVUumNFClffAfr5fZiVjlGu
DGu9Zs9JMJRSLeYGAmoy5ca444aNwGqWlfthY+OpVTSTQMrC1HAnYVmI9uqtz0Jl
ysrjBiLXWdwG7eYYFCcckI5A7ZXUB69CC68av9pdnv6I1GlPUFMp1k95PeN0NeCK
nJ1y7b4aocbzMnKeIrDwhhqxrwPqHHP63/D/TctXuSn4zt+zCxqcRvnOKRVXSbZA
RZT41VkHIM/0WLrRJqABINA7qQGrDlCJl2HSOVXH+F+0FWo2IF6ozQflV19cYTMC
LNNQ16yGzq7OZVDFXu7vI8w/HYVZDPcqh3UAJnaDjaeN2uiuaZHYS1l9SlgChFoC
VqBKYsnj4uTnjQUeHrJ8qb6Iq43CrwZ+4pINOl9rJoJBZwh+8/+EUmM1zn6fEWux
QDD58Hfquqvk177xRvEp+jENGjeoV0SxAy70U3mruZvuxdoQweHTJtAy+3WagPte
UFo5G3SMFxMybzmYRU6tFlI1CLDg9MNAh0y5tJFfhptJjcAVNYTbnzCObw6maoB/
vaJLA6kVCsP66z0uvUEASShC01nFSuOHe308k/4EL7fntYTiG6MliQnOup0cnd1h
1xOu1ewZfTxb7S7p3t+FetPuaptbrAp4DTuUq/JMtixtGJFM6GLkfsBjc5shwfWm
duUyMQ8CdWcCd4RFdYf24KK8YSuVcrhx9FP+t1wvCjpNcryhnIWem9wANGIpa74C
1HlngihcNSaw7Wf9L3CVmdyg4duMLu77/RnY+Y4d2omCkmb1Hk8sD6ay5c0HlUeK
6/SRvsveMPJfYlrTkWqOQAzCG+ljNeSMF/KAAz0hvSeFvhXmBwqWHAvYbXk5Rl+j
xR1zn87nh4lbfKT4iMdsFKjeVL1brSvtsW5RrchwL0LzaqkwE74U3KXIBlrSTrQD
OtS3OPZ2rJH42aPbM2a42j/GlPlv1g7O7fwr4Vnq1X8uOkVFeKU18a137oMCVJEM
VNG2QjGyTYHQXWRSx1J+SfucgPGgEIdpo6a9lARPg/wDySynCw0sGdXTBD2mi8Pg
qTpGcoU+WZHe+2h7LB4+dH8nhhgsGeEyo/sCEbttGz0PDj8foA/vapeRdXlN3TPU
rI6NZJ4UVAeni31JP/lY+QcguKMasr2PMAxwOltt/w0wUoFYQoddtw9s8m4H8L3Z
vgc5JEYGxVeUSG6ufCVly7RKtYhmGkxHzn6Jx5QAEn+QZljLaajrj4xpZWevm+ap
kFj6Yvsl2WGyJsa95X4SjxadlfGhRmiDK7ZxNk5MvaRD4KEUAXvTncLpCn3rSotg
DJp/De19/vQgkkoiJCE5Gv/dOS5jx1dZWGGuO8LBDvXPJhpA6nWcl77krojywnQd
5EfYTBzUwp+vJIb1u1d9oyChycOHQa4nYGtOO+9XDW1p9jj49w1/qi1tgPpSq/zx
2T2jXh6R/o4buYDs+A2x0Iu9betSWVWAthOXgGpweYvrHG3Cj7lsijEWZods2evZ
CP8bWhy4yqRN/NqwmqyaorA11yfc5do3enmjFxi4+HxxkujTIGQuvEAWwgJEqMPU
ocE900gbDTObfBymLfsMwHVugCxb2ulKgeu2lq2kHR2OaqIEYTTOvtblPHz+gUt9
yM1U/e98lDcSfKaPzRdEKK8niMDZAJ5Lbqwx2zlcM3cm6qJd8qK779nZZUxUBZsk
P/Oit/K2jcv5Zq+i8D9wkBksVL5tmaF9Seortd6a/jhxnJYu9UNDGdx6AepZazZk
H/egy9YF25PxajNu/vnHZY09hua3122xasY49fxpEB1ccPUrYWYiLWhRnHoMxzj4
uYloswf1IPHIXkjHHhkpIBzPxlGooSbMsMFnT8ki9PBUNTHmtzX1Oas+5EuF5YRW
4KeZ8cCl4Ja2r/kubh7O5iaZp32zO3s44xV+ZD59lVoiEOzYSb/ciH6Qcv5olgFF
no4EVgT7nst9lidmCtEn57fk5bmzF9ATFeYid9Y4msznYtbn9HpPRZiDQJSOGj24
hLzjS0Ga0Uw+7H10VjU212cPsTvbP10VQQfrbTx0DM0vEwvoJsHYEbRoZnEwL2ks
RrAm1p/udWXG1CSrRUPu9yUSCs8QlCzmY/nKBuyV7dxvIHRMOg7RjHMHG1r0f0HE
/fy7dleNQ2PgVUMJkZLBkn5nXa8FVRLZXztk7eN8MPAXi0pyf9GxBFoQKG9jIXRM
feJWHg+PWLjGY1ApwJKCsYhrJdHb3CVS8Q5rX/qdO4b1M9qYY4jPAjn896UPqkKU
/Az2cCd+t1Bw2qFkkaZqPbbgDaCD4eP6SElzVOLqsU0cDyXsQO118MD1gtG9LrB7
Wt6Gr347C7nuDuaQzoNVyivfDotAthifTJDEpE0zbEW4tSTfeweRdMt4Lfk7jCUy
Hc+lsA741nYzA1qV248/1YS4BP6jqhatqTjyD285Z1pgK+PUKU2bQ07E8H81ezah
QscSmVu19Mo0OQ0QLHjKm/lm/CmND7EDx2Cw6RvQ5pNChi6UVIyLj4ELpmYvDiRG
LPnO14jYL7BYL5BVVfdmU221Md6n46UWawZK8yhWU4oGuvNssnLs/DyO4JK+UjwR
I3gVxbg1ak9vJa1uAyiYG3Bkx15zeWEDA5DqT7FaLiCNVVyFnbw0x/pb55pFD81r
8KRGUO5KjJV0YdwAwtuLVDBsNjS5COLZkDmDddg7oLrau0Ig0N6jTYy1KPTQCUMh
6rlQPj1iG69VpGx+s15Qthe6stO/omqvAoM0zlq+FZOrc7AZFhw501KDNAoejEy6
NTJ1B3LAAx7prV4Ix0EYApu1QtUYYj/odJbP0iQrydmCvKmNrimC56WpiBEdm45/
VvyrgMJjGLYGBaIn7NZ0rbTNsukI/EX0fqoNuSwZ4N2iX7ecqb9jmVpcqVFXn6v4
57SlupAqM8A0ZSk2WA1XJrHzeFdImA6FX6D72bSPIKudeOdgE/OJx6Ll3OgJCnC5
SmGpA1yCSMb8TZiB4vnqZjEjguhyI0MPI7g+/xd+t5tnI1ilYDk4dTQTMTaPLyts
PH6d+IcaUmYLquZHlf2qHPkzSU87zEyzkY+KbTdPiGblckx755YZu26G9Z86+ufq
vht5cFLT2hmZXytX5nYbzYW+T9VpI/v65E5sItoxC9HlLoF//s+5znU4FyCLoMgQ
sPcdcrQXjQJE0z8XgqpH2yWEzvN8T8FxxO0ngJOrN9v1bFh1+AcHkoq9VgJtzQdA
3p9dO+DLMX5/vX39HstLl+0+S/ZOYcthSl1m25VVjw/SGi7fIMxRcr4NySjEZYro
s/2sOM7u6lBZUNK/C3qHVd7+q3i9bAdrv2xYbHGs0AiZuVfQq8f0KUY/dz2CuqAo
ku+Jzdp6r4+VIHKJSeburugx2p6Gme9KDaEIomKeouicAOeMdP0ElFRLYJ+WNQoS
Z/NotA1aVJCOCkBLENRTnTt7ijgHhe/lO9eQb0+1Ssg40N5pngS6XQpWvPCgbMtj
dGrXK8QcCADjrP2foHexJPr46ZWDI/62pLMlsUDM+Oh1qbsj0juA0ucaZwu05fbY
RN+abqh72TNbbAJVZ0/fZp/kDUXwqM/Dw4U30Dpw3bpzdbzSiwdV/IS3iUmRB0zi
AV9nDrP31Jx0SEJvSachC/OzY9mm/a7xMY7EdqLgvjWTdA2dX7KlfGns4hrXsaEw
58/MdYyT/nbtAI0Y5xI16ZOBoel3CysKCsoZqjBalRg2o1vTd+Rb00mc7bxaJqEY
6TxrB4dJcfuG4kxxCAPifbC9iDIomjn//3IoiVwbAhkNifMkLTc7tahtqhh4y6+O
a8d5Y7G9nGMQqtPklhCALcW7dWa/yQtKBZVweHEADDKqzTDNNBkNWFTpXHXfWn7n
pqH2D5xeOHaeNXw2wEClX6q5mUe1rnMtQEgf7TpoPZhmuHKw+Mi8ynKFn4/VfDpq
0qS5RP39esMdHNScJI5ZgrjxGQMzo/4ylocVf6I2dnPaeUfAMuIZpOHWt5i6yykX
DYN1KiPW2yzPQsmut3Hx2iD2tzb68cwynq+AUHIRhsWQNuuPx0yKaWnkReKOc6Dw
InvzltgI9lmPE1Pjt8EwL7gwXWULPggbr+p/kmRJ2GX7pfaXUgy1HYZZd+QG3ooz
BqNZWNkFkpT1/XcC+g1U9UM5uZbnJGIe9Ux3ihgiVyWj11clq9HXJpq4B4NPvagc
Fu/Rux36hJ5hWLwepAmQS8V+ysu5zuWe3QBqfuuBIXnbOD9mIWfmZxCG+UnUkRj/
lF4/9HZ7YKD8VvfgWdGShI/EcB6WrPcM29+yGSn5gNM1L0vYgMTWiVZ416/fAs3U
6cwnVCRRaNiBRhnTpcbNCYKws9duOEaxOMmHWchurO9+R1WV/9Yh3aBOKPhHLlTq
7WHj3SzxfuhWbv8vmxAuZhFCdRKRTCF30nHcZhql7ZuUwDxYOW1ZFf4vnR4nLt0t
yeoB9MQooC0SSVT3QHU6Ayb73arXGGDot/i6dhkL9fDIiMNKWcjoqIFuT1N9xr4s
davdLjC0NiFWOw7spyOBNT6nxyNukqNEWVQuEToscbgt5YO8kFckhlSPjV65LefR
d5h7khQ+GCShGkSTktlCkYw7nwdk8j54ITWk0Dg7gQeZxzBqvlRW/29dSp8+xzU9
myuI4RRm7IJgoi93gszymrK2ccBx+dZDvUXWlYYIRnVh8YoEMIqzKVRip7H0Q3dn
U0cULgPvWuwIZJNG62VhLSOqKl+ujoaO0XF5P6nIGu1wWB65E5gmCpF7zLVfWrgf
RAEHqcvlMdysAkJA8j25qcqLlXT7aGgqsWWHfXr0hb11GsVfhJtlchiIbq8w0da6
R74LZhnF+ziMcKpKSW70Wr5kOJqurfS4Q2ZGMyTVpkjBzAC3GwQMRh5G5Gj7neqS
QZ5QfIaCPmFQWGcTKG9xYsZGEUGXYX2OJkco/SGfHyolq5hVbvmYxAhyskR8B9ps
NYOdCgiYwrF/N7QksbWVcscoPBJcBrlW4kY7qXZByshW9fzTer+1WwmEoBn6CSYW
ab9fh/sn0jW7Q889CN2j/R7DwHkt8VjTI2F9LORBYIJaIZYj4cfVLb9Z7UB37/6h
zGS3BSiHzl2Tlmtxxm+sasafDc9/aRCu0haSqG2N4V5xrDEJYoFvVxMsKnWm2NWU
tZZyHxxRi/s2NhTWN9etEeUiaATWQfPhGNVq1bCnUaQC4rUMbymIVoOqv8YVSsZm
C5Vx8gBbQ7PJ7LjjWDAsfcTLG2RXoZzylT7eExCJKFV11gKzNSnS1iEMHZAkGoYu
VPGl2rOdoZIiBEGlKKuzvXcnYr9OiCSTM4XG251bk9BciAN2tAjY2S3Kgq2qcqTK
pWi1vO2A/xtd9iavEDjHxYIZ+zXfLtwb6oHt27GNdDRspaCg6Fg8PndTne7697l0
6PLv6QZAf9fHuHOqHSbjxaoYEiIVA23bkASxfpgg7jjw08eNAUgVqB4KInT5rl+J
XtLXUYHEMeGhtGUKipRxRGRpNXbdAXiQOBXWPgIMbrJB+3/tRzIMfcC6ux+8eKHn
TTUlEccTbLM+SQQfYt5q72w9euQ5gVNMwpHYWV+A9zbiOUoAyZCAPynxs8z0zUZw
aFAmzLMzorvnGIm2BOegzQOqba9x301ABekMKfhwYHMB24orqhp7ST32D8doRpOc
xUsPMlvAfPhDvfOqEFVuslrYPXYYSGBD6j5jmYs2ELbCWkZgcsR4F9FrB9WF6xgf
r/i94WaarVXsHsi4OcIuGld7I+YxkTnZbX8/yTqSpbxznqPIjRuZklxKs06DnSYR
ofuiqUKmtzqEIB1x1ltwQFnioi4v3RJxg7cabRK3cC1Q+wy3EJrk0ruuYyfwuZ3G
6URBq1jFGGx+mrmNLGhOEC/X07m9RSqlpk2aAJmGOpWeQ9rIsp1oMtB/oWrVxULs
g8+LPGALR0FmYciZiXhrtaN9E0zmUd6qbOCAPf5iyraW+xE8MPwcCwb1x9vpzBR8
vssXMtDqHHPuArUx0S+YxuIOG4QPTwQUJlNqmJ0yvMAu18UNEfzLRulPzES/GbZQ
QHW6aDSVpeMC+cminIkfMKxT2mJR7xV0FwCWdegQyWgDDpPlwTchKHAwk/2tFEZz
yr/itpZXuaCE3gfMQoSDQ9WQmzvj7CoQFOncpikNycWYVhJlJvuC5NkhyszafrxB
3lgLOFh4qSEWN8s17+XVoxZfj/67sjuuL2Pi161ol0k+MG+6KwckbwnoK1LA8dLY
nVk5Q7S6CKxx+xBy9pHOvHcwdkgaZWY5OvViUA1n22Vxi/IUbTsxLOIkpmAQ2bOi
V2xEX+TM8VNHs2EiyD94kcK/iqDpvj0Y1UDSeeF6qC1iZogI2UkDhy1lP2HlGRLC
b132eQlA6H5/SbCmCcsCu3Mt6DK54TyDQGHHHazMU5z+HA3jya0SMYnJgv+QnciT
Q/qQBaFCagbnSCm0w9uxAURhwmI4QqkJbgMOojFXZECAYNgXuKOZEG6ZjRVu8kZ1
8NSPLneheQcJfomCjJlnRVgwHoHLdSleLHr+463wxbU2vziOy8EpNso6mJ3FWh3U
6AaRlCgvZOAadN9FzG6ju/ULuv3jq59pGr583xlXFs18vxtvnhjFeMYE9O5zWnP9
kyymLWcj84Y657/Qjir87tdGgovInu7YtUJqvMsUC+oLxgaRsbl4+lNGOhn+wYwX
q8lxdUrI689WYfIRRFsz+WpHJAS6625LtYpJFhkhFRlkLnFMcHv1NCI7Dbdp0EL7
JX//OaMcEnzrY4pWZFqhMxjennxIMyJVyDcX0LF3WsDXOGffL22mLxl4g+z8pZzm
D9ONeaSINSRQp9s5q4L2pj1tHYoUKJXAXLoPVmj/MHB/jC7GzAf/DJ/3AOF3IVu7
L1Jox7MRfZnsXbXyX6Kt37wHLiW5xGjnuTuu9d+SH+4kSe1RR8/qJGrtUz0T4BrJ
klpr+cCPi0o5vrBk6qvnHF+lmIlTvrWybxRfpEo681k3uhMnb62BWb+Ze5h1mq0V
O4ySNxo9D6Kbq0Kuj0vMhnLzNyD1xwRX7HcMBvfOnYVocFrDTK+HbqnVNau1QGii
nqYr50NaCxTB+SMKxaarvAxb5DlfhJQUcwT0BHp9VOxEJD/XmeSqtBJG0zWEVVad
eG88Wecf8NDPewAm5kfBoZDMhgHqZjlnfiSDaaW+M/C8759FqMM79Ol/6t2gMm3P
qGrkDA3FZUmr/K0ZiKd36fbfcA5TLmG30nk4fddXLUV12KrqRNI6hOy2U4sfkuj9
GMNEPOP7EbhTiRJ7KiRvCEl78ovfgjeIpreApNYrfKAGCYTHgUQCWRP/svyZ39B0
ca57cWTI2cRcWejUQyg99GZKh5PRQOcgfJroDB4uvYNWjIhRCnW9IJgALl12Kx82
pMEze5aO/DA+hh2NEZwepgJaiXABwa38NxvG3rfjsuGiUAV/0NOHS92L/nC8HUwB
sdjEEdVB7vPmXzh5IsZULoAURO0sN/gw9Du/QfyXR2cYdUHeDGSVD+i49BUSV50B
22PBdvTCQsompmOnxB0BV6Jh9EuN1QWc+u7IaaaeaNfVrCGgTxPPho90mMzC7tA9
LUHTlnFJYGCoofFTKoNgxfznXmtp367A8o3HKWwCBmOLBE0hW41jPI3q+gSm83gB
QvAYyEt/5vrHYZ8lomtKFm1rfQY32cy0MiDvWw5IV7Iq1ousAhZga6YfUzVmDJjn
tmT/WSRZ7kvC9gJqtxCkdfTlzsivQPeiLnKRVJec/Uy0UWwyMZVBtCiBJBvgVcaj
2ZS0TWsx5mym2s5elLYp1WbAMexnekdxmyJXolSv2LDwcI0cBnVe6LORCDVXNjSd
Kuc2JK2kwZFCn6IXDMUbkmGYfnYlVmBzWYTT/2pGYIno+Tntci9NjxFWrzd1yG6q
L7jc1Pxcyk+j7oXS+XA+y63A4a8W41cyU7hedhxkI/comvDYmzy7h5X6d+ZUoFHD
TfKlHjyDTju18JI+4XN4K427wFAKPKgMyn/20zesM2nHz06kVPKs4vFVyJSHt9rc
wGLkd+68mvpEX+ey1z+sqyX66SxEKwpaVhYUsI9u7jkIOt9fWo8WOJo+EpdXek2Z
n6JeYcvIaSZHaUOG7uw4Gshzv0VjMfvZEVbnCt5/Pny7poA773YOH7wxkBZFIKyW
CZW9ZxLu4lenAO29MkoayjcMQzNORIQFukJjPb6/g75yP5S0tRsyQnwVUn94vwOB
v2iGJ3kcvzubTT9jatXKiRoeR49vAa6Tllz27xGzufuu2UW51aQpOFuVJU53p9XT
4UQ7MTKxXGEnwjqoz50azR3wulpiXDn526wPkUtG4UVpCK5VrL27WoSaWncZTsIH
zyxyMklNX+f8nIvs/mQQaah3A4wd020bRO9gJ99qo66frJlVV+ANxLYct12R2dlD
CelIUKoECgZBF7OpT9aRJZFF3REQOnz2ZDXd5BFpMMwI/ITYRApTFXQa6MRI+jdr
xk9xELysZiktK47/CtzssVniSc4tf/u/VWuoG7nzcNm5Cd40w2FJgWmvJETT+DXc
wkNoLW6X1N+hmw1U9WIST4yfg7DIYO6CsnzX5QTWsMAnf3d8eOr2LFiQqNaEIx2j
hk2ffysn3PKOOPwLxT/g0w01dIqQKpjRSgNueNc5Rbz14mUOCvufhbCpZMkOI+yB
w9FnBr1hDNtxP+46iNfpnMBpabpSgc366kERww4qmSd7DgIap53ZeHwOghgQDBAM
sU8f84fpXPBWV9F3uoBxNn4Uy9wsUG4oGlaZ8+kz+4RnEYsN/Vgbe6/3SSbOFkv4
MNJ2vrBF0Y7/Sk2XFgrP+V+MUDA0gFu7LsfN7+A+g8GFWCj/Ve99ukggPCZJgH6Z
miLAqrunDmcVypHq+LWO/jyXKZ5qyBr5XA7RZ/36PpkJAoPyEh4/nsdhFyYVBgXZ
OHCAjauH8cCpJJE++oaMAWFBcY/IJ13McPNm/FgexBSs6ZI1VcTm0boYU9ZZZJxu
pBc66kdvVPq7JTeHH0aWeixDckQKA3AasKZovILhvwnVu70YbDUR5TThaHgXbxxx
2Dwx2C79w3H+HkOjHlj9USn/lVQjY9cuIjHo2HVJT3YYTxlKPbj8/UUyVOQn4zZ6
mZ0fZMnMlp4X7oa4p4RArqS0CaD+BKtgMvY6ltpadxi/c+4ZJAbtD77Du1sQ4F1U
JGQcdORckjgDlB8oB6JFnGOjZNAGDdl/3AGrSrAE1Z9983e3MMrERNJQc0sqkIoL
pxJ8wsNIXJ4fbH6hFjLf9Q8JoJ1NOiXoySXphCllIdQfomBec/yR2iIyaZHogGSe
9jrBLxRp8iL/1PfGrMso4dFnunuMexZ98arRiQOaq1DCBPiwyTP5jzCJxATYT5LP
asQt5GchpiZ7y3yuxH8VDSmLpytO2u8yl/lq7BcrxQAmYEcS46d4Oata4/SvP23H
+Zlur6MLpNBLkPhRS7xf2HF7iggZ92BUiN4+k+dnPrC4S7AAmNyPRI9wcaaHzVXK
Kg80WsArjVhy/n+MkUS2NWiR6G3dGrwvTDZ6WJRzQr8LSOvkkVtkhE9Y/y4yA+2N
qz/t1pwsUkpcUPc0bFW7n6W/fEDHBYajDt7e5kANPo0qRVc1D7dtDZqdRsy3Roc6
28egqde2WhFrvTLDKsQ9b36bV4hNDp++uqiY2VNpwHSGoXmHeAonL0do+pZN6uCU
ZfnX1Nl6x7K6F+GmVBQxhCUMlnY0TYnwQM40jq1Hp2+WW1XChn8UQkg5+dHhRPbb
SNxtXXgKK1+yDTUkaiM0I9AKQ9KPrhc6FThJxHDTcReL/Dc1qhVgWpLL86g+p5PH
BVqgGFROCqLHgnArnyFOIKodqBYa/wJM9/5O9yGyTw9yHeGyLRx/EKvZQC1uX/W8
IDg5VnuHWYZ5fbCEebKlILKgdZowLAcXrxhZqaLO+1cU/BvznFcDWNNJ8Qs5VO54
Gyk1rLnxFDHeW9DHjcWcVfFeywe4btTowK54QQ4ybi28zttW/A6hajPReaa04HH/
BiVg8x+q3E94ChwNFjYcGQXPTXhhSDAn4pQZGMVyJd1y0fyOGrrJk/N/3rBjSSZs
4q7JCEzlSlYPybg9+rBMq/hBsajEdfzJkXFVGCazXtBf+8hE9dZLqXNgOFB9j5Ag
u1BFtQUkd0xWhJ5Tb98Jggvf0MYWvbaT8M43ZuIpu8sgdyNlAHRh91kfmSoCexre
t3EGySlgAMzfr9Ww6zI1y9gKlRuq2SAHVg32qIeIYsZ1M/v1egFbnm7oc9besoAP
CMwYH74XYtK//v+++unOdrfy+z+dMWB5PKGUi3J1rA66Xl83LtixnrjhiNrf3hGT
DavBlAOazYENkHHvf9sN275tSWX3GiQH/+imK9VKi5h6b3MPQIeWmuMEpAz1Gm9L
rKOg6DVVFhudXl3epXQSi5U7/La35J6HNQNOXmN4W7WxUB4rHRyU2+a2xvtOydtx
PcOZ7oMw5G6oLXQ5yzJr1fcX1DDj4RFM/XxutLQtWohl/w8daqtYSdEPUzSCZJeS
a6lkKB1YRRtzJCXpZnkOYZUMAp6ORbZHjMxBRtk9Lk3WVb8HSzubK17II+G8KY3A
lBAQDMaPnCDwBVXMPwZYHwdOmjgnYL2uTYGxvOWpxzvGQPe4FJkJhZ9p6OMENy8P
O/LnzUM1LlmbxyD6QYvdVCBoIjeoxL768R0bHVSz0zfViOtEWmbi7QoA7SlMHiJ6
je0TiraxLfCQxykwU0rs0R/VZcNNwa3sgvCb28ETjeu6i0yxA5nwAGw/Owi3Xnjf
z48rhIzXbfB2K0aPPZF2rkgICGqeFbLrbKAGXZ5k4VPgzSuntY+8llzGtsxz9FUE
2SuFFx3bC12dlqswks1OLJN+ODXzKGyFe0pgn+gxJlZH47D4n2qRm/2qteB91caa
eU4lOh7MlrxXt/NP3BsZXZOD/M+YSDf2LpbbpR3u0BbTfolIYELAE8U+vf/Jgn2S
0gyOlejFNJerZZc/gNC6Gn/BzyTeGze35VRTGsLr0mLDH/ivPOh7Q/L1uK1NQp7I
Wl+xe3+kYFvXp6Y60VhgF18S32CcEV0qM0sr5WHVNl7JMkZw8IvVF7EtDQm8b1Vm
VZiTAYFGzZQzkRlXFQYGxywQkQUjJ+3IQTQKCvQuTFKBoG5PRYEIbR9l0RtSOM6e
hR4BumgHIvhbn69PH/W8+O1teFjHVoGyVL4JxxZDxNkHmoQc+l4zWls+ZsQHxb9n
eAgjFl9j6S1zae3+vHku17TqRQL6JhCHsUreM/AUQ0dKvCDeSZUbu/pYJO76RM3m
TXzjO+kUltRydW+49dCPnptqf2gk8J/53oQoyz+xBYYWJfOUs8D+7138QbXWur23
P0oLXf/zCta4UsOoXXhUHHiz3V5b7B/kfSh1rMXMJPwY2HosfU1Pi5XtrFMy1iA5
wT/UGEs0SPgqG3VdYe+BN++OlJeJYNygvZhWd3nBuKCB9ypI4LqWOj0NUI8A0G4l
6Hzc/aphhrBhPYVlap6hAk1y5vcaZgrXXluZ2qB1ergTtG2bmGx92pbP+UlBqvmK
9W9ero3PeoVVu5Yl5PaQjHROAzYz9GhWcNJ6uy9uveDVIrXpcvGX48liYcRcbWeD
KuB1b1ddqvBrwYnW1lUnWXD0DOui+d433P4SOnOHP4XjLtU0E8Nmbb4ru34ccnuA
enhc3Mt+u1A9XviyEuqmHgBFiy/YMO0REkH9ujQFnTPrnDWXd2hT5oa8m40jK1FE
fLvN9RL7qd+gKrw7tjiKSyJ44r6020lYYyottA/7l5C2it01Ahgu1Pv3szo6JU2S
tRTmrH4NhgZgRj8TUhqe+xnLXRtvuPW6a4O//l0odwFe89m3Umh7zR8vp4o3Uoyr
I89wRsNU2abk0zRxKNpvkUCquZxaFdoJz5Ipcw36lFKA7fiTujplkcLUVYL091Dw
kKmZeGPlzQ8PEXm3D8I6exN0gJh1LwF4/W8Ma7cD87Wmh/VDg0twjU5qjJ+gRw+a
STxDATMQjeyjnmqYX1SHxTxVTJGrslyxVwjMVnSibGMVZdp5tOlkhGASA5JOk6nB
sPE4l3/itVjF9zXUSIIwYRFKk/W23F4Yli74MUZReNfihqXvozu4rVG3oxGg9mca
YA5Ih6n9JES82xrJxamxCkmDUJCa/6M2isNPgDvzZF4EQPcHZ/j5aTEtGLGRZeCs
tSH/z9GYqgA8ueoiGVqM/Qg5FPiej9JhQbWkGDv+6EfEROvtLqAJzb+cjiRfsp9i
QH865xcj56lDRulz8X27fgKMDjFsx8AE5OhGXU5EwlxKT9xjT5824kW2CNon9f6R
+ylLbf8Y9ddJ8Y5pvERC+DdNpyU2ts/7irpM5BFx6Ln0lUyc4onVRw9TB8M397qx
KarrmrKZodyZe4vePDn8rl4e6ChIh5/RUvo1IIJ1Swe7azgQhr1OpVR5GdHsLoJ0
D3v/Z+1OnC9CSt9WyinWoEDQ2eM/z5nQkN5YAQcoZSZx19mPt426wMiNft2zTMiK
HaYdlckOE3tmHPylpihWiKXET/4yeKTEEhl5PKYSJxFcfK+/5mfctQl+TvQx/ZjS
Qhr/gL6oiERQy+v6Qh2Q19ixdLPzPWYB/NHaq03XGlfgk/1KjUlmOi/7VFTTSuSh
q90kCVriPKfQDDTgX0D6nDH1KcOl+HOns5s09r2geJ24DHZ5pkxUhWVXO3xwVD4r
//yyn7VB2Xavm70KowqrvcRY0sMw0UtVbxT38ASvGSZDNi4+F1a1+cCh511CBYT5
LpmBXyCa9+Q/3LJpbBvj9FklMb154IyIw1bw5IYl+tZ2qVKSsYYZ6gnzIFYFydgs
RiU0xBPZNfu4kHfxxhYVYNEX3rEJCYyJjlhsUK//M9U9Jv0egD5Aavzx5xEvpk8K
XnAawQsaRtpx+bI1rUOrDm6m0mdzhLOcYFP/e37z5zc9XqPxOri0+oj0IK77rgdv
5z1a6RozfuJMKyBdMqoWe6N3Cp+chL3gj2sYk/JlVk5LkRGFmXAeZONl9oENa0IV
GF6bf25tsKeH/BuHkM9gb9jl05ySgTKDyHVB6DyW/cNE+mqvUzlnt8I/KK/MmwcB
I4fs49vYP508brysvzr3KZk75znacAeXCFh3IvkyuZyse57PTvWQFQzgbXyix6mQ
Gzc6k5mnpuXSE2BEmE/uayoxD3WGhQy2gf+KsfAAhQMyAms0UE7M0obeLFfH8kZB
dX8UXMuj3Oegot32QxMYMVOJDUxUrwpPKWS1Kq0SaNb6nZGeMIk8hhBYNbZ/MkDh
v9PpkOdwAYKpM5PJf1KoCdMmC5RZC92dXYwE0buFZ6G8UiZzzot/FS7qW0eDnLGL
o5jvAOUO/c1feX37O025nLgfQ03bZBTqpV1R4M85F1ThvAsA0wewklpOySx4Rg6K
mSzH9bqqQ4OuvuT8NxKlICYqm1VadqXzZTq1Sh1NyoQJ3pziX/C3NrQ++wo6NWUk
rg+JlHMaOb2hk2ifsdYAqL4qGdJfHs7uxHZTQwlroKMyZznjb6jvin7kttBj5hps
Hixb6INgNkey9UeWc1jt5AvIX4iSQT+vqqBe7uZKas+phkjlffPkuexKnHA2M7xb
3VVoCAWjGSxlB+in9jYtESzrkW7CsZqMRUqhZGdzBk6cs96NT/BdyRQvHLfWVGpp
K4yiZ516h5qJqM8z3FtcX0C/S1GhDJU8WIU4TVc26m9usUB7SexvKQ2026io2CtV
k6BGYDqZBfRrc9w8XByWKf9nm56fRjPe6+PjMUilndXATrDvcvrIaT4lzkmnxpgQ
zywLTUMcx4Yx1xgELGgY4qIZ7dzjos9dckdVD9EVawt4/4YJWIXoOQN6lbh52td+
sZnaGpzXF+hFb+eAarvikHma3xd5/ghGT5fawQJNKVsfQC7BD81hvkzbj5R2KNOu
EZ4Z/5mEg6lc2WRt8zz78Kk96pJQqK8Ab2P1MSL6b6kenoK9KecPATVbBXSt/W9u
vPcMqMyphcfudcKcHgk7YDvy+XSddBxlANIw1HEzWyatqpK+1zkrnBEBEy5NNYd1
h2+sPeGWLV7rtu6dLxXPQcpbxi/Uu2TwpjX96wsUb0kkRBRAfmJTMjlOrPG8S/Nw
wZaF5p/HddJ6hQYIjBkuBZPYnJqD920wezAQtzLNBXxgU8RwhB1UIA2kKA4oJ67X
zUuO5TqEzm3kHwSEz7cAAQiQq7JzVrs3BUkBnCE5njb/PmyZk1pt/ltrtmCHJLQS
ykGo+N0xLlJnY/chABfP2X8jXBzmX78dh01iEBZj0kLSMfaYKR4xMynC7+7EzSMv
d6O/UUUSVP28qaLtZDM+9x6y6LfL6jCmvj7eBLaxVvCQa1EFcz1wvnM2WrN6ifYY
833a2guj+Pm+6xAz4rW9AUvkBIAfAl5nyuDhXQsau7yuAfK/ZuQa4Oc+0Z+JyQNN
XvpvowfVDHwzu1aCIOHdajxraxhOzDwuMcKcpMnzNMc713maaae8JTufLERtzhiU
CqN1JALVefB+8Vh2QORSnoC/uWwnCL/mV0HKF5T2Jyq6u0LmTD42EptHGYW23wS4
/8B/UB93F7kExec18hqHcTKQ13eitYI81w/d9PicbzMCSX7eZEr0hhXR/sykY2kz
/y7GDmkI8XobvmELbWGhFEpXFBIWF6wCNNqNNelGX/Pw7jix9n6erbvnjiNq7qOQ
DNnfp1LiM25xzwuocyWdmxBts2AeZ1/s4gOTfAV2X6hM52Od1IBljNxgyDlLgDmJ
ql/6E312fRi1fAN6GtdZ5L6E2axIKcKwTAnFXzZK4oZD52iorsWCktH+pfnRpkLt
umzTDCEGyA27t1ZhqBHghBC59lN8X8C74j+gGqWDPgcJ/D1x8a0/P26sZ05SlBdz
1EbB6nEdzLQjVErYJcQf8a7zYx0YcDFE3mX+9/96fz5+nAl8UIWNWji48f7x62eR
yVYucuAkytjM/uZpPcqna7pUCkUV1OZFojYIM+0kIjo6dnoSliuPxqxf7+6akKT0
gvuHtY11ZhAno4IMMHiWAu8L0DiU6htfwuf2uGmilXTkl314rYFblH27gY774QuT
ubWYaQfNGXGk2xkPNBNDTeaMaX8oMD4Wfn4eElTHUsSKIE250c1Ak5ml0U71T4Mf
xXQui/BAwQdi9kyXXKIOTOB0sG4cKNGFpQZJKLm3cHQIIiNkae5MOGm2xANo1jet
n34YDVauYWWtIffLoUevgAKYz6bhlVf5jQSHFmB3I+ys3kgGgg6X8By9Ayonc0ok
popIjcf16uR4QUfj3rfe51JtRYL7ridgL/ncfUtOshl0mia9ybPGSZGaLjUd5s/w
8GhTkNX7z/a5m5X+fdQOOtUjqw9HRwB5oI5ln7qjn69/oUH7ctegudx394+RD7XV
TMCvvKxhwzZHSAyqhXxD7CzghSKSCUP107nngftQCviLUbmFjO5+XLp8STBSFl/a
HuVeEoSOKlj5XB7D/76mimuy30MvCK6BYK+VmlsM78PBxlWW6JfGLcKNYofhPG6t
T/tPl9iyPqVA1d2d+CrgCwSxmv+nW8Z/5fgiBHbJu520WbYn82dq6NPBJw/7bay6
rwdA9obF4pUrwNrJbF95GtNWDDtZgDeG3/gY2iTYRTDlfjZ/e8AWmh8aqYd7m2N8
8TK9vAgdHYV4aafSF9K4X9GdFnFlNn5TiTX/5QYKzau1cRehM8GLyMTorGnn+Apg
l0nMmR4Opyv0PkJoI8OouF+XpV4/HqqqfoVAhzz5KYOEiewSRlDvlEAI0q/u/BmQ
6pSb/8ea8yLnQlXbEoPTfuB133m6M+H8+AkPpJYP3rFAwdvk9ldFXjkIDB5xywSg
2yj827t+BbZNAdAntSrs5bXjDXqmzHpEhx57EU4WQHcSDwBJMMJlEPp3e0PFz8jW
n7VFyuPGdnG6kYtoHZXHouaQopQAtaDC8/Go3aVM/EPrqZprGLLDiJBjPcaXRl9l
Ou5e/3gQ7bsF7JiJYbtD5JHcW0wdxokzifZFRVQi8VSZIVCxh5b+83BscsCWXGZm
NAa6NJdIRnXSmldu0UvXJszYtcj5r3WQJAl0e1pChgQPRjLWkG15vfH35TN9XDLw
4sAvb1GGYuYxKAfOo3h32BF081LUZ9wdzDZQIjJTEE2oIS6kR3DnPP9tcmNQDGKQ
Q83dU9yDNYSy6FgFNatQwWO1lP6WF8+39wP2CL59k8quJ0i5hE8XMQV9pmCpcDMg
8kf3NfgAZwx3jjSvZCR4NbYh0r36vJnmLwiUAN8U07b2Qj4bTrtXmb1du09aHgvv
HaMmiuLE+LevphUaTc3eKB/s1RVzJvgvsNMCJKBrGZUAyemESlDVcSzXLaPwlfAj
H2Go7BVUH/EnydEeTzpRTzZaP2Igc8yPdz4e96OzXEg0zpn9jutUF/Sv9Il154CT
ww+llTM7nPtNPk/BfwH6qJCLYCZ9BRYkmUcE82Dngc65k5eoe4SdTIaFGRsXSZsL
6and4hkw9wBE8ruBnhoD3bPipEQia34ZQC+hjMVDSTkH1JBvizqyio21hYFduUmb
V/wBoLYIDydaGEnSYun77VJTw3CbRf02BFb4Sc0tN3fIsQK+Zzp6HV6un5oTJmdR
VnyIE6Qpe6yAVScspBK/1W8/c+uqgBE9qqqYEAWTmXVirg0cvu89GQzZvNfELCnm
0WP/oXYauc8HdPlbQn4yeuL3hjUlOTkn3vzAwpDcg2meyNda0rhTmju7CR7so0c4
uRZWozObDjktv7fD3O3J6kT8seXchoufMADc6j/bradHG8hdKNyjw6qAgkZshRO8
18oCba9791iR1GXssCt79+uGYMzyt95AJhja1Iy6TNs0MKlTax+XQrZhHYTt96cl
gZNYstEgt+X7adARnrjO4rmop/oPHHFl5+V+Qy8w+l+wwlEZHJVJaWKGSIcMxXtZ
QV53cHbfC7d0wkL1GvcWpb5MFVR1T01dcXhXPgp7KWLy6+Q4wqaK1Ys3efxsgE5g
7yRthh75mE/2kntdF35jxXAjmpdPs5WDseuYJj9GZsVggA1DATi9Ddhp3R8YjMA5
GOF0xSw3DgCIhbciONrpUJNsCu7M5B+T/Li5I3DYB2f36ZGf6EAL3OtlMljPUCsm
H9rNKyaQlIg+HcaX2tGpUDA7oIPgESD76Hxk3waM/56ke/h+8BQ1DCt6FRkQEFTF
IB6CnGya3ej0GBRHsDJ8nqglO9tMzMw5Jx9EwNushpCJR4JANHs6Y1OGOiaFCruR
iLZa+rrFlUOGZO0Ho9nKNlibjqPePYh9VNx7o+GKhRUxL1w/e9eLlJOPi1W5u0cK
1AkmsPAjgTwuAbntXzB5oYwRNcOaOl6cGupK1kvkNMkmzphKVokoarrDQTzV6zPX
K5QNorQkvP+gISCvtJEecIwarPUaxFdzcmUFQldm/y8/eBgNXGUj1v8AVb/ZPRBM
aHJXbM7y5K0WgdOEQaaaM5N6atvnMBVxqrdwgcSu06XCuxTSgIhrAdSNK4Y9BR2w
JgUikT1AnsFQWOAIiTAcxK/BjklKsWwSNGdhaoWLDSeBn3umBsFLfhovYHa3Zkqq
3Ac0lRBHNkbPvQiJ+AXKO1cT7nJnZl4fzmQcMYGvVtlcpqYkudKlA00rUNFzQQbT
pqTx6kJyc3FXOOM3Iowvl4yrfLVwaphQhkDm/0VEvhcwQrbMCqYAjyWmN9cLJpnA
d/NuIU62QfQUA3781dTwFXNY0rzxDH0qinx3H/X+6jhf77g1ggf+K8PqvjrilSxR
c5M2ylcokHe67iJZgW01xslQfbGjPocpSLAkKPac6K6+Q+YfbSJJGJ7bpgaoeCCZ
X9VloHCZzbS4l1f+HZO1v+H43D1C+UWoHEQlxeXhraxZ8XwRB2NZk+DxCxPEA0Dw
8WyGYkhjBht2+Zah1BzDL6TFHE32K5bYYRzfVKi4Z4YEz5cB3OiHO3BO8tYapUqM
64hOk9mb7Hyquac9VQDMi7UrBJW4uJstqP/W2maQ5nWmBixdQFKP0LEnwf2P4+cg
Xncib/quk2Vu+ptbAD/0z46d7VmTlmy9xpsn5dl2Jm9p5MYln2TL/FWYg0g1Pdry
Uod55URPNtH0RvyUBYOTYfbn13OBHRJdeXk3CibjpxNBWzVfvaSzm6XFbSf6T/6l
CaIlhcwQPoUBaav5mU+AJjOUFmu8ZdWk0XBbXDQM0DKJ6RrJgv1dAFNZouPAx+Fh
NDz+No2Tke4qlMUxdlprBLT2Nd8VuEFNFPe3fa/PfdvjdTgq8C9NuA+2m/yJrC/h
CPyto/3bkXP71sdD4qHs1CtAUbbdWF3eNbeLwo+Bpn1xmJD5hjISOIjWuZi9Bsmw
plirm7Wt5Mlcu1nnSHr1oa95YIp87L/axmInniZtA4shdJJSSzJYpT1ImMj/hmF3
agtxpP8Y5L2+UqYlxaGcsuJ3WQQrjZ+s0eLEWHsAWPoH9itIOIjpfrIfwAguj1jH
qa+XOhOyNOez8jirteOigPpn5aoB08MSt+unt9icNwCsWipdZIrCeymPP/L7U60P
futYJMQ8WiiWHI69xxRwDr4BrEu99gGprbdDu5ezC0nvMKvI9GlKd7Rc8x8VEnWV
G5ZzgM4ow8DsKIciO7dDVf4LuGy1Afu6IVD/AfyU0S5EhFVntyEkKin4QEi46ijQ
GGhBAE5Kk1d/rUhB3bOQKYYGh6BVdl27aTnWLkqKHLAtgJ3q9RxaiPSM73bDQrxC
43hHkVuusrMgu91fAqRmXM6JwgoI68hWRlJNB+1SLVzSe8vWsg+12y0YuFI6WoeA
cJPLQNXZG7VZaQyJL57Bk4P3gJD3DN9Teww7TP1seds4fx68DZiRZF3kKVey98Y4
SvHJg8Tbge8rbfo7bC6vrq+Fi/AgUO/cwgk7c5MDGqj4dTvfvbOgYCrjFu+KE11e
QkudzL/ErE7YMIE1QsJxG+IT3w+Egv//ECvJe15wmaCDzRSTBQaINOGvCMZQnHGT
TQOQK0huZoRx1Cpnvd8MGPf/RjiG0xEZ+pfccU7HOTs5iEk1x09fqNcfpQlIFRwP
ucks+ydjho6z/PrUAlGthwboZpFL2BSe515eQYVTrNnB/D+NDAqadqWEisEE24c7
LyaynxOj+bYr7zgvSm8V4rrGXPkHB4CK7vAM5qBSmokrh6d4F9kzzh+6ubOjEd+4
Zzf04mhN/ldBTp4N30KaEbQts+1j0lKqP0rFubk6Oz3tdj1e0b8d/Je1nIzKxB5U
TwCNTOXZ3GXyKtAas/Cs0tTdu/WAbSJQ9zPU8O70871CN+/tkcjtVBLYxm4RobrY
qUXEijoNNYNOoXniOxFKf7WFlmH8YnRobuB/wKPKvQ/KGtZizIr0LALtJmGRgVip
zvVj6aKqjJvsg0xh3D8JRKD+7UtPx86K88uT42NAXOsM8KI7eKJXDtLdkY7SgUBB
M+V+go9XHLLIemWR6TymOyi56BtGNDpqWBPNfpSm143eRhDAeVAhRakK0B6cthPu
ck3rmD9LCv2g8AsJwDccIxIcaG4grXLaSY+GmDCVHhRytuPu+12kKUUEKiSTga3R
Jd0pUaTLDARAl0WyZTZoVz6lafdXTealn7amzfq8T5mMpb1PmJiaCqQ+j6E7feTh
fSWVM59DChdfpsEqsR2s5VR50m7TwjdPDAEDG3yRdJmdamxzPpL+4wGUuOg2GF4l
jspEhcUILP5ZHusqPkMv/J9OpOjxC4zJPbDzkANpNeeX5HoAsXt8CF+4NWUnuRXw
44hKwsV2+DQxvNXtF468iCGkwx7ODxkY2aAy1bbWEaukOnPmOUkIdjwaCYuWCJmC
XjmqwoeAulwWINJHPlnN4Cvpmh2VCbYtdjQnyhxKzqXfaATYfYzL+npQedgYA0il
Qg1bloboxnrEqjP9KF22veAKIoEGbFuQwqY1My63C6E+u5mCss7NsPwhZHqb6SKb
zC+MolCpRCOkTicN6nRC4/O4cwir+8Y7fPS6tTJSAVVMBZ8qjdSjld5BA9voWzMA
h4Mf/UtrlhBXNIxDXlRm3ev4HjidbuP+6ttUbt8jq31Xywe+tojDSvhsG1XcmdGF
ih3cOmGsZg/rZd01Mh/oRXvCRsfY8I1Js/RnxNRANbWzlbJFfFe5+TY5GGOk2FoS
EftF6G6yy22oWrn8JhD7VwYzLwmPPQ4+7TbWubUwXlJp4dw/RU+OR4EKsdyrv1XQ
0/VhpkK/QraJ6x/QVDg7x1xoTIpzRAuzJ2dam8QiaUgc605TL+EBl43O2PaqR3QV
MCcOTGHllQRY1yRfI4QUEdnDEGbIzzWtefTI1pkldzrKm5QVDeGkbDX8mXHqaLd1
D4+/m5YG/GHlqXkqCiAscpiTfJCUGVUHYLGGD6ZovXk9vONvMkGua2mizBfGOi7c
GytDiObf60v+vaH2wgI+I6Sy2IrNiJloCJDB3HJX4jUz5O/+aU0kZuTahSGorOCZ
cO8WEc0gKcN61fhD225cHXHNbCVtAzl+iLhTfMaYG1x9KsfOp02LoHc7PCMaXVxS
MSdg0w0aVMGpeMn9u933NbOJxATow9JfaDTT9PHxELffjCg6v40ScL6EcVLte5eF
8bQvVmpd2thj+jF0KfXRXLy5PKUeqmFTC+TG7tOyUPufB0SSIW5l/agVZyyEOl3u
i8nrdj/fS7rNsp9sd+0N561My5kt6LI6tsK7nQu76fUcVw0Ds1EX0h54EU/0caiN
2ShDkJQzfezZus3jhO07cLqb988NPHuf/qwiSLF+u1DI2JU0MyU9SmQ5+rgov3cP
5aGEKTl93vtVwL9UnxAnU50zsQfVuHQtVLfCIXq+MZOgrqAb3lgILIviJErn9A2L
qOk1wvpm6mqNbQgxWfnhs8GsCDk6T2GjlXQrfgfl4HA23SNxJTGMcCPpzxV4/BcA
XPxZVVr/b2dOW20m0uL/QqDQPawVtz3KqN4MYNtue7ffi1dnA2zOERJYQaRhmHAc
ecvHBcUnety8E7rzbQH+z6GpLycKmP0yky7q9ZA9MJsqRJWIsui38iECb/HuKaXJ
xIIYaEPV2/GXmrAi5jNEVOmpZGgmd5YElAj6Q4vageqd/SsLANFOyLGENPtrvTDh
x3uI0FArPB/Mu67SwCj9keuEMm6MbmtvbRgeJLv9MQfO5Rfw/enveEiqUqNnlQG7
PdU2DGix8fnryPu2qygw87T4VfHYKCpYtMX6N0uAwkIrkJ9GziOimQY8SkJJ5cGR
QhP4/gwtCkzCtVVM1PW1q7fTOHXZlXE2CEpXrMDSatuDR5uNIYB/uueXGVcyvDT0
cf1VCw82K9xbZft8TFGmOBhc5OK8tq5Kan2EKU+lgp1fgK4SngVpl5llfphZK5XH
Bg2j+Y9o+7YFdFR47cr7RwBaNhoxFxB300T1+780UIEt9rJeoAc6RAFgASR65joC
9i3SzFjrhFi9TbVBxumZBdJPeE52/nuzJniamx3GoeFE67vf9aOFgB/MCjK644CL
4sf1vQEG5rkBTteizyVxrCNvWJeCdRoyqv1zF2uuyL3w/11BWsUpAN1LxdfF7Vem
LZf4fpBUQyJr3PNm4buq7kq6cgz1ZqDru1rq06P4NlTcgvpX+Dppq2DBQvDAuU5s
ly34gpskfQuSZidbBffSrN6m5wsSqnewNyRnaAmxQzJcfm7W+4XOjw+Y2aum8GTb
pbD483HiP071UmJeHLimkTdfe4acDaQzKeX4bdeXewxBZIfZPjGTwNl8QbN8osdd
8ccAKGSUxpw0BBg514RTjXgbRlfhQ+lHrJReCQvJzoAr8DZnMsWoMgNsLpqDVHKi
wNetPLMaBDM04Gv3eHwG8kCg7/cLYVVmCatE07a80hbTgiGh+G7dfmIDpVoY+tdS
JIsi8Kfpuz5tylH44y8kV+yvwM14OM9pZBni7XJFKi8Ly0TntkTcEla4Mi4MM01P
TkmQVqSche8H7kVoN6IpXFxnG1aWnBej2ksTLtRADB7opw/RlHImRL9gEAV7ghU7
jT2Co9Un4sHFlqP/TVZotDFcP/kW1zLSm5r0xemQF1BtYDSDKcdQDstMos/nMXZy
dckPIp1WAwuPBL3dKA332Sca4db9CzOTY5e+Wi7EcH2x+1c5Kh+dG6XtxdJ+/om1
hfynwS7qZgqbrFRLrMseBAI4K7aSV8bN58CWUGr99Rgr47G2l4bXKZbawym1Or89
2DCbVHWyS6NsUnyCQqknJx8VHSi1pZMxKs09SEfYneYBdxooy6iF6R7w24Astq6V
YQ2ka36ibitTsUilPP4BU8DAMqATQN0QtcxsSD3Am59dNhRT/hIPQ/hg5VWP4FEM
67u7OXygk+PNFrmv6OalVv5i/RpLORpgV3S+v6wEBV6LHNfHgz/cBnyg4fFymFLB
oy3uKdS4oL3euddletMP1J0tDJJT08aLWyugcijljsPyF4ieF2sF6JpUV48QasoQ
9UUK+O/wuT0wm6Ru1GQONa9yj1vN9kCX2xbDIF7VkPqk8yxZyri1smRJckvIM0rJ
0g6zBHJA5I/+qH5Dv1OU519VIY8ROvQHyi0Y9w3OxFjrzW0E0P7VYMg8DLE03UZV
sFoHlPju+8Yog7IKL0g7jHdLfPtEXMuhlU0CnzDWmTMW45AbMDSlm1RI2bUoEmiL
PWoi10uRu4Yeot0Cy6BS+KhuhT+5P0ZuPAWzHV9q0WRx4T5EvldqiRQM1ur1RVad
zi6jS/z3ZC/3o6d/2wGoPqfOuPxMXQMkbCXKXKxxSaUFiKPFfNZXa7amtsKENdQk
OGMiVgaLXguBpAj0A5V29LOOFAUN0+22incECMSpmMNWFGyfRi8+MwzGrJzbromD
qp+q+k3+JcKKOR4sV+SlFqhueAXIiBC57qPCBbkbClonCsdps8Qq3z5KWJDxL5rn
QcarMX9Q+Z7/lQDB02JBNW48h3CrvqfpVp5e7gQO8ch6Dk3LxWKbfEYfBpSRKyxJ
AYeL2m1+CqH9N8fIKupJdOpwj1TiWIW8rXRhgoasygQqOZOQ2dlmrAfEs/JMagS9
1dsR84vMVjH+8TKDoFoTblsM+v0p4xBx8NgWrNMDil1jqSv7fpaBwozdbOyOe1SR
tomeOZvLf626ymCAT2B/o+4hOFmpP90t4pz1lO8j2ez7r9dpLlBkHA3Ffrc2laeu
Wt5cz8Yk3jiQEvzWDPfCYlXsBM4QsbmojJYjr9M8p9VT1OMs49yAApzgfLxZ1R24
86pIUwxCLHr37utP6DTdD6ettlbUDXlNb0ePL/H0ZItjNDFRG89/0iaHNxqeptWO
6BAgYu+95ZHHLQ78btCq7ov5L55fJ8CDnOcyAt4QYW4yTH6M3tH803lRrnqEXQgP
Qb/RCzmZ3z0TIn7POtpSIT4OqGZxB9J07EESUQrHEYytu9a3Wlh1sQOwfcGvVznY
uH4KdBiTeCHWvM6XS0mkcHhxpUx4PN1TRdCPNO9hXVqeeujkE+YGHJFOsPng2Xdt
TMtUlpCszCVMGhazQXO1D5e+ZxekWIRGko0T/tQaUIj0huuruNyfmri4J0W8orCo
Immczk8zCVGoix8tQAxeoTQVqwNYL8v1Z9I89m4arx5OPyw0jCFCSxbGoVpGmPff
LcySPzlKqJwTPTQTFF0DoZElG4TqiAPGTn+svglV6S7oFNXjq3qVjy8P3Qny+tNg
NTdBh1OVZJHpND7r9td0A6WCnZYbOhQ/Ew66TcmYxYTicNMUdqhhq4YDvfdjZsNa
pxymVLwANlrhJHl+RQMUxDNZSV4/DT48Ezpnrow4fH2foq343jXjnLV1b5szmgDV
XAKA87vJcxRdcCla6MCAPrnQag7zhg8e6kfe/2bCZIWJ9gmsDpfe2M7t6zc9shIR
78NKDDN7peUCdnu7FgT+HjGavlDIWAn+ffPZxiJa0Ikgwajv9+aGD225Hnokj4Ze
keiEj4bYYqGYg5S43T5DxmCtualPaeZF9rekh/g4AR7f5231txRsZ/AJfSOwc9rn
iZhwlkQPxuhXitWhJnq0gakRiMndHwTbtFQ2ZGqwURIZ5SNh59QDRY8NwrIsBkno
TW4b/nUlqW/jsH7JuD+FkpSl02UDbg9uwf/xfldBkipuRAhjfPyajuW7koWbz7YL
/96fvsVXZ9at6aXqo5Fpzxhazp3Uwz1+UAmc4pPRdIS3o2rPCpIi/b2DMkc0jsGO
VAylsCy2dxVHLPijARBt83Ckr5FRZy7HvNjV/ZFjXzOC60vS9Xf58JT26RA0jjZP
CrCHssRWwu11I6V89f3GEPcOb8rZ73VOkxdSpJLkR+aPwhYc0QTG+PcoLAK6sefT
FPwi6e4lMZGW+l+Ib/XjZDuImqCJUfmEPBO82mq5Y+AwCWcywkLRh47oFhEAE2dn
3IJP59MKOhZ4+TAtllung5EZM1exfT0Cjl/zV7kgvpscqln/T2qqhvmX8uWFbtdk
EZ85AzQsf7oX8zb+yDNbqBue5dah+ySIHkmL881ZCvF8Xaeaq0KIUVNULMK6aaYF
tqZPuzlYu53qWD7HuAhE/hKJ8/fZlmfrR1r1WOVr1O86/Bfj991ezpQZdZJDFr9S
1N011BBr/RSJ1QF8WfN5LWg4LDECcfv5zSzwSfzo7awit2MiSXuB6Td7Iaqpt+ss
8qgCLLWWnVjP0F6Gd+hRyb7FyGrIs2VhzPzsi0Y35yRfgcjkAsEPvzxEBfDApZk1
R0AQqK+ISQpOiC2s4uT98O7CsBE15l5KRqMgi1CODymuNBJY7Js1v39B31tNhMQ4
soeilLRLRbXBG6499XfXUK/tKosITcago8AvhzeHVSlwYS3BfMrNbHFHheHBDW50
b6F35A/rJWg6Orx+/ceyb98fo6cS0wAdkiDq8IdD6L0A6aKpKmGeKQ7/0WSYPq5X
e8+EHZEGXJ2I6UMEc/c/rG+nVZArUPrGqcgPFSZC6lRLQ9XW1X2cepDEXAoIyVF7
vC310hb62YWOvI0dlGRTy5Dkw922HLe+quvTRVK3u/YdBKWLNuOI+Y6g0G6mw5zu
jYyz8McY9/m1in6nhfT9nuhserbvXq1KPcZOHZIi2b/QSaqejBHRQBuuVAcUbSpz
IEeP/X0JP7BKtiISyK7+nGGzUFGzFnJPLhO4zjzGsH3914o51LfZ75JeiZT32YMj
cgpVpNgNaZLAESZOnCS1I1ev8xrtcg+Qf3ItEcPwwrEI6k2Os87UM/g96ACu2IYX
evRHSZh24NoG9O5lk48zdt3toooVK8F15VR3LwrPzFKmVeTCoLz5zwtOzLAN+6p9
Oi+YwJ8zfXWQSCDrbqAoIEva4KHTe3GDeEGLYUE6pe/Pt7RGn1BIL2D9c3YpGvMY
Ze4vGOyUNUA52hu63UMvYD2ENQeupvU+XVV4wa24gMymXNmvExSvgZzzCN1QM0Nw
6OxShWkTvj4mjD1sySN0cesSGU54TW1nGL7U4iaVGKsW+8WHcbx65dqdtkiwrilY
38eWoOHtWpRJ/4qhuHqSSD9kzayh6vilSa2akXoAYsDDNGvgY8E8FBoFqyiwjPd8
SP4u6+CVhPyCK45VPHgyb/BirCgNZgjTzS52Yz3q/C9Z/IOAyZwwzHIr91DVQNEu
Cbit/5ERHXuoY1BiM7iCRg91gvjwTzUAENaHA5rWwB89juEtndGUq5U1rZrn5Kpp
lX8XXvkVra14le56lrcKH/NCPUsqdSsRk18dromzkPFOgvwoQ+m0WGoMgVPDkeUk
M+d/GvcphDcvjddeds9va3eyE5LcuMDnRyHRg2sVXT6TAPgtLtn4uczDIq/k51Sq
aSrtT5ze88S0WTeTfMyX6RdvbbkT2+BZ52hhpPuE+G2GTGiBEYzY9f5Py/z8AXfn
RefhgPLQWq6kYsgBrQMp275bX/ocnUUyGO/oU1E3EV1FhIDeTAGsxaO0WyLWEfTB
tEPjYfs8jHHKC2rpVWGtXP/hOBvENn+vZR4pkE5KXrpz00V2OOXTqfFU1jbqyhni
eQfUSeL5e3TFI5prLX7F9IKJBUscwGQvcrFTiqX0RAK5ihJ3kDznxmJrUM9cRhbx
f80yylTj4tj8TZFlxag7VPJq9zvafOm5/rtwvM8dFt4Opo6SkMMOtj85Yo/3j6Vg
4ITTaP4VhV2QNiT99UyBvwUQ/svjovuKaj+HGhBl02txnCzH9Y1WcJ6051dGa2lz
VyQrZUj7U9nGQlb+1D7d2icwFzT+uW6kCgqDTR6lq9ZWvu02ynmOHt4QxMrT9Wh2
i1vnrxS75v5fsb9rUH53PNrqWnSLAiXrin5C2k+legqVXKHHLpPyOLIyKe/eDCrO
4yQTpZHSZyO3clE0hCZ2y/KJ04PObheFAmQByOPuhg7sIKROyMjlE42Sxqmy9VJb
fsdO0/gfxQu8N2R514Y40X302sMWQpWZQobqIW6WrdmrwKtN4SYEOA+H9tO9Q9lR
2E1kwl5AVccAHlAMA+ERPHTvjLHEY9JtjUnMxttTluA6OjxFkjQLA6sYwjPNVPZ1
f3B9r3k+46JiDpR8pxxH4z2I01c79nzB7jB8bIL1HQ0rHp6/PWrmoFsXSeOHG0cu
NTWjgxv8OIuOrLCizDa8CUI6/jD5FCOM97ggZH6gQTBhGm8FMclcIi3bHD0KIGXk
t9j9dtrrtsxJDwmw2JovUvDX/hMhIhkdOJ42z10+58yYsJDINzbjQ9cACmm8hyEE
ApPqtcTRI60/GecdSJRsWwhcCYAq2spzIN5ZDNYWMy87MFOR+CubyWEa7zamEVeZ
M5V6cMMQQ5dMbdKt4Sphx9LpQ0P5hpvN8gkHSwFwR634Jf777636ezX4zdux8eiC
kgiBGzcNixaslT9HZ1AEK0CthyK4UZLTMaClU9hZyWXkEjwwuBdVWXExJ8fzXnA+
YCGqDQu9cXfLkIUe3ClSFQGR/hsHCxpH4SBo5EFwODfGb63Kc+jTXpdukIOxvqFM
T6VhGhOcEai6l2iPZrtbibJ8j+DpR0eZkcBfpsIvAzyaZCuy25M/VY+dmD+ug/jI
dUuXCNbrNdgCn+GML/Oh7IpmWtwu+4pPmggPpxnhQ4mEbzC0a0IrnDl8rEx6HV8u
PdwHqWTfKqauDmLYROxaSixM5dmutSvtFOrzbiJ8pWs5PAvN25b1IXaic9/h+zrf
S1iIrchGNSLkE1ShxMJAlaAFk/XOZUh86KYmDy/7TCdnxWvpUaKPzz/uDXiBjp3g
1kh9CXVq5b9xbADuCQeKAyvODn/Rl0lAkSFj/eI1BsTL+gxbvRAUPFtZk2HGjT1w
qR6oPeZEvAkp0q2qLsX3wAXS+eQ1/5xVqZZ2JFJSpHxWr1p8n5U9Xoh5Jjp8BkuH
89y6aqJvS/nPpjZdH1vkaIyp7UrUy3/ovdyqQr9dea8nA4zy6/Yu66CXSMg1+D7P
uJ8I5zcIm6f5ytMu9VX9L8+OqI+2/QzMbGOLwM7n5MjHqPVjbWO/9knXi1yGz3kT
fmBaQXCCS66NX8weJB17sE11d7FDI2FljABWXw6UpSa/cJ1/KZSbHveLZacJ57rc
aLP5YaZKQNgnGYgArcooze59WSCGj98o7LKFgbrgXfrSA5x1ICMUHzowuXv/oWUG
dThMbUEptfF4RoV44DJVa59DIF2ZanMAAAiPARFgO22YgDGn3TPPjVkABHYPxj3G
+VbZCUhkpaOcbLGaYGdVZc/qiuepdYoJdH4s1exSU2VTCgIrwJSjfDS1BsCscviP
6wnWaDVKvSNuCwbR3d18xvQWciRC+10F3f+NKDHX95owcOWgcNWAGCiMNEuKPsLP
j2sOuB0wFnm46m27Li/+FwUAHxfdMXKmS3q1ekFSZHlZL/RNqd3xDTSPhU6QTBbA
v2KJ6gfE556jzW1BoKxKiYT83yq+d8qtMK5py5eiY8ll50H2qbgKJLi6j1W/VGeh
dbtN8WR0Y09a4n5DaD+jIIAEs0xW+h1CCCFmDAYyC0CkNl1i8yfu4FXDSX+txY8C
uJOIeu00nXa8nxySbSjJN62hUbE/wbiWHuh18w1Em4WK7tMwPIy+JKLQbOgzGw0Y
XCmvZuY46CL3jLusBFCBV9N7tWT/OMqcZyPfdLDDFMcP7E2rlWijg4JQcIIJT/tv
gu2E/Z86jjqgB8JglsjasvRnmquuqcn6W7cnI3r+qNOy5xNZJQdoWgbz5CclWu9b
1Ltpyyi8cjuppI4FXpy4TDQKWEPZ+7jscY9KOn7TgNb1bnLymrMatGq3ymBXc8VG
XfBdpSSRSqOaNy1k6cmwhVtGD6/J2WHHnrVd9iFSP+VH0SOPQmfZWZv7KI8MIg3Y
CBl2r5BXBGWkF+y7/toYlYpteO+/QheT0le2RnhGpgY7xE0x+9PlswnwxLBPqvHw
8Z9nt+nP2DLSfDfq5gbc/2gIY40UozUu+d7tejm+SvDNRIW54x2Jm8dIl9JcNMsD
swOGNozSQ9V7F+PZ+SgzbvQWnU0ruPd08UwR/erDxxaPA6bjTh20SvXxdF5k+grw
+E4wbptJ19ED2m4Wgiix5Pq6XVE5dqkWNnSRMnqj8ekxywwJXj1F9hEKNsMcCXeH
qUU5RmmeOZbWdyCt6KkPFD5WifxJ74I/GYqRs/ljy4gW33J1dZtUX/lHZYzFRdZ7
SGKwdScmK9mmbVBSsY0u/ohL4x3/UOe/TEkNAVazF2VtcZNSmzIQ7TwDP+LTxieL
vijnySrrUrAa+CD5zuFy6RDRVb5eHcc8YCERcNFxZlCL90bASRJkzSvAh9Y2APbD
RfTu/3WsVrixHicghUI9EbRK/ao2Wdf0AKaxo6sjEfD3INmN1OOsyh6ksmdkQBqG
mFIcNZM1lA+pz0MfwwDyg+H+rJb+X0krX0Wz/aEirlezvCTJgkBVQ5PlvvsBOccY
3mJ3IswUaF7Y1cEnTIdG/tuzE3dG++mXBOQ5uwGRx32pyFVvEt0H7ZDD6JTa9tFt
MaPz/favzkWIyKCpoEg1jM01JbURHqLocxMzPMCZPW55MUvhYFkpPMx+4wLmtDaG
MPvECQ9iA9MuaNe+UvvobRaQ7GADB/7qLF7wIXIqdWBPorxafHWy76KleUb7rhPG
RouH8Anw32AoOywrN2QeBOltescsSNzBpTG6opVnYHJNnqFQPJGI81NEcEcTJsa4
I6NJeTLxHcxnTN98elFMC3lKVB8afpoCFdfCIak6O9SecvWa5XG8LFfLxqFDqTEg
+AyvogQKyIFP0f8rP7lF1Wnq+YXHNldFpO+fDroH4LrVYDxpTvcYubhwulfY+Opo
lj03fgQlvmd9uyzYeaPqrux/yb9HO4od/ZGGMSHxpj1J2t95X2FGqpG5nbH9zBGr
96kfGkTI8W3Bca6slSMX8LUlOeoZi1vBLVb82ASu7NrcShRtzLFUi+A1eFZ4VxdD
NolSydo1jYbC/e9LW4vC4VdPNMljGRtaEsnJ8eJ7NGNdVu0rcHsmCScc+SWkL4FC
NsrpyqEdXJIZjPieBydD0PlNnhEtAeB5deE1a7ThwPMASG8B5TZr3Ddsv7XDKl8g
pONEzKuAg1Y6twz04zWIoyhlcp3C6ihdJfWAe1Yxm71JoPzhb09cJDEV38rjfmgU
QzoAC+cnIvFhcaJBLoV6eTqrenqXL1KuzZ06vtdVFKITh2TC2riTKQ/bbN2EsJr3
7cXi2apw4mJCZfa6+ooz+kCxqwQFXrunOe+clyZUVV2baVh+QIOv4CoVz6gi34im
KmrJhE7GaEB3Gc2BG3O4COMf8s11uF7z0w3IQE2nvKjiSU7IcgEforCDi1KOAWu7
70z+cEUhSYx0ebiQB/9mS95V8AgPSkJ1ICnNIN8k9JQkbnoZjvGiwslVRDDSm2ZO
0Nuymuwd7LC8lwtoqsVQhN5My2LKGq3o7GtQKyQqER0wzlK2r/mg2/YjGps+VU2w
zq/7uM8uzXImQP4P2VjJwYp3OZw9r1zkkUhLDNDxknghBWGoT0YH6GU7cttpf80u
drYRrGvCbQPHefKkhP6ssYLb+EfbwI+vzbTA9KtfwMTU85BNg0dDh+8RHveFE1D2
t0x5ILL8/5acWvn9g7U1btwuKfdViSWSYWC95C8Juf8j0wHRFbd241JpcWbhN5Wo
ppzPe4scTJ63sZ/RAqN2pGtdI1JFz32wm2M+MTeYnrNZONi6CYnguFIycEEeCKPh
YEX636n6DJOpJVDZLPy3XRglOPH42a60OI+gvuiI1UBXaADbNEWV3G+2M7/GlRCi
UvvAhiraV162sf58631v5Csoz52fidbL8a0X2rHXCr5SDhHDcmMfQ7FuupcKAuS+
X5t7Nq2a6301MLc0DI6UvtzOcc1w669Hlb6aoR8VenSN7+3IyvtLpOSQT2jvZYLe
xRJVi/t4AzMpgVHcLCres6j9udo/5SLriZEAs25D6KVYq+MDQXmM+7f0PbToiVEL
RzLV4uf1pPE8KL0Asy2xwuq16HuIjWxmF3ZyiJvAI7BogME50ZsxfBnyGIhqFH2U
SDIoXW19zK982rqKy6qfHtIhOzCJqK23Ikp9yX+/KE5lwbuwP+9gPyAlkGANSFfR
YUtfO9Jq1FTTzRwvTFxvoY+geqSOOKMCuRret8qOMT64kRlyx0c/Y+kDREFW4ez5
n9bEKjzN+zZQc86H6jAWcbM1BHJqjJIKaoJVcLmVSLRP3TrKFoDmCKI3alYl+Ul7
hNf/9zQyASNWOFzwj2EUm/8fQIw89/mywE28OyR24q1PiKcIfChW8TDhLjqRGwh2
mmNlEC6jO2MdE5iLIWIhQ5makkaaAQHl14ea6BRvY6wt1k0fRRIqQ9RNNShKW925
mlMfzfsc172rKPm1U7GAPxlJULW09rF2fhQwez3X18Z3ASAQ2+2WNJNW7a8ekf5h
0MsoV+cnnCa7xDvU9Ia+eJRKidyRHiIVC2YK9L4hahWV8yJXc1Lodl6D6z/JVeFn
ZNRWCuEupVTfta0gYw2FORf6wFy7KTmd5yFxg09NBkawbMmtj7uO34PJffSVcACL
SXOUZDCKaDJ3p2hXZ1btCKX1sGBloG8nmJBqmcTqHBoNVgUulMhsWuWUHnFDWEu7
FIXh/vOq2QIDljNqez7OzQwnHc29cQHw8/DuljOMtsXvXNUarnxZ+M4vgFzVeNXA
X5VHYBT6aIODZF4QTRKhy4dROLiVAu7Xg6oaglgiSduYlJ6Wmmqlq+V4+YkxnNpm
dPi4GvWNH5UuV4HAx/0KE7Gx5V+I+B7EDB5d2z1qQqNOlpmpejybaGHwkdqPNuSU
ac97Hiv/zBMnQrVpRV5SFGSd9sC71DgvKuHL2A5WON4CNzMtBCN2zrP+oU52e+bx
r3prTPK+oTCxoK68WjEd/g3l1vaSoN2fap190l+KCM6U1l/GBXwi0R5NC2VICDt1
fb7Sd8JQBaVG1mhVeA9A/1m/BOIUm5bSwWwMORjEMpH3Imx6JnsF23v1+L6hTXQz
p37g5gxifjyXk03Qv69JtmmkWHiS/WSvdK+BLhbFuPfUS5s9RBodbwrJ4PpO14np
BL/zJGr6jnuKTsLXn6yYxZPp47mHVqDCei01hmRD1v0w0+Z9XwiNEblIDRmVpdsJ
FcGqQj6uFEFrsyfyYdKk6B5sHAQfqQU9I0fd756qusuIVe0XuVdz7NnLw21js5Cu
drGgm7QvWRACQbenORYfB+xoJaSnNOaINRinz4SOJsbRAYaBO4xOfbF1MQxWwNp+
itXzox+KSNyl8PDfIS2G4DrUTbe4twWd9CPCq5AjBbzvURG5hwCsxMuWc26PXZxM
uK0bhPDeJBmNZSP59vNGLCAbMk7GrwgzWB8XJkXaCfunJ0Ei4zmRR9wdWEfJ04lR
+lv7MGX9q1AiOUab/kmlO8ADNHZKwjnYoqZGmbDTq3c78qxbalDyPLyJugIfKN/f
lzD2oUFs+UpfjD/JtBUpaMb6yzGLVhz4q1SR7xhi/mWNIC40zwf6xZJYq3KAmw2B
4J80ZTT1MZuBPwwtoo6t5kuJ8atUDb7IPxp1HP2z687q3Dvjt8EmX/RzOtgzarWt
T2fWFheLkgBF/tOFeLh6jMylxekzGXOg2AeAYeXNibtopFJnYRhfqlAAWMwKm8We
rJG1w5rQz8n9Vtb5ni7UoeHgLDVGZvzl/mw8zCRhbdh05YStWTdzKW0mhLCObNN0
xZzibTifgj14ucWwook+raLx5rAu0Edbn9qnxnkmvY+SFZEyr+MLsdVwNEI0ivLs
T2V0B4nRjwCcIy1nCyaxPcWCS2zlsx7tS4sntjdxwm53yVDT3MHp4/hzoMIYBzD/
HxjYuRcD44AiKvpvOYmd4bO5A35yyXTQYb67tOVcoiF7kj9n/LvmWgB/YTrWNK1g
sJXsVQlnB9rT8xoTOfvdGZiKTFk35956ROORaXYQt4PRk9WpXRxpf29L0txaJ/Lj
PfCGzvh1jYVyrl6/PltTvRNkYHg9dDI2Ox6IWUGeEThu+WpptM/hESREWqNdxzlf
nF3h72/lYjRxQK/y1is+/q7WB0eJtkB062e5YEVbEyk6atxuk5hoIHpT+VuWTklN
sOr0kW3FQexA1VVQwnB6ulrwHIp/XvmMNCNSlNFfTZn1XQrx7Vrpf/P8QxtIykX9
vIFkA0idBkhhRBHgk7haFtlMPLQgLcPDtM0kAziTy62BHDbDWfVtT8OPQNxWpAjW
JMUFrRvcE6L8vsw8GQ4+LpezlFeBedNeNkI1J+YvfWc3jRqqdjAubwCI4+a4PskT
LP8WOZ1l4xztdmpmy60WD+/PmOoat2nTkvukEeeUj3UY+rEbLXqIEdOev3cUbzcX
qiVbYJYoQF2QTCLTG57xhW7O1NQFdsAULXruzg4i0BfnRl9vUN9Nl1ksCt4uhFSe
SJaVi+8/Vw0JHG12Af6eoOWAr0Zf2/HDgrRuMDXsZcAhNBpATcLqICOT3zvSY/s7
ZW8PaB+RDgariO7AQbQ7iRNwC32gXMJ3YSyrh+LnxKg21bx8PQmrKP+fydWoVh9h
vNfB+TjC3P3+4fhsA+ZFBV5ZNvj+2gNT61nE5Y4LITRkD4aQfCYafO1bYcVy7D+C
AwOchs8gIBd98vpW3Ve9/MQa98JiIg0Yz9j/nGKLervDlyy6to8Ic28+Zcwj6eoz
gHDeXlceYEDdVCkmNdyXAW3Fct9CLCTRUNA5KwP83NEBhnHfNrOf5tqrhJNr53xU
c31BVs4GzlP/PGdMTZr6bsK4e078einO3Sy/NuNfFAHXluTfyqjWb8hjaTh1xBkI
j7DmOKNOC9IJRzcHvMI+gOn2VBHxEOfiuXmk7UBjWXNyMd8dfZlqko7UN/2zduQr
HDz4yJLFKpBWbiUs4GCmo0+FQQcr3Ykm9IYmSRZOyfyQOy7l1nM/3G7LaLZM/QwT
Voc4EK+DfZEK2z7Hn8+w28I0udXgH7rYQ8+2v6yed3WwtM7KCg6lP/EGeZtzxdk9
dO1m5tyCJ83Gt/fQ8LHont/qA+MPaeW+nR6HZHk1VyOC3bNSKEeMO3klGVIF61Ur
beUPh/96NPuuSdxAy42HuVUZIsWoz1QalmmbPZYPsqMCt1MdIBdF21H4CZUWYij+
6pmtBUad3czZvvuu4rmqRen9V+SgEcW2GpymJ21Hx0mm1c1X630H0IDj49FXV7c3
E3Umo7CBDomdTo03TgvrWeD6MJZ4uPYh6QvBYSKf42/BpowxhXCQdyD7qAxOdYaZ
o8Y4cmSRiAqO+6ow8rYaVLEIgT25ln/73BxhjxpWcvg11FEyiG7nk7iZI93aYcRv
j1xxuGr/WRoZ+53IyLeYhTem3NItkdJRA6k/rr/HdSepxIOV3I02wntRNFY3sTyN
qwtdG1HK9kiKs1KkQRS6b5jjXzAW69u73jFYjCOEINgiWVynasAK03djrAd98dpM
WmaFKNAUHBU9cZOV4IYFp5KXgFguvnt7ELfk+U8dHmldUpihmkx2owQTceSiVTbo
0tLidgmQW3z8/mb4VrlZ/Gt7U3dRpmTpyp7NYTOsK27sGnQyAQd6dr30su1/1KRD
QrUWDhg1PczHHlPF+3ca1hod0FI0Q4P//BFFvHWznGdbTBm95JBG/riP7p48mR8x
X3XYhD5j4CqvRp4XE11iEZoD0LoMX3ESMNyct9mbx32WC8x12IiIIBUfE5NFeDj+
w0PgAqtBPPwQ9khqQS5PHczcvCvpTfHP2f5j8QA+Ku+UXjefBwK1tK9PZ2Yb+p17
UUWLl60t2ITPU8nUE2cnN4RabQz6K6BA7UfjBo+Fy0izgMf0xtIr/gSDP9JaldQl
jmO69lio9J0Kx92rUK+Q5pEjeprYSrZic2yvEH8G3KAF3K8DhNSxg1wzAAw94hb4
sOXG4MivtlLicEMYJywBJNvKacfK+2shii1bO0nZjhEiBrS39AZU+hf0xH/InXQK
AToA7FpOmAK+hRfd03D7IMDm/fiASKg62CNRQho40cemTyj98O1VieZWEH/M9iFH
wkKwlZiGgbFqZDIgkb2fQAF3wz4yTwgSNOshxto/lRfLmR682NCqtZMiZK5FPH1r
OqztNlo8j/Y+Uz5SRBpQinG7XIsXCHeLizc3SJS8w1a77kg3Qcm2/jxfgCEpAdqn
Or0mHyuwcFW3ghqvL2wD5N9w9eCO5MXODLiTd2h+D9ocCfP6++UBXocMxRbztL+L
P6V1IRNJ22WRYjrbEPenzQmu9BT5Ee6CgqimNN7kmI+xtYU7/OhwrWteKdHJ0dva
Wmrv2WZQQ3SKoV9X1q/YFKKeg3ZhP/yQp7pHCro2hprhXpQ7bt+l7DvcH8HmZYKW
ZmBMSlDX1xSViwmqosnRnlvCL8Ihio9xQEXQM4XwuQ17gis1WpxVyJmq7bHsDckD
S0Itx35Y8bHsk4KGQTPr6914uzuD0jbtpWj7PhNPALfCEJPaIb2fabTsS84wYsVS
yMUJg9EuKE+0K/ea/7VZK/mnMobS5VrFZXWo5mX5cnF8NHXsiO0i8obI9fPnxHwM
YkSCreXPbpSeXzLhIeSRHr9gY1mUs48IeqFYtMUyaMdMM67ASmnrbqRdVXS14N8a
Z2y757SYPFILZUUqWnro4UR9zDYdztm/aueH9G0N1AyEo9cR3LrqudUvU/piiVrT
1YyNQwAFb45AVxBJZI5nO4NlnE7a0Ks0U9Yk2jYrnyR9iGiZzQ6zDyy/f9ldogDF
+jR59yvgMYsH1TVBL0J1mO/hGrD7OMs8tYk+QUj4Xrsyv2SAtezfylRD94UXpYrW
92DigIjQOW9XF+N/nclYNFE1osaJLcgUwwHgXQWE/hfbeVysivykA0hPZGvFrhPl
DpJ3Bw79Soe0ghQQDN0S9dsarQx+n36aJZnT+CWMa77GhF/G9ZZcJt5u1m8aZHil
6RgLLBvCneEFcirRCf7/4FevZl9N0aHLMiDyuHp7vm1PhMS1DdlM2lGn0IBiDdIy
CsCVhVRwmBXTktoxF7HMZ0vyfOm8D6WRYoWdi5SJrRky2GdI0LDEKdLNVvpVHGP/
jXvWkeB4e4J4xmKk3Zxad9sGsATljAkG3l1KVwDFQ4vPThFIIs/NS6065CdPHNMw
pRw9odES3DeMTuMhrjF77pLWdY3YxmsNm22WVCRf5uJnGesthlkwAW7MbmCuops3
wtqTSGxi2U1b/39EHXbODQn8f9ZOsiU0VjmsVk3gmENii9GbPKbSRaKIpshxA4JK
ksufE2FBqzqXxV5cBfnUxj1FV3zPVifJVkn3hN6B+HQcRRlFNgH8bnDRbX36EpDu
u4LprUpMhLsf929if64K7PH5S1SN/mi2U/dICvLV+zvy9sAnbX8tT2OPQwMm/RqI
jM5aSIGPS5tP/LvpURgB8n0Hy96fC7ACuLm4NH6qzwnBaJDTEaTtkltLbuSjVQNm
V9ncH/9XhcpOu7KDqCufXEgxku0JAGJVmqJ+FYF+4S7EZdAQ19uQAUkPNorWZmTi
KADiuroCOlmUIyfpLpZfpd0v6KVAAoGarHKpz9vZela11jD0vzAADjVXEOfJt2Wc
Ru6RrbJWfSyLnyrB9YhC7POYfjyHd3KfZVDl28ZtbyW0wl2k5uIvutN7Badpzfjj
PpX4vfSuC6pxF71d+FgdmthOd5KVu7eFF52lyPDlDCeN33kakx8VBht+VnoLmbmZ
9yCxSE72jqPZuZqlWsO32xvp7jLS5gxBs2iDum3pLA/Q52EpQieWDAZ285G+Hggi
Cwbz1Kb9vW9FZbFPEAK86DQ6VTgjIVcmNOXh+Wg6czwaTG1td+dZ6eT05cq5Ledh
qIoTnYi4u02Xgu/x7+NRc34dtuyBtz28g9n/K9Yi0z8KWJ8Yer0b7YnHbTHrDqHy
f4xZkRPWfqqb8od+a1OUF+jqizBTrxJOyGSdJJplmqg4JNFTq3yOm87X4Ss2I7jT
YMDaInakmW94Fsw+IsS1qmXI+JS52FtY2m+LvEpQStvH33RT7VeTx3aILCKtwhvS
xjGTT8BeHW42JQ8k0St67IlyvNrSPitaFY2IpYlso4rMNFTkBg6ktK6NaMcIG1Vb
JKSnCwDeVrzMErTyLkPYjEvfXZyWKTu/bQcXNpIgVv+znN4I+ZZwd820VfQbj4iR
eakfRx/QmYg6Ux4JvMtJGmxCs9INwlFW4q//K4Zwr8D0yh5BMNJ9+oJe5LvVRhot
sg/lS8yPyBLRfzDPuYGDV/8GkjGfh71oe8LBGx9w1GQrMKtQ4AaHB8/gLMG36GXU
RX8zG/kUm4SNgkHpTGGDLgKJssnQVudsZ8njhvVZUV1KeLHTADTmV/eTzQlazyt8
WyYB5B/bIgnUHcFYYaLWqXjcDHz0Hoo4Glvt8AfWYuAp25+S+8+D5yvf8yJW+7Rs
nTIlcOTk3GhaMsNIh2XyUKdWVy0dY+6cyO41P0+V7f3V7tTvqVrA3qni35TtMESr
zQITXvLE3oin25dBWW8aJXIerIaRpUJgwpZKaTl3wBLpLjEkt4BX3OCa/b+bMGY1
vKFXCEmIiqdku84IUTh5UvidtnFAJVusvujX6UnC4qTw01tNX05Qw3v4hX+A+DyM
1aKfnYJ+FrWrmzOTsGzFkpn06nXCfFL3ithbzpi7uD6bEYobnan39o/b84z3JXWk
DTUEC/16mNR9blml/HzRmAqNjZxTzJUwISXldezl4CH6kiHd1rG9W1lGMs0qd3NY
ioqZ24QIaqApfoPaxG6n68dzaSTKNX7imTDnuaS+OvWoxcaa61wX3fo8f1qfb7XE
8ujOXNGRDDA4ZhksSxEHHudZWudr7HW9rVuuspvfcREkSZisqwFyoZ6+fM1rFF3u
DN1DY5jL6UlAhJo+H9iBPYJqlGbrKh9V1dSaqYYl30eQ1vdrlJzYFnf9OYWqYQnH
HkW/rscWJ7Wm+3yWoYp+Jld3oSG+DZEkkofDn/bVb736TQ0QGSPTyMADeq6paF3F
UjYadUnwpvWP5Xacfck6W7vTTn1JK2ISt2f4NyTaVl7vEJumok2R4BaWt77rhiLb
GelrWbHw9fBXkIiN9b95EPwwHJ9orGLHs0RTFnlVTggQiZPF1PTCZPXySOG+P8We
7AEXI4ER/dem/FEGDGyqxHIdv72q3jpN4n7XGvpFEKqt3dDZfgESizl1of2XDMG5
wpapLNwuPsZI9KgUEg9VURlKKYWYMjLBggD+nNVGKiJvT2J0GnQMc2Md7gLV/v9w
QUsZJGaweMhVfkuxeVHR1umI2qYLxgPKQHVKppw3mjIJ5b59pdzYCy24UNFmkp56
N50vCtvKKfuBEUc4GkrObg1I4/0hjVdK+fdT7hZS3KRRO8Q+0HIJiHNxpwGxwXB8
SyjhPm/UEjmGmOUXWI3l9ganIQ7vRnGkg0LIzj26PqfzP5XAXw0NPSbyaDLHiY8K
BV6SrzK2KRKH/2yensafOu5I++iieZHNna1E0dcvJKnaH6YY82ABdviBoJHbjao/
AkUwcDl003iMQz+jGeCxg0v7X7JhqIFWJw7CS7bj3v2+g6QaMuVLQlZAQm5H2Erm
tLX5QY6OQIgHYVMmUHhDBGHleiI9Cz4MJGKKC2RK96DrG1mOCteQx/V9edlqyzc6
ktj3whLas3Zzt0oSrgf4+L6GdQVDXKfkrBxc8Q8A2fyuPa0CoTbFBo/+gxxxCdN2
O0wMUU8JjWbhATXnihfl3F9U8TA3w9xw7xaKRp2/fVvY0RrnTrvDDEd3y7npwqDO
oVsjWyxMMuWnCSu27v1JEV9M0nmWNtlIqB7iTTvtPRTpM5zsEP1DSgOIR1BP2k3/
4s1kM0H6JoklXIbSSpYMlaeRosNb8MvV2MQPLHeP8i70uvn9p1GXwjmJPZvDbO7b
+MMCJ2zSfP3rBc++UHB/CpQc1g/4+xzKb7nJAdsXDiulN/jkhSG5vl8BlLhApiFO
lphflXoaxvZkVGqvez440lkLpIJHyDyjD9GWa5C9B5xiAGJYU9Xq9jL1fQe+2s3w
iV62FvGeuwGSfBVP05y1zWSpwkrdJdALYJ1mlxPSKR28y2DT9WewR+qCndsq6se+
AfTWdRdKGf6Sk/amx9emVLzl0Upbd+kA6kEGjyVvIurBDrAQCl+apYwTS1XZluI8
u7EkC9m2gqzlz6ADhivqiw7dfigiui5av4jjZxjSvLu0Oa2Y3FMzpyCJR/0T9J4r
JfpM9o1Lvi+6PqSkX1k10V+XvsLM/V+ucQuJ7ZU1FV7CIIOurWX/C/D8YLEGEVVj
Dl9Qz0UDwTWG9CFCJnrPdCNPgOmH92ayp1pMQb1Ga+Fi3qdXhpeUrfD2CwlBBllk
8OnajZ/p8zZ1WSTZAyFovM543pzNCoZWYaU0GaBZBSwJ/fFJ0Y9CzI3YNOvt++Pl
zPYq1CmO7Xu6/q/DaQnPXcAOq+SiZVs/57ui9Xl6HUL+ou/AC5GWkZW37UOPDKUI
JuAbgnlV+kQHdDuMG5AMGHEIoLRwbtmiriCmhwvJ0o71uOXIEEvAdxjWjXNmWHRn
l8kUmswzfnt+I2axaFZGd9Gy3t3xYycHIa792k9EPmTNS/2nZGly2Q6Lwwg+gOj4
j6cMY6AQABFHP6GH5kzQgn5xSqtafk0jV4G1j4os0T7zsm6kSo1oQS8Tp1AvXpiX
ZS/VoS3tfKOHiEVN0aw0iO3yDoLnb/A0MP8kwnq/OBceT/VmmP7L7r3EQfJgQ5+9
3A1XK5PK4BQXicR8f5IHGd14pdnAxJQ1OCadVEHKF9lGa1BjpR9u2+IUxXn5ng9A
ZXJDbfK+4vuajoX0xvZRRyybAZN3PDZmWhFAkxNjavSCD3iqeAW12cf9c1sgymIf
D7+nUeOKot9NylhO9bmh40+sNXd7RfqDpPdHh6aISp0Q3mSrVySuUJvhJ6shhmyo
U8wjf2IYG2UaloCU3DnM/FwftqZVAF7cAnEfhYw3N6aofsYZ9jZPX+IAWl3DFb7t
RQ1NaWzykoYvPqGvC08eWVq942GJNp3imEFCqAjLu9eOuaKXTkqAwZkRoU25BQ4W
oaFwLOdLKSOdmozRzPwNO8Zs4cAjuR5vdToKDW7QdiZAScRIcZHOfpTdO0cX6hN4
5Sjs3AwnxGGGgZqBf+qSzSx2XRHFe6ZSUIvb1t/DdLKwZAiAIJxxqA4IhrhyTPVr
zWcvkJ2x4jOYVRCCgnfGtQLZuRm/JBIVXJUBv6uKhvJ1ld4C2Dna0roah1W5fBjC
VNnOx6wjXR7FchCa/8W9ozPcRom+13UL/W7AhyxGOxy6mGk20qrfEwvlsJcO57Ry
ve/+jHHAQtUaTEq5U9uhGfFzvSgXwLyJAxh9gfro4GoakuAB9if4c++2IrZQWCEL
eFqoa09dyK1J2Hl5HKwg7g7M7hkk1fu6aF3Dd/ObLro4VfIw5X6mb/pcwAzxrKWT
GzWgHixwui1zZb9OjXqrpyJpDVVUyR5EqBKkZmK0qikIXY3BIsCVd5qTx13EGcQK
ZhElb8evvd/mID5xKbOIEyDzAkI4b4KA8gdXYSCGKq6kYtflbOu0+3HrkY86IvSU
4lIxfvVBEdNIKmttHjJdNj8pkoVMeAka0355ymTNh5aqmq8cXGmkIPXPa8BQgvM5
zCSZZ5lrUH9YE9FpC9mv+o1fmPed3MSl3liIT9UIsziE6le3UPcUJxSg+kdKlzG2
+ZBxcJ0ZJHks8EdRJY//nqEM808l24BvxQA+brtAmnTrtweh0wqvf77/zdLqqSSf
AO5A+XEy81yJQMhczR9+bCvmcC+FLsAVuPdpI9Bxo4OlzO1YVrTQXCrtum3nt/f9
GCsq2hH4zwPm0j+nv1ZtBC055Mftr01ai46i4b/Gny0Ue6WdPWZY/z51YUvjRZun
60+6azqEPKMbWIb8m8foJ7bXEr9qrs71HvBlGyBIoKdVYRcc/Cft3uzXIIPlcEqq
MJj1r36Lbe4aWXMO2V2yHdOjf+0jQO+gwNoVVw1Reu6WfX31H2422nK1+/7KZ8H6
W2PxDZ9ubEpuqd6040hPZLMCaFHZDThRqYQ2UiIcJ2HnlyIhqeh8L5JlwU0AcW1p
J0fwaxsRjEXsiTkoF/regTTsbibSfGwpIzeYRndVSCIIKhjz2ft5R4zAWn3P4t15
GcVI9Qjt5O1svKlf4mQ9eg1mDHyHwjYRmQjYHzM7PD3Src3IrGmJX3BfEfQA0Bje
32UaXyI08J4lDK1m5ajNSM6VOGG4Uz2LMCisGK8ueectf9n/5NzKKzTYZ6yZjIrQ
Kk2fSDgwHwcqOVRIJLk90LGnfUFEvWJesjGGRQkz95ntXVknRW81LseWbqtALTQh
5g+YVS1bfcOHFRdnnxfnhkuKqLtuOzvPCMtx/U2lFbRQDoGsNdkgVUXLwfyaX+xQ
FUTnAw0siyAU7YnKmJ6d1nCfq6GU5JyjyAa4Onrv13H9dXwwNNvbsnqnCq+RF8f4
9Pemd0qCSi7+vSisxYeb0tvYhdTpFoDDvbu5KDU0weBBCmu2CNvBXOIqTYwHSsyg
gKoZfcHioYkWGMsvZqs/IikQ0j+enA0TjLyKZFGdPE/OL0U8WElG/GhgU5zAoj3M
nHa9iIS7t4okoZh5Fz6UlhvBvB5Ejq4+K3Udx6hf7tNBnXdQu2gxH7S5+AVtpJ4d
5b0BHtUkLnpDGs+qSKMCCzwq/tKsy8kAYrzwafSlG9Wvvz5LXmcX9xne16PDoRMi
bG+RuGut2fj1XnXbCDcoiUgolPXVTXX54r3xSoH21zeQueXRdHvdzgux4+Q9ft6o
xj8wtFt6ROtcIpeWx8SUHXRU95Iiqkqh3zXqtuQeH0fSmPN8HLsNHHEf6Mzg6TuY
Zls2ZvN+cSejShp8Kqh20PNmoNRb21cTdrow1dORCRSQmDnoh/p6Huqx75ihgY+t
nnbWtwniLbdyq7yHr/o0Lv6Y4HzYhu90AG0yR/a+Saw5qPsKtAUbEIbL4kjffTtY
Nfi6bLcffnH6xc2Fr4dhjJmye+SRGvfknscE4i3b2MajieFXTgCjyEAOAguBCHEE
0fh4Z59Zp0d+1kmhcIV0H+ltLo5NM8ZngZEkQbxvq8k4Qt6PPAmW22nGQldaHVgA
FIfVaOYK//pQaZb+DaBxyZNMR9PC4SQIBagftNQt6Zlwr4/ePu/v7eBSa5PmgtxD
TYaTlobB1L1Bj7OLq4Syxu2VnuN8qFXZK8gmPk7jbyu0hNCZS3Yr3tfp7YBIKU6g
5a+zrOc25QvWvwjyKfBShsL4F6ZC1fKh7+jL2wlXETsfSF5etsj+BfxisWj7GVWk
ncvGGF4wx+1dB8dVc476mTnvHFhAvWfm4P9Fy30byGOI4uxaEdMskCLzFTxGjqzN
Vugup2KM3HQFiTA5C8cSPCWDU8L+OmAkOy27zuvHdNcBwX/AURojk4O5TDxi/wio
rcnBm7nYrPzaizZn7qMXFF9XIGrZajZEY5716fcDU2A4hftm8atPN6RZdzb+5Szm
XLWF0lkrmXF5YpE2y7Wx3axPVepHTfWD9k4X0aOHM69/pwY9EUUqHf4qsvPa2SSG
Di6FqbBfxu13La9mS2BbsPnOga0DoTkHVCw5RhkMS2LkpIAqaXNNFO5JE6LuGrVu
sz7iAZ3WTTuHHs/TS+SFVxOzf9HR8rbQJWOw0MfCgF3swqpm2G3Sdy4mjP7jsEy2
MrJQ/v8VQ/fFgs9zxbuv54sZP9DVpYpiyVAbO50/IS4gw2T/Nmw9kkz5caUrUSF0
QEKuiRvW3lZoqVXKEJlgJ0OgaTH6MtwsuKoMJ0m76AJIZuB+upQJjkrZtaSYKgUe
y4iAASNp5767ioFpSYR6ORyCFcglqYXBumm8Zq0NyMJyDa3aGMsUb1eGArOFeZJ9
qOb+onIrbl+iQCGU4/IKk18YTl1CJcJzzgROmT2mBzVEgcL4/B2CObnI7LkqnEhp
q/8jmuxyOTjtTWpk5MCsF57mMPR7acW5dJUS342Qe89VQiAZzya1rjHSlGYeSNKo
hsJbFlG3gLwTjg8+CzcPsvsmcs4F79SD5VguE8CKQrLqNlaEKw/fRncDlaMm7eZx
Ca8BVAngbRm3IAvpmYjWgUwIfo3a2d5HaSNVUulkF+77tYBPr+64m/Yyr6pCy5zr
A/n9p3vu1NkwI1Vf8wWpcPVnQpvColajO0k8r6BDhpn3Y+aP+ciM2p/eUngonPI5
aJ/QXp4NRu625sbbcMYqQgshJOQw1p489HQyEouhjL47O33Dmf9JWBhdmziN510W
zO+enqIPVTEaOQfgwntPE7ughgABxREWE2pz+HvUdXpNP09UDUQXw4FdppZAfJc3
LulO0C9LKyJAiXUj/U750zX43Fnl0A7lv9crsVBQ9mxupyr0XB1STUcv/kzueSlZ
nYUV1cj+yHd1w/ZtAf2DjZTJlaoWUgztPkdIakoG7CNmrd7QA5haWs31DQEqRkyb
7PrxMyVrNp+Dpqz29L1QUZYfCUV5RraRQLWMZcaMjorJKHCtxLXza3JnbVDZu0Fk
bMX+ELep4MbQxJ7s8Iny/QDraZVKRJANiQj63ABURobCVMFE8GhRm208LD33Bez6
kAJBkbCZg6BYjOtpkxeQGP1c5JXCK78e3VRR49LDyI1CKInuJ85XFPQxB4tqjI/4
/tQe+Q6n5WxPvrmwHUFUGGlX/5GGG4p0Tlcphlev+Thh6BpaA62SGhvih15AOG8x
VlAOsC0lJifAmpYBYlEPv6Fn216+Q1WQd1olBqWL+5HAI4R9IlC1JbRjgsWvbk5d
W072EQqK1urlOZuagNbMBZMsSZUVx2IuZyDnFyg2m8yRdKE32SU0uRbMDI540RiF
r1WzPQ2mYsE7ZmFRs8WphkTFGMq6DoY1ocYDwiRojEzEn3k12rfpfX+1YecGd3yM
GXJR2zgrbQDK10nHOO355Z2dXnxLeikGtRrhZSu6aJH0HPNGVVO3wGYlDYQvgOoR
ashocUh2kb/11gjAybbUcQ8yN7kRI4HI/UHcqXkkLa6q8OVMtMn2Nui5LwiVlNua
ljn8ZWzaHIUoWp/LweRqFArHQhmPeIbVGmLZDSVManYsqxGx5bR3Y3LxaWYtnIBY
n6UkOKzYCHFRT8u/ruyykGUqOMPLn0vPKD1WIUZHGgWdQmZIaNOsr03C/l+ERV3g
VleW1XIszadKkJhBD+YxTTOq5PVDQ5JWjo35hvvOEL+wGTJqYgNkep+FIg4Erqyg
MzLjqJPB3RNfIYzp/hL39bu4ucv5z3oilWW0eXljOxw9oQJpJcnEkV+1W9Ksl4Nl
IxpiioBx2aLmzdangaqTavowmsfvuRgDuKkG/7tPjmK+y6c/58mlBzf50VpV2V/p
FW8PlqGS22K8hy6+LRcyFFrQEaTTUx8a1zPduECuOBSX6epERxpucunZxB3gvFWZ
bP3XN/Hw02voCNUKX1JNTiejOZ1ynhIr41ttIHAdUMWA4m0JVMMAUgBQKDl+DjEX
Cjvj6rR6ljdLNHhafDDbYKcfp1/cD50kfGNZrq4pn/BO388HkFMz049VyFWE0ZbI
tTl6vo4Ch3yzBp+Yc7zU8G2g+ItKLs3uHecGI8ScW6wDBtXUua3i6LC9m/5NRHGc
cBv/veLy/sOtK1bvt1d6iWg6P0z/aujqWq7EZA222ZKx5edIROMytPDHM00inpu+
5d+CA+o/SCE4pU8if7AUpsKhUgvW0EoAuaW1VOSFLQnTIq8KpyEXvmVSFeOpNDIZ
GHeDSokQUx7ij4/ZhN+OFQreYQDWj/0aifKII6ArATLm10VTktZmb2gtvlEHSj1W
vrSEAMKqqFqT09QMVEDWD6Mw4MLj1pflQPQeFv5Bmc3YIxFWTQZiIQnKuugezQBU
IFBRw+69KJf03sif3MUb9AwWastSDRVkee6Qo6qWeMc5rJy4W+8YRxFp6V6SL9j1
3aCYpUjf6x9xoyzLzcoagWU5G7ZvxEU/Rya48TkvVqGWMnO5tAcDCAzad+9ZHbxx
eqcRFLgL+1JgPO8LsBx4bFyTieC64G5EyXLBxJmZIoatzaClBHVsclayfme529dA
QyngQXV7RPHSyFtxXAgswCGyujDDREY91gYk/Hw7VcNgdJJINNCMQAWtXP4GCSjC
A8L4cnDHtmSCFEKJFiLM5CwcqYT/NFZPH/p/m+zTNOu9dbw0Kg2jbbVxb/iE3sXz
HI33N0binJheJfbx4imxvq2BgUh36AA90lsdD1wYrfqvyVVkTJnWA+5TETqXnyVV
PK86nN4or/snwZ0zRN+SAJtRVFvpGKm6Wb/1OJwwX/hsZCeUS05UZzIL3ZeKlnAF
btYLGiWic+cb69QtCUy74BarHhmyoEXyN9G7KqqYcpcgU0969RM92R5GEW7U2re/
dFWTs4cWsI/M0sCz+U7q3wjHvVF2ROXdLvd0rEB0HKZCkG6sH2I0niugQSiCYOue
28VC45EXfZC41HnBPaIUgYvjcx+rburNClRII2RPJ4eGOALx6nvKsoUnNAGm9cMQ
HZdYXt1vGU6z1SB7/OcaF9Vt492kV3lO2k97WSpLGEfgU7gfV6sOy3HdVMK//Zoq
2kky98W+5rKpuJOThAzCdJz3BFhxoWwy49XHzlNbibOmEVedDtNCBJq9swYuywkn
/6BNWaTm9QWrvpzqIKxD9hMDHVf5tJzsYMtKHK3bVioQ5yVzcfLB+bXGRNpVAbtJ
+uZ1P37cRfAWpMzV94W+Hvkt5PAQn103lUo5yRZufo8YNhh28F/U+GDc0JesKoKu
ZEJmZwuvtP9n8IRn4+aLC/bftRkKzkC8yBXZOL71Dfk/jSFzKsPlpnKPE2yepq27
XORaxxTT/RJGqXPRJng10tzd5v78I5oiwKmc4TQpx2VvXia/+U70+teEkRKFTfrp
AE8m+Fz6se824YBz2nm+BDamuRGulxtCzCw+k1Q6lbzPR7QttoeGIjUYTre+6nbl
V4l6KsXsYaOpTow3rWe3JlCFIgxGVFmmxgU1e9on+jEBH1pyjunH170GXs1m60TL
mhRq+it0mZxlTPDPf5AvUUYkc/hbMeG24Jz9hFDYKcMjvs4lUXq1Z/G8AwzXa+Ir
W2JhRRHjbJpwIr4f3fN1Mu1bp3f0KVQxdW6Xkw5yKnoJia4bCPeXd6Hxcok+EjZz
0K3+F90hpqbZqBbORsB7ysE3n7PJFa1bjlzI9t5e4sJGdgpAEA41ipmXpKVwVpb2
9zfcFGuRekR4cpMGPW1gjIciZbUECS8Be9t22wBCsTXHqyQmI83eWHSj3hJU6IC/
dGPSvsaD55nYyL1I8LwW/SM4AlCS2od0mCKZX+Q5CINo+x1cabhspQ6sQA9XSEIc
sQFUlFGT50dXRs5vQqWxbaWgmfaVZdrWQIcfNONpUmjbv8eJMFClNVCOpQyDuFvy
mhW6GuA3HHt/1Lugbhu3zeTdISOF/Zm9/S7IDBxiGLSQlI19sKS8icTlYtkQ2L2y
DwVAdK+sU12Pu+JSWErAnok3gN+iOwtt2+5SvedkxFcJZYZTcsJ76tTI/sGcpj3y
X6gW90sEm1IteIgceX8whg0ges+nZVqI4yxMs/SDMcrRi8dhKLpI64cmhcYJC3hY
/A9VCseu+y8mI0NlB6IMGcr2hD5i4V+qpDWhjEVdvTeh2Hyuzzo6zl+cAe79AXP1
YgvWXmXLonGH/G86FMyCT0MAZTOIaemH6ndr0w0unmS3sHm+EL5hV/oOV9RkrMWX
1Ilx6Ddk38nEOEd+UJnV72Pm2zWndDzDoxhMWliy8da+DBHhXnnw2Tv6bw3ftlF+
0K/RyPBPLVumSUF2ljtfmEpJPWiG9YZZQN5aciB5EbD7o1ak80NrzRrjd95BUwn1
wL8p6gIU/18oMrIZMVHt2m2YMfUkD/ZQ8bMZ/gWLCXrK0ECfTnPPU62UR14ybrYg
D3E99cnom/oAxyfrsWfUnSxNT6IT2ix9aB36BkLqToxDQDYfwaFIUi4EkeYDHmZ8
QEPvS7s98mTHCmBBWsc7WIpDKE9dQgih3l0e53KD8Ucs+vYQmnQofrsBV0zm+0jF
mpukMyX52bULLeS/v5DHPFYIuzNljzSU7kQ6XbQ0qjklASB2sQp4ymE89nmqrN2/
+9Y6tMjYVLTCM3c3uQbwKw9jNN/+qMahPrwPhGKe9C/JKnYtbioX4iyPjdbfwBab
/xxweXPEjZiuZf13slxFM/6kclBRLvBWqkuA0SzkDp/zLGOM5kJKfOff4RWfd6CE
b6nZo9juhXqj9sFhkCbX940unWI4bw50/BgTCE76vGJqwQnlM6/hw6QfdIwH4GwS
Z83vYEk4E7tu6uw6hBM3s2ZYFHek2c7RLN0T2RUlioLJtrKbDwTJbKvypIfuDIwn
VgMtz9UDF5FFNEtsKjYUZid66oAXAm+SYYOwz2Hl7uTYk/9W9svpWw43+FyEt7DH
XDZ8PAD4SvpVoBur/R4HTz3w39iGEz8IBtI6RBxLZecD9JLtnsS0mtHUNa7On/5r
tCvqozY5Oxkd1LPbfnRjLc9JzsxfTTS0xBi5jK9WfrN6WXOK2Qx8sXAJW1rLQ7iI
R/ecXa8dz/bWls7YBsk531BMhSqwcjzd9MNJUXrX4Wg5K4u7t36jcODyndUv21bH
RYgj4nHC4TG6+dKNfg/7eGXWHJZcinbS9Ac7IQuUECsfYpOPx4MwJ+R9KTfQmWOY
T4DIMJi5D8WEaABsr2xsAeYHIrZiPs+VCUnNTRKwd6NtJcKXNvRm2bI3jKadwQCv
rFmqeg2Bmy8HFY8sqGZR8gVG5y4dx+hpdlZbJ7Iscjst2PbloFzhMqN6OuAfEATA
SjFmspez51i87hRARSt+tkG50gxl8i7hfoLbkJ/iUb4CItZ3zCeGQzsUtb0ApmMO
ayA2Jfauuk+MjyN9E5J+uugvE03gbvsaog64qLa7g/+2YwpptDmiESBxINvaKWOx
P+nxlXiCmZIWHr5X/B222nSUhkWO6frmBjCJcxwkAgjXO4JJ93ZIoLqccioj/pFW
HemTd9y2QtNTPJZLKdYiTNm2cOfanqvjya1IDt8J8UDp/IK410nKvAqymZSZe2oG
llc1bfR+4Eqlr8r6e0XJtdqeaG/3sUFalrwyCMDK9E1uOY0Qn8T/smBbSRQIcF0R
VaNNUGRsVQeIUwi/+G+oT5ztCa4H5J664l8qelQ11e1RBRzZi+osNlVjSwUAJUrr
4TLqlanOn2O/dJsWSQ85fWwjRTz1zM0djbvbz0LfJciOxuZ2n5YSKcJf16jPEvod
wgt4+8ShQqnltrDw3u5qLAZZMmcBHZcWRLny6FpJzK6p79ugrOFU2bvJbYzQnsOq
O99xC8VTho5pxh28G4I1n0vlO5ec0AUV8tPMx3QU8zq04shZFElX9qt6NxZ4IS33
dM02iWXjEFru8+EJh/OpGH+bCf35yXkAsBISNDe9m/ccXHeg7YvmE65ldn7hr2O0
F3gPPGpe9eiA3ieSEoSy2451YNQlbhvR8QCKbwxMeVqMSwQ2lRNzCLCImos7xRrl
TO5HV/mmv7mLCuiYx2dA9uW3+sre7zA48Xkzyss1dfqv0WC1s1Rvze5jy08OakhS
NvATDiMpc/az+14sk+wCc1w4iBMjUa3+HCe4lGuVENvWccipaRj65mxbh5WdRE9i
EXeqIl/BrdVGF3+fGAWKqGCe7yxpMVBURmkp/v9cI9BedhnvHm25dQtkdLcWTiI4
TlNJvTrYuPFeqifWhs4iKymaB2yhzTTF5rmR/u0bFwCAEnfAT1Tg5Bb2o/iqfxZ3
R3rEeFRJlh8K+Lap4EldFETHEAKaxUrKOkWAAo44b2zZOXp2jwf9cEte5eQlDyNM
OAQ+k4N4GuVvTM/4iKG/RDgLqfV+BPBVePon2UflhmcD9mOrH6X/ueT4mBk7noVy
MObEWCcYyL4B8+JyByk0yejbxN6+5mh4XvT7Yaztv0wH6DG2iWku/ruyjGTF2s1q
lb6S/v4zQoUSEg7qQ3NHCSaHnIWGSLHBA69bVaJNwRb6U/pudeFbsFv34ps5/8Lz
GzwCtYTnCEzMU2pPl8DCBPIm64ND5T4sYILDK4kAPxZwg6S445P0aKg+m+kZToZW
tpgCnwmzbWKmpC3p8HBYqQj4WvqNGv0ShaQR9S7AYPGWnD6r2DiynMIuT+JNNGmw
iFy8jaYVaJjL5KToHlTDSyyGRZVTPil/YFrElhU8tzGqo6Pgy7Aeph7s4zTmUkT3
dERvJs5bInz0xyL7oGZXY/Q3O5dA4/3dghIbpMkXH+9F2PYC8YKECRSSLfDlDO0J
5RMk8OqTF5IeJisZz1iZ+SmHiwAQCiygzpGOwOEcGACdOD4ajO4F4+QghizC2g7g
hHZHa3qqXS25lsdpHnNSHS0MGWamSX6OM8RLGHnLnfeenpd6bxFe3zpzy3R2h7SG
rLoe9843rVThD9DfX4V5p2s+uAcxlzqOWiUeS4tao/tCtFbS+O4hgHKFUu42QcVj
b64HZd7dP3cofMPtd4G/zTCxh74ri8K+SYFxiQ6PCFDQN4L0SotI09JR+s0zNJJp
jQiXO4J7F5+UTyh1UxbzttHjhwqf6eQhZaLGNZSAUiITR/U0umRyaDdCGNt/dfbi
+lz1WJiuQQc0qeNjxdMM60TCW+qNvUYXa5bT8KQgBrG1Eiim+PhEKQ1s5knIquIn
ZKjqF7/4MUv6FjP2yU/+OzETtoMP3pUC65TdRM2qDy8lCMeH/T805lPUN6E7lKtO
NsaIp77Vdsw21ROGs2Kzj7HAMTHq5IwQX02EAyfhXe2XljZvd68zxivDzf+aKS/U
cFNU28CbwCRo0HJfMAeYA4dg4ayVovH6RGyDFC52UcT3PW2I9E0UH7itWFscNzh+
4JsoLZ7pDwW+LgczA/67/cm1KOhNgADgrQ9AUhcZm/tO/AzXRMGPh4df6Kxd3rRm
/J7j/TD4FgnR0LZytA4vtY8nqe6e2VCgqJcxPKY+xvWL48n74hWtQlT6V5mz3p5i
pb524S4FSeaIQJdtmPuGFlUU9r7CBWvrlSa/ovTE1/2LKjNKnWMHPsY54lD0ahgi
961xvLMRkixgHfCjVXGHIAT/huVfehXu9mdkOcB/b30xxWaxov3+5RRNdP8Evzuq
7DnLH9sIUx9M5BT2hEyuLCXjj5mTT+eKmSCnoRkx7RacUi26TVV1PoVChDG6yNjL
tF7dCKxpHvhlO56f1C+4YQnB/m/xjsLb7aY9OcFag1/QBg10J7o7cN+LmwHzp5DY
DwZOnqM76UWBRm+pbcipZyWoOKp/fygqNsipKnnOeiy3wMC8wGfi+lW8U7jD/Sn6
7WxJHc/5qosqLVd+DpNiEPTgT5bQQ5UCXowkTWHTlx/ULwh+CuFT3CYLp6pdE929
Hz1kO4/8LauFvmnE5CUZp2rYGwBfUUZNggTLTP+v5EtBmNJWUI+0+xhtGkn3CjkW
W+YdZmDcuay+evwvfWFH6qTm6JtPiYwslezQUex9C5mH+L1IBGFEfMqZgCQ4MG20
R+3zIBYJtmVNqiR3s1FRf1F/Qc0khhC3eDiFArOAl5jFZk3u6BOXLahwAQMWATGf
kdYe38t3SKVyDpNHimMPzJiyReZc8i8BJMignpROBj2yi/2WWM0ozU5wNzlYWItY
i0azDk5JGD7Pzxh0dytZGaRGDRVYGoeaMAz3ikMRgCEJ4eofVAtUymwszx7YCrjZ
Yk3sK7EHsyy/6/Pt9SZALFFH1qLNj9YvCDNbnyIiQMYSlb5KmreQr7xyh9WF+jK3
22uFP6mA0lWol0Q/yx1Q1K1iac93Azy2ZlnXGE9+Q54KqWSUU9OY/KzE11XYVupp
gqjvE1ngp4iMp8L5LPZIf1X5oDuZP0rk8lufw2gnvhPYks1zdEZbKWYRkRPKACxq
hbBuXY26+Ik68C8w56up2MvWrw80eqJWTz8vtmeA+g1z90120PlHOLI43gRE8fsp
85983Ue9JmqrfVNrdqDyF5xGLr+POetskiBhhWx+Z1RHh+i4mLx7CH6kVyX70nxN
TDDn8LEfstl81HIsFZ7o+F28mhAjM/xDSski32bhN+68HSQzAc5POcniCUoQG7xQ
Oa+zbkk1PMxpUZBjwg6L8bFs9nh4Fej4FZ9x0ftk7tsdRbQHi//ZdEoMwnKseClK
RH9IKiYWxeN2FIb5qq7Jd4k25522Z8FrILCjJXLBzZt4EY62HBNpkTHSGvSdJC11
zI1dVG/BE+N9zzL8KT3gvZ0XWo4bjw9zcjNt1c9ZPJYonudB5VSU0ZjlFxghcRsC
ekDpV8J62fOBCXLv6m2SL14IbRRE9xSKmWrSorXKlYESnEa0+Mfb5vajvVtaO95t
WLjty/LIBmeT7NeHyjPDpJwv+Erp3X0qTf4ouA0o0zMePwuqsm7UkNFlzJE0ITzT
t3cR/StX9fiKi9uS3ChfnwgCIID1OjMfRnyPq+IjwkxX+tWv9cIcX2kXS4VKqRLt
AA4W+1e2b5DAoU63hfQbQCGbTYhk2y/4CL4taHmPKpid1ZnvR6+ZxED8JoBi1sXU
5vALwwf75OQdXn9pK8ENBnM+EqoBoe44wZSS+gEthXXComTU7dAWnZQZ85G3ZHsz
lY3pM2cuhZOB0FmtF0c5CqZ5aIds4npSxm4pAFQ4o7exAGqIFrisqv3548tEvtq+
J2f+uANWmBb3xSuu6oc7wzh5lPpZBQzBoR71VdHb+/I3M5Jp2pM8yeoGLZENcH8v
foE/ks1ZjDriyz95dcuk0ADwbac4TNkSF8RisLED8bH6xw2tuavHfxyp/Hq54i1t
ei3po7YyNlTqiU7lv6PnYkhxldNEB9tUlTlmjJgn4C6h9pf9cdXE8Z0l2JzQB8jg
u5AT1VUvy+6eHkXy0X8VpnTL6yXx+stO3gR2kLZaKFFHQ4xJi+gHQMslCPz6y/Hq
7K/FMEtCgu6/a2HCeCUr1VsOWfok7aA/zRGLP7rcAN8MEjCqh93Rjn5hB/tKEmwb
vRI/bYh7fvTOnl4E9wMtSr17b072iwRwFpZ44bSGGMM7GSdjOgrWSD9XSByLhAOI
zFA5HuaS9Ha3/ih5nRUB33p7BIVl48mAuqf6J5bbv3GoYl3Xeqr54Jg3Cn0zBweS
q8e5sbPFtQNxrLgBIykXUUiVmPB9WO4J1V+7Cvgdt2H7ORnfG4jMO5lg+lZmf0CU
nNqFOSZsOb0DsOWfdsrQ+NAvgAqOuOH5OsX0EwJnzhQOdLbYQiI10JIEumjPPtp8
6nFvv+uyWSliWZUw1YqxjD+TVbt+cXHW7rqNU/NidF7RI04os0kcpKjhLc1uNmY3
1YkiLnYyg+oumd0SK37buucFqSVML2jQAh0p0+LZ/PvCg58o4yEEzaPC9Qrf09KC
lpr76N1Suzr0S8+fKXGPh700LrQe7tLC0lPE9AihRcHhbvfClHnZOziuRBvT0LFd
xF+IRPj9gRX9sInhc2CRfDG06/rQYK+M8qQGRQZjsbkE6aYwoZcbN1eGUmse4uwk
i9/9Hgb7JvorUIEk1CXXwN/SFP9ZePfbtgFAIPCvMcNsq4eqLmqExoDOKZfZwK4V
kq3otmAFNRyXksai6uBV31zc9ynos4QteCp2P3NtqiKwLFe+46w/23A+m00QdScX
y2NIF/BoP0TIkOAdGnsnMd4on1RRQjB/IY2Um1KPlMeIn+wiFJXXZQ0VEacPyTap
M3axVlQ+pW1Yjc52/dC7fcQ4AhnBeTs+Jdt6RKzhzndp18egQYoDm/0V8RQmubYW
Fc3TVRh/ZGxidGgzt8uawd5+LwHIYaepBKbkSoOqJUHI4cLkX+Hdm1inBJFNpX/h
mXMGI86Mi3TxAhJMf1uuf/+TXGvhkMOsuqr3jgybIKGew/TqnJvdupT5IxgPlbhC
vSdM+9/74p60N8l7FG0PN5IeSl1v5V0L2D931LGjHJ3hy1jH3WGj2uoQlTRvdcOx
xhx6dbvFcTj3sf1cpKIyyzKIAmYSl6ZhfDFnimu5uG5SN9gNRC3EteBi598a9Ewx
l0/udgTnwPJNeMcNZaA0Bql5dVSVG3k5EI9dcUKRXI/lT6EClQ/V2q+mPk41WWH2
IbgvYUFdFUyQx484/Paag/Z9OtZ7G002+GBh2MyLX6KxIqyqRDvLYezbgdXnQp2w
If702pA14f4TFzUJcc2DuKASG2TzRIx9vhzJRfSHFPmme72GzML4aPZB9KM7ZxYo
KU52lSC/qp+aY5soR5zMtmGU4BY1yoo6NS7voectt5vXL3HvqxXOrvjnfi/Im7tB
7Kq5ho/KPt5+3KFfhVa8hOfs7LgmXkb6IRyhWc7WUa5w9dBz419rH/BWGYUjJE/7
0KgLA7hLnKeBGfjCbnQfM8OGWVBVAdfYgjlngXGYr0MspJWMfW3RL5+2Ok967Uwr
WJUnhNUMPbMU1MNNfgMiICLkQXYoL/K3PR+xGjv2w3kS0dROj2eEmGFuj2KFHQea
KOMhuRZdmYy1hzyJNl1nOapbveBfiPVgJzVsnjYF8mNygnlhnWUC8XgZgvQvNoA+
vRtIqoAd5o9uKAROBU5J6XVqAHnFME0nqeaj0a6rAkZmPRDkg0spHVhb477TLraR
b+uRqw6OBmEhISXfoj0yxhPB/O4pWLWfINi/RL17Jg8P574syXMLjo7+esrqM5hn
qOtQLH+wG+sSztCQPhln8Z/fwCewXCume0AlV/7vaYX+O0TMO1DWXcSp6Wi4Wdvq
TADLKHSbyGcwi7R5dbb1G9oxOzOLuXZU8ctgudaJkp392st5A+uhyO27yX2/Xx72
G2t+mp9O+hIF4/SBq3svNnR6931ugfdu8N6wj3wGMtIeFg/qkOby8joXllx+kCh1
ljakedMi015Iyo1j9y9fx0+J09O3wsCqlXpNl5BBAVtHb5eRAVzubrjmJ9G330LI
VNfo4Tk4Harb9MAY+VLwnatzfVWptxkWWU+hgXJ6cwu6670Cl6ZMUf8L1gfYxSOX
9YoOU0uSqmk5+eq3HrxTAfJL7cYp74fPYLwNsU2eGULVEfXbGmcaOT2jlkANYDWq
9WXaYUPYsDkybk0mTAhqZIOn48JMO5t9cqiKmoZVLZOesf6PUclNkFc31WGMp0jS
KQCEHn4AOvAw86qwdsQx6LRMi4tVjA/azT38I5oXWIdH2x1RVbvaByq/KItp5/X+
yK3jXZS3tHI3Ho5mX9+esXP1LHXNZ48yIDlMfasxTvchAMfYkHMnQkK61h0zPgmp
CRBk+WqVMyzqCER/OJsLmp/YEoCYCtnb5Wbjg4DJGQ6I2T1LOwxx1R1JVgqpWeYb
85kZJSVkhB//+jpbEQXz3Z9ojOWXoNH0Lc6OyeQlsrFNuoCtDee4Nz9aiyggX/e/
Pj8WbTnDnIDCVWtU673fw+jzme2oG9FblB8i6vyXWlKMD9BbTeKJ+d4GwItHEMW/
B2yu50Nl42Fle7T5U//+UZRu2cAz3kR79LFaJzFEJaXoaMjiWQH+WRXfRgMwFGpM
wwE7DfjGNo3dQKcuRJs4tWvYZgkXdZFQu55LMcWwsbnpXRnb0oXVKdW+C3sGl5AU
oH6+54dil5FVXh6iWj6hZtfonZAUVU9N1bv4SsKhI76bLtVCTfnn+EIi5A/rvhPU
oXwAvLkK3DFH1og4RE44arSoWfzpfx9up08cXmBmJL0xU4nayANhN7Iu8vX9MUCz
6h1buXEPkDOvxfDSpbaPH3tbKSWOHOFFBozHlS70VzzXOfh32sGhM9ca3F2F72vB
Q9gK6Q6kv031t8g/CgfJZD6gEdOfPFz++NMoKUFa3VlM5mtnMXYY6m+VprKpaHnw
8C4Ey9k/bbm8uZLu5gu+LWx1tT9LBlugwph09/nxE7GyLH9XMyCZkzwvH5QeR7Qg
8nB4HlStHXSlnPTwKvZJyGQ21p2JZhH10qGBWcHwytEmncnJrdWiZQK7jN5tmwN8
88JHp1ALU48SNgMkIpyJsNPWXtC1WijEDaNjLFbpPLgyOrz/ItAfMyxJKcaSFQIp
BN1RwWI/2EXMonji1QOOvdgZ6xhoWCceOuCIsPLc7hsKlBIQMzaD7JZxJWhJYUaO
9jbiLT/gZWvErldkl4/Kb0tOyRT3Fk2YcRK3EYwDEWKVXy26MyDtwbyGiaCHaJBk
p/bI3U9eIhbY+amyj9HcyyolvTsdNzME8aRbLNbIMakwlKKKwURPA9JcEZppzehX
zWV0uOhx/pOhKvhui1+JAmKz+vxGjn0A4ZgroYmgUvbA1QL85GWFndydweP0Hw+G
5KSb6ASDWwrtGYrNNMWn/WptStfU3DBw2ieA3AxU42uCTfjdWzFsNyVaXfu0XX5G
6HSl7kJG3mIGWJfXwkicHUFLUS/I1OB8fSnOZjrT39e72QiThin+su39CyVzSJij
vTtpUY5W5QzetWx7slVJ3ePFzmsWqcKVmmfepXttMPC/r1av5bb0i9/jsSMxwhmP
JKFfEqpPH4YjJf5mRRZV3IzU/UL6XsXDtoV9phtJYwKhBI141lR4GvP5MnFhCdFu
rMXHtKTsFditOq+7GfF5mHnuqSoLR3rz4z13vdR7x2vpaNuCFyBvEZfNkB383v2d
PaFnkvY0bGxRYN5vR5AuFQDM6QFuq5qC/jexj9041Ah3tEsON8XSuCfyLtYYismc
lHb/z/ujAbzo4H77A3TYzKQgR2acS5bt2YEZ8IKQ8Ec+dXPsmSR84CbYYf2GeWWS
cuvT4wfRqQscQRnT6QVoy6EfejbhMtCAgBjLF/EeZ/AhgfFq5cn87CXf89ZWFS/L
5nK1KcOOonegPGQ4brxXIedIF+Zlr/LEKFnGgGNbXOIkJIAsGlfSkyhl8nqGTmot
p/e0dWbCBmohDfN9BvWNcpKQqWUpPRZWHAUj6KHznsA7IhoY1hvZTBf3PVdQ1QW0
j8uU0XGHpwjcknt4Jk//p0XT3f/21JNfTw9jBpybpOP2awC/OdILjp21nJzg5eDU
RMoomAYKh9OaEiaEeuEwFX/MM85USGawvgJ21XHdZ9C0kQG4XUnB5L6LM2aFove9
NGsExT3hM02UvHM0hhm76uArqnhtFKkckR+Xf9jmBflAOR8dC/cOjCLOrcvhrYtB
FLuT6Pnbqy6x5M2JLt8lpW/e5IXvw/T/CpnNzXGUUxlpinwe+qOBs8yacV2IRexS
O74WJqBmg0Ygw2z3kURMzdXKJsQFVqbhVr1nMSinhL+ArUk08xZ3LjM8SXEuzJTu
s+Dpp4IB2fFFKEhP8E77FMZ8B2tDiXelNJ8a2A8kKT1DrQBQi6lEHVGY+mpdaC8F
jyRpwTBwSPk6FywM4GfgwJSvw7vOZYVM8cFGHDMBsU04CEm3xxz0qRRXMhmMEa6D
l7ADyKEQLS5G5fZjAt8Zx/7D7CnXp3D0wtI1OWo5mQR6HqdmpZ1qNY7yKvQbxasB
I5G7rSplYjw+Iwk0Wo/3OTZ8XNyQyc6EnwIJDTXMAPMqPDHKZfnn2lIDf1pjX2Nh
+mAvJQkQPq2NSRyQ14p3uoXbGYX2Y56jlyoPFjN1/T7OOXs1nDgC0ea2MMRuC3+h
ym266rgZGf6jELKdb7x0o0MJsQaP4oB9AbxXuM9YgMlJCB695PssbCrZTIiCnU24
ZIlFLwgdafjd56BNxsBu2M9/nZoJkigh0HmU3C23nPBKuxrY8M2RcEG0vMkwXW5U
itqrzL9x9gsYhPuTicGjYGsN3cniFeVIkq3MDofg1ZXGEjpULh35Wu4c41Qqjwwr
9UGwrTG0TeaqY7kDtwu45WKclR0eLeuQ3YmwtpE18flZzhSmjJAdNchihADe5vLv
pZkLbyt1ijYGFucgSUyAbNBI+R33gDJ5biygbNsz0HPnr2iVkfn2lPQhFhf2vEEW
zHCqfJIP9poVumN2HkoypS9sswwRSYftTCjLjU7v9AyY7tdD6wICl0QT70wBX1WN
IxbLRxScX48r1QcRe+p9UJpIyXqcpyShj7Bys5VLBudImV9lVKnjr4GlbNNBP8xU
xs648lK6h9HNPwODoo7oeibVLR3YCX1+s8UErG8aOLWttobhC2xkYb8hhtrFjGlx
QZjEukTGEzqB2KOdxj9otMNSOcTcV2bdM5m2Lunm4tbwvbB5VxunaqR+B8DXOYVk
kuPwsoZaqhyBNJRmjjjqBItO9kd+4tlvOViwPjYTf/8JHzNGsv8EWkIp5R40ITLt
blEjz/z3y+ItqSNYKVgPznec1wKzdVI0FyEANVpSM7bu72iahUvhSaRhklt3fKNV
rwcjR0UChJ1rOnfwDWoEyHIus7z2mL0Ji4I8JcYFRUaaxgCoPEHRnXuUjzsgG3iz
FjneN467Lu/PnSy0zb2QNMPjhMU36S0+nFZORZpCuMIUXGP57Hv13M6IVZnQHWXR
iYGdT2WlWb1lS8ZRtHd/N4Nr4hJsWuawWqUSUSJ9715lG8vv9uhg3RSJdNs/GXDE
dLdHK5eCOjdtvDekiAQzhCKSL/xozUuAGgUm38ZwQLX4Qni4fRT1x/QwDwrUm0Yx
Ok8wus+fPk+s/sMkMXZPUs2VvtUpLutHNu+ZYPbSResIprdrTvdhezIZp4KUWOrF
RT6uiv/OZVPhE9hYX8wsKEuXaBwa/480Y42JFLBBmb9a/ivVP58Hx7G+VPLCivz1
2w0jgsZfLb78/7b4rl+CX/AB1kMzyiSITApxwQE95QvO6o2ffNFSZ9vv1ZXoZC2/
5J0GH5ZQodZF7pHyHq4/jyCdxf9oGTdOUDMCr9YRrkZycIzZPh6KaJdEdKvnjr2k
fdQkgcIiLTDbMXGwmEBy1pbsMUHkBB5AuhxaobrwyKpAlsLdRMnV6ysMw4WBps4k
Emyfaw4zXxtlo8a3W0ZmxPatJ/S1MlVIXQ6qi3gQ8bFG+HSs31xUxYUHxucQhS+a
AQsrHK69xKZLiVoEd4wPNcaapvGmoG2pbQkNlYpYGN0i2zItJiO/4DqPNMLKlF/B
NpmnIH5oMRaKzLlsyM3+mS9JnaNyTWuMlflHhmizYxnb0aOy3FhapzCSH0CLXhFp
s9c+Ko557VWy8SAFaoOys0L9sgPO9ww1wCC2v5hlaH1eTaZ4a4eQQdolUdkOgcjP
WYShWf0TDIHIbENCvYaBuG5NhHQsDcMUrM5UJpAu9siONM8oplotT0sgQuD3RCiZ
exWylohXBNa/RMcl/m4rwmP0YBqDLk5MwqZKDT5jKfLiJIRpF7EKFDKOFthAKwiZ
/jyjHH/x8IYi26OQnC73PBTgXGd/urSnJD80iRpTZdd+BtX/zkEBcHWxynjkd6Vr
oMEKhpI2tShdW47XQe3AiV76AV5D5Eg1gKy5IvvYxEUFg0K/InHL20W37NvMiasl
Bj/dhSQmYbYc6IKUgE91rqWlsSrk669yuaLvW2ERwIsyBtO28tWPB5pQ7Iw7FeFu
L/PC4skysQ2qEo66+IUK6E6B4YWmjDieTzYUTOzNDBkdQ0AHKC7DE6Jq1k5V3PBs
qZc+uSpNEfKtqTQIOqYPtxuyI0aP0sKjC1CI4tlomDRuJN20T8lC/fZ5hcmsW9RD
UaK1yS+FCeZKm9BAbf3ZTDNulIZ7KL7GBYB9agrMSebjVjWZy1Qgp7dgYhhIOtcv
fwjuP9j916yRbS7SV8epKwTxmBVFKzLez+UduROTo9MpQAjqdHy3PrOVQ0Gi8dkY
6ty3bjxDTpy358yXcYxQenSYGU08JWtRuFN8XGkasxTtCl5qgE41QPciVrwkLSXY
WbbaC6C92aY5v6mdzuPXIxx7gZCgMOhEKkOqzfaPzVRTyLnDxmzLIrar3MM27m76
PZ5wufX0HSIlzBoahdAePM7eSzCt+EbHFwDOp3c63YvN4jaeDXAGpMS3AMviE1Lo
HGslmte+I8mWkbpYqKUw2nssIdF/P1genEDsdZiiqXAo3+2DHX+IEQY3mNEqNZtb
wZSoRq4xHP2FUh5Wgf0n13g5nL7+CuQNnp2HHIWUsXPPvAi7E/D0nWq4fUEZXHgP
4/w9O5y2G2u8p2gTObgM0B5szI/ZV2CqoSTOgZElnX5qoTWMarGRgXJfRK7IljTC
dZrfKhckOh8E6Z4EfTZ4gZU6WjzPPMVOjynlZ3tabAuFlXqkPvZ0hXUT929Wkzz/
GJ76xnplS4M6Wdr0yU+nh00Y+43IS+fWqBZPMtO4DoekShr32vCY97hHZoOmYoyP
/f9cyRgTL9S441TK7ga7aus36NnAKtllJMH3rB+lgdiaLSHMHldLm3wtfSvuO5lF
Stwa3J1J/vdb50SWMvRYD+lbcvJGZyI7qIzhLzxjODOyCezpiV7JTgtftNyLb9wx
fmP0nI9/N71JlrmTVgMIQ7WZBK0y8S21ZWEYiSZ8GOURA3pl91dKSeUmM7NzGGGp
HGMWqc/rZQ+9A71isub/unS/FkifToxVT+n8qvqHXZXcgGuMuACb8Qss5VfFbic3
CBGwkGINGYeAGqDEVyLvYGWcnVIb8Yl5SsCIjzat3pEpKfYcMHA9YWMQvP7hNB+h
HKNG8zTX8OdN54RsFdPalTcD0/URELBSLeV87Yh1MliSqKqaJ2CHHFPDVy2AZDC6
+MLifc81iEtOFzJG6ug0NsqvXflfpe0NevD/qqaUYAkTDd7g62yAyg2zDSUe0px9
TD8fTjdNDx36GonWt425Nly/CULfvqB4TJ/k1/Vo/Sm9hOZTB9z0RBONm8T4csCt
HGfoBroBqBNXDqJkMiMpvDf8JC52JlVBuLtnqhAM0YOr5Z/Gwz7FraaWToj8/3D9
S9scSzgbpg+KY4b/6J2Ck5d2sO/6FKKEVTVVKHCp7HGxfusRoPR2bAtqc0Ouct0m
PZg00zffGL8zAECnhyx43m7Uf/ZaZXnuKjAelyEl6tGSCppt0hMHWJFBkbi9bxXq
NQojHIgzW/YCsNPlXyWgxkvXRsq3Y6vD5KnKWRJGsUpa8gvTxt83l8NyxVQdnUG6
T8+hb0SOY01DJukD8qX7whw8vFiLR3VhCZ+KONSKVd+Gj5qIZjnAbaxPEHwYwMq4
4H0O0/wVaFHofhrV/vpAlC51zQFJAog0o1NZBgoEBvaOofbFqifxRtijuNXrUXqI
zc+LS4G+mpXHVbryMnBcTzowDmb4jPVooMFkJDbEdMQSCUPj3lxeP0WD6VWY2xpP
yzIA+mnc6ACaIRhu3/CUOPyjrk7oetk5D/BfTLvkM0RXAIPa0onybXGIbyXc9s8C
nndvOL+MLkwhmWcEoCcn2AT058eaf/2eE2fJ1YWqOPp0x36zyJux5Qk17w4JfMF7
DAuxldZoOfqpnpW0t3zzZjp3ZOvOu1kVjD/kyKGpAPRk0JaDnizAbYyIaLqP6NvP
AlHGIZ/hnnhymn+pVdFoO8nquJJmy6BEIMe0EsdFhXPvdFhtAporZ9OQyZQXbBIO
ayWU+FjOHC/zLJjaZXTBLT3ywLJGQhfEDQB2yVeusWVpF+DGuHqJ1XZ5cyAn4ZR7
NNUjIiLQGq7NDPEdvpLPepIMwsFVWwJWF6Prg1WdO16jFLxJwfZ+OYpGG/tgCIH7
wio5h9cpcUaAyIUPcU+2Mm2agfWCwaZXXs6kLCzCb/ju38irn3vp126X0As21rnk
35tDsD8uSgVtWsm681v7LVRhgkrpx31ZGI1yjAvDozM1kqWaj5MR2NsEu0/mvAtK
mqQef5knY+tFVziROKdFfSGZhtJLnioj3zndikyuE/ndiTitXPBLx6Li9l4lUCdr
Fc9RMBITuimBgN+z1/0ZXl8vLcgK3Y9BqGrZKGfBsDn2uO7pqXLiff3PDjR6/kSL
NeGQ1+K+1rfKZbym/WmyOr0LZtaU57P3uDXNZeG1ktkyma9AMdFA8wQT+mcKb/NS
vG2Obp4nOGtbOZf8VQ2tP3IGPeVMi6dhOj0a4kyuO7Jk3MZwUem+rQgqg0BQNn5N
d+nym48S7MO5ZI5wMMGVBCt2Ivss9OH8fH0PHWQA76US/yWeNL+KJYI1Mrn6iDcx
7ebSrxp3+RS1eYf/J+6ZE5ueDtsHuU8esxQPWhpnjMJtUYU3YlQ1tjvpwm7YlzZ7
4nYbkTR+6IxGknEb2++HwM1mOjlW4WIWzFiNLX5PDiIqEpv/I8p9m8OqK/T0q2rf
wO+yy4ffJxxypGCmHccAIl0XpFzT5RZgNwaxMbYOnjdxaGOd3YRWhg++QAwI5Pdu
crJZQ7aZDCJ0L6LP6p4hjprcpmrDvwG3iipUel3jKm1NfP10q1dLgh4hrr9Wui5h
nToTAiIfZ0Qk2g6264HF5GSFW2Hy0hXTNe4/wDqTa9SdS5eCj/kc2OC0MgfZ8OA9
9FY7YsChuD7SmpoQ3rH+ErVIN4SnJCrmKQ7pz9L5LfB+tpi/R8CGvWyAMjZXhzqh
Qfic+I5jGJfe+G+imam27kS4t2WCD19CURmiRVxF79M09v3YVhTFuyCkU0OvgaL5
FCPrULXbTdsnqjaGvyLJC8peJbogfOp7gTyZdj8H3jrYi+Sg6GIPLyCqW3Jy6Dct
8BNFz1ettnolT/r9qxEvHIdgLf/HBqFBdxm6q6AzSxO6b/+SvT/Ze1OlblJQbDwH
v04fcPGzUTiwP34jVPTdw1YfSFSwUYGbgUiGjrC3NtsAKolZJEZnWd1ZbYDs58Rs
ckIWJvns4Vl8SYqcYL+bgC0UumWOOxPigFnXmpnup7/WxTY0nipSVD7H/EX/dDFN
wuG1wu1wNzVHhJ77AjbrecG4PXZ8ywYLHYdeZ+d3cmNaJeHP+lbHSEJz5T7R+jv9
Y/Q8gOZ+GY3OeaQtbcpbq5UTxg2hn6YdVEaH0oVWL84CB9gTjJUAwEEDHRoapjI3
MbZABVNubZuHysYQ1ut/N6CA5F1r8u6O6UZDSd1GmrIEYulEEq4VpkrR4P9zG2fC
SJBLXLFrUC4/ZGqajruJyHrrcKGJr8HhZdnETk1ltLqSSQLTSoN4DmJZfBUOM3cU
Dw24Pkeo7jpLlkOVi8Ktm4AqROPBa2AEWUIC5ztiowsq8x62ufQlsAyEdb2RX2JY
B0sxRr0zw1MttSJBoh2IEF2HqA5PXTtfAGkZwpv9AnShOUEqYnyH3YM4Lc3X/hmo
8zD24udGYiTlfiXsUDnlws6oD6S+MXw6nS0BcsjKqbChhiFIa1o+uGKOHhnLb7KS
fXH/IeemQCSnuSDwLNHZ9u4fJNL9OTEoAPEeX96kw61d9vzRo1BeB3CjSdxIzfFM
sFQPz4VEj8nNqUJ2qKHfNUcKZkEFPDD8boe0T5GDkl/gfGeJsDiv6V7ST8ojTIrG
R32p1xlJQSy3KTEWAc58yJhMsAnGCFTAWiVSAMntivDPhS5t0qAJbl5gu0OxKrQb
V8f5APIm0x5Hpf1lw/Oi9yVHuMs1yKn5ODZ1nCUmIFuKEbYYBhdDSerUVTb7HZmO
Cc1crUZBslE3jQWxzV0BH/e2RNq/Rm4eCMFolwl5IkxnvbTzng6GcLqZdknAtbwq
zyedDK9UvGReCfwD8UND3isnJMIwLRo2oDv1+hHuksCVh0kG0EwDQTnMrR75KwLW
zYPCBOtCWcDEOhKj4Qmqvm1MMfbQPTwGrFR54efXHNeSVd0FZihrgZlrUKwsDiuW
31wkXTE+gDXa1awQWIkmHIq1sBbDH5lwvA2MXSHpy1c3hBhzoRH2b3JAkM0W+KBP
xJmOKsf0oH/A70lIWrDzLM2trx1+QvgVo466AfBByCToIg9tC+tCsDUbe2koJIQn
McLM/OkB0q78Ufm1DeORownl3QTBo5nqpTz0SWtIQ4VEU5istRA9//lgnOk+1s7R
l+Pz7jdrKs18a5pLkGQmItfzHkd1+qhP/CbNMDkbB3YDdRltLudwKE5ViaDfJY90
syBfuohgQ0WyAD7wR8pN8tHaHEG+acwbUP88a4SVbt4EWz/uozpeO3bsBpOjfAi6
BC/BmNEVxBzJ3JmPtKSSr1DEaaijlnlmjvgAjoJ3y/j2BkLoGE6nGTKr4D36M3RF
akzmmhLaQbB8myiZFOdm9m7NSTLG84aMt+i5d8NuPPOE5790lhuPGFxqqk6dRUHP
VlPnwrH+Bm5qOrHloJXdvCRNyIL3Ud4jTbUnm41Q1F5BgB5NJg2mgRIEWluEciNQ
4lBMTPq1g90MzLxUSTBliKYtMJIenVgqYQNUoAW8HLWDKz++mGe0vE+bmjrDg8nu
dc/wmJkTzUsdcPhg4hFJBPySIizpwZwOOM/72d7TfZRLVhe6qVXSr501JrKC/xfm
jaKtRBv9w3VZ1L+EkQzhK5Dnq3X4CWVU7vYepZRmDvzbnex6pvKnEMi6ytInQg2t
3H8ldFNuL386CsBaMSG9o6G+wZS3NHfTQJzNoWmfU59u/sg4IS4L/KKHE9eYcMHo
d9/R1c+Fuhy4jKYqfkJqHdzT85fyUaVYxFnXut9aWC5S4qeFvOyhi8EJiEN3JxFF
HwoP+NlfXnJZUNnWu0iVkqLNOB42BzQSJauv8Szr90WLl36oEeg9szbrC/LBd5lf
x1xweXkKavPWnLBlbVt1aDwzgMXaxSsvlv6072uaIsDPXfB5QTDDdsxs6wPegqSh
tlTD+GUuoM7LU6GS1yI2qzGHflFNVDSlcCl0B6Aw/LJ0hWW79NfcU6WpV7ZuguiS
rg7fK66vUUsi2ntrO5vdhzbNd+09WBq8cosef/P3JzV5nU1oq6LRgfdwcb8vHMQ8
bCFqaXMHmG+LSxxGP3SbhHUjfLAsosFBQL5uCUA7mrjHvUJXcT0uPN9Dibl2BMIH
ZaeZDF/hAXM2Y/8d3lS7H33U7IU6wasb5xIPL7cKsa57PrQ3OxEswubPDxgLhrVI
B5I7CYCanv/jGNz4rzL1UbqOi0tWf9bTW4d3sNU6tnAOpyrHKo2prJTBQEQ98W3B
SrUjLkGYoYcL0makXPE/9Ok2YnEH2o54QtQVhbkOVXNN7XaHdMpaqcfORZ03hb3d
FEHKU3DBwx0XcWDI8VyT8abo7Qfysiv3he+BweOXPuiyhWKPeyqEqGwptYSofU2g
V/LPq++LUMmoEjcWtgvM5MoDWEP6CcH9dsbbPKV1RWHU95xZJPsFzjV/vIAU2Z+A
JdSdHW3MVFehGfdKufpWkeKicUD4hby1R9p0D1fCMW3PIn4xnhskytOypk0/VzYx
yXA01tnqjgsINdP09AOLjwKt+ZQrsEkSi+gokheSO4ztUfPpbH/ILnF8MSB4Bp3v
CC02GC9Nadyx210baEhFullxgocusVuXjWNKh3ajyz8VozwS6XqD7OreIsYPSQ+G
kWKXqoUe47Zt1BdGhBAK0R4w3uxySUgyMFjrZdqoItrUs5uiAwE+6J2y5IcPB5u4
TKYs9bButUJng7IHi4UAeU8KzJOK3cwLao+Qkk6AbLObWrsaPlwQPODHx7VOTmab
Age2gJZA5KRxrEj4q8RZZEAMOMGL5OBucMi+dI/Cs+1P1J4bS0Hdjlzb2uU1UoNn
HQrNkyFMzVS//aJRB9Wdk3Fm6hAE62a1xirFxfMBbYoTlIOpsfs3KP2E62sz1bNP
4bT/YtN7YThJWVwpeXlxe7oUWBOUoQrQPIsIyyq98EiXiY0V3ZvfnqoUEn5cNTNp
2q4EDsmWtk4BF4S3J3KOZe7F2KkOOvn+UJllMKRLCWX2nWm2Wkc/UGaXQH7Vbisp
2ASgPgnGvGFr2TRT8yoS1ZogorX2cVkk30P4ZPsb7has6G+yfGN3wXesecAKQvSt
nwDIznJW8KCTnRvkJPHRMnCRwegu/0a0dcCg92fyeNjCgfC/oFA5PAaBRXc+np/7
YCv6LDe/fSzgqjZyTwD0Vs3b0H2Xb5Al33r0xHHn8xLoSsqmHN+abf1ZgNruSFtn
vRSz6fQ68i7VqKnmyX1gXbv63VTgD3VkBh+1ki11fBhMJ2Sxt1EbrcjwyeShX013
q3EoCSFXA78A/f5lCBG6GJ5sRQJqyfS7U9BV3sELyayqWsx+Mhlufuq32JYkjaFS
YdICYIbzQSQR3yMBaIy/siQGC06TR6nFfbiJf99tv93NdQZDb20/ITwZPpRy38bi
+b6a9ytfIaQ7FtDA1boL/IXBHv6xJERsT6pRyfyl8FKijz9zviK5ThoRiN5uIRip
BjbMCUofKUJ95UI977TjRKA/faxgk/S5RSJ4HNH9450/FAC/g0qC6WWtKSb8J1Jp
ecdbieztydRPKpfwfpEBF+X4BQ36DZN0A4sPwutYaVF+IR1BlkZwgwZetOiBc6pT
SEGkjJC7udv8OY/akZmFDd4LYX/6FtmDkgDV+7xuYEioVtkarLF1sH1f+1EMZHlp
Grq51i3fMsHmq0UV7iLsThGI6fHjQxAgdhhppx735N045D6sviD4FDqqDO9guqhh
UkA+F1YjD0zIPqJ7Q5tk3C0SfdRNPYqXZlgtv3tjou+VSLkTsP/SC0CVQ67gZro9
q8nB0DIOY9l7v/eFjI5DU+MPRSblbRnUkBE7k+IW57rMtT9pCzlBp3oO0Ex3G6+y
VDT/KtsvJZEtN2P4IfHMj4ENfyzaZWW/0xu1dol7HtwqRNXK2cmIlfLkuQce8l1y
AQyDceuLagLEL1+v/YK5oNgxs6Prwke7Jt6w61Iz2atEkiCKFQZsUOM6Qs6jVWlK
c/6dkfMigu2vexKMfH2ZXmFk4L1jMT3mIRUZDdibt27XtF6JJFpQ1s0uhgF2EiR8
XaOYFIswwW0DW/npeBC3wC1oamoebnz2ZiQ3M4t/sJ+cQvGATKC/ApYI7EznVei0
6cu8rHhSDAS2W7boFkGxYgtQmpU5qA0XEHEsNinw11ARLrUQ9MbbvgjXytZbV6uD
JrK1M0dB9sP5CiwBAsF0sWDaH6n+6Vf6PWamJyKLjZc2qAjzK5OdHNCX+b09Jd+q
LWXsva+w/BmmCy2RBYzGHrgyjnDha5AD+zcKOWxp8xlg8FLZzFVQvPOPblOxLECI
IcmRBlYC2C5v8QrI0e3hfjNewvMD6B/Zs6tZpukpaFCxv5o9Rr1meIad5IQwi6jv
nDYItP53ltOt+Ilx13+rl2suH8jYmF6Mkg5lysJ7v073OAtWdS4h9E61+yumbDUX
vFRclsFCYTe0OE4b/KZGddGZqm857/zjYV8nP1+3wGSn98t/3yziyP27pzll8TDE
texnJERqmeT1na3JKHrL4xLV1RXQ9SQnoXRr85AWKXhlaKZWIBF+WAoGuotlfKHy
6jJqhRpW53F34YNNiwVPSKOEnFqau7FLLMezw/zu25596umLTXmPuht5YcdqnXZh
SN5BlCKHTNccNS5nmiJvWmDLuQQojzVH+WESVJ+uC+mtjOsgAlOpy43mDMTjPGFb
rhZzpqHxmXoYI5EO06FVeDeUeDd0Vz0xBYusEECFYaWUOGEL2aFKfmDn5suTfDR6
IPh3S6PpkWd1GwuweFdWiWo+FSAGHaLMzdFpuIwpTsjVnT18nnRxd8OixwH0td5C
1yN2Rx3taGBZ7kbtNi2OQZifIMSOC5XYWykijBPdFETc4CNr7X+Ov/qaQdf5wl/p
3Fcpd4C5sAGKsa/2W+BR+F41A1YKQe87tlEmlvuiU6uD6eVcyGAmnRw8PwmkeZ3N
Mgcqc0nMmu1c0J0wni4BkgruD5aIwdC/Rz/X2qapotKb+gukBezsiecI6pwaUXlS
dvgGCjaH5mMXdLEj3oCxkxHDFjc2yAsayIB6ITpRZrOvSiXktnyJqCM8ovqkBqD/
8qJyFHuV6DRtbC40YuF2mPtxMTaa9h7EuFbc6+bvtopxK2gCp9nJyABlRFnMxayU
H8rNJXbsGWTRhBtN5DILtxdpJmR1DoL6kCsqAmGlWo/3V6k2GRUlM+mFGJJ5WZc+
Uo1OuRCH5GZkI879hjlu6b/p6We25vLmIm3ijVl0nDsrr0BVHsNaw6cP7uNrhzxX
ku6vL5Qj55g2DqBYs9dWQfrRczwJIfQqut27+bCRVIAB0Pv9dwxd6BayAfE0l/y/
6UQaNw/yBfYRpVTp/8HQVw4bS4KVCJt5hgKgACAYzNRCq0GUPCZVxCh8qIh2X4vg
kzmNhPD9dY/y9nkMjH/irYXxujMD7jxndhLIFyk3qHdK8wfvqlpz4tUuekfddZVS
2Kf2gTp/Nxu/Ccexw92D4FykD117GQoty4rBuW/DDSDplfFOrswl4NLbvEmXlqqJ
vh8ajz24OXIyk3S0vj3C+39GMAPCa0mMOy2iYheNx5YhEWEjXpsux0yBnTSaW28l
shXZwawwsKqFfjVkS7rLQQN6o77SqQzzADHgf127EX8Oz1k0+8HrglanDZODeqaA
Zd/M17vPQLfPN5WScNOw8O8STTRuXPEYn1u65Th1wqSZBleN6hNruuKrknXDnzhc
rMo43k1nV5duu3c3oJVouzsJJ9Jj/DwHAllraRms5RkRhvn7baoXiWKJmwID6tdw
zoFgXeJqaToAxTb6bD5ANnr/78HW1YfUNbQ35e2lMaQF0TphREys5/jTpnYSyeUA
U/ZfGta+z4BqCqn9JE9p+IBxdUOOipb7CZGfp3wZhOgswdb1I2G2TYWwgbqlgtvR
SQNh0JRiBttah+4MwPaKbZU9Fys9bqPDTviFNu9+uohAXKjDYpsPxlb7xG+OwQqv
a5TjAfO7MRN7vkFA6eCMjTXyy3GJmRcYllsST6FqXSSCx1lI4m1G379tO9ZQM32h
5ZJWRDnUlEWCLIg4cgSMOGc8yvFe5YakEhFUKlLbb1vxAxXi9IYcw8tCY+pFIpQg
vO3dp0JS+FNVBNk4E2/xVnypPtE/bwZ/DGzPE2s+gwD32fjaUJIKe152tXIlBJfq
1HRg2uT3nyjqGps4S/JHd32noC/XLrtAk0c2/DX4FWSUFDik6LdSDK+wDMST0sAK
vJSFTpRdwTVYlS8MiPvtXcwCo6YguE4JTfhJVNZIbyxHrCmvrh9Gzy4GM//w1AAu
sHJIgr85iObI4pAs/YLuaDE7wXpzACSuqZ6mJuQd+MgewDfNBLeO7WxoTQ18NEgZ
9SqoKRZcYzyCeZctxd09+vsOMLlGwil3W34hGIMbFIDE87AAm9+N7pu5wRJkxyNu
w+SUizy3uXvy30JCQ5Yb7W0GokBVQQi+t054MVKeLmjOV02jX0p8AL7mHJ6NTVnV
61B3Voc7Jr2jSK8xyli/tv5Xyf1Bnac+VM9YWdBGJR1RPXJzys7JSMmhGrwZWtXZ
+Mm6EXGinA6tw2iduv44qk033Xp7vWRzWgYwcQuZ45lFWkAMFdUMMWiBpn7FXsVg
XXY//R1R3aL2A/WXVbmbK5GTBWz3vXtuNHOIoi82PR4Cjj7jeP/3YgBC9s9dUNde
t1PFmdkFc1YHks9hwkZtG/oR6eS7G7Os1EbNoqZ7Mj5Riv77yLd+uQepuyq0snXM
gTnzDrmcZtVh9UoYmbFscXNUmCRMIAyAefZvJS+Wc5NEsHZyNA+Oh38aX+SCih6v
n50+Z1RrCUT8P9//h1ZiDvZ39MtSubmdyc5lsXXYmh/dCksRqePKuByckxHIvKMz
xCz4q9S2s8vm+0T+Ib0I1kCxMOoXxdJOnKgtS0+zrZBLwKWWZhgSRIRVWUM/PMY7
Y1jj9LTqX1h4YDH+BgoFFphyiUwtbfafg0QUJPRN96DTMfRdktEnKJIDMpwa7neF
Cun/T3tClp8Pef5ZHDMCwmEAsafRTQ0SZLqlO0+CIuB/OdYoyRJKI10MB2q8sSnn
Eii+hQDHFrFDY7l30+9/v2WQUrtr/t4dGdXstxNMGEDBf3Aur7sG9UuivxWXDR9R
uyOKRfrIsHNtGZ8ScRN37e23hMfodCka0P4IXannyB6JJs8nG77xO+ktYZLnhhOU
cm+lIScIciB5mAOL7RqzjyteSwYcqR3QIS6CSmUElNjaarF5Ifmz0uwL94cZwqJO
9onYDe9/84rRey0c6gn8ArDBuemKPeFeWnf4Wdv2FgDM61wD8ZgGiriXXFjV8fnS
0pY2nUMTx6g+0AAtmAqLonZLBWl61win8QeoFlgxXEIVkiCgVlhpnX7WWYEmuIpa
DzWuc/kZvbeF8TPH/xC/CZKIiPZnRQGdjN+DD2lHLBaE2fY0XdkcJH6eHuXcpYyI
laI3nH1RFz+QtyM7P8YC+S/FECaUOnfum08AaII/l7I5BQU+JDrBYt5ofpnAtepb
njVLEmOuyj2TY3cSnFd1ZWMTu9GoFS7GCK88amenGUyzwrOXQd5VoR/nlhFuPIqR
NB5KGYSA4Bj+mMCnbsACtrWAEHplSaspF2sQRneSffM5giA9rF68+XokemiyKp5B
wSeJ722ZgnBaxA21Qgiq/mzH2gRYB/FZpsk2IJ/jbW3utehPXnzO9LSZwdyAe8bc
ty6GCY4lnmnmOTOU7mwLPaIhHbJnlBwz8cayvk2SW3jsVr0Pj4xc+Bk2jZgy5QQk
1IOacKXuCJ600t55XPuOpOCIsx9iWNowMVU4i1Jr36BQpzDUqTDHY3BPVnGX0dy4
kjNY46e7Pw/HEPm9uAWZ7QuISUe83f+w73a5/xhYk/I6z0IiFWriShPjorsjT6Zc
M28wJs4RVjBuSVA1ASqGsKpJfZY+/wWVYCBU6qXtqoH5YkKieUbQ9UUrcIxH/DiQ
VOAGSid41fr4/n0gPImnSnbDhUp17qD8DN6feF91GuY1SDQZWhFSvKJwnPLixs94
gwzvvBMaI+6EhrbS7o21Np8W9EAjpvE2VhPln+0qUQnnJAQ9PnlR/DgiITMHV7s8
45E16rISF6KgVomcR+Bibl4AtZxsDfHeehTW3/B/PGBtbo5cQmAYZ4wy8UMtOeb2
AhUC5AudPqC8PTwhGFrp6Xl0SBgkD9OFBWbWT0wmFWGprIoubx9BXzoNmZ59/Q2T
iiWjWT1fgWjYbcd8QPE1pvqgCHgT2B+yZgytE3uNbpQ5S6tQOP5kYUZHQl69CP4r
+OcWdXQhrap3ggBGsANyq2WLK9x55xetF/CXj9H2VatRKtW/Q6kYLJRyqqaLVX2r
VxS83jwE2wTn3pTfpsQPq+eCd8Zmk9Owv9kOYRy8ihsASfQNbQB0csVlgRVpaM4Q
7oA/uPuYkvw2k46Kv6s99EKMf7hXUSO8PCakYT9q6qOSN1U88lA7chypfAP0l52I
IsK/J2kJC7RADybumYKZcGco4IPvEKDE4g2g+eeqvIEhJ2lf5TUZEZ3guUa2DdlH
aZfFmV6u9XhvQGkynWjDXyCZhU9qJ6FvCBHUH7qEGLHq/glPWCdjC9rTkVyR9TxA
e3YbO2XpuDyMFq14wauosiG4vP2Fg7YtWORg/vyVpp87xwPsfRbWAMCtoJiaDxvw
Ha9Gqhw7THA0nI/122WIcP6RGCF/hsSQVDgOVpd9Ke13dNb5a9lBgtKR3QeOaAkA
+dfzViS0O/o/cavxYO186saU7dMHC3vGsA7sN0pvPJS1Qcekot/w0rEBh3cBSArl
70Fq0jWqhT4os1XqhYkYZqiPn+gmedET/x/HncNti2267DsyuHVAHbBZ5Q6hXv7V
NRd2VwqSPu5YmKR1H7z4xDnvfMxkjd4BXMP0/YcRWDj+RP3YsD00Tj4Vtm6E8T2+
kgW2xsK1CphRuOakgITcoN6ZdDEl5iCY7oYVYbPWC37od4b8VTDT21pQRKoclj98
aEnsQJbFRxWlmgCRKVpojyHKFuBqs+qTlBk2EtnY550Imrsubq8gZTb+QeOCwHq+
loPPh3/bBv558yxgYw85Pcfc3lPQ38z9XaHsVy3mFoLrJ5rxuqKYTmZU1q7+tmiO
XCbdgipWkoIgiBfR3NaW6LQj3+0poNkStPkvs8G+rgZunhWYLpmUoU5tnJg4Fhmo
yLnA05ytVcL12HnHnQnkLhhRKlUDXsixnN10z/ZSlEkkl48VDf+xx7D4K5fBl4jl
dRwwfPtJAf3A7r2EdnwyLJ3Y9lwyJfSs4JIPcmke6Jct9UslrnOfqUHRNIkEDcpd
x4bVQXiWbJnf8g1pF6txnPvpicHnv9po1VwgVUlfvnpB2Y6N+kFrPdAxD9ciDG5G
LRT+AxliV1nCnyGT7SICCP3EKV/9NPjPopc+acSjCS7lpfBzayYE1WbR3fXKhYXp
Qny9COMzseSN4Ql5vinzuL/cNSamqrBjsV5Ki14GCBaH1bSZX7OWuuNBRNsojiAY
K9upc3ijl1Cwh7m4v/kEh7V2VqOCv9VbzMc4wIcFFP9JWh2YIITjy4thi2P6dpx8
ALyP5/Tl+cjKaaCa9g6xmiKSaILxbvq2s8lyKBgb2j844b0UaJEWCVQbm3GElVh0
NkKMLRL2SN0ealZ3ITLhNjUhR+00dLBjEL76qIClj417z0vTLR+61Uh4GWnquZox
bBtoZNRHH0IQmbjdBkRAMWnxor8QZCPf7jByOtGnWIzPX7TdZe9i2zMPjNsR9DZz
9ITPyWHu3mEYOLCgTUB/+KBudWI4XkkVEo44EJoqjoF/Vi7lmkiTH5Jnfh8U6WCL
tHQ2OprlZ5WFRn+H+/o5TlCpb78qMsEFWmYt4e9NAh7KDosA6c5aO5C4jFdg+qNn
J1J7yLTN0sg7dryqazfOs5LVjqkUhG8Sd36u2eRe4/8j/KEnYluHE94ntJnUi0U5
iWSvL9XqtyRxLL+p++sz8v8HjbV7D0tZl4t65ifERDtCLEOkYwcf2iFL0f1/hjqg
jNPvdgAvlkTTWMR4+3RhI07yQspU9gzEZ2NcJM2R989lWLWG0NP83QZ8iYx71itJ
mGjrHYn3UZX/3A4LP4fulc4/6xARxLLKn1a0H75fNq2AhGSbI2AeerJ8ucHAYDPH
Lz7F4GVt5ae0KNpmk+rVS5PlCxnPdYfnT6TOuYnpGBbABUnEI7GjpW5NzrlekOab
xFAuaI6Vt+o/viax8Lj0qvqdJk1GUAPyFrN6Iu1N1hXpToTWnU+H9982OTCDwzZS
uJGJRShegAZlv9/715GFiOZPBzASAquf5Fav3knLTN7nVtg6HEtkbtst3r/lLsUT
k3Y2eOm1i8GLTTK5564dA7AG+DEsDzfZSJnyZmNmPG5ggNXpeJLMWHpmoTDqJ+wZ
LOoUVffF75JeP6/y2QmbPL+KTGo4BpDJSQ7W1C6oYZ3j7X/viQ5eqz9ps0HDOHKx
ruI3e3u8cSQpyx4i6gqOVvMbAV1H+7rfROQxA3WBQztBNqUFuHcRiIuvO/4C/ZCe
SJ+k0n98TYt3H/MeNf3AhV8ViZC+T3O+lyDW9x4QAWB+O8cKUPiAB8RNF1Pgp9NL
h1/SUcbR49BIVx/KabflfxQKoO+5kAoEfblrxlIeFGPXX79d5ke21sIhM2oaXDpw
34xcJQRGiRd2IAoA2fFizTEG5dirvwLkYBG2E9tcDFh8uBN+tgqx8164aeJjpS5Q
R2TVJH++DJCfaIIG0Gz9/s8kBL2WW6Sb32NM3aGy25XCsMRKAVRbucdTulPdCa8e
mfdgxXnIRdch0Tbclv/qyKyFTh3TVuDz/QfsHiU0uD+y0ZDjmine1ZTXzx85DDyv
4jhtBit0VmBO13o8ZPYapX0DrtvqZpsADfCMzRn/kDr85VzDWIHaqd9wBZxjZ955
rCjZse87NJ0RoYQiZxG8RrDwIhGFRVihV6UySa6+gstoiXWptT2QD87WASnDEMQG
EOFCWTOQtm2xiju1YAjjsF0Dsu39VwXujwMX7VFvLpuC6ZY3FGiBGO7k/6Q/HDmM
tJxxW0xF8vLPFlJSUPbgaagSqVA+YIjsCa6tbJ1HJ9ekFrGVuPFvCs2MoKmd5+Vx
ilhsosVcQNFj2mEzBqKcH/qjEKJAOmeSImwPGxmcL/KyOg1m6YVZnifyzZc4D/3t
SiDcGi+BBweSBh5oP010EJdrToLbKNdtcg/m5ekoeSbzJ5rbYGzMo19xYcyF9jfO
TpakIruQ4LsC948zDdhLXP7fp6WaS7KbkYfGYoN64VzIO6Cal9u4weXxXViY/rpk
e4WYVuzM/z5PKshLdCTJAXlwEWnQIBnnx7pKhQV30idXcwodW1UuicmGdN/u0/RC
uXW+iNu+YMf+buBNyzVbTO+mvVJOC3oI+VYyrryifZEM3oCY8QNN0mZURVpRZi9v
huESw8l2gvcANMZ78CxKUjcu2FQD4CDbYTc+YNzDJ8vny4KaK4aUGbG+zkSy0xe9
vPyTxkN9A/zt6MmE928r2/jGB3nGx5RBjh4GWItrznuDnCtbdiohwN/3BQeGlWBt
y5jmi2+L3ge9elwRsfYKDzT9MsqgVfvnmFyQqr+yuGSUqUjco9W+SsFzPK8aTjU0
cWOg/YCxl1S4JkJaNJY/CoqWTHd51nlf60VLhNel3YRqBCfO+22HMrenQQS/P8R6
rUnnyGfZIZJt2EavUWE6QpbyLVYNV6YXY8PhJJu/yN/wDcC6GcBc3d5VBcTOT+5E
Z6uekZhb2QFLEgg1a0dTpGqE3ewU2huqoWEnRZpvZDf3R27QPlNll4N+V/3Tl53b
mEG04IGBH7dEy/ZbTxx1VPA8W9agN87hk2QGi/lzc0rIrw8xl2c+FbMouGf59/Pj
/0TsJpByunuOuaO5UIDdXu19+A+m6yt2LBV8Nocki+dAelPRLPXhkJ4K0vXATyAf
3RboR0hW/aS1ESdaPtcfieJ6ngz9mUHySBC2Ulcx5P2vDD7GproQ/LFEiVJZ0xzb
qMLhVX0N7HiH8ALHEh1bEfCK9pjy8+K05ilWr3b2FxDXJkn4SF5/Daho4FdB9Mar
HLumk/z6uHeG5g8Swd623G9/NV1Y/Qrpbr3uhYkdkx9L6GRzEUkRoNOxmgHnjQP/
Kgw6ucjZYjeAapppe+n/F0aR+y+QjbvfbKRCh7IUxp5Aktjg/vAU7G8eW0pkRjkC
G//Qf00JZkxefAtJwEXkp7foFH3mtR+tL/5kmfNJlPFupwD8UzbJE5FrxZZVgu58
c6Bo5HnJywTv6RSm9OTjNb3q785DtfRLdH00+HPUSjmZNznEcZWo6KSJLNp6z0dQ
I4X7Ws54U0v6nT7TcKsmRsKsH8j9Pm569d3ae4hcsOqAYsJbJF+4EaDNCdaea/++
qy8uJFD+b+QXer4Mc4artZ3sZTjJIjURZmLWAo3buJtnsm0XXgQvBV8gh0+qlNAO
bhBqSrKYjeYesFAmx/b4Xesmk8+LPOjE04im59gJ8wBOLldfI8vQm9YaEwIiEdni
dtGfzmajGzEeri1xqlXR6E6XbfqkVIbmg5oF8ibe+WOaiXpurGYKknSEbF3P+Hd/
Gdp/YXwJa0JwP78LHg4ih0ILYvEV5H3jZTEDupVa1cOkdIbc+I/ErYgZmcV9ejPP
ha99fNOTulz0Wu/FLCeD71LLQ3TwkzIreWkhiVv5o7HrmrrXji7o6NeVdSJz/VhC
4chXFkY5zU5fUMDycCzVwL/1Nr/bz3nE2CGWOwwAkkDuq70tyv3PiQt5qQV72BXz
YjmwYrpFiRSGyC0iW/XXEqn5CJJIHanL2lxu9/Rb8f3+LApBjlYw4l5ob+IuWnG7
wrmu1jkPT/CXKTzwMQZh1bPhSWYUKn6bnuN7py1Fo2GxCoQK4IxnVJywvlQD6dNe
ppSHganfKyI3mdG91h1XUq/AqS48hqJcH2nXCtRQjZKopGKHi8IpYM3d7xVxidDP
ffD+udSayGneDOQLHj/OhOpDFohSYfVJ+vVLR4IPJI44HdBlRcix6okLjhELDfMJ
YtaPAEyQTGS90GQt9fQ8lXWloIUGV0j0fZoxxKeqb9tFNCyBwvBkRJHK7NaQmSnj
3oEr5trA2fmI5U2LYvhwt8g97HRcG4wuewX7+Czv/99jS/qcaQH9QwvYtZ6SI/5d
vNTwfPdpQv7bOYoSblZnPX2d/MIgDMgfc8cj9e23kNZKXnAsHn5tvNoLLMa3RzKS
ApwoyeMqsDcg/R7LdRMWK9pnexsW2dzvJUJf4w3etvYn5WAPwguzZRHr8s0wcIJ9
Y0LHSowvwVyE8NVucjq1v2P/lLFUK4DxxLMSbnj2mDKUUpkiAMQ0+jFE70jxF9iF
Vj2fTlpk2GcoXQXwe2/awEsPD1xeUINb67pcNpUhwfgkwaWh/1WDzMvB88BLY+SL
t41F+LJK19TbIJ9LGNYtHC5NZEsX/6wCcteOzuQWlhywOpbOota4jfC2oji/arr1
hhHwNAlDP7LM41wKOFJ4pAoFHxn7QcxBOQpqHvnIRqUNtKYUApU88hdj9jfW1KM3
g/5SEco8Iyf0JLoT+VfL2ymHQ2gd7hIo+Dy6i0XL9nR0lMdH40Sn8w+D0/9L8xM3
1GHOmL/2gU7qsbZ1+oc0J76ilGxhI3QIpmUhQcSeznDbixjH92whsdR7n+2iIdBf
ssKeqb/vs65qd40UpgjWtsYjXV4uVs6c772filYJwHw56YI/3EyBa4vYrs+b6diy
6DZcVMox2qOuXpWoUqAhPY7j9+Dxh7beI8B/aqePWVRLH3Kx6Kxi7MyoUQagCv/U
EawzphiUMqoGQ9H4AC/92AMoEJkgzpBW1koYpmopB58zUYKGT+rtQth0Dx9ts2Sm
tJCp3QQ/kQ3xskojf7qJ+KJ6AXd8UidNrGeMXZ+RRXigEcRV1NSsFHE3WXfgGQwe
MWEU3nnHcUWd1ddrWuPldefREOPSOg9SwiPdlZdI7MGDf0p5h5FmL4nZhhkrOApM
AZjZ8BtjgTe+7ecU5wd3z1cGwgGsX4ZX4Vkm109rQHp7T+rVxGA/N+k50eL62ag4
NxoOeIzblCDMU0y0lFIMZQi4mR02iE1wcLQUBrL2X1lbH9moPKSgae3kQUe+rhEw
OEV9bBJSBdDk6KISxDAB26hmh+pl484oqe1CAoFC+UXeI5wh6qgaTxcITR6H6Zp5
52+edu0qGU4lkb0Nd7wMqqHaZ9KXse1zalqoVQ9KgwMxc20y9zjW7+qzL3xHh7KD
ZbCJDyk1wgZBRb/yKNINJacGP052fEZGjJfs9V5h8QjUovzLEf10OElDJnOzHNQE
i7f9M9zYvGEHxSyUvsRg94Yq8ktguNjEAiUzQeEg6fYgCQpuFyI/FvPkaYOqQyMx
ZNBULiBlPVip3LgnR47dh0cFNmyJfNL5+RPttAdJ5X3Sy5GPizkBbtRtdKCUYCkl
vdhp9wKn0LJGZXEV9RVknd9HNZjdvzdddCD4QzBuvza+MmvSaxLCj3VIJjok+kvI
YJ0KvF3fOcECjlx616ZKL7GYmXNAPNDq7AhvyfZbciG7hnYsFIqLY+ZWSWXZkHBq
KWssskktZe9XUhqhqIUZtclSEI863XcJVj6gddiwxbAFr3Ed9IWBgO627g6JgKv0
tlwq6eZmOnI5yFyff0etlSTJepg5zGmmaAuRqKKKlDFvsSFr/s0QZYG76d2hSXmi
bCbMsNFC7RMHJ+iLiarQin1vILVJnj6+4cMmcbAfmnTWanga+zWxjWU+Xt2ZXQHv
qGmp9nSh2YgpZbUIBim7h+rNSql80Ks3IYje2ZNSR5hoBtd9lgxO3ApEeYkL9V5W
ZYevH4B4KDIIEf6iAVYmDZC6L6IS05FHxrr+yl+Mp5NEs7MziYzJzoGjga3LkCbA
RwIkY1wva6BVHE08N2tAl4tX+90g1bVc+JxWE5dpvTcx9GQu45lqy3buZKkGlZAT
+KbHDDbAQ9Tth3Ke6JyVb7ujba7lwMxMvSI45z+Bfqw4knD9Bfo168+5MaXcXHR0
bfM6BFePKKNRA6zwL5mqdun/CyPQGTASeocGdzQn1iXt32IHbH+6G807Pcl8Dd1p
bS83IjBOu6ShBpK0Ivn2pspC1lxYtCpUmdkQBHlP2fQqJSiAa85HbZGIIZ63et7C
WwRIVrOf1Eeihn5yguReLX5OpOjB1Vun38dinRpCtTpoza5m4TIN+DVnzgV7lajh
R5aiv38osL4BMNnD/ZthsA4zIZua/ZP5iZCqE158AksJdhqpSfA7xm56GVyIAAHh
L4yEihtOmFf7HoYE0YU4UR1fJVYzFbEE6NUQ+jGCaAf6oP6eimWwg5EpwdA5tmvB
uziuSeQ3ksQ6ALtDpo50yJMQn6vWNpm5fQ+DSd+Urusi6ewDJLFIWaxzJlRK2oib
MsM8OZzNMMv6MeIK2/9RoIQm4onMtdas8TnDhECl0YxmzdJhtbItjhp8CRrDIjBm
fg7mvecZMbCw35WvILwdx9OPa9VucQgQcRSph6TXPxicYVvfGQLUMS+RSd92skc7
DPsgoGwb6Akq2e46lnyOYfdX7eVngsNq87Nui1ICDGJAXaCZSdgR/+9dgbGSUn/8
pOuKhld4NzzKZ4yhYCbME/NAQOZefUqjDDdh9dsLuRV5kAGDJgvJZKxWoRrpe8/V
GG5qPmWLbiDA7JpfriNJdyxIKCgfx+N70uo57pVgrApbQa6wn2jgPpggbUxCubhU
FCU9+yJLM1aOnpYFxxHFDP6E0GcRAhmrCH+6uvHWZXmc4L87s2tSpQRHrzP0cWN2
j0COK6IUI1fsS1E0hwDGcLzgF/mbAbOrJTL/SfPpVyL5O2T3AfFoKdlNAiWBGoAz
MfyaGxQljThZtwh5S2vXe9itUtNSVPCHCz1ckD2k07QZsf8huVvXyBQdjR1b+CAA
p0paktmFn6AUorEXqaG61qVQHR8e/MsEtp+nky6Y9oRPR8NcF879IjKSJbrFcDVK
ZJnsmOUHWPw4bhcnLkkPT+8spY+n/Tp/RzdbBLLuWNAu46ZEvlUcfBIJ9TYnqAU0
nru1u85yp2TgT3SvOuqaH/2PbK4cWlmXiTwkbBVzmqhcPvnZWURaqQ48/gfWJkVb
i8TiBKlcm/b2BASQeWQROYdgrjbCufwrkaPunQFFLrRHCdCFFKK5g0AOtl5kiQ2u
AtkfiTjCdYSotMYQ82jRxhEAg5N2JubTTG1PKNmdiIrh0+NhwOb43wUJuZ1ZuGVN
wWDHdlmeDYINYDUa+PUIHG6rV4sllHuJlJtLYnPuPRh1dkZJO2NsKGt8JI3135oo
NEF96+EUUP2fMLCn3lTHhoYScPWD28OoSJc3JUd5UVo5m6BvekvTtLjXZ3tHpmaV
0GrrknMkcdNk97EPlqwLl/ub4I59tvp5hftNpfoB2EUVcjb1CJMznEi5DG+KO4uB
vFlT5OXI+lxLaX2KtANdoScrcgjWWBFAMUmrtVi1IQUww8soEVk29WAykTIj/ttg
iW7P36l07ci7ibSelNzlqdbs2L2PJwtbVoQgX4UiQrkC8Id/GrBYSpqwLS5K+qvB
hd2Qxg5h8DZ+9PxtbqY8OrNuPQXn+RvDNIFw3I4KYGwIxdBNGbXY0fqxX0/GXGX0
uKP/9dfdDj0ZWiT/CSuytI3bOnmnKYyQXv4agxI08dJUp9BM5w3EIAyUCIXbnxnx
DNwYi4XvnnphA6WlD99h9Hl2j+RQZem/419WM3kn+ek2bWuPxSfYsCzGRFR+P351
v2u5f9avYywazUgkP6qTEr6WN0N5QgO/lP1B19AB6yIBk2/cG86tC48/sX6Qtf9x
HUr1wuRG/I+EemUygsbxRYeuaAcALkYMZI7r+vTHIYj0aGq8ybOZD2/PEKudzhHI
kyYDP9N2g6Ghof22ktTM97s1VBK9xxthjSX4u+M9CFCRo0MbVZ3p3ETnAc+mIgF2
v6bfpbYXwxCef/GvBXftPZ5acnIssgZu+DKP11uZFLSifZA4d6EzJ7LVklujIafI
bL1TTD1b/h47f2zh/ryP3jdwAycIK03F+I7YVjC4e5B9ILcayp7NNXztI449inYI
Sa+5ORYYFkL6/0ZOLLfncQYti7MvYlqZwdl8zWfinfBGySNIatbvwZB276yIn1lE
XFRmwHsdF8ouZkkxQvDMbUizZS4s53oa++V+CunjiIKvUY2v/YZRVSk678U8X5mJ
BRsM8XN2l0m5Z3B0kgA97AaV0KRYTUGs3+3s+f2Zchpi3Aym+VDBK63zAFzJn06Y
onfTan9Xsdn1MkHZN426aVFAkrOS+NMkJV8QLj3ZasRH07mjKwGq7PyKN43s+vLZ
CUtmLub8LHVlMOh7sIXbVRLtJTGiiirBsJiXBn/l12hhUynlAvcBUwiVYSFYPQYg
ILBKq1GWznl/xVlURaE8uKm5J1SGyruaOZ8zXuRjN5Nl65I8aSgEuu5UrkveWNER
c1USJluzgnOvafflIdYb0/YbDFe9YtqkpAykXY2qp85z+4D1Xkb5jFY3mS05bXTU
F7yGTB/9iF8wqE4b4edaTfdFyq3FWJ3Eh4GZtrhgVd4+E82D1KWZmxXpZVirT1RY
Wqk2KxV7VhETU6LKeTiKGmjnRZCwona+lyUnWx4T7L689iuFcdC3SIDVIGlUAFxQ
DposgbmIWzD48FBCnAuNeuHSqcJJz0ROsqmmuR9d9YzuPZjLLLZRxhLZ9z8q9im7
gJLdcBsZxqwfjppwB2aKQZGkiTNE2WUGEE0ojA/PshHTfjw5joTbkFlhyr7KmnkD
Sj4TbmVdnLz2xiEB82cwIEZzpYSjrk1Kqj9yC9WvtJWg7itdwCw6RHfXu4DGQ9OX
r4mnsX9Uqo8gjwv41wwTKibCBAXcaYRgftSyarKC5ehw0knuwya+y0GMgD0SQf4B
UY3vqXHHNz0qLMCIrS9qrPC79jOUxYgUJ35oZ/QOYPhoc6nIcFN3ExRhGyDN1J76
ZjULjjeKFCHkpJCjUVzchg1C24i7QITwPUoz+sxWB5JLGEFvSQtreyE3zEamqzDK
QSlP0GqmJ04O/WILuguK/HMNYlAgMwYp4jq21NIA5F1nJrk2s6GrNO+NnZt9MR0m
D7tzWtuzgCXRAgFJHi//kqKW4XKqc7wKF2qe6UUKFCNSgPXwHg4LqYfGySRCZw4G
qvvlYk7itpaQsXAAxlVvgdowZ8qHiwNXzF7W21hZEg/XVv0WQTB+ttqvHzDogEgq
aUxE+kxkXfJnPjWgeYfDvRCzL34cIZ2BVijIKi3lOnRVproRUJIr90GYEAhoeM3G
YnmTCH3XOeWjzY18Gvk4PdK5HFHQjf4vRFTC+T6zuAGLHCQoEq4tJkUh0vYbD32M
VemSnD8TswaPtIBL+TMtQth5pJTxrDTTJN3xhlbLkgAS7EMCppO+iLxs2Iamcf89
EZMw/7okFMVQrfVr+k4D0EM7jR9m//k34ggzyTVT7wmZnIClbtLzVKV0N2wCKwj8
acwB+D+E4ATxoZLkTSTOc9AXp2/CsP0gR1pasH7EgIe0w3S5X6CAVvLZc3gwYDUz
+X8vsi0DjNu4zYuoR4WtsKildAXYpVTZxZPQeJ8jlgVj4by8LYvVN/EPnS8oI0PJ
el7VP0gQcfOgVVV4w0Bo1jHZeE22FuNVSc6sL/xY6Ak5Pka8YaJXzEHVMr9BPTvO
COaBWVQp5ZRP1Rbt11SPVWRngBcK2qT0EsS7uvg1HVvdRjTaL0R/+wTRCT1KfWeF
pki+4ceQ64MQmZORXH1TMC8XeRnOoIeRBpZwZNI3ocTJEmYqtANPj+j6hJ9sfxp7
qUb/5YtDQTxEytbSDxqn0zPqJufOiEwLd6/PF9VH2Dl1p86zkb/gcHh5nfQ050Sk
bSSBn3pGh8u/Ffd6/2VzydnIEt946hbZh+klsqFMntzxG01Pchat4dtwAsiafRkz
WncAGAWIQ9P1ItmhejhLyIHM0Oc6I7m+xWXGCm39a7IyM49x89C9HB2yA9GbHre/
NUzBNORq073ejLwH7edGQzgMXp0QP6E8k/fu/LWguXYdslWM6mPhLfVTPYk1SnwN
SsY8gExyr39HllrfSehuJFYSQc8wBRHAqIpgWJyyCZem6p58tLjH6d4H4FnilF2X
unSdWMaQzUfLs+NpHzNCXQILfIc0W06pOKKS8Dg670DLApwnHQWAuvMjtr2QtVYO
q+HTCdsl56/fLFCAbhb7v5woeornU6KIBG+pObg/g2EJkpLUZ/8Fv0ioiA2CjN++
KE2x2r6uD0YGG2224r3k0jbbZISSphX8oTLnOlr5ZYNNie2EtlMOSs8SDypdTRo/
Q1er0XQTid3xcvfG2GTDOtwRp7ZjTeK3YVAywtPSrKvrZ1bGGDtKmrLF7/sfjTHi
3ninjeuxs1ls+OAoIpT5VEBfk8jMxU0y4Sgu8uz0BjdSBxKXvkAPwvX0CIEBEJN8
6dEXJ73akYLGxL/OL22hn7gRepKgYM4Q/ueXcRTrFRLcqX5JZWsul+J/R/JjzPpX
MD3YkEelWo6D9djctyS/wYdVmPWOIKpK0oeS/ePmP1Uozljjqn50rhHybi3QCZ3w
/iVAbsS87mHDOt7NkKdc8Jk2p4s+Q4w1DPQ5rxf2DGSUVp171+jyphQGaZAjKJ0N
ppsSJKbN/RTl/h+1zm7bBuN6g8T22FrFYTDXruelSuGXCaLeBzzgIu1VZbOnVsSG
xW+Ix7PKul9iCHmNRh7QCe5dewuS6RF6BAU9VMychcmHE2myUx0UeYbrrr7sz6vr
I7QLdLueXwJDjDhjWbsbsoi9S03XMHzGEckvLKgF66TxpMKWJfRGtT/p4KliV6MW
0wbqWZwMLpjNBtWRPvk8kgR8zofo9xV3MO0Sn6MJ8QLMR+Ush/hbevn34JGuRUsU
4yPnOg4UV/G9A7KheZrCKmjBRHfYHzU3VF7wXKF03hoomnQ2eZtUBh/Y9fY2QOi9
GyP3Oh2ZMtkaIgruio0NdryByq9PY6Idy1rSLJYmsk3y5y2r1cJB9TZiY7OPA16i
FsiCZ+vMILLB9T5ErpJoZireMWw3HwdqNZV7bDYWIPn6vdZCZASh4wursDptktL0
hWcII9RG1kAliyneKTCF3aiawg/+GZp8V2oTPD0ZAbgrE4cqOt8LOrqUxrsTcafr
LtAxdzOyJq/QLp06CgNOkj7+RrryB4EzLu/X1PBm8S33s1W7jE1C5dkLGOmYtDTg
iJa1OANd72CHpdKzu8KZivD4JbT87DVWHSoWu3ACHxW5vZT9BtSHHprZPOwgLzxt
mcdhMEyQZwa2sxT7ZDcFvaWFjShH7BWctR0QqUiaPh3aO1nM1CXigoD8dEdY2EWq
5b+kUd2i8zgKh6QtJ812xXnhYlx536mufsH+kKf+aWDhNSUCPk2QXktjUIeo39I1
cRjcadgFlOy7lw+5MV+yXF5kXrqbLop8nMFejGpA+eH9ZzcmsRJd6BBqQten1Ks1
Ab2EnY76bM2axIb6dzmLCMirz7XaU1ER1LvW6FZwwNIiuphXNFPlEj5cXd7N/D3R
CCf1hDyZn2F8LB2tp3kT8lvCeycB+F+jC640Y+Rmdfel5y8YNIkpgfkqolXcNQL3
3uwVJN5QkCX5QC3gXmeQPlxzg4zZLrSjqL77Z+SqRUsBW2lZN/Hwqqget4m99OXe
bYn5XGu5SQH5iO0ekZDlHhfqTowNwvFtM3VihVYBh2Rsw46/vcc8dM0F+nSHjQ/z
x33E/IPoQMGeTEBmNybg8kyMhWkBXQDri/mtUXzFKJpE/UE6R8zGiyWfFKXTpFxL
fxN0hc2863K5fkew2oE55wc9HastDQSsdiXkxkTXZE+gY7MQAY/NV1O+o8Z6cuvo
Mq0MoB4BZFeuoldVlFkD6GDedwh7IdEapHV3EbxuUjXeUsTxHl2KNX8f1vF6CEwO
wuJ8eyn7R0oebFS0wWCy3sVP3QGyE3u7cZrB66F895f66yO5gJbF32umbzA1iubb
wP0y/03ayPTamL7V8dWc9HNqeJtZtdM/KUSe0U/atjon1uENw8UIaRDFNLb2AYVM
bC0NHdvkOZTiL4IboQ0aUBU1+5P+WZy6h/ut1pELfgIhVOfGHHQL8O2DwTbFfKfJ
9WVeu4/tVElgnL50bjHb1Ik3WELQRnJwCXu/oJJYnPgvh9NpK8bmgXbM9qLh3Ivk
GzwKt96nbUbXRL/Dfd6sRKYoWRPLzjAwuBBLlrpzoxkUDElooHOEhOQ2cFj5LaOz
2gSup0S/5+NpanTimyr+zq1OR4C75wEYb6JDa9UJLIV7Ea5iWRPzKvS0+XTNXXnv
n1rXOIln6nGI2lp4ndrmGAEjEk8y3yo1fFRN8LfQS0wK+FPZRUhbnsffkx/XuooN
YQBZqIPLWGBr2lfXull1PbvF0cMO03f+89ICF2sU9N3g7nR7XPCHuauXIrkNGEJi
OHgtrp5UWd84SJf+qUmXi5NLYWbeuiTq5//ubXM8J+SIcWOUlOA4NWZ21fPTt7YE
otvnCNANAz59ikmcgpe07K+JWuAFLPLt8H4K2oK8hLi7k9PwYc85PVR84AVlX9Ks
Tpd5ILtvGsavM4NYvW/qjwpx5jL2Rj1FeUdqiwzfckXE01D/weVqUf4sRWOYr/Di
p4cGZKbJ39kdFliO6Dgbbi5UmB/5FM6Z6imDrioFWxRYdpLHWgboowlUgUC81bdn
bqYIL2nOEn2uc/UfS02YZb+ssKp2/JDAu18OKQXxwEWGwEj7lB8NKV+Q2xZowKE1
BdHxPE7Jw0I9cdVLQZQGjVwgoIVLSNQqD6Wo7MgMy5NJjRUlq9r7yjnzvBmlqCZZ
vs8otYbd1cv0qMXPlTkNKxpctpM2rMN1D2fpgsG0Icwg5qZdyrMfiyLTC2RCepz5
CvzW/0Xt/XqKqj6GFECZMA6suyfJHAF9KDamWRBdIdFlqw2ZMc+YCu8g7wtqiphn
3gXF9CNkcoOGxLC5yXUSphjR9Yf7Bs1wF0lJxDEULI8sRINr2iYD84scRZ0pnZfI
SXnIkGxeoEj7F/QiVnywE8XA0iuhJNdqXMTZvTbIDOWwwzNtgehaWYnXdeFiHfwQ
O/G4y5ENZ7Ib380pircIUi+DnCEkPPu/pRT++dPJnyxYJ6FgQLxI38Cuu4rMnA+g
ArqUV3t7rLqTk+4HwyoMHW3iZbkjiiJtMotlFPJzgLDeYlf+jawgqEW8DLNIhJdt
OPb/ao7XxNJBpcya7yKlf8mZkP4cxiVODaMdIrHxjsMRH9g80MxQvi7+c7+h9XjG
xXbd/V7SgVVy8U45H4IjxF7BFq/pfwD0oJoJU4IavjKdHwhYlRaN7bP3LOhoUkl6
38Y9O2hiCOy7kt840EY3nT6dvBzkpDW8wtuP4A7fL54He0523SeEM/CYPDSw9WlI
GNNGPAaY7Gghwy3ZxdUXEmrwWbulpyP7NjhBTXcQPX08yVRMYKAZ0n51No+bkGFk
GUaT9sATGifh5dA/WK2SbT7VyxGs7lj9BxOfQdUsx4whAHrO/Fnj5yoGGOfTus+0
n0MTmycdPSdlDeD8MzhcQLyOZlGPlz+2MdKXtQCXjfeVR5dIU2R6wpVLYXy89kve
1kUT61x45mj+1jXVhqQtsL+aZkKJd1SWfqhW3el5/4diRDYQbGbkpkwAZzn5qCJT
tMBnp2wt+R1j4eOGSkQ+zXQOjMbvA2rqNfgGHM8J9pOoBR5EMRAz8M0W6FvjeObw
CK+ij+W5m+8UYXQ/JRkXL4Y8hCiKqyDrpsbcm64J+ZN4wPlZ5Q9/bN59wq/1mIco
wZfMYsiOHHNjg+UDmsQFkGbLzJZE/rqBdD4jQGJlK4fOadAdZ1r47rd+nEJBxCa/
DHw6bRVrBjZwy5PNJ8/bRniZ8LPq8V0L96jeq+lxtjI4QnyauBbnaM4LDSpRFlJ/
JbcOtX2MCWJMlgc0F03yR1bF30L3MtWOph6HVCwaTny4Vlfl1g4Cbk9gebIr0g52
ZkCLMKiJ4N1P9nVN+Q3kIOdAhFiXddB+RSeFbN2oIzC2Qbo4HkpD2K7+urBIMI+i
w7MitqiNt794fIGCBaTiaJ7nIaSx82i9b6zrnHZflttZkv/DJuLbKKqmSuSiCWB/
7JUQCI8kMwGNXYvsYgfBcUewWgrp6sOU1OQAN7w6/kbr9ZjislIqLA8Wculsa5Jw
iFNxMlb9Q5cuxwU23X6xBk0MRgZ87cj2RE31gPNrCofAsR6y4JKUkWSmA4neM8Fe
xLPR7O2jlxcoaCWrugEQejcwFOX4oXrJoC8S6rjSEtmuTJY39SMVLvaMp2/2RHQo
VJ0o1C250MRTdZHTLN4gLh5z0F9yDwvj0nNyjtE+/I44D6eZ7FUygBT5P3XnaLs5
IIz3TeYWO8yIWMOL/oVqRjzX5AcwiYKLIQowGmUIYsGdpyPY2dKfGEjI2CxYt+gF
IkLAqXE5lsaIKHWqaIhBXMr4zD4fozpndHKmlX1uHo0nIIm8al5yRwzvDg/8IQLH
mFCale1cIrg1YeJ+QB/kzP1YUJsen4uf1d0Ify8lZsY2aLwjyEkSP7wiMB74/jQI
XAr4b1XRkq5g4/NUtVxtdCOzwDX+NeMdL3BYqFyVuJMEWk8VHtncheYNHEZ9aOi5
Q9SrVq+cPOiwgObD6VcsHeYPcrL3aigB+o+mAvgvtH1fBBXinjItP22X5/qenOK3
5idlSoR37WeM5dTXL9WPRdf1NpVH9DQ58t4ebLW5F9wIqImyu2SbpJvQ3otcMBcK
B1MQMqMpkbTie47GAisVnYm2ikplcYmyziyv484eI8w//j8Y8x4ccPaUKp4ptuED
x65Uvj3BoT5pvpxy4wnbFrWgUgt9N5ffbiSAMFC94bb2C82FA8dmcNuua/FhVWqB
hVt0dd7lAwPjbuj23M7OgAEZDp7H40DpFG4Gup5oSjp/sYjohrdtNQqDTKtZxU90
5iNE65x/XXvGxKC4oYT9g7lAaVCaAS/XFtiPKz2MyXEe2rzH8bJ7bmvRxsM54v9W
r2fC3L3YE2dpv7xVXY7O2lOiJO7zbpZTHFeiCW3yFqM8oK6dFCXyd6lGbk0p8NIM
5x3d+NXfMeIL1mz1130S1/8AMykoWeosEJ49GV3SML+LnnuawpNfoCMcn7mBkPT3
9B89H89RQFCTeQbONW83HhcZtxLHN08x1iQSr6Lb2yy/xOcuqQau+dQ1OCK2Cw+S
ccHtvnYofoVPOgJmWlC8HPUqW6TrPJHCDsTOpfCBj7z7hbuJnwzqXAyHAjLoUSDb
qh2HDuMj/WPe5hXzbMCNzoNKxkthuDHrK4SPCCnrGr4I9cGSS+eSXFpyBBU90doG
U36xopliDEkJoR5ayHnX7RdX8J4ymWC7SLlEWd9Sa9Grot8PLZJsb4Qi8+MiUYKm
WU664bIrTSHOYaDUvosmsimgpcSYQfxmfCcmSqZLWqz3Sz5W254dRR5XcYfUl35s
bG7c5e/O0+utVL6B8nrERk3KX+DIVNGCs/Knuy7mv7pASbPzBD82ZaajxLnxMUYi
Nx07P00kbBNoEJsFhD2gCw2EFc5jReRT8BlHik12bzJxEwPxbSPOSmgH5F5xuZHa
937BbdhhtZ+DWzc851GF6rfo5Y7fDJKsWTZhi7pIOf0VO5yrzv7UZ03vvC4uqD9U
dSBpX1qok0OXOmlhze4TfvoGxFvSvD/pPhb9Cu2RQxOUOgLEJpDybzC5zmO+/8gR
MAyD7hl6oLAJDS9VgQVpNzQD0bBkO+5AM/TV5Jk1KSu9k8MHbTmWhzl2gEgSvxgX
MGSa8izfVJcZqNUYBQEmEhVeAQRm1XAPpr6322vo6D2w3NHdzaJc0hrMbxWJk4xu
9C5lH53hF4vElvfTAKpxkRorJghs5xJg6RE61zJz906JZ9W3oKGrsRGHjKmbxF7J
pVq+WGeXh6sboI/gBnkYDNifWrig6jaP8DZaKRFCugRU94qqp0JAjVy3qJroP6Am
j4ularjx0TVICNy6ZBHTWhQBihUpneK/hMeRX5t7ceTe6UhMjktX3EbI76EibFct
AuoX/Sf3n/k1hxcfplis7l7nNcu2T8UOiMeCkXUjxs/IqEjNpHfpbqHPkfazWArv
92/qsoUaIDI94bm0xs1td4qkm/AG902nG30ENM5GupmI9Q30IbfJViIqAEflQe6F
0PbyIDo1B1EpWyIL7KkgnIcwLFJg9fVLw1bMwqIcNQ/vn4MBLP82ljTSXik4pmvc
YCLeER2pDFsyNNB1HCMGi06UJeGNwzrNaLX2bjNvddbhj5cXdjjcMW/+tgeJG54+
8a4e6EllRGbI06So9RL2VO3mW/M1ZBRkZF8MstAgbdO+uQ4Bm7VCme8EyuoSxO+t
tJJLea2JYayqmc5n1a44itLyHzFb9f4gPtfYZWEO/mk2MygO5WYZsJjajnIlLB8j
Wvtxmt7VtHcTBq1eMoOTZGkHgrRS3Do/jJTFV876vvpRbX8mCfGygjlMGJcvv/DK
dt9DmisomaT7CViPdWFEizkCiGcwPwi8ABLDmNe2H9rB+tmGf0ZSSxZIdwk+KJB3
uthHNAPNQYKAyNBAyAR73AJ8RI8QgGH3GhR4oRADI/kRcaHKggayUJh+kVPn4anQ
ObRxV0/W1XvF1C2ruDw/+6C4zukSzuMLmc9e+IwkAyXAzhrp/v1PM+1X7UtpBLAr
uUSOe/iJM9U40QaOL+WV7ofDietNKPntO/G3rKYoeSgvCtEYJlC+bZWEAcHxBpFg
I/XJAvzu0pVBusjhTgSqc8BGTuJzjbEGTM6Qajmg+4VOoI3EGAVJHo8LNBqjTNl3
f/vze5AW360BEvWzwT4BiCb6g3v/zMobGqpyRiKoR+KdfUCPEdu9pU9X5kLWxq1b
29MCP5yyulnSMrqBGAR6O8hdRGl5jLNV8TyaVLMbDWXJfHA3eonWIwrZk/0bSUD2
tXYrTkpXt/2LWeyX1FoTMlbzabz3hg3wfZ4QAbrAnvHyCD+uU4UL/RhOtG8QCsXa
RrTW2THSZRKYOw2ciRrTicTDcn6mn3iKbRJVvn+lBQgdueeuxTe67DfUtFrO0ok4
3KW5M2R5XHBBfCZKWGlTPwAwTdgPgoRIo/YrzCg7+5G5XNGq0OI6s0IyqKJSo4ab
R/kZiFUrGU1Ek3MLDKjUY4GM9f9JaPd4Uwv7NPPPuHyxRfnw9Ezj7pfSROXCcpUN
tBZcFsJ3f5oE4t2yZigd6F0zY+zguVDcC0+/QeWv/2/Kzi27aqEgcnvxcybvd8K6
jsUZwE+r8FJvqXAUw8GFSy+JPAsPbHM+Q3rp0dHmJTH8wWQKCiDeglddlan0Kmsc
sNYbtuDjYIgv5oHb+kgLVvrtivSRjsjubfNv9a4akmV5dR9r1nBlTL65GEw5CKb+
ClL20nFksYw3ojaG1vQ4nFB9Dl1u3dSP0A1egwRi7eX1XobSDS5C8323I+wL+xNn
j+ZP1GjxdUgsanCZvHg83Ma4OrM1NdnuFdrAZGBBoIgyGD7LnjqwVQkl+KM+s80F
iXfUuXicezdU6YMvby2J+B340rRaiokD7RWvqY5V8Peg2qD1yx08RflMG6ZH/2P2
WUfcTsqUMDXbtymRpWpzSGv4UGK7VXK4qygPwFtlBuX+EaH5K5OiIV3Uc7yepN6Q
2jGGoNbjpBqBhBnkNbzz8Kn57H0jxNAf3jYjXObcEOdeETgUjb9yUWgzMemga/zu
RI66oQJhozHTYJiJprY6UI54ZzDTP6gw00INy3/ehJ0yexiVLTvBwCoMmDvScb2y
oWrbW9CD4y9kuN+3/xlgMledeJ9SFGYeJ6NtuUlDU6h7RjA0I4W24UyP58T1OP2j
3hX4gkk8y6dWTPcOlvymaX6irP6kPp2c+9PlsTzZ7N/r2rEKP/ofK31ChYiqSXJh
e0M9DJ7+NfZnhzMP6sDwIQ8952r/2Ps51jMcFKuy0y07DQdvq7Rgwo7/4me5Wk1e
9tjSuE2D03P2hon8YQc7yX0F0LwTQF53tvNDpxhX8/6c8NO+LmJQVlFZdHBp4yDU
X7/+3qkkj6FBLR6HbGTIuKcdFlJMNlozIyeIexp7/pp4r9JGZ6AERH4C9Z/zFEj9
Ve0e3zo8jTW2V9HU5nBIWv6zSTe0ftWZqZVKYaxZvSnTGY/Sj0r013In648dsH9h
SvaA8V3siA5nayzTuoGNEgKNmC7Zm/S1No4xKVPF4JTPACmMibTBHwO/Qquffwn7
pR16JUEnoIUHe6ZCEi5N8H2C/ma+cmX+iMYiyHYXn+uhBfPe3pWdfq5epPaMJjmO
+BhV82AGpsBfWa2+Km5iB1+6TqJA4iUIX0gpcXpTBGsLU2UkhmKBSgBxs5E5mXJ9
5FL+mBPCjZwN7VasV8bJoJECfSKc9jodGwtptq3f99K1FH55k0okMiLEcWovGplX
2nvWygKYYFoQ1ZjzJgknlSPfPMSVNJ7KGbWbbLQg6UMBkG0XRlXKoM4LklVkZ7dW
nltB0+AMIlRWnQC+VtciFeUEjnR/vKpbzQqc/8xzlA5cA4IqpJE5rPv2WeIn9cJe
VLn2wmdxItVyCQKlo/O2GqjjrFMe1o9hJ8drhYcO7eTWQsbUZTkIbkXtV001eogM
144Q3oeS6YLB+STum1Mp9c5lFTync8GDH/AZYVFY4yPxanx3kCZiSyLH9JLMcEsB
e3DdhFYv5CDkg2pWt8mcQtamze0iGsavyAL+Dl8DFJAmA5abbxbOUMK3hG5ihh8H
GTPnT7uXs8rDUlxCp4BfvNtsiXP86oijSZdrj1fJT4GUVdtXaQOaqQNgutA4QvFJ
pUR+D3BafpASxzkT+swOiz2z43P32KNPu9jibUqkU5hR1A0jobDNoZBWWTzkhba6
ANDIF1QjsING5JGTvx3XA4ndafe780whPpGAfT4cdaEY7vSAifZrXSx/srt7928V
5KGcA1SYGWtQV52prOJh3cikMTItPuflts61dSue3PY9gLGINLzkROL00fCVtVTI
0yfIbsljQLIuo2hkdYRynFBl07AQfs1cUJWe08/Vkt/J17IWJyyooDMLCk+0jobj
Ot4UeO8HgJrM/cefbbWkxF3KhRbDorgF/pKK1+ZMTz/MqsP+m+tp7tUXXjPzkp1Y
lC2eoG0KYOpPjvVrU3KUTfqtYHyT7FyRXVL089Mw+TZTF8bWgSPP96dQ5Cku9RkS
OFhY6j3nqi8X95OLsM/IyWmvFInjO2zeOnrHjfBWQm47+mAPxk7HsYDB0Kkl8GAR
arqQF5QMx0x1nFvI0AZIBaV2AJeiFa/PWa6k+VN4nvncE5STDizgVDuTbf+24MII
MefThwhTAINOpMxnnHBdZ94V77Y9UvO4CD4eF3Xc2a22bq/QZ6CIGZHgM1BEzBDA
eGi535bdBRdRjGAglUMpFylg6RcwvxsIYQzTjnsm7kxzVMFxVTjz0/OSOpoZYEWC
Wh3yLODclYKGF121PWCVLaLOrP6xMDn6CLfileqdHOCZy0ZRqU1r2mhpH6S0KOVH
+njT3S6hhoYE3b/CSiqHyA7bMkC4vviTYdzkeG/qBppV/brODlY65nvKGRzq+bUR
DettWsr5pfQu3gJuUB25bs19R3oYgqI3DtIACZCNI61DLdg8h7LLQTSTb+Rw3NJ0
ILJGOJPwDpXhqRfYsv/dj8AUR9qp/JrdslzIRxVsQL+tW0dbD4l9wNDbrynF5YJR
I4J9gJzS8ehuA1gbPT4WERu+QC9SjjAgNXtv32aGY0Q4G8LbCkP/qFaGPspXYEFS
6tn66RieLQTM9oXhzzC2cTtwShfs9+a3MHfp9P2kdTmcXDUtAc5DvvcuU9PAVxOx
PwnhOkjqftErJwQnR71GaUWy9LXcjWosKSZRe1TjTDZF0C4Zs399bRfR6YKSmgwC
giKT0WGwnn/hZhtBH1Es2frPRs1XeiLBBD7HgSffJ/1M2wqZUscTt+IOCIWEaXhU
6O34FYEE/0SM0D2ih021OfNLkbok/Lg/1lJvR8eXR7GjtR2QvjL80+/aiPvN7RdH
2OTfjpnsHZMWHXYHkkrdaUy7DW2f6a72b0ZaMpwFoiw1n4aSTy4afeJ78YC4cAgj
z7ARwhBV7UrjKIcIQwbGeZfNCLQ/0lG/MLWU9X69yj3F3cBtz8JU/Gv8D8GRuheT
9EQ5nn56zFNSrpjz8mYUbVIg+CSfNozN4yQkontCUn2wO5uMfbaQ/9nrb2/VVgGS
im7QKv4MMqehp0CH8XEao/tUMycfsvAvdkle0hZkrzbS3SWwE9GBfV5lkw2KbxDL
AUIwrx/44zZLc37NbvnTRChP3AA3VZ//C6X4weetpusjuiUqopkkw0A4IEkIZUYB
dG+Oe4oIf7kRQP6HPbta7StRJkyhLtNuRlzSLAjCPVXAhRB/NOPN2+MlNZVW7wzV
pW3RBdRtYFRNUIVM7pb7RbZb6UjxzRRNesDIDHSXlWLny85Q8n9mGMfRSgQe+LIQ
EFA7YtU/yrncK1l8WstvSEatNKbKpkxerNhpcmZ8gjq4jVhbjTV9tAKZoA2P5aaM
YbyUd/z+Sjt9HaAUsYd7FiFND+9zlKSS7ls/GfPknJeeVgZpnhQVXvfvjN3pkxhU
QXCaPXFhuoB6AyITcqtrCHpY4IU8hA8H0YpdMURq1wikqxHPUeyQqN02YcT+Ktx7
he4atmJ8SYTnUqdyu0BxtJaoTJFBAPYW1DUE+NcpvG/ArUFIz3B6zA1+sKTOxty0
lo+621B5psBbs48p1BVkj4Tvuv66QoljZhGNUF69x0jRM+5Nqv6QaoS6SyHVy5e9
GVGcFpSJjb2/XPsx1LtH13UcgWqLnb2hzWb8xSR7taWiHuQ6H/IKYl/poNESwx/U
QHbZCFRtWl4OrxFnJhx+PcvLbCut9qEcGit0tWZboZ6fkH83AF6x5zz79nhCzgQt
7xIl+U0yXOxupzuad/THHwov17JLW4MZFW6vNKJ/NCnA3GK/5jqW3LdsQ6zFdDvw
cLScDgBnmTUod8rjxpoQcRxUZM/Q688VNsKcIsNtLSHkvNGk8YnAvEIQDcrO/qjz
MUP37nB5fd7naVVvdOgQyhM3b75JclP7vRxmwPIFRLnnqPyaqt+HQ7aaDkoX+5ig
wlhfHALmAwRoCATuuPYzE+YWwsX00jj8uwd8lqzhowclwUN7VV6JDAXTDDC7hxBR
1H4oVYFzRsRWVsJ1Dsv2fb7srInYS6oupNZ4+XF6Wt3qWZErolsbMcgFcETqvL5y
zX+VZmUXprhYHFwnzGLY+TIQF4VrG9P+lgoAUCuSRA464vSyu8NpiFaVrA1G/LN1
00Nooo+vS+mDn8TKMbEXCUS5u7BG0DInIQgj7GWR+KBXgutzpxYBo+RLxmfGvKqs
TlZnnMuv4ccGb11Hih7LowIJpy3Bl7cf3C5abZSY3BcXnQORWMKFvxHGWHugRVEC
w9G3WlKjhBoo8/cwlaYlAP500CUsi6vqnOAGUDbaw/ZevR4495g4fZPaptvaaysi
kUO5g2pP/+TXiZPy65aGbFbMBro2u/eg3yKpQ8bYb+gJZidLAFh7RXe3ysksljY0
od9WtJloNG8YZdB1WHlfiSFpRwZpb66rBKFHtZUWAH6LYALjy/NTvXN2rCBuZp05
KHtzrEnSZdDCEiXi+DgxRRovjYa7US+SBVocs6DcIW3Sstx1TYXjFSbUsm+tigV9
zogPIG/LsIpaWq/S3uLKy58xs4q/ICUIMKcpZWsIXrh3imgi8ZmBGhsLe3AqSS/w
XXmlTHYxztnlMchIcpXrEVhBP0uliX20fPwz66QAx/Xswo1qHsn16x4FBVWfMF2N
xnUGrsVMhkigeBcSy7HfIsFggW9DjzBt887+NVgRjFBbWAfJnf2Dg79YrGZ54YMI
UtFGcUfnhxJVXeoLGb2XHuGpV7zifATiPu1zjHRIMM/V5WABFfhH27yvfxtuLCxu
pRcYbAFkhHrL/LNy+o1GCV52/EVVgxXr6V2+heg9aENqKiytqym+0K1HX7u+VI1D
Gbzp7CS5WpWNV1X5zO+kILfSY3TuYiuEv1Sm1Bap8p5BlQpM2rQTArus1Ed+Kz4c
yYN01aqqmYYSvnI3n9Tx3hh4R0IkOrMXd2Ii4j27wNpySRnyC28DWGxz+kce4jjl
xXfYMWA+fb5di8bIJf3PIrxxcn3acVCFA7FhLqPebRxgmuPcLQlYXesxej66MgnC
ED3B0fCOMEX4iu79uBYizd8Y6DaOVIKNJgtoX7yy6/9n0NQkjrXHVk+9tZJ5aDkU
vb+Cl1oFBXcrzpZPHtiZYomv7AifpYvQbc8jAm+pjFLf2DC+mhl/HrRyes/W5Kog
gQvNJmpbO8vax/xiAu27i5u5qDYEFwOe8oDSQ8RmHh0q40nfFc900j7GLipzbonQ
UkMF2cq3YGiJP/AB5NfobNjbqhxCd5F+3tG8aTqdPvfWo94JqZ2kBxdWSx8EvuSR
avkVjT6PF5gW/7VBnB1UvvrLPtDWE5BkZ11eJZDDm0HvvE3AV8EzCbnrHtvU1HIK
3911A9VXQSnAY9QsMiuNruv0yC5JOFn0C3yOCrkD4qn3x25dEokrxmIb5hvFPCMr
0letaJu7pAMix0r7WFrXZZziLcFaW9jSMEboHQsehirdhJMGy9qUijjlZ6s0G3d8
+A1Mfp5P+SeLs7QZOKI0y8aoYKAdIlnbxIogxMSaNuQ8G/1n4V3QqTd19ovHou9z
HzYNV6tVILcfHQd1iLGwC2YCAbaXoteF6Cc+3NoDyHMxrjmrPuIknktDZOMQjt8Y
BUFoYB44T7HzeTM/2SxHYGWBlv2/9bCZ7gUWgV05bQDkPMAUbD8L2dN+e+4riB4o
td6yOf8ysJs8/7zSK50I9xxV6pMWxx0+1wjP5lUVWOTzwWJOephOq19CxW7l4Z3p
4mAXFn5FkuefUbA8Cihax9QGJs8BH8ZWoZtfR7CHxV5vcwZTlFyF2Qoc0rWFqCr7
IjKYFFvgipoPvlVzzOw/raX50IFjvrz8ma15rj8Q0S+uG9BY8Grazqsmqi9A3Rmv
yqwNfJUYfsogBPNZ19Ffn9wmN8qbphHdUVF6GBAFVJSG/BcDoROt7EXUkR50RMCr
a8ZYtkRyFiYw34IRHYtZtQvFQSRbXgCF8cgaYjo8T975l9/1BzJbVFztYQW7Sxh9
yhHiUXmIROrCQpeauu1Qy1xc4v0XXt8RcksKpl0WYUJnrAU0W34t8ULGLhCf4t2D
oxhUdc+hJv/iA9Kmb3CSfBL+XkzLRkERG9mKby0KxE9mvBE6wEaybVe2PgmkKK78
4erVGTeG0RXcfjfjwKij3Q/xe0tJdbKmSZLUONTNuk4hiNXWgzUlU1va2JUC80Rr
Lb/mS9iMvQuTpaIPqqMcPsOgNg/Ff+ryy6dxImmmsaCWf52bDyVBzk4UgAXyZZI9
sZqAlRfXlRkFuvLJFQLO/gjxKN9YoESeXGS7dKOGu1ngbOSrrMgWReKENKqa2H4b
Vv3vMb4REmePLT0Ll9qNjmH/kdnDP9fONJOHd5KOWNv+Z7ksUug8ojZoBT/mW1xY
2kInueX31IgOfDbeVaq2heiZtR6pKefuLCEEN1x+/spXp1NgiuF6pTWXebCPCBmD
tFFgcxjfaRk4smiMaGlC8/WRmhvwuIyDEcFSDfb+zYAFEuihiuYSuFBewTXuqH/s
zI7h5e3BqZ6HKCrLykkLRbDkx4O4b2yEVp46E6fIh85ahIPhOdkBFEfql5OIU0nL
myq8LRyaJjdC9F8ror484o/WvNvUS9YLAGJDvJrtMH9WVQoo6EKgrAwLy444BNIz
pwYoHS3sf43e8pBTxRvQcy0H6h5hAIz1OtigLB483bZszKnbP22XrA3PRpMZ3vfB
gnYE3XZw3/4B8uEc9vCJ2eCbLdid+6x5jrCIwWlpsn/zhJp0Em2f/r6h2l0Mh5tB
qSXihUWPEALPPweD9jjny9S1ROkNZICikoVEZO2zLFtvK+n6piMBAq+jeYN3ygAi
C9kbrxR3cyobvPBdai7NU/lZliPh93wEIlZdTInuEv8dG0PBJJ7CKuWrbkuX5idA
HyM31Og/diFBhuZAWDhnSjI3hKAb/Do/fYdu3yiclEzb3ErFzy+9RFCwWO8giIBA
TPeG9hbGkHjiWR6Rv61DdJ4vPjcqBXwUuq4fjNhEM+QYK3j+v5RRvmUZbjCNZ0PP
ul/2RAeL5vFeJSNg472CEQGmr+19hJxbpVAMvi4ZEJt6oaeOKJToq9+v5rHOwA9H
1F6ST1wHx+TOgEtVQjUKalhbIuU028/XbQ9HfoCm7NamKKIAGNQDhyAtXtf4XeyI
MBrCWXI+yReERJQGPFXmxvRKlJOFqtuWdqbxq3xzYmR8zR1IW1vbvnofruy6iJOp
gu1JR1xDJGnBtf+Kici9DG19trZR2AXHlcqPnLIkmt9340oxUQBSrT1KZL8uuD8h
OrswD25U9aEYVlegHGmGaoRJCHkAebbHqnycA2DXwmgGGatiGLS6suTMwa6hUFHR
TXZsrYrClqJ+ZIguRArKnxUiThUasP4Rraa4H7BDd08vzSmTuGclL9E5Pfdfzhuu
19YxCN9oEljlgK4UngsTCYzUqPQXUZZmzVPF0+BPJZp9Tp95NI+4Xs3FskLgYYXd
rOWTHITZ8wihJYuRHNvHSiVWd2BpxHekx9kMGoxEfpj1YvSSinabPXkhI7CcXOyJ
r3MuEufczdDvdHJ2mq0CrzU8ndwRhiU7A+FoblTIgr7uqO3NxfahuVWHLxoApw9j
nOfTgrphd19lNTg4EXpBcxZzsQQFY/4h5AEdEE5t3HAa1FcPylPG3cOB/8G9iQ6N
dvlkzBlxor0j2dYR/dSGsCRXO0DmdP/wipphnXV/WxkSuN4AH9wSU2EYrDMKFJaa
jsESvCoz0vTj3FSmDaIpjkLuLd2OA4W9Nyrdk7V004rE4TRjGCyKZ6u0KUYgaEGf
Eb8sXUyeXwsBwCqDyjwtwegW8zaG7CL1ph3KF9WqwcC0frH5XlVuHk14gmQXK25U
G4rHXfeupgZu00dyP4eHNI7+vh6BGVB4SIAKNM0d4xwICguEbl1m4+UHCdX3R8WQ
5ZpjUvdPhCpI4RY9DCOf/4yw6HQoz5EhqmTfh7Qycate8Ic1bHbVe3D1Qs+gmd58
5QQlTzI1CYzWB7z2DXlx1aDsqfw2PEVaj6jsN/0W2lDR2V4g4qkAli9B2qgYY51+
zLJSAl2uXuUTaPKj8SbeqvRksNsDoVFy9mzGzZqupQQ10wyIyzW9QtSJjV0LQlQX
PBdyHslYj49f3tJjQLA2BGxdWD4zAVOIEJ6anL1kMtbCJncDTaRKixIKfUBNKoTv
dzJkUxV42MnPehpJzgkIkPTG79iHfC/2Rj6MZx1wIl3PPEM/E+Ll9d8Ty+f1p/7e
4clSEMc+wpf2t94EqG61ZCrBg/2b6Tq18T1jOCjAgS/l5dmg34YaimykodMo2FYw
2LtcrHLzLQnB5K9ndobB/WauiTIvB8l/TYFb7A62rkMHYWTjJchEexhNVpairjG3
ep2Vr5LUrIAAJB8faV5MK0N8P2AtgFG2GhyByqPQAKfg1N+5jPzt6FI7bU3OQ9Bt
K7meJIZH511QTwWASozT7AUABM+tXjwfXveDFaEukCJsxURDez7FSFeBMWbZQlOM
KXpfVpQkUtIE70o/ZFXpR/kYP3iD0a/z4U47lyNwjNMPYjzNCivU9h0hrQhfEKYO
uy2MhGWelOUaqPhWyzooST2C3L2Ez55pB6zwS2OyLsHaeWkR+1QUzGnx/dcteFSf
gdYVS7r2G5FqTFTQ5onE53XEUN3K73QxGNujLK6qnXRH7DjqxIPNsQ+x/lhjrDqz
crjvu7AAYaXbD98VYZC1B098kWgDZy2nr9ZlSVuBFHSh0/+xGxs29w1HRwDH81Pq
6K51wCMP5eafN7dwe9fLbzmN4cbsmWKfZp4di+aw9zbQAw22/Bei9VMu655ibkmZ
RkpIruEEKveZLb+dX0istWpg83aYoyXGiZhaxFrH4kQdAOTyPp5vyI/PbeRq+4Yk
yzv0lhEIlKRpNz/AljEo0YoovVMMxGhnJZGZGCx64Rsuk1NMjch4Hkg0IvF+Br4h
419I3J2B6hcKxVZ73IAIhgNGoWF17IZroSt85FE0S/xu7syTLcol7xIS96tQ5Bvw
cJXZreaVRKlqjOHbDkD34GWXHPrT1pKXclkGHSlduazMb3f71H+eAzEWL6ODpc3t
E2f4MCKjZRynC+IN7yzoELOugCNVa0v1clyoSni0f+IPpkv0H37MJLrgFYYON6Vr
nYJYwx2zrq6ZhzufiD7zrqL0Le3kVbNx3oM7nmbsJrsMD1wwndTS9kJ7nWIFpyjX
wdv7Zb4VUqisFJ4hWI5YZiZqUAiUWlRMGL0TStp6spk2Wdf1d+oh4B65C6weIqDF
6NvVAYM/SesUbSF60+YfrP76EAz4Wr00rMA73MTz/W2XkBQ4tW/ZdZZwOZtrhupb
gPs4u3cRBX6LkGHjTOxOl3B2b1bEnN2eNAEyM2P5rEuiCfqWCeP3EIB1LrH+GvWy
nyi1mOnzVF8bBwE4xv00kzvsNGszBor/FhEh4SbQ9EhFED8PxX2kDsQxpwSo0kCw
v+/JaUemmXOdvqKIAZTaAlrgIm27PysnyTBDzBpXkH+XcrsdsFavb0h8nUfK0L1O
3iq9nR+s+Cxit5t8qJfG/8VQmksX+NSKrKLHpbuIX0nsV4HrkMrvRMuVT03iku9I
L8UjFUH2rZ4ZCxYiqkUb731Zz0+uJIRrY+6sJrsxMmoV/UHRYRt2sSCpxClO6Q9B
mm429oGN+/oMpBxIJIzceq91sV8TjIF3rrWwubqoeGrPSroeTwlKgXC2n3mVJq/t
J7msyG2cgfMBr/RjyiuqWpEJTVUhiv6TGXjb/lcNKNtpU4RaWttnpgxxqm9t/ZLN
UXhS2OR4oXZuNqxhsfSlhvjTQs23UZNZFhCSbwq32IGO+hgfJVEtdyjszKZOCFDN
woYr8+43hA27kE5tnzl+Q2i38/c2PM1OUvznAEJr1WJsf9GrLrVvr7kVSVYYAi7L
tH9/0mStSmJkriS4f41IvyAYPQ/pedLOBreJcEzvmfd+igHp5NFAn7/Ew7emvE+p
YjrfECrs1ZyiwrklCwGlvqGQWJzPZC+zawfRTXJTfRu27Ee9Sk7iferELVx4rhjP
39Z2lkFYy4PA16kkJuUdcBDMVCP+EkGaHVadJ9uFlGhQycAQQQ36VLvaPImG/rTk
aHRhhgBO2trR5I+UWiZNaed9YkBOHyB4hqQIknEcMOOGfQm8lUwszSpQXU0v3mWH
6Ckx+7SbJYdG+LlDMqX4sazqiKBKFfKRTucrmJAkdaWYdm3V+RxrVEBh/uUcC5z9
/UK8O+HtfrG0SRKoOsQoCW4mKi4z2uE5G5OQQUNw2HTG3L8Po0Do4VtYiij/i0RJ
7Um/Zu9p5LZoALQkdEzNSZwr5Kc+x+ES6XMjjdlrJZP1IV/IOsOzHzc/F1yB7JQ6
3yRCdRX1vCRlE3GUde8cnyxMsYXZSYVEz8WrDjYeW0tkLbYNWEnzw9Fhgzpn7jF0
oux6stibCxLpgxyjcxRqjBwVPkYItIiPJ45v3RUhojLZpCP9bQNvd7Ekfariu5FW
xir5yrwTxaV26RlXS0j8GQUCaDGRpZjNrVfARjMEZgTKTQeuh4+fcCNzK/RU+yKv
f0ClWTsT0pmK2Mx+W4ymk4wIca57umbq4Mi6PMvJa0bkAY3dQY1hsXUrQBq07k2n
ZdU0nnCiYp0ZORHAEBiwoTTv3zcqc89Y62PiX0ruoDYwj8y/RfGTgmmt8m5HXoWD
5zDEDCTXay67+gE9a4gym3tnpd5OyfYprYSLO1s0F5dMp7wn5SbH8tDPHt+TLHzk
Pavk8OwaeRknfUVxIu7UMt3h/MsrNbFJYSXbT9E/bi4LqtMb+zbYh9KBNBPt5FIt
XMpHLKAUr0euItA/NmuSwkk1bqZhjJyVDliIt+1FeNzaa+v6AJqPAWA8YX/6csAr
IX9yYMblAymE6/MxTrASAZz0cCwfOLRlqesorrnhEBVrAywv7E+HdMJOpxHPou+a
rQcxlbY8hPnRCqhYfGQwTzhaAoEfawAx0sxjQE97e0vFUAibAO0WPtJB3kSstFDD
0KVXTvt/s+k1UPq0w0psIzKf5ouf5FWIaaE6z8oRt7eSs+zRdOAD3GhAU7LEcNLp
rO1G5HIJgobmjCYFoF+asw1aMIzEvVyBx5Jhroc+JoqK95RdIruhZlsh8M0rw2xL
ksTrqDhIfxvtPueP+bP0JMWcl6KPwHctP3iHDCX7hy73SURFcdtZTgJXY9Bo44VS
xddByNwpDvqwYrGWo6YM8c/K3/2Jp6BGl4pET97pR4DqVrplrukQGCzrQcmDKZ8H
AB5IhOB6mnLv4PqppF508PKRp2FJFtlLOlkUOBcb9qz9V92VoIay2es2QcgD9E9Z
Kh5gVl5RHaakAKe4hBH+d8RKSQGnPcGU9k1JziDo/xSP2T7+pj623aQlo7v01nHd
vA4Ev+sZ4B7T6sLcaQf8QCFth+smNUGu/6UioNaTdPidDpGoXzXpUKY4ZDIDqUlv
MROZeOfsWWo2f5lBpC2UEFStj3hjLtQHhpvaSEfTe6wOsoy8CaPvaULuIeKlySUx
pz5xBqjKY4OKNQVaWaMbeZU1e2Mkrl1odNH1JniU/HheaWPavFc2xVQ/rKtnYnS8
O1W592N7BU15MFQn8z8suzV4HdtK5Gy+MYD2zfl0Ku+slJE4gVUcRzPeen4XiXH/
Aiy/mhDntzrvvjUCx2AA/cxuOZveoNurT7vPjnxB/kjbd3ZJBJWvQkF/9aJM3Hh1
npyV3jKVINsfK9sE/zfTW+K7r8FThbMqH8E2VVvjp76n4QEp19dQOqbJLuRirILC
KhhaPgr74Hh1CR3ifONGVf0Jktv/7DkPqGbAI1z9jjXC3/EGFK/kgsetjvWxqI+m
ZYaPtCDXdhx4EePfb/eVGVH5Y7Nw4w89yeJzxwZ9I8EGjrtR4QbMfgXFhZXfOH7N
bgNDRS+7CRGC7khv20/iiLDPV8k0Hl0QBF2FVLNKNfKeHrT7R97bwOOW+YVYkhEp
LjNMmwXA+LTxYNrEbtgmQCzr6BTPq07kk2VKLTmnobWrAAWNGl3UbKVaQWmphqYA
P3EpZ1TqqeZh10U73BYRe8a5UCZs74WV+Du/Erith52tobbOEHt7oliSUto1UBIF
QOghz2BbunxPuX9LDYAP3JwVdYiNjYzb50HG5Szhxi1E3VecgrlNLeoj0ZqIPQKa
MD5YuVtK07g35+vYmMTESZXYPhQA/Ea3djxCQ7ZDlU/eiieoQu6d70zTuuiezsHk
0uc9mRncclskYg6cxUfNRbGtPjTwLeRQu1ZWune3ub3mQ86gVIG7VKroKXbHWR3p
uVzOR+nFwDbIE4QtWpK7cAkQtdi7ZGN+sDIUmfEtk2M2hVgagb+XUHEVHzhXdoSj
gDCub4Ao5Z559RMJ/2LC6sPjeyJNM3QOTMmT0zQ1FXkwhRTEQ0/YmCKYVOVIMubm
yg5gsW2wK7MGaUjFUk2//cdEJyZZgRTDmJGk6Q5OZ01Wy5+pvtOAvcq42TsnaUvD
Hxvis/X1vvn9YaqI1uspukCYd46/F85Rmn2T+7RWsRLOuqoEpRv+5RtPKAkhjUAg
ZGvxe0+8l3fz2pg8bxKijXVKMhQ8qBhxd0umzPQ7LiZqe4kewdK37ID1KGnokV5u
KJH8KbsqzNCB9J1yIbLPVcActmi+NaD5+j8Jw6craci1l/sVosJ/jFL49+kGRrC1
/CHBhcRzJU9NkKF6SbaPF/vxoliFHNR0AqJuyi1Q53B2LE6dJit1EOXjP9cJl9L6
fffT6P4ST2/Gys3m7NStdfOYXj1vgQvbk7XRbPmIByEQ4OL0/+NngoEpJLuFUNaO
NIEKu6oUawZ0gU/K3nZrhMJqc/enlpUJLEqOiqBtIJrCfJfQxMADK4YZXPTBckik
hni56LgLX6G8cYhC6vz94fFGTwEDZG3v2OFpbHL2RFFKyu7biInBG7wgkw753h45
D+NRdAyH0/stix+dOTLlYV3vScGMVRTWUEubrDLqJ1WJBT9Gk5ibbPPYdYHCRXLp
OhMzUrJbsTQGiJnrBRRxK8LEtqks7RRIRGMl9eWG9YpiV5NtpKLY3w8keJoARGYC
HV58RjHvbEJ13+JMEHC39kkdxjTq4jexT89w5nzwRQwigYbqYo6YBkHFHAjC4yiV
Hu6UqvxDXkYLOqtk5EdMDOyMbWuX7k4TJhHVfOYbfYYCULLOW9Q832AuVEncexJl
bNBrXWHK1eXdr6MyPwb1dPLd1QjlqavjYJcGwa6oOpUBa0mf0GpEC5xpg0n39xp8
0cFt+kCg5J/nBHNvTO3BlrySl1kEFW7/SbPEhyWTcmPanJ117QuSIubA5Iomk0Rv
bJnnwym9tg8qXVOUUlpsWZXJXempxp5wTKmdxQ1eXO9fsDACQRrsjAumKST21dZC
jVwN8hu4VttGAYh1JnXpnTyNVO/Dt+MyzA3k3i+GPt/j1DbCV7cJu32lnkfduiUk
Lrq3hSK1yR1Q8doR0Y1owcljIludFqcPDD9H8vdBJA0EvJrt5qqqKZknZ5G71s4w
wr5ZHgeeUtC5H+6fQH9uSOYo2b6avlYLGd6r8oWDFziowQf84yxTdBBqK9O2Z4Gv
4540Bcwmph08HtvONlgMajn3sz2OJ/Iq5pnwyxQggd2DdJg6Y3TCfr7b6GqP3Tsl
ImQAbJxTE96hza6fI+tcP4CLhO8Z7e3Z/K4xSB+dh7vozeYQ0e/0vzjQ18KCEyqK
9VjyPFw6kZUuBXfjntQ/t8UWtGUqWAN/8QFeOjQWiZmhOt23J/bfyL5BtL+vx9eQ
O9ik8i/GrfL5icH42JdUL+HtVTqKPpSTGBq6EdlfUHHTXGDCpRe9ffq14hJcxGPg
HK8ZII0+y7kOo+8jaws5OSOHJq+aqmTit+t15K712e9tfpCd61ZKhIsXoTZ1cNm2
10NVmk6HvmWo1+fajbER/nllTPxUpRtmqjCNPoaNZwBj8LQhOoV0DncCLnHIUikn
hXoKVITnZnN27+++8eLl+UcKA5xuFP07WVV51CiQxtcMEL3wAc5mG3u5CjRLCsd2
n5axrrE92jjs8zyrS79C/ul6XhpRFBB5t18mV4BY9V2IoQEJor+g46q337gzV3p5
skJ8ApYBNCNOEkUG5yVfbWwfxBx0/je4GDZk2JM329Z8pF9S4cCc4Im1y5uB5dxZ
KZI77C7ePJbIBTyOA+x6XUHddqTZInTpULm0e0glX2eEQiv2ZHvUZCkaW56ZsF0w
ufcRnOHZfK6WdeUry6Ny8izixdP1GqL95HvVJJUKMz9mTl4BAVMcf4APdjjCRCpm
jQsoKYq10JvHJbkhQy3y6+NHQiuVq7SKO3ab9DER+HvE6+w5VlfujeXjvDlhGIME
2g6U2IpwjWQv7K4l17PCtYLMEK+TM0Sv5xFnbV+vylAA6e2rt1COPGXYjMc6ZUGd
usW8upzUwYozoOkngAP6YbXifpiWURlUIU6lCVXkGytehyuCx4V3+91MUKL3us+N
Ub7W7wJ0dG5bcgISuDIZ4bLCP32I9LrsE/vPbyyAw9f5TNL4Siz1bgRM5/q7IoFH
tkPpUmj8o4geuAG4rnvbnSjxU238nf9hn/s1etrJ9xv0PDr7hLdanbhpxaOxG9Tu
nhPBJw03flLTF4dBAtMDmxckIdL8SR/WqdFMBOEgUhzsT8eXG0dbf5kFA4H5RyHz
k/+yV7a7feUnCm19RTPCrLcCLQea3s/5gHRwpyqkFm3mhy6iyeJQuziuTMrKu3q9
RgXkGHQDX4HykZTrVyt4PdQMQ18wIgH/9pemvwzpzxV0Cvw5NqieG8H4E/q5gEn7
F+Da8voi+E3V7olVd6oD5Qw0rdFLSdeyteMu0pdA7gch/BduKcoBm1RQ/u7fYK9J
nh5JHiAZtN6NjLff+XlWCaK+od3uNMMh8vuu4JuHMQzQy6XSpbVAd1GOQ5TREnHa
lTZAxNGlj+ZtJpuT9JsJBer4ayrH1Ig4lBNRgk7D05fWaJrogSyaIUEtbP8eShfV
s4tse8T+LF1Sjp5Yrtbb9yuxWM4F9+/mcGeg1HPbMq52jrQOVb0cHk/NMHV3xohT
CENbLq+GRy1xEs5mRmKA5XGiMBp9xT1gIS3VzkfOFF6feIpAN+aQtCLLH63GubTp
cTtJYvqS1tPfla5x5XD06YnP9iyn2uohdbEVJ+Kl0AX+dVUweQ+Vk9mHPFMEs2fN
JvYabVslsmfHr5ZrWW8SoETHfM3QsXqaGyYWAogQRQ3o0wyNtdeqKQVyXEhHzVD7
Zs77I4++TSiPkpg8t+fBRBBFiHwfGpzgrLEw4+Tap7qOQaGCmFYRnDHXMZ7ElqBd
/XyG0zVdu46SFiLqPhR8uAajA0KpcoEhBxL5iBcT7tHikkHqEtcDmigKGvMda5SK
M0aSmn5iVY/0d0cfW1g2CgZj0Wq4T8oMxfYHN6G7v7o9HJw6yCgoxLJd3zKRZIFX
c3TfOBsi8RAKKk/tYmx1VlbWnDpHpnHotvtoc7iGevB13P2LyRg+q0PAZiJ6OBMt
83OIZR6w5jRuMplpWGgwydTj3VvuRLbHoOubuJJEYfb9BJIqtFGgr4YQF7Wo6XkV
RVNLDXvbKaqkr4sroNKND04XJh5qZb5oKqPGtMJOluDUMxYP36RW9ikvUBTivlVg
9lLJl2SDX/JJPmS2O18ampRCGIMDFuuIl1kX+6wONx4qzSJqaUwPlbhmPa5xBDeU
N0g66JT0p/Levd5bdUPunIYAY50YnA0SjIL5hgj6Ivs536sUsfVS4ygMF9BNiLoO
qyekNrbdHxQhH2ZxM8L+iIrFnp21kiGYPrUCASSmA48L7lvnRzB3Y+hRlqjZ8J2M
xUS6IqSNhGNnb4DK/jsKZQrSRsof6A3zL0SI9HAYJk+oV4tupQFCaE8UH/8Z0KNZ
AOx9aCqHZAslsxJiK8mESa/Zkzq0fzZuKlvurCZOHsWQjNATosaqN3nk4ppT/T0C
aGLuRL3gxJ/uRZrI8CZ+s+50mZ6SyZRiyj/5fM7JEV2NYLd5oiLfapwr0/i+NgON
FQ81CfJrCo9YuCwXCce93dNR6TrqTzarSPgPeFeV2L1rzbSJVNtGrqFNuXUe6tAh
6e+IYrFvMSBcgg11eyGCREuEDX1duyfmMQEiv3XZfueBSukUyHXy5sWevCK8gEn4
UxqJAam5AA7xt+hMkDSK6wsHYiK7RbjRVWg0GBk7R3D2GbhxF5zb1T8PeyudOmKz
7DVcFYA1rTcAwSGFDTpXezaWu7B9HY2IkTo3JA2eK08nzusPGVMgLarMICTwSepj
ipdyquS7gkh/I2p3yk9cCQkJRJT1aMevnR1Yn+0kJI61vEcDXfPsSKqa0iKA5YZ1
x4RRr/z3JTJ7ZhARS+N3O3/xL7XwhPXAa2bYbwQrHPEpruomXoOMjmcQFk2mjwYg
XQnwsPluqNnhvwlRzgTYRtGaxdeGv/KQimKdpfWTugOkBGZXK8R7GT1nJ2ATLu6+
UZvEmUAwrvvoSerOXDJEozPlwsHUb30p3EOoetrZamcoN2ts/zKPponDZYKEMXS+
pY+H82kP6P360lbSPh88MaQ10syPjQC0lI2FFxsO79nOR8XuvDKhcX2B4MfPAV+R
1zC/5rCumVV1RD+HHshi0tsX2YjeRuvjWwK0FRBLckocluiQZnP6llAoBMp3Hvi9
tBrloc8JacQiQ35Kl8pX+p1j9TZzHPAXuYPtRJO7ckdJLrpdTn848LSIL8i8na1Z
l+kbh4DQaDQlYHG/II8QpfrCeFjWmHYptR/9WrsaltM/e1EfXENJmJuq0wKUZ/A6
5IpGRFTpY7cd71tAm1RaDz/LQdDxgEkfyOrvR3h6i6wmooSjdp7tzxA+W6kOqJwq
vfbRZY748VjMrZNvzsaWLI93g7YlEaf/0WqyNZh1N8xg6IYInYvnmUNqE94wog4G
DoiujgQ+BAnVl4wunBmjxffxTlxXMPZ16SNlgNXEtFjdjUqQRlg0WbBp7S4QBXIx
pQF+2t9VU3pX/E4+tGSITsxBmYb1bWQFUOcdISXmP9bWPgAkT5eUg0WIMs2fRQho
Dzqr1Eq/Rtv9BmisiQnDEMbx+dMsRTK5fqJS61hSDZreaM3zDL1H+cYZYyjod+x5
hd7pxi7NUQIvCi/TjNU7CnJW5nikXGrY+V32LZeFvvoUgM47NlniZDzZr1Q452+6
oQo4U1ZWo0XIY+/mxzv8AvRHo2ZHvh4NQIKbCyJJXwgNFSART2w6e8uhj9pS2Kh3
yaTZG09uKQPGkqmgXwP3/e3gLlyl4asVqCXtvgs7v1zBupRV8jcCdtDvsIT5Dt41
yt7FD7rbgeodjNGtmnIDjFcY7v1em7MgpG1NX08Pzve2eWT/kKa2xOkhq+WfZZGf
gJoEycRKivFX0oWK6K3wn8ZiSBkSYHrD8xyJTciuVbSPcQphpb/Fp7sFvg5y6GQj
YMBe84UBmAvXDlrXkr0tdyXDFY7SFNL8NmPLIDxLP9gtGis1sbCMcohvdB8YMxhh
SNAIht0J0iOXL9bg6AuoKaEeXpY7nClOaDhybUIM/LDytI/P2JXTfLHx+PzVdvd/
cyeDzkja2A+K6k09srV6JrRQC6J96g93mDBS9umivroMIJOcEPjYo3Vuxx2GIRau
ggWhm9hLP1E0uSmz2Kcz2+ua4izeou7QTgNn9YOVRKihfJpJLNms3uFnPyZ5fOkh
ZCJkotYPTu77ffXpZrQL7rnZdc4zowbaRClixiSCDsldbcKgu7wRGd/Uxlg0Jwxt
Ow//trjCvaTX2S25pnCUa6gX7Xf0iUXrVJ4p5z7cCNlj35FwOhZur2yEjfxbqqD9
gIH35gI65XBbyEeU5kzA85UvfumaYDjEX1K7BVU78ukAEIudO23fNbkniJTS8453
FgObXpVo3aso5eMgPqr79e2P8G0ArkuBp1HysmcK+UrKq/FBlgVpWTm/1MUJ9yHH
R472QX85CXdiQWSe4DzCqDeDQZTOjeUdtPYQWzCaOdi2xATe4XKBo+rF72yEYvFo
hWF1pmUcgCDPJLebLAyTQuuNjfIs+gT8DhaDsxBXuVQq3ndt+ypcQmDlhe6/fAf9
sh4h5NBGivFH4xnZQM33F+Ebfx2txdIpYPNXxIKIhnYtFWin/3+XZQ0ixURWHmay
O151ZXFXzfRJmXXUPCphq7N9Ak8MPabcnSTzT6cPYrdQsO89WWlPySywp9yCceXc
FLuWVWqRwMmdVbnRPszzna0a3WOwjiB5vkejIobj3T2aOFFb2yox62rNLfuvUJZr
EZgUEQ03ujlgghG7HEr542CIgtDz/U8yAB1+XTpUkQPGka6AfVKhqYYAOoHbAvrc
JDq3eHes+ElrUkElTb+uZ9MXT5SNlqqi2nCljQQyUapk/GF3IeVqF28V7K0YzUwg
iu5SOTwIB63JauqProHtA4fXNyFC43LTU3hBezsrNRlcsrOWH1ksJeeyMO6d/Aoh
Bnbd9KCxUXltFDCUpQ/PdnKI90eloTIcP8rQpP0Ln2XxxvIuHvWQn0bKAungiTQv
W35CJqoM2DR0cLzmehY0plqopvT3vA3DHY2eHeNMXp0NxqyX/nS7MtXCrGpEyfzN
jY7tN09wduUGI6ywK5Xi/4iH0OWMb6t/XN+ztDsFM9dCXdS/T0ErSKL09UK+pICo
ndzh68BPsQLIw0YZ1h4u0L/nZ43XeXxVIyS38t3zjqxuD7xewXAlo7AZgRBtS1vU
6iwpzwuQ5ulw5h5BnxlG0rQx5RWKZZo4c9VaewdhbdYVK4ETUeww74B5F8m/nqSx
bQrBcQRh5/xhOSThVitk67yH09miitrHT1qCHHg21aDVewn4sWtZ3Fzr5Fj+c1LB
THUTyXCmnkplYtORkInb2zaqV3hcUS4QMKnQPVSuw8B3vQhUuaGHQN9hQvyy04hq
h3kqLK227ho90ADzZ9EePNG6smpd7yfKIYxB/vhhOTpU5BxbtgneRl90pbGr0I5S
gf7I0M/1DaYF0cgiaMuFp6HQu8wu6L2bZH3jmhOzlUTQZ4ALNnqT0EwKjTtT/517
s7qJbw+DAvlyZmqPcYxF6ML6c/KpT8NGbUrGlTZsOJZH1pz/YV+tpSXt/gRiHg6S
ASHoN+s6JlgfLjGZznCi/D78/iqfHb4uSuQxHgkvSeamBOUqJeA/CeeWwoSX3uEN
I2cUBq/kjFH+q6hzUYAFE4S8Uy6WX0rn2GGHeiB+EqKZ6llMt/8pcC7ulHssQjqO
vQa2qos/yVsOKnB64xFvm1z4TKWQJwNnXIzpFmaTTLOMkf6eq/cZ7eRf0yrUsxKi
uNj1ydFWWgQjaNuDlRWYpTZz2vQ5k2KSGd1L7ct4A/YGmLK/aj88IiSHM8USPy0Y
xlxRFGLo8ZK2+QR6kJYhyqHWTOiFx9MkaJaEROlW/jW6QuDy36C0v+itR4LxwwmN
rRLu/WEHimOonAGMPmNVEDVLXvFoa0t9ngx/+GmkxIih5dcOPFhTsO4ZZ7OYtjfx
x+M8R9HWMoIu4gjdskRTdzOMrwjCE3F7FTxQHLQYMEJCZVRP6FC8OUrpdA2OQQhL
YYg2+6dVE8g4FsoZ917+bP7jJJndXKADqshqUXZK4MogikqUSeXMUapn6ck0EBw5
EPCIRY2UflY8QPBpZe7JrWKXMaQrM58JThtW6WxNHD/HnEHsLPelEEWiJBaXFMTM
ba8tkm8FGUT+3sum5jtJayLcyfTHG0Ori0a6S7L48M3XhUkM1DxDxpvLz1636E+D
v8DMhnedWMUuLnVXAAIX3NcpowfaPXYwKZu34MwZmWs6inSDP6LqtQ1IjAQipgXO
f+fD4sUPoZb/dzu2eA6aq8/NietAO7Kfej3p295R9Mmcye3DpOf4wVfAC4qzPiKH
KFVVm/raLcSTRR77AinwQ4gfJ99jARHebtWWN1coyaqfz/0dO3WuYorP6UOMLlzO
qEs7RH+kopJPoBSLXMKRNdzckldFGgmZaPL6tcxXUSRV9bEyUYlpc/HSf/HG8T9E
OhN6nyoh9wvK5D7ReIOND98jAntEBinRQCwrlf7n3Rz4pZIw/aChxQhtXAi4XXo6
oRuZHQpjXneG3BO+dfMF8mjg3n1xRoESS93uFYFfE47v7EQWEXpLlBtSAaNsXpbh
u0anDJS31d7myS3a2mzmZXm+C+XjUed09UIsmEgi0RjQpucdaQIyPQVu4YoKj2HD
9fFbefQ+1meZ7MJjHX4s2L/sd7du7FdLxBz79bL7xq9eyQJT/Oo2ugncphDzPAzH
rZ54z8/X52qDbGurROfBFpjrxktlj2Mv8u2E0OXrUpaHrvQbarK4Fh+uy9AnOIHx
OePdFKUDL1soGBuAxehjNe3pBnGajWGcth8400eoYFUCJs8/xpm8t3aTn0F4WJoD
dED4rm+W2YAkpYdCyQtY00+GHw4emETbr51CdktKr8txCUd07VvGpbeGyaghf7vE
/rt2pHIbrXjDDGuPPEMmIOqnvsugpZOKNioW5JGL726nG6hPHd7y+F1a1dnfO2O9
8o11RRgRyabqF+S87eLkEYtBLJ7aotaZ/ISKJKXVmnv8BgcEPSJhMyC0/IupzGmY
rnPK2gXgrbJgTqDD+V1qbB/j/3k+8IOdr5w3k8ioOZvKJMOT8RmaAT1lHBaGIFNn
a1u6LAQrq2Ji2MFd/oahhUbfohbn3PlZGtGH842MaSx9k2Y80hgM3R9MnCmJpJFS
WI8sWJKzVsFufEkG2eNDEJ+sLk2LtVX+l/Kz8DZKXGgTEZvHCulFUnBBepWRNDkk
8M5uFmKltZ12dTrhmwZbWtvRhyP2eCAsrZmfRVbw0Ix7rV6ogVJp4IFU/mAawvXp
jSIkJPZD2n2TVvB03y3lmk9OHy4DrjhM17Uz4z2dTlruhNT/yBuFqkptBeSxN0n2
EiHQrRJnXskjfCEMeK4hNAlH6drUtrCZ4ZDgo/zu9Q3bK/zZA3ZmFaVEtNp+HIKL
Fj/S6IT+fqxhZqmtWOYfSoXQLS/TYiibF9DZQzhkFhPIvTOkLJlbqmnVkiByN34O
pDikUMZcJ0CkFPuHvAY6/EVMHvApbZAlcpgvEfuBKKWYCvmSbP30cFcNgDlBUp+z
p8YguG+L/MKOjluFNevHcFwnH3JCqsDpeL6j1yZdzhUKXr3qX16vEmS9aWKELSad
7xU341kedje/U1drFfYum322x+nu1IjtXRbRZeaHzDBppjiOH5wkIE6QWGi5QZSC
7yAq3qIK1kX/2trC8H7ZUVyzIPdYd2LqGu8/jfS/NiL+zZpasu8NfUDgsyLAYweB
tteXAJwdMSDZCF/yhZVgiYkYJi9jNBxLHOdS+HYOxikYYEFrjvanceSq8GbgHAxI
s2UggYuopvChK5i8ss8YbonBtN+DP1Hk/rj5jciaAkptK7yBRFg7GNI8XNyRbfdT
9QxASgfiZEsRbW+mruDV6mq/mLCWnCDGtVturlxwgy8aeDqx5wR52KSAevvlvrVm
IjJN/64WsOjjkDSIJA4Uq6rDTUmeIXYBbh001MQf5Mp4+Jdmu5lkw8sSggN8mp4R
y5PQCnixCGIKu4S1cdlkVGwUYUrlFnA51cMUiYb4S2WpQaT9SQQ+f94r20TE1Vjd
fYTXe4BbAUT9xkkOJztr3FdDfC5ZK0S2PZMzSfFkMMGrt7gYOY/pqvHvUktub9Ul
A3y2M2pEYYp2beF/7sC4aI/65FmVoeSjB74CAhcLvy4gh7ykZ+/Yin6vKT+ljpAw
HSugDkxRPNa1dx1epqCD7O+vj8HSvX+a09D84Jpp11rzYQSu1CnByGhKYP2b6+2y
HRBn8NOWrIcrhll5U4M9jmc8Tgb5aejHEp7LDgldLRDbrU+aea30Th1ZTFooQZrD
jY+8AabkyRzGQ0sJiBzV9ve+sssKDoPVlpfAvrDowA647T7y1UrcBzQOMvQar45P
NhCy4amVh867A2jZ6TL1r/zIp8jMe4O49cKG7GNkWPkOrMaVGZnxJIA/kkxPF8ML
AAmRMAdKKJwFfL8gBWz4kI2Lm0LwddENIr6N59XmLfMoats+7epV2Vky/TlrrJaZ
hO2brCZ0qvZFAWIucNsI7/kY10AATjsAlR2vL+dObl8ldo1N/NBdbtoPxDLoqMhM
Aqum5rJy30BliMjAFqeivc+mSA3iqd1V3/AMlb3ISi1TW2pOPvy/bD1GL7snxRVb
Ig+HfvrGoSd2B7rbwergYaLI6iqN5CjLI/XZk4O+a70B/e5i/ATvIB2oZAYPOKIv
uLzQEjLiIr8dUzm0tlrW1+rlc83wpZbQFWXb0Rd7uMqR50en2I8Fpf6PLp3qwURx
g0qOHmBSsraCrX9WBIBgpdtEu+12x6AP540KA1U0EgpSKodFEsFuW6fh/fzkRmHh
THJfNsWf1SZQa3dD2FkwKEeU8GYjq745+9Y8PW1x3kFtc2qh3cmdRYIBI4YIl0ej
RTNgx5Ep4wezIuvUVO78bc32GysSCcW6iLw6zDdLE9ZeNwEEFLBveycVX2GPWF2W
uIBXLNn+6kRXG/VTiHicjRIQJFqcYI/SBqiZQuLB1yFvhwNIc9KMDWagF/X3EWrO
+6ZXZuxgsVrNwVIlBQkS5/QABNsj+4tMyfi5tBXlA8hwVkpKt5/9S0dQ5EMzr0OK
CSWxHiExSpm0yH2wP6S4lXqAf3GzRgHNaCaKoYPwzKFm33E9ISxEI6ly+u5InPjo
dmz5V6h0ZDeErBWjcyoJVDqQ9pmVTmyXzVQ8a84nG4EewxhSCNvKxjwEmEH1FB8z
nOCSbsA3lqX0DewCuN74Ofvh+bxcQEVnManZF9qn3Kb6lYc8qp2kGkR37Wl9Eydj
334a3bE1nimLqubts5NzRtkFwqjv/EDcpFsT8DuWdJF5Fctrz5ixn39P24PP+Dia
gPHmAJecZRUJn7sweRWI8T+bSDx9zGCDDRZfDzr5iSYo7zn4BsWkw7xb1Can0IAg
unDXJZ8L1WIbOx1lDOaKtuBcAUrlbwXeI+hqLI4x5nqqa7G4W+bBdBtApNp8bsU1
yYtY7LTKHVsgV9aV2tdE1y1Zrm5tCQ1cB/BAeqzLxuT5eTxlzNYMrmPHXolNuXeo
TXzghevIRaSp+peFc5BJZgfVp4dl1NeYXyHN3eTPnFzFTfi+mx0PdDRwwO+pUgQq
O2sHa/lefmSh3y/L7NreaEdhbrUOtv+EYWCBiFW5NUSFcH36iAehY48P7EmhB8fZ
wHw2cMz/vy8IHgQ7khk8QNBrEDbPGWsu+805dirAaubHEIKe0XCmS4v3AS6ZLS3X
4nq+4GcJ5xNpO/1tgsUmt9RuizRZpKE5mqAU0/MtIyl8Z4/NqERgQcnUllOi7C64
2c0XdYae7D+ZZEq3d7FYZh17zF4JazSazPOLezaL50RdDSRL7pFwZFTXzDCj6G40
oZiPkOEnFR/yD6HM6w+5vExEv4pxgyFgNIG9PoN/ZJu3UAQpzWXb5AcdKAeKguxE
e+h7jc3lrk8HmAOZifaFU+Bn0M+frnBq7ra4Pek5LNT2dUAiKu3tbAs4lykKobLF
l1WyYDX03SnYkscsoZwRyqxn+4g7SldH9Y2Nzlb4KkVkMnwN2v/HJuYCskKIrFnO
tvAi5+Q9l8Fo4+sRsZ2wlUhTmwK68op5PaSc1THdNvVjoayr+ZixKmk8sjr1xK7T
mRMo0zLCXOAHEo7/Rgxfab7nWyICuFRpBQeYNmI4AfXc06leEVa1uZbhAA56klhr
O66MK1O4tsXOhtDChMhOwbpbrvEDL12r0I/gQqPijadV46yJGOCDo7HGeJ3Lyl8K
oKn/mNgFt/An4K6wkOsAQxLaIwat62h/NtzHKcrmlcYUgnAkb2bxlAqUoNNSh2uZ
sc+pPPmKF8EBLjXmnGNdRAsexvZ2WboG/6BtG18OKZxQqtvHN18gF5oq8SW/1Bcn
pFZYB7XZt24bWmd1wgri2c+W8rxCIlRywgeQsN6MUxqi7CSnr3Yg1vmU7DVd77aX
yOM9uX0aNX16n7eaCvElvaciX215ekX/yGn2khS23msHqo6biwiIqRmKKCI+ScgE
xiEm/V8WVjCa4vAEYjDDwNEp4TL8xfIZvDJFqbbco3Z6HqBqTT+csuTkqLgKGUUA
daazRxADMhAacmnVv11sV3z5kwjaCARUOaFq1EniZwrgSp4cDndvScvShVWaOzYA
KLvIaLIyFbdx0394KrPFDu69S7kvS4880eEZdHb9uO5HH3j51quCnMEA6WPS/o7c
7Uoyjc7zO0CcptdxcHoCB/c+nvNcBqZNj+84rVHwoKZisunTnx+UdynzHPPobRba
j+7b+FcU3i4fhzJz0SVg4Nl2E2yhhTqDqUFWBzOkgRNeqYNtvn5CSusxIL7nBjZD
+Q2Kc1TspgvCfLK8VzfkW5bkOb01ZZ9gjeXe9CIhmMPMYzO2Nx99kRak9Ujsj9Gx
6LRZNbz4DUh844bJzcV1F/JHLJ+jFEmDgIW6i5m6jXSeeELU8ABn6JxCu1Zgo2jf
nSwZHkMKjRjb96Uq8iftDbok2Fxn2Y3S2Pe2N//GsA20p2/34cgiU2bT/oySAJ/G
08FQagSsQp5CE6Cc9U7aedqMOlu0trdu2CXt3mKdv/a+HdOVBMBG8lQglBYgDGH3
siMn4KVSNX2cB/+pYKCph1pMlsgG8gkvjAJgyWuozJtWV4+/Di5VpOqnU/K7PLSO
rFp6Tfy7KaT0moUee3PjMImsYM02IwEu2OoNOqxmUmd3VTaO4MAI7xLRAC2P9K6N
8iGX37aYaMNSg7xg7coFCx35ZTopTpVywBzDvyRWh6XSbT4fax4Q2Fi36iMOnSbC
zHWBeBITUEgsZ06oPVNm7BiiY+myF5XgyIgYZCkFao/ne9Ce05pvxXjqYT/Z+Thh
TGMms14nSMUGRV+7dE9otc88JqS9TAfoV5bEYms0hNv4YSAFNhLkMarEDUPCkkfc
/si4L+meva4xefFcPv/K+Obbe2DrOfzw+9slHnSOUonL2/i9r8QiiFnkCXb8eT9O
AUFo/0FeQDbUdbVMB7LQEBwEFksRQm9xdPBwsqg86/sqNugO8j4Pm6JFpk6wChXV
eZrNznn7+6Id+vYqzc86BaJbPzAAvqyAqwGnWKgAAk90NGMrnoo5R72iXp0d4i9V
bMjG4KI9JCEwfdEyT0Iy1nUeNt+ty3YjsZeFi7LO1c/YuwtS9y2Eivo8E2utn2GQ
5Ii1B0XqHfjUA1wiU7nV1COFzPulqH0AvbNMev8HhKoW37CCn9fPWZRQ7/Y/tSWY
CRkJ7H3cKPFF4Mh2Tjpd3gHkXP7XHn5cPqQGK3wuX7KSDOHTtwdnltdoPhY3huV+
b8fCQl9y82QLKsVpsIh8Hj9FT1MGz/OT+7avPS03SEHaOCE9ld1duVLSsJtNxNd+
rAqGO0CoDgQLkQjGdNRRUWYUONHSiTS0ko7GK5RsTpRIB0c0nupvJXtF8lYR0wXK
STCA4FuUR7RTC70pVel3nEMjDZwycHQ9jWGX7Qc/kqFUnUvx6HEIGwqG7lxdPmuk
7dU5XFWiun5sTGEak9IiT0bNI9UUtDr2DPQO3D0aMwcqlludurwpO98fnh/CMoja
q0OmqMP+RdpoCZ/5KjtlVW3vMQrK+Lk8Jhi8f5v9vYdQiyKx2mFNAiFD54b13DRZ
21T7G7KSQ9Cr/GvwKdcFFLdx3TN7vPjd35ZmEA1VC9BGAd5PxRslwJ/uw2nRmTgL
RF/MHsRRdjxFNVfOo3LyaDCRGpOwXiCsT9jSUqN58altSZC7t9nOHIhbds4REQHI
uK9W/2uMJ3ZP3y/z2imxp/LzVaMNM4dDSOW+uXxRsx5VIwHGKCC6U4dOlukeWUXJ
1xs5UqCHUu+6o1PUmym3KrviPsn47z8L8I5xzjZKfdlGPucuBnY5cYC+HtISy5CN
WKxY+gQRjS7vwfuP/1WagBI959GCPExT7Q/Y17aghwElpMugsCSIEJA9C0DfcBi2
avVYpeg81ww3ll0sw1nvhZ1UjgwLVsttcwqaO5M+TnYNWxSg4c2+BAJa4AwNlUNW
aNd1tMscoppVFKvXdC3/5l1RW//Ivoi6nHr/1TZuRnv08iaHnrWXmH422TY0l9r0
aSm7q+DZeWzDKZbPVDPVmKtu1+JVY563fgEX3N9B6B3VgKrk+j+qXaWq+jI1HCX8
30Pp/MMs8cc0so9VV6r3YqgqiIDzTiO7K4LnrNlx3DuLZZaPc5ukwFb2L7dWb5P4
X3K7XShhI6131LuviTeC6LXJDL5jKJpNltsn53aVkuiZQBCUAYq4yZW6sdXKGfiF
rcqj2IJwMs2vmmTm3svilL3XdJd+6Ukr3l6HIqvF2FLGSR2zJXRL0N3jFqmdbIL7
fS1GqLrdioq/czHPsaR38Ancyw5gPLrgkLNdvAsi8vDww8SDCjRQbFlZDagLE1Rj
g6PkKNv/hsfsvoZJb66i3rkCyhgh6Z238SPhsiqhGmnfMBlm8Wc8P7TYfc6wziQT
8YSIlsWjNlNf0E4q01x5FSZxCNVwqldO0avh4Es38ouHAmzEPTGmznlCEttGfTY0
vqdx5rUrMS2H8SZWoIqxOUMpftYun5kkiruCBRs3Mo7YR90gpi+HahsFwYmHstzo
pR40mAasNGbGe+yrCuboI8TaZ9jaUGG76WsFE8ufwpI+lV1IhbOvFerT/pBcPuO6
PnMsLCWWoHk53ZrF8erqR/QGBDFoFx1FcSa7FGKok1biMnh4gvBsNiHpCcgK7/My
0g5P26qIqjYZqNHwIoQpTgo34hI7X2df+CO4S73iH5r0/Mqc9LBfnAr6y5oC5GkE
8NcclUYYMF+2u1+zKmqVK+u9xhDCxinoQxDAGCSE+W8kbjzWDF/pfIqa2DC3GTF2
QKYvdHAgoVlIJj+2qLV1Vy1TlKa+tudQTEjk401GLnGaRdLepAZ39t1o4ZOhEs0D
PVqgeoxZJagQ+fpAgKxgLUYB2cGGMz66DJQadPz3kB5sEb+SCrirHvwiheiw0L9P
MIYDdY3IX8kws2/M96LhU4xI1+GxAaQBADeduYIyZD8CDmPIxWJwFvrgawAfFRTc
N11ARNfB23Z24WgoigwxFQfu5TLNPZ8Sf1vxGTQoBh7VTzEKbVsOVbIY/BYgK6LX
xhnu/F3iABUkWF81WeWys1fgGiVM15U/xh0arkD1lyiuk7PUfHNEEBXEpjIRyPAQ
qWul+rkD/vpm8GOjDZ+oFSr37E3bDZ9JzGh0ygjqs1RrgKa6e4e54XbKIzwz6meu
8SXf9J2shxgWr5TPW+EmUq913ympY8Cw7YBDXUThnAsDNuU2/kiTBWws/xltq49R
AEbQmBanyheAMsX5s++g9tu7zr5wWq7mXQiDV+VOuxvV06ajDhLyP3WSUamEdop4
kqrfyXPhB5kmdGKj4NPSa9vgY0mmWeaSLvx+VhvdOsWz0wPScG6fdCaaR7LQTYrB
PYuCdpUsYu4txln6wHy7N2/TH3ur7nGTrDNP6wx570EUb1gwje6BAXhjXvgGih1W
jYa1SquwHhz7I6ncZNShkDFOawIjnYPf7MJhAYjh9wFkUvO9yPI3E4Ke2qV/QunO
gGr17yX+dsYCgnuaGPKRaIi+7zmEpcT+CmJK/YC6biRLQTHDXpXirriDH1PIo57N
qNSv8cplbys+RlLDgh/VO+5Cq7twmuvUbNpq236yAIdveVFqsAoWJcXmGuDjAqOj
veZSsxoNQzk+IX9YHtY+kNKrbAVi/MZ5ahsS2k2e59JaGjbEM1CeidhSh3G4fryP
akJcZ6QDYvRQDBAe3OrLI/IcmnFjps8XMGgPvec+glbjebmZFzDzXPN3fMwVhOGd
iUstnjvExwy2eJgL9pPiKHioOiMRmIc5RbCRo4w36+baKo5jRHJGDDKAgme1/BDZ
2uXt+MuYaegYdrdMDJ75ZakhHlbR/xanzOP3if8jhHwLdxBwP5wvI2tQRlfH8U0p
Q5XZaTS9RyYuj83bGsLACT+KQ6JbIo6MP1R6JvTRJhj09owXiScv9v8ljm7fSmmO
vKYlcLnBtkcrhNf2mrp0NP2nmGoQC61JgY/svkbFBAOe+rR/siK7hYIBfGUdx7Oj
Ke55KbXmfUT+uGsmRML0XnTX4COcMl0Mk2WJHvz1liUEDPNiR6wdt2L4OvJ8ki6Q
bJzzfdwFc3JFA1iD/I0xJO6yF1CzGNW/qlaa3FaRzM+xDBNRNBohR7oiVWWx/SCU
AGj9OTNZMJwOY5sdh8+Mzu0KFAMmPkzQuVJGr+p2d5p9uArtAXJTQB8roNpVpONw
djKuQkBIpH6K5Km8b4VtGoMQ2St1opzHxHdjGGU7rzXoFza49xq/g0Ag/MFX5n1G
LTdgeiCuEhEdhh103Kr7iNRqHh/kY3No7Ji/ENR3NhRreYPIxVqgGZi/r5rCbqMx
yUt5FJEdCAEX8PTQBqT+XowF2U6dHnWVaDO2yyKTbYaxEcElNWAhBo8oY0+mxq05
VAiERqySe1cpoBZE82Oh3pfvlG2Bud7nJxODbkHb38F57VH6W9GWtGZG40UVJWZT
avGVa31ztQIn8Y9G4Kv7Q6AsAR5eiW0efTtQd0cwN7q6COypBHiD5LRm2cYIwBb2
w0pnOpyi1SgLIE3vu5P1+XJicf9VPlNk30urnKJbj+9N2ZGKKPhmym4uHlPHdoIV
9/Fox6sW4OJX9eGtCWyqBFfbvVU0IZ/sIudZ2/Na1hAz6k0hnedz+m8iWYctWv10
MTzgXB2d75sT7FQNADsPSpUmoHTW+bHkxi8i/f05YldjPNcb1mRvS+Oaq1Lvt5jx
IpX+O7DqL8ThHKzhv8OYDm1iML2mA98fihyeN6R7G8Au/nOmjLpOADf1LjttK7Wc
O1H3SSbTwOMysNnZFzj1BaeSoew6DbAdOG4NOgxHhrW1d0UwTPVS2MpNrFuqGn1r
zooQuSkmFK4Qwwby4zVPPiyxdZihgMD8spKUgfuKsnZQOhfhhWgnT8afPB5t1SA+
7RlmUMBm+Bs0qFHEle4D9nWwSk2XtRxTQg8jHx5ZI7lBBPxWYHKmSePI/HyPultg
uXNv685HL1TZdllKgql1pJQ1xYFY1GdlwPfKamCL8t/2/2SG7RUm3BIFLOynBdVC
Y8ydD/yHcWSAqC/tQuugxuUjc9z5A+th4APfj4wYa2n7HAKwtjh3J2Y52saAu+CC
a+4yMtjAjdD+eUh5/GgKLeduyXc6mENF3JGtlWgTovgJy6in9VGgU9Jh3nqio5df
HhvDUUkhzXIySZcpkSIoW3X6b+47uJxpkddwy/djRV9DmkbIMBObWN8u6vkC/E/9
X47qEMFwVzcmIcM5nxEi/InmV24R++fzetr5q8enLmswTjqfMT8zkY0jdpDnpR6z
viotmr5kDZNYb6KjGWqpNV1sybd7XQpKDSjnjGS/psQgCHQRW7cL+qfD2F2MyVOh
iPSxEF7rFnMuz2CyuAGVen4AZ46U270up5WilKGTskz6Pn4p6ki++hoEeZTyDEt6
3H02QsLz/qwfpeDKHQgWMz/MYs9t5fJobuQk3nocB2Yqe3IjjMCgd6eE23oWylea
c4U3kKeLkkzRv5oY/Hj2cZLMdQrhT6JUM3YLm8dy6kRIvd5htOiS6+n5Kh8ST+cX
BLcNdC6ETQAiJiSX9zewgQRjJs04MW8ncrOnuliVUPCZPeqS81jNz4LQPP9otaWq
F7LWb4ewHadoXRVQowFrXqbnLGX0f7JUUr9VhS+f6VWVNcJkwo1FjkVVjiNJJr9P
ctc7MwzBk/4Xq/8K0oIktskKrhBUfRJwG8jW2AM19QZ0JkxxDEzp2Ij6aeXaUFXw
sEa2i0DFwXWGNBk6bpaTbyAhLBUgsnVEBgYc7gJDYwW0diMULrPsFj0f8fl4L+wV
wBtxMYgVGD7TUOxIKdlHXkvMWzq5VtoKGOpIHXYWmoAq6F22aiE/oEvdtsgVHQr5
AnPeGvv3PFPQlnOO+/QufudcgtE5mdIoWqKRHv88h2hECvJp4fZcUfiRVzqntffd
PfPuqzr5o3Q2xIzpDYnaZFw0sJf/JkBGiMr4N9HoANfWRjrSGf5g5o4zn5ajteHx
4XTEb+2ZAVfp7O+Ojx4ih5l0q7gy8e4q1koAXXKrGY3pC4mZSU9I78vDQBKkHncH
Hv5k90PPGIArMWFAtty7bsmDC1j50m+qw/7AWdKWwsGX9PmHktlg7ynCbSSvOPt7
n/kWiQXwpaMRoSYmHriOo4h/pjbB645aa6uYFfr9b4kUE1LWUL7qDHLLKnlEBgcM
xpKZNZEaEkaDudEpYh1YLr/usQ5lbDC4TeDewYPyN+2AhOeIai0Of6MeNlMACWLF
IRGVYtsle1YLQUNRfegfKjSyiyvK40lp7BQDtQp6K8dkCLAC56fv/a26VoMWgrjy
4BPyB6MuCdWxcaI0w4Ztp+48m7jVc/nOWCp3v6jLrwAGrZqzVfZDV53QzORZ/wfT
ePfwdJI5w3luUphC5REmq2p2rvR+0z9w9LetA9VMfNTBgZXq6GyRzCuNjNptX1Nc
5TB00MV8CPJ4tkUhKxL7H35xS7STQbErZb4pO1U8vt7w/8euxw/BalBMzO4CzxRy
AEIUKOPoa1/r33utC7iC0aaA0dXAh2AKHeC80zOA+YagW5iLyYGdCTyvY0KJxfp8
pMswUwtuhiqkCMGTCJ2rPNqUjdUw6kM5TjifYbxnPymVIHG43Q17S/IQqNfK6TS2
BhBFpcsbdDGPDS6nfk50Lc41b3gOvxRzdYLSU39Nt2VqqfbfwwXQSMoE/xAOuWku
NBcTHs0W7CTOY5Iav6BSlo9wYmzV1ey7CvmXu8I9g+CZXbk1yCClWo6a8CLN/WiN
1qNJNEJBcY2JtMIt7cHtRacvi9KQAJJ/uOMAGE6fswkk+nbdGMQYd667cBGMjQFX
kXjRRe7Hm1KLFxfPLlXTKfF76HouGT6KEGJgTlKmuxFpY1aD3zSMLVThzCogR52x
0S0PXyLnM7iNECVis/kZpvR+QH6BQFyX34falLGi4zBG09Mhqp3nFcYJSu78PEIs
hV8PgWdoCDYisCG/ALhYwveKHCFumriEW+h/O3IKtTu1xEJ6MU0gDAHYBuuL3oVk
XK8Z2nZc7Wspd9Punf0C6quL5evIt79ZqrYQooSVTRXV1LQo5GhuZLLDdyZrbutw
2zmAkYCNuLRvmjFtzGfVkq0HXFSTRuQpCSaXxq4kjKlH10gZuxUms+sFo8a3ehbR
ePIZpofKFUpm8GdYzZoJpueAu2cGJzqawW4kA3szJ2IptvP8SRWLyv3vRHsFxT7f
vBbnAp+M64MO5Uinhd2jKNKkWJ5ThBdVTUi4exR2idh9J4IaI8bgu25E2xvBId28
BP70iwJtLcKcdsBjyN3L1n8rDZMGIPRHH77spJqxuSgjbiVJuBsFU7pYdhLkcvXx
WfJTM1MgTckis2tPR1YqBF9Je/vqyalXvqiOkha4agM/SmuS8cnhjOLtNWLJJ4va
npUYO9GLgEbUzcLN0vLY660390q6iBCmrXGzwSQyOXqy/8tlXhzPm/XLjd5eZN88
uco0pASrJicL/dBrQoLpdAcmUxV2F17lk6t+0QzrpFrxmdpuv7Q2GF0+YsnJJ/Vy
C6lMV2EXwIKRnHf4uPu9ZQ1yXyO64Pg5hJ5cN2lXnj9uV+a4qSAPt93LXvrNbQMg
SJk+/DGG7F+i81ih77GNBUn7LkWocVxApLzeztOYJF46v4LRQSPNg6vb/XlwsF9X
Mcrp9Rwn14VMav5LSfEQfNhEclTPg7KGpzMPKiCyBcoG5+yxAWsmT2sQHlvQ432B
qBlF4MXfhWeX1RXI1AcftxKXiQL02/SesWKTJA2ey+xPdkLNvh+X5Z0Fu9o71dbQ
Gdx8uD/GjqRK1AYQFV/IxuFbJ0TgF7OV0Xp5NpaUEAGyOSlgDSkqo3S3pYfpnV34
MXmbnd+pD3ryvQ7lqUA5u5EqK3isIPreB574c6Rq9vVRUAG91VUTIiycW2k0Ytg0
qhg9+CX270BUylmsaREXmiNm6n2wf1h8qNJjBEpGy6KnXlKjQWtYeNUysLWwM0kx
+k2XAXHUpL763ZNJ+HtafmtuMeiK6XD2ZSPZ2kryYSJxoMOaDAoBWQzWLhvE8EC8
84wu2D9ysoxnB2hjEwP2rcVWFqRPYsVTtrouWx5RDDnq9K0dPJ1veSJPRdZIBZY7
ve17JioDiz5gzeuf2OH0c8okOsqzpBcxYtRLGGOLneiiM/zS5VuJ8y1dD/oA3YmC
QeMbG2GbHyyTD24UMtNFdfzw37a3EYPN140lmp/a5PDIDgfHLfDmOn7jbA3ynZkF
2yrqMYRibPkR/b4Ju5vYaYMwDs4uWfHmZ5js30tFKfFWO2aKH3XfXLe/+nue3gOX
xRyEV2MZ+D5KyPYFddxMgYki/V+3HDxj9TqgmgsUlIR6k3XsqkReC5OlQB68kGo1
kbvedPLFeE0fDWg1vIkNpHGFRkFSkWd5Y17mYAd9jAVCDi9nVgSEMMwBSvSLaNZl
8JCiEffljqUH+HsfjkDvtXJrdKBU/EZ5DgluDVF5H6NGg81jhShs9PqrrMRPlvdg
YeBcq5AAFnZspqd+XYcfE4SVB7Uaz3tCU+rTWchLnpAc6b/uJT6abkWmhNIW0VHY
SRRL1CfU6+rio6WzRKtwnVURiot4bbq3/yvVrzbzZ7etj2dNV6Gt+Ol9Nrh3+gv/
T9ecmu8aro03ggK2Bie9plQjN6S4Z5HP6F7OsGJuC8oCuVKGPtZF5ed6oH2gYqaG
+JA2M1xvyN4Pc3znXy5uRaJL9S79jQXlcrNvxTPsBDLLoXInOQ5kwMCV4NYtm2HM
YxJdqcJkY2j+awrvwoN8CE/32a7yq3l7eJ+XM4xvwL3bYPd6yYPjf59BCiWxwoNC
wxn2k07vhRbzgaho0pLiFa0kki/qkgzXpVsOFG+GO+/EeW5ezPn1ldEpdFclwiSp
JJnxZCSz3HWWmp3AX1YDO57Gi/1p1oo0irqxfeLgGTy9IOmi5VpdDRP6PACrwyCM
F2TFyNy0VzyPa6m6BLeIfekgc7/m2U/WG6IblJqIU6TyzYNDrr8aIkaW8X5jobDv
/3Lr/jgoRYDcKDqKBePH1Xvq/aKcPjygOnp8oiI7E+uLfqsbkDNrHXvTOzA7mnoN
o9+RJCweNZiwZvVweCyyNirhJlZ88SjBTccuphzRvI+RRZVwpPVkkrAT0STs9DVU
BIHNK9asGzLoB8i7d0JB+OatsS6i0xnNeE4uhSv1zISQRPOSfgAn7g8Y/2bH+3Bi
iOvy5yYpgk+kIkrS0ug39+m/e0et05yGq2fP3Hg1UMRZcWe5Xl6rI2b4PZVV9NQz
hQ0qoA/RCP1RDZ1gCNGytTYY7Wyku3fWiF39V3U6czVML/h0I+QqmGhhTACRCI9l
rPj2GDsNIyW4uK2R0GzLTGPUenJ8iSf+X5OF84buYOSsj+nXIW6niUdMiOh8yJu+
WA5U+ENfiY15dHBK4P7JxDNghPkYpMEEAGyc/yeYKeIwBqy/xZT+n+ngGzjEBvnV
OqbGHuJyXEKYQgZX49tokBgDe/iAAvhzjbjIxUC412QoUHHJVW2DMvNecfu+UA8V
aDDMIIKCbgbKnGg2XQFKa58gV2M+tQo90/XbB1lbL+AgMPvXVym5xVHS6dt/zOiF
SXt0E1gaCR14SEV+ss1SWsxDcNl5gtUiYF+Eg53ljJU1gf1jdwmRf+/iT9dQfhTI
aPwiJ45LpMISEoTagGUwB7KG2TEsdyDf9Zp2lA5NgQre9uFQLiK/36cNwz1CzWMr
n6BxlkYGdC87qvrMlFrGZxauyJsHvClPzJb4Y+PhUYt1zB2mUvXiq1DmU9CykhbV
Lv6PQjmnHHQypUQs1kD9cKHXjVt2u6K9Mw1ZNimIWlK0BC5epiQnjhkAc1+016iT
0eqpagzs62x/+atbjkLYSI1zjMyuWt6FHxwVWvofRVLN6CKsB4NGGGl2/8zkqHjv
/VVX3aZqHl65B8u7lTAZw12VhI92BFNDQ3gb1528B0qxJcv5ZB1MbhyNhF1rLiTi
Ry5jZwI2ZDcxxwSVuAxg3Djrfyq2y/3PdxhWjGnPeaNJcrn0gmJEkLyRBbs/5NCG
bJ6NhWai8oK2vQBh012q0oHwcz07kHEc2hiDIgrfExEOnglzN9oFB5EL6JsQpnHq
a6+Bp9tKSn6dmk6fQ3LsT+2VO92WjztQ8B/qffug6J64Nvb5bIKjK4c+OmEXc8rh
LjVjNpX3uDqMBNQunDy6TApM92LYFKIeLY+2siyN+TuZXHuw3DkbxUVIdPZCiNwf
Xh00BObaDL8hIYKT4qzqbyeAdIhVI29YiYhY14wlvSw/s+D2jNO0Oa8HSIGdLX7X
g1v6HLgmcEZDoVi8Ye9gFz84PPCmRCKT7manHglIGwwa6yHyDVhj5bGahy/Vv9l4
2Xe+j/hMOD93QHccO98W39kvlezkHngEf5+OXNOMCkk5vTRgJCHF/BfnBOUQqmSu
MzvPMDsJel5qlLnDSmRX3fWiByqJ4Vqk5tudWAeTt/wk/8ItwTkg5pz1zPUbVBeN
o/UvY0NfkiHFNyKXH6/iTp5dHX3IZruMzcZfGdASQyw0K6rhiZFO7iqXlM4ZTIU4
f/lAQGSNObziqHDSyHdhaLKZmHoXw8oEF+37kX6VR/ZL88k4P+d2JiGRdiHtRfx9
gJK8mWILAn1qGy4Tu9UAC/6GsUDnm983aelRBxTnZIn8zcrT1XoLSQ0mSWRYMl0a
9YAice+Tof/4qh5uegcPnWR5QlCjh8wUbkcnxx/uG2a1aamDcQpqSbSMldOQgLmV
bIkm7npM9bGg828wb58lsFqZBvf2b+6Zuk8lisjGWGuuDx/OGsHT4Ui6QyDQgWbE
d41AU4N5vM+p0KiNC7rk7omoWD9hIopHpfDU6FU+rSxH0jTSeh1jAbvJSnBmmjBA
3qBiQ3HfodEKxneKJujBut/c8zG/evamXw+M26ayKRt/3kJ5vOm/+mtCw1LPyogN
8H7yZSwgfE7Tb/788joYbJrFyMM8BDpcj6DynKy+i6Jt2zCHuA3hZxcUsbJFG/ta
B4p2Gad/uhOR6vb/K8l48r3SIiBbX2W6xvd5zZEcMAJxcDb/RwUFn8EssHS6Wil+
69hJFQyHYuaKVhQMrD4lT0fg/pS4BRjtJb7zAM9Ia91CtHCO5Tzi5KAurMov/oCJ
ogMZz9pqdeX80DTrFTSd5YWPIjAUTGimPrm52WIGVGPBV9YHJ6E6ckLebR46pzkC
2ZwDrRea1TaF0y8eOl8HCYIEyMu6Xlg6Xdmi/mcyQq+o5ZXxR4R6aGKugm0uP7gG
82Yc+1nKj8LfHXT+gjIYkLXiLU1F2SvCyukmm1e6q4eOWT2CNQ7tHlK01DzrXHu4
3n/H9uJBWOri+ljZc/NoS/uekU8HOqwr6ENtKYagilmAuGPqzu1ETDfRqOB/WJfB
ys0wb8ZjzgNth9/Yklb49nCeKk1WGFG64aP/dcQUHivyG6MGGljUkr/z/Pyw2RuC
FykmJ2iPjXJMx1NajzkTlugoqXyHTDHGz64+Y9B5/L5P3FgjvPhHLt54dT0mhy8b
wlzhhY35L2YIC4WzO894tS32BXSAj5Lx/RCVE8yweNTI0Y2mDMkrONtwF5Eu2d8n
wfb+StPdLV84BC+DSLoEtPVXxdDtdLOdZku1RyJ7BAvZsquylzBEEHIyFQTDtDwB
HGGhhWhJ/MAhdncbsGAeHd8BGZ3mRCyLN6unBmAGY3D+gZmV0uUanDY+Hi0TqooE
FkrK+bJAYreaf6PxRHOg6yvprH/lji6E6x+1TeG//+oPOI04fMJM2qYC05Jhkjip
53esvp2kII0mi427vOrbKa2NXOQwzqtq1Nu2b3g8XC4N9as0iwC8s26gHmPc9Bko
aYcFqAbbC+m5kSzgVlnctxZM/7dt+HYnagNHGjNAu2oSSIQ+MTR+VrPXMxro3K0I
zv1xuQyFhqYEJuuimeH+mHUWQt8Z6k7xD5IJ82rkPVjp2kEHrCel9O/lkt+6wNHN
+Ra34X1BoChm9N53bfo/c1IwIiuDfSR+OOjkUXwa8tHEoWEdxw3ti6M3CwO14ZxL
aZtOCrQgpzcZTK+w4lUn23FWYnRJ9bUPrabKoSXyW6aB8o/3iboK8NSFjc0uhKlx
fuzzzUjE3WtJbc+ejLTx5xWsBqE4YG3khmAo8UtMj2z+pBV+QT4n8mCHUaa9+7uv
M3uOZiLUtOcBexb5bE1R8/+okeL/EfAAIBdwcRUeL9RCfLshifADenHnXSK3P34N
qYz4odRTj7zHJeWhkjIVUb1Tfb74DYnwXsSQQCN7NTnjpia1/JB4h/RK0X8Aesku
NTx29TOinWXFGV+4KzT/15A7SfcfZbuREWDjyggbQWjplu3Fw4tcB9P6lWTy/6k1
A0nPNUv16CmS0NHdJb7dJ7/L35ZvZG19EWtLqNbYwzijwwXEdKXNz+vgfsRwykVu
MVmq1LZJhaLq5RES45wIUTFa/+pyzt+Jt+btQfTMGQVX8V/2qxC5H/QzHCAjFy4p
qVx+56mR09vjzeqgh3pU9hG2ZzmM0KDoUrl4ehzpDHYzMLSRjoz6fowJFc7YL7D3
bFXsE0dGUqqhJWrnfTalptdyD3Oqo3xEOJtyVdXpkdd1BLZJskk/dIDpZmNety/5
DqHOcypR5xHSP/b3IaCnXnBrRMJtV5tBr2pIy92qPpxRPpEVZcYJrOr4G66MkBMt
5e2OOCd3a2ZJkObmKCwLT6qRRmschfdvrFTcNE2/mrNZaA8il+G4FiYLs1o+ymg+
QUdmcWHQ/k5DrX610PFUWCcyvuQrbO5syCzyN7G709BshXN/RlnuCTEjhmd7Ws8U
HKVC1W1Au3jyp9p7pbpv207PtXc/iQ03/5gl/YqqFmo0ORzpfuqfqL4FrkZP6hrr
LqzAUAcVgBNO+m5zLM10Z/4HnWPBibDR3nJzXdkuy29q2U/wgoK8NIeDCJUGDNzb
LYKxujcfMhzNKvSfn8ahYOCnfLogSRXX0QnGNnKImRDkpR9z2J12w6IU6u7/ZsBM
KhSmtuQWHp8PYDv9LTqO8L/KBqLr+LVuRMlffi0davAgf9hh8X0G2YPRyYSOb18y
3QbyswWd05zwSmlZuPHIaYg5TWXLQ+BOMC8PgEYBkq+RiwsAqPD75tM3Kmp5CqFs
OBREULZVeoXpNrMn18ynk+c9m4VSmg6e54SqxEIzH3RoY1cJMGNnp0gRj4ycBKpb
FPX9IUIphRjKU/2u/8bVao1LhKXJtwHb2TWd00yQqcnlj/pvUI+mpRwFedeHodmw
9gyVTk3LbK4CPsgONDy+TwfU2SQOaKR9eUNxAhrRz17Eykg7WEPs2TTIbqs3T61G
wRCLXzJFoc+vdXTm1lqD3AgSXLmUZmJ7+++zYHBfm4og+PVBYM293bHY+3Qj6lxR
OQl/DToYYeWvJIfhclmGFkuFtAIxyDrAGUc+pGjn6FJm5KhNaJTNaQYCH9TSbGnS
eFMtV4SwHsieYu9eoCqd5ypN/udsWzKfKqRk6p3rjYNrNHvKKN2v5NfHIdobg4Ro
21DqbEYMO515V2Pk4hvGBmc5S9OJ321MyMHT+uVQvcfcM8jk1Ytc11L4D9aQ8OZH
MYC2fdFD9tXfpdAgs088GN3YiwF1WZm4C3B9X4XdzMfYhsOl6b1ATEo0uKAVUb3m
ihMExrcmBsCx8BxgeVmGZd32OgJpsEi632Ehs8PoHlc6M/WL51qyO7SyKCgBuLSZ
8/87cQZroZ0/NS1wyM7RPX+S46wDumB5ZAD9/fNmG3jugQLcSDTmYEgRQXoW+q0X
RwVyX/QsnURkjMjbYvP6un9Gn4mbacUFSZWwp42+tPfc2QUQrXFbliB58XDp3aPX
xY2df6Q1iQqfauVxuzV8VSw9AigK4vFjdn9BRuzvE1//XOwMJpY4tyBXk/xkRObm
ZoPhYexWLQwU+MXTqbMHWFTSXEvk2fwaYLebVc0OFagPWQfCHpXBqSO5rpXIuOna
58ifxMSK8j+XD+aRLleAyQOTyZMAgZrc6Uv7RiyIDAlDIJt2G02RxaMUM6mkotSl
Z0L8hn+SHap81AOPskZJqi5RI8wSD7Lzwj3JLSgO+EGRFLIriUhioVqssaxv3s9b
8kTKjO9MbJeR+yKKTHC79EOjX7XNMPIXETfrKsXJtqM8+fTb2m+T/kVO7NLZgS56
eiA0H8Nfm4SsY4IfYUVXj4DTPsfDzOYEHDNTu8bQeaUCY9WKmqezSQ8bGPyUf79a
xBm893m2OZdCKrS078GezhU5Qqpm3hrCYrLX6RM/jCxMr0BtRww1oTRsYwIUZ6Gw
Y5TT0+vG5QHFR6IYcBJkfMwYUa74/Wfk5XHza8gVTNU5ovKyfSjxtPBBNsGgk87B
DJI9WcDoFG3Fp5JzVv02+jbJ2mSKn6EAKkQK5BQ6x4NnuCA0SUb7nRXtGC/6KKp1
876SmVhnP58gaEnKOmrX4dwfIyBsNGmsZCJRxK2W7VwABaRWoTjod/GmhgbL3F9h
id8b4QjgHhRr+zZ0EIfLEuEhWlrxOJpgSL18URk3p4wsJH/JTk1K9CiRUDVBmyE2
dV+tHX5qQqxNxb0dHb8i3XBeGMRWt3hX0yKQxDeuRnhtrcAw6HNaIsT8WeQ/puvW
dLDkmOnppnM/b6v/R2lfeLcn2ilTBzRQLgWiYjR5xj36gMOibWR+IheZvjcoqPhk
SW21MDzbecFXK0S18HAvRrsn8SMifq3lSz6YEsHCvCb9gwjO2lM1WSbBNMhRJvel
25Y0JjslzDuocWjgGP9/eQhZfbGFpvMhFci7sn4ZFT9GKwuMtHFP8cCMH37C5zSb
TRYhy93abUk/walayOwOq/kl9ThTMEnBF2U5F2s4ONtjyaDhF4kn14t40Msw36T+
UyVQIyUXB/lpsGrvKsIZxowObC1dWqY0KzV97UCJ6fqEUlnSUFr/Qy7hPCL7MU4V
JGmFkE3lEljhcNVmxn9BeUSnuoEHsGtDI7Y770ABye2qDxuyTl4nihUI4kXA6v/D
SLOWueDSBSpc2Ki1SC8dkf/U2agyaOAb7F4MYBjclV6LJa1sPAqpyz364jz10DO5
PS5ifeBMehBphPYz0GD/iQzoocKqeSODbn76xqsgwG/2NJ6rHbzX0ukJdUk67G4Z
8kv173ihrYQjI2rOaBWVAfNcbabAWRVU116ekPGX2WyvqCLWYjlumuzleCqdUT4S
FClvoSPOyO7to1su7pzBhd97NucGWzuxf/Dfp6E/rQahH8OHlJoUv1SgT8enh19D
w75yeJApy/jKpvWmQvJ4lZS+okfk2dsndyY0JcjTjnNH+XN3Fqm9lmYhP+We6Du2
szgAmiEpfEgxfH2svYTl4j6+KRHKkfAiW8jMK5odLEXep7kr61ZQqTohuz4vBTae
NymcA5wsRWjEZiMYwhzDDVdgYPZbpxaRhhzzemu2l3Gij+pfBsSpkpa0t1l2Y+GG
k/OvZfdnkRSbrSNTEMOJDO7c1Q/IoDAJlgwwuga3UDeqWDyUOTgE2BgyZsw482Kv
Hez7+XuBGjFiI4Ikjmfzs04pvGs2beLTXFRxLuCgyuwuMv+JWvTmzaEdQYFUnBZz
XfqGVfx/TJcoah3tQciKo4ktt/7R7pmZgk/rmkX6P94ypvZVqpkC5CZ7Mp8Z0lV/
KH0zICzHbSIVx/CjqYcmT8S3fI1sQPUJeV6gIGfiztOKxB4xELl//w2nqW5IRogM
IxYYcxpkZY3kgW11YxhI+EkorHJQL3W4vDyPq1CK7UvdXXeo4V3P0qqRA62eOi9G
+Ig1T2mlJOHmaVQUIzQyTEgQVdjmzu9LkxOwXSpRzktpkOIr538Dr+b0PJn0VuKU
ektgRGQhI+IcD4w1vl2AIoWmyoTBuu+Vc/AygJawm/oXorRoGpbf99OFe2KAE96D
ZTLN7Or0m8YUPlMpFIrdLkbaOJYxOnZXEcByYGjw4bekdp/25/hDN5gpx6sKlPXv
YjjDvPyO18BqrN0u7Vh9BNEfk0fx3Fq5LCBQ4V0ryS+De12BMnQtDOpXItZW0/Kk
xWixewltUSY8NhNsxR7DqxwMgR1W8pIY8CB8yVB2KuRIijb25sqXtRsnOKzWg0g+
sn1Ld3zUgTqAfO/LrNM/xsR0tWlEJHpJqVqDysO+zm3DWgUMrxS+IDBNJr2U1+Gh
Pfc8jJI9ZSQjihvokpmxt7Ah+TVD6z3tln0vB8or7I6OeViwAZkeYGCuVN87sSSD
Dds4gkofnAGs2CvEJi9SC0UxO8Odq/TCOQSwkpln3YJtAOhOBP8/XAAalSv58hBm
b8XS76bZSRe0/tJ/8EpQe1MaEvMQ+XPdh0T5sjND/D/rabYCIV0RKco/0XSQ+1Ao
MNxh+KmWzKo49jCf9hUALO8Yodu7s4iHOZK+85NWIRY/Ji4+ClHpdw3iwpBTtZsK
W3qRqNuitrmLtKBWePJw/U+dAdjquRCiRW4LLGUbuOQJ+ArARpmvgeOtQQu3TWT+
/N8Bp4asVIAZMCY+XPsm1TlysR0nDf3zH5hmnjZo1ISMJ+4IY58lqUTXtDBL+V3x
te5UZDgZWpE0M8G8EZTX0OF9Tm/vhLn54pdL5tS1E6kYkwu+otHZZcElD5WtJ76Q
vyDsUWR74qF8AFySveb5TPNmXJt0zCpb2ZnTaE2j/Ytc1QmAys64s/AKcst5n48k
hfVx6RoNiaAO1KXtvgyxoJ+P+P2qgzXLMD+9e+8+C19EsZjbAjFTg6QpKs5mNju2
MIrYCW1VOtcPn9gTaqyDangqbd+LteOwcXzyM/5Xo/uCAdSiBkg89OZMpZc9cLBT
ZVco/1J7DeLqlP3Nm2U4m0QYdiu6qW7Ng8jhzKNLD0XPVAl8hc3gGxHxsP8VFhdf
NJIG+0knEiZ0+/EBSQ8lJRvTPhiKC8LzJxVUPoAWmQS1fktOTjr40JCCHkaIZnJH
cxwFWp0W/mJ2ATIuEI73MXEIiXWoXi95aiczy71a54p+2m9imFA6h86KK7jRf8CA
PRWLKIpDPDUjHKuNltz3XRmXCt0A19H3eSUJoXa9uTGiQOopnWgDD1Ajl6dhr3hZ
of+JES+8IEeilhIcSQN5Ri+pUYcEWEXh6Brfo5dQxklOCq070qFzxh25NUgIRhZv
XrnsKH583TO4EPHZEVC1o4Fu/0JL2bq7+5G+eBKRqzYbIu48qFHOtknmdKzx9VmI
5D55yesJIMDcTysJqGNcolRWPUrlMwhv4XplsknhokU1nTPrXXn5MAAtaLrBBVP2
jxauTckvvElSYne+CN0YZxkTbUTtno+Nl6iTCTczRdRvyFXF5gk51tdWxIxxaa2S
T48Z4eHGWmqQcih2h5wmSoiti7kr7/WX1fmKeNq5O+tIN83j5/XPey+x57XSlexw
/5PtWX41Yr8VeSkOh38TuBjAvN1hAd16np8ORxjs+U3MW5cOlHL/arJxh19bxSg4
uBSo2ovetXdbx8/DtAQXMLpqAanuqTBm2DDtJXNr9I+RR44tQO7cQhg3ie+lisQv
iDYuuvt1w6YtYpQR+PyT4UcsXeZnriDEjh/EKVfKNl2oSrKA9aCuu4mIEBG8gdLu
LmIeMYQm6J1lyQih9X23N7FpNtSMGi2amj50cZt0Hz+zDOrkPeOlAjwUjIH7CYF/
RI6955yzJdDcI7i78yH5shkp5gtDp4m7CLSWRRZ4I06oHJhH+nGJlOXML0ScIeCx
vy8Vfnq9n4cCaDaFdnZ5OvwS4mYI71GP5RSRqi0/tZo+09JC5okQXA2YpN0SzEO2
TCjgfMRnfHvk2IAWpI4akw/lReFqHrDRbXbx8wntkquuXdIIzlAB51sUmkGi5OWT
a6YYAs0j83/TqAJqtQU5wUb5ISGlRuFti8vY+fzCHs1EDA5BCs7n/rl1QTR/4aLJ
+SDtpZ/o7vcnCbT6SKaD+3p+HoUaSU8UaVGe0ZptKNkukCwGuYt88CSRbUULAs7c
hCMibdY9tU0YD8umUgdunwC60+df4AfJZfXTJ4b9ihrOE9nPdzBs5YPbtagaoG/n
fHzZPaidr8gKmOP1q0IfkdCXyv0XUsErHAnrC/XLohGx3pAjDbDCkruWjM4UpHjI
P5EZ8kN13x3FjpGZfuoBsCPituJTdlhuUTpzVWb/xtuJ6O21Od9MYBhU9aICrXn3
lkDgUjBYlGmk0JamzbpnhXvZ3yGZTcnE0Nww0k9AwNRlYyodu0rnmc/AJJgc8E64
1xdC88uF5RuBJzhpvEww9r3KymzwUvvLs+futzEdO6sh2kJMZ6lvAj0hXfmG/DOr
hT/tUBV3HY1nG27BATUlz5zUxMyntCtX5HQ7HT2q2ne+f26itNYB4m0P3Fhd36JY
iLPPxXyhc5ihP08QOt37pMDdSC+X1kz8VwVLpsrGxgeCL+Klq+K+GHZk4qFomdSS
nZDQBypuupcBwFERVPfVLDlVnHhSZ2bQKAe0LKMmLPdlXBigrlN4z5KxL2Jxrwti
cPnlGT7MHOqmAyGbJ0h3yJiw4WLJeTaijBWdnU1Rc0Bt56Bp0OKGBvfG201ReoMg
F3G61uKd/J9xozu1LF9DTtwsQ8Wwljpl8nweW0m428kNJI08b4wF5iHL0sBYXY92
5jDJoEFYbTs8wZM11HwStLPMhX8eEDmanPMiQPOSdiv1laaxVHWf8XfZ0BEdCOye
pVswL0WqWsYoe8QP4dBoY6Jtcs5t7OB6Ver7roJfDJOjlBHZdSx73vgX8JPfT6P5
uk0b/Ca6gC+MUDIaFWz5j3mOe9/khOSeshtqwqlBLanusRORuV0fpNOZ3qiVX+2o
RMHM1auTVND1tsowJBrfXeolYLaQikOepCN+kx/Fv/idwMLRUx0WPXBC0FXcBJYQ
OQlO76r0MBJA3WKybAfaQVg6scwmMmfEj1Oh9Wnq6bWI7Mt86lF9RJA8aOOHA8r7
M7nGOUiG3mcmQhbN7YQKTw+JUcmUkZIJhFlVFOGeFCiHrSe1Fd8mCAmhKCAa9waf
efQXPHA73SbPAvaKeyES2AbG/aJXWyc34HdwHWFmPBP5IrjvvV+H4FHbvbv5GLrA
J5Bj1EKqMxTT2lnsLZEFQnnptFiWpjVS5bvJ+PUoTbO1sOpOTczbigjGRkOe2bbD
VXm7CqKPziF17n2ZQNyJ6Gf879dGOyCBHByul3LOx7b1ZcHK/rloeWH167gXtQQ9
bXYK+W3GAraK4ue6f9QScn7DOt+M2vOpZ17K4KFRbjrIhkcNRGT6N3v8cX2ld/w4
JKowmgdjkIbnjxDfnHTwJpGSH8seP2RJkS1dsTbVe6TIAfpQqfWRsMfvTAcAvJhh
eA2AKwHwLPgvG0ElIcmMPUEtWwjwOZx0lzPkGtoLbuo7F2gveMgGoJinOG1NX53V
oNFSHiSQzI8y6Hd7wA2JglNHcHPk6U4tr+MehGGq2zqEQp+ky3P+G8TpuYAsJCKw
qy/U9SIbW3G1spRELEdlDdMzbByL6Gi9+JZI5BIC4LToanvmNVS/XKejqB+H85EL
AXTUc5Xy+29eCsoXoAprhU1guLmE929+GLUE5fFL2i2SZTzEQKVANjJWpjOpcSBm
6RoYZmQKTNLtC71din+HMUrv2XO5JUHA+lG9ZhLbNNytNR0/5MzJk13ESySzu54g
DGBs2VoG61WB/XXm1B/AHGs1TRrUk4KLtG6okage25NSZQyFk4wi6QMmwTht7sxs
1yKOUBNNIZ6d5nCQ7PNiM1BEdmtKc36VCcGi0F+xAJnrVk32XAGiSuTfHJJRv4a0
XeUoE+R4wU5DbU/+RgoAqsW/El/mpZ2NwDKWCk4w4yCHD+1A6ZXN4PubZVij5KOD
orlxIwaLg1REC3P2MeZoGtGQoQpWz0KA7j30cjBvXr2DW8YcuqrwrQuPQqhg1KNK
nBsExaKHfyv/pLwG9HfSlAZltDMGki1ZW+1qQL62ukM5qlL93BEx/HRdKBeCzZOl
CB0aYXU295HkGL7vYbTsFC84/bio4vryaeByGYmN5UqcSkrerqPcQBpKtBNg7PH8
szIJk/D/+++tPFO3GN044hpybtLEYh88q0gH2qR2s7d5uzLJ8dCLx2thLAD7zX9V
ajLdag2wnkU3mdjuYaNUr04cvAAgqqR/AB22z1rekgVFY6DFCOzGNgsejA/Oqh+F
S/u7m+94ZfImS7Y9uOZ2waWKnJs0D7jZouq8E0Peqk6C2qL7wloIBH4gcqN4n15S
ix0hkNjlnPOlSpLn2R3t9fDXVJRRJHP9y9BDQm7FJ6fVTGPpu/ewdOlhYGS13J1g
TJkL0WoL8In3RQV1mkD/HOTPgtiHE/Uzq0Vw9aHa6bCqdUq5mb7vIKXz6U36UnjU
U/JSosxCQegXC/LunfNmnhzQozA9M8oh05vBNLBL+P9JAw05XjpCQ4FZ6OmAW+uj
71dRhcvyR/adMXZUY8cRaLaP/f1qpFAotEHTK7NZPL5+RTShtWyCj/SjmB+foRZn
XA/yfHcNXwuouOpeOnvYu/Dl1ZRl8R1bUzCp1TqK10P/Wa5vt0ZEmCGpEeiEbuS1
BXfV/MXEIdKw+TZWbXSmzjtapq9SiFtq7bQbjTTxQANAANue8Fd3MHZHz53yOHU9
jMAxIlLlrn8auIqNxDcM3ZlrfI3KPkAtdTkgToAEoH2xD4xSGxxDbE8LRQz9LIA3
bsPCgh1pzgv4BRSosIz6yosAGCe/4sECaMzMNpf21G7lrcAlc4fI6ar3J1QCh6YC
H12xX7sEdHGbIpxvlcFGW2XMNe4x8NQJl3Px1DnvUUGaIPhJBXMpeqVGIf2bL3K3
OZ8McZrPA2KBchEet0b1hwwD+MthHQkdqzXGn893IDemfImmtrIvjYzjoVSGMNOJ
Uk16ncjbbnYk8YVxZAyxorIoCPQ1bOr94Wps0nTIBUpkruAzIdskmbUpY057Obio
FFtKzJepnZNlub9L+SWPw8u4WZGnDQLtdBXMtFPMUg59jPBzijRviWKSE5tO5Ngd
rdIRDpO37Js4J9ac05q/zEOaJS51yMfxTMzgGMGDTBCPwzilKMfpMLE0P94107C1
/P1MyHc4/wbsVz/kxDIK1dULLzpcaZWVVjV5vKVIPo0PpbLIrgscf/YtFUiqKL2r
0c/O9G3t8KjqwHSjZhImUQFl9t3H/S7fKi8Ycz9V6L8HoOjARYJEeBypcS9n10Ze
7I0qy/TBkFSBBN69G2rvOz2WhVrWtvlwqAgEs2r1PSF3GXkS/Lr5TLmf6klEiojl
Is6HBiDaWR/5Px7B9Zquu50WfmK64XQJhkvukCbqQHBBaCkBlxHYypONQOQr8THo
9f+JTqyE+YuXTsSPNCRxnIwlzj7RCKPNvZwKsUV8AzoL3/uPUl0V9Y4p3TPE/5nb
AKs/YJPROKE6JTkrrHFm0A2zwOG1C1f7jtcwIuhC0HbpGREPI2OVW6tslgih+/zL
WsoHvsQ3YY5tV5OY+6UlhiT4CQt/lsb0XDMRhr+ububHMwDLZVDoBvrMzMbcQ/h7
T1y5Y7FtL/dlloJFjF42K88Pb3NwkHkB8vcDBJuYflfRzW+28Mf1Z1v8Ij5z/uiw
J/uu3pH8Lvd3zRc3HYtRyTWf7wFgKrXdPiCyyUiCBgE5gFJFHoz4XMsY/XVkDvps
c304tFh4drVD1c10DvRSYeu9BnzrMsO5I7gi8/HScbJeXjmrOkip6ZC9zVdtbidV
MxeYeejGOxmJuID6P6xdyi/PxASVlLzeQB7D9zqJ7mrXdAZ/sFjWjY3XLNd5xwFe
nud8FBirAitzpK+00gOF+z2FnHw6V5wBB5LXZP0XRqU1IWaJhzHmh0RlL9f64Qtg
5CbQX2qutv5Xx+brHfzH0VC9BmrDV78MIdsvseaWiMKHZf6tab3SF9cm/keKvrQP
Gty4SKHIL4eVLdVC2fLgfx+rLsHULCZgBJIyJTIRaDrr9cmZP/IWXTTVgm1v4tQj
txVay6yahWHGFGlJ7m3vH/laO3GpqZO4mm9voIKkBvx+g/ePbfpgpBXWT0TaSAvk
PKhLg83LMhyupdHPpLly3zLdT1mY/c9Uq+EiRyx+vjjVnhN9INzdPNIlu2AI3MxP
y0WJkxgmmkH/0Zn6CxsST3YUD2Uypo5rf9R+UPRTZYZAO5TKOeoSOT8bJjHhOCP0
TOuNsNAbDBTNEOVgd8ivIR98mUs2zuDp3auG5oNk7bUOUanXCZx2JmPOU/wkLyXM
tA+P3hWc9Imtd4y8mMLWa8oi6oyQaJe2UJO9pczE/dAnnSD2eNtg86gd7w/+CXBY
oz4Tad2beeEZPq8zLhaGvTf0A/Qqikuuwaet1On2iuiwThmNU3Ys/LeuOzeuaL0t
qezSAHM/Ah8/VwMDeTg6gQU1ZfiR30ctwot8qRAabjwmb/RYOYYPaFXSX9pZyxFZ
fr7pG3j8G5b00DMF+q+t4puXsZWVEuRA1g8m6flLo/qD0mnnEdxsm30KRxqe8pJh
WZ1LN/3Q25OmfrU3u8QZYdVuJAsKN7CBJ2fTanmpUfKk96x2L4O4kHfplVbPbqr/
Gx8AKd+EynnyTf1E04x/tD++qGSNPnSzv79Q9tdKwBNH773d0+lRuvUJPGxf5nHI
o9VsflPjj1p5FkWaW/hS3NswMOVP0c422d2zftHcflBlCFi5qRfXAfucAo8O9S7B
rMzNkiBGv2iwKHyLzuxRxrbDnhSH7JD17xPmwbcKkj82Xky95x0rA+8bogEyHSIo
6GCRGg1fGlwvkdpF24Rm//4+9g72gwvpu5hOJRjMa2K6yR/bL9m55qOWtNAM2Xi0
Q+78mG66rOz2+RALfD8bdTHxCfVhFF4tDn9VOaBGAt0SP/cI1aFna4XmfxHDl/gj
0kMoyxKRRvSqGV7Swvw4VMI9GKJDnFvyaeFaOoyyjRiARSOzcdFBRLyUfA7zsgvb
nAuzxUMmc/1erupWLH+eHZYokgbFdH0wkQvpuCdC/Tdb0uCdAbkJNcnHO5LQ29xF
ka+EKWuNrBkTVxyUvjqj4kOQ1iL/yWwJtQfx+nvGBvqMUvb/pFDxOoywXWES5Hf1
GKdiEZhi6zyJLlk+yxhc4LdAH6ZMq60CXskgRfh1O6+Lyn1wYxG51o8tMr1J/+/F
ri4Q0uAWoL673SzSTLbYa6dnJJShs+hJbwSjzqyRZh25CcLkemkWWxtgkE8DWIx8
uSOi6I0oCvsMUovhI5CqiL7flJIfIAhCyiF1kYh2Q3B/tSMpXgPCdKCxg6A7Dpov
oKDog6dUNgy2uIQJbl4JyMBSEXm5S+f6SVZc9LnAmQ0R15QaDAxcUMdd/gGznd31
n1KvwyoVOoti+IMys8vZC6eADrOL/QmCFQ9H2/K0WsF37FC5W9qYogaZvSFy0LbD
9is1EEBptReZwt9qvG47jJlejKoMo3szvxmMo8thKnGqbb4Vk83WQ2dscHMALcr9
J9hqmXTPZIz1FY1vgF9q3DAzMKHwR0t4rVXiiKuQR+GCsa4eODZT2kZCLcOjA42U
FskkkcUmO4aesCrYEdQLru7cBYAOGjLzGqq2Z3Na8hR3iWtummqKoYN2Iy7x0C6B
ToQ3dfE2axMkVh8j0GPA7oq5FmCfalAyhxxoPXgFOoR6eZKhuThtPfWjCHu9T3L+
Rwtx5tlqnFjiW2lnMuB3Z1W1M/Dia4oL8T9VPonbLaPLDA7q8kva/NB+1x97aogD
/Rni6E0iaMPTzEozl2uxnJljt+T+O2w0cpie59WQakwhz53ugWV6QoQlCpVw542N
ZiYuJGn1eKNRgMbd5pSuCtvB0qZ3A21qvOtBAhdX8qTWmA/AddiKYlrzWLMcPeB+
tqy60arZSkc/pPrOwVmFm5hTWhxVTVA1l/sRFslKw2u9GX8XfYdFauKlQjC4IxFe
KFwS0TpC1Jh3OWQ2ka822yPhs0hAQc56EjFhbEQ3W0RSxKKB/mteuPxFwhb/MCQW
CJ2pkXu/fJIfEmdsM7ryxnz/wNsGIxx9NIMHrLyG0x6Zt2XigmoS2chHGHqgRWCn
a8+54JkP0PmSFVfk/MdYvrYM3GE/cF558HbmqJt5wudbNWmuYcZnXWiRmSHuGkVm
omV7+TWrCRruXKpYNAypZwDtwA3J5rsgH7CAQ2rc2BV6ZmV8IJqBeoXv2oJ+tWHs
23ADGA487+XjTe2SDG8u40N73s2NHfVMr26GQRyGd9A23cwec4O3AftwmE2E3+TX
lnX8DZYNoftw/lfFFcTnGGLq4KzyADLTD+wqw4clhkNQYDBDG2tlVYjmFwpSSq68
C6bZgBajvImlwyCEWf4bcV0kTScQHQm9EuVdf7X0Vt3BRWwkx0bFXj53SCtK81PU
P3v7g7bmozUJ67pjsETUfnM9rWlgwcgHYLwPi9ArLEyPJMuzvxQ6tR6ebI1VjLso
8aqW7s44wx5aYgi/OlChllP67tJWDIPOFd6xneCEKtpRSPkySYMAQYvNgHBZv/Vg
q4DdPudUQKk5UFshpBef2Ukyogy7Ccpg/qESeHf/8GR2RLOY6O0PHAnBlJVyR5pQ
/6oBlsnyEyOO5FIjNOqKfsCGDF2h4X3vghU1WAoInxaIR7/tuMjCLi3w5Nlvqdcs
GTUjSNgW2diTLaXOv645CQEqGZInSd+eXzNpdjDBEYqjxEZj9FzXwbkZ0f0PCAqK
7uqoFcN6g+6ARgMlS/Uh0JZzh5ZsogNmBvWcXOZqQt5q5XuxhJ9FrECOSPci+SY1
f6Ys5CsS3XB7/9XCNMd/ITEfz5kwaI9Tsy3Yk+jQKCd0sLQ0hoBR+CDYJ89z6mx7
3nW92/XgI9a9OGoXpqOj3TWArB5l1jCDGplMYVnxukMYr132LDjg+sfJS3vL09vJ
D8uTgObcYy9FudUHCDG3hfM/LUQ2Ex2jg1LNFnjch91ZJQ/y42n+fQpjkOFlh8G/
A0NpAKN2D0cb43U4nry3HphHQ7R9y0yrmaHVuYi3GT1MWbkYlYER+n/km93e83/q
3ZgqHvzhUxK1EeIWTsQL1t63L6v4pHxWtC0n2sH7rHDOwiHnEB7R0uObi0iHebYH
ZmW6ooy6Yip12Y09k3p6GQTGo5gJbVM6+bpbn6UYwdtfqOVDUcO3LW6QLUYwwGJi
wpDcRCnv0hYpJ5QuYDFk4DqrYYsvVnqmh8M2Gpa7EAChAbQ00LQL6McHDArgtZBP
DeEpXrOPRiD8W1xdpYRWqWZIJKq7ccEhyoUTpeFSgFh+GilOApABXNHbnCiMsDSi
F5JBOSbe5kQBtllvaUWoOU2poaY9L6KwKzrYUAzKlRW2UigGn0zt2fVqKeMZK5LU
Vk0K66j/4PilUwyuFs7tBfJKInt/kebafGlt8wFXaDrxF4WnoSM0KAHjaWXBzT4/
EWqao6X0IzH+toZtwNBf/6nJMRo+rUu7o4ph8yeP5L987SgH5Fu+bqyirXWzahxC
H4uVB1MVm1fitQ9C0Q18xwtP6aJ7QYsRoT26oxMU3ofKzs+ko1Cx3uwD8HP+lUTN
UiMnsOCKFTBAyXuRUg9hD2Uf5NUz14+ZYeWYA0P95spXZuCA2zqCKHu1ZMUewNUG
yUvo2B54JIDx/ksZzuW6UEJvm9gPZmh1H7um2OhXmuqt9DjM5OZUvVCHozrcqsqk
BEEmI7OrqKKRPfBaGVVsiU7Ti/ZiFPXCce7xp+Z+sPMv4i8DmdfbpiM6WozoGOZH
ocJYC9H3RR4J2dyETTQARQ9ZbGCC6iddvUZZZ5eYAadbFqZY55faR0CbhNhyIk8s
/JTpmxuAsG3yyDsuqTZIBvfjJmSpawEXkI59ntrcDROo/+JMcWq3HubSoWlc46jm
eKpyVBuc4nJAIw6JZZMRjQbpdWwAKi9jMFNr6A8XVeLsy2DegVipflFoBgG6KIJ2
G89+uG5YIfAYRR6pnh9tGt+MgdiO/FgN/x2zEaiuL2JOi/oHZBsQHs2fjPhskU1T
nfpH5/STSASVLRxhFGEyoztSrkmRWlcovWhoC6jwQvKM+7YF80AidIwUidf1WGuP
tpk/kO2/YZ/E5MltoM6gwcgAghlBo91rRx38Nb/9jRKHjNj3a7nPzzP/O2LOWltA
WjRfWiMPRdtmPHiOStv700X6yN6qpU+1vsSRp0zMh+gi3xEE00z0F5a/3Xg0vPHZ
LrV3pvwkojw2SqNbmhTBeUfjZuOxis/i9Evg3YpXeBJ/rVarF2O2jLic66wSOjPf
gWh/7trRRNi0+0Dvl6QlWdeXVnmQZXVJhNpYH0T4xo873ZOKTowfOh/Y7wUm5nSd
gBLa1oG5JPSltfG3cYaaqzrblY89UubQwcAM2ygqunjCHpbUr1H7JS+33bkiVeIm
UP41CJhPEsd7cDlNyD1nEalwDCUGlsRvaQwkpdd6vLQKF0bO8X/ShxeG8OJj3BHr
mxWhmloBud+M0tOkFc0Sg53IbPxR1Ra+8Rwy1rV0u2GzR2al4b4Z2X3t5uKTnMrw
pwZ/KAePMG9koXQ5htCFsD9OyIbcPNpV3l8UJjKgJCr2Sx05iFBCMPUnu6vDcu/P
8dzl664rwkJKdQKnQBD49cq+KTnb3LK3cX/1u2CZaKZSFos0VYAvc0N0B5lOWpZX
G4yec7qJHGwsPxQ/ikwFZqlMcwgtBEGQ1rnS250OxizFsMYl906nKQ6SR0iuO3c5
Gua4eSKdH6EPyl6A8C6dk6pSDU7DKqbNBbu0u8SW0pNGQ/7MkVBat1b5swsT9kaL
kySCh0pbJc8A8v6uwi8EtOrzwIGc63BHg+CiY3RBSsMi+uIXfGShTXWmP6vZFnx4
mvqbdi7sQwrpR5ftmwnFmq19np/gv/wdIz1YGB5RajfqtwTq1HZV5s7zeL2ieH8e
fBUVWwiiYU6JUhSsnnzxyW7I6XnynfGmDit1nc9KWnq7psj4TqS/S5oCZP21cwsi
DHdEHzsjWL4JVBJIvVw4gV+SdqCoSuboINZrKOZfSKN1F/bjqhTE9jueaZpe485F
MTYkD+h6XY89stpC3c6V1OwXBTz6mMBaTKpY2JnR58yerqGQmQX64XUEtGRsgF6V
gp+YmKx83O4RjvVpDH50S7T0WVJaS1xUM5qeMiCATmX84DZUXRDhWzCrbqhZmnYP
tM7cWhJYep+OTLpW5TRavu8fTAJKvQ4gSEzGiLI6Rj0cR65pkw5bTj/VwJmZlcBA
9xQyaSkK9iFq1DXTic9Sz3tbsAOgqlXEHELehdtlGZ5Oo8goJeLt/85RAQwUE7ie
ZxX92wFdtdw9r9fWVGGxql/l35ycTJULMXabZms3rvrztVb9NLuQH4e3BPKAT1lK
KBvmE1MiIusHiDBJ6sYg4ckWXlTe+v06QVd5/J0+Sy6m0acZJvEAbtjIkydx0c1/
Tptd6vp6U4v8hshXIPDcLaX6PQeWQ9uDbCikZqiRZ6EiFE3rjZGvAKF6ULPSxcOS
P63CeWPTyEC/lbm0PIQsu/SII5P/RZpzegbldTUA9ho9QJuQnlvfEmfMQvqUM01C
Vrh9tZtEs8Anl2XMGwTIaDIZ6tcQQeJ8A5cV8X2lD+n4qvYfGKksacBfEhQFiLqj
1R0+XzUee8xjzs9TaQ8qegRZsL7/JNAO0HR76o0hEePcv1xSZoJbOzBYsNvU8kqj
28HXI1B5Pt8qKjSOl1Vt25eocl31tiHPwxx6MwQlWWjQA0xya4RL72d16XYpVjqN
KUZbafWnW/xdjC8f99SQMs7r/eyMrLPxd7KKK3i3j7D9EGJzTLtEdcwCLv5SJMSB
4OMTQO2QNUnEuoRehyt8cd5KTTSQ9kNGrzaSeYpCZDQ8hQfFO8d66QWifsVQoIyc
23iOhCIdYpv5MIqYUCgIwH5ZnqLjx/E8mmMH998ltBNg820kuaaeMKQIHnoVTm1q
s8A9J29EudCuE0HI1/XVG8rNFXmYC1ocHUXvlsJZ8UuZBQatjQ8tXEY2Pecerr+A
UrupYIp5jYRRqfs6rFN2NkxPXW2rv43rNk0m9+sjL/avSA3cS5Ow52tDh7UyiQwh
K14xH7Pkn0aVpobfpBOboGEaZy3x9wufZ3MURq0+nK7thVDiHtC0aRWbpb+Mxq/t
CIo1YXhutCkEi7VWedmyN+rFgcFHrNXZtLq+avmTM3VEnPeAEDSsTDvCu9s+KNtE
BDueTiq14qpDwILTxL/VoHhztqmsk+n/2dclNFS0nxYWJCYX5O86fLEeHgk/7IvT
yz9FUC0oICOAcrSVV5w3fk2PDLzpDIB/6AAnABwVk7zYDvuHHbG6ymVi/Iz45115
HxOaFo64EgNurWOs7cXrK1bCjMwx5/nV65hhACFxbnAFKMP0FhmeVF36GURMbKOn
NWI/h0kL8hfgE0Cemt5H0PlLXMnr1KX77iQHhOmZ1m1Zi3N/3mzRtFVBzM9Uyd9N
NsArsKxUTtzf/2PasGSGymp6kKhBh7+W8UhQqQZtkGq47jMDjncnov9fFuWOlfKB
6sT39NIP4/iWAkh4GZ0yJoJNh3J4Okbo+PZGToKC/xQSElMCdbZw7yh/cVmbBeHR
SBQJadjkL0HiRAKZ/eHIJnzXh/xr9XM9JF4TYH8HMdydrunmAwDR3Ez8wRQ5RpN7
dv/cecKy6onQihQ/fuKSIvpsFm4RWIVrAv3KBEh/8gG6hH34ssbBlVkZi9tB5WL9
D7bTnV8gZj/ajRz1wAlZB+u9A2TMSshxIwenv/nJYXh//EDzx4hvRSuZgd1zwHJP
6zMT2K+UMGWrmlbQNNkyi3GrrPjnlRtKYhJJWQrwDAb3mlrCQfux3tcfgTqdKNYy
1TqQgCaPwMJQ9Xs1QUE+2lhoPt8yx5vLg5ioYMshl51Oqr39Swy8/wNKAymT3tjq
QaK5orgnE8/jIZDVAoIIEuIEcOsxsUnywlJpaNsaDwBFte/H9XNsOVd0IBFHv7YY
l3o8r6Au7/m/RpLhz+42IGBxZsIMbrPcLZAXY/AE9z8ibTGmnSpxdiPM07SNpOa+
YfQdDHsyET/09HcDcMSTq+cNiydMRj1EJ0EXgE9+Vhn1elep2pO3JmBNwYpG3OlQ
gtKGsU9zMB8ppQwkbgaVaO1VU+FxB+Nzly+Fr0L7vYjbUmCOh2cE48pUIMFeDyQ9
7a1dtubn37Tr6rcNA7unj6ift2ymX1HTsdkNrWZ7yBK0pNNGdWWff17TQ+kysUKo
O1oNP5AH0+h3AhjHez94PfOzoMcq/UrSrN2ZiAkI8ITm5FUE5+tV8IKAWh4VLkLd
D2kJPi1DlK9NhxNZRwnLsE6miucJZWx8isU9Xhs8vRVdPyN5/CKwwf2z5OsfJYfm
5xHnQQbDiUA/24n8xXRL1yMRyZjx2sRoRWN2ZAh4rdGs8dRJVkrKnVwkAPKLvoH2
hvfEYWSjAPQ3wxa5+IxqZb51oy8QgLCDKDrFJKnPslyUUwlALG8n/ifTxy10sxIu
zspMtrSxCuQuwnzi1uOp2mSX6+GBkfbgjOheq9Sp6zylGuPm9ZzWp4baTXJF3HFD
BHVNSPy3N196xEzmbSojjLTw4tgznbOYEyBeSBFBwZe8FAv8kLCp5SEL3UeECLPr
6/+4/ZsxhS6bnF+dy+111uJyEJMdWYdG7T983UE+jDymnJ1NcVDfgoLnR1IPadQB
0ngG1PX1pCQze4NlwSXXeAIwnst+vuOEwXSLmXWScLa/ffYguWcVt0J5Hp0mjU++
JaiBZTf2XNcC2tunniUdCzjzG4I5Svs90MQlyx5fAl4P+h2las4vHI4OZLjKIrhZ
lcZ6qI0O18L4vdWCNnqGM5v3PU1F6jNpYTvzKU7wr/6q7BCNotnHWXxPROinnGJ/
weQd/4ccmUqVEXSMju6VKwPZ+VsMv8YkFnqzOSIklsUAizNJ6mId6udX7rOKTqUe
Gq4yhO6UhnbiB8hwHwY6ZY7EU8qYnOhAhv7Fwt5eVIZDEi8pyM5SKEj2zHW/5AMr
SUGMlzWd/IvtqwUxUHSBZDWd/w799ffFtD5rhNP478kTQ/TNb8UHFLtsqKI99Oa0
60jbfBNtupTRiXp9QcNk8NipQVNAqkGDLPMtNgMHP30I6MHuiBU4av9xyafDbbHt
i2OiNAx/YeAzEtGadXWoRaonJBh5hBe1eFE1LhWGBhCC4ttviylb9hifvPO8c3s1
DW5Msezs08RErQnPUq3V4VP8ZSIbfAybuR3ElWp2TeO17U9NHeoQtUOgjehAeAz4
QlO0n6GrTiB4QwZS3xNifD/v0HvHObmvXpgLEhr4KiGAVPlNGSS5/3os3Ocu2A0P
E5YKw5DoTTjy3h8L/r++HcOYppLVWnlr9vFmdFiMZ8VfjcTLK3w/To7IQMTzAjgu
WnUw8za84gFh6mku1eWMFvXYfzXIXd2tdITmFHwajjYamPWJ/+TYHW54FY5LmQds
d0m7r74EumbWBH1WLHu2Oi4/+6fHWsDlXtCJR3Wlw3+3OgqVNieIvZdXso9FxCUi
lDBx/rh+kFnmJCJHuJBEPKa43dWFUrGFWVYK53KrRvms/VYVGLmbVwQob00+ALjq
AjwSXCEgbvX1o80ngqCphKHoKW0rGxlcrB5sQ+OlDwz6fe9YN9gKbZJKcE6PCQ8a
5NoSIDd6CqQ4vd2rjQfyL9Z9RshzNlKmc6MAvfQlM5OlLOUp0BiqMHsosufAInvQ
Thu9qjtmKJSvMt8KDk0oqOJ2QBPZ+NAUKTRr+rZjvSOVuMkmB81FQ8/lSYw+LEn0
Ots9SMwnJAaRYh5CcONcVDG0FQT854Ch4F9kWZjM3pUacAzuc3VAuLNK2z7JQRIo
J1lXEcLkz+fmJ3CYCRj1ICTvB/t1rSJB3BkVvYeNoOJYOudjFER5p0h/m7GbGDx6
+HPUBCRvdqwatmSA+DUW37BOV/UVnuRZG2fiaumkxMgugWnmy1bdbO+XybFQy9nh
YYko5YbHUfI1lkRux4sDrc7oxM9EV6TClLaGxAW24V3JIqarWMpv0Gym3deFlzot
dKowQkhtddv0HggeXe3rMcZ07w3iRID/yab4rC7aUgEawmb5nddOWh+wznBzUyNe
cSOuSUbmtowqfPA9D7xranCzLqbfRxvXwQEmIfk6U1276qU6zqx9pAsaENwyXJ9Y
PqM8fONNKHI88q9uhX2O+Z/OnBjWY7+Vit+yWvmasuXUnqYUIRaK6UAHBTdqkLIr
g1/SzSpTqGUFTLhj7Qhr/UiknatkqLXyENcASGYRuOE6GpeLDWYlE/fqVrvDSgm/
1Yyj0E0aPrCxP5GGSywTRpF6JNWXw2VWkRZn4W7mzQrNUUL2+9jfScAyKvxWCGQl
edlubi9UACeSWouUryuiNOMITgtTk62N/K5+q6WID8ycobQxy2JUVkU2VtGlZS/0
16HvgXxQY3nYktVdR/SNOp32h5KAss2pffkWxU5emq6NX2d+eG+Rcd1hzM9sVD1X
M9kk3pP27Od/H34SFqq59NEQ+Jc7+g2vXPVcT7ob61bq7C0Xzd4f7cvCKVHCuTj/
aQMuIAHcIz8dgPAks7/fnNUdHHi/tLd3PvVuM4yLKNh33jHV6Si7NDTQ+5ZYrWIs
yile0x8FPh0DkkibU3WQAkzylpT5bI+4rJUoGy8YPkMEaZtKJBx1rZGG7QWQslFA
F8HDXjHh6hGiqPdWllkBEtGa5wQ/ZNCjEFpPGdA5YtZcM+BRbRlTHkpyAbsoYnDw
8cvCjeU5fMF9s1bNAXJFV4yiysCWhhFjqE2jkfjjUwwlxm27ZAKoTMDiSySpRxjn
o1XIKudoERngVFf2lVa1778Y7Y4Sr5IqLZaHNlXrvqtLfPZfLHDXbdcx0aHV3CuL
WyXA47q4OgSqT98VqJeFzi9Q8aVTLqHbss0S8wmGWkR2SB8biSfI+lNHR+0RPKTX
7YMdsuGdRZ+DcnT8uFzH/L4Ya9wbpyPvaM0r2v1L30jL49cNFry0AcMkHEeuaW9+
d8wi3XNn/lFcbKcx+VKjYHnl37yW5n9xHRSHYwjWjd+M6QiKko/qSz5zOWkBwP2K
tGm1XOr7TmzUpGOlBvF+QQEBa7+DDpZ+k8UlYr7gc59EP3od7MWcZ4PyzQiQwDvl
cj3jU9+Zty9jz+5y+5xurLLlitY+FBrOipyt6Xph+PmfOeQM6x168p7IOMELsDES
KC+yTMKps1VONProwXDiOP+sjvpIuijXZtaRg8IN1AoIFb+DgWDqQVmSyUzfEiCg
e5m+FOrJ5rSrh8c7ImTZqYB6fHdedXnVxDIrf3ZWQtiiIsQVej4hSBcPhn2x581r
RTtYlbZIQJJ4+zJXHbnR4uyhZ2TVo6bLMDzcUya7uJTVrjcHEpBm9IBFbu2lrLvd
I9RCsncNtsTdUmrMpXiVPTNeJuKUOs7I89bcXECkzeU1poSF/2Fga80Qrt511EVs
B1f4P3fdwfruySeuxxoFb5YJEgYNNwjEblL+PcOcLA+a+OG/6gK+W23578CXBcym
Bs3fFXab9uRpyk3eujEVx6DTx+Pswvq7z8p6DTBK9+5jMkK7RNegUfr6h+XR7q8k
AdJZ3ptvCwTXRzjgJA31OHSkPuBLIH6juWVU076TtTEjm6m5Yg6yGdSVcsJmOHlX
59sfUwpoYC9va1U41fGdo/lpkfOF/fGhnjbYyzr9s+WqALxYtjdjZbmnVWRpsHr3
vPOsH0SAv86iHbKULosPUndYuIBfyQIbZthf6kt1ckM+YP7jbP5NLxclwH3cpzGa
svgu3iE0WjY7QThwzeY1bSoSTz9LnyfaWKlg3qzxZaAtSH78hyoL99E9h7bdjYkh
5CuaWBFgbxKWB2+LhAhuhUMScuoQywD3sTi+ZxX6YlTrIVx/UxlpsubTW4Yi6IF6
9YYzEp3av8E12prw+6/vjYdw8IXVa/FziAbXRfm18YhC1+BsOCkwrpwBaWMxWDT5
/fcXNpzlq0ocS9/67lW8juvzl3vx+466Ku7QNr5f6QjyVLlSCpUunOaXShmi2zOG
huekdZ3WK+uNlMeywEcIvVi6RNueKlOWkmTW8z6RuASeSyAKFkMALl+u109blacC
inVdzymKJPqve8/BN3j20+eToGsslO9yXTOtCo6RwXFrrFb66o23aAyiCkq37BdX
Lz6B4TNGJsNQSgZFb+tTMS2HgqJaGJhMo3Q2nTTGneNStTrlnDLHk9u7dK10AC2m
cNMC81fc+7HWgEZZvwlbFWyE08El2ZroQNpLgYNPDXodi9MGvlaVWV8rrjgn/RY0
1UHDBQT7lwEpDk4UnOOv+YtQ4G8S5MOyC6P7xPcXOl32skUMhS5dkXeIs/M5dfgl
attEqxufhepJ20CP3V882m+GCnjXyMHgT7SapvyFTTc+35Ane1SM6nMoHW4+tuw9
R4I/448N6VJeNw+LETdk7Vqq9oz5VKrPMKH9siBgMKq++oMcgBDc6Twl+dweUKIw
H+YmFFjBD4146SLwrABjll16hx1ixx8si88ib2qU81HC6NlKRwB/611S4bsRu2wo
bx7kOZb7LiJTdms43wBkNEqFmnujcqgwkszNfUNlEV9E+/+UrugZQtqHKhSn5l5O
lWcFn7Sw8MpldyAL17RCuN6FxPXt8vi2REl4m2Ob/v42O9Bz6qzLKBaIpOmSHLyi
Wjse9kqA0wv9KYKA8oBGQiCObafLkvycgsR7Rx5RoMgQ9wLgUnp/KEpGFuLyZANd
KNWgWXkKtXQ7jnkGhFmcQK0/GDzrL6aBrSXaA13T4lYHcht1ib8bvDVxDxangv+T
PVF07Akb0ELs4kHklKk4ywvDi2ZiMQBpxxbADwIGDNsvJTEPVI6GBegVX3FlTDs/
b3IEE5kRx4voD/Tyyq6h4ui33ODDYWIOazaPw/Tf25Yo+f6Eyi8hWadOGkLO5LI8
qz7qe40Y1vc//b05RvwcyCmRCz16/D7EXxjN7CEXOFfw4kWVO91Lh/pDPt9Q3BE+
i5Dgawxapuezr/i+lmYFcpSAK1UaE2sthc1L28r121wY+n5R8xedq1F5QEPHvEmH
6kTVUAZ9WKyV/F6kjE5OkgAUOdhlsYfhH/5w4x49O+rPxCq1XWc4B41+ZZg5cPen
uUWjehu8f1lx3wI/m0oE16+ekUs0JiHfZkokdAfRUSPFoMp2AxrWUZHR8Wo2T/ax
X7/QxR/AbeI8+t+TSegqKoTcP400VJhJkyfL0KvnBdv75lu+hgip78JRXr/duoEm
r3Rz++XxsXW8oYHa0h/iFLkYzkTroCmNU3Ewp6jF8Nv0Q4/1qjV4n9QXYw/aDukA
EeVGstMMbrhQl+vYMq1EW2/KFCZeiJIhbI/hP8WfPNVOny3PEWE8ZHTwIfw8M9kB
OPRaVAZ2pfJXA2KDXCuDa27CQCEcQ2t1lVLLKjpztGJahaiSXqSgXIEVGAjdzZOk
XsTcTnhuu/fqCd8ogRpmYHDyMZMz2FeGGcExi6jAUQ4crmWNn5LIEIlSqvdkoeLh
Gcjy6oYTmC45OaXKXejPtIG0sBf0EeKPIW5DyiWcUF0Q0HwmBFPTq0KMPv6JUsGw
gnrqjsuMmNt/4ELnl6ULC77WCcLMsbHlSTAOwPoMoEFCTfMajqxyMbjHXb6OKwIA
I1zLbenh+0YCD7LIbV3d8A1R4/cOCGup0MO5IbRRge/+3PNcexXxrOgqK7LAaT1w
RQFJd368gda6sizHetgCZeyF9nI+of5rzCrZCQmxVSK7KNUCIFJGdnMv33mIFs6v
5sX7lBbN6us6lYbAH0+YQCr1EUVXqklotiJpdkuptoGhUCJL1CDGD31rHpfO4lvO
blqFDjDUh/TBQgqTshil40FWxWijRXyfo5039exF+DNhSzGgOiySbGWq0tLwyiw+
vg/xAPaywyWsiGorEYfeZ0QmO+o4rYl/ONfr053G/hwhX2AkD7JcZQyunUQOTR83
YRsOT+GhfMuZ408QnJgk4Fo93x3ahsbWlibseeuNsxuF+NjAMPRvpFHyPbawwdZf
u/QdiYvxYk54yV2QbkHiovPwKx7124iDljPLWxJ8LLWxV3THQ9lmHZNI7zj2c1pb
+jV/o6rXJcFNSV6Pw1Q0RNH3os5k/ePBsYEx3sBdftvrW/F459rfMBX+ZZ8tfKlV
yqcMFwWwcBXO1oET9kPS+Fpjd7VTk6759PkNYAbPchildc77R34GygXFwfI5dMCO
tcPj+2VYR2XwMg95LbkkWZPOyS7f+3y6e2I0Ry2Q89jxtiSzpEWMzGUiKMSkUuIM
qKd8gFOu42m1Z1qJcxoS9EdlF8+fCb16Y3GIy5ikixpTQIcfRQuvC+ojwQr0XAeT
81SbW6LzFcsbWf9gEz4iHU/C4FqTuPb9hA+t7ukNs4MipM+aGcl6am2FWOJvbAT7
2KRzVHxKWv02xTKhL+lFM1B+dkydB+ZHpvvPfWbfjMiRg1GSivasgDpk1irE0wgA
pRPez8fXXNKIshERqjGHZFD7xFMut0txiu4hJiswrCevO2m3n1dhadxUjhe07+D2
wjflwWkNhBoSXDSr1TnoSxvn5fs3CGHr2YBQJht3StYQ1FDSHRotjCQHdxBRGovb
lWAcuaXUbFk0xQ6OL4uJGY05/qn4kMwjQELhjBSN7HLwn0W518tgPZ6y6k4jMPxz
X2Cv2ggRvB7pBmcKMxhEs0RaHREq2fBruvrl0Nrn7NKOk5+O3k8WLamr9hs6J6aW
iULLm6hWEBBtvNrrB9Wg9oII9YwuVaj6SVqihPnAWaHuYv2tzzfB+gdAk2KhaJ+K
47mwQIKOF+yBV5nWTTAx30YoY8cKv2zSUqyPi/OELrqurDGLQV0LrCmcMnSIZoY2
Q2uIGYMCVGNgthgSmENb+k/czEYUEu2OUQKj83OqeIG9SR6ffATAggMlDKX06FhL
8incoS9Z1goB9qpby+5SAl+Nqk2ezOjEOFFbZ7HQDZtE8YfG23CCbQ+xRUgc7tvt
aGcszyyq09OfQWfMs1oIpYMoBy1Y+sqPbXKazILZjdl5HrLWHOILgNfpA738Mod/
Efbh0fXtTmTg0OKCeA36gN5/Va3BzeQfSXXTOUsqo30NrT9LjiuGsiKAjDqaktdR
a3nJZ6nuHIsO3OsXwMTPz2K97wzElsuAw0sirzYNdni0yAG5uSgxC5Wq2RBVYloJ
H6ELHBUB4WCbeh5GGZAl0ehuj/UkzNiqz8S9VauOdF4WDkxlKETzOxx9a5XWrNTg
bpuee3NEeWip21YF/y84vWLLQqL3k1YY6MPWFo/Dz2bUKhF5ZvTnPHNDNYqZI2nV
cCumSaMnbfD3NDEots9NJWQ6G3tFMUblSgHMneFOWY2HSJ7p8xt9Zcvb1b0MxGzd
ztduYGlkyUV8oXENxek1j20WtXp76aqzR83Ihr78ck6SXlobVmoGdd7cv/iu9nTJ
m44sCo9MqgNfF0T73dImj/DC9N1erthaDqvWYuz0Lmc9q3lmUCsq9wpkRPV94JtZ
tA06CUtmi+0TpS/xx4x9nN/VYKw4CYwefiUD+mgjp5ERs6sWhHx60szAaEGCFKVo
dOQojfD95A3gcrd3M0Z5AkPal+uk1+31qDY8B+QIrtni5Gq6p4lYcA4+AV+zrwf5
MYLNhfLlyxLLuT3ZNi90rdSmDIUiSJ0Pvdwir9vMFeXBwKoumRuelC9kEJpU0tV8
wOC+P6Tig7O6wNF/rdzcOITp+knNr9mMHOHJ/DQgWm+DEsJZapcSNSQ8Ru5p9qO1
EwD76yYHDSvIfpQ91lFe5vPZo32MXks0tZUOzBMrO3/WEuMDcWLKktx9GMFx84eq
2nWpVI+eCJOCIs828AQkc3OWn+vt3AalsSCQLA3pRa9MJVmlGv4pufGAeNTNmSZk
Na62MQsKmTEgkjdmg2aqq+swrw9FkD8UVXkg+h7kFoXEMabod623dKtTeU86tGnX
KI5USLPjIYiZ5MyX0s3yi4kyDnWSAuHUbCQ4q0gf4VdKdEqwHIRSjcWTNClkiiHS
6tjHMt8N0Vh1WJyGnXEtHv9LjWiAAZpt/ebgKfO9ZdCYE5FWLgZaDGLfhMTCtQV9
swdENysbBcvGkEUoaLcITs+P7WJ8n1h/ml+OFnECCi6Ox4LA/ZpWX5lIa/iw4lID
qM6SmsgjA7inXus1wjugQi2O3BVBev/HkU/McD1hP0M1HAz/crVhy6l82XpFtUuI
R6bk7Du3Hxhvnx0z7FbDDnQn1e5zj+/1YGZRvjMsU9ZhLCSTPlbgZAyknCrqFhs7
FBflgpX88u9GDlz77b9fFmv1dfoj5sGztjnu+PgR3VF+5Rh3QzVhwZTOg8+7MZpE
qEOdehIvYQshKRgphfdTDM3kBN//+AVInr0opetVzYO/ntWxEK3wzzHd9lHN70e3
cd9GbdiMn6+0J7uRSsUvMKera99uwMc386pRH+MK7gQ8J5MKV94WBn71I+MR/xTt
KaJ8GEunvQZwnnkrwY8M7dUgqa9GEbugSqPYCGUL9+XOnNUMEsGe8m9Mgi574AQF
dYqAYu6qT6zddRyZL3m1NkXvZ9TkOZflNQNxYnMvDVq27iGt9nrMLWW4MCs14h19
lYDhQddngkjaCll5hEKV2Gj/KY2LfnYsk3FOeL4nejckIVqu0zBj1H3RB89ndAC5
v34fHcTzpfiBBxE8wt3bwD7adkEvXuUQgvGCWN3QwfR/FYAF9bKzXrDZ/PtUe2np
ZD7iKcITxG7018OfjYhx8SQCtlzcq/OTwTFUiva6gIxs9RZUTsY7N4yrNpOKRTAh
59SaszlzxqoOyZwGFm3qSd9jSu2RLqetRVQyLOqGlbGsjbr54pC2MB7a33BFY+lL
jzHktewyimjnrc4I6fMd1zdonAbv3oiSpv4JT8Zno3/QBHQcudq5IlczZKGtzahn
dDqDaNTKlbdF57XnoRnvvyQ15Cv6YJgL5DAtT6QuXcviZ0LMwvf8WRSkrBtUrlJt
5tYTIKtJF4BBVHRF+eDZ6eBu9HMrDNpAmpLnN3AwVZxcvtuOXdG+M+4pLxmHaWCL
4Wg/wAUmxKc/snyyke0KEoOfj0IinydILr3xq0JtXvYh6+wt3cWRxzTaWN8WKvNf
mnXKPVAV2GlZkFQ3ZiVanct5YQKaT/s6aFStTVGWIVeiWSguzmaEzIX4L0mhPnbI
uMSRtTPBO9bAZ4BJ0b3HJa/fgD1dt/rqlawAnJDHkOzr0g/ZPU1Et2EOyu5yyJXb
PpwW+8aaLCextvsGkz3g3EnpRK+51jObRTm1/P4m/bfHnzEgU+h7jQyAyEBsXCHQ
vBfwwC9InuYlHaWZhxDTvwaqfgwRoxkxX8h6TGOEZKZjLzaHIZ1SBMhYlt3hbifr
PRvLzubAKwLfJ+F3DlECjtsUh/1coaGaHIm44iacop9FNgj3KHvLX0rZOk5keCw9
RI9xKDyHL1z6Wy60FOT0DW3hrCatvGQMSLwmioWgqZ+ojiiJI7ySiTIQn9nnIdUR
/izIgmfBda2jM0q3b/rXyX1Wth6bo93JzxZjp7oGJFCPB9Gfn2eUvrF77sdR9PQn
RuadEZoeghkVD4MO7uMfyuLtJh29G/sH50bioEzZsyIbHcoyWdCuaTlGc+eNERsy
k0JaJBIHfd11A3mVy70pXNi/lekdsZ+GsdzZGSDlXbJz/3ApVGC8hTlrCCZXNZnG
kivPsMFbC3VtQZN9ot5O7CWkYmjqZscC8hOnqWpIY6/UZpeO/uzgGKd2MM/ZXeoq
WLJPNFD0uHHb3wNk4RAu7y6Dbm59iAjdgK44x8tGDNOCdxtfaH2GkcuFt+schXO3
jIXEb/2cNEJ4zKSA982l2mY6vCABO/CxQc6gpG2g27/44zZLyTeRdcrnwtwGIist
oa8czo2N/ea+kocvE/XslHUaPShQZ6O9gX4N981O4JOwjyEu6NLMTOkqSGfHcCry
Q/NJBg5K/Mg/pRWoKyCY/IFcN40WfUx1iRc4PJZDgk6NVAHfh+xXizj02FAVhp65
8yUG6NX95v9Ilr6Y10MJyvwCD8XGEYFokZbpkpTkljNeHW5QI+1UJhsQenqB6zLs
yUZj0JJb9lU7OQXxYnbOA2eA3RiKfNV8GI38K08DadKyRPgQVvFJy95Uh8Pfafyy
tDSez8b7gfSrk2Q8bABiE16vo3BYHPOjIue1BMfLyVOA4SNx1aguh6wyFROpYs0K
mv/pCoG7iuJIR2MLEowMm8q0o3DhRCnJw2bupeiDZLsITUq3DmhOvDarxAbVuFWR
ke6uHHh95PDNVJzMGbbMcnGnv6L9MUeN3SX3gnFF4p6nnJ30ikNMV+6O3668HVZ2
jeS6Owvbt4OleoyK/V6Vvv0eaRBTni6D2FHSM9KOtsO3j1gsjvdryYX/FYcCgePA
IxcQua48jy/lOXpab9oYmkQQD0+1tha0r1TOFdSuArjzcBoGSPdwobqaDWi4lnwU
SW3AgcyH+n+A+C7CesRJSw329P2e6a5i+P4FtUjhaglkKwJLK3hgoqpOYGrck/e1
JM9bQVU+TJns8IBgPAc4wnOAJrvdfY3y2RTFTK1HqpaucwgxwzCwK/I4Zlo6h6mi
bWvcBZVMK9Q33xoLLDXTNsSkvaLAOZjmS+ComFvZAopj5fj5cEKl4Gq6hf8j0AJT
NgckjyOD6XBMRZXNhhWW9WjxZ80h4m23UQ5Rxo6mybGwrsrgCN9rr5gIAS3fVFQ7
wkOvm25zNPKWwU+Xt61hFkgcz2ocM0pHxi4ZaMJuY+0MvGbT5o0myxv4AnEYcjsp
4Gn9ahhtui7ywWuSA5glBSfFMmQa9nWU5to+gNMPWTqtzRDO0o1UWEW0LR1k6YKZ
8hBLjtzr9nPZbA7B9YFohkaHfUWQJ1aA3xMEzx0q+20rKK0x1Jejznh2bpgjnsmp
l2zY5lNN9rYBZZmN2w2sgzY44NkHSvJOU+oz2XgF/jLERT5csPd43NUYxR8h77NU
r+kqbMvispYtm6pp2eJ+tz9sp75WlbKM9irk8J3rI3HSSfy2uITxNYUnyxY5I1bH
kBIMMJfP01Ooh/psvI8XslUP1KqV7pwMmOn12DYMfzzpT5SOi7Wvv6tqY/C/2d4W
Xye6wCi2qyYuwdWTjY8gnBJ1oIt+axFHmkbgv4CoXp6Zela2Ji1GrhbABJ6HHtM0
ckknZPXRbnoPFrzN8Tp733T2KO+z+Cg+041UpVxsu88jr9TAz0b4ZEwlO4Ze3v/L
/vW40IuNVaY4C+DG/ZxmGnPcuNqtD64nTNt9Y8yAS6sO2nlrntt7yJsyp0xOTPNw
eFPqIdL+j6tbyfG38F35jte+SED0qhBxL/avUV0lorKyza6dGkEi1t6ihJugXzzj
lfy/qD6ZRShrj+ca1T50CzHpkz5NjVXNe0K4f0N7+GdP12+kNNshVSqiU/Ayafso
uAtsXT54HAo2R5IpzTi5k0pdMODRgys8MJZhbhl3ajLmxa6GfcnOrtHDDmylMYZW
YUF1J8PAskG168Y++GMraG9X36pDJlDnpwXIfQ77UpqDjIxwpQHJfKcBVEWTgQS+
oyookVx3nxT2uG5dFgew/gt4eAJZ/f+aJzQcg72GI/t6IARwcrcyCKpJCrh5GawF
Rcuqe3tCexB8bRKp9ZXfGjIQMHCQCfUr+M/yC314D+GFdaSNYjT0ch1Rf7EOWSD1
r9esiHtZGvdSmMq3m0ATQlHaBsgAYNYtmrM18hbth1G/QPCa+yxqImImxIUzZTRH
UIEn05jP2ArlyMkaxS/P8/N9K1sn4PkAJgv1gMR7+mkFGbBB5WRtD5rp0yZIXrnR
yyAqiycoH69yhDqlrjTA356dsUx89aWnGVl3Yk2a0t8z4aaBHzcvk+XDxKDYprev
ehzt/D6cfPqFCgTgD439OcvJeUzM3WjdMJceCKpbvUqmcN04Suo6+f/AKprz86ni
FqYG7zR+aSwG3M8IsH6f4IscyeZQhoSOammcPLbp3wPlt36VzPK04EjICBJFbCxU
YQ9ZBasHWj4M0nV3czAU2bXt6EwCjQ2lvrs+t6CIbmSwUkMt/rS7YJdzGsknyFwh
8EI01Ak47UPCSCueBkTXujlNmVDNJcvIq1W9Z1Mi0jc+o10KyOzAdcogLXjpXwrz
pkLi+lR2l/5xMPSrJOWljhIFHl0Ef+k1qWi0YfMsvAMirwPMkEIFtkCSr1Inkyc9
vQQ73YiuiECoHQ3o2MAHoPKXUayuuvG6A18N95iGLSxXwW9uHxAzuuCtsd12UrYG
kOPux/U7zKhvLRt23IWDozy2dRxpq0LHqk+aNZI7PWJVnvvIGOwEQDltuLURwTTL
sq8RlEfd+jVQ1CfJzwdCbH09B0o8DBcvH7ba8V09KXfQxBVmpmD0PPF6zrbXCOsg
ScteMKcNexx5k0yP/Bo1uPZ+MuvHDFoeDIMnmiuKI5pSviNapaC5D5rnImsbAuqy
U0GTmUfS9KMs1L59j8eDYICIcBywO//dkGEw0yc2xUWXJ64pKDaljE5448PRwJ+E
t5FBN6Ois5wHI88vYAMThMWTQtTcOdgn875aP2fUI7Zdn7O/7AzO3fvU1mPkW+ci
WD9rasHeyC00PoqkfjPCvBZwC4QPQJhnCcTNt0yTp84dJEN8aJbKzJskzwOJdQmt
hCmwc/3OOv+UuXM3R33YQ8JK+RUX1CrEO4Au4PVmK2QpWQ3o2tsP/E/GzhfTloDE
2ZbXhT8PUydIEuEZ6TvVDoNDAi9taWWiCK5UUhgJsm9x7gWJqUuAymMXHHshSvj8
Aa6kUeVw3EYFniT7Rcdm/ADttRUMrt+TarUTDoT8AZS18pCDuRluAGqfz3Von+yV
Cn7DRR9bUenU2WycrZQwOt1mzLKjT+YXSYUMaGg/AZeFO9Q3kjcQZViciZv5tJUN
Vuc+NHPSvR9YjqJ3hj9s6su5N+1UMqdv9kNWsw1PSTUOFUEgts9AbvkHeFk1uzWU
rB3pj6KIh/HMnSAo0KiQpbvWMacQAbEnSZTZa4FDnDuO6RZLjQDxPNwBciP62ZvE
8vJPS7Zs2j6hRr1cL6jbg1grOPC+VZhMvRP0pgBaAvu86d5SmaI3eULV3OqSq+eH
7+Gb3TzGBdizoL+D+Xsm9NPUPJJeG0+HICiNSKry/vqtr3qFy45OP3f+G0qOOe/O
Fao4WJk87x8fQEuZnTPfENYf7AbDNZSA9isstuO9bN8H0e7rw8im++Lhn4M1mQgS
cbTMnVgpLkaHvnwaf+I0Rz0l2Sc36iJZ9ZJJQmuw1am/QH3ioyisKuBkshMC7886
2AiVp471LDdkNcABX2BLVciS6C38fQwSmwGrGYqHGmAR3+ZgQBKJ2UpXnsSyTlmR
OYD5DkPkw91X/VIBfsftduVn6QKp2POqnd0e7A/8k4RHmTISurLhlRawXDn4GmcR
qcvOwJjmcrmCBn4worMmNzc74yPQ6a3L0R4ptVN/CP+CnVz6tray9Cg/5tObZdmd
EvzbO5TzM1+vbKoAq8BVKkJ0ZlmAVZY7ktuCGUQrp+qz9YWwqZryy4poO/s/Mkqe
8AQGr1YXO+s2wkTB5agU/BSI00HtXAjx/OSDwLObun0EgNN6UZCvtfNPQUgsOTue
SeGVZP0qaLFc184Yh3SRVaVk6ILFE90hi3EYNTaz3UO9qC35mY9QJLFskXJQTN3c
AxZ7hdX6zgQN3ozRFbYYa4awfUpBCSaeI46MRStCXcWeXhBHVzJf3C1H4hiF+eUL
WlF49cWcc2ZDIMm6m2PNGlyvo3D3Uc6bzQrquK6hYhp3rxUWtZg8WfcTT+bA66Bt
mKNLLbk0xiLRXpcBHXv7fgJxYiIz6laAlYYBn9+UIU1q3v4MP13DqJBAJ/knPdI4
H8Zt8Wfh0AbGAFS3waqCW/KOjtKm1rYXI/QQxBLvwOMJIfaVXl1x98smI+Ea6XBe
6OUTyGnuK0C3q7oGP/41dLZe0wYenjVyDVLZL90tFlLLqhN+3z9LewpQ/fx5wiza
WSohlYxw9zyYuAdGdLiuoScAHQMUVfgI+iv0j0RcfyM1S0g4eAXkeCUwcOdB1k8p
Vdf3HIcuIYlTSYKHH2o4TR7JnCh0TlTeiHV13wEKy3wNHOysp3IV1UxSGk1jEM2q
WpDy6cqpisleKZP6AjeTk3HeHU9hzDSXLH0MlSj+T4jKQYc2CXB9JtMPD/QVacmE
nWFras1uEz4UeSRnmgNusQBlp32x+YN21gCqu82qEC6ApM1hnX7MJqpuaC4JZuxm
QSkpOaa/XwVgDzy6nbdjXW2k5w5uJPnLdr7sfhEOOEmtZKrqLy83NGat4d3+755Z
Li41JwNottHND9hDROnVTejvH5Zinb6oNepd2O4UpaIzLcWCOKgKeMsmKWuXNzDx
UMyYVyQmVQaZ1CBs8R6WDrIQucELZiQwjKqWPlBfBZDc9t76rMmZEdmY6J/Umspy
6lu2g6gLUB6FtTyQGUzmXXQi5uBVebnkBuqlOiYGE/Y4NbxuclILBOYCSYtM7n3v
YLR+CxBUu8lZlYGaGDFNX8M3sLjn5j9a7/rYtWAOj7ojaOKiA+QD25KSd/+XKzDm
hILYXvIsdMZGa+fFDAD0WshZthdwNZp9DG678tToOHu8hmErqFVNrQGW0q82kOcO
yCT06prJswM9pULoG26qkGTxSTr8HwUgItex2SAfJdmpygtdci//xkWdgAwqKgv6
KAfAo+5ZkYzNexeenvDu6PkYwJJ3YNLDsXM49Gowgkk1dYbIvFhNfFB7WVhnGtyz
2xBaO9sBhWaEbQLQsoM7dMa1wKwmf6spPYipdU+Q3oCKqjM2T0IoeJ4jZ+a2zeET
nvnNPJoV1FRzZ+v9tFfx3AZU9TPhVzDKVA1YFhEw18tczmN1h453HK79cwAoOouD
pM/jvrukywwuEEHFJFVyfEMqfAs2YpONtA2zFE8RGXYQds0j9XnMJy3YKGuZ0GM2
EaySnXsDtUN194yo4Ag86Nyrm7s8ZH7XKwT/RNe6rk+PWjxpJhXyqlCS6WPtz9Zf
bhfslYidcR8L9mhP2SYuIb6X34n0ga1RbWY2VXslXUB8Yx/93bBhURF/Vt1+bkel
OB8+n4L5jHrcLDRPSxMtLKPOyfv4XpcAK5K8MTkpN0V/6SqtdysPXTbqmZ5nm05F
ySsnJ/f1NgxhUlig8zilD0eddrui2XKwQ/sB1x/4o0RB3v1OCsei6afFhtx5rJFN
mr9s02p29YvXlxSsnwAyby6jH20cMLbQokqZNUkLI221TxT7hL220iZehRMIm0qH
n87opeN2/IQoLSga+gzY1e6dZy0QBxVK4sy8JW+FpDldx32AoUGAdaj8W1cie5bO
WN10LpWQAS3P5bSwye6HPjniL0gC6KhMGTMoj47197bdyJrucGvdHQ2G/TlAQuIO
u+teb9K+18irw7N/JkBPnfPhBf/UcmZ2aPMPy2AcGkkSkVTNvLz8BnuPgI6SqV3L
GN3zkptgJTViG32x5Drjwfy8JjIH6salj8I6Pfkv8nTkO4hEFTYtwm5c+yXS6QSA
XkVhCAbmqOUjPvIyP8AwaOd9p3qjuPSi9x9aXWOBcMMDNbwkhqOIZqzSMxFdeR4L
cbQUu7V8IYNyEYnThq0gn/5r9k/T5Wu+pyJFrmNIfj7YXNmvMMqk1wBwnPFKzN1H
UFqQToyOtOSuc8DR53DEIuTkgslQjn5kTU55e/EGee/HbuqwBq6BpCOmKbX8Ztzz
jykCdFAw8nFQV8csAN4638jOLxF86MpeMFiwxWkHBW/qxuEtm/gtBWP6W38iceAB
yUB77CDs/FYeTETd+KA5VNIk71k5yPw5XO50gm7O6Lx7MFkwWso7RTfRBWnfTY9e
ofyTFQL6PHXbytJCyanxSPJmSYvX/iuIzv0ovI6EYxriz+FOzEF4igIuP64NHtsw
WanjAUQX+13NTBBEHFfNe2Ys4TgUfj1MFTbY9flJukmGH2a9bLwU5kccVrje16qN
rSVwoQUCr5YPFuYJHm4gJ9eb4mpM+n8VoPPWbX4/Lpadzt+KTIelbj8gCKrgtlO6
b6Hr/L7shwKAFaobIUHW7qT6YwcTVin4bQ+G4usfJwsFkQvEUuNgioKuyfjLxHJp
3lHV1WmaS3M3Eggo8RJK1PeG+sBmoRxuNDm+IZ0a4Skn/+LAeyiBDwd+TgpP/ZhX
FJWv4vxNxzOMt2o1slNrbeXPZ7RuzbyYc2T3X9CXsCK4Kw2tWl7cl7ocijDZWNJ3
yaiZaKpf0AghJqBQBUqmKH6JNUGvm7nv7mYASVl0H2g4+Ul5flk3TIAU9UXqXV/q
RM/HF+5QDp47feHUCWFLCTyEbxal/7PI34pShTwbXz6mEG41cJjZR+OKPOdhMQl9
7sFxDLxu413erWNRacAFx20rc6+Iia1Np2FRz91mJ+vCmSsdozvjaySbRaJMEYh0
+53YwFV2lqbk6KpopbPJAazgDAOy4R1u7F0erf1tyMGUFAAEX+Nj4IXpx0vlAVbH
Xtd5oV4PYeX0LI5j6TXNtkTJOvBZuHsbuiZwC/aHqi6WAqUrqGi3h55O2QP2mQZT
aOhTtoyqqACvtVfzcHKXN2i2Ftl7KBZbv0z8Z5wHq3QMwk+yq35ATA3P6jBVAUvU
G2H0TAUGBr3S4gDrDLmBk+j3OPbqSg372i883mit+1mGwG2M81srk04Kpv3nli91
lwMUOUogm/iNzT8lDf/EkZFmCRcxVGUaZulKPOCpa7jZVtXTIsE5l1xgoRUZ3R0q
iJiT13VZ4tmS3GOm5JiHZdHVnG5DRfwX//A+RN/YqoZRk2D+bk+okSE2nF1X4vja
Ok+IIQQ8er1IXHyydYr8Ku8ueP3erVhnJy1TKbX0osE094WzHV4IyI8XUOxw6093
em397k7k/9hnOWU3q08SKtry8mv/k6BG6VcLrW22YXICRj5dllmAa4FOWIZpUmmJ
oLdscSk+muIgEb+7q+czvqJ/iGczvac9RPPvz582ifcUAM86tzmsBU2fN9VK4c4X
AgIOINVezYOmXE28eoXys5/WojyKONz6S0uu3Q2ehvCaT8JeHBsvQpZ3KLezEGt6
g2h6dSQe42UdphNAai70epNoEmG/lP8mD7WFgSJ50KFq7iPbBH/IwLXiBY2eOgg+
PonGuRiaCTHgebvbVGStIaawZ7Op5QbI+3TnM8lCiSIaBlsPNw/mIdqjjr8tpBuE
UThKGPObl/rFQJY3DYtG6DpIr2SspaR2NP2Ca6ZgpVdzbt9GP/FELYqSs/HaG4lw
QtwPdp7PfUuadNx/0fhMoLlf4cvdZ8dCCbvVAMYdiwcoY3cfNTryMNDp8t2t++oI
myzjn8+lE3KZid7JuFvRQRjAnlXcT7T5vZ4iwPL8o5554zPS7dGo7Ixla7wWdGYB
vECeX7m4NPcUXl9flW/3YDPx60/4Evnu+BGOPKeEGNmQ10VvmUMiPuZy4cHs+RNf
xhCzStWDnI4azNuIsFvE+mePnbTI+yAKXzR+fgdlCjF9GwjkmTBG/DnKrfp9Uk1F
c50uhy/rQb8jwfXWXHd+MDpY6bk2J5t80fI9XtFH7brS7AOe6A33Tv27IBypzRtf
p40mpQ+pzxVQ0xO/auVzGV1sQ6QWimJlPxtccVBo9ULF5yA9T66ayNkqfK5dZGZ+
WUTD2Qg5bNxYp8noE0IEaqAGJQQR3q/rIAbLPI5LNaVDA41BQ8Qzk1qZIswzTW2S
2PKKuLd0xvzrZ4T3t7+AcT7jqInaYFAA5qBRCWvDgf1pw9qr2l7h+rWc4P/KJLzU
Se8UEqgZTrqqa5g48Ybhn+7Vuu1lLDE9xOI8RhhNUuvNNteknyQ2UkWHnP6hLjvO
yswrrEqTXIFSodTWuB11YRBMolKqkwmf9NDYVKq97PajU7kkdmNPuLG/aCCED5WU
RV8ALx5HFk4BRRvxvqCxWluRBBhdCxwmTeZNnvtp/ikPJcWF9WVq+LC2O3vv6vRw
BAticMbthyaniqrsMb5RCXI6xvxgUV1JXEz+VdtCwVqyfKaXlPsq8KQXO0P4Q9bm
LQtc7+7AzH9y50G95B2dM6Xe56vm56jfhOshUzlC3kuJF8+B6Jn6rjZPstsZI+dr
izJD4RnKcaMgcIhq+rNzSBAwTMAqarrJZbqpMhpsy26mEJ5GBcPs+dwFKP462Jgc
LtQv2j5njCHbc/8GRInqUPP+1bXTR1/4iVLI/fPJIk9qTPTv2g4aygda3qnbgd2O
Tkjx7OHvTQiBPrDwyCWFcmfxHU4jKsXVHgsmeF/f/3MKCZTr6f6C1O+AC43xoEi5
5gQqRXw8Qb6e09jM8Qp1311eDJzjT+XaXxnib5jHT+sfm523iKSNTZyih2/gpAdE
Y/PyIWvpuwIx6DfLjXTsUq/CxIDuZ9hcykWzx1pDtx5LseQ78c7FeGQ4TGLK8Zwj
ovWXyZEs9Hui/jkM7QSgEcwvz12glEF5Yufa2yF5aGB1L2RgFuLzBrkNOdLBI9eU
fVH0nhKqBTYu6MPDjQ6apA56Q4ZiFtAsytv2ELWQzWF935rpR0vXHRx2QcVgwQ6x
96BIXAgrFlA2TeTaPDUmerJUz+KherVhxs/OQ7unPdNe7plppQ4z9ytS/fwyl1QX
PdicQMc5tEFngSuA8aWQ+DWQmy/2eKGn+u4bzpVTwDO2GBJbuJslSKlf/kNBUVJI
W+RsTbTMbRyr+xqIAOWPDHsJflBdrPzlzk+1ygpPtfrICGwSF6ghQ9+HYmdWfKve
BS9RGYzx7VFAuXzfqhwwlvVXhoiuLV/yvde/hecq9E/3noAy8VOuKFXb4BDhpuqk
dWzSNtJyTygt48W+CeAduHxkboBcMareKrhMOlT0jL8/SAyGVVXELRqZ/gf4ySjs
2y0vctMvW1lvx8ZaN7MGijpyNfcRbTC8VvTG7Zs8lvbpZJ39rIVIBjj1SGAC3hS7
Tn/MlYJGPEFhoheSOvM8DkD/YGxJNQ1CVJn5htXmWeCDrOGb0mM9q9CKbfzBxqGS
OW8VNk3GfpY6bTwEisMIx/CyRYvlhhQFpt5z9RIeL71fPS/Duupy2LEkvqJ5+Sx6
1sFumq5/a4m63o9hD8aeA4fI6o29gWJM/z/RoSbvgV0HYZ8bytzTSnvZZKcuClvF
f8jTLKGMe5tj8yQwXwut6Gd9fTna7fdPd6lPcPO+CyqtgSDEMlcI8OC87iev/ExC
ezFdNGW/HxqJ8BMp2MWUwBMRpQw/p6Y0acH5+G7PZKD8Bvv3v5uo9H6V/R3t07Vx
un0Z3xyMxYIOMdCdhQiqfJgyI3FEBq2cScoDrYgTFfQyM/mGqq2ezn9uq4qi5nN3
GQYFIriCU6WeoasAYxBUmVCaBBV4BsOkMsp+9mY494kPJuwt8iLPQpx4P6L+dh2k
+7jPh6oZ60TLURk7NNuAiiRn2X7EDQqzlw8ioz6GRlGUuKDqG0qFHq6faNxZdiy1
sfLaeLN0XO3dR3rOuaj13I02f+J544diUvNgLtTsCT2mhwP48aklWqbx9MA62BV6
cFaX+0Sl9HL78qfyUQLWi43vIUqbLaY9JEOf/UBjZIBnQhUSi1YWKtCYNo49taTp
sc3jm3UtLJxdb+x3SAfYtgYCGRdqEJhshRz+PBvxnhgCfN5I/KrA/+bqMcWSF9ne
8vWg/GTuZwoE+QzrfsOUNDsbAWP+lFoe8RHErKXrADMtdIMgwQOz1cKmewsZ95Tn
fZacNLtkLe/45gEldHYyNFHdClLdVsM0miapc/Hx72oCjLRUySRXXHuaPQtjuLd3
Xn9Re8JkfPf3PJyAgdM7gnrVqKl+8YTVc8K4HZvY7cy8O2DDP46CILJKX5T6O/Bl
rDKL3dIECIQYYrHKNw2cKMQC5ZLFdIcaoPxyGVkSgTUJuTej7TEDQjuNC6COgx1G
vGZHrsjBqJpQeEFEOQxOGNLnH1zWcj+LiBbDOzMB5VjabvdZf0sLhKGOSqe7Hiz3
8DkG8KObI4yejKTk0dlHmwGiQCdqDI2YcJ0hn2q35Z0oOWZzhjM5KO9SZyLbfM+J
ftRREuDxDtLN6l6BQAvORrUpBlJLfQX0AZxRy18ynxVH0V3wRTbASxfc+mcJmSeA
4KaxPmgl9Nyt5fhL3HNMju+0REDGXk+g0TIzPHnixorhvlijDDOS1bqGQXpp8eBO
R98633syFRFGoqPLhg1N6BW3GUqcRwzSkJCPlO3Wy+EVE/lYtTPgyiDlm5qR1hqn
Q4ny3Pt4d4Vzo86xBTJ7eTsCCXhhAZPz+W37k+bGksQWgFDg2IF8MyIGBsN8YagT
x7TR/IvJuHd17Wjuim6t+Zs6L3eIZVg4VMYO3x1bsWydFHWDPu9CW6lVMDyFzLHc
9+0+oR6dfAarsaorFed7y+xlMtsiaRsCrgYXREKajRqKAr5u0ok9N/+SHkqOm0IJ
ywSz7Sa+v1CcVT9eJNN8oujqY099eL6gRiZUuGLwNb5s9QgzYaQlSOrRkKmhu3JK
TRoby6C/svIqucGYEXMK53WKnA45tpiJs9rYYPUU0y0IraMonLJTmKJGUUH0Tt+V
QBea888FKz5w/Yzv89HgXj5Xy5Kf1sdGviFEScw72g6FASOAh/NigrTCMXb4Cz9i
WGOhQg7b5akVyrjKa6Xq2YsreU1hjA3YWrS2BQSDYKIvRNfEm1B0B7yFtNKdPObj
5bj8elxuYeGip1rm4eAxBVh6H1187zUaKtdee0DwY0eAwSoRjpsGPyDPxiNteLSQ
UcVKb3PUGXG2VXQBwvDzmzmufKmGL05vlYAgjDjMqTB8DahuZJC4w+B3FITq70iK
51JTSJN3g/0/UKqL5ZokvSUIIbksz3KPRijCkVWKmXfMjja/ka9rsSgkuYZVpnYW
MrYzy+Oddoc5ogJzgpMU6swHLpeiqqapIKuoLS5t0ug09a4GC+GPtzvH0pa9qEsP
RF06NX+tbB8zGYg24aBMQGF45mJ4yvkh71P3AlI75OJ91aklXXDstgWMtcsMFZjk
EaN2G4mUoy1u5nB9ty32VGkoERLq1sMtEE56KolX7iD7r/VSaEsfepmTpLW77jov
0lrXbgQG+cvMiI7YE/vMF92Gm3Bp+VQH4Ag7q9Qf585FQGAQrO8IJFOGvcknIWDz
oU9XqW/LjDps5XMWjiY7/w848wr0TlcgqVzMSdb2VW5xm+Eim6PQwzy+kxOX/+ix
XiC831Cevm292pOrhae8VfYx6eMBO7z9n6De1At1DRGnBPNyBlA0adU/rCG/m88K
bgnQcEojCHJEsxzubZe7SznLJhhirn0678zPOIv7VzmG9GZoYBFpp1goIvcJ+Cj2
BxJvag8TybaboPd8rj8hNU6mhyaHOrVMTUSJ4LIxXKH1MeSlwVu7rzlLc9yHDdXa
ObwMTPUtgwHSSv2+iVGXlBL76JNA6oSLO5J3uwK+h516JnLwLqa9PX0g+n8ZIlAz
/zAjtgJ1MadUhMDCiXWKmR99iq1DWZswbIe5llME92OeC1XpawEZjwvmwZN4OIt3
3ytBv75cjQXXmULrXNFtkO+DZ74+n5KmdBIwciztvu9OBJuPJylCN+/m6TMG3FCR
KJC1PBeQLWm/xTzdXDSRlBnZaFPjO/3hNSTxxu3D4Ok9LGVZKY2nrZYfyHVLA51d
ph5RKxw29lVbgKYDm0YWsAFDWv9nfdzagLZcc0HcIeCixf62rq+QxIf82mVU6FFi
B+qaidnVRltpJmLerEy94RW6uDDkHh4hkAM8wx2ZCWvJbS7KfdvybHwa7tITsf57
xCL6JP15MY4qR1+VimbRO56TuZdyCIezlccnEk6kGqcWBcSsW6FgVaGxvCl3TV8i
P26M/s3rTbLNg2OpvUgIRlL4fq4Mxr/oVCTm1dNaMv5TNCQniCUp3kXiyIYiur3x
D1wfRcTBI/4HWIhA/FHLEVzsPkEgApBBSHitq64KtGuDasBlyPJ8EuDaxBuVON7b
T7/7vksTSuEpVSYwshXwQvMzP3VkD/SOkV05edDd8RtrkvMPjpi6OnvxuwOoBJy2
Ub0UnicTJT4+oqYMFSWZ7qh7i/Y8NeWszeHGD5Ugg4U8oMMEkB+IT37wxQ6ut1rf
w3LXXugNBbLp7E7Vnoy9YxYBrvwMA2ADS+OvYfW0jC4BSN2dmASPwCWcSMYfaLGM
gGWedOdeYiRIMYBi3W7yUe87enaOxNM3LzPa+nAdXJSNurYEFwlNBOmZ25VC713V
3ez3UmNouRoNovnQPwrllxXtmIfRWeg1OcFL9a5m49OdZGXzm7Ej66x91MPaegOn
eSAdEXrsYU9gH+XiTy87IGlUTOhilkv8HZ+Pwyynir0ySU4cUyuDk34VK/4CwL+1
vp8+UVPifo+sBd76ma13O4uc94/8l8QcV/oW4SN8f3ndoKrT596BgAa++o5Su+q7
/lFROEQR8jv/8Oxrgi8Nud4hYAKeRrhuMMf9jlZrgtVT6+2hwqduDQMoktRC7XpF
ua9eBqhauhhIdA3B5pfrab79YAjHDs103XY+LQYsf2JLgpGkODvh6dbOI8ywDPdr
nRlntlc/B+uOm4QUbMmm8Xxq36aoJicloX/fiTWV5iU+YKco8mnkhFTaGAXavelZ
kDyHrKmcXGFMYrAWzV9QRJ10zFonO9pACdSNPQKqeleX/aakhZ1RziShAdjR3ial
d/MOiacGnqla7wFZxmxcQIQ40Rsmue+PoJUv9+Ev/+S0HtufxK4SbrbLz83YkL+R
MS/+W1eNY6ntDSK+hkuHAuI5x6VNvC4Cy2GdTpKlHVst61pQ6/qLmmEI+fiJvvOs
Xg4UEmDpWeh3Bv+XSKZAjtEtsLrZ4P8FaMR9/eAOl8e52lLbrHBRGU/2LEkAjF+Z
a+sAiprFhvnOb/OaKAg3d7kpD3rKB07weEAJuEek3dz32Q+SZsRtgB4H3AtIJOba
jpv8+vzJTCnBcmpULtrcaPdzMcauOggaxonPMHu6RIZeScu6LCMtwOMguhwGvIvW
ckZlv6XO+kHfVWi49N27CXy+7tDasppfCd5GWWFyd0YZsNWIrJkBMZWqNmA/T/+k
VghLpy0XvYxmJ6veqxqV4K3AEdLCNabhqYuD2JcUqiL5FswPDp6ahWisyDIsR1iY
UGg2rY/VcJMY6vCCe/4OK2cNNYnBDfazL+f2+JL715jHgEmVs4owUcgCQbX3PpYc
Vj/5Ep/60qyXYX6R56iLKZAnTB1bXpJtw/ZWuwcdP4KLFISOouAkPByI0Gvg31gT
ahux2QkgiWIr+aiA1SjRlmKZrW4VcWNjdGVoqtR3hM+iRulXvPBXi6/KDPij7YpO
8UiEW9FTFgleaNGpulrG794KmbpVGPqwOl3d/+KETN2QXKHQ0VTOleAjbIv1oBCN
mHnyRbEphdnkOpwUcZCVjmAq67YtbKrEta/m2vHVXoLm2u/tLSQ4zc2N3W6Pn4ly
3dyBx67fHMiR1/x+7ocsPWCGR/LHG7nAcxcZ7Cz/ku6dXlRDY4/6eChAwJbTpq7A
R/ja3uQvyGT9FtqYLAwFwpvHmTLAH2MabUniE7Z1HrbGLiKFjUcnVFpg6l1nPraU
DaYS9lhZF0dE0DQtfzsLx6exP1Djb9kTaGuk+Hsmz3ZqA4Mfz72WzYhHs/5RtoLy
N9/c7dHXmkEImHC5ruaJ9z6wHurJeopjeSrloUb4wX/TP8XSwg7tEeJq3wzGexcS
1emzNXIwSLk0RO3WXTpFP3azqz/aBH9fieJhb4gJERppT+vi4RPWcz/s7/H2nf4p
3YVV5D4chZhcPTd4Kc7J30Nc/h5PcRihgnNDcuVcUOZpACVi9k8lFn1ZQl0fKYUV
sJ9fiVh7k2dCfdt9Id7Ni01eNiE0txgNDRjSzAPneMpyBUl/8tU3KupynAHbW7Jh
GwZmyqyF4+L0m7piTrHcdl+46RgSM9LN3V7e/71mx3RmZmnjAhKKEe4LQ29IxOcb
kCEldlkaf1RLGDtnUguWd1EzNuGg4H4Ms3liYn607J1Y7rXJEmfYy6K3o9vsgszv
UCMh9A1MNFSjh+XNeEXDQAm4zpSv0ufSbcvdFyD2AjUiy7lPzlG2Am103w9QY4HP
pDumcy4GYCIi5YhSeXBEYD1Dq9J0zcQ8fmKo2LH9WfuNTxHKdFriRN5NUm9mIGtb
Rl4XP+iJLJHPWxgYaMn+GGeYD2uXm1eO2qRi26STd2yZjCg1fkSfvgbUQ42fW2VH
Emo7cZwbGBlxfbPpGuE2NU0ypS41UJiAxT5cMfU++lqKw6cbd1fFyc9uhrR9Fdm9
O9sESJNlEMGt1lUrxUNsL68gVIUa6F9Vl6Ss7AMuzfLta+yYyjgZcit07MXuRmGR
7QXCH4tjNx+Q2pgwppczreu3DWCaFZpkKzCuc0jwXUgavzo5VCmf4UfPMqZLb+hR
7SJb7UhboSyE8x4rAp9MYtymPuQbFC9CTTxPsm4WLuoRC5yKIbfLBdagHutu3cd9
yqY+tk1COn/BY9YuXj2zf7vgs885NanrzsYTg2I1ZPKsIfaJ5GcnKdcUlh+yRvUz
wYviEGcnmixpZmPemxqDOhThlP8L0Kp3uHwlEWETbbSLYD7CcqP3ijvnIlDW1RVd
rT5IFSl3fIQ//GpQ+pyfyFYnEICyuz8bjRkDMS4kH7De9B85gDKBB86u+s2mAJu6
VwYBMMck/+r8X1tv2rt7aSMqNz5oxhu2LRY0CiGqm4b9EcdvvX654SX/K/AI4bhb
1q1eFx8GkyuNNM1aS2Lpr86nRc+7nPZB22Ai9mgoSzi0detOLQyus8TiRQD4HKqX
4Q9rVfNsF2nz+hskxgdAEDxjm3lJUKB6qMRqlBgxwbytWieR0paKYuTSthbTKv57
qYtgzK4HrMdSPQ7FfD4srMJNu2IIco2axQp7urKxMwpPdKz/e56g/kVULQ7M0g8I
cpuqmKdMltanSB7nBaocJFTcjXspZQZNpzNhsihv1iGSNH0qD6X5KtsMyQYBFM/b
FdAYFlG4sO4ZgExJLoipsH4Ka0UZR8sR+GWg9s7eAomEvvSGEnNvet7apy9rvtsU
TkrXkv7X4wJdn98gtoSfus4wdBw3QSQzwhHY8HrYhaqRPglxLUNQ/xLbiQVh5rUX
Od2VOTCKls78p96ai/PwSrfRm0YGwYv4ogYVvoRVoOjm786tVNV+/q6Nz3H80vMV
Erzcm1Y4UP2igsYJ7VIrBMJHvfiJeqzhNrwZxqVZLBDuTHXN37iST1XXLrwHKvNi
SG/oxIYKMr36aFtDe7iSLeS2RBlehzYgiyPPLj5PgGHVdy4TF+m09iw4SF169+I/
W9qMgCEXha96qgK6ZUYeN7b+68Xnffy8ydqhPpqiD2O6Xhz8iPdgzA84VYcwxqC+
ded2VT0uR2L6qoNb93+Kq/N8VWdltF6yZcUfVlLMhwepCJAha+1z2tbL54Vti8h7
UQuOELWtWvexmRnhR+t7K8vHfYdEPtmdCfVZqf5E4hFbOTR1LKNnpiy/X15Et6dy
FwKE/1AxiH5tMjZtGZk0jrtjaj/bnujdqdaUGbmXzv4/PH1XmCklAzzU3hYKCgYR
qPUf0GIXCM8kq1HmEDHimOdtW2uY5b1mdO5yKWEooRmUZVVQ7qr73SJqTcQ8Lhkh
ihVT49rG9vmXZ1albPUSWqIwKLFIn1fYiKP4qvK/M50XfHo1zYZYuxSRT4L5fOhH
UhTmvoasplWFm5zEnu4JeB3NabL37iZWXq8a7/maiHaf6kxbJQQuxFpofHJiU3A1
c0KDKY4tmuvq2Nlls9UU3qDQWWsW99go9LpGiX1FEYGN3J1XNjUmWFa5GMFDvY03
7GGMKeZOz+tfy+27QwvqQsrp6WQA14nDfQZ9Vpjk3/5r0qL7pn/b8lTyNlmuoffu
5eI3yi7VLhxJC+KaCjs36UdlWfDe7RxJMk1+X3FoSJ+fZKy9RKkuTMwtJeoq5M+5
Oad3tI7upuHdY1z6p6wfuJveYkWFWNV6zqVkM4J5hYj0T/BeuiIcHplVCliT7D5p
JYJZWmwbptr+5qqHECfnLHMa987osKKh8w4zKK0mjOikjWIEPd3S/HQaWo0f+bF9
kUMCo+rMy6XWsF2XtQcIvVUH1yoVvnDIUA7LcU9qZEhKFnIbhX5SkgHS3znkvcbn
RZ0excKt0apFVsL9xvDES4jt/6h14reyT88aI23zx57vrnUYytbHM5ePKqc7yiKb
k5RwD38/XB337qZEwaMA1Q2T/tgpW+AbWFZYatsR/k2vvel4boZGzLDjRc2SYam8
q3rRvfqwbzRWpgZoCly797TNyL91i5MoJqBTywMHSCC/3elNXRiFaRLlLG0aifft
wEW04qnHOPd7zSoRt1Isj7D5NMet2dmiqSOnjjxBd6GsP4haKFz844J7apN+mFyO
AKPU4EL1hKUKaswlUg80h0xBA1cdJVDD0xCTtxxHLP68I2yCa9w5bvP/5Lj2RD8c
fgMQkXyaxNlK4+LC4rOoF//jMQif5cCseDsmCoRV435mH+2IjbDibNUgTkfIls6n
RRWWMAUGzpex1qxufrJKGxwJWAJeTRNaffRV2RCooV4FnJIF+YtN6D40LFY5f5Xs
2JkJ8Zz/Jhrw4RVxuuoCtR5vBxlJftmOkLj5OTGcAEdPMYS8WyOEtbwbziinn4CS
cCXYdS+CFFetPq9VwphPBOHj5/AjzCNrH7syIKQwcGK34rG1W9sHd1YxZojcaaae
X5oAnExba2o5KgjbkaGZJIqrqjj+wNmmz7HMiUiGANS8s1nmvK5G6WhvAanz0ITK
/KTl5R6yEmEW4J6ZyRRGgohTHptbfebECq/OubJp6qp9B8BtxvUzfgy26lwWo4N1
GH0NDZXVInrU6roZSVKvpiBxfBeYpj5koQWgJ6ebV6ooSdTiaDQOWiEN7WjEXjSz
+jtZFKe4kszC4gqpoD8jhwMF7xtBVSFbeO3+BxGr1D0a7pP+lc8GF4x/RjSNBkpt
UUAgHOrkPVV26dyMD5aJLaWrz54SPDneSqVgKTv3Qou9wMra6fK2XnZlof/18UfC
ZZkkEOD09l4AzveQUHirGNBpc/8A11nOAj91WGcwCuRBy/DN2E3SKXtjOyHXVk8u
6VXRqP6xH04zeFBzi16xcKI1uiXqxUWaHRoIpsBlJ931OvLedN5hxt54ss7Ic3NS
mZTYG6LPsTI4t3zHCOhz6qEXXcQNgwL5nv9Yb9H7MSxLzK5a55GdSBBSrpIQbd2/
7yjdahlOqEsZBB7W28y0FxDHHhqntvBvyoLU/zwf2bYy2lCQkktVWZNyK/ZT9Tk4
fphop6aPfMHUTpoImryjnAwY96ftOa3Akad9jjnO6O0Ham/O7SgIMEWUEhIJmZqR
bjbYRfmXqUHOzvqZgtW3G9nRXA+tqrPqws81pS7C8TG+Swm1wo3G8ZecW62CAnQX
fIgLDjqbR1NmuRvZiSlkrfv97PF4SVL9DiJAr82Rc9HQ0BxwlONdPt3VQGk9HEKm
BNxHi1vMWIvFIrptPhxG5iVrccpLPGHa/c/CtgEZdm/Q/1sxXjc7zwynWJgoC7eu
oX1tmPzmmML3hCLFdOD73AWhQQX0bswXqLgmbVBDLchOcWpeITri2+9ubRvJVHm7
Q6nDDf4kew8T/7LFMZmcLtXvWLETZtXrN+Yqc2bIpoR6Jf2KmHYfhC22NkR1CAci
m7OpCNlvPjBrQp+hXsIcTDacqEQf+XoJHysXdJ7oP/VlIotvwXSlNBvqOn5UNU60
upZwSpAUK2EtuU1O9J9bzMbWe159nqM4Px8KSo9c7AjM2TXv47RA6QJEz+MEBFM4
E4uZ19dB/4ycFrlSX4sO7UZKWTq31JW6wmHCNItGhmuXpCtf9EA6oap0G2OJ63Ep
G9ZSJl2XvF7ATEeP/U//ZSBVrGGxvvveqAmgKZYkk8PovPHEFgVC5VpDVXbXiFPT
m19nXcd6UzRwn4mh+ptw19CRDO93Tvuzdt+mJQb5KH4N3DmKQaiZJ94HyNLtzyvL
SrNcV9weLn9MC4Gh6B375lnRubMXioyVYlJ/58bLH9Guy2CM/m3dHmLtCc40QeEK
V5b04vhcOi1cZSdLMZJFm5GC7ewNb4aQcUK1IAxoegukjVCa81Gw7jxuF8g0p11c
Wwsev83Wf74/llTMqPT2BuLrsRUwl7afvX6znEO2BPw2pIUc68RYNgDEp+QpkLlH
yCHsLLVw2HHOIOag8rr2cOGkJlkMz9lBD0H9GFqa6mU2vWZUILfSRr8uopSPJWIw
JqQBEgx91+4D/+pX/LuCsMEsaWQKExONkJdli8D+yehy6BBheWxmQ4UH5ilQvFUr
lqM1/nu7/1+mSZT3Ov9UjWCFfhgWM1wqhOmlJiBLqNRkfqRZwPC+5vDmrtD1edFY
3VuJpnp1E9PYcW2HQU/eCZbUg+mB9xboUcZZWLoE6q0X0O2ZxjPqfdDq3EQ9vldN
3UoaOvOvat5KyZaC2URJHYsm9yg1pCc+Z2qzLWJNn+FFYmbU3F2LhqQvEWNPlT8V
8zFraO2ULggVS0JdUZsKdob4yUHs52M3Mqqb1mpY2AyFo6Baym2OXPhARoobDcty
coBcH7Z8+512jhireJLjFVUFALXAzjUFD/IAWIxuIhlk9i5mRVuFxDn6RcJGgfs8
DzFQgvFeubv1GBT1PCXnKL4QRQHlO4F3JoXg/cmZG3DjTTixQSCwAlZmDJ1jQL61
PzC+LvZIEa1lhOiN4bpW1fo3N30YJ/T9gCojQyJczm6ccgEzv43jsvdWFko7eZR9
iZng99j1BGwE3pw0Nfou2oZXlHFGDyV7yCh2QNj+5rE+AxE49QD/Jsb0NO5sg+0I
kipF20ScbulGV2xFD/9v2ehGtWW8p5s2xYSv6cDURv0ojTkQZhYZG24ja7vFHKQ7
sPasM9OBwj+7HasuC6hxz0nu7joH1XUqcCsAUUPjCEjH+kXeCSbYMU1nUy8Coldp
PJHD1oeZJh61xFHTq0Bgxuzw6p7LYcWJRx2pKIbQF+/HQXEze75AXhnty2LVb6FR
mlpHyTV3oN3xbrcz3FW6YsCu2ZwCgP5ddYyCp+BalZJ5C9rfVAcVCAT2G3KyhYPX
lQRuN4bYUPREjaAaulC+2/N+zytTlKrNPuteHGFDFx0KxCOpnaIBYWyHBeRk2Y8y
rJacqrBZFrv0HaUteVMZypt1YLgrUDSAhp+r++/ukZWQh9VJeQ5Jd23UW7E2KP0R
SrAbNQ4nHGGpOBlZcSF5SlRgg9heS5zDujjluokO1pvdOCG/8hcMqNsRSEwNa+Er
mNIeDVWBbfDMjI8G0N7ZexUiAky+qAZXWmN52xZcF6eDHRfVxn67TmGmkqdidrT3
xFvmnLIYysmej7XVtsv21uEZX4ETSgZp0fdnFslss79Kgeoeea1Kbzbo+6f2aLMv
QqpVUNTJdxCMWDX+o1AUpndNfoQoyz4jmw+oc+WZWPtVZtjTFeAsWQJOr1V0xR3h
LYhfacE+rWz00DahgfrbIjKho36pQZ3abb3iE2wNuEpXUkFYz27y/pn+UMahRLJ1
SelkJQzQ6+iFIDZQ1GJ+0+3PvkPNulcIKThDNOOK+3Ps1b3mwkgG+cxjvYuNrBup
O0+NaMfqibsjwpsSaxYN3B0J0PYV9IeD/xEPUZXtzFU9bdS5qY3Y9VPHn8urgyj+
Mw64dGXD/+p7ZceLUIzbZaWULUCBc21JuKvjxnKJYbZVGn0s9bmWc5HpK682G4on
pszvhz0rBIsOGHLFvlOzfJZCFVrQieT++3R0bI7b/AY4aPhdZCEcSMnwYO+kj8I7
gVdXvscvs4e5c8xMK82LTPvLb9g4xmsiKaBcWxSLZ7fYa+I37wdScSOtbRBxyYYv
PdSIRfsv27r8Sil4Dn+7p0TTHm/kOQT20kmfkUHO+0XS9Z0L1oSbQ2n+BvF7sLaR
88FopROORuWrem4Qk4WzHRiIC/A+3EgVLlB6meDhCHiUOodrg1BT0zWvq30vA+eb
xn4D5WaeHMjPvV/0KSlByrOsVPq6h5pSCNgW8grefHYXvNuA8Oj5BTGDOLYiwcha
RB3zWk6TX78q/cAHjNZ9mHl3Y5YjA8QTnEIEputawVAm5FYZ6BuRyT2xEjtXdf0Z
68IWm3pdrBvAggWyzVbts1kXZyhaKorR7jr+8LENKkmkmvezH3X2bVUypDiBnjNH
kY+DMUVlmyM/xsE0WxXD4hx4rD2vIM+D1FlJEA4u/UQk9U1UBZFjj8jfxRRVCD9u
eSGwNnOnWCFisoOquGmrntwOaGbKhgsOYzskrm7rehIIag0ZTfXVKnR1VtwsvhW1
EltSPrKEoWYlTNvhIu9Ytn0KgPiKDBh+A15qPGPKDm707tk/zlEegliN9T8Y9Spf
Y4PK+OCq8uURTknczeudPjbndYo/l00GneJnwSZUDZYHV0k6iy8JEHgfcz16m7aH
eHhbpbRnCd2VQJFaQoL6oniGbD97Gt4zU8aIZFcosCK0UeCU0E7qOFnFY0GtDKSw
0SYyCNp6UvyNXzNmxF+1Qt5Dxr1Q8zfMx29S2kd7tGidW3PS2LOLwPWkP1pZLNzr
Y51jgkOTKzg4/THRPwQDHxMW0qcPrgou6VU8iE1eut3bTl2YN/iKPEYf3TCGYrr/
IA8d5lSOst7HHHmfIWbIbq5qYHkihS9oZfS0xsyuobwGdJ/gQZ9Ll8FcZ1L1Y1Xf
fparZzXoJ4K60FoKI34zfZg6aI+efvS5rGq0X2DigbzNIgRC8juPWB4DuUXUSeQZ
6PZOc4aD4H4piwWhR5Y5nFCwAG2p7IPc6DVItXWNHyYFeaCj9onUBmD1F6n+8OAC
l8cplagKyCvBy1hw8M1s3ObHTVtybjA3s1VULZxhdEVy1yt4MKGNUtLuDkipBdn6
JkUU7gcGEJKO8d0q/KzLVOZ3Sj8n45aY7r/5v4KsEiZcIZXqTCo2UexJgNDbZcfo
4ydNmd4Okn+mg4+8QnrI5yjCFOMvehWVDSAt4QKbaS6e5hvlkW4xn6i1bIYX3iWU
8VSI5b9wlVhfMrFfa0PzSOVmP4WDCAsGn9A8XQtdo9l4wZzFfgGC8WaInQazJovO
1OP7rn48I/ATP9qjdBroRXvAJ91Du5uBmqtWwL1cHT0j0JrsNVJ958uzbYGwnCWs
zoDHzzAU/l14JNhoMZ6DKRutFzIMYCrsUM/BrfDPSgwPL3qFuP1ai1Iejvev5yC5
9ruPgDsDH+QMiY0jeu6vehGWcBbo7/cgAsip92YZ4SYIR3ugwfWqMSrwb3d1zJFO
oyniBdF9v9mSGro/KDPILji69CJFlGJU0DZI6ZC/vLwNc7onxx8nvG7n39/wkHSZ
5sjm6KxwSwW1rQYqR8MgOSA45UYnWgv6nreMt7bs1oyx24Yp6yscGdjH5Jz0NUmD
Nxa+XFvIi1TFOfLhnLq67Ck7QFhleXBksIHCnGW8aUAvrh9JeIsEQRRBABaFVxMc
kV3q0jx8yffdnveWw9sf9R6rplw3vZRKPb5Fh0/8Qn7zui9FispOvnN4+iditlk+
1drGxnV66XulpvvNgJRQdYFzSLlACa31proenXtga6X9y9eKASHnrvAziS9C7XKr
y7c1sIge8zrMNog3NF8hBre21h4Cc83vwkibB09xj5pFJPKWKy8/kS4H6+2Q1kE9
1DEjyqtP5wr3pjSfx9nD/bcwP4JNAWYILW+1AKyiBAU7Fhd9hPUqqQm0/Q8cSErv
BcC3doiEY9xN67Jm2e1cQUTtlXTI0dum9TE6QoownfngYVFKRM3rYLg0NL0xvx59
hfRhBdyykxKIQkYfwft1uMi/mzA3XqHW5ATKDLBLBzHiyCTQDAIZzE5+Keh1ml7B
14MOv/zM/J4k/IzFMXP93hzSZ6+vu7ttbChHTUSaYFlqpDAz3Nwq6bgIDPIcG59w
bf67Dd7aLyZQQb/5gFpc6f+V4M2bFRoK5gR7ezbkbNLAjBRmbBXwUqbi/uJY9bxg
XckNhIAnxOXn0ZPRBmzASomc+Yz7IetgIZTK1O0mcDBzErZoP/CrycYrA1//QJDk
68I0NtHkIBkdtpjwr2odfi32s9HvJscHSfrAfOUjG+yytV5vLy/MAHX9f55LpcVA
b1bbI1OPRyi9xHxWXDPPuAMHf4092o8awJ2WlHzFB6ix0U8wqPs6vmb045PGQYNM
UuIDIfXLTW1zAxwoz3uw5eDLFxmRvI+0aIlCg7h11fGg6F3c2ijsBP6F4z3UznbX
hFBGv5bFKtzju7aGyy9X0Pi4QF56A6Ns/w7UTzMnyjbOPuh8iwVMQcqtFjna8imL
cr1mJzoa+F2xGBFyy2/4Cyotbyfe9mXLYv9YftAQUINf3TUVE2SxOTvQb591hbwJ
y3W3BD1Btf2jH7/3Jx44E/t1IMLA3fQq7PpmZzpSMZKyLk3gxrnB4Zq/aDRRIwKz
+kH1gwo33IZQScg3MGLe9NJV4E4h+gl+Yeww57RbyBj/ZlJ1d1Lv/vMmMTyT7N7H
hYvAEjTTMK8b8zDLmWaVGPEch7xo05v8vATae20G2gJfmRULULfbZZLwDPDNm2rr
CewqgZaB9jsb0DbJ+Kh/tLI020sLmjWIuJfS5ZTnjt4OuCdcR2xmmW/rt5RTn9Ln
1bYzyj92L6q5rOvZYbO7At9lAgqfFiKW7RIOn2FPaIGMMoyzlxz+qYpje4STGrnZ
GNGGZxtKQoObqNDb5zq3sesFTGtsUhP/Be69T/Fe75ooUNPnWJpvXHDpNVYv8ACZ
GYwnI+zKLeF+kHokUAfkHy0ofRAZVpntFGJw1uhRddKCCwKTcR/Dwi+aLjR2Nye5
aG9vKSP96iRla8S0oNA5OkYCB5vDPGgoJbFnC/59yplnf4u7zZILksYL7vkOfLsu
0W9qANF7ULZx+Z5kJ0DFYR44K3CEdD4LTiqVYnCy1gfss5qYWALSClBCl+Vx9SEJ
DLpFQEWjWIQlfty8l4qexlhgR27H3neTMh3wSj1wVjD5GmAMcLeO+omKJKGU9Eni
8pA/yAKqR4sqRKNC5x1/kKtCR1upM1OlFEIRDokMUMEEwH924lU4tikPdZbAJbmL
osDlFO8pYweLuMbG2z8SU2HphDXXg56eJbcWL9vobiAE8FTvGUAHYo3xzhZ3bUZm
UzWZqE/CoXMA5whdHUD/LiEXQboENIu5SVRjJcXEyYyBrl20bD6TeqNHszgODvst
sB+ZGnpVVXUgsxfhuUzLcIrMhvhzgjqMTWtRbMrSvNWILP4AJRRNTIxlmlNIfWPA
BfFvrMMJxpHH/9pJRYHVOPo77ZUWXwC1qweK4DBeSI0u4VrHUYbCV6VxO4BZQNAe
yTD/BkbGdydb6B9pt9j3O5njlRB4ltSNcS4i8/XdkCcSt+QKVFwTmKP3SdZNCZTv
JiCDeOgYzFW2PH67v2/+XlqopBbxgCR19Qz4rwxJAGPM2lf43te0zmdihnAHSHS6
WnxROQt3q9zUOjguoDm+WsHSuSsiW66urUoNCqAnI5DNCjRe3QJnJVYfVTr/ZEXQ
KhLTYdeU9JQe2BgSriZx+A6x+4NEfrTePoVAGz0fgABDhBOh7AAzJrmLRxYgT7pW
J012Mk1bq83lQZ8BHHvxeKoWpNWrsZ6C/GW5hHfrNDBctnOsjSC4obeDRslc5jDK
EV4KUpeI7mVDzQO3fslKlLfMgHpHpW0QlP1CV+4rtHwlYDySXAtX6vlxefI9Y9Hq
iDOfgpXyh6P1nvjN/zBJSckjssn/Qg0aHq0r59xYB7xuExMIUikiG0zAPgtU9tr8
OFPWR8WuaoCPVVw/JJUWXxxbm7ZeagUUUwNjlHCi98xbGyDO2y4w6L+hig26lB3G
ZxDdovyl64qM6SkAezsoH3V9DAeClMoGfCkcGyfG4WRD6AzbxMcvusYFCESvn/Xr
RAMe5vjZf+8/AYs1oB3UgVg90MHfn8K8jgGem4y6PNW5AmZ2p7dISDx/s9U0EkCt
n2/8fDlB8s/w8Zqeg+lqnO/hCgcnAVBFQi2ONEGbGG9oULquTaqdP9/h197ADV/5
t4HkwPUIscB61w7sZlDBiLrNvR62UdDqKw5DUkiv+hi9lB4tIZyyXYF3pQ25iIUP
ejHoGwqz+DjgEaDpIudhTS6ScEmBjuDypd72iVUOKIMp0EcNyK/WZsvsRHKOIuyd
harKsEjudjkofR6ZlQLj7RjW+RVy3Dl4VfN1NNBAqHBdK8jE7GEYjdiAeyN6lDya
qbCsx+hEHsOHg9XXXgxj+tVu8NPdmqFXXtvdoQPbxJx4B+4Qq2+mJM54QpV6u7fh
+FOfAaC0CbJrl4WAY0OiYSewe04mty/43U1R6qVK5CPTA874Ds+w3PQ4K7pkw62A
VpKDM8BE+/06eZNbV6GiDY1Sn2odHcgKL/KkV0ferMVk7Vx6Fw2B4CxRlMdwYrSo
ONwV/WcjSDGitNb95DLhsczJDYsfeEbz6mve7KxUC0N1LBX4XYaeTC67Npx50s1i
/4NqAP44g7ribAi6yVyk/3L5DGnZrNHSAHSvk/QvU82YZoHC+7te+YQ4QJhsV69y
9GxMLNn2A4cFdjx8Kdf0a3c9s3wiKz8rA2qH8Rt+PZz0P8jvevQEuxhshYA8kVGM
4JSF+KmdFcKaeMQ1OraZo9x3Ezu7YWwp3JsXP6AC0E6xd5TiA9ihhVNKAOVcfCde
21GrvU/3kmmsyFgEDaYZehWY4uun6GOjNfZxKmZWZI7RLoHSlvnLAF6vWOstmi9N
zLCS5jUK+T/+ryps9JUCKwUEJavd8eeLMKk2/VrewYzYTWT72zLhx5BDxQ2s2EKo
WZr4YY3ya5SKB/1hytJlsiWH4TW2rz4x6b7fNYwx/eF4I37PyXKXUSRIotJFNYop
/n2piZNLmNFRWlQjFSpW25jvL+OXieFY4VR2YPL+phi7eFCbl4k8fgTZ8MzN5pGo
B2sAowbt+nS54Sh8+0GwXe7Xc/OBSbM8Fy4chvZnXttuf/MznNGa0u+d4NUOyQRn
RyQPndr3e73hkiOsU684YW5pr3zpHeG8QRasPiDIKwJ4DjM2wWY57BBMiposIc8j
N6mb91jBFRborRi49pGrl5Q8jLCcpYieH/ztA8cFjC1yIhvqP4GOLY9nPEoIy26h
8ZK46vDoG+MidmioV6dqerBfM4pm8UMYBgoWpUMrbDyiCtBp7QPp3FG9tIABVt9J
8az//jid7mnO5/lIV8VXLriuYdhcJOaHw4sbX7/bXNOV3G+gfhGyWfOHJb3sns81
9tfpVIzuCyYz9EY+761BO3FICXXP/qJXF7F8NpfmOckTVK9GPwBAnPWMUFztOJmr
BdmsV1KZhrslCRpP46bAkm7hejima8uKpYbVEIBdru7J26EdtjZnaPUGlfzWip9C
lFzGxVMGI9ucxyukctXLOJo1XEhWJ1ofWYnX5tNok1kWzbAJW0RGUM+nPVJJlJSo
PP+sy4IQ0So2EGye/oMGyopPimrt+I3RfvB9OpAIBJb5+ILG66anMV27890J1tDj
u2jSt8tbMagHRxjcwuj3OI1YNGLgHT2TRIMuKmN5xZJvBUqHecDmdROm9Qu78VDV
7zTE/3GJhWDSFJ8OljHxT364CD6OcXCH1Nq8GZkv1JM/0QZryVtJaLIvntMCzLgq
zCa2z2pPX3dbWphRhTxdLImEOJw/2lE2PiyYyCyAfJu7Atrh7Dt412PFrHJ4mvWS
Lh48px7r6Lii8evIkhqTwd8Sb2V4bO7eJ5p0xSG5Ba6yosDuh8kZv7buaWxfTHgY
W/2uKM2jxCSSB6XhxdgVPnaklylSGnGjAD8e9khpL28U7Nt6joXzWaXTbBqYVFPD
+W7Pen2YSP5sclIgsPMkG2uq7m5CwZNrUyexkm06aReNFFo6ffgyg2OlacnA5jWF
Xf1p9Jbk9RL2TNQEojLMFL4t605HZzG7LNf+CSCCzHs7fCUfZvkUzhrgiPpJ9dZs
F50hJm1BkloXSXq+SmIS4k8yF+qx1HtiNZ9VIJgMeNgOuMOYhihCmu68NfquXwDe
BYdZOLyn1/K2lVK2MP9bgdRoXM+Nf41z/cL58HdhIaaVUHmKOaY0sJHvNOULkGt4
Ft00ewIg+iO0lKE2f2Hls+n4JED7Io7f4xXYqOVgkCJFX9PnXhlaOO1N2IDS9gcI
bYgFXqprzMCDhI9SWRpoeDS0quKA9xKmJFAn3UH2EtwxW9yOyG5Is3AQOQM7EI3K
xMrQNbCcQ0WbjiHRf3BhzdlCNjEZdZGtDcCbd12EAHCwL2PaDjmST8FQL9F2VujF
6juge0Tz8RR+flQZsIyYNGqtwR6jcKgKAxoVUyfPiUJimipD1Fs2/co6R30/ta47
iAGoyK7ydeu4bqOmTVyKH0Bd/TFhWFoza0bwQNHUDnI2F+wCkAQRqndhHgY2JvnB
4cWoNLN+CxsFpbzBEjj31zJE9riC3DSU6LathFCVxFyHhyL2W7oh/vun7bDPqFna
68WD0B0gWrQcy1mcj1MCFOW874ihTGaPHjBw6KVjw/lh3bYG5D2HDpJAk9EvqA00
G9ZSxifB6V/UnR8wVGgt24bHYuMT42NBMTIH1n6u2c8tGUqH18Qnb8pRWNo7nLv6
bmlBQ6yeo4CTq764eWpquFn7dOBbnQGghAib7YTnuPJlT/I18C57cg4xAkrUV+9v
F6AlLb5qEyHl/HatS1BOwU7XydPZizJK4CG0T76YIrATLAbpxdha0wgKcdOcS+7i
EwzOv2AhHqwE+bUUSBk4JWkeC9KNOgfAXgc0UaZJPHzVH3C6Zxkj02esdwBRMo5W
kwPqDqqeRoRBNOnow8kTGslvMCEvrz59SwNpgT1PBJvXo/Z5pWa1RQ36HYftiECw
JnEZj0XGNVBYlsXK1OaYnCgOtLkLFcuBdzarwnxpp8wq0jqE5t0/FBu3A6BZQjp8
XB0AoxbZwsAvVcwlUx5f66AOxO4qR1yvzUOCbiCKBoTDBoQpA2OtY8jAfuZhUx3N
infY8lseHIUbHZZxCc8Zgo7Gpn24eseNHr95jV9Uk7vfueCUeKF+Lkrq9J3+MN9l
bEdwQ0Gmw8AgsqV4RlxrTeBEDikgSZasxCfXXfq0QH7Dl0YjwU4uQGswyUtUNjvh
oSK/qI0hMgTAcmaftzlUXwm6a+I6Ia/DpSsr99REWYo/MPTPKdeqgljak7niHi81
5cPhOlKClQYDyX1sCoslkBAcMZAZYZSEjSv41hWkUP/3m3wAW+O2e9/9dQNaZaA3
powdhBMJ2vBLnvBSMKlpcynBLxyVXHd8Czv7xK5vBc1b24PGbSCF16htwCSy8k4y
a9Z9Pw9whRYrrY2NgTtIM7ExM8T0zsWzDg5uwbIgSLMolF7rz7uOHeBuVHtaa/K2
vC/l5Q+EEaZuJX0BOjPsxOfIz0qydXmD+epAm6S7qEF0KAYHaSqqEhQYhpZzk5QG
8aO0K5/gb6/IghzlkGbxBaRtlDqiyRb9mb6uNcH3UFfzrX2SYzvlsy5/WcjjxGii
zCQ7j4FXvMZxjM29av8x/39d5jTWhMQ0tPuWtHMN01nfhllM6JdX90Kho+fp1Kns
/KLC08DMKufXMgPsaTRHPuiO4igFy0S1XsFoBeLtdJGcL13IeWShU7LS4unAEWLJ
IBJtRYYtsX9iq23amwPJEVpTGr0SxZqLSgxlpMykJGQxbr5ES3q3myb4ogWaWrTg
rx6/+hlZQdjn+AQe8Yy/1guyhlICaWY6YcPcuWUPa/4xaEqxTQ9MJGwPSbyApeZt
l7ANsHWPhv150qzdQwqluAduTMOCErMnuSn7w1nz9gj34akOGN8ykJpok+YiAmsR
lcPiLhZ3rq5eQh0rotMqrPA7Umu9KynFH3WBcwLAbYkyV+sspDom3gsGsvtyKC5t
Z2JUGlFvL1pTMhqJEGcmW1b3A0/SjZOtTR4f+pbe6NUw93AmjXP7LsnWcwJKNfNe
w2Pg3qonIKYzlCRfrbGwQVf8wVnzy4jyYYElFpampHWlhnOBJhQqD7JOdz6r31x7
3OexoEl9iGh80JLljnhV+f7Cg/DdDVYsNXlTV0IqMKhTjYJuTq/C5PFkMyH4L8H5
L/7pcQdIubNFsOpOZrHWAfLTpELh+7BMrXz/17U/n4uq1G1OzvZgQLVD7jyHInzv
w5j/DH4FPqGZr5oG/vkZNCWxyN4dKikvys/MUTrHOnsfAkpVyT3K/1KCHNe5OQ0b
NT3YUe0zRW/r8zR3gEYKDn239iJt9EoGJju1RmemZxPI+JVsvphdWfhs0cOGybsl
mmJakUQN9CeHmt57ZN+CgCZvdWV234StIlCIeTTBFSmjJV+HcuXtEgfKuUq6ZeIK
0jYo+fHO9CaynHcAKB5f1vl1BaWtmCsCBqweqXpnHe/DWO3PTpyZOFjTkYnHbKLG
/v85FLdYoMNl+P/f/dVgF90R4mcBpyxz871CMX5yNfQKVgvALhbjgTX5cFuryGDT
R1MneJ0bqdhN60r4dghj1wmdnxPMdNLR9GhrT5PreArO/YdWJqYgNcVu2lXzjZo8
USATCvq5iSH9I9iaZsAeNtqrkAL09lAJF9yZ0fTg37oz0AKiCGr69lbbXlZgh5Xe
FCK22HTE5YEXi9WLQXNieGOMS2V2ZuE/OoJx76ifxVVI2RJ+tjzGhIK1jQpledGN
F0bYreGwKigD36JsBeaz81fKMyUzLdYouMYz3RikyCaETdu34YZA1gXDOcXi2nts
ca7H3AEngngbMHOT1LNz+fiLoU2yCHjNQJVP8VRASAcNww2vjVJzmw0HNGONXWb6
zZPWl8oj2+J+EMY4VjOqFAERD5fLJBeou7AtuVJt34zxDENPL6OetJAJExXH/iHL
pTGwejehLM44sYkC4TkWPNb8w1F/fwyKmGCXGzhFm8BnfioX0m41Fq+jwu6NqTWp
wDbGzmP2RTzL6i+2Fu70ZfneqbfmnQtp3m4LzTwy9vAP+qng/nSK5bFVZjy9dPJz
POYHdtAHrvInDFq0SJ9VwDqplRhuoOobjogx9VUsZwPRyEv2VzQdAo+5egN3zjxf
10bjNL68aYkqJr981ObqYKrar14NHzWJfOFhLIDdt6BR3mQ6sQ1ZVGOv9GfKx/UU
7LmZew5iDJDSBVKqltvyr1eIhXZZ2+qWZ38DUtOG75xsNde6TiIoEFeAVcqBQ9bx
DIsNAsdsGFd/VM9oANs0YgqbdZq1W6l+rv6i024NeR1l+akFQex/uxBSvXT6IJGR
+P5fN9CYwFbkO4babmqBJI4msoH86+5fCrVkBBQTleie9CkGcgM6NbdvDUpo+k9h
XzzOPoxiWVhrwYOglLx8xsVbcoadlyG3sx5bVebmYgTWnfQS74KncxMw6Msj9QYD
pddHmxS00ZZJEupf60Itq43BAsKdyP5Crx3Q/mqmgYQ4sNau511AVbHdMg3RZzW+
7N+sfuss79MFeOtTsSyyufKdJk+VKkaTt+1IjZSo9xm92BE8J0hAJAfgpKEZ2lKz
GXGppiZEFOqkrOZXx4k+IO95AbSX8nfIP9mxeQnrFTJ4sowpD9BiVO8DUy9lcutQ
RQURQGzNz43TafbJPwICWDgk99Yku4tDR2/FUe6+aWm40JIHS/tCPYYUMZq5Y4Vc
5n/F5yDTT5NTcr7/pT74rAPOzjvu7LqcWIAQuTUJ5xamjb69qEHc5lz998873IBl
o4Igx/HqlhqP3V8LpJN+ajiDE+XElnZOkr6FbgsyqjVn3PfMad+r2trF5x7eZA3W
yM8EipLBTnSJePOyJVBGeM+8pFwxWGo/U/xLh1sJGQ7VX7dI07QNd2Q0ldfqB5Kq
7rmbEzxLsfofQgEbkyuF03qTLdvOIvvZtiS3ynlbeCdUcYUnKRqu6oSjNEzdIL3w
vnkdZxVqcazJyeuMAWXBqu4e+i1Bn7LnNgW9z5IKt/Vj+8iTC5pfVtUqVeQNh00X
wL7HQw2cBFzfep/s8Ov70vSNMKeJwml+Vkk50cVRFppjb5L7Gkas7s0U8CObu33f
DJxEIkyYTZuweqe+y1v37gSgvArtKMfiau3blq1wN8ysMjQts4rs3KUZ7nGPzgSw
cQcQ6x4BByUZ7/Jt2z9kdF6WrXqFWDJfAFQN1WHHO2ZbwQrXiOeD/XoEjG5qpAw5
ZKHeKDyg+Z9sT+ZhV0cW7FCKTL6JKUZ109++GLLu0DA7b9hQOIky911Q/NTwA9yT
jVEdFrtCYgzjIYKQJhv63fZNi0hANk/VWMilG7f7GQdEId3MoPmPVM/PKSNvnzcJ
DOX8rx1jh/upQV3lIlPu94HwlHfo811YEqU4OPXGh0AsPe3akJ6Y6DFrtyOWancV
NXqPinCvr8H9SqDBLQDkeJxHqW26kwCVOS2m1lprPZJINb0zQUnHAOp9L2P9KqU5
xgMf+tFbvVjXmMBGTMAJVzwXBrv05yd/dCZd3+wE6f6EEsBrDc2/QV3XECuOnZ2K
LtAT2P0qXOEzlTvikzLiW+eXpYaUDCOCdghohcEFGXZS8II7Jy4uLrRhgfSczEf0
ETFZlzvtxdctuu+3U90AEcC30n8+MDamqNA8tsfGVhify2SdpeO+y7oxfLiMN3mI
fn3b9rHSxdc+iavpmMKHwRqZ32VczItK3nBDUpbWyWcZJQxCQ0uTlVWJ1Wx8O9zT
V+LFT5N8JyccaHPSMBvFLzd2DsQ6cWD6zh4qMSMI9SztwOqrS3e/pT31TSdQbQ9r
pYQ/9rs33HmqshRf9SHS9l4zSroD3sprNV9sBTSFgDdSsBcF8TV6Ym4zp6tlhibM
yd4Xbt8eN1StBLgdvGkYIcsMKw38p6e09vfPyimJFJ8ZQFMqFqBSKWXtnZJj9g7Q
j04cxwSaxaZZjmQHG31G83tdZSr5GH9TPNuG3D44zxz5G4ogv5bOMZV5COO9/cU1
F9TQlairOUnsfFTgrE6JfervMVXPKU6OV5t6T4yay1ztvLmJ064vLDg9/HfUHCbv
HIrTgTrSb5y0yxCgoBzptmyE4v2v2aG6bWmuLAUJyM3AwfM82xsb4ZPUWEVWRUV+
UG1P93mEn2P0M+FPGqyOFL17C+Uw89V4xo3rk4M7zomjghfxqu5lM/AJCBy8Z9Xg
NiSe92KG/QcazyWllVPqOX6bnX1g7k1CJNmPXma5/ygk4a4wZ1JsjvBx1SitDVXu
SPii9lOEDgQA4CSKXsEw/mMWQnqoiTSddbKvLXC58IetKBwJ+aBf8akOliCkzbCN
xn9+pnJI91FGTvASbV2eWovzPW7pg80WogYrJGcK70JpdaQ4i0ae8GRLfnPxDK6P
TK4YE3lZHIx8wfAsY2WobpdyVxachM/1ZXT7SacL1WEDqoDROH7YSncVFoUOq69p
BzhxN2JrRAt+XLGc04rLmwVnWg3+5ZmheHQ9QvFw7vEihXmcWVkkB3n/yf/96FAc
pbcOz1Qx9zcYZ9M2LSlsCvwPdkrB8DfL9+xo7QwWgkkxlVaxYGubKV4N0CShlskA
DUYOTE8NnpVdazpmL19JYtXuWIKTqF3mDL6Bhb9Q3IXrmcLtmgv2BuaIv9D5pqNk
X29VJ11blLp5xoz2aBdfeDrXn6H5Gj2xJGNOkRUCUx0QpI5XJbBphEv8Y9h6yi6C
hSyKxX6tLJWloCvqalAnXJbO6El1GQk+uGfjz3g/7jRI2ffKThW2O7taxu9mqku+
K9XS412mjfgKa4N5rHCt/UpJtv+FzcCGIeZX25mZCY4Ga14NOAq+7Cy2qQhhA3uR
db5AJIcyLUHyLZ2FCQ+4eTZSES57CmZ67UEdESGCJ0QUtKTNZDFks8GCfD4kxI1g
7Ucxjt4+0G5xi4kpBbUInDl91Sveoa0e30Pi0ou6NgP2awpVMpr+D0+8XTXdQIs3
OpC74EToW15VwE8Fn3mCFrysFpwLC4xVG5uVk228owE9uoKDkWBcTuo4gO9KX2dG
rk2aCYSJgKkKAOyVEsMgZ70bVyQskIvnagwFifxwM7HEQFu9jheL6XyH1mkQ71X3
qxCg8G33mCtbB3i4CZqpeaFuaTBl9lI2MXnPFqCohSv6HFTodbOMkt6co46ZVCRD
Woh8Rx/VyJwM+5wlC0VPGFvuqNTFJNlopqxLIdxIydlcBL1jtwiN/ED9bSCOBlDU
ekLV5X9VinpFPoCZqrZF6h5X3T1lomaG9DnahbHcnwEnvoqOj9sRmH46XVqPqFlU
UUUuuY35a8+hWVdBwMP2T9CBQqY3mUV7/nn/a4z+9on1bzk/GOFMGefe+28WiDFQ
21RwoYHyYtcSgHr4k/oTrXHJ13qAQco6xW7jfo0lWJkGsXfd9O+EHYSVyhb+sBjq
P+Zwt17ciBZ19HS/gKQjOB4P1nyzskDp7rE6IdJIedbHs3WFEQfKW1RutZWBk9ez
Ya5RAmrNWzmBpDvt6M+8THNdXabMZRxm8BtD4BKqcQlYHoSGYpAtgvCzXvZSkHc0
0LvqKt/EKAQSlqy2RAUhvVNsC9+tvR/+kTavFLasUXDrS8WOZFWpG/1BtxpXRPVG
zErX69NLgTbfwF/+FszIj9xXLP7EbrLS8mrm+xjjdnDnmaHrr5AWz6HzwBlUdTw4
pBXFpJKBYS5s1qPl35cw55XnMb7vZ3IH6JSO7BJbVtZ62HLhmJ8A32vpNFcXKd0O
Oy6S78QLDy9wr2OIjQJdMw8QZZmgmionQz/abybnnGgho52mffB6m90GaVp6IF+S
wBWcL9gb9Z102OlMI3l7aCxTcRhmMBln+tVotZvE/xzKKnE70yruY+kYg6vwUNDw
g3BLhJmWevYe5lJpHQB1qe+o64SB7Zgp7E1QFTpib3oguB2n3+nWnEI1pYzNPlxO
+ojq45jcaTSOlwZRlmf0Z90Fw0us2cV945xv4KQcpIqpAgyrMGAZl8zVthe8W1tM
NAjEqi7v2p/FHsIQxDUP5+ZKqsZva3XW5oAAXWNh/aBpoPVqBB+tEp9EqG3NpHER
i8OFyVWqR1QUYEgLDXAvXHVklupehJ0m9222LZd9z8wCrNPOlC8FixEUuzF25HoV
zBlfNL4JqHblSs3vFzpdc/nGs+95g55rlyqnO7KsX7uveIUZBHnt9FItOO8ytczu
ZkFrefgTkDUtocQulJ9+UibVKQqAAVIBXL7CzxFeP51ERLqfwKmRKX10PvrPhF7/
br8cZmBrOk5EW9sdbA8ogFFG+bv+kRSb6+kAdE+O3sgKk0oTS/sc8lsiep4lWEpc
KJmPV88gtJoEz3YnApVynNk2xQ2iQ401V0m01VpqsUUOI5rOVt7vIcEbT9TkAcX1
lEc/04POXJmWiVPcx63pfeL3Z7tCYiRJSikvp1bSTf/DgrX4iwiuFAifuhNsUoUE
xnD0mtYxV+ObpOzaeDjocecgFFXlRBllR6YW8tJd+utU2knIIqHibrlehtFZgKkM
J9Z7YwEhSjTek9XHIFYzBMXecG3ZfyDntD44B1VvNw2+3lscvxfXrDe+z15hnRl6
dJRKVEFeAHwpWEahuCxIs7qzYvMQ0E7rXpvajv9or8c1xeJTcNSnL7187LQ+YBow
pofpXhO1yauN+OYEkH9GR3vD8VHKUxMGxdjJ7ksZmspclBNazjPadf/4f5loZzRe
YCwxr5IVvVNQp5ELUa19gsQcYVkctLYuw5VhrQ886pAIAXh3iEfq4bm90bLmiKUi
xgd4JAtnOnLiCT/W11D9zbouZk0I2sq3uKfQK0dtjPan/UK5rvNh9ri53xYPM2A6
cJTDqr+GQJE4sYCSjLxVedCbuLzwz/i9GWTfq6TpFWBHFd7O1/2AQWKrx3BJJwFc
A4NFQWTl5gOu88EsouNK5fF0c9OlODg/uxWz87MXOmurKP5mpUFTQWW+TWip4Vn1
+jlyUu+JpamQc44zKN0Yu+mXZy56bvemlCNJzq+JDFU+lCyPYIbl7aQ2+UHmwbUb
+8PEvL2dwMbooTpyEaAZLEN23pg1piJA0uOmS67WhmB48pOFO3bBZBcGzNb6U4zz
1iYrgfG+UXhjyPGO7xJHL7nlmVG0HiZl1qSo3rMtLEHkxUKm+HRDSU78rg4Kl8Qq
JSjSKJFeTeLXJceqr6efyAjKsTgTPzVMo0U7mJjhmDuB9jedQSELZ6zKPKGmHnNv
3n5+zxXJ1UOpxyCBduObho17NRTGF9yDcwOFSDIfRi191tRYLRcLy5tQqiS/e18W
amwuv+ZVJO+fo0fG2Hei/2mVIlStcZU5Lx1+37/qgxmRWwPHcH/9+cSeEPyTCUgm
9imgaBGY2iYB8N+cb0HtKL00HPz81CSeXOmIoLUcRaDW0B494JYiEiZmnvxLRN1n
P1JS2t0qAplVEGMMaYkfXPaLzvqEQS1M/pZ92DGSHZN7dfxixLHCrLcmkhTWw0Wa
1lPWt04/sHNAi1w7djVZtok8HlpEENIi88VK/3ZB9unpeIT/5HcrvG0A2yJqm0v6
E9pCfa0dpwM9WYqjdbWtww7G6QQAd8ptypFg7JfvDKYLckZ/DQzCVTQmbSLK1qWc
1Lh/GqdiIiErFfrmwt+SzH3Xo5kA+VJyx5v9oUsLMyrEgDNwCf2ouyG6SPCfn2Z8
rpseKDcJ5OZkTbp/6heHn7mqycpbUk+3BKLBwVVZUm43Nn5VyqD1R07Gst6toJI4
VUuAUxTK0ILyS95Yn1mZTZUCiRFFu/kJoMkIlKJE3SDX/sRsc7JPeRYYVBTZINBk
mZv8Nb+ysAAfSZlXVRx4k7BUOabvdC/+7BuBDJHq1rAnLZ2jDidVtk7j4iOVPj5Z
CiCH1/jp2yAsJMxBEh/iI1MzY5qLg9ZzV6EtcZB2bkjYlux2SKZbJ3IG9sNFbF7K
zCFDy8cO7tym8ULS3qazRXkOZAC8pZBOyAqF1ydeloPwi4VN5ttgq6sUG6dMw5qC
9mZee7GWcFqfi1acepzl+JJBXiVv9wXXWyrP7EFgIWidi6DLaS4+dQi32bjmcUSt
a7y+JGqKTySX+ekKC3AiWa/w4v+yotCsiva/sgJG3x+TML2MAEuNQ3w1A3SAnF2B
NPD4qgTvJVHXx6Lse/KnwcoayJS0X8em3OOk+KY9ASmo9RmsPdD0kF+eygp9eVmL
xfTc9aJNKElz7B9eku9rnEzZm2m+nxgA6RZ7CB5wzU0u2+YsHvsOmkhjIUhlPZht
xxMj/tL7fI7OtpoVBdWX/OEvGvPGqLkWRREeOYPv1AZqhe3jjSYvjabWKrUEUN+c
jUTv/InGjHrT+kS8icCFYSDQ4mhJYlTvOXeN/bnzVU4jcuIxKtlq7L8ci7ObHQpg
9fSJ8JQxM/jNEHLNl4thZxPGZ3JuDVrri4wkORH+kCKf0K9boz0LSIfKq9kzFxzj
Q5gekCBHrtNQtuhFsxLSPByPin0ZLd4Bu6POWXdTjztFMijf1ssp6T4ip6f87P/x
lCfBiTs/MS7/QysFSXLr3hxN3yQGO5PqTZrpr/9CBcEMchQQ8La6WIBMFIRpFZru
6yN1/NZdpeB+s+8IbpmbRJdAdrJMoaLljnXrOxkQQR0l5yNN3jkWxIPbi390k15t
wtPfpGVFpVAF1uyH4AHXhrreAQdEv1Mrh8NJsnR20imRs5c8e2xd9gDa+Sd//xTI
kCchl5woNhQYZCFXQ4l7SxY6QrQxDkyDSGqFz6OnnQHrbkWlM75/9unmh5Qhxv1O
dTjkCIEAMV9e4NEXbFPtZOqV9hctu8XQUWk3eTOunpgIFQElskB+DCar0twWKnnh
xJCMlL63WK6osh5DsF7zR8yIdPH3AdMXpCF+pLcd4xU4YQCH5E27E3sbjD7YQCA6
nDPrYbudNWBfz2NnLNVFDCIr7jMZdlgGn9cGPRxiaLvRpyoxCXTlro7TMcP8ovy+
CW4BlFdYn1/Rrolu0oAk38N6lFnO3FnY5sO4ny9ATug7WEcoEjT/0kDwHrWFDcIs
gxQ2YKJSpZ10YGNmnrJoRY61Hhf5PIIhfhx14hki8nJ+9f9hzBrdXEX/BHHm3FkF
PH+o/n4qmCqjrsfabLA0mM6dXX54SYe4bS/GjCri3jTEkC1R4n/LJ7ZIvtqQAxZZ
yUnsewrggrJnYjJxTEFp224zqphNkKFufjZghIjMOqZRM5GrCNaHPRVv3Lmnv58u
BmCfCVaBPPuDzDOvvqNqqt1NVLXJkEs0uDabg2DWSecSo8aicvo2p7qSXD7TmvDP
KBINJ6hKiOWb/k4e4YnSbgh6XKvlMkadrDZD10UyImZmkMB+B+QSCWjObJtz7ipL
hq/taYPFSVQRQUqQfV0jx/fHoQSDP788/6yoi4AoLL9Xk0yfmVszBfXwT8mJGf/I
HHsk8INH6PytzrcrXyI0E0BCmjZb/tp5yQMM3EfHx8fq5ao66pOAj1Z82Ash6cEC
xNUC2BPRE9uBwgc3oL6G2M/ZP++UhRZQo6rJx+mxpooh32fJ1lH3v2QvnKKSSx5r
YcLxocDlGSaLCjkb5O72KXvlQaNEt7rQmBLvasLgpUlDNe1SVS7E73kM/8EA7T9s
cbXR/16ij4sluPJ3/y0CrWe6ngXHRcYBSk2d6xXzVd7J+s7RfT6Q1skwbzpirUzw
gFhCGAa9VNLLtjNSGWqYZcK9A1wJt948hxFwZPln6jJAVm/Ku8kGrvjKZ7HA7kLm
fqG/6OGQ1k4uHZA+ZX92SN2qVk9NQM9+Xn5gcP1zn7UimGZa4uZagZJ00ZJeVE/+
DBp0GmTnEvmdHT8AenCoplzmXayca9rDkzr+m/p+CFirFhD7yqWhVOPFsMysIcGS
eyOgNP/2FGCjbtDPnBXprXom/MvJl6ZZL6+OcW6tH/Nuc/hjfQRKjABfmzVhhMdV
c9xT51ORhSZOUsvvzs7+pNBlRPr3dalwr6OfGEbp4/+o2O3zDK9HGoRGU+a714T2
GH3N0am9rcRW9umtN5JiJxIFqmDSc4X9LhNndou5eGnP6XOM/TluHfCWJLV3403P
v7nHDnV8EDpsSJjnR7D5p+aM6+pfg9sS6IJ27N4S2ph3qa2UEgG6mrCLbTep4HqD
hByyQUHsPrdz9UtCuQP144OxlH5MrPyGLnUKOeoniPeWKbq8wIXK6mcYRGcwdj6J
OBq41tQiXdYb2A2RXdAY7Wm1HvVqFMSeChdRS33yypBkgT3143m34KxMKAxGLff1
BvCuJeJoe8PLmleEY3IU2CQcKuJ+j3PeXuCMIK2yKPyWiWA0wiB+Xd6HiKzG1XW7
Sz92gANVw2mpIaS0bBCFiZJjV1+De4tu7kz1+D4ubLxx1cbmj3g9dHuj09A1n89I
MwAuqogrRK/EEaaA3jrr2FR8L3vBbLYdA3BKB7w3+Vf3zS6xvH+/UCnHWSrWywcx
pljo2SM6nom66u2OBvII9kCWCvD398cjbRGV/hxy+L0fjT2zNa2SEmx4fhu8rBom
5pMXBMQfQsP1WB8UxjBJ9femv1DDISQ4oQiBH15uY21Or8erLFT628Ih3rWXnsWP
K1+maadpBiwCsHW0gTp2tbhiz1HFUOSZzpPiXZusMPPZvztVvaDLJwPtMpxnUGJJ
WOAS3WjHqJKuFq9NkyaLOAGGYmrTWdOzaV0frK7poYE2juBVd8pCrX0ffYt298Ts
Va7mHmV1Kq4YDAy7Gx4wV+IGYz4djFvOM9oz/Rnl0NUN8X98v+gP9xnFYQChz8mW
DTjq9l5ruSvmLqgnMTV/xpQY3mcPWSk+JCzjJP2sSbhcFb4RSFhJ/cruaw9ClECA
WFRpon1yuZoftMZ4nyHFKepUM8XYQarmdVw9Bt/ei6ypTWFsdPAkOc7jgDujyU+2
YkwnLldj7YSy+E6ST+2RlXEHDzM03Yl0Zw+hwfs0Oupqez+lVvjxGdXJjmKRKYs9
kVU65lv9/vKCRhAr1Z5M0tqDTWk7d7s9Fi7+w3w4PLHeXXfs2cp68ZhFOzep4hsi
Wuu7PpEavBdtWlRFAqi0s3nAcvox2iZ13vIXmg6EYdQzcNmhU1LYGdIo+orZZq4G
rcs1z+vNx/rMuEeo0IBmSMhmObSgGn1gT4BUEd4JxW4//qWDZLuZaVVrw4trB4xP
igmF7vuT41wb8d0R5gNQReuicr655EVzUEINVGP/fxHsqbYwg1oNa0OZZTkTkl2k
eMVnj1a5eVOII/qwQDqPZKpbMP8X24r6GKVC96IwbT/uwABpXRElLe5QJ4oxtpOK
t8lybdogdwNODLVJFMZX9WpU6NKucUOx/VFD4VqHMN0IO7e94JRL1Cp/vcdAfE4S
DFIE4T5mjU+s6aUFXJP7lDuY6QLDoCQenquDytKEg+ePa74Vl9sA0ax4KCcl3lu1
DFtb+aZqJvzbv70yn10BTh2mVOy7g4ysLX5LUSvjv7ciVNv4CofWTQynTuF6x9tr
DbbDFFZjpfwjk//RqChHeXgh7XUJhasDJP3LEzBVmD+jCF7qCAYqbwT2oY293nc5
V2pZxOuL5FPG0eRNBkGVlUs0Pqa74zxPMdB0sbtt811EFWek572EBB+uTxMu4Vvr
+ja8qj1qiocuwBedzzUrPoMyHRAeYkudjXE4bZjAEopliGAJvkB+D8XAY7SjW5j4
HvJuW7DdjhTm60NQgl3Y/jRB5CP11+bUNtS+Oc7xdeF/CmrkwlkGF48yV0U/6+64
fNjqttmvVC+cwLzLkLTaSvde7ZlLMXPWyetU/MalAzJLZyw5DZZ6a4K1bLAloiT3
9QDigoPhlgaW2S7YwCxFlYScM9ZGsuWvV6OJhAdwkJLI6dyse/dosbMiUPjNzIOO
Mut61Mkwp4Tsg7O8daQWq2wHyYvlmJABUqFtF8OvQTJZN16ppAEk6elAjIpexXmq
3PfzqQlVftWWXp+nglGlmk+A3CeMqkmX7s5mLJmtbycEYbllRXhoH1InEd/MbvuR
a/4FlgZEjGiQ77hYRQE6WPW8XfoeYXqqW+ffz2URgL5Q27xhyIJ7s5lAKh0xb+xM
fXg+a58ozbSSlzf+lVgeBe3EI7ou0B5yB7SWewnjv2a7ZNWKZNXo+53yphSmO7RC
g5aZbWhSaCjKdMRzCPCpXHBHnoLILglKL2xQlDwcCSUyjDVioYjy1OOw1K1Q0d28
fdRQyvzwwsBMU4CQ0O3VceQsErytkrEhEIuE38P5U2BYoSyXSh9/fll/zi07sIlf
fo9BXcUBxd02cdv9c++5W31l32LNuLxCB+V2PBL/ODYQv4WZb3AtCSNjxBUduwQO
wqfsk0kDxgNal0Ts8Ru1nAuLr77FXpYh+4CbnubybPM9gOxpe/oh3Ur5VCi3URSG
NtMSLGearD3CWG4why5W/u3kVX+C0QA3f1qSYTW/Q0UXrw3W2xjp+XZ0vAuamXPA
n4UuvcEhQLEhpTFkSMIlthv5fNClQryVJyK9Cy3vl1V7PcgePqW6V2/PDLde0mJs
it5y5je/iGswPwShCXE5WWNX2KdKPN1daWfbsVYWsdu6G/lyY+evqfalds28jfWw
tCwjAGBTBvNzgYfuoZyf5p5nmx2oeMDg931l/BaVEh745D0Bm9A5skMw0eLvjfJV
ky7S5tVy/rVNGCQnGJ3fsm0jDO5/FsWX6WKFF0WRk2+sv+JKMFNUjLGozPxzYeSt
zXBOwOozit8Nz51qD1rD6ZOoJU61J3JypnT/5eiBpashGBSYw7MZR+sguL04zufL
lHFv0tjfvJu1dg43ONbQY+Plxhuna+ULd2FymKJzF8Ov7H80MkhXZCtiNoKR8Z2W
1yrhmP8fs3JLZyRlTd8UhSrXx8INsgt8ULrji+lY923GXVVghakulwk95s5r2gaG
rI/5gwvorRjlxKnhj/TNVddFVHI0qYmtGQMbdYNzMkw0hXW8VjkUUHWEQP0mhdnF
uub/Fbmpjd9101fwIS/81WP928fHFCWZyjjVT/q5MqZ/4e4AMBalj8FNBCJsnKaF
lotjiNblnMIU1SXTKG1ubvor5A7flK1VlfkgDKlmgxs0yheRba8Q7CtBV6m/tXfV
YlvWnql/KloH7czO0grDPqduMchw+GNGbPIje4SISk1/y8IVAg19tBDAT2U/KI3i
WH0X38TcBoj6yrHqt3Oahi/ndE64u/MF/sdr3RmhnJaJwPOjRbwjfSUdDTE7+h3c
IebNALzpfXCMD2ljSogtDxh+EDyh0QTc3/H7ewPfOLu6QUcqR+iziVBwyRE5q+F3
z95YOF+cZnBpygRNZgRWlfMf/NSr0AtyA2fbodjM8nCcfhRIC+oDnRgG5rO6v69H
uvD/7FzI0WcZ7tXg+QTY9kVevgT5Kr3nP22M82xjBH6IMhxpBpzoSnm4ODgqvt6b
3r6X/XO1pZybW0JW6XUm6a1sXf7LNTz2Zb/e5Z4N2wVSohXvKCz/ewCWrcguORUI
fIehLbLWOwtWqz2qcE2McdXSYOetQYg5BuGqXNaUgjb4hLhjFe21VTe20F/iRUWE
f5OHbql+Z48pJGMWmtFi896/fr/EgUVk4ux/BnvPHQh9pkjf9i5vh/+TYjK5+P3J
sH4PtBUk/4Cke3sbEiRopzuJVM53p4mGyvLWc1Gqt+vgICcV3QRsxnt5JvbXGmEC
8FjR0UYuf5qRK/qfBT4dSYBA5WJ294ZWVBZD8+rlLKmPaz2uXOwcylAPHXMHMWUX
gD3Qbf8WYDfhDP/+Ll99lhNxszWOFhCD/BS8QHtVsLI7M1cc60iAUH8AOm5FURgi
c4Lzw42MnmrWW+JBTqkZk5O8MjdwVq2REz/fCCzkadjfsGU4tFJpcgODF15c6wY9
Sxa/TgaVY02wzqZgoCLqVRGjAaW3Ult2xq+B2JLpA2TfoKaCGWOAdsXCkBVBX2J9
s8FRSmZiYC/9xjAaDotbWGc9wyqiHhRBLkLd2CKtZshbzrCq/f0qZXgPVkLnds6P
40PpV43B0sR61r69Fe13LkkxEYzhfcFpMFo9fdMCky7sv4/Ian+Y9qcUhBbUqLrE
zi+KuObiWEwkPjsxLxE+T4gxDWH36jTrUcmU5f/b+yizaxj7y0LoC3l8nyBfrSXL
pYbBQ/MdK/FyG3Do0KqygGu/iHp6YgdZO2h6JKD4eU7Ix/fEvmEh7wzJo6cUZToM
R5c2gn8sWrAF9oDrZ5zX3F8PCtvm6cpycZaQZnpTbUNJspYUfSIsh4yOiTltv7h9
5C3zJL1Q//RuIgWnTUZqPNVUmV6uzK7SVPHboNNUE0YYi4OrsgYjhouVFsayLL2n
uHtx0V7kf/JBMo3OhWc2emLPQUote6eyAA6A20tIx4HjRF9+Y+B3zpsG1r/bfd8w
SruaU5pKdjnsK+KeZbeJBTP+nn71DiRIlyMax1lD7bf5yLS0vUMKG0qsQlBwfzq5
rxIppKHTpP8SV8gm8JnA28usEPNQxciZbswjTkqMmuXOzPTJaC2ynKQKQ9ooA/yt
mU/jb5vQy7XDQdWRE2MLu8bqAYsz59a3PP1+H6X7aJ+DgYr4Pz6mSAjZbaXRmn3C
jWdmArkhwr+t0XT+l5AkHBqddA0UlXoWlsH1u2EXKw9Yw3seT2wLtbcD/hbjwDjF
YNIJjfITKlOgeyMKoPKsaOpN5535DQCIYlwOEJVvpckO4/og17B814t45Grqjy36
LlIEdu8iUdDm7RGeMAsLVi+RAZ25sF8KJ1BCJ31zjxM6MijYWbYaje6SEP1KNY07
UDGmke+zgYscUiZDy3Y8sSMCwMTqHx+FSMaE9h5ZfvHFZGLiFVgk0SNPrI1dZe8V
HM7/Uu05XAa1kc8/yO3Bt3zowVc9tl/GNhydIGKLcEcc7gWfDmaJ6rodOXUcs2J0
ZFFTaVKsbTVRuje1V729SFsKGLpc1Q3QLd8pBr0KsSdT94XCXS0ausQis9UBaLAu
lcWP1FgRMOuNuDFzmkcImXvwd7mZ3lzRGueu28I7S61iflU9PcKALpqKhxyFRqcS
sFYMI8ksWHdwKLPHruWZhyum1zF9rK6njcuTjWSJj7C08I0IUXuMw31Kfd9pPYTw
N+MiQbzAO+97Gwn1o1YiSIwOPKOzmDJHTCrKkSP8XoGH8dAxqV1mpkmHSHp7pSy4
NNbg6BzshPAkvRUgZ3At6VCm+Mx7eHLE4WWVdcko8Y1BhBAgRNNidqIR7e1sukni
9RhoVofYvcev0/K8a8Zg4xRrbHS0ntXJ0M/P8XQY29S7C6UHQG9ftAMXhL2T6169
iEw6HDSQzW3T86MFlLFKKNLqHfq4d8l17+iFDUg089F8cIVqMdw0/BjbhUuT+n2p
xrJagMb2YHQNKDqH/BBCQMlKK891ug5r7DoEmcoPRkIfCX+DxWfG197SpCQ8tAJ9
3d0II2aJqR3VGxUDp6aRIq4X1LDIT74ITO/XaNfRp59euUP03k5dArCvj0To9DUF
uop1sQtu28cJ2cddIPHQPlNClcUF03o8giQEbx2HUOEv9gkBAtjJ+fKNZdaTGaiL
J9tUee/Z5mfVMVoMD3rMY8LvSqOfuisO/N2uo4TKalc/uYp/vGQl8yU6CmIHA1Nd
Qjva69uRFgfS/xjjzNBtAuQBoKQqwMSRmgnAdmtACpDyD8eVrldOSL31FfQn/+dr
C9gIxZCFhqczV/MLwAqvM3K9sVmU86xWNWG0at0jKjhNaDG5Tk7YDzuhGLqbNaCq
KRlUUXdHoqgUlRpQbhUPAZX9nQia2PcAgLtGHEK+UddCaV6wnskiLLFWZY2WuJt3
0AMiONaMoyS1HKJoHtDqxvsxHwNXgz4TBEJUeYTZHoWVYLqRTMeUD2oV2PNdamg9
NFNs1izgiyl3c7x2w4hundgbqVvxYpl3xVEZ8eTZiyRcUljmzOMn9pUF4Knj58kh
JtLsjdj0RXNgk9fLobY26xYseS9X+8qMohxlfl1e+5rytNXhyJmKKRtWseADMgy3
LO9z6lF2ogDSNH45SjVjy5zHGi9fV/1rHPBcztqXkwZ+5F4/1tztBzFKrSOysLrW
skopULmJgqfZkLXLrua5/uVwbs+64dmKzQ9ab6xXckKZ9M1bkyrruMppQjjGWrG7
864ShpFBCn3CjhBYv47ix40bosIljeYaHcrzXOJPrep65pDmkyKsQb6J0JSPrJS5
UOOUsiZ/U/WTPsqHT+YSsqrZawbqlr2Lk5+tl68s/6Ht9Xk3xagl1X41pDNLfEIU
DvL31mqX6iJH5BNH776LIaeV9QAL/msKCM0geLsfKMQ/plh2Hb641klHgLnhSrLH
yNUxS48WAZSaN+ze1xMLYX9KE/ATYQPuyXJECy0En0pUP2N6/qN3Aghxx45RAr81
+oj6uY+IwiBT9f1FlZojnIaBL70JoRvEivSz7HdciU/LdoJN9K8YFMS9+w83myEI
2Ze+2dPDuXj6BCRpED9ULws2n286ry3MGvCBvQ6oG8yTTfGesFFMb3+pCLXe9iDG
jo2gYlN2xn/dhpFW5thAILgLLX9Hyp7ujhIynSf2bT9vB0fglMpNq523GFjGtDvl
FQE8Lc8JqdaN1uoSELfXzZVgtjl+XF2maDFZhgTkKHdZv+ELwqQBqXoe95slPfCB
hCM98W8uExlbXSK0uInu6EZg9vwSXRQttJDlVDIdRoFFiVlCNcU2uuNlAG9JEy4G
1LSaU/e2jPcrJpuMQlGplhpd407FAnxBIlLS7TE7j6WSMs86wU5lw/uxZ+pWGpmN
VOMwpkrRNFAJe7DYpI2SiUWMcA0QChDfT+V7M3VI8MknSEjtUN8Sn+Fe+/TmRuf+
20B63jO1HP6OVcmPDAgiYdPXJK4qrCO/KDSt53kjxfXByK+6okUYtaAn63yqXLwq
EFp/ys4Sul54u62K4FCUSiteN1n8ysmOogGZAiLncXw8B3sVbpCVKpVf/WgCznY6
KfeuEwEY3X3ZT59ZMn6Us2HroybS4i0PIBsA/xb8XDaAtMI3CvoaxPJlkbVr8iuQ
ltY0c3Tl1+b0DFvzFzIZsFUXKJePD/wtk9z2BxNLMh710+EXhq0dU/B+jj18Kisj
VS/bBQakZgaQEn9JLkRLJqfNkZ4YoQrAV4qpbksAxCXBxBk9vPB4jr/vdycGa3qU
D0IGPVaPus6Bo6AQHnESslcID3r0Ee/LXS5ZeP9O1+zL+S4XHrb+pLY7+7lDzWos
kyPE8VwA8D4n/3BmadZVlCIPGGn4H0AHHoYGnNB4QE4RxNJf/gSjgn4MXZVTsMhs
2FC4PFmeNTPMc6HSFny1I4z+dheDhdq10uj95XyE9kDi4iBnYqErNX/cZMn3X9YE
90EGBclPcT2zdCTY/sLU2yfZOCFLaDZtxTh3qERan6MTG0Z0JeXN2xEjCLUYU9pg
NddggRTYM+sN/oGRbzCxfDg0Vnpy1+JCTpsSmuP63TiBTi/Q4cG8An7SVxTuwnTb
CyaZQDtnHnXEkk+ttZdgDiUekZG1shD6Jrw8X6nhOjjLNWB10Rgv2l6OY3CRz4xK
hWtG5HX4cdLgsd5XBYrFL1wJnK1V3etoABhrQ5aytE4TdcnK0D07dGvTjxy7qShQ
CSr7J6cPGiE8ODJS1YmDJ22sTMnc79uev8H4rJj4FNM4pOzHR7HGsib6Ph8cDkzp
6wpvUoEwS+M8XHUlR+q7ZtI9KMWsO+ke4ukg4zHNwdBiZv1qHONJzD1uWXzMI0ae
SzVIleon5GwFAOODkRDs6U97+4+0keb9GpAlX1NSa38cToNlqR8wwOgHF51OW63n
CFODHQTjcdi23+VpSBSKsrG8hQJkPAUhLBJLV/dCC7aZ3EprknjdxINyanUh3LfL
FKBfSVJNnDJoAIdhLEG8u5Pfzn238w08yf7os2srCxUm2/JXOzK43/EsrPyupCRs
wHvk2Zr7bAmVDJbYz3NmHJc9n5wIx3bMmigxBnUWqvDn20YsZl9quiJySLz5wbYE
CcZT3X5fdvtNWYxHyvFbueJWnPtBbUwDV83vEbtG+luZIQn+yByO8R/u1Ui1pcTG
tZPzX0GA+GQkkTPXfQX3y5+WuSLmf+UK3RHgwgdKQ58HsUL5snYkimGPphjJtOdL
YvcvzffHzVsO1eW3xvnAOA+zMrvo4HHdKY/t232/ZR8Lcmz16ybAWGf8KFavrstc
bHEJnH7Q25qhecOSCICKudJv5vNX+/Rvui/hvnwBa5LehPWZiGgNW/ajYHK6PP+K
GUorxELqBZQO9tf9ez4Qe3ZLa9wImcy48MdFovHIcd4nO2CRQhcHueNx/j+fbh8G
f/M1xtVXSJ41bzi+CbHy+SBOrRbvZgamZmRe6H/ke+pj1hLp1jf+Kctqdq+c5c6+
4b7rcLknFxgTcUSNbcB+baXHNnq9zCrYLhDzIPIA2IdHgxsfg/2SaK7vGBfJDV3y
IL7T2mmU4MAvvD8Il2E29gKaRUKFD8TgJcu5j5tMWQ6sDn1IJty/Mt6mJW+SD6WL
NHOr+L+KxAHkwmezkKX/HU8N8AXvwOG5pXo/6XChDBjZXBG7YhY4LvzjiGqhtVNd
QGxUZjNY9TaejcILTUKrkWfYCe2x+qfZTn9/IrIZtI3Ld9w1ZBU2znAu81UXXotu
MvKeOtkJL5Sm2VLv7SoHTn0zcqPzuesTsP4zm+nh5LCEN22mNJkFFh3+KpRxagH2
Nw3B3k9H3m/9d6idSJhzrzIqb+hP78sJnmCDB0UUz1c9s4mlfBTRcGL/0KYTVTJ9
G6m465Go/OZ7zkLKPp4tmcZW1824aNY3lxOfgPtb6bFw1zZRoELaaPRfictREW7g
l9XyIXPpNq3Uf2fgVKmEqzq23E2aBJMmc4mLXXQhJXsJGZwCL6SCU48EDZY+OMhF
YKo+930NW+GS43L56ewQlBjto6GnEhcRKxs7VP8VyFf5kjxQcGzIW4XD1kkE94CT
dt0VmxJopFXdKTXrgD7EFaVvbCPXzmxx5DyktGq5JkUbbqTq0aRScftEvbV8biBK
dG9UWBK9+yvMKLiAehcFxQSTRuiFtUrpSObhhQYOSWO8eQVCtR4hOSNER0/6MJqx
u2oDX5Re875HvWxy4bv325TwmVsB1Q/0IAgZar04CAVo8ABiQyt0R+QGNsuz2I6i
pET/l89Aprf1olmvdnaY+6OS54u9le+fzoGXoE1ldN2ZaWNWamZLhNGeN/tVfleu
bx+Ub5eaXUZwtpA2zOy3BE25P4mTkjRmL5lG2NHn3QNtuOETHMR5/bk+UlgxZRdb
54xbT1ktPpGKM6QL8fr9Di5QzHBJBmeyJt+r0FzQ1FXl1BsHT9N3GtnbQpKc37Bb
zSY/MsNQqyLRa4wQLU07z1cJNu+Uleg+vjdrnNWwmw0IhbENTThq062JIWba5LZy
UMZZnclfRLkWZeLB+ol2BoZYmgn4Z/Hiavn5OEVSAyuWvt4cNzRXnjdsNfPJgIY9
/nbeZP0b7vOj7LEt1UH44EknRRioDyMFdA1wIZ20pmPSqOLYPKeRKHAcAgbzQsc+
J+2yab66Q1tgIhBacaaO/mbbLs7JH97jtVdOCapCNvv0efHmIf8IFIjuX2wNDDc2
DMqGHMCnFBBh1Z+TDWwfOtj6ShspeK3r760d0Zs47i7hywZ8qQgbveWWuRhtOTO/
+cwfTUKEDWcnaKE7nwvOr4V6WbVUmluMehL+IGV77c0B/RRA5FO9XSV3MjI2anKF
RbelhLW+dR97f8iWvMC99BmmKMS3MtHY0FhUTt1Q1ChgAzs41l9MVnRBTviHTvlN
mSNUKKVDh6hH/NYcS3xpAAaLYoHMAv+gkFDQFYiiXx+AMUPzuTF7I88a7+nZzrNP
3YtlYDmwrH2L42gtuIfrHbc5GO/oyQUDkuXl58LVsLBEkF5H2z/UK57R8YfEgPV6
ywlNkKUj043/Kp1ySei+7aFydNtM1Ecb67E1PfxLoXF2F8ZX7Cjt2zwD+5I5KHft
c61RrrX29BZgH+uoL4IELwBV/Nf3W0csVLagEzWCFXZyNZLSTB76DYsrvJA+bRXO
GkGR3sXwpwl4bj17u6rQSDkdOXWFrl5DmlfJimWBYNbhvu/PQcUDExkODGPd/1O8
AEeLk3XeGW5n6ZQdL/diWrAB53YuqM5Awlfm8cPgVci2Tdr7RkdKS4VfLAxlNA76
nyMCSgvNHCEfbeK4VoC9beQCLp3eE+UTGjJnU0PMJAKSu851xk9aJTpT+Gzjv6+3
5XamrupPWOjKYbFhmTdJ4KHb8x1mWmGOjJliQT8M6VlB3hu60qFT/V2XjQvjm0MI
2wMCnQAMtRARmts/Z3al1rM+rnXDQInlNUD3d7XYNS2PFRQYFVx3GXDS8rrbDd3d
nmUbCGN0IAWLsAt1Mhd2KJTJibPFuvhALky4wK+9WRSqpA29ZTY7Qq5rRV8BZNIk
dy3o6zspPSb+RorEWT3H3cCeLS18bCQSBIhH4tzl2ez9Cm85GkTVeeknlq0yQEU2
06SMaV0S3BY1UZRhNDUQS5B/12fUshwZHM+APUt1H2FLosZl2QdThY67mo2ZjNzg
tVaKxS1xjnzT72WZAsY65K+EDvJcfwCgPWOv/4/FEWDfSuwBxsiIbFlvGN0LDaYz
NNnz2aoZ95hV2EVlngR6cZZIvonxb71BQOjVz3qxUfQ9Ihx0JFe0e2y0FMmmySen
GYCGS8hVA7qh4qnQYhEkIpyG0j2tnkD1PmwLAkWHHd+nIPugkks/u2sFKo2zKjk5
DU/+WnDd2KjSVgdriROIlrlRtYfzQ1TThud1Lcx9RlHxVqIHKSOhWAjkLq2kKitc
P2ZKrR4lKMEgKkJzLZpmLkTk8n7TXPtBizlBbtO+j20ggEGjwQc+zWThH/1H/cyd
FUZAsbrt5XLfiCZ6POB1nWkX0Amg72KbPAMMDIR7NNAKufbscRAektSAONlUV8ie
w0ApZlYQTScUa0o0wfDiPkueLwrmFrVKW2MUGrVgkInRKOTv0UAHzjeQYyWG3DAa
IBuxM+WBWvAI0nZ3RveqbGUOyj77exPg9S4XNIzudbVIHIypBdX+4emzhP4RK13V
Ws6ZClL5g+GT8vNzcSmOPL9+orJw7DiWldY5r41iBFah7SFcAJLwEMSMSA7vtN1Q
ixtIs/ARwWupMfL72sV1Cqf7/EUMm8ya9gVIWAU6k4D5zZ2H10d+mDPXgtHyGLJk
hNSWS7hLSZx9mJHLUzK4avtN0g6lcqm49NIv+5Hhw2qtPkDpCsQiL3lO6NVVUOMq
DSRwbHd3934oCbYYCfcp3gDXBynTGUUz7g1LZhr1oNWGfF0LwC5RWvv3W00QLn6j
C3tnECiq75bqE2iuZk76PFpo8I/BYMvS555mak8g6McqTRZrFdL8RaUmbe1juY0U
UBuLJrcxp7bccg2bFmx3tmv+PE2uVc3UM/cHfwqW0wlXr+qbMLEIgzSrVTFWXwsK
HwQ9doGr3XJTaK2FVqmOcfGHItZ9znjEJ/bjOgvQkAFjdQG1kfiTcq9fv9joQY6l
eUZeVC+Yk+FNfOZhFPep7jRle5SrTG9k/EHzgQmJwJyGrHj8nq0I7PQLETQHZFjj
tSf/JVy0a2SWCYwlp4c7sg6J5U0pmPyJlatbADo/I0hnHrcm3bVYaD5sjswtilD+
i2WqF+9UwmwydQ2iGUdSovksPpT+7st556G/pRKzWGsY9t7bIfeSG2JDyoSL7JcR
3YuOuMM9GiP4nEX+L4dK8E3x8F2/5A3blfA/X126hsfIZ0lKFmAT62y0F6TcVxrM
l8Dg3o8Izdv6I8M3wHcf3Ho0Bxfcu8tn0abUOZGcZutQfZrhRDWxVFGHhLH9wIFM
IGi4CUwkI8Hatv9+P64bl2pNbqSabyEcqrCuEr6Om7j+fmx5JsLS1QEswovrtqmY
9BXqT86Ka5wnG+aZixrm459yL2aCGyH7kWTQgPeZnITuRdboNsfgw590cnfVwjUr
gE3dId+b0/d5kuB2XMXFwChQd62/3+2I3+maL2dHw92Ks2j/BhgS06Bn51HDxt8q
veMrGdrxUXClsaj0ZFHmMbvzl02qUURVkQInGud4s+fezRZDo4WZBQLoCkrS5V87
FoPx8GDcPRqvs0/DtxA1yDfjZCB3Pv5EpGxb8hBgzSQmIJ4S8+deUfWIhf9Gq1Uy
uCXvY9WD4u19+iRcWKDGZkQPHbPYjQbGECACwJwnqCtWRrgrNoEzMb3UyXtUMd2l
zCfMMdO8SutYE2nTKgTm3AQuazYAuTzzw7ACarlXme5z9l/KwysnQvHL86/eXbGj
tBcPSx/f7cOGdtf9Se0sfmJo6w4KJLvKJ+GqdCOPFati5UnEyI6NdJ0PC3MXYWW/
cq0DnQij0qmBygp9FcAIlx7eGCHBMJUssSEoihnTjnesx+qHZiN4zIcYjlgzyXAA
9QfVve0/4sWRYpZfLKyxSWyFMrHAum9V6Lcfi1axGJcAmIuTp2JTZvQj2tDkqTST
U9O7ptlhydgTWUImlhtn8vlyAO6jKSrhEXxaOJpbyWj6Y/yMUD+7fyXQYxsXtTGs
CGPunIlQ8aZ8N+1N1Ysie9Ad4k33mRQxN1zI3TO++QqvFPo/wOFAfF8/LRQR2H9p
O0I+TW7usVL52DDFFJUzVceHb0mvyrWWrCc+1BohP0UzhpjRsXFk8qFmWPcDw6i/
hJtHkZIYoQHqa6CHcKlikz7z3Gpg1URri37NXaPjX2tH9sYFVpJuVJrSVWlz6GuV
9YAQAvfnauoFlkKURfmRM3eL/wbWZszYYZ1Jp36sNpSAqJef4UxqVpcn+acgMWI4
Pp5KQlDLTB2jz2h+GpiCOYyMy3NEtLIOfWMh+jOkjI+63HTJ0LX73oeEjBv+IH2i
UpRS24XzWZKUmu6VuSI3bKvZ51/zIBKtjkkLz9d5EQEYjq6hYQ7+UjjbCZ1d9Vj5
u8ZSj2RBijSwwCifxd9+0NkOHAmyNSeIoGgxG66ufXU3TK1qAeCDI6DMu4778rVM
9O4qHW6bdaKV648HvdbwJAE5mHWFG3cznQrRT+cMZ9fZNgtCIoIUVhc80iuUSy+p
EAn01ASfkcTc1oCoLkKCqRwpGd/YfkONkjGOPkLIPMbByRHmbtFTsIuFMA4Eb+W3
yDoLMG1+XYg6J+1s0D59flBuxoIaTvAf+/IL/xn3IttI+/3YrfAtd8T5aVaPoNs8
l8aV54ESJ5iDRf5fKMB6aYkr4cpJkNnLkLzzyCoI0d+PKdhRcsocXaD/pFKCfSpw
pIfld5Kq4Xwh/sGveZRiUduoGOWZd2DYoYromF+/gQcgYhm9yUbsm6138Mzr7wq4
UQZ/VnpUqXFETBQLraucanjguF475ynh7j2MJb179tbP+2rvoYU4NIV998fRFzol
GAD8rxR8eVOX9BSklv0X7g5PE8mnuei+NkHgOBcrxFid6TXsK90re/Q4rmAC/Qul
/ftXioQaPhCChdwBhBggF/qzbdBaBe8k/t6ei3hpK6tExkMWr6KNxop17Hqbvvcr
4eN3tUO662vGHzBkht4fRUPxSmTDehWLDgipjElWxKM4PMjjPGIbvx0jYoM3UktC
N+j2QrxoNLkIPDNKp18hHRzoKt4UOFRHeVQC2Ba9n0T+Moq3iC8r/P91lAj2nNde
mlyzoyPaOucZw7KdDVaDlzGHmxdW5rBkvsDrgbOb8RV9/1Lc876WhnSKKNRhmVVe
N/zZ36S46fZv30pKvjYWhdpYAVMeblkodj3c7dMpC5XPbJqWcDhkJtel6t4VbDWx
d1xhklEc/25lN9XJ09/ZkWJRASdt0WMdETtqUgAsELIjLzWULd5bRn5BxUjeEdH5
QejjWIye4tsUgadaHJsHlccvfWgcPiope+uWBYi5yOTyaXSiJmx3/iY/c2WDAcii
1DouJhmZOWNYuWBCraLDbONYnXxef9iC0t/gc1WeUlgBUKfp1hzSm3KQBKQ6moc0
g7eTZQy3EaXV7AiF/PCAEs4a4DHQy3488ixHt+xdfn69rtgS6WC4JANO3uHonlVU
9c3kfXocLGyPi4oP7oZaiNglYfdANjQrD8JGsYHbG+SUpYhLz/KGrPIjx33hg3bj
mtFkNK5PUQhWDekOa4FrIAVwj8lWSLhegUPeov3m61YUlYPlzh6yRyzXMipyrWi/
lM58PoU0+x1o7uI/g4FLXI0ToXSkEth8J8k0RrBJ8bQgz9FleRIQ68YR/ncGuNz8
POA+LnqBTPzcfpKBW4CBtBex+2v8qslUArZAsALaHk3WwQyoNLTHGnZaVQY3iCC2
ry5upvD3Jaa72SQa4X+B3XItnU1ptZBGy1J0EewiLmdfy0wMKS0sdNeq1aeEOuoc
ckQqqvPyrc65azO7cbtOZl29/hc5M2abX2DWVzJd+td3/jyZU6u/Lfx5waqg3YJE
oWLBT3Zib/C9AQvjOXYIV5eYFpULwWZF9u0k4EjBdPA9pmKeCWRIviBP93OZXU22
qivbvURI1qcmhm64QijetPisdaL0WhPHHJ5NdurlQ6OwlwQbMja6sYltTpVMwR2Y
j8mUDL3slw8TDn0v9FfogZZ5e6KH6ziugnhEOF0I4u8zA5lHNvTPp/3kIypgUYJz
MyzZfTrXtm4fNBOFvkJdg9nupVvMs2FJbW8XRa1Y0k0gbkC5CCV5a0W/O+wFW3Ia
l74xogpSQILVIvz5qFMdYIEAMS3GDmVEqrLQ60r0QTY7EIZgwFIOPlpRxZwD39O1
oI+J1YKsA0H4AtZ8qjK1Hxg3Psds8AHnKnqcnMtjCQQ68dEbX+/4/eCSEvT+kTSw
JGcWeNF/Amr2JXoloDQR/OUgx8Rt9zQDa7IZkOSM3td11ZHj99oYf+rY8gRStqRV
bxU+rIhRiIb1mAvD3nfFugzOkO1GmrKpaJFGB0tAEuinaft3Kb3x+DTYVYiHTWZO
BLTDzVDGUhAcfMl4duiLSQz3+WatQeKr46TnbTCCP2s3ScjjKJqIJ4Hwdf6adUof
fu7p9hSwLH7vFaTrnIFc6AK/u5NbWWEJVeNVYOHVxzl6xBE32rf8Vpe3cAXkOr8l
vynKK14pumAq8/XrLyjLyAq9cS1IwZejyfzJHPUJa/sOzxm+P7d5If1gDymMVCAQ
7HctnCWGbfxpT72XoiQhuJ6yOcWxQJOc7SjwnCWGsfvEoXG2It/f2tBPompGNc9L
BqCMZoInt1s4M5+cg4Ii6E7pgOBlVqcyBupff2p5/1IyDZ8PGm7bDUYLy2F7hSIo
mgoYULMtViUwnNW0JEmnOx3SnLP5fc6Ln9S92ygA6tox4YV3asyfrVVxqJkrii1v
A1LKlMg3SCNrLoCg58Tr0DhFAbRodyIfRHLuuhOwt7JxfhP1uaQ6DdkFFzVRA3YT
hWM9aywEhUfoqux8Q2mFfqCUxvNhe8RrfUeJNVKnDuMmNqiNH1vJwZ6oUfqKO0Qv
FAE323OjacoxERQgtZmHZbhFdyEjT3B2SrrRaWDn7pPIeURsZproPL2H0goYVjiF
8SJJ01m06g3TEvaytOsDJ+j9CnYbSwGK4jiTTGr+4oNVCmlq83t8+89dOTFS9mPe
TSM3L+/og4Abk90Dn+EFGC3Q3bJix8xUWnN68ZDzquooXuUQywlc9W+a7VfLXisn
GJNfQw8KEAFwtTUZdzBbweLuBMknTO9Wu91FiVOjwfeU1qlUsZQfb8erUwLAXexK
Fn2R6l6ZZojdua9Jvj17+eGSnmqjP8bEsKPR2vjFiHjdLvj1c+wqyWmw2mwH12eh
JH/o4Xcbzr0RPyFiL8ngz1xlPT5dUfoMRHBDfltRuu8t4H8yk5SA81cdFHQtUSfY
E26OtpaxRmwn97er8FD/qVcoy1BDoP6j4G7nS8wAeZBGLEL1j59s73x7H6T7DlC9
HYrAidqfNKwLLAbFMK09V6pXrprAMBGroy9jOJ3PUUGPz7GmU1q7Zw3JY1Jxm6is
ZLMpv7BzW7/pXFsEbLmwjMgD/DxQdmkjdM3a0DymArwA8oV1cmqJioyMDiy7rTTJ
xHMEmgBQ61MFRJVkxDADzyIR0W6XSE8AYHc7g7R465vOMHUZK8KGxyZ0KezJ6kIe
RznmprivmVSn0GteMSfR2Td9WwybtVgXYuCyzUOyiesL3jELGCjh/zw0STqH66rF
5uy9LoW4NTVC/NZarNr1JJCLeeHXwP3CU04TB1GuucLkQhUk9Kt1BNkTc44j6wAY
lsRdC2CaR1ip76nJ7RDZpZPib/Ey7GLL4CNVUbc/rVJbCBYWDyUbtBiy2kdEfkVP
kGQvgJQfh89Y8t9owhYx3atKrOgnDI6f+87LcL6EXZqJW7CE0+AolNK8bWrn7BKw
bPHJVAg+Jku4bPAV5WN7GPq2Yy8BI0HNE39Mf5/Kp2BgOPsWtGK4kj1xvYKooHkO
m6f9BqRxfvSdCWG6oxBURii5GPP5srD18R221NjPLlriuX0b3H1XpmZIdwKvHQFb
2AJreCpUZZYMYAdYNXihI8hYB9QcLoDZjaaohZANaKQ1VMV8f+ft89Hdu0Zwy6Dn
gqP0YRR2pbG2NytmCPnxciae1d8os1pnpUHTcm6IgdhUQHa3bK4hKfepR8/kVROR
lQzgf2Ln+IBa+cRjCyUsp4RHgB/CzWD6FjOng4sYLV120xeb655lLaWNOjJQIXI6
00IvC1ZWakwYIy8RJNG5bzluoF2vKB0n8ogQWFeE1lSOHVbVohEcpEOTa++zgo3/
FXohZLYMErurHqnZ1G74A0GT95CWufaf61cA2zCo2lKpLWfmOElb50+oRX/PagPv
/t8mdHJ9HfM7q9SrwDTynByNK+ELZXYG3GyT036njbJtDAxiXJ4hJRviI458nOeF
U3M1KEQyCY66/qwBuaRoymLf4G7Pd0FuvulcjkXQFmEGpusL7mWHO8/bzXLtLfcT
Vq3Cwb5tV/6PB5noX9e2/kgGqLNlCaX9fbS2UHGR3q1twAAntOwcF6UuJjQZXDWY
9UKkOp3r7+00v1WXKzhF8ydMYEl8skuHhH7xmxMQ3KjxQKhxrg9HweshR9JGtLj9
z9WRPB3JRBdJTrbPoqZ4ySulXDGMbguHBD2X5f+z1iCigFbAseD/Alr77iUGxFtE
9FQR324derfFQ4uXO6R2etOShBUFwzznH1V/XRLr8xxEaXNxdOWBrHY/cGaEkhNw
ySgj+RAJ7d3n4RCv1j7twVYTcPyakucxIBpuT8pHblyJFJyPdm3aF/66ZrDe234A
i0rGBtDn1CBXXTodwlH3DpNFPyG/2xsxuRjJosbxFAbbsCb5FOh7BJfV2X3B4uY1
OuNPcSLC5+2az5cjS+SXevF9t/hnqFOuXAgRz1T3UgqRWA/zQCbtyxKpglXjQIvG
lDUYAbj6Xcs/E+kSB/JtV9U1k1I29v10dIejNnfwgI7Duje7dOHk6tCD8pR68bsv
p0xnSabzKs3lN02QMU9RZrA1sCmJfRzyiaOybJ1ov/PNzUVbsdqQim/e8e7h+BiZ
cnrtg3O0ou1sXpaP48TIm5VF+upay2dBJmGWMLHWHUSaaFyth71Br8LtAGxArYnh
HNh5nAweFsuMw0klGmcI0XBKEOgAFKA7worrFllmeg+cvmaOIfxrIgIKnK6xzsXS
TlVo2EKHQFL8V/7haOb9CR0T6n3F75vdA73rj6nNMobTTHgoadcRQL502obHo0I4
ObKPzducBe68akDtJ37r3av7kUrH1myCC3KK4EYVv8iO3DfBPRCNBDU0VSChfQJN
LZ1JUTdGuFFeHiBeLiuDWjE6WdFBfaFPSE+Qn4A1FJu3rvn3D8weNYmCmqdH/M0n
4sRbaWcBm6VccEzQVOaXJhqMPVjzPNT9UI3h2Qj1k9zjVabk84n3kECRd50wnlCb
RQNmZzC277GURCDtbImXVKa3e9OW/IEX/ophj9peqd+w9UjlPqZDQtIEEydJqser
0pTC/vNy+C/CHvfntdcaZXllsbpCiKllyYe72aHUyjFzjfmXJgZlPgFANdfzmLh8
2FOrKTM4dGWpxnmpur6robUdq5dYaUkAzV3W1GN/pjYZ0CBD6jvOvTTnDWYwGd/J
d4GMOyCpjmFHiJiJytijbQsjOpQu4RAz/cdjZuczlYcKvtEHiKEmFYdfg2CSXc/I
qKMDwIQcO20j4ZSdWxA/QofHdhMx0MvOEAdTEefmkZ9tN6IiobrsFK6Iurjy+x+Q
y1tD8Ovf/tri5zv/6VkcIBrzYv/Hq7nZwZjSDSbxdnOUC4fLiKPyZinukxaT3Y0j
XDd5EBsHBNgKiqjrte411dXms/euaFsyCAIq5fYVNOQgsHmC3MqTaSfPEDLaPHNL
iTrcl1W8VUew0Vm5cCi1NdOFnsSovjUR4u5BrT62Qeb7eHWt0voQB5mqnH3AET4B
dTjsnhb1nTW3SfkSHTHTeFf386weIn+kBBMpVYIgzAN0dflQ3KerzkFhlu/XlKdz
O3vUNeLg7mGBwK+guErz4t1bFJ6P9FB7hf2860OLFukTB9CW2c2Q4ZFWyC0mKQeq
J9okCChvFUUQB+2vCoQufwO0YWStSgtJOiUlxskpwbN0OnpokHMZqih1EEFFvxoy
GTc2HMghxnPvBmRZx4lW+0xwuxwHcfulXz0U/CoaEprfrlTUm1YXfMAt88Lcq5Dr
weWaFRKbfszrtiXiitA6vi8zio/zxugeBHpjdy1nYJ0tPGEDpowmRiw3vt/zCRLo
WFEfXhnWztIGb/H9gA9I+Ibd65loKXEvow0q8S5tB+Folv/s6ko2aYCGt1JaVtjh
0SmOWW11sN7NPN6B7LO19NuzgITYn3sA3liedTAvfzBumqSSyeUPf/hlsih6GVBY
iJnNMtFtYNq67C+CIwyhRKjIj/xEtocxGp+EyKYy0wpFkZsqvBud8adEUSn7S7az
9tycOI901VDcep1Dz9oLJhY6ZtXwdcaktem9+g3/MmqoQJIBecBqRCVDn1FdtWup
YwsXKFMcYjbq++g4yu5ShgplS/4pAF/M2dGnLheAxI5nqvilDUnYtZ5lbSO+yCWk
tkI0UeycVN4T82tJg2IccmrCPX/qaWI9HN4oxMiOxWg8nhwbpaRpWrk4TGXQ4vQs
gGxvgXHXhP2XdqbHlszdD+jBXcR4occO+Cphv65aaObn4jKeyITPwJTGyajKbP9o
Iyes96AwY/6lNTgQZvHUc+Ns4fwjuMiFFvPsMGxB9I6BpyOobIcmNte8zaf9Fqi4
kJTBYQN7uyyzr3vcWvSpfE1TSWkPpHO0YxNqkSfhZ9JPz8VBlKVJW9HepPpHVoiL
pn1H2yKnt8zjnTssoxr1DaAdrH+R4mCzCoiJ8WjEG9roqcQTRr3/g1erjnMurIDd
JjXhPfuyo97yHt+WIGwbOmgY8P8kcjHshspOUX4XElfCaKdYC4Aly+wV4rNCPQbG
iG3oLocLmxwb4Z8dPr5z9A18YoQTBtuayplH1wa+l9kHl6kM+A2g50RCxr4XerTA
kangtafyCF+tO4sGHCcJsEvYzCxeHESGozMO0LaRZdjHNNutq4jjoxaLHlAuv0M/
ZXDzQ9olA24lCbqNAzBfSpz6tl37IvD+tjjxGnk2Z8Ni65KRegwI5+YVg6JRZAYq
qUizwiMCRV83w5ubp/p3DfvqhUOj6dBEw5wKmTKWyAKpM3atY5MVUTbTOKzWLkYg
MMZ/SqWMgX6B3diPZPt/LOoptb8wY+PPTi/dLFTJkqadr5qN1XTTjNeg/H+wXgE0
Grt9CknJ2XOlpHVhZbhZ3cRu+E1ZUBXZGeSh+MHtod7ON3zk7JTSSGGX4O4/VPu7
d1YfUdqVsUVO8iix6ATEk01DR/7dLiCDUwIq68b0nIOifnOi2eXejkiNsyezldnq
v492MROmfjrpc52f8pj8FSgvgTfRElVXSu6vB/IF08TYoBSvtYcv9k0gVlHv/Rzv
2COJSrK93xtD+CfmLLQqS0TiSeomGrmq99xUNqqOV1bK4mN1/sE3bulPrp1MnloO
0PgU3Lt/ZuKV0iMpz19+kYHNxxxhYG68aesK/n0LQpiSXm4WnjkIxk8QvuA5WpvQ
RgPJfMY8RH8f07XOq769Xn22OnjRbh4u84K0+VTYu/klTXI5mnQdBmgn7+SPspNd
369NkwFX2lhVeiX2UFakPmVbOk7qNs8Gtu7zFRbG30vxBblHGJXzOOK8Yudt5YDE
igRhRQuv9o3KR7pgY43+xvvkJGA9UvHGYghiUQiZSGFwdhS+BuNpc14z25Iq5Tno
eqfrMa+Ps/aGgPHF9qRZeJNOsgRVWNk+bVxJRs99XQLktIHnNYX/hflZmvlGQDRU
nqkiX3Qy6yPAI5CHIxfVoQ+HO5Pl8UgrJS+WV88PhQQbC/k8FzZstbUxdF+q2xKu
IseJJOdRfOiPz3ylKIeSTYnGu56LFxDt8twdXJPRMHjHQCKs/kedN/8f5rX/4J6F
hnE1+Z4mUJLm4tsQ1v8ywxYp/4kuJ+pWfuAGQMqBZtKthi2t0ywGFQW7knin6Dm+
+7y9TLdKojAX6+Y/OpRjFw89DfAiVzOPbkF0K2cGrvFtkIFLT9Y+6nF968fnqy0N
E/6CjHAqrNkzhCATyCn6bpsIXInYRiCw3Yaur+SvK5Jc0xRD7XYEPPCBx4YITe7V
92tg4mlUIoAqLMb8xpCtf06YjHSYvjY55a8hOyQpFFpRoyfIomogHII4549g1ho4
JxcQhccXlsMZPeCxv4Ax0yI06GUwRHXYtUmPnmy4My82bJ5rSTGS9xVLwE0EdefD
pIn0NqflEHqxiYmq5AZMZ9mCaq+4rmop59M1IcAHjBaw8MHN7SFn9pfqGVUy7FTA
aq9uAMZ8Mj/NhY37DDA7nBDxPValbqQ6xOcak+PypTo9+NzUzUjDqJllaTiIwV2o
OS/HwfEvTUPw3PJkKVZHsQxLDS0OvlzLG6LNL7Pil98wrqXjsqq7L9OH0pzi+Hb5
8x6+81/yIfSbd9CBy0so0tV0BVOVHeyvTwXBt/X6aXuZmLYYNC3GENaETSBUrY3q
BMXlSlvTQklT/IzgNNPlSdLU9jB3tAl/GUuSta9aLTcdWKrFNwA/JJQRmb0ehQQl
6Wk3k7F96KR9ZXbrQfqID8S6tqz5Clnj6SYpLM9pbsFiGwdxBfk8yhpeXZuL4CD6
Jj7xiO2OAzheId/6TRDxO/irlvkD610hsh/3csOd6EDji6YAVIwHoLkfrZNNQPzq
OvjN9dWLeuwGXHbvyAsX79wm5fNv/nFFF5lspjwU0XbrYpYvaM7KbYPDVBqNEuyS
TxoxRjdlQiR/eWt6CHsqW3sGeu+NQY+1II1spGdKXzWJ8vhIcD/Cu4upNJwKP4FF
ESm0Ka1JQkYBr/15tkTdjiQkuzGMIEhzflptRbz6x4Dp74RCHUQsPkbzHqqHeeMO
3gnhNWxfbD6kbxkyiWHYnxrmBaEHHIQv4SWnitd+YpaUonfTpV898ynUv/S5azp0
g9PTnzFb59jZiSNJcVUovCTmwRvzKPkD1zBvXp/X48Bgr0euKI0dC7G9wwc1UCug
5bWSAteqAeRwPedtdYHYKUmw3KAriCgWQTxTMD++0Yo/xoVuTonZDb1DkjnYwnO9
CWnUF8m5YjVOoFLhDCpkwHWwd0Hag/Y/SvzEKgvoxIDMawep8wvAeQei+yFifzEm
vxNGWZ6JH8HL5/H9QCt9wqb6OV5IVR9R/ibjz9QP4TBX/+EyBCYHX696l08/vvAm
22sxIsYpY2lOf2uJCgrhgwGxRjm8F7KtUfIh9kXcrz1BIjnDJWJF2OfchvMbsDMB
/ZTy2wPpkFMAuBrfXZPv5dzXEgNJ+s3aG3NycdB0SrqeCb3+somU/Mw/XZJaIaQv
WJY90LANlkor3Mt/XplXcfjqxxMw4atxtFIsE8w0Dy9NuhGKF7iLeAssYuAqX9XA
OzePzIJM1TSOKFDXSnKCKfzVx821Pa56q0k3DrtMJlZC63l0JDYWRW2tioP4/AUe
SKIzNaYm39yRoSMEBbDXTsDQPmTSuZeVphzZ3bbK4XynzFObDcovV86DD6F/bvj5
NkhmfLIZ/yd9SM1o1oESWYfCnljjtLYe/cI4L0KFD6sLiLqXAwL6/bqY6K7M8NDb
FmFwLS9F6YXcHG5ZHT5rRZmQ+3cVnr5gS0DCC3GDeytqlgvvMaLEhmdlf0TZSjFr
IcGyUBrko2WYEcx56PqGyQFjsWm8QANIWPnsQyhM2tg2Q/43xi6updeBhFcvQttQ
EXRu0eLZ/nNBaLEEmZKlEz2zi3QkWhPjhZvA+J6GNJ5surVNWHTk34iIEDNXdomW
1pYwPFSAz/HTiQMJV/B09OMql5hHSDx7NkGhxt3NZd8iF9kyAfSYHuoeutDBjxy/
GcO1Y/K/SZfff0IYEqGc1m/o3RDejCDJejcZxnhexlxjk67Thv4TbQmKezsd6025
jz93BHgs7Q7Uug1NIVyE5SefyJNJOVwv+32yVKgTM7439fghR8Hwg5B0Eke6rIEC
8HqyfWK4tLgksJB8w2ac+0KH5mher2vcal+cXmx+9XMt1kV0LPkFhN7z2z5GA+EO
fT8PRx/G7y+MGqd4QA2ChyputelUDgmBsnmu0lF+yvHRPzArBaMOhhsMUQxdI/lG
P0auTRVuGaovDf4IASZf21myR1Iq47qlcGTfNYdwvAA5szzjT6H102iSMmlNiNId
ZEHY3cDgXfx6MLAsmaneKxSt5AMRCf0JYtubp2JnPy4BeeokYRCbWqWqQFMtKMX5
KyabVObd/JiqXWHtVaWCHdYu40C66TWa8ybMKc4dExUr47744bsOdCFwXjBBgPRf
Wc+eucWwax8QE6OIeZlKIiDzmAEr/mWKwL+3aPRir+zk9v9CtKtKE1cb6Qnjo7QI
ChoXLZCKi2OGaVbB2RExve0++cIRnX+58WVUOQ+zj/1U6iiXFG0EuFOlsAf0kP58
ERmSTCJ/pr9q9+Vljpc212xjU+HByRj45xpSRrLRpJxzpYeS24ywqG6xw09jSLrG
MtxOeCCj0czjNOQFCLYQWcLelmPzHOVmfvFg0QnltRH7TvOJAoS4WFpWQ1D8VkNn
nFZGp7hwM3sOvfMYFtWbBMJ9WywW7CHTMfS+p3LumlG1sQwasKtdldK9wl1vhF81
C9sUMVuf/1fCh7iPoprpyAgc9fZAqkzGtcQgRgU7QZyzy/FHQDi0P46nyFMUak5O
l0npy5N4+++VEHeZ8jGRURq+AoxR51aZ2d6R0kr5SEGBMKsCYlrs8sxZ1yzeE0yy
i9qtpF1/tQo+F3VMe6qCdY2heWPjBHN+rMIxzVXkpuNqY0dw661RJwv082RD8Khv
dCBAdXbIgmUbxOoJXsFjEC4YCGfY7Mv1sgL0aYvwK4V478EN1Hc4XZpO6JLZa1Io
ZhVWHWWQqX2xQyo5fPkx1yyyNduUnNp7B6IfalA5GIL6H/JtsBD1VmbhfdrebNYc
j4QFkYGrkJQEmZFZ8WoM9nHld6x7vEIufmkMb3FctaGhrvx5LjWz717rDUGvtmrS
alVw8jUvnPLTamdFYtB2tzK8IIOj4oU0Q2uqp35dNrXwAh8rSAeW5ELPVCJzswMB
KGIbpVcCiBTOiqJeiT3pUJSqEVXk49zeXufdbNv9lGuv366X23tWyxqNDzN8X/Jq
Rw5jP+entRHIQ++iiyI4Y+Azl2rtSWovqP6YIzmJ/UtcC4A7iVFyy7zDQCAgfISu
zooQWpdEMuzJFOg2e75XHeFAsTt7nqwxFKe5fqMk2Tku3KyBb2kz26HkxHTsUl5A
LwCxu9volC07dgAqD6ZccLJVsd7Y1rzGmQ2CBKe3o5r/6VLgfAaYsUbE5aeCWBne
mncfhzTPUr1+3zSJufwaSoiBEJE9xXxNxPUTTa4yjSdn+gk0vnYnQSrvQIns4PSI
0A9Tpznqguo+GavM+h6P8Kf7l2/aiKsld6UGw7MjCEKap73pyn6aStCRHEkUbquO
U3kKA/7Ar5Lbjekl3Te3Dxjt9xoNqlQWDxsyq2/khTPTEEN/I94iBCx3f2QNfrVK
HkwCGer5s6eb0l88fWVImUvg2cbIl32SQ/WnIIxQi0QDRkD+NMxOjFduMzp07IZv
vbKieWtwq8q752LY5ksRA7hHF0usIxy6KZXP1r4JndG/dlPFIDpDwMxKEVJpt6KU
JiRmUfNRNB4R7+apePUn10DtvePWiXK5QBPdg7aHGG1KmHyNGqNoRpLxxUkSIHvO
qavcL8d0Ehfk86EGFfkhVDtGcyT7H3DfEVAXv6w6jixyINeg9QFuzIFRV5tJlmc3
4RwrX4gsoskro7ldXPKoYN248udo+xS/va+19QAFlnwzlmFxTHD4s1gyujlIQC4y
l+hj8BK86hETPNMmWtaN6OtNFhNZCCMXNy7HhxJPfgFNSSmmxwaZBZVgmfiw0jao
oGSiA6TjDS+v0ayLhXHlDuecY7wLja01QtgCbTWtnOwk5oum9XClQFBH4oPCqcdN
9mtHVazsBh+biiHQphAQ7vf1/2KJXkiSqBW1FhBlvMi1XCisLj4k/u9HLoQyNe8c
EUKrVHRPZyBRoMgDGaiHZDdHGAVyo6LHAQt9ASgzw5/cimakFpE0PLXBuG941wMx
yQ8aZAeWKe8vMTwRSIvs70G14jcSqTcQ4TTBr7RvS4YN0wzlpi6oMFQGKi80iu0w
fr7rFKziRrCnS8hqLltY9HlekRpFcaOuhWFZ3wIMg6Yvx4qsYrXl2V/iUiDZ5tzd
FsYURcA6FJlIH6hAFLDO7+ztKJ3XO8Hu9LXJscN7sXc6PpHBMxugXoRZzUcXweQT
wHxGCwM5r0q9TwT4PZLHUP3kZhY8LYO0XVSxTmzATAqhpS+rFTECQcMYZZ0cizNh
xckH1RnxeDk+LjX/smB1JFbIEg/Pxw1ClsRVHBCcAIU2NdzZEJKqEk5k+yIptFux
7rqCy5DwNgIsyjCxM0rCbtNQGGUvWnHq6mQgIsHDdgypip1gsOdKaIh4cj8KPAsj
zj1IeKojMWhBqBlLgWXdfERHU8v71yxRhgX6aeGg14iQMPgu26UQaUwlfoyD2904
ifAB37CqdhC38ud9VnAvfCOhaKI2sJm40bnRENfrM7qLiLaOq1+LHxeF/OVn3o5m
og7XemgaplTCZuitsTRCqk8eBb/PD9mwgkktHTxMb1t/Ho9vnuAxsuFotYRQxbf7
RndxphRukZHgKrVpIUHjHxZNfv7W8ySPXc56W3fRrz6jt2rGwag2CEu6XL7qQW2w
+1Mwl/VqKXy1U97DgosH/OMSWUNPOdhd481JOAxP3+HXDozt3K3uWKEOO6gFr+NC
hYKCGRc73nX6Cp04dSMoNo5ZRpxNivQruHqLyVHXUXV+mTuvPHse6OJDyPd008vc
fwflrrpYWOa7NKvd665ec22DOLbt0QYUMlPvZ5miJjQPMoycCET+ESgdKYx/vZUC
/PsNR6OLP5Opi9BEh+3ZjieJZLFrHH5S3eRs/CxtTJw/N0NMt2JP/yGo6to082j+
PfMKBzI4nlU/QeDTiUq6mLOh3LMXNrpifY9YybNmUaPN/lwBhBb1BWj5EWzgrJKC
BpAE1eDScxxd9+1PuYNkLW0/DTQOr8geLCWKjyzszF2yWzKEPuM0xNZOoCFM1Mve
Yi6yMzxXRuFlxzKlcBgCNx5d2D73N9vqE9GY7nyfQuWrpoUSUI4eLCqZ51dmxBSb
+CenrTJws6qptzH2UgIJkFJk28SXFoNcJDxCdEIr7EBV5E3gL6PZB4PCQkr+7JI0
CB9Jcun8uKzJb2fxq22Mf9gR0D4YlBCSMNFQ3EdkOIzmGBiW4RSfRHVtd8DgyRV6
STwbcD8I4atOZLx+NXAZYCf9ycxvgxWaTvvEqNqdexGuK+Eu/D0U2nE3dS+F7EXY
TBRCmGzpJZXP0k9s5eOtGRLgp451xQ42GYLbGkDqdvTb5ezPn2+1kL7cERk3k+wK
kZqmkrHFvxG5YrN9hzX0ccFZyCDzugEhKanMsCdsfW00IRKmCsZ5XbCepDUbYEoG
EAfDqZCybiPNOZxuEBx3aoWjjuECBJ4wONwlAUoVB5Kntpu1cgAi+rDwu+q/3yOl
VvQNUrD2tFBtDItYqhGDgPaR3+iKnbJ1/bWpR08hB5mzsQpdz10R4NUauSSUKkzx
hh7F0RQ/Yr0mEsz58qYJtCQKEqhRayM0bzbWdAJlCY98MEtNTbwyklUGrwGEtM2b
yUooJ3gmK92p5mLMChmb+Maao0O3B5+wUC9lUjvPZY5bEoWJmPyY9ABeDAA6qp7n
Sre55R7ZUB96TQXuhxhkcpDXK17t6Sapyrtnwb1C8iYcoRiRpK13qLG1CMOJcdZ0
8N2kByE52PPX6JLqzRSuxl9Fic9O8sdpX9PgxS/zqZsGmgRSOTPxx9ACq3apyjtY
qGXtGkW8Atm4y8qcFKuYo8szHpyX5Nx5mko49LxWAF6g1ju1VgxQVKsZ8tHxRyDV
2QdD7f3UEqgTHM9oh7QNtuSbcXLSU515T/XBZbD4PmlE7+oybhabmH/47jw6n+G4
kNWTx/ZIKh4hsfOPupuB25+zbDR3UskF3DjigdiWMOntrQOpcGgZOox/PSqW93S6
YeyKUypxKrOLY0lh35sEcNqZ91sOaBQFPyQiHoCecHM9ZBqU0r0bqA2E5thOzS1d
4i+hCzp4TbIHRBra4sRaqozRepGRZkG+FO2uCwC+J+lfPL4xskIwpQDc8msqBDnz
zBOlwBS3vX928PRDthwNzse+8BPK+a+tMacVC5U7fD58s6CCKVma0xMzpPLL8vq+
PfePiS+2QqN9vE7COFgufQWOi4ZSQ0L05zwjciv0v48wJnwtlL3y80zZ0wICYMoY
rfrXwjGBOhkdy0iEw7Kn9UmtXjM+61Ve3l37jz9Lw953bKUbfm5/+IkP94AhRx2P
h5T2raRy9WDLW42hklIg37heaWOOb9P/dROZoTbjkpiA5XO8G6WL7Z1FbwMUpunn
0nBFpKwSuu8e2+GNreZUeKDTwLuRQm/hBCLke2RRWiBHwew80uXoQMvX7OqsMkBZ
2zp7XHYBr4BDemKJc8AASFQrqRC79F9weC7SZip0be9ivjSHeLcPD3p7gKBeacOB
Jws0JZyADtv8GE9zYWm5tztK2EXtjNIFjLvX190EyWVfo38KxZqGtnKZ0WJDCEAF
5O6TvK9SFlEg4ytqm6g09I3UndDHrU4qEPqfeFkkctkN1DAmLXI7KclMDIVQSMMa
MJJ1KxLl8R4LKID3PVfUXAV70wfRQdwfIPX09/tEdSIq9R2Glw4oz8CvfWgRSOsH
15PAWz7URSGXV/ryMn5Zi50l1Y+VG0IOz5lrNnxOdhoLtS9N7YxnlhdsrK2hoOPo
FjDVcM28NDzRHd5BImpJMPZqcoa/k5BCAiR3x9zFHT81LLVVnu/HPzWybcDvgAFq
8Q2ht0rT1AUbfQ1aXBt7511Eht7g/B35CQsBPJgVLddjy7pTu6meHdjKOPRqVCW5
52ELFLryULCK1eyuAWg7AKM3ahAerfh1gTycKMsI3+rceHuUgzhAPaFHCxho1Yp3
2MeiiQWIrm0CqZUspS0JZB6HvSNIgUmazpRTB6DEtbCgHBzjkrGVU/+XCIAbUAnt
+JCCg9/Sg5IalTCog+yHEaGZWjR3dYf7VIpIDLg7l96cOxpvD1c1YsBUzMC8zx9K
j/s2rhkEGA/cUmYwJGAX0R9tR4nYM7uETynkcSSy5ILrdhed34E3Cbi13baxiZW/
jlekycAcSPlnRT7Ajkn56pdvIKDOOzxCc2udQV4FcWuf8yQLrIMAKQQbaNo/WifN
pCXPnyCqE7o2Nv0Fw+DuXrg/rXPqndctxXQUdSTu5Ls2o7Mn8hK3bZf6NNvKfC2v
rk4vt5xrYa2Nm8L+RSk+SD8BgDTK+62r9xhqjQ3aqD5Eytf8GmqhSUDRjqdVphqM
RIvtvVwGFw17P/4A02h2MHUQtj7X64ddDK64CgPNa1/QsckJDx5B1E8DlpXt592t
qAjtScUKV9KuXkw8aNdQth0iQ/QMVsJQH+PUL6mqvMIB5BgliBw2//cWlCsGBRUr
p5jbQMbUfhdS+LsBZfPIIszkcz0Z/i9lBxnEj8oGP1a7bYO2zAmG/R5SQ390E3qe
WbGtVTJhYPRnuCM1KRUMan2BbQD+TyYGH6LlEZVkN+8Cgb1TQnWxcAU+FvqpSG5M
BDfeP3Ptp1TGGT2ie7pJOUU9KZVyHmPH1vRRNsuICYtZ6Ll4SsTNl+jJNzl7tZWq
xoqcfSO866bDhr3mw/u010BeHqVFWh3SLyst/JXx19KMJY4VWseuYFQMOAT1f9QS
ZeHZWt+SzKD2bYCm6kgW/bfxHLAMf55q+rlC5xBzKuJztp8O2n7WHHE1zI7UFCAe
d2qKzGEvVfhjrv864xhYtlPW38PFvDhm0X3OyGrlRYUEgSYShAcUUnznwmggLeFF
5GTJOAYy8qnIw6TotndnaYc0/IxfUqu5SUgIVkNN6ys8xVZLUhrHi72dbCyIdb0h
liOpxv/ojrS9sBj4V2ha87zx90Ra2qp83phr7mvTQK4xVmw6XdXIikXmgXjYIl/p
HbF/pIXIShtnvmma/Y2AXkqKE/zaZaxxCnjzcKLgfsxSJdv6lSM8sWOzrinFYFU1
Np3QTfTHIfsrQqzd9YYykMGg+LWXt3ig/+FTRJgTJ0wV9vbGtaaOC/IEPhyVOLFn
GIqR/e/5sXvf8+/+0BBDiwRERVDL0KFFF7FAcxpEm04bdgssO9qvRKjsCDbYjp8x
EIwMpS68pFbAwGj48Cb6Mgc34iGuGXcSNSXgEmJFidcFnlECyo/IG9flKO1hY3aV
oiv6nxoV3EkNYlOX7MseBlSmfmzmxu9dx8WHehFu2sLin4T8TwZvLX0SYJ4IxEhd
LaP+INkcxhJZ7homoTTz3UG13zQHbl4Y0ffWxIymKZKAouXonszbpQKx1vL7X0TY
+VrxNluhHlU68fH9YR+xc0Mi9gMxS1hgKqeZZtieeXAmjQriyTs4tsjNfcJh2jZX
XHnnHTqo5RAja6k3DJGH2sqKk9/JwTDhkDLL9eFqTVm1128QWWiRqVJfpnUnbjJ3
VvF7h35ZDQwRNDXy3wTM+ggSlXX/xvnsfjpr9IUbLjT/z2lLWYX3CvpZy/rCKj92
8IU+I1ZE7nV/FD2qTH14mDTUAKo+HzOSW/qieL/KrMDGE+tJqPk2LLB5ofj9SQel
jP3R+6aSJbDkPtNQSXpA+zeVGZiu3qIAh4Wlg7P3Sl3onLDy0U5rlVmfjDYgu3ZV
gcEDyrqjwymU3GFIVzBnntinaR2UJtBycO8EEp/TUBLWxZvU1ddsh9w56DsxiCEQ
HvqsAhmBfTqKTsddiUX4WWf28/hCke7txtfR3jLY0BxYDTlK1bzckvpVPcrckrDw
IHc8gn6nMIIhf7qopwDB7zQ9UzeZwMtGGif/igbLagCiRa1AqDd1VI1X9UxDdjz9
/x6nQ7gspPskzkve6FHwqZ0u2KjSRoF24BZZWetx2DghsZ96uE4M4+gWO/sshsCR
4mL7dSELZvLbsh46HEsWHya7/3X153OEciQEYVnBruFW/bE5WJvceLxOWd/9BzU2
8ifBofncNWeNOZ4PN4b7XNy5kIC9MHy4JSWUeXrX/OSpOTLvnyAvxWNbnTcq1Weg
yxNF/T2aZt1+owVcvaqaBc+gzJZncDNck6c62JS0Ow6RJbV+6h+xqhLoMfD7IRad
sIzGlaX26TBlBJBVeQ0JSCKatquW8FGOUhbPd5Ko6T5RT1Ic8ImpjzQqzVkA2zyq
KguvEfmGktrIzsxvvNzBPyzp+449YLQc862UuWhF70EyiiCbJQKMaGgxOC8A4uim
fkDfsKPLjVOR5drilohOXkjtOWGnIL4hnvJicJ/FLlG5F86DcbyHEDIErqvUQvMZ
Hl4B+FNDGgNR47NllgOwefEqA2amvkvGHQYruF8m88QFASxii+AOi2z4XUdeWtTw
qXIOpRrsWnw2enGFuIVk5WB+bA6NE/uUXfelDponhLhk9WbRPz8JPBFFrepGw7lL
8Gegtr9Fa0vjieLq5zrLw4qqMVGw7z3faLp94MdBsGxo8pNypEqtX12JakkIQkmc
cFmZu7hrD729Q0mkJsOQaVIXd+g1PN2J52faHZ3D937W4dIMHEfZY9SNnT+Kb5FI
J3viOFaTISLw9K6dC3ANF0Uc6CFU58y0blmOHi/ynh2JLhkDaVapKViRQ2GPzXnA
v/sZvb5NHFBo1gRIcCwNoosQSCohY/0ri1jczVgkqCg5hEK9iVzGxm28yK/pZv6D
pa/Fb0cRhskxE0icAnVXqomp0f6O+lgmzeL55GT9/rpUcE9zZyXJa1YTzDz3zaHm
Cy91niadyl8ehVtjbMdbnp4jcHSEwQQmE8pDYRUn1CbjVHM0w4LRLZxv/P3ftTgM
yG6fB5/utgzhrhQp9Zuj3QisDs+9P5XJcFZ7+d5p3/XUweInAkvmYEjudhnvVIk4
eTBypge7n8gNUq2QvvDrJbJ8YtfoEICrYwYTprNWEbxJyEtm4ZzE1gCqPM00Ov8K
eFqCNs8QiIWOsUvFn9ZUrpwidAJtYyWW+trkRKds1hMpbufiM3b7kqlxqH5Vg//A
0YI35VA4yGLQNfWrouIO+YIE9/YEeUJNSPJqX2o+dwx9fzSstf2dgie0K5h7wYNJ
UbBkdpBW7wShiE7q4TNnFlws+/rIaj6eNmzknfPkqjBKoRo1+dMbiFCvtrBPPCt6
r15uVXw/8/NY7SM2co96LBgrpRRv6BxxmF1wl1jitU1TFmFjugz0S/tY0516Hvui
WJOh2k1yVC7aXrafhU1sZB5tAJtvFbwK2ZtmiaGj0N4tyJ3K+IXiOBrFuLco7DFp
6bg1IkCTiasoTc/5/vzQuspRckMOI5sleoeQb+A8N4ixdbfqzRiHhA5a6Q9rwiAu
FK4AKYTHDfzFSJTsKLf0fb5rXuKwIs0O6tAnfDJ0ecnmSBY1ptOXDmDLbldDspIp
q0SU2SX5AmlJqg5/knXdQ7b7IqmLGBvhEYdwC+orXJuHNuxsTbbV5vNTfLdJEKox
ivpBn1GZ1M4T+2P8P6dFM15a8HgAAn7tXni6n99vY/hyAYZLISfqYEiVLXvlZSi/
D2HhU4vcnOkPlgj9+mG5omLrx7XSOWg+ZacB1PpijBOEuCwvwmls921eb8SmAI9Y
cH1zttMHwEVqwtjpQQGDSc82HTfn2MnmbvTPCUnPhAj0sbALi9XaJryD+TBvZXmt
PgKgjDRkpI4H66khmUZPW0/umx32CKahcwJZsvSEsWwQ5rovNPuUe0UKh8kp9Las
Ec4EPcD7iT5RPN2fQCs5WxrHPwsJsyebttXCjAQYkcXt1+3OC2UKrbXI6WaX/V1e
CmlGzK/Xefk1j8OmP7IGnSjARpH/6CKnjuexHdd0469XuSrMrWI/799DvpBROKLV
qF43E93Db7AoDalFFCvrPu5Uh+TkCujiPdwW1Y2t4W8PmGXgGw4e8KzDT4Pvq0Lt
IChV31xJJaFULOtM1fHUXuyWhRRxL8tkldhbLANNO5LYlKhXCnj0oo7p4VqtIbLw
TVEkC68hRI59XHRDfNLw0LncIWuuAdwyDUvpTVl9kgaSneSRHt5YPHEf8BTJqj5f
oe1jnLJip45w/KYxe8NBpk73KOAjx7esNoq/234RWZfzZwWLbUIp0158mRbnr/Uu
a3XUKbXbRMtWuikvpgEr3opeYOwN0/CwBpymq1tZnTXo/7Aeu12hZPOYpFVN5L2w
q3XRHuN5ESNA83tD/66U+nNZzBybeZl+inG+R0v7nGDJwGbImuAaGeiB1wmskvwZ
RrCbhvYnd9vvoMBzZyVm2fvR2MoejRk5Iz/WuM0M/CgVkITNLKHWysC8xAu9wYrT
qXcFQjmx6krQXmpy+tdJ0ISWckFURB/daE5PZ2kZCba53133NhbRvWLt+y8wSuFh
DSIa2GjgLnmFwEtUUiOcSImUtTDfFqCK2xijb3T2nRHJjXEqi28B0SaRt7f8XxOI
DWg2ViKPnKZO+6N2/jkdMVJ56ploz5F9thkhHx6NwUoBycoyGy/9Z3CweQj3fnE4
2+iOOxEnrRxaHLxWdbTbTFeA9cCyc29syKsNpuVCKtoU53axWqUr/yreT5MfCXk/
BpnAs4uDoDPqutnN+j9KsswZhrENM/nj/6WwPpe916JKGw66oI6VypMTVJa+bizl
hz6Zp25mPCkh0FoQDhF9/kTSSTjSo4FIAzCvdQirNSAjdLycwF73a8fBfR0OhIHd
+SC7KKnUQI2cbGxQe9A4ZmuwjMbG93oT6EputJHM3tgzHeneixh1Qr0D4NDb7FhM
IXmEP3I1zXVq8o0hKWM0Rn06B68G0A2npIQaX3ZwJqi1v/+RbPUgwMs8YmQ4hcRS
r9KG+cHyodIbHyzZedzvVEbfKiwOwykkkwetQavK8R+0XlSAgTTTE39u5FLxd6ik
zB+qQyz/DSN0x22mjs8WF9fdVVHdFpg26p1DIjayRrQ3SC5a+lQAfwDt1A2fBxoR
MqBTeo3H45XbMSBkmsRpX7vv3GMdbxn1SfeXIR86JR1GCB14rs/kI9aBhSmosjRM
w7h7l+66srF3lbLrh6sfvMzR3xEnzymJsvGsWgaftgJZj/5CvpJHTPtvyd0y7SHj
czyiaZ3dijM58IVxOp/OQGhQg0z0uQ/tPemPVmlQ1jfp01Nx296H/NiwLyGq8smU
g2dkaY4hpt5rHVWkUhImnojG/cgpBHVFGf9sXPzcw4tnQi3Nm6zn0F67cA477BYy
j/EmLUiqc567Y6RcVAIaSPSEaYk5MAkUbQIFDy0RA47gwdaGs68EOFK+dy+3PMDr
eUvu//OEG5Qzh7wwtPio41aM2rFRrxoDpV+wJehhItpygrTaa1inHct9eLUd20ZR
hpFVx4s9CCe8ZiuaWyEvxCgCw2/7niKuySBf1nELGZJLJ5SfGYNO3mUoCgPWqodr
ikGMEMu370b1+lKRoN19lf0UUFPqt68WKwOa8xKbkY02g4gExY5xZt4WYYayp1mR
XUYjbNC2KrWYpnkCWCtyPymL6WCB2t4DYKloi5lwY2VVDIhZFWP/vmS2mirwmEhO
TdG3x3WvsFIfagGInYWRBGLx4NRf4SdB5Y4ZGlcnzetoeCgSGqWmy2Z0ogiM+2rl
83vRq1q0SNUdY6fOyHcA/R24W6/FdBwhlocIjC77nVQEJiBqKLFdllcAuojXJCcN
vCLmMGI8NmJzuulC1ns9jpEMZwkmbx3T6wzjLn8hzk6KSqUWTnegMYKeH1+Ba3j1
Bptz/WlhWdXj/s8UBql0lCh3zk+7mmlUu7e9qlOLmJ8L7MxtKAc46VD6i+coZB6K
P7EeT+gBbh/oQnx4E9xcd/lnO28mHXdw0h3CSNJyWAI3DWrGpKtidloFCvsTOm5B
q9s7MeyVX8lnIyR4O5ITc5GmtyUkextrQNPwKFIuMMNEEEyvPutR5WUc1smQH9gY
NhM8/S7kIltuuf3cBD6wNWiYGUAjYlvwFTw3+KIfPdGP4OFzPpOWshOesNM5MBoa
XoqxCNxlDdcS/SeOZ08Lm5WZeEyYQ9+DGm2fhtGKFFbZBWO+5+CLVhefuzBgwVdb
3Jlt3zixJ8ogoT/bEYas7F0UlY2HxBJMe+lIivR2Bju4bjwns83n1DAHJI9C3Xal
NxPkubK7kMWoL5LsefnNBjkccpFzI2sNCMM7ye60ZSRtdpbqTa9YD0HcjKp8wUQg
W0tK0aIGj7H+GFx/41R5tiTEBzZIqkwQfT3u3i3TPoEItckLpKCcqPJ4My0y6IS4
Ja/5oTbE4973JodtpXYUlkwN3FcirMtGTgQvg9EktVd8iQP03iZ9M+4Ad88A8NC9
Jzp2FWTDVaOfPo0rmjIHplrnFIUKPgs3ury4heeQfYmZxw16zl5etLFGQSZqFdFg
6vtOt9g/OGxH0u+m+5i+yj1gz3DAAqckAa64r7Pfl/X0h4BsTb0mcyISKOfnJKY8
zwh0Q++NtKnr1oKlrfctgC78Goepho1Jplk5mHXIyKr0OheIVRGun9ONYoP3MlA4
Z7M8ezG594HLi1TRATsuQvsmbNm/DICGOMyykUy0wbrKAzmIbGGkg5mTRA16mabB
M9AF/LCRe1DNymbCgBI3uxSlZlpB4MqYZvIZu41CRgQ3RMaOZIGw78p5TgdGSYJF
j34xwVh+X3GALl9UN2nsBrIyf2sLQ6WZzktKpa3Oi3R+l0y1UKRxktd1c4Itn3BY
XHir1/zSfWet/EZ2jEwJp/1OsSDqFdHKxdLj5gNPEqP6WZMIQ54dXqyeQ7NcZqK5
o6n1UgdxTEANe2l6z9XDGdpN5bWr6IFx8EtRYR5rhA2Zif9JvBjZQCMXvztKnsKp
ld4zZhYMAtNLje1f7K6tJzfZk8sSaFv7h0yTZlWMsaC4lXcZWNCuNf3ghxoD6Arj
ZHwY2auKVUqDuggBeug7YMOnHXWFQKOd5UwhB5kdIfuCVwQDbvrUyzaPxsCNty5l
4Vmn5jsoYnZiDtEalLkJG6YOdxeBLZ4JbRaOXlbKxwnqXvPzHu3pNn4V6R7Skxbq
ZtlNVHFcxK333rnzDGHRjDbGJcaCqxhV5hGHoZ1+v4N+FRVM6JwderQ2ZYpPvwgH
Eohw0ZkBZ58txy047OI95FnCXHJjOYUJ6W3nUbyhvy6rFeASF18325A+Ow61Hg1g
8DpzAyBzIJIbiv6PZjdQPsTk+UzRXPG004SGITbkzeYtUmJQdju0rDN8roKdtEAP
Hi8G7/QDUIHq9juTHCR7ll7qu9UkQ2Uk32xhwGqCs7ynNhGK8MrccVYD7KvbfdI0
qd4kO7su2N3Pvac9He8YYyrON6UGj3Yq/ZceDxaUGxuICg6wjYW3KOKPo4s2sM0U
A9eV7wfur/gQt3TzKLkK54VhKVQKTR2rhKAsb+43MQ+MnVuMZ/Bz47zfWGJ0cVfJ
tqK/DWceu8/iVvY/eLLY9+6xP0QuBFmJr5Bdh4wvU69v5BeXbVVMTspHG4IjIX/H
Ee1Bew4xOMAM8Cp49ht1z8+p4UIlTpcBsCIxflCCpo5LqczWXGwGr9e9y2y+uCGZ
E4TtEhpJVFKNs1UxMnMwzbxq1LE7p0lcCQHm2IVS0o8lg1dnBfXhkcOAlT4v66K1
fNK2X2oLhiRil5H0HI6vRLVYj8DuDq8tm1yN4IBIGVYw9hAGHi4x3VU43+GsrUww
fmG4gjwuv1V7V7l+V6n4Tc0LkohSas2DJVbxgzJFFRN87bYEOuJHXSa4AlJ/5pmk
a1mxN3srW7TtE3efXczggh2mdKg/uggKP6QMLZYPNSrG1mZON+jJGdr3ahwIfmHf
qDoy5vGaMg4CCgJo7SCGnNV+umqvh4TnqsHH5YGqL3qUNxpGEYtCmeNcG/G3YME2
sQiHKE9XZlxBGK7XazOIUk/Hx6Q+zYBjcvtZjDgmWNkbn/h0DK71nqTQu+9DYqxO
n8lhFq+wg2KAgcwkbywvvMXtfhk/1NL8SomWjxIvfp3vdDp6raabLMH5Q4GWGcAQ
rJatf74XaGXbUPZcK66jqXwIEMCMhrpl0Evd6+4WWl5iBSfz5T6mTB4oQb8/rovx
yCOCphE6y+AANKNrsJ/jaV7PP37CNTYz2N1hbaE/j6esagWfojwXQc8+HA0BtrYb
PKJFe8tY5wdxZVJqYkLLIeAusPesrrItns5iUjFTIcol437DyZGcmcHZykx0GU49
qZsSRjA7PdkfyFhTxRRm5RxgBnB0Tb3e5rMa6zjiZJKn24yxwSKeFlTVfovnhmTC
9vwzhAPouktvoAom6xwF03DNHBpjqHnrpEizfOJm54ewLUQiyqwO5DAhiTLRyn5D
FpH1h/uRfbgs68l8O7uH+qlvrwm1BWJAu4RxUn4BCAh6Qpj+NH5zq8snoho9XHwU
JKi5MB7nJpUp01nKXY2L7O2wfWgRUQRmXX7juHaH2jHd5YBVpDly8vulghE1Wplu
Lwm+5gk5g4VDhqR54wMQ/eIjvRGTwxb0Aq8FV23yKksCbQZszWxwOfXsQG6SCBl7
cQMznbIYkF6wUDRwKJfkGTxwwr5sVQTq8qpZ9E5el8s10lni6K+VwbZMOtSzSNak
KiwOYqpiJmh8dOn/+1L/epZSd0eJs8uaK/iXPuZfrjny65sLeC3lYPJNUjixF78M
RfiTYXI1iUoM8vThUk0LLGAHHcgdVqQ1gx6wW1TXLlcp39iPKXlwAVMGNMz1fd2R
seJi7XWFAVKb4hO5FR5BenFXWsabBH26o0wzrl03CAWcgGWZTg9RijrE8zuT5+Ae
0vk1Hf1mlZIDG34DmblntjaSng9DrJo0IoxXkbuMFkbs9RXrokfROz9XVYxfy3AX
HUsyUB1qrBswF6gD9f+QQQJAo89iSorMggSnurH9IfWl7ktr7ZPlGxo02i2pqqrL
QTCKIR4ygRSuQQvw09o1AlBe060ix3fk/VDMhglstjdZWAZEbDC3kNu9vSinLDtu
fLAeNjiufUJFkuWoyDFd0xVP4/RsmdIn/CIe8cblu29t332fniYtoTSwkRrwVjWv
Uhqkq9yZ9YyfpU+Zy1NZhqag/Uh4CrEyRnKGl3zOGJTHkv3t45jZUFci+nUysbjv
VnX/6wFofsaKifmNodxBOwBxcci5t1jFf+9odSOxDAtlsB7ijN+JZKkVJrN1BtiP
X299ydST0D1X0rMW97zByUSRmSvuEbMLmWUpOgzed3b122CMI+2c1m5Zri6UhrOQ
tTjvD0x9PISqa/n3g5NO/kZZyYq14yV52qvPnaZU9aEgxiUC9hsXEiP9rDf+9U3+
VQmUujNzObzc+tglmQrtI9YVhN7Qw2aZO0kTVRJiA7KumYxbdJWaS883FTF29p6F
aVLTcRj1RwXNMiEDxmtvZ5qoipgJPmLL8lcjam+V3M37zPD6pvr8qq66UA8v2wfe
eMWnI42x3T4ehfSrHwQjA5FQ6pv9eCNEVZabS6tKQWeU5OjzGQmGpUhVM1t//qs+
E52qlvc+VVHBguqOZO7+YwxbjXUluJm3UeAaVqfIfaTGs3/deTFKg9n+3mGAlmHT
UxN09fAAoziBVtTfJ0tnnajbo63r1TaB4EYU643hUt5uEl5sbQi9PefpcuEsRNSy
aTm9NPN8euOxhijUsfrEO0DLLDh5ZY0jrRTWzJaKabz+G7PUE6r24eB2ttaxcYPM
X9fK3Vq1uLcOuMZCBGviHSUwMhHV7QQ8XcrJDg815yuX36vCB18YsmqnHOkn2Yr0
6bjGzntZQLKSkC0hsWxWeEdliPiceEHiCGLm2KZmMvxd50FSi+BzBISqtunGj9xE
iZac31Hz/qWlQDBLVTO6MMKv0GVw0lOrqH3uvOjWZ/rR9+9xxgjNChXa7R2AbmT3
R/z7aSvTQYcv+jUyEM2oypMy/WsuqlEqis8utwLiGNdV12SMoWJhrwzxgtcLCeFF
31B3z91hdnEKJTJCbFp0rd/bMI48w+ymzN3CKuEspTIUFMYQi1TT8p62ZAxw6CzR
xygCU/ouk0i1QXSQmX2BFJfZkmmJpW0RzNwZJBPEXbTT9yU4kGL+dFuu/IaJQXnN
SNpOisSg008+D0zkWVKf6zuILp/OAwH0wK7GG/LjFempizvQ0PopcDNLTWhK9TVz
TgPDn2eXnX9uW+u3UfiI/zjE/0XbqbF2OdJdtGHkYHAzdk1XUrBYuZ74NqXo/bUa
PdbtvblXvuEJUrO82R3RW2uxeRLxLr53aOqw0fBTkLwu8Q72YQBghCp+5pZfuBmN
RfZVeH/dz3FpifWC/lFxlb6GP6ztHrX7sCd3v3KPhqWriBEHk5DqNkcxQkKuAIl0
4HGVpAbGTcF318HliLIJa8GSzs5Ai7gCowUb/nZUmspB8S/RghyamXKKmYGvP6dl
o6kLyMqztuEx9LAZGHkjEWlTvWylrR3PLAypX1VGocH51H5hIqoIuKYFo5S/TxOV
Ywfnoq3m9rxrf9i7ySX5B/J80LzoUVV2KVETh6AWwtmpU/Cp4kCvm2O838BsUzKw
7ovBXEG6N51+21M5aNCWOdZqHXulRdlmjzjjjVshwk0Iq8c8CNTbZNe5T7pP2qNy
eGhHeNmtxuhdxFPIYQg4MRE3QNBdbRWHpNeC9inZt9KLWwhCUy7sTFI8g4RF2MO5
q26l232GdXK8VXK5pED790Fq4OU6FohKxdgZ3RsZNVkzLJVlve3/Nx/E5XQOm6Tn
gVC42a/cqgGplolqOqU3VTdvimUTzbFgaKkRLh6KxiEYmyM+QUouW11KBs2B6LHb
JiR7kBY1ykR583rARJhNHhID5IMqV0/VVHi5WyxrgvRomd1FFHpG3uIfXwcQC9dB
1zVf5/C34oL7Cz/0rAB91QfXzelmmsjk5T63FgQ1eTIkSIROU9nJSo6POJvNRD90
xh0qbjIkTYL9QLZ3VtvJFsYUE6A5eYrFUBjKaDBoDNDcI2E8YWrHxjztEyuMd7p/
zce2LP+xM70j+XuxOt4qT+RbdzHJWdiATgAeHFjqEPg0v6aFzObOX2BXJCsa4H3J
1jP50ZR0QDH5ktDS6e5DUUFXOMB3aHdaMAwU8sYfK78I9gKqq3iker6Q4QDcULGi
htG65VEkvRyQgFLbPRcy7FH9OceqK5qCuWE09x6aXbhOtc3k299OJKUFNsJYf8SN
gGxxqSQDU40pkN30DpMwL11E8eR7n2HaL11kWX27S055+LOt0vOPptfcbLLmYaAQ
F6IkiIzOmCzHahH9GssgOuDIAQvodjvwMy2Lu2DpVl4c6EhwJslSO2SpJcgxpEJF
ZV9rRM0yETWN1fAWQUkm/TVF91KNZB5Lx46coItzUOmGUoRlnaqHTg6LcuLrApge
+z/kroy8wl4DMiSPFzS2gC5xH0+2keVz2UcziI4Ng2rPlz5xSOY9WNeVC14bbYni
LvensMEsrJMyrW6qPE0JIN1jijpT48053G7nuXk0h2n0O3UPO3YhGy6fT8yO1SkA
gd9aD0Rrsv1aysrsgCq6tsFepzLgckm7hBCmn56TH46Mwmg/ESgUbbkVx4ll9X1i
HChZSTvY9VE7ZEKi0DIiUHkk6Srt9qqGlxogvwL/EUWbVfZaOSNSgzAi1YeZ/C0z
ELHjUiVBsPTjX0zRTvN+SoSqCVt0xiHeMZ9Zh1WuJUlpbm5uqbmHfWjfioW0+8y6
R2FElVLgR/VZZEBNWbRicdI1yhSk/AcWE5A7GvGrG3wqqyyJWBZkZsa1tQP1n75a
aer9XpC6syqIsxKbA+VpR7arhIxz0Wh51KYjk5sv4GfTKLr2tNaIeH8Gt2H2cHTw
Qz5tv4QGant1075Gh4rnKzxtksiQO62LH85HWh/RvnT0Xv1c+/Kd0OJJka8aCdFw
rpz5I2GJ0BqZL8Es6IWzQr1AhwVjB/rxHuAmLLu1iuFGNhBJXw+fLKrtfOtISh4J
cze1vS6TOzjizeSdr7Uz8wPfNXa2+FWTbaPg1baraHNBzktgXR2ExLdUlaZqITZw
9Q7FyX1VaI2TKuc/OskuZNpfupzo8jMFu8HnAILkV70K/XGxZ2dmfiGxmgNAc+YM
iAShM8r1YMo84NTbl/ORpYC5GwRR1PXHU4leeLuqa6LwDFLsnmPQUCKbmWP4VjiE
i08Ms0IqEOK7SNo+Fn02PL4Sl1zV8vMhhX6c/V3w8/6hkGS/6YEVQX4olMPOiu2n
fM47uxmml4qFIVdy7kCEUnsRNPuAaqq6rDW9n+QFL+4p0M4QIaT/GlLLt3uLAzSI
F/3WgYQguNtsmD5MxS9QhR8GqkxsB1B7NXab1uRsP7/tSp3/W/+L43XOnz5A48mB
Rntsbg0Smm2lufmhP3M2DiWKDeArJp9pcXtEBbdabBWa778QRcjgAdDE8A0tzW9h
9rVjmcMagKF66YI8q2riYqEcZAl7xLtJ9hrrrNDRc6yzNEOINUQ9NAJXfinV017t
aczsm+VmSkuoUPr/UD/FbX+q9XmgtuUASW6IWbGK2tVqYfe8F7WqJte9DaJ9cm1/
N2koA0sMBowiOMOszIsL64nFxeCj3y9rRXLtrnJUx4072BFH+KKIQmj6D/hG7umj
0xYAZ4mLHBs9JbGT95XNpY89p6jfFarIyI5sEH0qlg7yl4admbSD+Jvhg4WmsqUV
C4AwVxQ1S0GXWtZyDzP3skX5M64DC7mkp0pKCndNeIu0rP3s+wW8hLot/HP0zJJX
nmj6fqYmtjspVWtrbtFhwQrEQyf7nBJjs4wuI2sx3zpaYSelgbYz91llZx1xWcAw
fzmwQG4YBGSwALgPJ4D09tLvOqYIUhafhvTfePMGJvz+GDzXQPpAS/ObSSqTRyWw
LjPI0uGbLyAaLGQLet5G8QjThXKdArQCJyd6ion8xadfTkrQPCR9Cz0x0xWJLMs7
7hi//vHvN00t8u/Vc4e77ue0JIJB2W8gvVHXfGDqmYIdtBnWiZkV8P7Ou8rfmyWf
7iBPKYv0kRELKCRfV1pjBsMQ7Ig3kJsxuwhbXgxYBJkKlW2732ZZ6K0Lo75VKaDe
HjgVhoYamWlZOBlSoghYmsP3tA/hiMswvWFvKyyY4QbZXZgaapxf62MhKq6/WP94
8VgL4oAqHUIcwzPFPm3N4xPY3UfrDMUZ1ILxLjXLhu+HPvY0UNlH6twJwL1Deyl3
DB3UuzWxeHqDRsEYxztHK5pPk0lDo6c3eT7q3Tmh1R3mbOIQkKZ7keCaYPAsIhFd
0PRVbzFnqtcumA2STnswuxyESA8c6PtSeXGIK6b5LkmhCcERDuGA0XYa/Qxcw1it
2NZAF6ROMOcXQcNVF+hg4gs0YCzaq9Ks7Zfg8Nca1I1qRLE8qW/rad6UCoDfOVlH
UOHFwlUXn9PNvvYM9IWtDrMnDPNxkyHhkMJ6dz51olk3UrPITu5rKpdB8HRfFTPi
r9PLzY9bVeMlB1TEIkGkeYec73qcME4fd08ST0bbsxNlmdjcEfNz+sZXQrn5isgM
33nlbyViRIRY1YBJp4efcnKj9gkL0RywH4KISHV9bhv6hHxtksRQujUgn+ezoven
+oDAJB7MJ38Prn6D84fOlbCztW1IwWmKQs9sAGs5XNrTUcFcrS7gvdSB2KediEue
YWfXHkerQn5uXNq3nsKLsR644AllPBHzKQHngxF7o24rqMpzSy+Ytb7cQ4Pr6yUc
k9lMmedjNnOxU9DH/6hicjqzU7DoVBRf8Ds/kv/v18y5NzcEBA2khAr8joXGtGAk
0FsyWSIkR7lCBqf21BhCf0lYqDct0+1dgzcCrNZrW63RGRxUVwCY9jYmwkhu/DEB
T0U43WZf/PV4KCTWM7Qh6wdwDVx/opbHaZ1BDfJX74t2/JAV5d+S+ibWISa+m76E
0YIJz+K0xa3Y+pC/j+/Re/mlNYBq2wQC0wkha1JqGxn7MJmVS2PFsRDwFxlohGBP
HLGh7P6hsE++mzoFZ/0wRam4Y9k8VACiLY5BHSPA8MIq61KgyJK3hrFVrTD4Qj+M
KYB2SAv/0PiQFs5OKoWDutcR17FkiFn5Wm1LV391mCnX9iLW/wl7Yi91OPWjyEB3
VKnCtHhDk32Io67EjY0uIx948ZY357iu6UT51BdOxxJWbtac/K5gus6j+eLRRJ+v
6T6ODWttg0F8RD+7rJeVLgrcNyDNxS6Qxa25/5V9cp2fPYoUI75djh/9Wd6h56xW
/kcMjRclpGoHf9XsD9ZICP6ZJX6hHek1NZWR56isMTmMtjzH3xw3GqwU/iEll45S
RIH+1igzfQQ5iiYL0IeqsBfJFS6nU8m+SDq9VQWSyp6wzCrmq/1E2oMLLHEohcFS
9ucLLqnaTR9r4bvThsZ045PqacrY/JecPKYvI/KQ1xi+D8VzDP4KXlsBkRLFF6na
EZY8WljG2dTVCJzdaEf2WYXNdizCSY4VRUl4R8A9mAdwmRWTUBdxnGDnl9mBClF7
x/K8JjUirfrpnvM+5p9n/CesXRqZ25uxsuicQcIxq0mD76RyL6ZmbvDr5XHga3h/
otZal3ywO5a0ccRYgd2BBK+BOk5WuxJeWX7dftrkbzVmgTtvJFaTxQiDOzfPaP98
yAnkFjtlE3IvJ6+wh3ovv6mD/WMoLDtsHT9DRX2BUpVx6z2RNswjWTFpVWpvYQHH
S16ZQT9OYB5LjiukTObFtPIu2Dwm9FHJPQ/svw0D1DG+o6/NhvBFxQhd9GovkaVc
JQr00Rcna3MpjRl6cyN3/II60Ny9KqedMpMZmEVIrkkSOEsuNUngihZow4l/gCLI
xqMtgodXTEx+TCsjN/yNRi0flKbTHlAXhWLrtFGzyUwgemblHytKzZ277VfsxMZ5
DYwsHBJGksaVbv+b5jldpHekTIgJkAijiAK/Q4ySIekYVmbq1+iBi/E1OkohzUOb
+p207gC17Lwcsv77w3pz3y5PR0yaVus0EMHGUy+Ye6KNLJ3vz/lrlrwFPy9eFFxW
T2aGWw1G8GbL7fvgusGw6ie7kNNvcdrH/QJpf4bQp2Lr8jC1OmoqEgP3kJFRMZKZ
LYXfbymwzd3DTOUewbi3aR0nSKMoDq2y7KQVAJy11aUZcC0zGWtlY41/y87hL9B9
bmEo5uQJdpgLruBThf4+9YIvPRBnLiAZv4V7Bd/6Kg43yUeIoxpPU6s/JcadsPmb
2TkUFo7rJtga9chqg/g8HuDsuvEfxqp4KLZCc+xGjEGqJwsM4B8yeD6ruwwvQTtf
7G0cKI1lef977Gk6JYkw5IBLFs+PQaNUFS8uFrzvvxmTGMi1cr3CEtHBt8FcXp87
UyaaEmLzNnhTRSfEd3iPTT4V6R/G46QemzfTdg13BGxX0dMWDwcZbwyGBas09GHo
Jkd0z8rpar+af8u6y4EhQcUuuj2p+xHDtpCoH92pWtUbeQvUf0Ho46g7Gq9P2U/1
ZoYhozId+v6LMC0ypo0K+oWTNet/jqeF6GciEk0+V7CH44OhMeUjWtUnm2egXy9Q
F3zW8LSKUKzQH3tJrb2aHjE+TxnL2jcXswPuQ9konw4oYIejA2yLq66XMRApf6Qm
rKIqsDt3YXd98RVg7jd+g9m76zhHNrHtCK3OAOo8BgopuirLpOsUlQuMR2c8Wez8
z+0LF6wQi7busx9BpLd6Ce9X4KPHvYOcavR5iqrl+Ra1esGJVpqx5ZAZ5ekbUyN0
gcLr7I3Qj/S7AOBzOtIgOvK+sfs8CB0X2CFm0Ed8epF6MDo71qVJh1EJhwlivs6+
/kxbzQZeraeP0v/8atJNYjbiY/6D3NzCpqS04zPEpd+qdwponPS82BsiDJWxR7+L
4p6PXu8JzBJLiUcuJwg6H7NMHCrZmN7/ddhBvDeDSS1Xs2j+QCo7XY/itynsE/VU
40Y3sMT7DxyRuhGhbmcDlExELjLZVDOgCYgyUGxoKcQYx5g7+Sgh5rpFJuRizoVT
P++eJzjAMQa1RbaJbU6loitrYKrmTzoztL4jrW6TP1lGmrgoJrlul8tOP9uQt0Fb
pUQrZnraEcdGn+Fa8D2tkGybuNrjNKkR+gxXIbruRYuLYx0B5rBzUkKNWtf5Fv7V
ck2oi38576i0sPkYw3mYF4IpXk9vSuVnH446gRhpUblfLGlTkS5Tq5KdbxHQKvYg
cAMjeWNQcWne3Au9SOYyD7Dn1VutiQtXlumjfMJkDwX/X2J02CCuZ2eKWoFqwR5n
GlGiPDoYcYSFKnrAWkidGNF7Xw6SX1uznbQXW1EUlbnZJ9xamjv7DQdg86ZqlVAj
jN7+sFFCPoyQVDA0AeFPAytFY/MMkjxaq4sHcBccMyCNPSCrPDZq22V+4araAnge
gRzN0K2rpIi7/TcRumsrgS9X+gnU2k2ruBjEqFUtAUrpHg8tZkX/BTQkJgo6I5Ze
JatFDg4Wm3l5bKmY0Z8qrdcmkK62O4OU8jUcJ9vxPwoH87SydEQ94P1Q1mDpaoOu
e9Fb8BIibhQWVPtAdaglL6qtcsfKUbje+G9R2n4afDy6UyLvXwmNzpPyratbl1sV
+jXVyaD2bmQVqFgKxLGmEXhR1zDMC2Xj36FsAm44+1eCajUI4MfmSwOnBQnAFLsi
5di+MFrUjlkgMJLt9mTR8TSg+dE7PGDK1OmcaQlNByWYfo2af36xlOUYx7z6Sa9s
VaQ96tA6gz+trfFRHUuwRJnSV64yULaCHT0Y4LA8KgUbxxMNjAus0n57sKGYwFVF
Z+bWPdiY3KzpaucHFxzZmgu9cSAexW6oFpQUn1b2VYPPZWW+ogp9L8KT0+cECP+W
VzbEVRrwVQrLVfzRPXtlfS0xpsbyfH/iVHc9S/XcY5JLGW/1vVn91GNLIPVciFn1
q9gW3+Dk2IoL8wnSChCSszj0A2ts/VHER5k6FgF1nRdCrllcwgKa95a+uIiHe7bj
QocvV/6KGplt85nMXOPkDQ6hFbyUW85zFgcqleks4vFbEEXM8u6umgpzrBm1CEx1
fZXLJQkuDm7/rtmC9mqUAaw6ui3tORK/P/g1unYgXe8TW/QPM69ogshiHDTXMzaA
Nf9EU937PMy1ORpCzyHHU7YA8VwcjUzk+BuV5ArcVTx6bQn739v7oD2VvdPH3kKY
ECtnukTBiqhe6HeMF0J/YQ4iypZkUP2gfvu6GShRs5cvWltD9lPTLClXmuhpuKvD
qWDfQxfzsJiW+G2gsjsRprEcfroD09DaLjkQ+vTxsiz9mFcARh2j5DszfNSdKmsc
sGxOzpJ+fp7F+oBhtjWK8RnEmePZoFOr7akv0WUz4VhFgIvy5yzRXbqW3ydEYwjv
6H8b4drCkuS4wdYbTYIRpNi3tAq4DtkDsPfMxOqDbF+4lTyL+od3TeoixobpSDzV
4Xk7wP34Zd0oAT99qRYtzHuASbHDov4qOoz7LonF0ek1i6WV/fthq9CrfdD66glq
pfu+PA1m0ju0Hs3DveZOE3zAbR7aaAzFqm8B/8tcuZ5jg187Wr+slhPCDjKrNFKl
XE5l47QrNR0Xe6VNAHFOXS/tVw8tIdTqEwVVPDUunQ1OEiQHwlLar/Y0wiHdMxX8
odoUMxQl/chfPm6bHFu8HZJRW0pdbooZCHZOHRx0ft/8qQQm85ZzlLnR2/aMz3Tt
ndnHfajhp5/yCXKzRUn162a85dDxN50FxszFoYdubsWy+uMMnpEMI/ru4QJf/uEp
75oRy4fzdQSl29Fi3YjV4U2fkbzrM5iS9K65ZFfDbt61iirRzeyOk+bFlypzkl0O
1BvolGYM90LcokDALYBGcqArFsMJNt52pU9Ww9jDoX5ouixrbBlsl9Svs9Yqc3k8
4BwdtEiTtGETMxg/3AmzwXWPH246gLXtF13Mj/1zUkbWgSKcEjHLHb9VY6Ao+HvX
cpWK7AfX/50YUfBZzm0JiKvrGYblPP6U8V7j0lKRxkrGhApZZiH51YgaQsf9ln3t
wP65q2W/1ZQhYxhkfBcddPYwAJKBTDzvL1fyaY25Fs4UBZ1k92RxAF6KCVmpig/L
QNRwIhQBfJb8QZIhB09hc1/sbu9x8WYTY1yo6R5ra83ZIc7MxwuLuVJbuZithqnQ
WAvJjSpYAOVlEH/vkysuDx8Wa4TjroPwvR0U5vWYC1iCk2vNtdsDx+2lVwy/Unry
p9V5jv2yx4N+Ji991wdadEV2k7PcWXEXniqQ+lyDLDYxTMLbBFUWf++IERKOQIiY
2BvTx8010tydPo9GnbG6I2EQYDRtWD5wr0dJyxdu1mAXjFEB3l5LgskVZ2MDmnsb
ExERB6m50Me5MPSPWxvbF51Allrzacp3rKS0R8008b4EvQbJEHTS2g3gtC04GFl7
13oPLKMSPlq+DAripb1Z2UERTV4vt/hUOj+SDdp69c+eS+JkNY9bs1GrR2hBwS/Q
VauxxiIDWmRt6u6JYjIVRlPZBhFu+4pvHZcp5mRrvfmX62eqdz82BNlbpaBWRyod
CK01Nd5uwNOSmi5pkE47gpnTZCcQm9M86zyRmnKsRn5QFH5UQZCxR+hGU87fPiEc
k3R65E8/FkQVoiS9qdu9Z23bVixf2A1q6HQXv60elDkCBTHDim3l1vzql8Z+r7+p
WTwFF4ZIMQ3PXQ869vO+czG/0g9AJ6e06thRkax2FkIIEEs6Gr1areW+zCpmiWju
Yc6N1PXMDM2Qqi7F55fZZ3GU3r/wKgJP9NFZbwWfk7AwNi3L/SKvHo7EonhgHkv2
NBtRab1dnE3miwfGN2uMmWYCindSvtxI/YPQE9w/LpVbiX/tQavVZ1SZLz1qee6J
Pl1O5Z16cg/Nloo+9e3eFOQlIbA5wbxxDOM42xkXAAm4iGrkQK+4LBBOnYpz4Ss+
2ZBl7Qg7rS8sdac3Mfxbn1lt/ABfrz4hYmoCm9IQDQbbqlEWRFCJbXUiWUIV4M8x
ui8r/Mot2c3qptdn9n93Hz77Y/sPj73iKYQyjCq5qbX5VgK8QqEe50EgyA+QxXv3
3MIT7YACCPAJjktoNyzoxmWqZjCOxI+pKxmJ+0Vzo/PqAdKxMY1GQF9g6UIbqnXx
Gjwsikn+QYnxMoAOexKAVEmiHpWPrrulIFg/JK+h+QJ8d4X8/M+VNoipMgJ91E2B
fkN+kpUFIJay8Q4weT8qZxdIPZg2aYk/G7lhJenQ1JQ2ZltGY+K6x73tsRq2V4oJ
OFsiLDkQQNeUp4FD8ov7ydvcz8U2tB9yk8NUggpA+r18dHRmju6JvxqYsLCQG6aW
h+r3pkTXZ/bBcCJHzdhX74D/Iqgl4pHsC403RHI2vAr9VKNnYZ9Wfwi8m0sj5j4V
xlkFiM9u48hKqpALdMmZS9vlHWEigj4dbPE5NagkSBPwi0Jhb/ydqqtAouuPpYBx
U65xkGqJMOQRFBTDSUE2wpBbmQa82clDKLMP1POsSQ+wyXzd2fzDKH/dysjZSVdr
h9vKrYmfCHs792+ZrLDZZuawfwdG6B/hTVbf7+xC/nVAeJT5VNu4HxD+Xu+X4GZu
qBAjx6a8CGMUJA6hd9N+pcyDUsIPgnKkN+7gam5NOg6fKfYp//yXD9kMovPFuIEi
klcHrp38HqQwVpEeqJb/97nx61NlkRpVCE8KYsYo1reOK72rnL33sszNq1JfpJss
6zbLlL5m0CaoWv4GM2FkWxvvuZ7ggZQg3zDSfreA5hKzTYH20eJDQPBw4zNydckn
dZPN0wq1f1eJifTPhBRfnI9X3bLaYNa1eATj8dJsvu/8bO0rlNkJjWvqWcXPkN4g
OZdeWsyFsq3lox8BDnve+i2F3OlbNQ7nzCR+KGsEyhT0/AZd3XYITbbKlFZhQRbv
aPStZjKpul5ebejVF2dMguX0aUaoJGthE2puJhqrZ7dtBTWEDp6TcudatBdKGjEJ
AZoPwO4K+cDGQIW6/Kc0jhdzExQBkhAz51MxJ9nL0r51VEH5cnmmq7xBzH5TPQAr
NeIg0DZIyZgZaQUUxNhHVofC0ptvIIDBEsK9g+iUMXknT0BCgXCEKlr41Phl6psz
95jdnd1WnBqfoZHD5aafEm76pZ3BgJAt9WC3+hgiVuAJs9XAkxJynfeOiILzNZ4n
GjpV19DznAdXDK0hrpt5wB/zDTd3gJ6xwNmaMuyCaqT0EyNIyOH0dzJ/b/Q6spwX
atfJvMDME2l0ia5cZMIdtwyQLk0NfpmuqmxdQSELI1ZI/77VEz1lRCvlQgwxM6KS
P8csqiJUtzdq8tZH9jVqEfeABtA93lBQNv+o8O41rT1chBbPiU2ycPtcs53dAEcD
ezerS7prVbKaqYfA4exk+iVhr7KTfmbFOULT8aIQcQne+QD0sO47q9+CK2Ut2LtJ
+viJqGzAmxdFcfSKdsu/FILZ1i8USlX99D9ejP1l3vMZ3Elvs8s45Pqodg0p1/Z/
qUBVpdwppEfijSySA94Yq7DTA5zSx+emsk/Fv5o/4GfkZpqtDfIVR87YFBwvaBgY
y53TJkx/daUFSeoU/1jzJxRnDEyUiDcAAIeMvHMop6+Too0n44nyy56MYwgxN5wF
UAJH52mBbglbB1x22EqFgfYX9r/EYMjQKDAJd1Gxd+32oEi1qz56WxjFS636yVAt
qdLy6mDVbuNfIX/XhDK8kf9FxGz7odmQk2nddX8/TqOGn0VgnhPVpqqaK/a/twYc
tcoaDGG2FCZXEnPaC/hMaWWM8wkREzegZsi530KqyCnb2Y8qwm6GN6ndq03T+tF4
oEJrAiz/MbI6f/SbOfoeWKDu7LbWnxHHudPbQu1RZnJABHA85VxjrTPTY07yor+E
fYhvmsrMRHMXUrVASHEKby9a9d1AMeK1d7fLhsKohDowLFPd49ZUs3flS6zxUwwk
87aXoyereIOCK/BxVYqJ4QT7e+dCpadjQvb3xKvIzjYmzMV3MV4hSgdSN8V00VjN
UVsRZIl2rBnaGLsbzkSur3YxOIH4MzHr2JmdTzDaQJOxOHa4zbDf0ZgPoD1htps4
tZHz+FYojPTnLgwXXc266HaMPKXC51WjQdJP0nzqGhXXOJ/y1k/zWyv6TjFzQRHO
8eGahwU1VxDLFbaT7d20KQAaVpa5E19qlMw8yzbVbvEdwXW6jYAV+Abb/aq7oc8q
b1Uc2VNg9+70LN+Fzb4MaAI/YlHWL/rYNMtnvMjvYJzXSnE04xtN/1iTrmaNQnI7
/ZPBY4+Jz8E/dtAkBg0jjV5KPAZjpLthKKXdDbV9tGJa+WyWrfPB026H8Xgwm0ff
LGr1ug/Dj//q3PeKyJG5ich+ymgnS/+mEkYj5wKLSaA2KBLbfU7T3VpLz4NzcvU6
OtcrTlKV8X+wd5Ou/aA/bvmyICN6y0zLutkx/XaRylR4Ms6GkWmOceLk5nSYt29G
zXfWzfo67YSU8tJIZSvlNHXLhQwAvSN9ypICGtXPM5NEMKFBMhsnDkTIzOMJF4Wm
Y8VeqB2VddX88JogSWA9k97xzvo5qvku6qMET9VviD+CVU+jcs2QsncNyBV1YnVg
x91zOim9pbO4k1KGvz6x6LnQfEPEGxzpvS8cqjV05b8e6BH5z9ASaGmFEsmE9iRd
K0Ev6F13keGFNCnMecNnvGUPVsaq88WDOJZBoWm55kWn1OI54uqKdB4ldqxMGt0O
YZH3D5LbRU4uGhxDeV7saMMY88bRB6NN6wUx+yaOBkU4RJMvkOLy6HLeY1zVEbme
kadPNLuUJPGIsopaGLcPlPHhfuObXa4zoAqfWqxVZknPfoBOGZypMxxDxviWptWo
GsmCOxwxwFQ6o6jJ1T+IUMlBQpCzM5YES9WbqP+ajzej7MA6JbL2zFZWiCHDB0qt
q9XQi0ks6eOU+moNjjBrELl+SuaaZHtW56rJsBOHEkT4Qw1575bmbkcau6jXc2XT
UYp5uYuDWexbG692r9M9R0/A3drNn/+8W0nDgX3zvaA1GbRjajerm1CtlEsgA96+
e6+OwmEaYuzbzTCOEAvKKWluU8JlXtjUsbHmZctYFAS/sJzYZDgZ0HbqjXdin8Tc
dhvTK0mxRT4cdLp1PkPw7lUfKsb5JYJ0RqyvW9kAGiL5uC/uIPbmz5fHPfulPE3a
p8MnnfaWOawLpeWYSBNIhPpSVM80uPlAvDuDYEqStAtajHf/yNM4ety4Ykb4aTtZ
Zxw+VgIsLA1/F9d+bZwIP7S+dIS1V6ja4/bh99OUpyE1avCetZq1rVyeEbhyJvky
nKN57LQKIcKD/JEc7i35oPIEgUWdBDs7sE2J5/PtPEYNpZ4gQJOs6BlHjJcUUSXv
xXYZ5Bgy1SO4WRjP2KmNUiNCHDI992K+xO9h2ZDfEl7mzX9uRwke9UjuCtfNrZDS
RYebDM4Q8k9mfnhufV6yq8jFdkwciFswge9pSrsopbzK0VE8oSlxzVxc9nQEqVJQ
F+1CQDfzHwomDyZYw4qHb7WAdp+2QtEyrGw0rIW51NyBuxBImwUwIlI5AQmSG0ni
Fxhe42+CuL1XjS2H90XjuWPk0dz80pp9zZ5sOdOUxL4bXAcOa00eEqLBuMA4Cqmm
OpgTTtGrjj3keUf3tPVsqommzalHzRzXv/UI2IM2SrU5XI4U7+2TU21HTaXJMTyd
BU8kSkwqnuGWstxQ1yen3bOhEsBUtLLgH6SSiWUbuXMTLxM1K7J2sXc6hX8Mg1Es
xCrwflvSoZcDer1tkmcA9K04rV/OHn0zkKN4lPf9X3y7pO5VUN9G8k1Npgd8X2yD
U6krESEOMqO4an6RoFfQsGPooNzdzkLM3c4R8BikknnSLoK6uzE70S1gycoWdgWB
FIBSwLLzRkXEFNFwbHREcFcGOtGmnagwVUa4wZjyD8kEO9aA7B1o3QWDcvojCQI9
95XLrPjvqlFo+7Sa6xp0AjM5bSVjsS/XYN7vcnFUCV4QtwU8YGjqQhQ+Uq8lj8tH
OHoH8tSBt2fVEOPIvJL3U51RNNzwfAxanV7YgZOcqoqhSti/fy55pul+Aa73FLYh
vQfYDEWCH3nnGtw2aPNU0/72hkpDJ8Wcy4CyUYMDFSD+VI4LLufdcJImdE/Vzmy1
yhCqwCmS8qqVQJvyH+w03GXBu/+Lf6LiG/iGC3IsHLrdPnwonrPa+/nZBRVCaSoi
AOSEdsVJj8jZ0VzR8jfOrpP4XlfbyOJjSOl6mzepqc41gKfSXGUC6Tg5KekF57u0
JB77YXwtoiNyboWGGtnUJSMS6FAlBEL7bs0MRQTmyYPHJrSKakM5Mr+RGoLf6lH+
nkeU2rN+si3/kNB9zyMlCfzwTR4V0+JH7rR2ycp09xC/dpjBdcQaNYHOssVZGqed
0lE+8S28e2dG8zbr5OtaYfhJjXc/tpvQO1algntFta7LPsJT+1Bjp6oUBlZ72BMu
HINpmMvQPrXD3r88EFz5/xsXBXL7KExeMOnF81hHtJTNxUev6DtBv1VQFME0obfr
ZHlfSs0DUFL/AXBB46S7B8FAlKltBoGsRcLXMsdv4DqdmdNH+BSJP8QKklExkaRC
EZQqvON3Apocc5NPhruqyFMrrwfXgixq0/MGCu2x6CkA00bxfeRUf6hNkjvQr+pj
fkIlMWzcMpUrAUajYPqxWIGVuKbq8aqO1HrOu1GzvelYikoezkfayk1GqcRpaGs9
aStm2gopSEv/A6uOBqbDC1Gtp0DDQHChjB0nRxJtGHcGG5mqyCzXboKCGZrT8RTw
CToGODHePm3YdKsVOGVCPvJJAa8Na3/DphQ0ei573RGC+G/ZV2MOGG5hmllCySJy
q9bApyyMsm5DiZzvs/nBa/mpuooNUb35P0oI6xW0gGcol+xIh5fiJ6aFoUiaBkiB
E5LpZZ1aMBvd36RfmMxntkD5ThrcqzEdTKo73ZvLtWkHt5B1pRHPN1ClnarT807j
4HfW6v2slgFUjYk/dgRaAXfMRnR4xg2wx9xwhdnFUPHSAO1LNuSPpoWwa12+j53J
mqnNDvlYx0/vO5OIxyLuJnvewjWq8m14tR0khIlULMG7V6Z8EvmYKKMLZAnZFnG+
/VFsRubLwlLKT7hMhmAoatEJiH53UVYSsicJ8WZCZz5cX1sqFCyDvGf0A6BH7pa7
M7USByCWIof09HGXzYA6QqjKqruJy4TMQz+6mJBrHB9CC6GrocjWS+2K4CXmYuyd
VrRFqQfFClgKTfEc+RkVPVM6Yies0nDr/KKJPah110sJ2m3xCOz1FwjLcB+6zULs
8T564NqeJ9WeeKuGK+odiscvykwNS/ARek9D5DA+Ty9H1yLmLggY+7AadVOcTm6P
Q3M94YpLD2jvRUu2EKyR5oFueC9krJPt+pszh3nnRAtZ0LVRdDJRC1aQ6rXJNxky
5J9Fy/rl/J8R2tguM4MEfGznEWij5yusjqX+nJ/xUvVWNAe3O3eIQgDv9qkCaZ2K
QAaGYffPCfiwqRtdnZd+f93vq1stvtKKj9+3rY3JRybwhNrSYatfMgnc468uzWyC
FxMJ9bwY4OqDs82wWYTrlmSCCoel0T1xT/MFji5yBAc1vCjL8T6DBmAbN+W5lLAa
7/V7Ilar9idZ0noh7nh6VDT5PguD+wEr0IO3F9FZxUzYB6CiMc2cBnEKe3VeiayC
RJlSJ6gvTsE1GmCGeHaCRbfp7ujpc2wtCb6/72TrhpFnq4dOCV9+Hs+5ew/tzo6P
QgyQIERnEBbWC60zJEYFZCjx46CBtx9zB7z9X2It98Vq3zbdMgqaka+lpb73Dopd
5S6rLL7h0ngeNB42isO1hk6VXj+Bp4yY0+kZypjvjrqshxL4PFEIrEnCGsFuKp4W
f/uEB1Z6t/DxKMzwBuW7hES/oiBhZlySiaQu9NSAMO++QmPyOG4ra2794ddWfVu3
cAC8Mt4atQzu9LkMwUd9X0ZX6TbPZiyXIDCJrw8jaQCx8B5YHRZTtAc+Go+R6YIk
xE72NcyWSfXvtlp7aIAr2pysI3fP8/laQTbq5WB0F6SIckBItuQE+MUev5gIbQX5
hqPkxv4fhwOOZMe5OMLN22d1eS46joixNI6lWjXJ5/AWBCNmAW3HSbxyIZ8kbKj9
7wcckOlQH8NZB5/FKZ2JPUJLAeTEEDaEZWF3bnkkeI4Db0SjF6towntWizlVEfQP
hzuq8OXhoT9NGtInRZ1HimKcPxjhCa0fmC3pou1WtbpVuGfRD3tZ9ar/8oJSTHU/
iNS2BWsYmAwjpVtK+KZZgYwIk4GWj81FIEjx8ZOqSnw95FvGG3wya9vY0eZ1wXio
D+WRj1/y75SdAznFXFFPWCnWDrRNDFw61Vbb8MIx0xOhSpwaz/MWX8mAHFW6s8BX
U8ItJz0YjRngZkJbWI4RyRfPPzg4DGV9Kc+ak7wnpJ7xecs2+Jq58FyaMCoRHE9B
bJLMtfcHsZWy6/S6e+QriAi3Dvp+EEZNH6ZONUASOiQgE1n5jX3almtxI1IunO9I
e9jsmYetYzPd2refH1wDi6ZBavpl7+ayoSJ58IxMv/IJM8d7gow1Es3fjJt78qwy
IufFVIH7fAjGPdswimnAlCWd8BxUcydnRhosi728q7A3wqov7lQTOa8YvpReJF6Z
qgHiId81dWSc5U0t5fFGJLJfPa4S/bctqu/RZrQ+40Ftcyc5z58GelYo+dVBhQMo
W7L57tJAM7Ji71e+IonAoadquX+rBJjF9ZBrfS8H6AXbh7HEmRTMtTszay+izzPM
PnEqgoyE3o8Gm2wCG3q5ithTO4sS1s5M9wFbavHRU2fQUJp/2ck9tRSu1IcSupVY
icz48nh4dlR5yrejF+cRxwmTgZczpvIVicKmbt0PYSktqMna2gJXBwvj61J57igG
i9Blo2lRhtrpn3gRuUgDnYGRaQE1fcPz20jlP1loo2y/ZHgD58ioFb62spA+8h7J
WG2341/i97c7PT1VWEaxuDmLZP3+UPIouoTxXOGQY1UG6N7QJFDvHrjy8FnCFM/9
HGe05gG1hVwIwd0hYhP32m6UecCfGS850bcLkBGli7M4rTv3dNDGa4phIvPkTKLI
XTds5R3Gpqus6CRYUGP7WANAh9Q0hi3ZhqmABz1AEW7PG20cZW+vFDGXabXfLU5y
pZmbchQya3Iiaf2pwKOs122h55T1vD56D2THRih+/AjRaPeihNmG/11gqpW3Zpk+
ddjBnsN2ULJnrIWKdmGi3qbHiiCvrnjRGD5AJK3ZXIxInBfefm6iMC8XCOFP9lPQ
8NmAje5fRKyXaWrH4by5LJ7C5IK9r2dMdiH5K4rHCRVRfcIqZr/Uf41w47qEDHWW
LU0/3DHdSIsL9ZPxE9g1lDFjMQSQu/y6bAKbMlpH45Hmng/3GwGCQGKAWoTcBk6I
qdo18ANutVtJjHvwhjKOyjmje9mH+94tJk4tPMMRCNCQ4ajcrWt+5kabcuGIDjf0
0HxzeDIjcEa46GfDwuxsqp6UvfxE0EzO4EpeP3Cj+9BGqQtu+SScHJOx723J5CAn
lSmEEekoTu1x1DhQB4rfqNuWIm6sZNPN2IE3EXsDhfDf4X3GLmnTUa52hRq6k1vS
kUhm/NT98mqcG+ng0cpIsnu+VHwk45NWLmISJdJJv/AsG3+5T2RTebCS4sVTdFnS
4LJ3M1N9tiU7PgX+fTggDpb8FY7NRUdA3JrVZsrJFgg6zbgyr8x8+tdS5qngLLD7
FZ3yfqbnvKrjFiBAzRoHNCx+p+hmHrcYozSJHNOYGr2jvxtsD05bzpuB6ga/6GtZ
Figq5dZoPb2SfracAYQelQ8vSuXWFOnNo/h5HMx6NUzYhlht1JmFeQ2PE/EB6qiu
Pba5Q0GARUA1RNwtpnHuNhasSh6miUkPwE3bMS2qLZkiOStHqbamw7sRbuDh9I1l
N3Y7Mg0WCoePGZnL5ByxTDgwApvGz4L9lsBODJlV0RW44d1FYLH0M+GEFNWf7SwS
8gAHMdWFkZvhCrXQpVBw9rdG2NCYcQkNuz1aoL3ybNOdrRQk6p3xdZABJMcTBfGR
yud72XqocNanevXejq31s+isp5bYk3Xt062zRFol6c9OVovM2PKmPrHB2Uruv2CO
oyBCxj13b4MGJrv2cCsUq0iPAgg5X0Z5MAvsG4altsnwB6Grc+GF0BIHknGn/7/v
l5Nn+y1EbC+DbdDLCwtsA6TqK3zwheInuyaBcYvn8wsOHj79+btxkMI+zIQDYm1A
BWZF3lD4SvJO5dLUCYt9SiE6gnN5ncInvES3WjscDq7Fi4sSRCZVNange/8U3N6+
L/9vPQEEwUzDU+r7z7gcilscYeBHgR4+3iqJ3IJoLXNuIEAMH21AyExgb4oB7nJU
y6kgJTgkfoFoKBMt6Wral3k5RRYQm4ql5OD+lAPO8OfSAH9KUXYO7AV/WOsopxFV
RNK9FfU75q2bJSHumA5OmDBX06ygtxBJHVBXcph0A9GULPLkTXDKQqQRd67OryHM
aR+Xsey8Tt2mItToxy7sh5LNHbxByrTV8Xpay2t5CYCZsm/PWbpxXNjQ8wEn48eM
QhQ+zYKQXRQw37c4HHlyy2iGFg86nhdt4kI1IcUXbAqOSyr7h9t4XCL7alPFL1aD
DjojM7JdRTpErs1dV/ms/C5W7+9Zs/2a7iN9I1gDCDNHI0vH1zeSIRsi9E6AHn5b
a25piXdan/sJp3gUe6iEsuyYxIowntKGqcIPDDHuLhhkfMie29FdYyaB1+jNGB25
LSuHBs0A9Yf99oc5dGmA2uUdy+W05UwJmlr5ula2VVy0IFILWpRkBs2tWKPupO4Q
x9Dp+awnGKxgcrttkTXEieYqw1wN1uzH2vMgEXDqeK9gQ3FlLzGfR43jW065kHDC
LaX/kwQnujhLA874xSt3xLCTlEuBbkZOIXArnKI4zg0xBoqcWTKwlYNwKK/3I0wN
ipyIT3eQvVnN/zlIi6nwc0nR7t6NvP07wiFjtN4qrpsvwwomoXmp04W2+Jq7OZJq
KZbvoIw9mEiTAidOoJKmFuLaW1iFFKsdcX4x+jkFA5HO9DsvX5ptJMFXOq4QceFp
lt4l/hp5sjUsSR1z28foww8FDnsk2NRHhvuvGazX+EFMvPlGd8QR323TXiF2MMne
UXY5bOhPmk5ESPzDUchTRN5BcwncoYX8aS1JGTcSonb6OciVS51vsF8YHG2TdY02
hTui3stf2HFLrWuGmcujfWrxZFIxA7GXRjXK7VsT5zPzYODyPOFltYIU1J7sKu3B
1UNCTchSI5+5UpfKmxaOhr2p9XKB8ayJ3z9DaFWG0WhF+OiOnJJDH0c4NCAp0H1i
G8BgrhALjkzQdcrq/Stqh3Vgk69TTuWlLeJJ8PH7b5eGrBmhyKBEb40UnJFJ+1x/
b+blV07i9BqRsQ/wkBMtYKDctGOqYLLOJOFdB1b933iI9u4188mwR2mEXZqP6zn6
kk4Tq5LkZuJw1Brt4Ogw+SRIHyOBCM1UgTpAfYDmAsO+yMPtt0tvAcfFG5KHlzGw
gGnBwRHCKAsTpKLU8ZA/fPpU9yOkeH69EYvDi9n/ZyGmkE50+sVVFz2jpWAVkLs/
flCJBmVwOF44h5pNUumx6ruhL2NuEPkpr7sws+an1fO3zBbUhauWcceAaNX3xLLF
QMeL20AUGilVztUM+zhU9xFqX1cdx4YBNivOBfs4DSl7j768Zuh+sKI8LiRcXGdh
GUVwg4/DeEQ8jSr5SmL54caBuYgdB05jgchInjHdkKwYKOurBxJ5N1EuPYRC0LEB
aO4g8VqQM2Yssrm7CLEy0epR48braElNt5YIcA+PdqZJd3lzZ1WHPgvNAwHNEJwo
YbFMnjFdi/XW+wprRok5/uivuRLyRRcPNmf2z1yGAamkYUtpoUoEG24VwAm3B3n/
Ishhk7IG4PxNLuURCyk+IJrrOu1rRBX7HeCsMSobHSGPZyfhRtj2C9lebg0S2ezb
ghZ4KtLxsnGocHJepdzQ0xuylUkIuz8euyNWXUFPpEz6Soc3KmVJosCSea0yx49w
2UOpgU1S7JTGXnv9/TxrNdMLmLSCXke5c2x8C8a0epCcvnHCZBYRuZZEGw/ZGCXS
GdXASVacEtQznIN9xXLzU9f+fQ9UHT95STHbhPiKIx8jg56OCc/g/bkiNSATHjWT
L/DJUV8b258lqSlYu3GC/rVyXVHEMYWPKkA8Ptgpp+LU7TRzjS3SGYplrtusTLfW
DFzP2X1B0w2omzNG0MIOQZsrvYCYeqeh62VzXypSU1R3ZBoVsLD6ELwGRnGL7nAE
vGVriacS4bOO2FPHzEpFw5mFh4UQRLs9HBPtacBr3C6A46M2+Upt3fYuWRTObkQv
g1eVQliI1kihFX3+eNe10CbEV/bvYgtYq6RCBs8A0U0Cb/jsFZIEsULOy/ifOebC
/51RH8nIcyWymPYzaodylIFG+uYXoYzWdO8R7nYk1WL8/zGHDVSxHRPsK2bfwLdQ
xO25HuS7JkPK8cikntHYLIBoERgbrrvnyxSjwZJU0mNvDQIpykOr+ZYf3/UOV/VV
TpTtPp2MrlaBMZSpQJ5EUtocK44j+MkpvrOHaea0f+Jc3WciCaHAoVGiQrCh7sxE
xNiH4nu5LAQuxdhiR7BavwwSaF4LYOFwyy8kbo+rJs1UN+J99J2TZkLLxJ71qWvg
IO6NUONEI3HJlIKaYD5yqQedUN4byheE0upFqT/efVvKuwfnZl9ByGhTAKmS8aQp
8rH1kUEiu3LXsYVd02oncJNPJM7Emh952BwjZT9QRskuRu3RRomSVEu6r5XV7jIi
mwnFyBN0fM8wi91pd+qqBHIHcuNhUVkVBQp5eLXL88GluPaFEdyczcvKedeL5KYl
thXW1OfGpdChOtOp3JYG5sBKifHkDysytTWNNNusdTxkv5Ao3IzIGjkeb46Hb86l
KhGf1ypBAkIlzxD4k76ujTD2S55ZXq4Rp+VN7myxQlDNVR3iy+puZvtBpGmVYeEl
/xw5CzZpRYz+9DbX1GqA5Utkg5QmuseZfcinBxY9ZiVQfq+CAXMsjgHt61Yit+Ow
BBnltBs0lFAKTtTfvsjgsPteGgZSJWhTVrgajMQnTe64xKMZoZFgL1DdnhxXodFP
GwmLLYA+GUh/517znDWwnfHa33+BvDTWXmosE+Qgl83UmfAwxN2uF1CVjSIewsAI
z2FBApEja7ja3qcUsQwIj8otwUYhtzbXh4kFvfKKeKoF0lhkD25IgW4BTsVN7Jzs
+LqOcn20iFRPZjclOFDxZsa4G6xNN72de92m/lnJxVidmy/5Yzad7zvoxszdfQNY
JlqoscN39UWADXgn87HZswkWcrZAt685CalWQLr0TjB3DDuiNPt3I2SPdwagzB0r
kKMqQu3yd/f49HBsynHBBAJBk7bwXVhrXiezoiz3Ie/95MMZtSDQtdpI7+lG81py
GMbUfeK8NYCSRo8rsKMvsKCMP57dE764KTBQKbVmwBcxH03+uDHy0w9fS0ZXsuQG
BNqoblIzyt09/4ry6Z4lsg8QhpK2zBAkZQjtX3f8OSCDM+rtfN1ZqhsPKKKvu8Lp
BkCiQwVZDH8e8dP4meKqXbTNUfH+c2LtHD8YGZU+ft1odLCuWjUoOnZ+tcHZ56oV
KP3dW0/1gcIlg7bFru3e0Ou+1KnEd9L2vZoSKbCC1+CfYdJ54DywGq3q1oxhtqPf
wHSV8nmGKeGtzfyAXLui1OSWgD/mthE6xWne7OibIE9O/ITK4+TFV0kAMsD9YeYw
YM5rN09XXnbF6f5MOsYMzzxGMLnx3TSrkVebih+YG2L7tCNeLjylKp5clR8nnb+l
jezXda1Bl8ARY9m1OzjGJSV7Sjp0vJaIOjSRUyiRgR5p30jBxgQvnwDmM7HaPf2/
P115sVZObmtTRdYuL13dt0/5hPkbJdZOOsS5hS14F9n0Nd893moQxjQq9qbriLBT
u+MqRvclIn/H6ydMmLIsMiIPyB36U92IYVyumTAEQqdmfQ2KKGvHppmT9qFwbGHV
gIoFNJ7VuD9isB8bD9kcTlGr0yw4liLEr5G99ZF8ZmE7tcubceKprz2zzVrVNGLv
SibGV+ISTKmwcp466qPS4dN0KZpC0BwrEQmpiElJP8IKzRgPGPzlKGJNjCXAdXIP
VBVRjoPhT8Yy8Odz95Cw7b/MkO7DHZPgfAEvhC3i8lSWF1xbqp+RVtT9ODH5BeS0
3WvXtlwWn+diodENazmFN1TWQO6/YpvyHGw/TjOQvua9TblZa6LqoBTjFtUxhCc+
8x8nit1PFDF3oYvH5zAYNQwTQWswDItTJfAyr3DniNyeNaYdHRitPoMcdOqotfpV
ek8/v6ZkiicxDLpQfah/QeHQ1+HsZ30TxHDCk5NuZFQuBOAjFTBfKZYGJ5ZvqRPW
BtCldPBS0iL2fKoCbAiHyHeUwPiHUTxj770A27xMB1oCaIxbTxOkJcq7xm1J++zf
YZ+B1r1UO463/u4Xii7qXWLUJv0NKnPkiNn2nk6HDw24AnV0M6zu7JZzJKzMaxX0
OmlF/namv32t+r+PRk5ePf9TW84UMAtkZWJSaNVLQYCiUHASgeACP5Ks+vY4Rv86
4VB9DQPTRM2AfIyzdoOV8HH35mutL14rLiy3RXbZEWbVwfdt+3Ac6gwS+64E4p71
LHYAZXzloixcoU1KOlvUzE+M89xc+WQFIv4a8Z7Nw5Pw9BIdIkMTdrO7oU0zXkqc
RhrJ5hZmYNHCRyG2lvl7HChoVaqP5PFvKe5Z4UdbRv/oiBMXnOTTYgtXm1ag6+SO
W9Fb8nNRX8i+qP0uaUyTD8km9O2To+JQGwrRGQjQI2muaIM5E80X3yhAzehCbdUi
78i7cjSHG19kmvXJOR/paEI5f/pIwfhlIt27ueO7AdZhiHdOgld95UwYnL1rAqPX
43vytF+FhtK0osigKDnrpf/K9GwfneLIPvgIpUxvpWMbxi8liFM/zMwl65XYXuec
61w576vSA9H6VgyinlN3gd4yxpJgsPMN+hMWr2KQwq2MyUPecPqKtxL9Fr+5+oS3
8lzAQtn49IDxCPpjipiyY0OYCXwdV4OL8gHMFldN/bJyqTA0V1iVNmYu+x868y/2
+fXSM+N61lQoXsVgF7i5xpENjytbpWiUlQJDMRq97i3KNAoF7A987adYvwEqghEG
ZSkMtwPbIVklWdbRAuXj/x+Fop5SECRx08QAhxZcpnKDSEOzWbFuMf3Xy0JP0tUt
hmnDtn9MSeuz+YkFKykEdPvVKbD8s3E1jdQ4x4R8p4g8fqyZsb/1usCQQHTz7GYY
soigQFDbbw4qVPciOErYBxHMekQwMbd/UXG+pQKt4wLnkdNk6DxwTnhDvstSLwAF
5TKJ815lAVLl5bkkvLbSm/VI++QUkZPkib27OyAcAfpRVk1IDG/deTu3BMCWhmcV
Pu8pff9VvN4YONVzZcOSdwEPEK0Pjnzs5rJl1ST8s4NF5FJmcCgl1nKILlRoNlV/
jXpVcOPjYFH2QPii/D+WvdV/vcQv/IZUnhETPZchZuI3evj9MFKP2r1dDY3WwGWl
7wd7g+5lvS4WXv6QxGKsjATEPMFtQlSSmDbUbFLa+Yhr5sUigStzuUKgAukyzq+B
9Ydgje3rZO5Z8OFMRQafp6lAf9kfSTo7/srLhchAkgH9Iq63dcOnziiimv/jKZMl
auX9BnbFUUk5zgNTkStQythBTOyyZfNurLLzEHcFXb8CYSVYaxOGt4G2vJBzJInt
ils7fkt3BOaLQUxNrMrj125kSJS71mzDOoVMpGxXoLFZWgCI4f2s8kd+2MBczFVP
uAKkde6AhgREycabq9/aLbiInmH8NHnDp+MJcxc6fZ1DkTLvLN0n4KTa0nsJMlDx
aIVEkzr2M++ZrtcvOB4eHkPHJ9/2+m/lrAXpySzhLu3857tBD4wgcASyEgRoruJq
iQeqEU3J9r5w/Ha0pjLF/xTTmwWH3mhQfM6AquzFfomA3MnSQBzZI9NIamoOWsVJ
hqR5jQw13yKVF0HuwfjyHNCnXyO15ofRf0rCqOtDTyAGFAmY/2vOplNY+D9zsynm
bYztqkChP7KgaJqHp1AjlXaqfwPFw1j87tmmI/96zRDRHhi6XXedFEOSAiI/yIv1
8v/2Rf88BvNaBXZmMUB4zPpZbpwqDQc64+6sb7vXmccacpBNmyqm+R7vSwgCqh9Q
fWny/c5IAFFd4/56P1j9/XwYqPsxbY3r+hDuI2oPLaoE8+7mZhyn9oUeq5cxmQdj
7/7SBgiUhNSTMvW5D57ZPtJDgSkpIpFkxOab13rA/C65W3t31R1QhQJ1xsDQku6w
xenkxeM//5wzRM6+8PE6ndU49KLhfBYhaXgrlurHLp6yBMeoJKRJNJ1/o5cLucN2
EMuvUYDAUCn1HR9IEhGws7Un6IWpJlNn8Xee87ksR7utBuLfJRc3x9Pm7+Kg1GOl
jSwAJeM7a6tSS2mNIxhT72wF26VFBpC5ES3zpnvZ6/BCLpM+Ept3Ef4U5UxSt+68
32GVb98o3tsttStiCFcBBkd7OeKQ5hABhTSgKtdcKBrGlDcARdZtLgG2uX3MEKmN
OsjhK9M6NYuqfDZ33EMgHWYOcRyRyHyA9p6H7385qWurWgnZzeL5WHCNRSD/KFvz
lrUtZLa+Kgp/qPKj7jXBbD2tQhjNkc1qazGaMdbEBakzIuOGZ3RFj2eJ7YFEDIaH
0AU+YRlLCCfzGViLn6fnhWyLHKyZlEJvaHH/8AAsIVbn/0rJkzCWqXPPMbwyw6HM
rZpZlpBOmQpQFRaTP4fkNyhOwxZ4WgEjSDpUPcr0WJBvWLXsaiiIc/k7TPAYNM5h
zNIYrYwZFpI9w7zwkmZzixQ5IxlUFAuC5iMllbaUQXfyZb1+CGk4QqNkEoiRUvVM
l2RGLP1ecfFVSWeJVKJlF67IV85as+DzNvgw0YKawb6vPuDvAsmVK1b7to1ccyNE
Sa5agL3nRcQJanWGwwQVrPFicF2z1ALDGsUNsaT8nrp4V9idVEWOi8g4OiQMAAoQ
rSdPEYbJfsaggFnYaetsM0+RAI9UFCd1zNW4ZIlBR/rScxGFW03wnr15Xko81lV0
iOEFfcN6NylKkIi3Zo8EyJGtNYL3+K1nf6xA1rYP+svqq/3JBL/o50rJMXjaELzt
FMRI4OIv4M1LmoA3/kYN9cGNYTZI4akNBJB1YRWYW9HrdJgHw6rh6PPOPHCIR6Mw
UK07FtRbabJHmEGhhnqQ1hCi5aI2XH2yRVOJD3skvig44fzPtZi2V1IfTt3u4gaH
0gmPVenhiLf6KRi2HBhWfmAwykmyV7paTZ6mvUNxMmDsxeSmp+NoIgxegGtHZaB1
mIt0a9ixIs25IvvEpN4ElAfz4VvVYpt7usJvDGal/42Y1VSvagiX9LcqBAEMMET3
7dHh6IqdxVcGJSdThxrn7OwKGXeABzciCHD4ItbEnHJGZJerTVvldz7hsKlNticJ
yf4SZWRGbFuJR84nIxeHsjJJa3AsQFx8WsQ/mta07cy8IYRl4yf1Y3Fh5PN2E1qU
TIRN2dk2vA7yJmAu+MxQ08vKkjVKtRdJQ9sAOujzp6ifwQUuMZp9qQ8n0obek27c
A+WbmpHewGx5RgfSggrYJL/7JFaDdSeYi9M9rqkuhwnD63LuDqDQdoHoLZKbgvsM
zQ1lr0DNmmbdbmx2cVB93IrB3fgWKo01Lfz/iKipM/MEoKnwH0sObfqYS3oyzeJg
a6v4BrBTESX7jdK3rMIOLv1fAYyEdUrQR1agqynkaCMsxL/qMqTvrQhyncqQggt9
J26pcgpfsx5UBZ5FoS1lUzi6N+956T6ZhcPkF1O4lla5ATR9hv6IvZx2t1QJVpv6
i2v57Axc1cseqBN/aPamwVboclR/ISIkdbxy4MemAv4myaXl5Rw62IBx0rv3h5Ax
/e8Uzm9kf4HYmW3mX3Y836wO6RqGbB5+Uj3qocAcLAhM0jFihPc4RGY1SN2eBKVJ
q6auG0XbEWzuQ4h0+ybMDzGytHzFPXMTqWHr+uR6/x5XscHPEchFyorFiG72Sw6f
9XkTsIOzgHqam228TfOJdWDoYzzBIPBVhokM7kscVm6uqU/lmCT/d63bAd/LeCle
HR1zfm/Ts8AX7oYpH7xhFKKorXNg7QdMr1xpdXrcAYr2RPrg+1rqCpEyLbgSBsNA
MKQvDxSyZiYEt4zJ46kNP6cKTRmg2mnrxPnEiDDXUon5vAq80sWVouLKtxgvSyAC
ilhL0w8C/O07b9O4SCdqzn8nPNnxL6QvlWqh2YfM7mcWQV/32lCFdD2NOvdERXQ1
Zf/KMI0DpBED43eaWRRXR0hsVmOkH0mHLbhUUMIYnGk0O+lYW74c7K6IEtf6zG96
9cip2CIWAHNPJGRc2+KRakbfBgLdlE0AHu+aQLU54A9BrWFn26r7E6fvOFrtMujg
LiyE1n2yvA+4wBiAcbzg1CWhhSpRe8oXQzeL/X4LJpjS0DbaMctLVHn0neXuksGG
rnNxb4EYUj/vaHj4HUpyo2e4AqyvJa/ld5T80mPFEN0KvGzefvFJ1Bm+GupVNiHb
Na94Q7zNN2XFAFr0Ci/6KpOqWsd7qu0ueF00ZLI/3+NNEsKeBi0sGk6CYoWxkeVJ
4KAR+CHJULPbHAbNuiTiPxFGApxFKcWjJ7hZBovLZAwoUZtY0aTFjKAD17b52ZYs
MophDYlfsNlS7tIBreADE89kiBwZNM7Cgy0m+KpKnZPoHAuxrRo5ZTeC1/tz67GF
+48ltFxoFdsk/S/DgDz4ZJHRXjWRQvSMjRW83HDhlA2MbiS8jubO40FtcLkovPqb
Yse1snFrheTAGAnmKz+bbno5I8DSmkOla5bqAWNB/iPa/s5a4rlMoMqkKaDbLiWu
+6okjzKSd1ncMn/t+JUdGBIJ/CbOOt2FqNGDtyKDBkF8dfAJ+9v3Eexad20IA7Vu
8ghdkq4+yM3SeiYGfWWBtI6/bWTO1nkCvz+fOaIUMhMkIZZYq6wwulK+YSk0iO/m
v/skrWxWj/F1ibBQtZY6LPMVeIAzltX2HkL42+pgEzzMSq9pJL7hgarMpTfXdj3p
wvY15tKteCOqor1eY5IqGWNGobYBFWq3oFFlGz4l8MKjDhYiwvZ7k4JFqgDi9v+q
7oQBgs1WPkMyi9igsTB85tOHVMvuydz1HmD635lEOWDjCfb+gx17rXcDb1pcEdJf
pzKhUZjCL6VSgyOxIKpVXXBpA7XpInJ4snKAyatFO2C5YrQ+YnIqJ7tlFBk5jzcb
jRlhdL9GMp/ZtVDoF8eev99wJrQtrPp9G4LNJRpm1OB0i90MyeI//xym/Vos9o9m
PcYm9wSgZh2GhrIJja7hj2n3r4537z8Nof6VItxWjcFhjZi8esU5uIJJnnahkDs/
1YGFgEvfKxOz7y5f5grJUW/ptHkJo8S3KU4kmVZoIUbdc4k7nafIhkPcllM3piHM
DPPaTReF1dr/vctd6ELcFmlcolASGR1uZOYRoTYTB92hfrtLI8TqFJrQCKQ0rB7a
Zp0YkonqWLTgMKOMYwz0h7wN6TOTy+WXO++0cw8jdRID3eJZsZc+vvhDssxD/3PE
VAkHBT+JeuMdMnq1lToVhtHPnZZg0K700tcgb6K/sd7UEEKQG/cDjZlMstn6SIpR
BU6E2jTBjzQYG3bE9ANsaoXlUCfoKNrVFZrlF4PRHFZxWHcxOLsvbvVELfyU812C
pLSOiiLUztCAXLM/a7ERKtiRpIPWqk4KMZ4tV6h9EaLGDTOIXlO5YmjfOzEANVH5
lJ5EOKacCOjcD9D36JiamU62mE0WihAlQl7Vce4KWK3AmDCiZIOuVBE20oeOs0FZ
RIqFmcc3TBvHQ3+SMWSFSdlEjuFTEVLmfdJ/Hs7Fs6Th7vsphnUMEI4O8c0/TQ2K
qrWBKeNUD65sQHBzXZWXE/cTUhtl9/3w1DrdvNqqrI6iHxTJhlO6p4dVocB639W4
y7NOzzrmHmBC+W5yrXvqPGzn1Uc4SshN8arNHst61kI+yfoGssuh90jBJZcHSb8S
trOFlyG8SEPbipYz+9O7hqAdZbFK12sjVpiAZVClcBjIvAhd7XFueTK2Ch/VJLCY
nrRK3o6ebjt+1vgniLidwRWGVkr+dPN9kxa1+6Z1laWKbTWrGq7zSbOn/A7iBqWD
YKZKcQFyql9slXd2tSegfYYclyL7tPzp7Zng1g+PDBhlemusBgl28FNMy3zByse4
cQ89RU+F0d1wkJi6K0PDGZLNyBurqeF0f3AuWvajQB6IkvDd8eIP4UQaKaOsICEn
vxEO3WF+LAKn9wswD1d+lk9XG8uZWr73xqvLR3Y1UpfbCtAyMxHPWA+fkBClBFuF
/vr1Ky/uSS8OD+pzVpBcYu7ODo1ourZqSalZCb03PnYBeiBT98oZIf+qQbjkLaps
y2Pq/hieFD+kFygyPztp6lze5i6uNivrQHW/zgeVEutEnai7lh7ID1VLWwELDwAA
RgCdLL42x6PecYAP9AS0aZ9Ujiyho6tcEiyB2L22r41be9y1/0PqPYk62jnzIeMP
khkWZYree1n1D1oUt2nWRpWhNq0kW5Jh4o519E67DasccgbUnCOTz0t9w7GoOEr1
BeSEvz1wcPWzBfoSoyvzO/NnAn4ckCtWY5+bF47/xrk/n8HUwzCM1mJRXJk1UU6x
cs91vOzBNG7Ikj2Hxvt+4D1SjC8kijA3WqoTHVsRDKhHlPOnLxuBTYXbN2nUgeM3
VXxRV2YPbxjDgxnbAXOZx7a1nW+qjAAioLb+zjJcJBEE6AapPJwfKqHHmvABn+Nx
xd7oZl2l8Jjon+gLadot0C12BNPDcFhwYPp5GzSk/c2WEyvnhdO1OVU4tRQ5jrhc
rYarPBV20EfHMFk2SGIoH/VZpHim54U25Pzmk505kc4/xcVEcnCAqoRe2G5ZBYFx
wls7mAg/UbdxpoPBigk+BKkxyxZlBf0gZpLfNtM/KQRtidKJ3bDXmNMKTtMod8CC
sVeRDD06AZTqTHqesbmJvT5yBg5z05yj3TfkzShOH2pj0RDYg47ZzHP7mOS0U+Hm
a31L/ABX9qiiKXykK7v4a4XIbXb7E9Eg6F7N5RsFNZBc4Q2ebmLnR0MtQtuKLhy9
J97nVXoWV46+ZKy+Le1ILq54G6Q2LyoRTygSnvdtn4F93rrPGSneXa279cCpDlNu
9KUNNliWc/K5N6TbV5qXtH/Z89aX28Ja7SnRtXd2R3L5hwETM7FUP87g+2JvbHOE
AF8SmOghUiGB5PNGX2sb2cwnlE2iOmFpphEDehca5NVHfux4eewJQbpCzpXeJOdg
gbkFyfaFjsm1Ei5ibmOQdTOLG7ocyQtgYpTGQLrM0GzIiHBist1HzD2hDzQhebKQ
13xbXRdwJCCPuFXrrRVyG66ceNK9ZRtO/wHOOviNAkVHy+Fq/8yS6B2/mWKALa6R
9T2rVsqTznV31XU+OP4RqG4BbF9ZnJblCT87nXG7xstKEOoq017M12TSlKb4eIL8
LRf1jjcHFYtR8j3g12MwUAIwId8PEpl4UwnEtyX3SSCLlKwJi7zVrvTMwRp0O4BU
t9DPnqCXoBErF7P8zzfiWkk96FcTe6tEJcBMc3BN/05HrS3BMe5vbS1PkR59oK1A
WpN99rRTPymPCWpXx6uDGhpVIXgr5m/nB5gRZu+TNNEIcrwb4rz300MXYP3pe7ZS
vqhZCbVAq86wukUZXStN8y4IwDf7HNXHFCqzKAO7v1sKeVUS4FqnM7RYNjk6al/9
KkgbaImCj6kDmfilaIY+yopYV8t3M7KfE0E2pBvNFAumDHg4pRZ44Ve/acLotQ2v
LBLyeUomHYxlGcZyLy1vmcX2DvAZgWGEaQkg6jlY+9DEmzXQjYhFBpmTuaTf/h8Y
5AqKCQxjL5ulul6FdBn/IqckDBZloTntbL1qzVYQ0ddDB4Bj3ynsCzZ9bphmta0Y
0v1f++SAaLfY3OizKGuOR+Hjn7LDI+44c5fMo3pY6QR21rXIEiyqntxu8gfsJIdJ
khWj0IHkya2fpc5yA4BMhbATElLNH0EtGisNVgQCX/qKGpUfvHQ1f+S6cuP7Zz6b
k62w/GPloIRGwuWj58UQLiHcq19f7mI6qzMGlAs9O16HW0lnNtG/WrLfrnbXMzGC
ppbbUN5/wWMiekjX5OqKRJxd+Nb5AbAqlD9iSXxvXskyWHtN9Untp5P4Iv0bdKBe
KOAb/iXkUBFQmw038KKmwOqagvGdznHr1ryMUmcO6HkULdtGDmbJ1oHFpYnUP5ZW
NchNiaXs0NFO6RxWTY6kdejy6DTUQM46WBpfGry9mnXZO4fd7uGg8Q0RN1RykMPe
EClH139yGrGro40CtEhUvLiykza/Kj7gszjGHTj96gWGAmnY5IOleOKqwKFXVjJs
n/qgcGn0tQkJbEnTVULCaGv1gS7Ua3stKDoO+5aSFWEmTgfKcNnSWxUO+1EqPVjF
hI3855Yx2bb3DnOlqeK44qvCpuUinirQPeJkH2bGV9RxGFklkBD1gnxruhWGAmba
I1GADyJEAiVk4bHdtKLFfvqMtqc9RKkpjrDK15K/BfxCZQgvtX+AiRqK3lf77kRe
TlHAQ8Xy4ZQDQFMQ14axHqrfiDGR0QFp1AQaZ8kEDLtvrc1xw4inK8kjW4gKv07x
Kgt1rbtrZnrFk7mtCBGCCVW3kt1Jlow3oBjRNL4mAEifqFcIE8BsWQch8sgNJnUc
tUxJcXrAjY/tZI8jMuUnvHHoODl/mnfInU8nwzC6fNvAvBn9O+fJkDrbsYBCvUXQ
dGvfdJ660YcjYm5yBTzsuzl3DW76K3pT4OE51pI45p3uDAmmWkvaN9D8S0pBM98o
qO7Dfk0xypY4/dcMNkfYgXwbpKg4k6XBHjIRiRZVKylEReU/M5ubETvY2Bl080lO
v1Sw5S8N7MhofnSpv+9jRaixIELACSEb1AnfY2zsHkyTQ4ywIUgzQSus/Eni91dZ
C+ZGjv9xU9/oOLUi5gk5SzLJDEWL61v0mBovjoBw6BoTaaKIpWWrnxr1Untm5EvU
CcC35+ub44rpozW35AG5caxB7vZDMSM/EsH9SzvbXuPdkAl4dlCqYoEC63pFlnir
GkLn15Duw4vnxmEhaqN86J95Eg5WVb1vrCXdCd5iWHdTt1q9buQqiP1mkEkhQLAc
9lVU7U7UN4+OBoJrs4JtnqHa/eyMPM+9h1oLv4yr5Bf8qtcwAgZ/Tl9JKpnGAZql
hmo+iLSKYS/7a/VanEGNTRWyliXtJq4j39sPeBJVVl7iSWbblM1cfptF/mlKVxXM
k87FQtZTIA4JfN+txtU40XROEzHZOpuKe5TyT58W1Y4SvumNtPEbxVYUcuFCqEnR
oUDcSgvZMTD2MgMk8ZNgAm4Co+b/0cPjK7j1Hr+RPcOsHCVqkb9RWkexPunjlNxb
Dzcr6eWIUdFKndQsojbiHQ3cBXBF0jYdmho5SfTW/c+JAZMQKl8Oj4VvIUtqqDyO
xIqxQKP1QMesOSKBHqoOJ8Opr1GGWknvC7gv/QnvzbBwSzWerZSxTD0l2GlkdVzO
D4601hYRJTq2y0Uy1RCaETwyf0I9/NnR60u8R7+jLnBwmEWh818zoGnXX3zhAwjg
SfPrBfEm9axvSfME2Jqa6nxq/S4H8pmACU39mA4BnVoCdBiC+6N0Hf6wQ0xyMAaI
1segr/1/ovsvY37ULIMX8wZMF0aoqdZYG/t5j2M+GR7he1/Qa2eSNSa48twuppLO
Dk3RWC9YwiPQEOuWyuSllVdupl2dEyy5JXRCWUAMCzddxDKlAPU3MKh5vENqqCE7
SnGfCwmUMi5oSKOmFHxMEmQ9+nHmNhblYQjpcLx+Cf9ENkMYIgt/q+ZQafsywohc
i3fqdtsrT5izac66jMa600AWxVCz6xHWaUmcvy/TLYHj9xEpNePnbUtK39nNLU9k
hT+H2ZyrQh/Udjs3lX5EcQGNhOgPEm0sRRvoxKLUkWLc+xTRD6sswaWyP+sHovsd
rP0/H2V4IF9PtUPWG0h3yGZMkDc0yKkRVQPZpsJju9TD/OtRSaziF2XW/tX+uAcr
9tlEAy4Pd9mdfM1ZLPBCookcPMez40O5xiQAkBoSgheAh/bXImLpQO/qzrSMA1S6
w8k+TdP+A4ULBhQCOkP7l5ZYElJSDXhwPJf10cpiUiVYn9qXr4vkNIixzTbz0oB3
OMr22TTeet5/Cvt/7sSDYDh2LShHZ/cRsonU6Ve8mB2xG/51Z3GpyajtDCH1kuIT
6tmQpkrdUo9O3Y2WlR3B2B0B3yZy0JYl+/EUiR6OaZmLxFRd0FP5Q3Pxt5wwHjOo
eL5tDPJL6sB6liwtzbQKAaqJms1uY/zwz6sLahEsKQws1ToF+DSzprYdz5EVl+N3
NIu0VnSpbKrfP/cVdRGRF9Z58MF0+DSdnDXR2W9ehp8BiSfE5geLJ9rfNukzaoMp
JY1zUhkwg8dODbHIrjLqfgpMu/qZCVaoHhfj6mJDtDt0YIqa1ybCewZcOOocUmeB
EZQdPykrMdRv7tpUvng+QZ5TaSMH0gHpJqp49fLkaIagd1Df2072oH/aNpzevo0l
2USE64DKZzbT9MzCkxKWxFcSfurIA4PvLx+O6n4P2YkxO7ko5xnLLWKJFBFAYNzR
i/FQPN3mpht19Y/oeqEGqp8MfFSB7C49dulP6FYTgNcg3YRR27Va9kYRXdRiB1wO
kJ2IFd8liATE+I958aVgp+7vy0szsJvs6sP71UdS5XsthF4QlxXVDA9qc/0DzHBf
w7OcsT6pEsgFHqOVEGkzsGvkKp4/DEjzOrp8JU25hzRVygGasinRRMDJpusR/nUf
xGqlalh86jmkDvVsXW8PMGilOZ7ptLjwqV/JHSCEL8NdIkjdHvIr/wEWJApziayd
85guhv9xI5/j20hX+LpMW3H3pFXVwHQhPMq2wHDhi1HWO97wtaBncyIOD5sNnhJP
UlDTmC0h6RPLlRJs4R+GwyxbAMCVg8ckzgfecS9+LUMPc2s2QUEegz3EF73iR/Tc
1M4ocbnf3U1LbiCTrIdKao+6fhsS9RLio85agP6/Wtrh72G2COTNUct2ymOtnyVY
N15XG9RtLTadc4tDUmbV6PRAQ42NLPnKJIK7krRKHNsDCvTHIMeQO135r3g1O1Iy
D0ujzvMFoAgLLJJYWr/tZICJRZUu0Q50y9M6BdHp/cQm8CCEKOaFo0hxC2EFHCs1
op0A2/+YjThqmCH5wjXiJ1LOPb0UArN70u4FzLDuqjlU7nPFHj3Pv+TRhrKZZg6E
jFsqEAvWVmq2xGeaF70jLIcwfu5NvT9UYC3sU4gj0NZxPJKUJ/pCMa1a5Xj2avFa
ZAOhQ1hQo9RjUlSTLWRfipx7204J+cuv9PCu59AAHYIjb6V2q/MWNHH640IqtBXL
TLWmOQ5UPyAgxvgEDDZteb2RB4YKi5IeuhTa85K63whliydouJDzGIdLAQZCbiDS
1EnqrL+YCAV3DUEyzmF/CpeycR164DsMvWKJbyM6PLuqC0SaZueOhrxgJ2KXU7jV
g2UVCgWaK34aYJLu3LTaGZ4jGFVP9NWd8nCOnwWtiCYNVzkK9AqqNarHh9pJc8Xv
L/Ypz7Y9s6bFv5QxaXdldS2Rjp1sKWeHxVnQ14hvKqO3eYeMEkaynKL6Bmuc+zW9
8hLY/y0fxt8DCoVeGC/g0sL7WkDmvE6j1p9UfmPbrrvLLFvJvDegxqbtWA1HV+ke
D9wJmfqMHgh3CtDip7Ae0MFkkHD3Kvd+wqFSOB4AlJRmlcPkQFtI/o8reH1M/jus
u2QXGOA24EVmyixM4PujvEnq15VZklu7dmFFL8yXlY1BptQMmaU396UrTpuSvu9E
Jmleg5aGe+FIuo7IX0G3j65d5l7w+HOYmQSvEfnCloULQIpR/WqSReQ5bmwsUrcj
OfcGO9I2afzlA3JgKxd/yRQuUU4e3XNImGI93I3fwdXhGTEga3ImsBMLjexZ8U0O
hHj/gzGxDwXIwInWINBxXkkOhFI890dtYGjgk7RuouyBNqLVxd8Jo+EjSMw4I6AL
ZienUJnGRFMG8fMFP6fYjM96+ZTroDJ+hcw15N783XrNp3VZbEeAUBYQ2Sjg3B7q
oyYmf5t9UPCHEErX1woI/tUjRiNgVJFBeDJWdbRicZrWUBnM3vKoWqkfSnSRIpbl
F6AGF3hYhVgaM3lQ+eftk+7pD2YuR9D1+HWJtBwsDEdmURdtCajDPYvgoCDkuwta
+CWKbKWbq76GROBttIrHD1Me28PnuIUAFrzUscbECh26dXW+ll1tkVA94UUgo95Q
XjHTnbHPOWkA2xXkFFuHwa1EJLlOMK7AMFeod0lMeQWRYovQswC5CzDgcjmjLABX
4cfR88QrGAV09y1asnrJ90ELOb7pxaxGSc+sAQJ6rumaegf7dbPlUQUBd5kBMlb/
gWtfeL+HzJUyvqjkIyxkWfj9vRgFZ/EPfT9tsPQ+HDOZgUsUhbmmukKfQoKr6fix
iH5TtZKJYrlkeEwOgF4QUp/Bgqd99v1bJO+1WTHB9t0iBHT0zf1orcDuNlrXM9na
N6Um8hdygWYLY9L+YAFr29TfmO/lYlprk9zO6Edp7ZfG9PzrpO+/ECmIcHlhGwVS
LLxwJ+U+htC0cqyyHaLxm69XNvv7VLtZYd0XZOzm9NAIyjEkla5J/HRf8jvnUGxT
PDcgn5E46F+6moS574vWJRb7EcSnrJV5s0h36cYGMcbc8k6WIgMmkRsK5OHN7upe
FMWPAfLRFjD/GSQrIXJf9rtV5ieTopjm8YiC2KAwolPIiSky7V/qoNEwGXo5Neqn
0t6+tGBJ016x1ZD+4FVFk9pjPv/TYT3b/2dIRosNOvL3b5W1n1ZHZe39byb/Wsb/
B/T9JwVTi7aqfj/iLGkQnxn46stBeyTh/7d+VbTXUx3zN/pvQWkPE/WWqEwnS+eN
d/SRQpF1l2OgnUdNgpX6S6PgPMauYLmTASCDGQgujsjAxcceA43PFTBGJVFQCKoV
+Da588G5St3hBJsP2xXQapwUxxn3+QxcL/fHNFi14Omo4nnDS7NeibuWZkpf8HP2
rb9yT85W3zu/kznSL9UAVzmsJ5pgceEy6lk3cj+4D4byWLqplHufc0BgI2mbY3Ni
/f0ImNkjc55atQszXq0BfoGtdYZiIYF3X/8Bozj1/kx1ZmYT6nsRxq7DZDEWU2QX
DG4it+w6hCyucpywwg6z9mLr2KQwA486P6EER7HqMvFHf0Wv5dW6aj+51ukBzbAT
qNHQ+tKDtfwAbzTAdlSNlycgR/dUSm51S11GnkQOgZy0ZmYiUgBCGdXEDC0HUrGl
e1IsplSIqgS9RZLNpfPHnCtH5zEC3YQv3CmLf2qPWZ5WaZBiyFZFrEIErQQwNXJB
MKCokQ/C/yiQbj/JQFvRGMH7IALa5deYoK2k44njjFd0+24JItlosAKlVrbMv9KV
dh5vxftK0HxubeaSr+gndb+fibgowmsz1G3JeIjC6rwo7X7j5F0XWnku0jt+XlAu
bBDcyoDY3pmm7DhahsucuCaRPi8L7oPuf4+mrAJoZSUMz6suO9Lwa5gN7b9P/svW
ZTYwnn47lRY3Cv/gaCJoHx5ZhJxSXILrBkb6HuIxmUVRxsQG8b0M+8eT0otgG9Kx
jwJkd4ICW1bvWOYiDPDmIxHZ8j8fINwIdFPYthuEuay9bvZipSVUCp/Y67v6zONJ
6XnjMe3tiMG1OdRJ2b3HAt6jxAFa1ly/RGlee57ntt/thq9jsHOx6+h7gCBcU8eb
bIeVzOpy1e3j85EwrOMv4VYG36VmXUwu82sw5HmqGiM1HhHFeyPTc/qY7n4omYJb
SCvWsBbzVDb5Ah2pj942YXK2Y8MqubwoC84ieBl/i3x27/eNtOOZlRDKNr69l8e9
9tCmUNYp6AsFyxx3zrfkPzrrozeRh1Pwrtu3MFHQOf8VVtBEo3nr94KUa9b0uxy5
eyo5tGKrjg/KffVQ8/c+29IaFLcOipfappuxycctYNQaT3RcoJxwNmmuhSMMkLdh
Vfo26nSFZq/FsQWHazGfFlibSlzYndXsZcqpbRn6WBm7Old+2uH8ITa6SwtJBCZU
FH4My+JgOYPLqPa7UrvPgC4nn2w21M67COg/P8kvMRLnCU6WvvxivjvkTKRp22jO
M0xsj6TCa9P68edY/tREObT0ReOj49WD9C85ZyaA9yTcuuh8c5C/UcahdS6q5umS
b4SnAyjhSe/LZHkfxoFSpWt6SHT23iwIfkxhCJdj2k6PvbmtufAzw3sARMc31fQQ
DMuwjLzgofdJlhhv72zECYxI85s1N/7kk/MpvjoKsZ2uAMPAK7sGLojOtzr5WFhf
csGjmtlsUSG93oilyPqEF05G6Y3LRMTvfGliheIXI8mikWuI+LlN7kgqA/T8nRGm
63eh/U21WetocOonvr797hP9pOVXi0VXeAe6gD8KbkzuI9verJLm9N8jTNxhbKR1
4UuVVINFTb9Mqhfc6ciUC5FO27oD/3fLkTBnwx2q8QAzy+rszAev7q8wtppFkLw4
K71lIF7F6JzIz+am5FuAXh4dSZzCDilNHNOU9/+EQDURjo6cVjSXpf+XcEzy2Yvw
MM4pFjGQrIDygnhB9fbJhufop7AhJ9sguLvn99oZfmTRQm9vajfojqCiyqoO9rHg
hgpYu6DwxCSaqSBFFbR3EiaaEd0LYv/OIjiGbA4IyHC3x1CyccqxOINYGEoKcEfW
a9SzHBrUNKFiFcFHfHme3o4vD51Pnwou+hiMpZJPlOKgNAKyJ3bKXmfimxILKXG0
dOtHdnhP3pO4NmnA3vgtq4D8GGg2FVh5L3GgLmIJiVQMLXw1DZ5uGgZ0WVlwBcdp
ibLU0ltDoI8+1CvGkkOJyLWTpQqEzLYESGhNRt9Z0HzQKxF+WoMK86ckFV5t451v
yDMrXz+DQsGxxR3vVNyDetEIBbxE4Q7VYhVmxDwPdUEmSjF8+qmtcQ+STQpRl8sF
eBNbvnLEFy9R1PsAJdZdpSunWZRvgIwEerDGObn2hLarKlzAH/DVpL3cQK/3FlTT
rDntAQwBSWfuDB5s6ZPvtCqrbw/5eCknWLoKXOGqrW92lc9txVYyemRUDlllX5PB
D6zPs2mwAwVKaPlK+5m4C/qyPeOlCZjx4i2zSTBaxhz2cvHMuQp5jq65yrRb8cHv
QvqFpGxmp07WPhO5GRcmKJ63W+NIlKprTDfDyiNTBg9vOYYG4ih2VShNbRqYbgTC
hDIu6WbillB8+gfR8RtKwmj5hTkXizmOXs+MPzGc4bT6kgLn4BA9QMh5fOyUrtn3
Nfa9c8rxaBAOVST6FT5aDUgvlU2sodMCYjraZp+dWHE/QastP/s6bMghBDmxBuj2
Wu+RSMZMiDIh4mITOX7tgm+dCJznVajz+XFFkF+ZFtL8+E8mT+Ia5a0Ugg+58tyQ
lX6jcHNuYYXMcNGQMkXYJOQevWCCcXu84/8JnzoH5Z1q7UBxj8sW7CtLeQYImyCb
Ao2yBCpbZTYD+6b9kOyyO/Fz2p9MqdOORke4yMHLdiln16tNCEq7R1K3O4J+frdO
Os7Fzi/eC11ryD1FqnMqu1oH81YTRzz6qJxeyUjK/Ryr4kW85+MqQPX2lx1x0uuv
QA/wsB1PxS9+yFFEWgGVfOPm68uNTr3FGUyK0vpvpjpM17tApjfrnY1FapdOuOZe
pf9Y/t4JDiBGsz2LiBCCyuTWK0AFmKKvDkvVovtD0iVv3TiqLzi4MjnLpB2ZgGAF
LcqqiUE2Crc5hBuqpna90BNVfC2FYbc/O5aHIsjrIbv08H5BoN9nBLFrh4AfEY27
rOcBmxuYT8J00UAW3QDWhH3zPgzcsLnnq2q61oIoQMpi19x4fRVIMDxMdemUyrh/
pVpIG/rQWeyKXvqxDCP7zHCTHc6TooWL200wpyHqglRBhuicif9QnMvuTHxNuAfc
y45pwESjxwdf2SNz+csUAWk3wfrcFkIuFQiRLfMsJ7w1ZNIYoS2vtPxGFHNGeCQA
mgX8wTLZOnnw5JBr7U5SFWAKmq4q5UmSqZ4ohnAQE1Hcbg+EdRWCrKzKHAb6kc7h
7LjSSIz/oMRnv08eYYY4hvwlKCiifAiy8+BuJyg6gyM/Cj71z/fAd3UO/I4irh09
QW0z4YkD2lJxaNCPccWuJN4sSDBeRW2s0dk73bNCyw1EWcXDzAojOrRBStXGDxVg
qv0FwkO+2Ouk6sNh8J1nx6wkx1+7Pa9VUgWX3BZ0dKZbLwh8tUj5eO99aNlpHoJv
T0YaNCJzIedtuvOxhCiMIFUQ3ox3lxCyUux/3XtfN+qmPRt+w0GhSi81FBLi0a7/
JbXBTBqBreZnJJstcYUJ3MnmAVGiXFoqpZ4uP6TwtXXqOxmaXk9ThsEB7z2bs/+e
feyUcTclGCGb0o86nV6q7GwwmEjLNIQ6FzavebOFbM8O3vmgJ3i/EEcCbtF836LK
NYunTh35U+iAD0GmynWKNZOUxDZtL54jy7eErX3z57p8YApLOWKAVKTuhIcom8jG
zMefdOoy0iC5jVc3oCbo3/GzwtIkugH8KmFsMBPSwuHf9SQv2Vl52nG+BHitc5LR
TCDZgNm/YWIqcuVg8oqJh/xhTsRBwMW5BHZ9vVOlJilI3TfNL9dCywThHTGFsur6
d6sJaCENhmULB65A4U2LJ/eJ9ou0/F+GVffkYLEeYO1i9eQDM1u4Nm8XHEJ79l+n
C8UU+Wva1aiWIu6VLwrTpZC7kIT74WENVJrggs1FkGj1Kq3gszkHEzvE33rE+1x3
txGdkbSCCNRsbs4A9D+ZckQ3jGN2BKo+xWHUvhUnAuF22VukZo5px4lGF6k0Gk4O
9VSL3Cp5L3OqpkhfSkfU1mJx7RuTAPPxuu1kFryINo0wF3E9GfLm1tR1bzS2oeiA
nMLlmXa9UNN2isIW+lO1lmWJlHG/+sFgbDQkO42BBFJdAGPsIVQphfUA5VbR63bh
B15kqkZL97zXPjX8PCsPcnRDYSm0j+a6Pnqiq36C//H+ZOX0Yu8M3uEEoMcxzY06
kzscpHygsqfx7pNI7SiuKqKSmc1DYsqEs7do2FT5HmitxRbb3w8YgoCElXAQXo19
3OFFp4IAOSfUC7ER/+Rtn1zWhXwKTFL2eLWYCz1ZcngItwIpymX1cxhfXn7TeLL/
LJH4JtM6WSEeRtgGSqukvGqXOdEoslqPBPZd4VAIo4zJk+/v/zWftRCMLc6NxJlk
xkjzSqq/2JU/zsoSHMyBOQvBceu6lO+fX7vGmRB8XANQIjm65a8do8yhZ/VkItPL
A9uEKb7HZXZhuCjrgXSmkWJo7ztXgMRPbIdVhb5mqo92XvXBYiLuLRrgP9IwbABV
CcrP2QUvCAhmK/f2SPBHlDdnmcx+7fDWgNhZXqggGgq093miGGsQouenWlqEb94V
uwhNf9aLyWnUd1LuTGjb8KxJmem3YPWf6J2CsFNHlsCb1JCeE6En8FAQ1imP0KpM
mPMaUOnMDTDaxyUuiGhUj+CNpAonBzn02N37HCnM6fkEoBpN6GQnbWAgJbwyAZWW
aMh5Ypm+4U1D6CHmQoJI3IbtQzOp8LGFj93iEdWWDWXBzUnFucMSq9bfyTjjC2aR
impI+BrBILfeHwCxwsI6VXau3tYDr17yqd4w94CamHhSxyfMXYU/6PAYwBEtHnEj
+tnkZrT6dTFdXL4NQf8Jkw8ePFIENsxK/RauRBI8Bp7YzxbQOITa5vWYwiGg0xyw
pyIfF2Bng18wsgdHTrAiKfbIXUTfVU4uu1VxKuI0iG4nkTmabgvCKb5ujr3VKUIn
yhxXvq3bWt2r+GVCd48q7wQR7jWI0y6si7AVUgW5Hi6qCeEEMhAQT3hhakZEApoS
uoRd8aMEn8OFR4oLgi3gdd94DgaaQGygfBvrbjEYJKBdX45CqtP6yKQ5tIIWUQHF
ZBSDjH4BlvzP0a8WDWuUoaqxqyIBVlyXuxi9RJLPdrxd2iJWOcVx8iG7ZjYHQbsB
W8EuK7U31+QZaJTSubSFXkvT1oDzwbB6OCOJ0QSQCDFdMbeKKe2n+bamf9PJldNj
ZnKScQSqinXfOu1KV5yCp/Km60uX3WxafL0d93yCLGydCb8vzRF0KZt/1JLYbFtA
tD9AsafT1v5wZG+nqiCuJFBBvg4K8YPisT+G7jBqdnURTY9KoAu9O/rypprZ3BsZ
yb6Dp59bQjh+t7UMfSlbYkloGFN5gj+2xnKUaCpUoMm8lXMO5kCG38L5p+vOg5Zb
Xi8mA+rxZU6dTAUiC/lF3EeF4E54LWiTWTqhf2Xyibj6TlJ6XNb2nak7xqaT/yqd
HQVFiT9aFdv2VBpoLLO3hHM75hnM4jDB5e/pYtRLYKWvAXbkjr/96mAkCVOVK6dk
nq82gnL3sMloDY4REB+bOGkeVPGguP8hCJnsdr3uoUeIcSKZj0TUmEq8gu2eZU9j
BiSRVil0qQ2YP16GyF20qrM20sm1flibd6i1IWDLFndXwrNa4KPkN8Mby4oXcvZJ
BEd3PmKf7TekDpTpvIuU+xh9a4dxdwifGThkvJuHJMz4xrLtLKdIGjIJ4EBk83Gb
swRxUtX12xAudd8epP/QSmsYLFH+iKXmxQLCwGtXqw1oJSI0SV+w4MfuMrtJCj3c
FPiooQMcCx0t+6lzUGRB505Cc+MGkH8JmzHjSYe4cE+NOedTS2Ie2V22dUu9AkSB
RblxvDKflNmc9SRMtNTXz6EXQCsvjI1EgPd6niZwHeGn/z2RK5kjVkSw3lOiX1CB
tqYy0oRLRkMqOIoJjR+1JJdjAZTgiXOKfc09rvBQUQz7nxtiB7BZSsB+0EFh4hdV
1wzc/wOB01c4kcHmMqlt5/QDh2wI3nQy1d4lFeMZKZ+Fhmvc7MHthnc0aejUS/Bh
GMTZHV+x1Rul/0X60VacI38GxwKH0t1sgfjG8IVwFvYwUBQAZgsUB7DQFuYVQtn6
Mat5zLPRDSXzH9tg+Uc3Gw/pGic6zdEpbfcl6DekehjcKnuCIM/mCrqAmpn1vBYl
JGoNpEgWe/xceAI/ZldNW2B/D3O/LOJhleHTMLdnmeeBmt8P6vPy6qDqzRoyVK3m
ZZohk266h0R17U0XWS4v8ElgD/eAdkVB7LIHEYzy8jnAUC1bFzte+0hCAYr2KZlo
82Ocq8C9qvjV7WkaamEl9MmqQ78q3DcMDc7wsbXUGScvy24C7xqYARTO5VfvwsFQ
cnJx/aFI1JcTrolf0212ekKLcvLrxyg6xAi5cQ83yDkylFLPWY1WgeijwNMgeBUI
yr0Yu6mq0WdM+crq2MFZQ6TeNnmK3vBdcoNIBHz/Y3eZSIbXJ7qaKFEuq06Vt2mZ
94NgQKjwNel2CByCyUV8QXztJjvQs1ZThOcnjSL4bhcINDQIpApWwuz1skrII83F
l7GNamZPwcBNSdCgP9JGhCkkq9JSdU12VpCyOA2jwY62en2jbhykxNT62eTAAODP
kEWTVuyXSbQw+nyZNKl5z3qKFloc864ntN54xSqd7uoU66tewc7fr2dz3ZhH3r7z
USNG53sOvAO7tMwO+mGHn5y3hvP1kw4aa73w5dL6QLlQ0LLBB7bwq34uPiUTy5Ai
FEScw5DSLm6NF6oTl8d2uajbFTZkTksj5sweHL1NwxVVjF7zGcg/yMhPqj145x7N
K02oT890dX4OTmolZf72fSuA2HLRV3zq8A+Ggc9LG8nm0OjLbzDoZDOKWALIupUw
MPmEhGc0ChxIqeuAWyY2EEbFwL6Y/pnnTVZlG8lI6ai4DqOf0mmO/ca3rbPkZxFr
f4DqU3/RuiylM6APFO9DtlLmm6VBQ73d4AQVBEsaA3KpKnNYd0Dp+6lqMfjEEKlw
xifWmdR1Ea8Lca+krEn8VpuyiTqwijac9FV6WuAJMapXgpVuxQjebeEG7/f03lsS
d/RQYSRa+GYtx5N+pNpYDp1LVWW7GNmkHrX4ajvrwDlF4MnyGGn2r6khZMsvKS0I
rBDcsznsUM/1yMB1G4S9IE31TQ0HE6cO8aoVAogtLpnwDXFDd3Z6MLRxHgwA8aKY
8+OpfszNImjx7JVw4Ex8RAA6HKBRdnHwPeaUq00pVxXLAGAoYKsh/odhKacqEuUX
b8+lsJNZ8mP6EHaPz+rqt+P7BTfF2twUpY9xpP+hseVmihQZ6TgsJNDyChww1IKi
TkTVJSLGKqYO9xm8Hxa1i8XRbWgdF4uAi/bSHRRiMEeHt2HSM4y1LqLw7PY9PgPS
uI1EdDKphAe9HVY7z5sZR2k+dwV5Amasf35n8YSG0ZdJhkCpfqDu0ofC/7dsM5Sp
MRh8HBSjR9i88O4NsCwL+PXCwxsHZ6b73vxIr5DiA4uCZMmnSrh1QkZI8LxkJGCf
bIDi2QgRke+hG36ow6LLNCLHLoytzMbv2QNlI7fE3qG0mztp8VuhdyF5ZSuAufJL
YdPtRoggvzyGCTBCAD6cfDzSsE8PtVkZFmvAKEb5oymH4wGcr1wN3a76VD3tCowh
UUfDSRrvkjpdlAoHLpJrcMNtaqiEVShbiL6DnT+mQLk3G0P96zkbWdvmEZ/LrwSt
5JSYKxHA4x4p51EcFW6lvG7NzigkXWmqHrsm2C2kU9vKkiHoOaV+5I7SsK+8A5u+
+w3iuDWxWp/2UfcCIZPZ38Q1z3GCPCIOyj1NHSX+wN3xRn9CX6k57BA0aMY88EOS
iGH0l4PQWrJVU7qz3xwTE67bIdFvJSMjHktTZxQgXKRZkyaViBL/yT22HtYEib+7
WPL0ckwBgPxTxpp9MbLhZ3+t57SCz9ifxlcIFAgAb7SWAB0voXaOBDHELlNsY4tM
8VF4+l/31b32AN2+BzsIhCQJWG1X6+PKsqDYX2Z8S2MLUsZVLlDxs/KfliH5TBRz
oKMP0qxG5cU2Cgg9euK87qhOnKVw937JLKdIGs4P6zJw4ZsBcJrT5j+6RDZTuUl8
jck3JepjuBt6IJGMvRzwrR5rNmNjdqDoqMlDonEVZKST4BS5aiaEenm8pikZbL2o
Mm2FCpODYdDx1Z9Vm9horf3pI+BfdD/0yR1lzDiOKOMGLkY4xR/wpySzv6+ywl8u
2arFf5ApfQ2SSEXUe8zoNXRRJtANnLGuIFY9BF2jLyg0jA4DkzUFNXPGPgT5ViKZ
dERor8ZJAQEP+S4dt1h2f6Umds57q47bR29CDUfnGES93wrOwOLJZR7UAlhORGC0
+v9jKq9y4LuXC2G+qhoDJORPrN7k2BcNvkDxLPDST6QRIzCiKCBf3YnDjeSEt+Xe
9ncH6t2DSsksqzkVdBxvr11EgSNGb0YQKkA9q1C/qdThdE2lL9Wv6k1WoewTMmfC
DgMSuldOT0ZiPS1NegoA/6nRQu3M7mjUL1sXK8zlcjCnze15a+dwnAwTeKCrYfT2
O1m7HuZ1NtmALqZzqL9JcCXjk18Jd4sZLwATE9jmszwKr1HJi8fyeoBhekEPvG+3
Z+f9KMZmKV5fnaeR3axJlABB5JdpHEHDmWbk8GvFP4d8WyLn8dfLJPjbmS+swZDN
/eIHYrRRWTnXIv5gJZCID2BO+75SpV4Ft4qFHiDLZtz+HG2igg75zLHqad7JlADy
KN/DCd80ysiW/hxidxRkorYuIal3xZS1vHTU+ZlsfiT0CVa0ahrDqvwtUThDMc3R
uBOCo6f2xCvnla7aRtRj+7UoPyF8kd5tF3VtkzN7j62Qiufyi8LyO2XedqcutQqV
d0D4LW8XOwZcgIOLTt9Tqk+BGPKXlfVekSooYhe4LclX+1wqSw7CbUad+Pg4f4ww
Co3HlExk2rZGvq/XAfrEnKTiD3OtnikhUis+tolfEEgFdnULGsF2t7+j7hhWg/85
IxPzx6lOCCxLOyKxtwI+PI9tmLErZICXjAVM4eujip7KwAOw94gkmU5voXWEe3OV
xDdMB9geAxSd1moRlLojKb154rsHkNBENBAVDvpadE+eTDI50Y2XqqkYtAe8JxQu
c2yxTJXjQF0afEefYbH08u1OwQzrImKLMPTJ8VJuMF0QLqva63P2qhifylmPray3
GbZBR23QPxZCKV0jkTuUvxUgfYy0sXhTRPYpBuN658c8QljPsq5Prh5PRcSJA8K8
dx4WxXKMTP00q7KHMnkQ2zJJL7zukBY/Xi/ZsLwWGlkRSynThwqvIGrkczo1DTzm
5HMdqKDZYlYUTe0KywCZm89f6I3W5XgViveWbh5iAPSwoGi11O9IKICeIQhdMQEL
sLQy/kl8t7lYATCC0NZbNSx9w52+DBtiNdQB1EZGm0QXqI07PL2/EUX6bpeu8z+2
X8vF6L82m/uNephqaNs971MybwebYTkZ7UbTtWkUHiSeWVxuFYK1fGnfvh2BP6g3
jQIhz+oVtPYPiqAyGbeb1PDi6eV46xnXWKcYucxDsd3f/bGtWZvlMbjv3+zd5Vzp
PV+258HQmTVY+1uj3794ANXRz3OLVO37JO7H83tEvWSZDmLQTOoLYKRJznbHsWWR
4PN9vjqeSXgwqVvcFaPoovi7T/mth2bMFbpUMHDeSIcD7zqLcsxQftEqX/YedTFV
hipEoucCWGQWY3D115mevW+pQAmMkNKejAw7cbEwIec1OScFRdnIU7nuiYmp63YN
S/m+u316m+hYNuQLZrEpIcrcneq81Xw+Y8Mx4NiDbNYL3W9gGzk2xUbrLM8vZnTU
DeZ7VBmFMhwQPzUkVJxRkZWDnoFn2pKSTluvc4Ivj6uqb3fJjZ3uvfGmu1C9AY2l
DnvzdfibzF2ah3BUnvMPq+GTC8LGROcUcFbgyOkDToFM8HAWD1XfNg/QhBe9qRj9
DVdl61hbyvcGSZGpqoLUVm0oVCQv9l32qHrQ5A0adGDm/dc08l+aoq4nLaVijX3N
h2kISKbaNv+o2LBPVxSmQxvKsJDQspIHSBBemREvTuo6HFjpYNcZvI0plAcjdUzv
lDlbvtliOPIQQTWqSGw4W7+Mn6ZZxi7cekulp4ODl+kDidBH7QUqHG2K9NHvggaR
5beaCdWy0yvz+7GmvANl0cFxE7Jn8qpQE8HZ1GXwGNDTIM9Ey5eIjjXwj+RLjqT9
GMcISg+Fo69tcPGwqrja1c0IAkmgFSC9BPRj9S2cqB6Z1fxh4EODY5lq40QzWnkV
qXuRm+TYH3WWYfc1re5k7wnMP5Kk1Qti75fakm10YJIM2w842ThvPyKt16lkUGZ0
rdKCCZFPAFaMWldNzLRgykJURBobwammCg8StGcQxtjeDkwS/SxVMo+R+47Oz463
ebJXnNEDZ1isEyJfOU84vkL8XO8XbX3KEB3ap97SiBAWjwjPeThdrU/W4q08Tk/V
Ojiq9mU+AJpC50bD0mObztB85BB9kjZG7SZAT21Yc4Ah9SWo/KuapBIRMjhwWegh
R2DA3UgS4H1eoIe8L8kSuAXThVBkjBh8DqtfR4jJ4+gPPhGL4zWUp7zpP42KEy6P
H/o0KIiqw7Q0HF20TpqCpTG9QJYQyb+Xx9fS5nvIxmStbd3369J/X4Y32R+ZIXF2
Ol3I1BjKPtj+410AwU+PjGmFY0CIlpUJgCB0TeomdXvBrdkni39h6e+r8CLOI/LS
m7sFjGXYy5Us0wM5i2Eov2P3rLHqgZ2RXcsgRsYi7h2DKEGBc7g5aw+eRq0693yF
s3yodMUyFfUlMdc9zx4kvLYfNZPuT2rb8Xeo73mQEJpxtSWE4X7chVlzBAwObHx1
kqrkfHe3HdCgirnYzWej9zSuSp6E3M7xzL/NsNJSS6mQOlRLfecj9Bz/wk2rfDpO
xfkDlt6F0zF4NpP3Zlb4FfvvoNpxMmk+A99WDHeSj7yUiUnsxLph0ZtzautbhEE6
EaVd2UseSKXAxzrsaVdwsk+auvqSMipam2PbwdxV98xUyDJpbhLLFnBN3c+/CCDq
9WgGPI6Qf4p9x1pCtsewbeMJgQKzT5I+68sUjvLE1QhfakRK3Voc9HCLz5X47bKR
BrWZU5BZeyq2uVK7qG0JxyNDLsLsNjPBJAJt3n8PYqoBnU8MuArCiPDSxLs2fgA9
TkPr9bBIBnScZiGACgkRXvJwekwP7CldhS5soq0y0u6yOSKokJLxyJdxPqb8W2+l
Ev1pRP2zmqvzwh5fCXQSqWlS6myaSimOCv3iaAWXQ36lYoMF7E9SJVhEvjO55HVJ
NiC4wqTluWuavYOKEcE3rHISUNYe4vV200JIqOpXublu0I251fmc/F4VZuOOrbYe
ronpoK86EXeGqdlLj0+Q6ZBaNXFJtrOr0RtYglBgkUIcjCyELB8q0knxgpqh/eKh
K3gSMEAn9AjpGxusyceQiXoRSvxy2o82t2/KZx2pcTywAS/Rw/iMOOlsDHZ6YPkv
LcHayLyBzMjzb/d6MRAQdV0kwXWRMTMAJDqQfn75pnpko7BzLJeO/GidUIkhJiHl
gOCFP02lPSHCqbzC8nUnVk5jUEztDfGCJSXXBGaVJg0J/IEbPEq2BFsDGWrFcxgi
FYQ9bevOTLnfpxFrUsTAev2gMhdZ5LYUqS2Hc1WZ+S1U2An/UMGVwollyynE0x5y
/pBLa8xC4ar9vBRyvShp7kqQRmnCDcCHY6+b2cb04WFKGJiSmsDyAHIQeeJ/nflv
sq0AfV9PRrxxlKaq5WYiMbrkp8t8kqzRXqIdvESvxNj6FF7iagPyZFiyYWNxzZWa
VBfDRzbl4lAUWLUjHMKLKkagGwKqjEDtkOmIxmuC8xznJD0XHd9V9+TdlPghy9Vg
6+bZ21o8bbfT6jZneawTTiWGWQoO1gB9mUF4gWbBl1kPkzffVKsF4GsxE8aX02O+
RJnUhRb4ztMupMCpWHnCaRs69SZy9q3oyNoBReGyNf05IOyJcruO1STsAsycNzYn
rdj0VmrSY7Njghp+FYsvP+Te0o2cRZPE+iHdu5KgiDELLH1qlbEE6Rh4T0dGlH8l
3ahanXW/av0kLJI34EoEhu0ZmV2RWL1G1mXyD44K3APb2tt47tDlbTjH7IdWcyKo
On7m9YZ6YtNQ2xwjQiaQ9AIh3xoZMkOtdZl3zKahZ6btvdJJLCPSXmnWbi+26UUQ
pDMUVsDwD5mO9JtcqUnhfOU3ArtSnI4DEkUZIZEf9jNHyN4CKXyOVMkqG15hSKyE
gdPSftEEvzl+zX65zBaRiWoL8pze8HZjmp3LzxrQVWfmeXREwbrGEmNVMlPq3DbZ
l9JwFmC+vZqAh8xhx7oLKpA+nuWjnSKQ5SoUXJpbEJRBE71VyhDkHgWPICcslBc/
ASkXTToxypQEV4Hsclw60JALleA5lDfjyfXcKG33WoTx9yv1RZMxjNpyGm3lJzCc
Gzp0S0kh8APrL1W0SIuCxuOidNb4mfvHe2T1NcPp22XuvErM0JFe2xWkjaM+bPsX
cm1SzC7zO38WZFsSG28tMXsKjeQ2k4zB981PeoqdOeR1Lkb05oDwzxyZtOcjVdxk
z4LVvAR/KCSxZDvwNL2pTTlr7o1R9588aqjerj8HEuKPg1mZc7hmB0cEe1nptgPK
4NeBptCcg6M6hBcY6gWrwnuo+Ydv/I/BfEguPcfiOYkvHi6vULhaud5sf+TeyTyE
bd2aRtQ0IkD2mPQzDVc3fb4xOXczm2Kgszju/kuGCMwkdKVtKijdL4uR6/BLLqJF
ePRX0Iy+wcwxS4G7oJ9zW27SZwok8OBIoNelax0Mj3aSCXT0vEgJ/vwoEhMD3ufV
3C7Dhcrb+GHa3aIE0A9AMcPYVQMffKvIn11xH+welEU7Z53KDgenawh8TzNwK/oq
eGS2ZamOzUQk1WJHJ0cJYeId45hI8olqPpXJ0y9fPxg7fOuf0KaNxwluxEFE/sIy
rmhw0KTwhYDK4mcZcfUlbqxf14bFR6cqLeThLkWBKI0s0ZW7H2nUfFN/d9vKE5+j
lral1fPM8uk4tc0dLcKF7gV0ShA5R1pskNR/HpRn0CzL6IJZu1YJJcuE+Tq1Uryg
NHt+ibA3bSCvrOTU21s6Ihp3deqxSXWc29Vp0Gu/nepNmfY0wrKSAsfnGnF5mjLr
GqKn4Gb2qqhb7FhGNqrdO/2oYrwyzEw4w0aL8BqUTr1D2coOVoU4dLbUQLR8W3Tb
7eTZ+2ku7jiQMtMggKxuPzLQ2OI0ceDnJKYUZkFNp0xJ3uKFOIoM529d6925vY3M
Sek6xk1ZD/i08n8AwfZZ5VUjs9nFnQmaNn7YLkINjP4llqx4YCeqBNEXoCY4lKX2
QL1zNf2TOHBlzYrbRZlO87USqMM7WQnYEbave3BpMsmQRO4ujAchI5H6SpdoPEZp
CPNRp4TNb9t+bxjlJ7GhIUljnGb2IcoOgIPuZgdCcXBp7H1dV+WyKmywGvq/elZ9
OoSBk47pGF4G+ZHiN+9gUrMPBnb+UIAfamUt8RighrsRb8ZYluhGOIJi2/WYLrGX
Z4DnGpq1ZdGyPhgSFGFXfHalvtSxFlTMUD64BRo+Ha/Gj1Juxcg9ZJk2U9+22py6
Fk/dsQuH4247FgKCAaqYVV5ovObEv9KLIJ5BHDmT8/yPl2Ym3rz+tKV//4gRIHwt
Jd25DfwZ3Bw7tv+C4tWWjZCUl08z1JJzxJzdcm2AC0hn0ene0iBt4C4eoF0Uw2UE
vUj3iTc/Uz/5pDDIt/Xt1kxU0aLp46hHQAAoiCyH8mPjWMAVgWwF+Oad1zVaBO+0
k925NloFkdtT9BbgQfr1a/rGLDnm5pVorcsYK623xEbhORTxsdK3aFyd+52qsRT6
YdrIZMiR2ookRKNUUu4bCn/oDq69CH7+HQnN0TyHx+7EphajuwBbh5kpC4WzWcIY
Pz3hjMrCCcXO+qFjajk81uA+u62qbxBrnXsC4hkeQY9ylf0Kf8OZKwTASxE35lFE
4MgQMRwMGE642mQHQ75OQRmzfQuytB6uOHwZIOQGwWHTgWNQFEkcB+RIVEfsaCkI
Yved+vdxDyyNt9DON9rPhxXT+grNNkCS8OQ0Xn0+Jp1mv3VBl29hLc7dTgX/A2Tt
qT+hHHxmk+5MXejuuWWF3auwAfEYACEKTcqU/MY+udGC7B7NVbxW+6dL526ox855
41No9V9Tf8lm11Ke74vUKhSAy2P+fnz9ekDnCxMi73Frk3mafzqVjYJRbSpozD3z
mY0PRhun52ZCipnT2aj2LONHxZuJqjsg3ugqWTWjdZp0xgifIMSCDX64b047Vd1M
Qm46y6XT75RuaJ9ua6FnU6lf7Bm1de+0tQvGwHWjF+Qp+qzaXY5BUXHdWli6iJbt
MxxRN95nctfnfIo3v6nZiC9NuVt4mwve/KZcbvSwT5v3ELuVVEogfes6UESmYAcl
ugAX4Cyk2M3QQEbMsBqJtfiEn1PxLACl3tRP99o4fSY1IOmvLaroKgxeQFV5+oSg
J0YxpOye9IeMeyVca4lvkVaflGS2fi6G5NVZ+pyI6CL1HW+2L/2MX3VHmKvmrBbD
lyhmFogB1crhdN1ZAvQAb9ANaZPSlshWx4xc0+QiAEnOLy7TN7pcv/qCS7Rj2HOJ
vDtgh1W8ecvOyglWk5Os5xt2RE11KpZe6CfdJgSAWhF6+1vLHFF7rYmiowoDSdRQ
YNJ2sQL53j4NZOqEU5DgHMX3+7RmScN8KpGhRH5EVGsiHaofwgvJbDwKL0SYd2jJ
akgNEyBNpqggUJ0w/S6XMUreh102UshEbVXk3qkiAXjDuUTgehcXxgs/mR0YbNn6
xE9ieAxgqm6t3TGiWF7JyMEP5pDvMpLUf2aLn4J+3gEDmGWAxZZ/h2sn2FLEbLp2
AYciOHQXdBTQrtqaF2ESgeAGAbPrevuyYCIJUDg6bXsrB3hhZmSYi8CodntmJpnP
PgKHHGIxH26Q9uig73adLHMhzS78i95385abwUZgm0J26B9Azu6r7lSlkq5+I8c3
I1u5wS712QQMvliA/tK1GTMHVRKuguWfDUHfwWFYEwk6ZJhJv/g4XuaGRoslKzCc
mcF1n1+7aiX63wP51Kh7ubmae/1TyN2zdwMITAqUMKtAVUXLlVbpZ92v1dA1c3v+
GN39Hsgak7gpF8NI/vq1TjxZXAo8pzgr7TNhjHnAzFp+JxB0Q+IL70bE3B7PGk9w
3LcaN9SNQpPTjkVxO3Z45KPRWMIGUAkc48WG/kUE3/nvOwCKOZ2lwuOEOfrkBZi3
KkHXVhG2VWS+y9oJ042QFiAjA6BXHnJyLjjmeM1reTIQgJz/mH1LYBm/k/R5J6WH
Kilfx1EAQfgf8qzSTVQ00fi5Zsqp1iazYdxaD1Ekbo/oHSGsyp96Stu/uXwqYr1m
liNV5TgouTxuC/SALY/V8Wpj1NJPD9DvRoK/uxIsju3U/Bc31vcjxi+HI+fnWUjT
LyeDQV/f5EdHjS4UsJgJvuylv1Bzm5t8WSselYHLwfue8alwiWlLz4izh1CJhF0O
b+Qa6IbH8Js/N+RCcQVPCZcB1nV0PyaHKZlpAw4k53mcOsFcc6UFxZzra5952Qqx
BSuo4Rzp6DgvJIhFYC7lYrQCWB3U/ndoczz0t+/9XHEp5/81NMy35cUzc9iNZ6wR
B5EEr1A7Z3OyiaIaNAKA/MtWo0hnSIgBur1ykDB1jBlOCKXvospRn+abRnZcrdas
w9RWfhdefT1FmLLUcYFkCk90hzA3uTFuPoNS55A2UWvQFMN5r0p9q7sZxzQQIkdd
1tUlEO3uzEoVGSWwKxZKQdm8uDx3ILpknFlt20f7ZppURTeqiT5GuYtlCDkxAera
VFclEt8TwyU6h0aiWz3l4hemUsRnFUfMl4b5Z3SAgswANragcjd5+T4RgepOtEdS
SmYk0Bk8tvqHKEkBhobv35aUFIutEEjkKBT6qXa7u9+BFf4wO3PX3vKdeK4ZCADs
bOaODgDw6khJQotQ4EiiQ+2ObZDyHz2g1k24CzNspujfx8D7fnqjxltTlRbiLtgv
w/VzbzKiCHlMyG8I46M97vcOo2dV29FjzAWrIkPCLN/Z/A97mkHLbMM1zrpxPMmx
zeCGLc7RdfcL4kEAaQSTh88WftoHeJmOiAP3hdsm66EbiPLCX/dZb+RBxDDL4G7E
DHD0/eDHq7gBYzR4XW0I4Ht6ZylbctNLt+fAwVcuUO3h2AKo71H6daoslaaxoq/5
Ut0l6D1Ct4We+e1vl+oHKm1EwkRp1Ey1Ofdp/mTE6CmhVVKLheStDUuwRrwxtej4
E9fCSHQhtqm4VtCrMnNsvakwUZ14DvppUmdL7tBxkGVK2rIgAS+CpmSuXouRVJhw
c7RZIdVNesUdTjKQsTB9tKpurBdI0/KBHA5RgZY11hKijKbrffUZwUAL1AFYvnrf
CMzCqm9QbH9piHjul8/x6b8V4ZIZdYotGGLh2TEsYZkv3h67Ukzt1tQGoxCuVck6
iCKibRQuOMKgps9M/zsI+hhJnVRok1yyxNxjL0cUJuNqAlxKFTokdET08johGVP9
3fVj9BdlUMKkJYVb2hhquhv7h/JqD3yiD0ZSMl5Pg40SDqEEOcy7CtbIIAwTX4mT
Cz7caemuGsEdEU+SfKdCtGSw2b2yxx8QXbmNl9qurf4r/LCUC+PTiObjrpPEm07+
ADEmzz8ROZrQheFcN20i6w2Uu/s4I+LrWp1B4KUM0uSdXsRaEj6A4eUpnhwKmX+9
P1Idt5JiFMN191zLLY/DjKxp/vx8Et1jPEWXIhkvNu+5/n3epIPgChtA1v+i1i7q
7tugSclqZW6UX3dz4xveEwZd3moW2k9fJN/TPfwnwpt+g1H8L2Hqg1/C2Wr8Uuqf
lSwUhUJZiE9yk2+mIhkt3Q1qta6+QZjbk7NhV0RbKx/5sgkFkpMl2+XMJq/2lQIR
HElzFHVaz9zjd64BmGzhkTX5dR6l+4gqXMsV8zQ6sdkvLxolX/ClDzbWcDtWG+Rp
s41U4BHm0xk+9vfwz9ItlNuYXgOl9qRAwSfH+BpxNVUmye9p5AUH+TXkuUJ9pIY5
SZQY1o0yOz9f0aRl5zAVzw7F92uACVAf73trgF+F14KQpoF3HKJFXvAWLWx5OyCH
p49pEXq+0K6VJkASulfD1JtWDVlPhwX33O1FvQ9vkRn0HbqprWkJZ9sgR65dAoPr
z2VuXVLE1cBMKldCNP7vHcRKwuNTohOB+cDl6yTK3fLXCcyW1VzEwpblYAirWKkP
/aRl4E9qOM0WqBFCpwv6/Kkec7qf/OA9W16BcKD5DXFkb2TTQ+yjy1CH7kewu9mr
/jL0OvlJSuQlRV8SqBjlaboDiVtznNn8Wy3+YgJfzcK0wUGIgFQl5NP1CZq/68N0
32NMHHJtI7Fn2lxUgzzs1oW0pGYIXlWTykI/ZiK7Q1fTqjpohTiwuKC1z62G3n4V
J/SBhxH0M+gl+SC0SjW0KfgpxdRm4LaQz7e1qZkpYjW/oJ0L5/tOX/PdL6ni2emP
UAaGb44P1XcCisS2ZFnTcOoF8W0vXGU17aeOgHc3mC6UD861z5VyWsBGMyosR40E
Rlh1h3spkXv51IKmsrvCoy+vXhU5fbQZDNcEUPCQpSemhAIcuBwn3sQzeZAjD8Yk
156O8tovh+91JMcLCSKPgQlp/gH4uihGJjS+SlXdTAhZaSLhLjq6gJy47n6seEuP
x0OSwfWHs/ZKGwfBCoZ0dEXpIzmi9lMRXlOK56X0zh5vt8qN0F39YU4qJdKskYQQ
Xq9DmX9A0acPYnK7fZrJQZ5cjR7e1YlJLUoL37/toPFUJLcRvUBiTM8O5Nm/c9wy
pNq4SGso5gZl3bGc7bkS3CdFSwhMtetD6xxlOkt4f3Q/FCJXETdXk46GpxrndRim
PN3OYM6BSxqsAztK53vhFqzaxO5m4jJD99TAqrJ1SQZtwSB/3OpuTj/6/evc2MsR
3J2qSbITJjTCGVNhDK/DHf3IbMgUdCz8+FDSp/VK8hI2kJuN8E/YMXTuoJjvbT3B
yJ2JSo+dd3VZKy6KuzRRnYudXPWifGALk27bdLsYx848JE/98AS22EtA7wXpRgqg
imzfjiACFOWrEPLxI+AKV3FJf0aSzCs0A6aQVpHk7nVD0kqgxljDkrHy56jD+25t
KiC9VI/x7X5cxmKkRmx16SfNLwa6BrZBBYcb3M3HaO4gKylQppkPW+387JI8vmXT
vqfAbZ4YZF+Merjga+ibo0muRg6jPLljT3AVjIkqO3C4xTHvz/+1heFstB8IV7i3
rrmnFimmJElYdVH+Qtwv7Sn1B+tGQOzCiEFIRz0fo3IXCwS7XEr5fcYaFLacHRsP
mgbOX3XXq5LlbSjVGXUGnMlx6cwNt0D43UGw3H702xZXx9QqIpLaj9r4/OMEp7Vh
gVq+IRXxMaR4z96KR0IzbfdaKEOQBDZoxAxt9sh79D9YpwdD2iKh0sE3cwM7zppP
11GLDOXUzkUF5OZV1OyUy8+duVZ7/OW0dJSTmuDtYIdK1OVcibwVXlRZ4BawSlUm
fSHnbaphTPZPRGYtb4qwOWGX5cTNL1fy7aNjFPPMnXPoiEaPIPgtZ7yNlz9xtsS4
aTQSzUEqrIn21KpFouHBeG3NzW5GTnfJ8cYZQUd0iWrRlwcc4mcgQt8VdwTdIGph
CTro5uh8bvOwPSKi1LiyglDpg+NwrKwYM0bzJWts/WK6GeyJq5VxmXkke6Ln7Z/w
m1NGAH5vK1AW3YhzHUzIXy9Vwbrq8GWzn0/gs/9P7+njqZDf8kBqYUeXVkzV3Cny
QSGJby9vPRVYHTxyx5t5EY8MSa6RNJxc0GR5/S2HVmygLygNdPSJe+Jniy/FR2x9
TzS2WPtEA0Z00uSG7/UTzw5Nss9YPJqkkJebhiPMdq7TJgsWiFGp1uOrygA2n5cw
XolwI5+qu1Xmmy/58PitIzuunehi5sYRtXciatokFG6iTn+OtvdH0nONkfHbyv0y
Aj8Kk2PPshxxhQ+wvp+IdVgZEjtVm+U6vhpxghul/pYZoOxBAok/rCNIt77uQLPj
hDJlCDix8nXERqdMD+VITs9Yge4wwBiqCx2HnDqw9jW+ZRwizS7wM/1Bjs/yMC10
YwmOGXZ/mbOi6FqwqxBfRJmi6Yi1fXkap8aeF2FBjMZA9TCdviGqZ/c6CifrZuF9
6FxP5NEYJQCYCPN98JHdQrFz0iBlu06k3/ygvWKdd9hS1gHwp/Ds5XMnvoFXONO/
Sg3AuhVVGlPwVZ6ShDBOiFKnM7coX66fIs7wmkaUS9+W1f82a6YGwbFelui8b7B2
fD89dvenQTHAsHn/Xnh1rygSGq1C97Z/L9xORXZgSNiNdusggjsj2FkrjFlgwJN8
wLphuGTOZOjKmP0NaaZFYOtWYsQIpbwpeXo8NWsVsw6nS9tROt83Gvp9bxhOsYFh
MBSGYR+h20jVMYOD+F86bKxYK9iID/lILIDlu/maNIi+kjOzj3pwfqHhMHPKaKuQ
rukSi0Rnv4YDDdjbUmMAb25v8JdqN/ORMTCuEXkPOZh0LyQT0iJL3USCjb/BpwVZ
OPCTVMzfkP6yOYa2ag1q9QJP6H/mk+eDlfXH5PjGZmURH/YEfIBoa6J4Kkv4+zE3
Xd0DhhnbKks67nHBN+6bCYSH2xrYZuk76Hp13leZWmjI3Zo9b+tBBOeU1XHoQ7pc
SjZJPqhD98yARJxqIt4gieppzUzPUYo/BbDs8Gl6PnGWgsDenrkekqGpHN1AwB0N
UfzU/HZvKm87qa/zfgkJ7dLafxQZmFZh6pFnZUQphxiFUxoY1tx/YAWOPBTEBREA
fsaHuulNZqlNrUWfBPhRKTVlKVjfVpC8sxlCU5eJI9gylhdIR1xk1ELe6lnNQ3ve
r7z/0K1MGHkXoeg6uUklv9iAq9Ha3XnGi5q9xjGnXNvCMCN4YzqyIhijFzqs+5Gj
E9aV0HBpB/7LxRHjLO1g8mTyCU53lmzgLjr3BxSAhhVbcuEhtKKK7Iew+RFldEhv
iGinn1YUgWrIq6i6KhHb3n3+G3qsBoKCMiZyFkweA6boBZMuh5DA1hXK82ARY7W6
evK9TadXCJM1TFXPAHbnW+1+RF1Txm02Jxf0WbtX+ChSpORV+7xVW8mKiTSehGG8
vV7h6l6Qbo10ygn5jT1kzg6TZonIVzfGYDpHzrMe80r0/pYUkqocQMgrY8u5mKo2
/Dqi2GDxClLuYdAKIKS7/wDVw+4mjctUiVkt/bj7vDdzvr/NC3KaBfm3BPDcQs3w
g0oTaSlB5Htn0Hr7WBFEQk9Bgtt4CzUubf8/2whI16HTtv0KZrbW6zRIejg1oaPy
QMVmrGJb07D62BwsD1VOZ9GPiwECXdoDui4h1KPmQnV7AnssKBdkvHeB0Qgs+OzC
K2njwYvy+UfsvodeR9e2YSOcPwx7fjnqz6aaWZQRGj/YHOBOJpLpq7YIyJ+N6g7k
lCDmWCaubnysFavdRDMv7ar99iCTSZW+zpUJ2lRXf5IJRnN/a39FxaQYGrV7Ykda
YCgbjQ24rD23djKw4FTU5y8qhl7pHvxC/4PExCw1RMcvrSz1jIK7dJVuo77iFwtf
GXZH5BPtQu1FtyIb7DvLS0p+5Gs6ym5dipjBRZL+HDO5e5dvNzIqE5ZjcUHuZf38
hCdP2WyAwsumWpyJVCDu0X2ybeELXPtl6i+jdFSniqbrhoErpGPbuD6ZVmk23Fp1
ym+fmb5ggtHJTAYveiviGzL8ZREDsNqMbO6oACkZPgeL8i5IQVPXj5RrOnQ+luE0
k4MzR8569bTT6it+KlePnvgv2TEIPyb4X7/i4sl7mISEA1N6ZU74y24DrY4KDHX+
4p6X46lGxetL+s9eOh6x5Xco89lWE/mv/v5A/eSVHCzlUj6khhbe7OLzF4l8fhHX
H2ykLIsI+mCLuENcu0ihPyEMJga+YbU2m0VZNXm+bw/w8ZFgQwCdFQoaPrMazd6E
bGUlYh2p3KjuSP9bCaVkoe+4ffKPScFDIXox165rRHoWryY7VEFkF2BJPiNkHrgE
E9qzLnITH6PZvatc+Q8oGXIxnBEHuidoQtA146E7rfyKBPDCts55FUMM4BFJOcAx
hQV3QirOM7Nu7lvJr3Qg/7Wl2ITEkatPb6DV0+XsbMvfAmf454kkqj4eQvSz9o/b
uSDbVuH5csgvV6FR0onfjqrlaRMU21+NNMFeoOVaZLElvNNcpIbJjcrxF72P2Ma7
4RtnLcGeOn4+n/ciMN8YUQRP/TG+Ug26DVXjxs7HGiCeIiE1STV1DHNDuTTztXGJ
e16VX1L9aJj2IsjEOM2rylG3uTL1ErFi6K9w+GB4j302e08fZf+tmO4avRTYqsrh
9vai6RznCG1zdJVVWVKviKajMZto0PeoNaiTBRbmslF7lNhsvzlLMsin/MI0+3sz
Ob/0ZmENGdCil1MONO5glsbG2XhvNWH9uYBFyjL3+ASEFmL4dV+yID6KwAOw+JqP
BxMqS/GlWDK0fopMsVTVKSj1/6ndG4ZYZS1NF7OhWpPZZiYzh4WluOjvk1cczJdd
aro8Oyj9Z1V+J95xjnL03ugJc8NiVy2Vao+dkt6WBCMuiBIwhLzPwEuQxIFKcGbt
xccTv8mKBL6WIZW8hbESgyvDkkHZoIOnRzqazuR+c8H6EIBo7QqYZ0pR5dqVCfXe
zKim+fBOELw2HihYXYVQ9sP6YBtfecAWBaV517VekJnK6VUHeewSEEz+6Whrjb0G
zRy0eQUhgWzeFjkOp9uMovXxgPQtuct+3ZWgyfjiuWHMS/iyesYIyuOWJTZoPzox
ytxeXvY7ocMkgfXxkiuokLTXizioV3nfbcWlvTAMSOS2WbhuPSY9FSyAPyWVn35S
v86+2u141woh9E027Cm5aEgFD1wB7C6UuX/sskYyjrmSw4w5WsEbx7G1gbDG96nn
BEBhz2DhVl39CNbkblEu09njm2u9uVueZO9C8pap8u0x2KQY0bXkbUsgb6cD+r6Y
aOckXHFsNrJ4xgzbj+1B5FgHB3ruG6IZiGj9n8WN1W3/SnekGPQBi8RM61jvwkCU
BirDof+V9b2P7aWJ/iqMM1N4VdDWCgtE5ShjJxL5sZaJzOK37fawSpHv2N4beH0F
wB6aulK6WpAbzjcbLcgZe6N+Aa9IzWHvGxPjXjMIGk/Q6W1ZZKYWYhCePqCNzTI/
DRREroI/Voqjyvxr5M+mDqTmAw2/X3iUDj7BwYjhnqzW5C4DRQ349OSQ1+Tv0vqP
3YigRMcKXiKbrKvhJkjDZhGKt9mUky2OW+/6WSYmM1isbaglhUZMS66uQ9cKr/li
cHwbL/ylAmO4Zh0TXgNZL83O9JePhm+cENzA0/Mk23Mx81DG3HB9ykofDpnysZD0
QaI3U20dQnTQy0fQmLnM6nHdHyDKbD09+lqp3MJUkaUoiyCrZca1vOkaZ6ijVYiY
ZQHclVzdl2VSrwLcurmTTF7HiAwPbHCkgkHs0Qozc8p6eCGbOdvvMRzIw++Wbuts
b6MpxBAsPPJEUDUsQ43gLHO3wytYD6/gGWztlhnd+aNxR0OntoD66Zx2ZBBAhfLp
DR6egUk8//z4/pV968OiTah/J0Ph0u8/CTqIlCoRMcyiHmzql9FcwhNHIStW5x10
gKKnncDns3my/dvmOgv95yE312c9SUqOFmIWfv/eKDJDsF2NZOE+EbGXxhQtjopR
ZA2a+srSyubcVG+Xe+c95ak3s3En2adj1QlfDeseKvAUrqRqdIrx3eGzquZxzMKf
02eNxJ/kG6ZcaA5iYtQGGOJ2JNDZm/LWTReIKXFSw2IlhSSwyoSax31X0tqqsMGz
R9wJH3574BjI5+9CWzxSKGsopHFMHPrW9lqtEEjssoD5dEDPBv3VMfn+yKWLTnL4
xh2KBc3p1EL2w9tr7wOPsbiab46AvTiiPHut0fabvWiaoWoSD/BdrHvYPIL6l/18
+R+JK0gaAZetm1qOSRkRCRx4NAoUPhbJqnuxW90UDaHKf6z6mrI66SgMgjQPnkPL
d2Mq2paFoGDkNwiulkhPlspbNDysrbwOV/pbg1uwN7yuZ5hJhfw/sbmTu3ECug04
IRRrhhIcrZUcPWzyzlrGGxL6cWncu9DsE886Q8uPbBYa3q6twag8RAAjfqWL6gK9
mBRDDXO+DGwz8GgJpmuc3FG+5EkIeVd5y1F+Sq17ddsyJrDeeH+EuJFjIaBljTnO
6Au5GYE5S3dJXhs5oHUJb24Oia4iSOGSJIxUIi9ab/Ep6czSF8SnlFUyQNnZsqjI
lfUd8BhDgOEXDYONN17NcfINT8dbssIDIhokkl7e9XfaCz0U+D44CBF4HtkwcKQ/
4CfRwMgeHz1eTNxMlvH8Pts6kkCNdQELKY9eZ02A6sKgixiAKH/CAcUUUGStVu//
tez9JgFo1W55IX3OxT/ebLlzEmIwFGv6h3TGJuG+BnDOmoxwhcIbEUXZq2EITIuU
0kZ6j800UMYRdsn5Yij4QNBtmMSKE11uMxbLKw6fvNApzlckWKLu5XJ5ZAA6gUOs
HKvgiashY2ckFlBeGRJxxd1Eh1TO5N+xY/UK1zedss01UiauENCi+NJoAKFF+hj9
A6EpNO6Xq+q+fB0MV/SuOT07kKKYlD7JhQhyn3OHKMLgDtoRc+mtrfmTAPZSCuHE
CoAzjcBNdcHjkr/AjwAX/Rauuw1iNVdabtdKOMwTpP1P/glYLFFFExyv0qsWqwLo
4Wl3Vyx6gKTbhtsKpzQ0krFUuiUMxPsxoG30GR/VaZi848bsMvXC69aGvWv+3rtg
KEhE5kI10MJQtsACDTWp7IiFqhfPIOQd5yW6aYJznX5ODg+fSlyo+WCGvXz7XWmC
JjNbV+2lA1n5obffWrJWLKlUyceeZ9Kt37QaJiNrze6imLoVWt8tVONS2jzEqzZC
9wRLA+njjNHti58SQgfJYaIs/4NQmIMGAabYGgc7rvumc29bGKfOt2SDl2Kvhp4o
BxPYKi1kRAWcXUGQyzXXaHDeshr6cnE3LO512GXTE4tyoaQ075OtGnK7vBJlomOU
Aw8XK0wQ/RHBYKZNrJbfJXzEhUArhXH6IdZl8SubwraNdm00sKhRAxx8fH55P74x
L2juAPMYUnpQOJCIMTarhV89AIw4NxoIzjKcrox3NI7vezjFScxplPFfku+M5GyZ
Nqc7k/nb1kQFGbq15NtX+4CoMMGHEwEdKNMYWXpIKnSRGER9qRC8dLSc9Y1oIk1/
dhmNadMn97/tzZGMYnwu8L5/VY0zWyyG6+YdQrKPRdV0TGd+mLCgcqCekKbrWGvW
LotwouG9jhCz3FgSUXURpPqLeOA2MuhhDRPbrwlGHFh7dX1kHaEbmtnv6pB0d+Rk
u9F1Iud5GMEpeW5fF2SXv+QYizGM+6Wk+MjdcgBM5Ziqgg9dcdk+tKWyvBVyGfAj
n0o+XuQ0adqaqH1lXm0iYag4lqPmpIQ3djtA33L+9qiWmbYbiM+GEE0nQUfim2MQ
GggxAvtBS9c1pVsCMZ0KBrSLX//jDq+adHehDXng/eeQFqx2NxA9LIxnCsZyE/bB
+IYK7wX5iUhlayTkV4j2F6wCQB1qjK4sQ8qfOjFPc6lg2GBBJInGmRogQqAqDD7u
T8kbl8Iwu683CRBZ/9SkeVIw0hEiiZuRlULFp/Fw0X3kw25N+HyNnKGIClZHFWxd
XfOVH3k/vj7edI85yYLSh8Y4BB69g4OLkubBW6K9O2snZhr3AfZPx0hA5Pq9nHWm
7aZqVvHyCCXirdjePatzvp4oyQiRb5ECIbCW+rxThGM91+OCPoUg4tFKAenkhulH
Rtb5S8q1Q6YQKSNbBWIKR8tmdk4J+5orsgghTRrxhWMz9EJkP2mmTV1BwFsT/jxo
9A0V5ZoPMyZ99lvlQtzyBv20nPr/W+8bf6YrGLLnhnkOE/2+zFvyHKaPAVQheiiD
rw//GvANyEN1pIouGDi8NNHo9c5YGGhTPF9osrPPz9XscR7uyP9zBwdux4OYzkLu
FmqyX6QYsAZwdsII3AZ2X8UxUTb4yQgbpbOK/fWjRpHwX5UaNCjg3y2MCoiYw6JH
gb5uQrYYiglTtFRqr1cIUWaz8D7r3awGMga8+kt4GAjAC/3T47hVtUeOSmJ7ZNLd
qlhecLNPMHf4lEBKC6qu3nri++etB8hpuDGOq3sLFq4mxqUEVblYROxPlAhIQzuA
s8NJuxYgGnsj+/clb/SRAfvIE8cBREv4Rn6BxDWN+gpzOiUhMB59zT1DWdgyNq3D
AT6rzP673zWgiSN+b7XcJx8jlnFroaHR+2WR2HYOtQrs1oyF4rLBYI5ngM01XFyP
mDtnZsHXyLNpL52rfKxGWZF7PKKtAjm+TnWwCuzj+LUx9B0tQ+YroGoWbfDh4wlB
vI819Fg9o6Y0dI08uBaxL34jLV3uuYqHy/P0cv4QhctK915kfb1VNDjez2jA7xWj
oO6YwdJCzahbCAliaX+iBDPoPM191/6ULgTSEoZQ+Eb2NYMuo4unHZQGli3zaj7d
735BAkQ4nQe9ZjFPSsU4Mm+GBtv8EACPg9rpDxQBvSTskAfjz51qPp/t6cAPo9LM
Nu/X1Vxsc+itOVCHN6rcPd74IBMcgUV+bvFfONqwB6TLSZneLuaYA2bGD6IKx0Yi
a8zXM/hzrh2tkuRNnK4RxejFvWyYhQ8kW/+vd88Mwz4Y/hj2aRzwZjPzxWqBxrr4
Ht+817U6Gli/Jc3pluOe2cXlB9b1EM50wrGbb+uQ6imAqhRlW93tzAzN24dqUzIo
C/GbwcCJTYPPKVQcXlPIBZeZ2yT452rIc1s5k7O/gLykPfcz2YS+97bOtGoGL/Rw
ZUXUe1Jy3IANmpUPg5ZP28mr5+o2qJoKzgtRY8cAyD8RXn3SmM8+Q0HVpn3BinFJ
brRH9fHQmo/WPKYelNoqq4hBvCt1Yl0dFyuAjQ+uRmjs6a8Plb0eBbaenqcvm66y
xi2pC4ywxTU55v7qm6c/GIBZoPWzHEmwqPUEOMKpq3mWUYl6pwgktFkaIgsS56tI
zKaWAtCin322Wo3oPPKz11Ys1tZlEy6Pf6aQxiZ3H9FKKIjWSKOm/dw5qEeWvbjW
N+JCIx8Kn9FI2SbIh7hJu2HOVgG0EX+sLWiT8CScr7TBDoMctpGu3LJd8IU1v6D+
gGqf/RJnI0gvexxrA2EnhS3qv0EK0WbRrg1EBIGngvOzGo80belr8/EVEtVqgGo4
shS3NqCwX76nmnycC0ZU7h8XdxE+LyCB/TNMBXtu8nHymimNRSY5rtGDp0Zdn3vV
3A5VyVTH3nk271gTHc/zDGXR7/FTbphNdN0+W1c78oKo5QKX5enM8flyDEm6sH8p
4XRUWKzY8Lg5ME4GBYD3TxtIiXYECBNtTowVE4f3BNXaXCTzCeMbmH5UA5kfJm7K
A0IIz3E1aKySq1CfDnBSL91WIGw99A++U5L6vbUUJRUU5jrB8QgD5LtjjHUsxwmk
yueukCouV2cR3TkV2tOTevSsJpft3Hb80bUwVxDnm3tELEBL4KDS2v82a2XUlpOq
c1geTe1DDX0EseaUwY5EEkBKD610JGO0v3HaAm/3yceGguIu+yDzODy1mITFLH0W
ByXMPoA8eZw9VsfpTqXrhiUAVoFx9lvpA1AycXEBh6CSKlONfjIE3liYQ+JxFcqv
S6Q0OfbWwl5yRrhKdSK1rZYsGcWe6FkNDQjIklLfwvK8f5GJC0bseIKEnQbsvgjH
4O1SBzQS0o3tTEKRg2IkjoKPi+TSHuyHvX+OeXDxZfs9OHT/7XLXRPeviZUVJNTq
Aue9bbC8m6TxjPx2qYSuFUgVSGHJXRi8xecdJmMqN/MnxUVk7xAN+Qqbk3V5J8YF
38R779ZKyML9rg96aOA+zEo9GpQmmpiXNL0MtN9pql1nUPydQaMiNfn841X1P0al
6RRevyYmShhvyKiBtn3FceJt53UxEOdKI6+cpGV8Ki6UE7Yy/FkVTYlLG7Wm5gOe
ujFLoPumrB9fB0ytHh18Dae0Kf4wSq/StrpyiBfQL6GD+u8hH4htUMmRT+A7qpsh
F2ukXN7/2KHKkBP74i32vqGv16h0DYI5Ow8GZ+VVx9yngy8gLt87cM+a0OO3ceR7
75r4ob956y8szCnZa7wCBbXNP0ywR/95nLud/GRIVrUmD+uy3uOT3b4c0tk0R17T
ucpr8BLh9PakNbKmevnse5cOZdr7JxGJL7vTVENyndRPi6XrcraeU1uUHaoFOA/6
Mdli6aKF7LDBuU1vlUuEmsp/2t64O5T8ZJJ2JSoNgjh2+4yxTcdVsR3FYOoSJCKi
JbV3fQSoNnGy7CJDazLuB5qBq8VQ5YBL4NMrl6zf5TBCUQpabmUmr0M8cP+kWFHg
BLVNTjpiIN9jzomNYJEEUEp+YHBg3piPJlwINBOysaziWD9r7HKQw2Hftauu0LRZ
zwS9BbO31snin0l2Sdijrc+ZoHyqaB++8w4ePdVB04p+DxU+XtwcdMH94ZUUNQpv
NyN/uKmPDCSYOnb8KQoWkjQX9ivpiSeMxlZi4jlR8LP2KKPLb6iXuipBpAnn7wNR
k8HX5J81DpwkP9V7gGUCtPwN+hn2W48bs42G+gh/0JTQeqeyqy5oUAejZev/OqDL
IEamR5+QZ4gsODt51eIAJa911tRRHnmVX9gf2XBm/fApMVkRNd3oFC5vHyEbrDvY
QmPIaC2ka5Keis6oGXsD/nokHoDDCEPReEYpgTo/dWU5MCFzuvWPNF6SBanx1Emq
KFzDx/egkZk5btd0WraKhevpsuW6vSxxYVRrCe+XwEwfW3iwQXnaV8CuNRJR7iWm
6RHYhZ5bMJM/K6Sb38MuX+z0wEFBIXtYKjK5U0w2ZBCmGyhN3lW6HIm+kNbzI8uD
zu90gjgImAA91HbIB7T04GARhqy9QQtweOLKE71H8c73I/1RnK0zaMXjVwswXQMu
Adu47I+WwOakfAcswNeeFvIkkrOA+HXDzFZW4+/FrJU2nPou/DjzKa38jrkYPfya
18PpVlfvxaLtKKRKG0L/paTXjtKDGQBOh2hCHaLIslcan1h8pBIH437o5w28ZdTR
TqihuiSEsszetHLeSs6QjM5XnEW3bVd0/nVoy/C7rWkOwXfqE+lM3JkkalS5gmey
F8RVfqgxJx9o6/NZTUxaUrFu0k560yuuRJMII3k1moF6SZhBb8WZ1/G0Kha0Ge1R
x+x7hAcqzfkwbfM1Akarvt3HAhHEOlN8OEi9MwmfyFpJrKv2FxZgk1QVxThv/TAj
zO7BvlNgjEjwmvPQWoFx32LQoWrW1T11Los1kdORH0zkJUQRJKYsh7SYUDUeQs7u
U9ZtGMWWJMUVzdpNaoIPImTpeogJNZXAdregYnQUbxZcq+jM9JyOAZlV4oOekssd
RcO+pqesupUwbCtxEIl0OVApc98QX3URCTxtf3GM+OdzkJX8yur1i4KMrWAuuENW
OlJdKedfDEjGnSrrVuk3BSrlhu29IbvmhxAvSUR3s3JSbdfKU+D5S1hZ42Kci29N
PmeQg8Bk0YPBFAAkEcufSNfMJ71hMETvRgJXHgasmX6Cy4Rqi900SctJ+RY83hkp
nqwzo40EkYtf7It5XonGNGK2ghgtlVbUxzEQdQ8tt0mbvjWwBh5uNaDukaMDBRYG
k/3MWhgfgOWB2O9mlwSghoKfuA/BoyIiHOEouD3czUXyqZpMXLOF2ibQYl23rERS
raqz5s0mOdNlIejlGCvhDi3wi+3Gr7ksrSWFJ0fZTHDJiZo0eXgsKT0lDwHb385x
kYBDe3jVjiR/xF2rFUSlWBkqjcJetCHw6pj1teqkQ4dNhB99vMfOtu0v9StdIDIL
KHd5DVL1u1CI9tsMNqWPc4ObZay/ncAnbtmdx5vW8eNyQ78FH9H2CX7X6fj7Rkgm
q2dIUZNO+P7cIK7TVANkP2ORHizHwvZ+lw1GdRrOgH6s4ShlmZkvmJBA1sFM1tXy
wI+16wCv7qeds9yck8CK5YldlXA1r+hIjoLzwbgM+zkj0ywWHxkVWQbOMdivDbgX
6cwk8Iq46g+TEzcvpxYzN2GYxYiP4zmOe7oMk++TSWS94kXTTBbYYZSy9kev4HAK
Tv/LLX/1ETazD7HbDv+tYMdw1lUs9ItcGTcDuIDEHwFV20Nc9M7Sss31KYKJR+Xk
QK9H+FVBSwtbIiZr/s/4ueRLc+9ibcunJX1/H8iPLBdt4WAj/Kf9imoxxICXD0zI
D5PzDFHvgzbbKTCyZ/Ztfh9zuHxTdbsSmwlNMc3fJFTnL7WHhQE4+MbOvLrxvx5c
MtqX1gVJv2oqUUrk3q6ulATm7GS7iYFDVgMmryUUXOhsKAfOv9xSKktC/xpv22Ta
iHIGmbBQPzl/dk+k3qwt8yjY/qxb1edXEJC+G/qAb7lhq5R8X30dJeIrp3a0ZdQB
luTwGmfXftQEf0fh4eJCCPCNEn17mKbkCgdkXDx4Ewf1Pjc7/Z+/xwxU/2kctEPR
5Abfv5rqwyP3puuwNptnY8EMuqxNB3P7vG5IsnVSd7DyvuWtOS3/hYgC18a1CbFH
Sr+oXZ0awKa06+mdLt9epeabfGUepuopZ5FiAMvdUMdHFQ4WmeEpAHIT7jldkwAB
UxFi8ejHU2bTJW3qLEk4iVARUWbKRqHj+y4xeXdABdWv1/U0U0EvtlJPmiSV+/vD
GmaHuZt31EAbHL6Ur7NvNcl0HeVM6kKSTnJUBJslK1rWFzOp6H/BuIjWFNwkJRGL
lmHD7zjPazvOQHE0ESeYBaWXn1+SUPCibFadKFtCbH+Jjh37aWCVoRT0FaXRJFr0
uI8oYHnpkpd64Hl5RX+l+WFMQsfixrR3HVD1Ccxq62a5KC0+240jtMyjlGAH1XvD
6BTS4FfYkUK5jeUMt+5tgI6eNUaiPaO5U9oTtRw3tT3/uIX3uZtJfqPjy8ppphwU
UmAvcGi3pmb+clODFh3gzzApFiKGbZuSiwHf2C0LdrwgvHg5a7J/OsppWcYZrqtb
m4mwk5Zpow36fXqcPkBn9IQq2NbkUeoFrg2V+AUbHrGsewpOkv2MgExVKcfnX/4n
sAHzyIX3wzpxMa62cj64A1rLUFP8Qau/SlnVDKIt8rxw5bT/jEe6Tfp8NTCaW35X
DckjDWmKuPfbQkCimUF18Hl0lHpW6Z79K1UYz1MH1327RxyWFDyqa++qPNOT/KxE
h4H7T7qGr7X2jblE8S2R4iAaE4Mtc71pwceMWKw5fYF/iRbaiiITtSYgPOqnQHrE
KPnFM3Bzj6mlB3u+ktbQTSiq8RlE6Lln3T1N/8SZjN8otTFIxM7DaVhl8+YubCrk
H1eh4SkjM6JwA24xDqcAo5bGfzRCh7y3SnqPS3/SkyI4DusohStqpBRKpU/2O3UM
b4KzamaTrEBlb7Hca2iWTd7PWCNoTL57+6r6zDXhoUTm3evJzB6W9eoKuq68Dbzq
lymWLdWs5wld+r9Pmm71nJlXXbhAdNa1UUtptPRF0+T+KwvwwSkrUMIh/ToQnR1C
BlYsT+NLZxJ95BBljyK8nI/nBOrdt6DtBRVcr98Drdc8jaxgq99ylBo4B7VL8p2B
ulUDlqdyomxdQg+EahhgJs8Nmi0j3oWeQF8Ls4KhiJgqjSYWpfoyHFwLtlUcI2d9
Qni5RyRn0xijrKZijvC7KNSRjL95iGKiYfBPWIUvxt5h5VtSg8RNXZYMa4dZpDlb
O3Q4QdWsjrYBDiC4kr+pvs0PsThmk9G6VA9s6qOGU+8rV2Rd3C0ATp6sZczimJac
4Zf+9ACkVFqQCM0QyyByFM0ZpbYJRTQAwNQVAtCMt7sHCMM7Vidnd+vKlHNmtFw7
ViOPNVjojpISjEzwYx0reHGvY/UZIPx2hFOIKkRIDZeLV6jJJc+2bFlA18UNkg5W
NyTuy1iyi4fhdlHrtDc8oQd5+JV2QnZCSadBHvY3jmC8hYw/JOEUHFHqjXQsVxCT
645UIWB1sY826HzGvXg3Thf4LYQVBPO23numLW0aHgq2hvmU7T1C5qCNwZ7VQnF2
tP5v/3RuB/VLklIWERO6LU3bsF9VduAiYa6uj7fSJR+9HjzxO7hAyAN45Gzfi3xA
E33K8RKfYUW9NMI9ZjbNsTl7T/MzxQE7dC8KAO7xKoMwuAFF2tPMfEQCAs+lRh0z
7Doq0gWkSYHOQY35POTSDJMifiNOy8IqDrMToRcI0tLSu8MPv6eHUj1bWL/3nBGc
STp/+eoc0kkKwtzBjy100VAIBg/Q7enx54ymUKhpRjNr0fxy7iJUG6TmW+WZBwqL
JUs8aDjQVuYJdA6SP2CKcYy1Tk+vmxGM0gXRUBdng60u7wRG0lyU4tH+XSS7h3O1
F54HGERqqswEXY55HOqu0sb8iW44dnemel8Vaz22kkHg/HKGU4Ko6j+jDgcOpxaA
3IqLpQGUE3zwpaFlZkqYIhQHNvQCWnfkmqg3LMj2I7ESWjKcJrLMbgW0z+YH/Ojr
3v91+0piWOlSlkxGoSug6g0O5Zpo3JsFw3mlo3e0slLukkS2sKSPKb651gE4U2fM
oqOGDivR8JNB84Fxziz6xRrCbPT9JwLK9HxgRJPf4hsPPcnlSf1cScL5T0Zt3c6o
gaVYO+JMN0CD61jrS6TDwzlw5QSTnpq6nFAiGVZWzasx7mNXth7oEIjqUsYpWjra
NVPOrp+cTbyInyniNUJj9P/5/52Ht2wM4ikzEDRWf1RKiyk+kujlM7AsJookDhDv
PMSVyeI4ugMZ3LkHqWhfMdrTheJbFrYw2vzuiF75+01h7oI/xcixwvZ/pJZiz80b
Sx1J2QrY5T0pStEESp9hyVwg7VBoXAaxTAVXpqZWVUKA7NbHlAH+vZteDFZCjDW5
6KNhmbAM2k5kGrJX8DkkWQl+dO/LtCpQ9pqWucQlBb7nMEBPvN77EnVUyaC7txLv
zp28vPGN+AqUnctqkjZ3JT9PUQ7JjAWbFjv9/pqjHn379ZmejrYLYkcj/5xtveJe
YJp0cueWlMVQasWosaH7WcoXFqxKcVfJ/z3lUT0No3E/pYcIKkxqdexhwgvQQCQj
o9CZc8xsNBkcNM0A/IihQwynz6HCRYP8uEs/bTemBuU7Yqfj7g5J3zZoFDX6dfK9
RpQhMI7o+lJBmz/JCtjIeAFUWoqsB2vjPZjmVH0z6Xk3FhXmBWjYk2nDY/7FhCTG
wmHhWo8BLCEc+0KXM2YSzvFXvjmL/8xGU4mzJ6iNp9saFv6byzOYI3HL2Igll5ls
6zXcD0gu+OuMRN5nKjRnJg4XOEZ4Rm/ES+zudkSGkbUThqpEdQfLMR0NAp9ZdvFo
IFY5KosLX5WDJmcDCd0SfWnOEYEXCQL8d296rnpFT+anoB9g+3fowG0beV6JiLIn
TR61osiNoOPYuf3gowQ+LS04qs0yJ+8KK6BXc7fsHNKBtUVlcEa3UroLb6wCNbyl
IPE8G4wlSSr7FQDOWDM1Rz/XFLP4oSQGFjeVNKeg9matZNvBHB1iFFw8SaSFsw/F
gD1KoD0Y9ebC9H7pDvSaJyg8UqeVwweLQzmQ/CRpQ1oDd4ra2Nnuer1meliqvJuB
Xkzpir7LuRlVqoBwvpL7uO2pwja2YO1IpV4n2zL0YTKF188Km3ylHwA3DFgJjAHD
DKZOpEIsuZuvXpM/Zom9K5SjI9soPzlZfSw+JFIs7DB3XQJDaZ4aFKSzblB7e7WI
xsE7LkmC7mNcZsx1hXWs3YfdBLLJFpvymXdl4exBvQiFh333XryPfGXTU4CGM0X9
MU78vz4hzgwHliZnZxNrlx2wBKl2aqTMJpxuroqpDEy+IZ6d3L+0eYVlCy2MNbRu
wdZul4K6zRQ5Tt69/D3yqs4kwv3OjNmkCo75961lbf3CWX2v+vPEokIfrm/vJ5qC
pGyRJdxVXVix+zNDDGbxfscbYwwe+/DzdYMiFMX8xEfikML2V0QrhaTiWkhRX8h3
0uTsdELzCLcQ1IjzhzImVGKpP3qKZGtSi7Jfdjt0mgTPofUYSNGTmF0FPABmdj+3
iatklmiWMRxBtsG3Ej8fUp1S6bNDUFXY0MV5YJYppDqB7tL8z1NE1egZj6zEXXoT
3XCYidGlzQoRaSLSgDmbulUcG28NoPZGox1G7LATtv/gRkiK7InkkF+WIx3hGPpf
IfcYhmnluBRVFAHl+x45jIoA9cJ3O8qDSnnVTZ3TFq0oWZAG4yanlwFTMLWypogv
BSA8vLepqyvnZzqJKzyeX6rqeKKqRmiQPhhjalSLEMSxutQ9cw9SOmt/8FgLCu6O
NogGutaWZH5Hy9eCqtWAtYxFQt7nxqBxOjVnkJwhDU33wIyxfcG1lJZUndlP5E3e
HxgFNRkCdC2NlbUls7hJ+k8EW823RfIN2PRWSd0xNkquk60kFW5DwAmp3Bea8DzL
QZEVpKnNjV9QgNtTlgiuXES8C/NCAHTTzSpiELmff5BX525cvNwHWtsh7wRl+EQk
LrsubAH2z+AG+4pJ8fKWR5gnHQHP5ceALSekh1Dt/9pmdjpmHpXXZoC1+5wyol4W
ULJVWR4INKpSGdu7TsJdBFbSYn+1suGwDqUmzPq21NnyPSCVoXZQ8cCWwoh7Kjyq
gr5XIAYuJ7juojkRTmdO7N9hCiotLz+IlEOm3e1f7rHwWv0jWQugiNR6QBEXBKor
cEIsc1Rs7VTVCBeWZ/Fzz+0ZTIPD3z6s5ymVsf7ixgLtj5ySR2JEsKamht8SEG7L
VULjswwCMoDPWVIinb8y1r343EZRm+UpR6zxyoDn3PF9fzLn1NLCzYWExZ3tlP8Q
buqmV5M63S9E0BBJnuO+h6QG5sAPqw55q/7dq0VAq0kyru/CRO3V3PsPxurqf9jW
Q08LSRxOulCjGL5mMKIntDNQTXHMQ34ERdZ/OHO36LBPOCRSFZYxEvxHMY2nBXbA
cdcKjOWvEN8x2+U07kc+UxGz7tU94IltoLmMATP5WRySurA1Xw2R9nwfw7VYX1kr
1Ad8SZSGxASUBK5BwGY4AQH95SQomYxqMogMQnBBSHrfElbNCRy9QzBVaJ0N7/0v
m8ctA44TItAsybB2myt/MgGALbCl54n7DJYPq4Z/0m0NvgDWlAaD8VkIIp1wSVLY
H8yKW9BRfwA5yRXXinMcqagEoGm11agIMT6kOcDbRcoT4w3wnVjfvrf3ffqbBMgs
UPqaNds9AJI7peByhObwVm6dnoXGLV/nTtQ+dFYpsVQYuWH7Ml+Fx9dtYgR+AWc6
xIM/2mEmHlCwDWW+qauzuFNQsdGq+l2m5GUJyW+GngXYBxR+eVXo13gir76rIog8
k1tGsKbzHhf20hoORmiP8VEBFjSsqmGbdjD6DqzRBktj7LtZHkg12+dynvhvUNJv
RirRzuovOBcLP6boqX8ViVdhf7HsOb+JspyAh2i1cOQQ+KTU+V56N/rKoT8bM5G6
Bln/jFHohl0sDfCScz1gWLy6zY4MKa6BxO3oxuyM8WgpfOvzfjKLu+rnGcA5Lzi5
O1DhrWVY2MOZKLa8r2cevTA3nEFmF1/0hIjAb8u12f1afGPh96oIyfDaNJRB5EqG
YKgSVp7TaOOLjABtpUe+K1bcNFxRxruOKgHwDtjRPTPd2UcX6J6yf0laU58V/8Dl
0JHmdzYFuQMbx0PZUO2+MKdOyuY83XTL8DMSDeECXDKUJY+sTwAqmoP13qmQ5XiZ
Jmx17wz7r1tYsLpDu6nKs+KOV31GG0AL40vGqYeKt021syN/itTvVKM/vA09fvj4
nKxFw5e3OgwGL2ZjxIWjAoxONC4EhyW/5ra59j9NJSUbW65cZKH92Z542Lgi7ijL
sgCywWXChmmjBCq21+IMVa3sxg3Vh7j9v5FYj/8cuMSXZci7lf4hUlT1432NeS9L
dWzrmMkk/7N3VHcouVo1jpMnAZF+zv+BtCu5cs1TBllertscBqmIH2KBszeYbRg4
qaiv+bTwxhLb5AZaAqcLC/JXfa6xMqmJQhW9ADXm+BJ1XdLC7vMnx3VWKRzwjomk
+V6jSztZOB9o8mx7PqUuX8Rua13CaMfABnZ4OCDPQFi+Y65wPc0EBvvBtYyi+Vn2
aw68ztQLBrTBYVkSm3/SBC5FmBSesYYLsHcH4IuqIwlDyhpG5LbawNYFxTS50j/D
qc71eNNu18yI7+1FrutYg9XlUdv2EgD7mrpiXeUVnM33ZTCDEHXxSNHxgQhy28KH
OgmfR48Hv5Ei02Co6U8BRyW2hNZKS+boZDDmwpRaxFyZ/L2HghsoIu4xl68jk0te
tbQCuUe5Sy4SK/2XRzDAC7Kc5QHO4c6gNRKcLcvI3lqhdAD2x5Cne43w7JJuzwbj
pjDNcbbjI2iW74x5PllKYUuDNXb7918OmQ01U2h0ve3XI/JS62qHzsWn0cE/JKeQ
9KhEROKj0Rl0qP/toRV42disqyS5zRsymiXsW5N9Tx2MM3qKzhvxCJvNDdoO/lT1
RinK5lXQ06HNOEKobeqTTYlvY9be9ms6tvSFNwN5WX/7WNL5ro/3yeKb7LcUenvN
40KwmXKQmTA4Fsmgq0bbMb/YRx2DDJhquLTdMd+B4EJb7mTVeekqnNDrc7JJs/+w
0yg7oHC+2dXXSyAJHKHsqiPTiGjokvek/6/oJrgpDNxqG8DK4hJntXeFaeTNK9oW
7+G9k2yxl74sEKGPuc80A2J69bAFVzKDOAOJ5bU0hQwCFUueowkSgx/9rrvAaP4h
itVmtwedlcw+B0NODV8A0LHXJLqFICVFudOrtl+hprZPP85t1YmQJSRop5LD5J5S
YGj2q7p7/bOw3L5XLQZe/G33YDN8sBbu5IWQ/OWLijRJh1UyYUqs/LGQHM5abV+O
GXk38N78kMcEcqzWMYfPoEw20sopslR2Eg3lWzSorWNlKwsLgrJtylD6+zghgXzM
xrXEEvuJwYK2OWxmcCuGiLdUlP9uRfgJKLZX9spFXnGwMLGvup/Ay26Gzq9SPnIa
zkSVy1oTk0s2yWWRF5K2H0jfu5ODBJkJwFvz2ewoXRt6m6EJDyL6h8rlaQTfgePI
wBPEFfmjBwu0I6Pw9gXIFERdbLXsQdEedHXEkc0eY4zcsBPizLvP9Jl+dYoY+b9/
cWlvjBC+k8/ozXMVKYE3gzd2uQktH/C4E/oQF2Awh+Zh5BzypvPByCwvcivj09I/
ij1bxGtVzdmsFnUHQVNPnj/9MtYDhuiu9iBd0RWF2hzfTULzWOq07l38fnBgqml6
9cJV8u/pkZJgsc8XUU+uY8zGV/KO8mq+swFEvIJkFY0Z+/yMwpntuSmgl+oeqdDB
f1yM+7TQGIbdaPFYW83WRcnzvdTnQKj0McziKgJBgY2qEuE75oXJU+k44qD6RdSY
5sVX7aGZqOAq101fsEP2rv2eMxWLI2c7K2j5FJoM/JMtKCG6kC5Kwi/zcEuA56bL
DazSLb+LgygHqAUKeo3NW6oi9Ccl/G6Jp6g5X6fwj4foZpStrp5cDbqs37mWtCGr
fRfzMqrzEeMtoeo+VkTun7G3v6pIB+SWZjIhPOftza1Gx8pT2DrxRQ9hi9dnluOq
xpQFpcG58jFlp3xVfXN7Zc8JHobZyaBphlUMqtrEwxJPEsSlLPBE4S73jXbLQdpx
3OZtscgyktf9+RKdOi9R51Ja5ITM65psPYKGs1y1XhTFTIgznt1lRIpPeJUO6Gls
l9OZWULwF2A0l6nucvhgqXFLSVl5rbPIVYOc+2gtSjqASdKCl2SQ9BJINtQEfUrD
RxBLzRgkOrgWsqiwzlMfbDNAgBFip2zcIzMxO/jT8i/n3Jjys/kvi7LQXF1PA6pm
A6KvkAya3UdWolvOiIfyddOq8kYFfED66rpXjiyvfz4/utKO7ZOslOZDoGlulL5I
IwpOlAGn7a13F/Wro7VMT+VDjcyTdFGQYaT6R6LYuqsucEhzwAd2MGNXS/Qmm8lt
Byp9uCnNnq/oiPM9YcJnVL8HmMtvjeFF7bGFwOSk+Zy40oi/3UkiRX6j14VfP3F5
3MqRzJytc6lSKPPMXafmbHJYDE6yC4l6Vq5eBRFGTJKIfPBNQwwJW0GbJKcRE4r4
fjGH1tvBHz9R0+GSriPu5D5U9e0rpk3szrGk5IMcFLeRRZ5sfZssNP+NUDLhQbue
W7J5rsk1RPZ4FDI+EQ0tvMutjpTp5OguWCW92Hvu+Fs6QXxOAx5d45zAnHhLZg9S
iS9L+C/6iXBOsX55pOO8aT3Ppxlxko+jLZHfUIYTWg81K1n9nq01pK4pTgbZoBjF
qCSy05S82b5DO1ao+Jln6lLw8XoRLFSXWs6ieaompYhksPSF5m3+y82bfbmq3o5d
G6iXu9eP5YOSxaOIJAmczMz5s+Ce+TY58/cbNr5tzHg0/foygEfDGPL0n1BQTllH
jMOvJPedcnDiazXuvWZcMFot6bPriVxFsrgTNvc4ergeCBJyPWL8nXrTJVCg3V9D
di06WC6WrGS0uTldpw76N16veUf/l6oQ9lxa1HDYNJitC6FOnuSTzxpHlL7gA13j
qAaRgdjGN7hSaQgpdNYeXXvlNQEzBparnNhLyJePDmNxZ9AyYZjRgL/Aa0iYdhfm
fxGnX+1i9ZG89YA6ov0OCT6OKbMo18ab1m6BLlY/VjvhXt8ssVJ6Mdt+odIBE+Sh
6MoEb6st/S427imStn2EGJ9sGVWLx1Idcsz+DS7Lga1MX5wYlWFgCR0vhakbzHX2
B5lnUonRFTHQ9TXiWRmQUtz4zQMapkO7wfznlta9Eep494GgUsaFPRfKjR6iGlhC
qcjxSdzgTVy6Sh8TyBekhHBAxvb/i1GrRzhO9WOvyqWJHfcdlesBxxa5l3qnAj/U
l7+mf2TzaqFebsYEc8fRL+DfmpOz+vdFNSZUhj7gRCUVDsStVBqZV93tyiNVUJ+x
Rk52ORa3k8nazT+WqbHp8RY+45LT/X9y5vFRIapBKRp2wqXolg4e8d0Hc3H3IyMi
R9HtV+9idCbZVuu+tCK2iPkxDx2LnDukuxPeTI7TKJykmKS7kzgCim3cCPKJE7Aw
vUAUlcrsDeB6N0uFO0vgIQMOJTqK9m/R4rRIPnjZ3I5/dLMA+S+TZ2s/O2f6uHq+
kvnVMArZ/RjRJg2q891EFNpH32gzsjTJY/PQjt73J7GBwXbLDj/X5DsBhLdVTrbX
K11caqkfuqlBF0sfkUpNweIcAZQW0MqFZbPInsXruGl2kvsvwAVRbGk69i88rc9i
0UbbhrEDSnHLq7zSeNwHcansuX1MtnPWQXu8KrItG42fos0rqV1Mtup/zktOvCpO
dKEicfr0aQo3myVrxJOo/gC5xrJQKx2b5sp20gJ0ywD+GCBLYJ4vVuDZycVOpuO9
e26ZT8d7lUogjbQnuC4mXBHiwN4AuX80kErxDJ8wmADLae7A3+RInOf/e1KSGCdw
wD2efiOszZgUZFKFx9PADF7Uq4tY5lWcyZu5E1Mp6nA0KXJv6L+11S3l66aatAWL
N7gFhs48yGlZcacxVfQ+OLmQvp82MsOB9wChMOk3lKgYKfGdSWLbQgPyrgxkxI7c
1JO7cMm5B8+lPq+THlzfqS1LMO+yuHiIKEWCLNLjlMbT0XB/bRT1KW2ohYX3dz8T
AA5c3v1pC9Z07Btt0hluIQE8C1OwKvL2L2YD3hwvQwFD2b9vvt+xvSFmGjM9+wau
XzItvgXynukeAIMsPCzCGOoJsohi//tHzfSb40YjJ+crSygpDRV7iE8voWznfSWk
VK2cfZP8l7+rpB0ZDeSw4/gkD6Z6D3nyObod8qibnO43nfJWytslmeDLIDhvHz32
e8QYBBm26bKsjIHequXKwdPYM6y55fPlXezD192ava14+T/5s0mYTXzHEvw0OaP3
gs1+mjxiSXzIGZQ/v67GV9naYcRxf2rEO3s/7KyIYPWKWuAVPUfvyJ0bwxR4mrLi
WXz9rUIxocBUxNxR0GnerXgIP3W8vtEwzNKLgL/FKLNWQbNSUvhN6TSOkRi9tNYp
MdRi8LuqOYVWcLRDNRc+0B07+UV1vBh/9HJGD7o1sjzJA0yEojZIpJKiFsdMa4YZ
PAHrcY+JTrF0Ej22mje1vsr0gF/pVSbC7IIG6TCx5QOywsljuDvHgxnLSR9eFgPv
5TqEuMigDv/tZjYsEltpmj+o8EWk7wW1CKd021jPDpjv4sqGrZd8G80erb0DiHfz
Y0XisQ6MK5ZsiVibu3qPIcxnOGpypwODLNPZEmOuuT71aujHfnkHSbu7iA6LEypN
UhQLH7q6oS6w0HSdu6ou3Kkvamo7yhW1K8Xn2gzGNG8h5z8qybdYTjMeB33tA2nZ
sICSuK4ExOUMUXvQuipBHFN1cZHLvErh0PFJZmYOHXPvnQBXNDGeJLF5YAmHetWZ
aYgWwGe0QV4yrv+LDv/54m5tOLCvOl7P+etIm/pUEAsobLLqzGkmgLM0J1KuD9tB
8iU+RPW82dwE2+QLH6of6I/xPgcFJ3BmbgQN9FjDosCOOdlsEtbCJoMVcLAxDahp
it3bdBPu8Cp8AvCuRN+x8YbBI8TluyBZgxL60jMkkMgUOn/IeTiHv78T+sQKQqRi
JqVSkI6ezJ+cd3TVqdh3tZtzSxcHs5FrtyTxlDWbrYmsrWq/fzv+kdSLBIcwZ6bC
XkdoxzKOut0JJ72NMKXlpxrmAJWd9OHAh6XMkycYx0l/WLpj/DehsEVUOJX2PLHk
7cuCNQChx/mRsb6VlN6zQArukB/FcpGYxoX3IG3OJ8ksUpnJiwaOpwMsRGqZAOjM
/aNpDCo6DTwdvvnLyTBkOQF5sKDzMRKDileTZurmzw42EUwyltmnPvibGGFpKSWK
1jT8x7IpT5pFWJPoqTv52rtJ/IjX3Z6yxpZOErjhZ52XmgSu6hOVNDk7CL2FcDqB
Pzh4ypReRNl2Z75MxNMaktlR+TQTa/pT/UdgCQEqEumjZqr7dVHVn9tj8kqpjbh5
7mjjCp2IeBwQ01Pk9aGdtztuy4OGsDzxdQtvIvgWoewlG20cozPm8Wot8nSa9pDe
5dilkSrjIdkA1FYuyKu08kkl6MmZlyzHe4IugiCsN4fIkp9Dj0MwGftEZgePCkse
lJCQeUW5RNTzTe2lvUheXtYXgnOiZCmPfaLtvV3q+99kW3SdHUGI01Ke2weTX6cH
fDQZokkWMvvXu+3bH5FwavLkz43Zn3ocl1CuL9JyLi0wIvOJ9mMXYgNzlRM4ekhA
ycoDn/ObZI85VEtN4JudDRCL9C4K04f1kd8+2kjFKQW4VfZlDe4IFdQj903RgX8C
tjgTlUtQsIUw2p2FvRNhAwexUnIte09SZYoqJCBUzBhJNt519FwecjDmpAMsu0nO
Uq9+sMJw+E/Tplqqpox8eWbarYlf62hk77uwiodz6Otq+RP+uv8nyAJVk4dGWayo
znKPExbNVzb+21sSEHpbZz/kP9YrJFYtdl2vytD08xQgTWloFgeCo2Sg1t2aqPJP
2OOSYxBfP3Spsj129LpjrfawWDi5BvtnUrogb6aAz5IGb/o2dLNsgMKRc0EZ/Xf/
MqVvxNqcxOzJtYuJzIHJQysPYpn7RNJVi5N/BhhYRc4MTd8JPCt78dhtCA3DayPF
1N5HHZ8BpJqyGMKtQxjbouzic7IjkHbmnDynWHfFOXTGpa2246EKfK/aEBo6zm/D
sLtsaHWE7nrCqQ0nl/13GewfjNW1qmiufk3U8JQBMB17EA/VHHyKPio1WojFLM2x
MvoK2uRY7dI2HPps/f86UuP9isKVGu7iXI3FjgjJMGEVt6AYiLZ15DFM/MwIdROM
6PybmlC06UW6J5bxDy2+CO2TJ21MKaWWe7bEL8N28uAVhjvBPIJu6gpADD5cV8FJ
SkQnYxn7iqob35G5W8LaVggqLPw7aD3WRW2ObJNFZ09gbJBj2GXDacy+hnos8iDA
mPF3J+RWO+noJjo9pBoNhuLaY/9rIvMlZR56ruMEreaROjVf5T+uf2gvfoQowyAL
dSEm8b4jk3XtaAsmjcNElKNnuUExr4HC5VM0O+DYuzo/sRAG4Qe7MNGaYV+SbbEW
wcAs0av/ppnXNMdAwXYagwhsExQdunLOk71WxFx41qCjQqQ9V7+q8C0pdxSTy/e/
08PCHxF2xdlRFjZehh/peNZWMo6snzJpS/Gsyfp9E6ijxOm1y8En93p5Q0KDAA4V
yK67ktk8qoLp6Z8AnDUMDjtjMIShYi6yXJY3U7g/H2t9D6jdPqifhWKr8mvaR22F
lEABs6eorKH65CUfmvVJoAN1qp9ezZVRGsyd8uEepsQE94qoiuSW7fD0bH6DeTbb
mpEmRMCGTTxERzff6CF84RLD+RrijYs6JYSo4tBqOJBbBgfCSnTyYiEzaw/ofnzF
y3MN52fwXi4CuGnPU0pKpO0wN/46zntyIi2f38LBmmWfzpEn5ojGMHHO4zak2rNH
+vSBL/TSEG4amXWLBgdLUwUPvljJ3nETBQ+ZfOQT7L6BxdBDLWRzWF8LFSou24Ol
OMxv5d7bHFrF6r7W9syV/gjX5Sh+xdothVTF5q2HBhhZ8l7j4shCieR66I8L3sXP
3PMZ6h+2A1H/acDoO+RZ3sOYmA1o5OJjkTGSNM+Lt7bEiQeIrrs08Sqtwsy972/T
l3HS9ydEBYYHeLd/IhNZ9ZF/aP5b8NSujW196SyE6hvL4hfu3CTSnn6tjmifZ+0i
7jsypO17DTFXY+6/VvBe+gg7SASWT8o3XNlojWwNOLZDWQ5+19V40srHLoOZWyfx
Fuh9g/PPh0vTqcdYYToxkKPJ5fp2kNviDk9+FGDaZRji10zzElA85IOIJGX/T+HD
23X95pEWBxBqYBmeMwbz+L16A+xdQxyNxCZfLF4B0m7b2gJa9+UfruHvkNbf49Wm
AvebqeP4C/gKO0XVJuTbbGVs727fYAFavUR4uZ54iM6YUJmT9pLEX1YbOJez4W4z
oTp/EffG7plkIqrrzsFXOca/f7q+62gQLfshSf2cmsG4sHFmXBGRIzQJlZ/8h+/R
bGimzsOK2s0GQ5+4L4pnXD9xYHSz8imGltH90Z6G95919ZvQUw/brflKlYW6+T3P
3/H2ktrPLvOrl8ri5egYQ5uKjvMDE05Y+W8pLF9pBvC4k+ee0yawB4P/ynHViSYo
mG80gy4bd6e5Da7IcvFX2mF1fGmxIxCJtdZVo17AOmTZlmTSi5TTGrrE5vCRLpUH
v7aL7lo1l7fQW4ED3F8VdKCQPj72+PkbhMSDvI990Pr3+Ce7Lvk2JdvWmcWazhY5
U3Hgf/vJ1vqPlbzCKSwzAXjxWJo/vWfd8++zNKW6gcO0r2SVkYP2vdqVOHZWU5lO
dj9Lx+7FRurqfNvgNfKJzILZVQr4K8AyY03pQdriHcEcy0WaNMX49cwxUoTxq3mO
8rQvEGtlIfSJGTU9kW6JHRT2nQPDPmuME+Ta+3Cg5sHd0vxPQb3xUCueDDnExGS0
fUwYo5vaZxhzI4lZr+KuQe3tC9yRzq7gtwpUPsua32a2K0QfLqKI9rseo7fqs995
VwitkQlVobQX+KHRAlR89FJwowvabm13/fYxv0eEkWRMhW1bRvUqKEKWAHSJajOv
o4w0AsmMfQtqTY6869U7ZRm8x39eyP/W6BCr54NZTW/7B7qXKbB3vVrvS8YTOE1g
PznmGpduvx63jPxawNbmQtyZYiPtAUlGjDRGr/QjoRgsKaLKxoIN4VQ7/Bc4jvKN
H7nsrrbTTRlVzaC4IHvMBj1eosScycAUL+axM1IVbWXgFSKwvGL/9al8Pc+Va9nU
7k3g78D/Agvr6Qog/AnNMo02dx0MfxmxgKSWqL30dENa2mPNb42xBOBAetCv8AJM
bb0qffxdauOEH+ShixsjF+z2fqbuitksloadsGUC1JS0/2jihheZETZzxbUBv+iF
PW+Eh5T43MjpQuY79M5cPdXbypdWjyWI7Vd0ZQuOqBTUkM2xjTQ8iA/Lp9AzERbD
ArmeOYk9wa8rLk9VhNfHN45xmxvm38ZS65KSGoCdt7YdHHunFpRCSuAOvuZgBBv9
0bTnaFF0OojMBJpuL+4cJgyGhXBdDbFeMzZBRYbki678YqzRKSn3/CTHnEwSYtlg
3vXUpx7KLmCG2HWQAK0AuEkIaXkXD6Q4r2syL8x1mZoG0YP99G1RAXSrbvGauhUI
rjKqcAJ/k5FPosExfDMB5gH6jW1x7vwnwpgewLFAG3/mJqxufcB4FXvlSbN1qOyC
7dwLalndpVBlDD8q6apyS+9kyOgxRjiha/XVTX6y9OsplM+jknzZw1Jkx/GuFmFY
woGHkDiZEnThBB3ydYeFS5I0qH10Mf6UweoZ63Ox7D5xgMlGwP36DwKMHNzKiZaQ
GKSsvBhifrgVwi3dpbEm1DnCZxe8VWVeSbOqCA4cb2qOH9pNX2S6wCnBAbN1RCFl
Ck9U2AF5k+CC8m1nZesoKlNL7+eYlxdN9MArNRF4cjwd1aoWzFCL7bMJmVgb9bHQ
Yk1zFuzknA9N7frJDm3D0lWipBeUeBraeIknI5U8O6kVaik6XsMW8Z+qS4r6sAHF
XGcZKdX8YjtT6uMYqtdsf8eK9uBT1UFKwzXzbisK9VOVYQIoGbaI27NYld1Ejhp4
PRwQvIQt4M9w0T3AVdbeD6/1bPMOiR/Dmz18iJYZn573f4IInwjK3o8lkBakZRwM
1Y0AnRmMsi9nH/50vfJSZBj0o8DlZ+KVltlwqTWU5l+8DzvAh2NHOGczuXKJW17f
WMCJZP7MpJWfrUnMVdcvx1uCvz5Qz3ibj5IEiHdwy1zglbg/EON1ei/Lp59N3CSU
7COlv2H2gvWj7L7kL4Z/8sUpBiIjPU1lF1pmRumj5Q4oUdvONu+pNleDJJbKBt8Y
sHrII2e3AcvdXMFGZ8wFX808xLFPwpx4gMTVIeVyz6sIZIBaolnhw7jNyCRwBuFB
uDUwqXHXa2haUZPIvh0ycBHUJycAsegWGnwEfEmu/a2nG3sh2E7jQJ589GwKy+B2
ij12EgpZTLwIilrFNW7YgbDN7mdvRJMximIQvOLMGHsgCuPXwIWwseA78Kw6eRXL
/TqojmfCgydJMtfA0FcRSNdz+3qbJtlVNkBHM4Y8OVjPslhUvSJ5DqHLWSg8s11e
h+x8//gZTKUfCRn+IJ6wtbva1ao8hWaq0QAINz3K01i80Ri5Vdy0PldUml3nbS8E
NTqIAlHRA2bbzhRow+a5MPRffFF2ja9LtC7ZmJ4p/vL9LP4njTRuZkSfxq1KxMFR
dZD5T8zkHLnhSd/Z3eGBWu3QPkZTkajNntRfyP5EvBrfbtHwyf5EthuOfnivJdMb
uZgPJvNO9bNzRd4tJSoKuFz2p83eANKNSc0glEvdHakX6Ua/JDXmeFikCS/Oigkk
Uxoi/NXDhlc0G+BSx5U7/Qv9EaEh7/she7hV8XIBiJdm1slup8vTnot7m7Sg/PHh
veJ0PBlrrjj6v4FaoB8J8Hasu5qx9ihi1/gv92UGmv90CnOOIqC1eoNhkFAQeyBv
1XDGtfosvVPOrFGfe1G5e4gwdRD5dMMXI+AgPRATS4zHKnsPmmsi2ObC+duJOGO/
V1yrui3m6SbUNPtDXiF+W75E1f8+/IsgKAMWbv4psoQKO9C94Hs1nx1Mz4yNupui
r3VEEWsm0YZF5Eupfa1q9iBQIDo/2KHsAU7+7MRPdz7FiqDWfgCxKr7c7pInuebm
ZanEgQ/IrLctPScsvPgDFWcG1d56QOmp4JUbhZ3ufy7837D/60P/ptT0qmrJDLqN
3t+HE/WLHxBu3HZ/3cJMJa/SWZ0Jd9MzHX5dlmCX0Sv6109ZMtrlWbdc0BJao0Jt
dkddQfVNsbkjbwkdzSVyojyVRKH5LOHJ1AXRySFkWgCLP99zjmOI7+10xqa6jkD6
5s4jgUX1am8v5BoY8f/ROK3AA/ZA13EsQETvk/6TlUb4nF847qzLh0KRVNQjERHm
k1P5G3/klWqks72rhG9ZbcvWC8ljInH/YzEchjwUGFVe1KeZc/FQrdE20gawSsvA
hUzgDmkqsySvpxJhTfONpzNgRRqASc5mCrf8UgFb9GmJ8BVsXihONC77+jihZ5ae
aZvJmjjyVIDXPun+nzlRQwPQ3p2ZRznhjwkAsJW8JOMtRrBCBXla1dWwetlffjra
nR97TyjT3ggdwgygSbM4DQg7s/4XE0HK7r+uMxQxfTy5P+HqAFCriD3txTmkLghu
kqw9M3DLUo70LeP0Rfl2/wyxtlGiLYp/0eF5LGIwjS+rmd7e+dmdKa62VDqjrgg/
HsXvEwmprfZEGnZK3YxxquuBRmKzX9m9J3KL3EX7xHvyFPO5NcxMAUx/JxQ1uGcT
VrQ/rxkBf2M+b2pqUuXDbfMWvtZcw9+Px1S0ovAjzSkq4rMdb1ic2rHptdZF8NIB
AgN7txfUCHS0TWQD26exyLPKmula1awR6remRbRBasZ1Za7zSp/wXL6UfxI0Y6nq
eM4HRVGAGER9xlVF7EPLHOh5b40iMnEQsCB2yyBaWdaTdpDi2tUpGfqxVRKIJGhu
oFb+YU1/3aXzipeQH81wm3qa67zr8LswHgqUni5U1TKfssm+rIkhZTDoG9JnKo5Z
K1CtiY7Mt35Io1IZ/aTJ8DzJBOdHip6WQ4n1AaJKXh9ZQ8T6BTC0aWeq8GLGVjkX
DUTzbGjIQpeZMLhukjjC4RGAWpX8r6JWPgMxiHtgk7LSkf/rou9FqzHfrqdJtfR9
+/0qzJ1qrxlITcWrqd89hXy0NynCwIw9Se3N2jAYkuJE9+C0ciNQdOr+I1xh3ESV
IRD2xOcm1GLalt3dUfzURSVwmfZDQfHmKa568xndHPTdLLfJd6fw/RcFWarhREPa
4ChB/gglt6iFOYOA6C5VFOyhTpg8lFqQsgY8xmyG4hzx+9eSJYeDNkgRVs/5RUW8
MO0cND8BX5rBQ32qvNidttxeqH3Anjn9xk6yJAh2TmoX8SY/ClsI70N0iWOuZM2q
ftbkTsgcmeiov/E06etNDQVjnMgiZ0aj4URANBsjSuXxV7CFuw/dT8FN67POug+z
vQFtmMd9WgBc8FTgTux5yDO8iyFSVD6DjyCFBqOP/IP6gyeR0dmFwJnjzXMTqlYp
ea2xCuGfNeNUb/0+giynJoW66QbX3Aet1ARfGarYQ3qHaG/AwRcDHRbcQSYOFsC5
yqJQfUSDTlf93erBGCf5oYUPb1K/QgrPlWUGBccFYcQ63K2OUylUnNXITDkaABFp
cNusZF/4hP7gCI6GLpdjlUD++EujH824OFv/Lxv+xSHqj1xg6Wk8B+Y9tboJS/FS
+AQlyqwK1IsO28GHBnYarHXAIJkyhqtEBQbt2KcwZ8JMNn8apfRtYhFcK0yqPVyj
2xCbLGDyigK3osy+v1qS608sSaVLXDR1SpmcRRUuY5XNKcO2s9Yg2r74VAXoe3IT
b0Wh1fXiTvqrJxgNDnytsOUb8zLNj5p96gmxmx628PfC1e5Z+riTF+hwS9Iep89b
g5OzKdOhRUcsp0KdWVUzEga4s0GycYDjN+FshbOT37Ij/SS9oKIAwdKhu5p4AwX7
NI/nl+k7eA6CeU4AmgImzxkJTvutWkvezSrhGlZm/NW9cBbMv/5OiksT5ygBHijs
f1gngmlGT7XTQ7PVF+kBcmVFIrlIy6+iXvngUxhfa2TXNWTooP9B+jIdAf20gYnn
K9nxwfWdvTJPlFWPjy4x1DsmYhejH8TRGuUMVAQn2N54X9ozWekuUwGSfMV7jWW3
yR2oVbs6ZqKwR2rf7psbYcAsEFv1Yc7weQX7fpZHzoH8qErjvuk6YZh9RZb/DLY/
VE/Ix2OC/xzH5wJXPwSL/5VAW0R72LM8PN/ENG7J+U7b6JnGMaBPjAqZWSjF0A3u
TOHBWhl2EgSKX8p7Lg+DGiJng2NzFzFFEmolcTNbb3VovrTD5l6JxkvsNI3uJpVl
GpySOmanSttcF+zhcstpz8d0WPPV70kLeyG6NQi7wzvHREvcc97+v2yx8pTYzeBE
teREFqxUSqzAORGG3xOtvwqNSxT9qFIuoA/KELLPIvsHt0wxN1UADlooU/4hyji1
bW0ZL+2NXZVDUHL8aXi7c/ucbTxFWhbKyNLjd/3FJsGaroIxroleqp0QahD/Yc//
5O6+2Rekx11eVs4mquQtc6/zNKO+BCpVyY8sE2UOzALyIlp/7lrx1n+Pmq4cnzI3
7QSBGb+7qrYs7++1qXWH9pvwNiOt1i0+uswGGYTbxKh2WHjneKEBJuVD4enn+Pye
qy2V6+8XbTA6tnQRiSl+bFRGJ6mdsiiU+4UeANXexsEiS0LKNKWXimEC9D8kLZdf
v9/4NTMc1rIWTtIimVki/o8N7EV2wXgAD93IqL/+N/ANYHEeiEYq+ajCyhoJQcbo
FL5b5ZjkENk+D83lETH8IiqfbXFJqIGICrDj/Hf+8qk+GKjkzq6He0FPOxOwjLtu
WXbAi6EduHIPf9XEhDXSVfLkuYnSujSIXj35ETGVIksrEUizIcTvleRWplCC6q1U
be5BCCoV1eO1r4yiijsQtAlsBvtg//gQHyhp1HPZHvkG+/SryyPd/PC5Hin2HCaA
5tMx83yEBsRNc5jUyF3IGTI7BFVat+cjUI6gqiN2P3dcfZPePlwU57gFGr0Wh/QR
q9tI82UtJUTk7TVmLtC248D6Uxp1Pz91gKlu6SHrlNG+yelCEEzjxlyetCCPs2Fm
cDV4/D8xK8TfUNLhlikno6ajk5/IVLyTF0yiD1YFdInUiucR3ZB+19hqwVqPoQMJ
2d5HShtyPEtnghyatLJiaA2h8mxA7aAbO3HNk5g9jqZ86r3LgUNNRQTBizzHUOlV
W65z9f8EkHiYrUOfQ6y3TxkER7oPfWuCMiSNjdmLmXCsaIGrVG0G7bAopah/DcFX
ftN6ubgpHrZF+mm5qCnI9JbZOjTd6dUFd/UegJnX3UWvNcl4uggISVXlrNNTBLjs
Gtra7Gtv8KnHnnH62NMxYVW5xKRi3TVNJnmLaRYL8N1nZ+bd9UMZevL52OKnu7eD
faYnT7IAbG4rimkYltdldK9w2cv82Sq6CW22Oyl545YlrHkrM+TfZWVpyBBLTD6M
uFJsVTD0GXCSTQ/av8+9N9VZKMeTPN/ohgenAlnp1SJw6EH14huksJNleDmf5Jfb
GkiSGQFMouR3k5DwOeG1haV+2utbPX1+RK2dB6x5ADrQXiBhO3CKjUsuk56gt2i1
xc4TbMnvXJAUxpm36nsyHPXLYKW5SjgL0SVrRZ1XnLRzmWva/dGpwZD9CkLtuPhK
oqAQiOS8iyrudL9uSFpuwAMa+yp7MK86Z9CW0NzBY/UK9ML/42LLC+/x+Km7wDQd
WBT1KLB0AlIL2IMhxmHn70/OzarK1qnfk0jP2/ZySi2L6vN+u62gzFH0PxyavPQE
2YLODFPwSDJR1OG+73MlAzfsesv9+LpTJtK0ES2lowH+tdO6Vd180VGBeLXGRqdp
ylITUd4jrFn1WUQQVcwHPolflhRmY8wtUZIJ6lt9ZtBs+ejjHncWl4LdEt6PXyLu
/lfR8SQGPJ+BHvqwVOTZrAbfK93l5zztzC01TrjCnXRrYWwi5OBNHeyYHoN2aXR1
M0z8DqMM1jpcL91stVFT4ovx1Np2nll+y3MAqaidgJqXj02umy06oXepZbSqptI+
vwHGzZKE9Ylz3t9uJmDx6U1TZtr0hYrqFHC9yO2lcbmoMDnPEq3b++RJYaFkSlxV
U4GE5Ag0VO4X9LDQQD6Rk0cp3tca+TtXvG5OkgYBIfqmfw0+XEzSm1M0tdEqWhf0
mkreXhUtBkblcj2KqpGJXVSjygybrrcFl/pXSt1U50/24abRiIGMPwMx92OD9zgN
oBouGZstREFQfZUo27JBmHoyjcoIhpDNvUXx2a9BVmYT+09LxROEduZhQktTbEIP
Uz99Oc0KH+xO5NOOMJ3CfoNkfW9jSIhbyxC3UqLpdVgXWSTeOTz8iPqdPA27PMLm
hOTtUn6J3ENzJeS4U/bmGdsj6ZyNXbujDeULH5oY+zDL4Ld2uizx6qWp7li2QnTo
plNpJiYU5H2by1tt5jAZslvoytfUudTmok4qpkti+iAsnVq/vPv1bZlsxw/hwYxw
fDFaiyBgzXnEnvYL3kYgK6cPpq+rnR0uc4x0MWeeOEtLgQt6Fo5bOTlAJfueyew/
3TIXjWeoP6YoS2A35EuXc7PNfJZEG94XZ7JpR6h3M1bF6jodLQ0SpWnm3H8CYLzZ
Gtjigea5lvlcGQEBq5oF1Kom2sCYRhJr7Zh6nxr0DkmRMmuZgezvavn/9Wg8nEUL
MuLaKNPH6C/4K2aTLBVsR7kWDCobYJu/GEwzoln2fYMulPUTmriPI7JxCupMc2xb
pQCeO8zd/6p0f+qbbAffgiCRn63mvgE6thB38GKCTavwa9hthPR2fUdOaJm8IoPb
CXxDXKOkb7lBEYu+Z7oTaovL+qO2GY2gZM4C8Ah9C2ddygxPF7713sqOIQCpIkBx
mSYOXpEXlszKR5IYMQrPkx4HS2S4uTG+o0JNQlZIqnT5AKWN2uujvMCHPWP0ljVE
73uyhmCg2SvspHGprdm3y13cHrqMjT3GcDT6xwjisPuCp/n1F1QRF7Al6bnfES5T
qXrQrOa8R4qH1U/cdKJHUYvyIimmCIB36f0hGjao9HVSpJLdPFZdeRsI1107wH3S
y0cD5u4lXmiNRLgTYC5ztRnoSv4esoMxVdD/MsSSqk0i/yV/IN+eK7pYunrsZIKI
TIy7wRS+/DMa6xpT6OIJW63wgzVwIiIQCVz+N7HnLaJEmUX7YWoDpZLs4uk0H9A3
cUzcwPfL0tQ+1Lh5EfRTYgLW81wjhMDN34IpeuytZBXVLQO5Iqau3WhhHYAxgIfA
wR6osvWL6Fa3gq5KzyymmvXsKAKeflwChxjV0IzY/74RyZae3HINE6Mrn8sG/3Zd
ghHnt7I90F6JEFbMePtOSMfgpFTnd0vninHNEKr3j57fE9Xy4byJVF0/QwcXRUBk
6GAeRIcmrLJP4dSLYmx68S/668b9mI8+PFgg54BfUV1OptTFKRdiEQumGpYRGhBU
nEBgoTM8NcpJYMGTOMa6+XHgV0H9WX1BWVEJU9we9yWB6DL74LgNIesqP1xGqUSa
8xBIiBIDc6QhUqBQwX1gZft7SjDjQ9wbQ/UfSKGdjoHaIjDPpVmS6cWtRRdZCmDS
FCq4esorUEAECvkjTp1NvAEHH5QqfQ9+xG13aqpB6iSKZyeK/9ixpD7uMw4SpjL+
YLhWkw928Lg2PZHRe7dttw2ZxnBV5khxaG9fvfnbNF3GNIxF7PJ2OTZrf1PeHccU
3zOk3SlnAPPbmsSQWDTnLHfAWBhnKopNQWMYAxjWuOel0Ml1m52e5pqE/zbU3BId
oTZFZmJ4RLnjmGPJe895xAw1MxuZ+TPQPpTTZFt6lezwhO/owsTS3IdrnwSY+LWY
ep/Sh1XmTdGZ7gE2VKkpdAM+jQg7qLUWBGqnE7Pc2gi3OxOl/T2GIowDfV1XO1JI
qunaHe7n0o4evsjyTKED+DisBvX8KOAF16PxrQqscEpBIyJkXrRkTPWIhFklBEBD
DEwm7YTVEJyPWZMsqHC+wwmLYiDa89EM4jidPr5FX2DFRaAhglY6oVbhnz0MHfyR
XxvaKd/HO5fuIkZBrJHX6gbSMY+05t882vO6BIbj1iE53DI67bccCNpTnPiLppPv
GxR9ReGinoOY3A1T/DSBzeQb0AVNTj2h/IJiZeoGNVFmSog5L/3LX3A40aE2I1NF
q9EvuF/KtBvSsSkY2eCS80oHXBDAK5XOYyui8TZgJA609ln8SpkLKFO1TT2MOm/e
/gWPT6tQBQT7zUzdISgeZ7VGvEP8kLIBvDsHbqgJW+B87PWjCqppm+tS+uCHdHvu
xXWBamnI5feLbFsU6iTFIBwXFpBbPqGZCzZAwKhZ6ugcWoF2v8odGsXwP8i/fu9I
pbXkq1LtsMKOzgTodE/hn+bLVo/IVQcciDkLPd2kwLpA2g2P/AgDXZ/7K58G14lt
sjwBxpcK5+QvOS9bDPHGwyOn+LkgxDi0M45EiE4tnAV8/PnaFR0T1jC7anqIWUxH
9FeGLmIrRHeBbME7nzL6Xiwyr9tKfugB4XaKs+YGpNjQslIdTAFbVdYH0EGAvBNU
WLUDaEwFZIMWXsa4JIg3Xf8qdtfdmHHWWoHf6nbKirXadcboQW+gGyAgQ464SFUv
Cm8VWUMDdGrVd9bR2wAHyNWZI9rq71e/XVx3JMwwlhNlLaLgdS9jCU0ibpofDXX9
cK+N8t4pwLZFLtZEInAEkaJ9c1Gi4dFxdw8VnbnX6YOaKQAXg72YS19MlJQ/lR+4
xCc0spVQbTEHXxKWv9XQ1fgfqGJIbqYL8OrlFZOOTcDUczCShaN7TB50RRGn/aTM
6F9R1gPw03UZ5hVqb7KtX8BHAYGUQlBSzXbQFOKn55PE9vxh7fv1xVtTzRz+0+vf
MdVurfrNCghHcrefdxGwxdm5E9QPyuC5W9TJ2Rv0aXk3o+RUu3ztJA0qFyViad5D
UwgTbLADAwpNYtTDwfQZWe0YefH8Nnt8oI7Z3HazSuq8OjGHCFtjBPWPaOAZBlxI
Qqk81dnRWIrQj5KITv94K7aiLQ+/zs1pM9qM4LjnkNKZekT/r+m+W/ETRk1M5EFt
YA8TlpFcg0NRh5P7PAKkrtzMm+WRNLOcCEmNYG5qq+A5zNKWW7/P8fkiR9m+2xFp
p9sDxXpKBSEJqcShbz8J0TCEpD1vLxYSEIQwJz9NNPhotb/o6oNXoFl5V+Lhwbq3
b2Nt21HLRqpzAZBOp3N+z3pjnZOXi37gi0Mc/QjR2Dx+dZoMlr2tVsPfloqsAdgm
5KsvlohYo5wqAR8ZNwAhJM4tcGkGx2mgqzMpmrmHMlM10ilj1x0fKMEdi4odsRJQ
nPgWlPHNsmIRpsvMEuE/rodPjShhB9fPHYjRTUW9dlk65v7/RmP6tkZM4opgS3IM
v+sEz2EHPcO22trQ09t3cHv2nE6tK526vrOxfuSwwSauvSz0IZYrmCtZ9IDLnsRp
uS+BfIxFdTn6Rm17H0xGj0BrVM+4S2yeHecLlII3d5FAgVzWQSDOMgkgkxhZM6NX
FUnbDJ9ncnEfjOS4q4GGsxhYe6fa1aVE7CORul28VMS9ABuGlwLJ45JM8B9zddVS
x9WhuX4qQdxBbZPqDlU3PPu6EryjzXW4Io0xwLfSfRc+CXC/LFFxN/4EU8GGuIhc
ySmjxOhoa0WvvXHsXtvmOEJ1PNxeuSVCbt8hfySn6MtqZvHqdpwXFhadhr0/9/hu
zBr89ecxT2XkP5MRmMuyIGQ5wSKtvWSc7H1+NYk3b0sPUiov+WX5gx43hm6AVicr
g5lVyczEOLrPT+l8nLAqHSLBqLTkcW6flYzU0DMtIyTRtV2hZeb+7DzVhuxufFJZ
nuyrXz1crqHJqmxNgtdWRmWlClMFMaoSb8nfM7PNEWl6toNWRoeCZhxB0sTKcFXZ
X0SK9PPRfWTaii/L/OHAstEyK8el1ROOg93SH9JPcW7MMSEiREZ3GHTXxKxsv3b3
CCWpVYOz6YMhbJRePNT2/CS/8+Ss7yUvaAr+HfvLA+VFfNpdMxpM/kqsjLMYwerE
o7YP5JMvniBUQRSDP3NpGCY8fv6H/JT7s3J/Ii3Awa30dE+y6MMjsquAo7VZp2iX
N+bNCYczHVYZofMA1vpXb2LSFgot0IgPRjoAg8TZtvu57tjY61blxjxSRH3nOr01
4iu5EraC0xolWSqYvuMLm1mZNPSShaHpw7x4a7mxFXpPS8DgEbRwlks4sfSqRurJ
O3a/LSkyV57thNrvZkWLTadXpPton1tEgSS8Whffd14azu4GV3tm1EXu77e3CYlS
s+cxmoySwRT1bXUPg43K6I2tIMX07HPOVf8dcCK9dU5vRg6YR1BD+ZluFt3Uv3l9
iv5aVhZYFdVEYZK0b+zeP046MX09YRDo41pjfD17wa9/kIBAfw818GJElIA0DTLE
PnG0cBv74LRFfeh2a8Of3F/MFuDC9S2a2dbWWpQgj2F3rxGBa+E75v1BmT2RuwAe
lYIjXyZfNYNQbWsRAPaI9dZfwR7z5ZiOlalmcbawzx2pIkneFdjHsl/foF+0NCt1
ZXCPZ8hpeN11c5pGdoM4oBkc1u7QCUeESmaicfdQfghgt2xJJMJUEFTbWC+Km2jF
tf6YBhDLRJzV1phkIxse7z6EyjUuz78+pCGoW2lx0TRnCUpYYkvW5WODrMNhfhfD
Y+RiUAqvAjALFtzktqxJwjdiRN3C6rX+DnkFo8UHjGiZRq6ISNchTKj5Gz3ugiFt
vgpuk9LuKNRdNo2NRpyDlqMfNZhtJo1wf8f2Okfz7u6zbhZHobD2sQPJLMCVvL0W
siJu/hfk8VhqME/sSdI1Xc/VUh+I3MEsBj9TfWXGbleL7KttDMmQonab4NrKWJi0
VzerHGjhfn3OSjpQEcYhShtGM15y4pKrVMDgWNPIpcE5y285M1aymh72XIOdSApC
0oAD+YjVdMBAYVATxwJL5WOI0CMe7DK9eC0TAxx/sGM0piYNd3VGQ/OWSqXqKzk7
WHctezM5bZKSrI9cur86sf7Nm1lo7n8AGDBu+2sQQ7itbwPYuPjByXkVmwFzKGGe
PN3Jwc65jf049z6pUxXWhi2Ka0b8axom004hBmzfkZk3GEqnP5XYyvh4qaq5qmW/
GLIGuPc/Rwmky/z8QFR0RGUpaVD1SrXk9cE+v9TPkoqljr4RnqXdRjDtoAAqreW4
KKIZdMwLOrJY1zGHp2soP6tLD1R1WwQr1v0DWe0W7Nzq//cu4Aqu3IX9y759ydyF
lxqJRTkvT0TIze5RXdi/oiOwsODPkC0WbTAAqZ/HeyYKhkZ+3wkiGdujFZZ4Zfet
v8DIDiguasf/xBosiGxvDX1J8So3DubYhFNgisMwxmwClmwJM+fWTeOkwE1NXQ1j
qcj137pTHxRHPokDolnLrOdjIYA6pmnU1LpOIXMgLgrhUGBEjSQZT6EVR3EWOaeS
4kI5RdGEVpKX6SCRno/wJwrMykl2qqSK9zW5UCdsf7Ptq/EltrEtfk6PplXd+wzp
lOmiNsep0+SEm+A0hpG6iFwINHPg63cX2Adi2Oo8Xs91CVSQoxWoCjdBjBQlVfTw
MP5VJJETfog8RLsNZATIux9/VTQeai/3hUe1qY7er/aka9eu0fd6euaBhmYfHm8y
CS3REz4S+oph2lrGBw819RR44q8GKrOeYIZ4D0GxtDJjY0OyhtHl//y1eCkEP5jp
d2JaYlY79fdvCrwvP5moxiEnEBqhWhtxI2hvE4/sijt30R6L+1fpNOheau681k5w
Uk1U2/KVIJXTUb3Ic5OSyorEBZ3JGReATx7O8CLlZoQcMLhcFPhPZ9RXjEKd6cRJ
q3GsED+SZtp/w64wDXAD4/AGb+gFZO08K7qP0W687BtrrVdXCcV0z3efNa8oHhyN
75P0dSnvKhrPfXFYhDQyroXpC6e4Xy1AONKwBrVum0cfagOH8SMJsStPkFg2V1He
O7ekrl9Lh1Yfz8aG9CWLy44Pv8Ot/oz08Qpf9xjW6ARgKeNNsQO3uXpMi1XlspUB
KkdXvDSeV7OftI1jO+ATWn2hLzQeA06HBPILEc4Qylm9KIbdXJiWmrrStuotFb+Q
qL9M2zN82IHdgJ3NooV72FEif/ZAE+J7H6BvdWu/fOhiG5aoxvH62+UKIqBXQ46d
agN/3DS5+nuoweZOhC2AX3/yJzxzAUnWdfbfPS3xxupl+9ftyMuu9ULaZAMgogU9
NAupy8YYFQz90efSsb9UKZSyjRxvcxo9uGIZB1FXJja9WNYqWBdr+QLioC2LZIE5
J0jmfUi5VG2Db5GhOTLPJiThruvzqZ2SPTg/fRvFwufedWMWvddbUAsR/puNTOCS
ih9oTCGhrEapLfvC1RBuGavCSl5IrSJMC6B19fjiRMj6ZZmkPOq/CyQX6o9rKz/q
oMxOCYNYzvPjEV7taM3HJZ/UmpiYp6nDgYXh6K9tHaoS06uH3RtSS48Ab0dHqjs8
BaLdaEUWpXQzIze/tqZMRPqjz7mbeysTnVU77Fj2My/B24L7iS6kU/TjzOu5TKr+
NN2Nk3SbQAWRO7lppA/m3Wv+FdugEp/MXfiP/GXqqegMSwDzrq55ULxYRgvGHYLV
7CMtMioQPng3fJXFYGtnubZ+0rg3AGTFVQa6gjmwQM42SIPEBTpzt2Mgn5pRIqtq
kkVkhFk8zGdRECKvwcUWCsIeern2Su59d9yp/SDBNbFt39rz9zJnTMK0oA+dRlBJ
Wzo5xbA9Yhublv7UGhG7GXjmizPkspcuCja1PVd2o1EM5d6bUn4RaF1g7lA7JQ+V
RN3DO/du71hduU4VUI8A4F2zUEX/oakRrBe3iJ5uAg579lrZOXhTC5uVZZs8ymR0
DtmJCB33mSqRBbH27Z2gGvZfuj3usp02Ja/vHZIhGD8BYKTpGCx0ITgX79w4lI/p
FJmJBsgkNpgQA1eny/qO6V0Vk3Sk4XHM1T65hT1P4kw/H1aN3re64QncY8e4QXHB
vNnChJX9w06D/y87Dy1ghKFGs0tCTiARIrwJ0rQyiwR+azi6SFqkxm19GBilfHvI
qzr9oX1QwldjsPS5Kib+za+AD7zjd1yynwLb005/FO2zxyxx8Ygija0D9wBdwkHS
FmRF4evmUgP1BIxYG6J3rETzpVfw6237QvZtxEWI7q5bIzChyAazNx4nmRxrmfmA
3wWeM9bep5DhHQebz38KZeg7EcAzy64Yiwn6HfcrnmTFgO8MQT31mODv1MEDBBkY
Ad0C0UDE39wlugunpz1Tet2xUFfdscn3iVErK1rUf2tNwnlfdkG1m7bRzaWU3RMB
cul6WeXbpWMcxKiGkwXGZ2YEpmu/laAEKrAbwKju2aFY8XgzJw1Rz8JPEeyghXYz
G/OClLnMQIubUz1nT6361u9trEWOrsfegCp0S1Xc4xXvHN40Blc5An0AX9T2XHNu
BvrUNdfpZq7eikqFzlcXSt6XTWbqeXJq/h1f7uUjzvxxM08QaoUv3HpHNky91BpL
cAyBls28zLKrxdUspC70bELq03BQ4iHDyvtdTMM7VExtJ+QIExygY6025MyL6ty2
j2DnmnWzqRScdIwYpOshPmp1SRBQziD2rrvSMqYvPPsk0qixQ1fCDcSijqFUQ3Gi
EXXJFvrXHnpkpd43DgIBN1F9aCrjtSYC62vHDbxVYVCJDSEXSqVTVuG1HvAgDsIe
hXxlg0se0eS4i1INSNM+kMcmWf6JEdFDpn8zISE9bcerzOG0DSo23dPEopSAO/LR
V28hIV7bqAMO/OGToG8TaNNJbrnsfN12kWdF9i4mpcIp3Vb4eI4huPTCU+tyRraP
FfQpB6sKsmXG7rWINMJA1LmNicp7uDnVihrD3gKO4ie9eHkr1PUduMNObO7C8RLS
/Sa0rzDNsZWeGJagesI2omkV+e0TQkTToSwqgxQTo21p9mBOYDW7iywsG4euDSVV
MtFqqLgrcwLFY6TlX48Z859OwB3BaKCnm4iIqz22fBuBAMmDerXW8JWELP2g8N+8
XfLw1zFtedrPUgF2pWTqiHnPFPT24sHgGgyQswvBb81nnWUmQEaiDWB1M4efc5Md
/wBBFgk0Dvoqn4jyi9sQ0x5ekpL0hSaUwi41lSorv68rCRlqAk+Z6uFc69597nRe
wYltWi9aU3XzqH5aUeK+HBlOEiZC9LDYqzho6d6Xq88DD2D3CeXKA3gqpaAc7nfR
WgQSgolrQErg3WATJAryYiaQZDeKAW/43wX3SJSotx+WVXuQT+mdPx/vuFgmRx0l
z4eVx6ihlmbTku0p3n6as6Yj+F3EMKp0f1nWBMQhCGU0h9UdOlNtxIJ0hOh4f2A9
UfP3uXBfRtfx4lcAnhoA7dDVIX+7u6cRsIc9kkhp2/D4FJj5/xgr7dhZi4bh6cKk
q2wdVM9o3Us8OctkAqQ15c9jvI5aOPr/aw0jllV6qwoxlNerCF9tAZQE7/66BAn4
A2Jhy8qmYHbTKKYXq19x5yzWQJG2Ejah7BnW+XP6UHXCwgXszo+n6WJYhODbxFNQ
jVHwWVHvY5o3e43pg5dkHK3AOVn6nK+7vc3VjXVaxY/jgmV3QjAPI7pnQd+7JjnW
ZCOuzryps8/G1ni9/Y23C7dC/CHDx6mFGZlqoUzTIGI68DyGp0wj649YgPJRmNxG
hVAhINlGoAV1Lf5Pqnw3T2uqhcoMumdGzWhlTIN5N/0S3TXmjf6Bop/b5PqDR8yU
pC4xfJzdCH6PJP0c3rZIkvmUErM7tRdAgFPAyhFwXwJ5/xxgv+4yM77ii1l92jYV
oruMhD6mvNN6eX2caLhUv1YCgjEcgHn7Hbf71HHaj/l7OXJT4hbrFZoViqYr9BuC
FoGdtUodsoNCmHq0NXJOc48z1Pvh01j3PRHDwbkwB9CTwDRFAeqKqrGo57G3pPnK
V/MAeo7us8RsXV/rCxNlVKMhE8Vk1KkX340+bmz9ewSBJNshv2iz4MVpLUamXQ9j
x+5EpWFQA+Ha5rd/tPNiUpg6Bs0VIXphL3SKZNU54pabe4BzqT37QThJnIv7Fuu0
8gXhIP8tC9nc4s/RBGCG5pFsDdciQIxb45cOfxVu33+ze1gTz63ZOXgIeJbuQ3aS
aBRmbBZ1sDH+CFEeNI5eJTREI3SwwpTgFjLO00rSv0nwSegcq74QRk0oIN15iksC
WCp6Glw21NUh9ZwAtt9SRdMIjsyQvH6iQGDxqDE+0+ZnnssmhpSfdEvUTUGAaLzb
lhRqAoSPT4Mp49ULSn8K5aC/DOEsxkASN62913dlwoNwTw6RPZU44GxgrSysZZav
A3EXenFbxqEVntcc3JTl+cgjcrYG83jJwTNXcXGrsO7bl04W6Zi2LggrDigJW+Uf
Kd4XayGS+JAP3M3nYHjfGpnYEQlfAYXnQ+siX2lOsLNaCVuS/aU8o01pPjp6sMEH
nXTtVXILZB6FpJetA9ygDgDsIGBzwoW4q/e2QtCTbLD4Bj80MY5YQsPqQ3cM4+To
l9KcuWvSIoEk6ly6O8SKQihb97hcOSH1K9CU+4fCeElppnRiCGdIJBhq4xSXjLPN
1tpAVTz5teb3DuzqlomSz4DqeSEBTRsOvf8edByZzARbI0Yq70Tc18rdZDhUgdpJ
fewP5I1/dHKRnlrWnxMVYhshw1kxL1Ja8ijwEq9Z0cJ0axX8ClwxYT3N/hxfLjAc
thGMVYThnJfX9Har1B+UypMvU5bdxvPAWTJi0+IQAlFrKJpXqhaPLjEtvBeeX1e9
4goYIBVFlsiWLc8P9H3zQLzi2iPylE2SV1QPlHaOLx8hNeJa7Rs6DJHGopHl/Om3
hqrOog0ga+yPLlrYSacJaoV72xAp3vNLptLirxdu4lrFvAcfl+DRQnyGNMPJrTLd
t/jfXFeWvziQqj1YmOsVtogJDd/0aSkWsExZq11skeuQNF+cf5tKsB+HAX77UuLG
/b2742tmK9LfyD4IFuSAbAERbdERPyUJzoiBITDSDvBxXfc1PBJXu7oHQfbk3+aL
j0X2+D17A9IZnUpSBZtjW36lS2gw9cmVOQJ0ZyMGx16MEoPFfUsw8Br2r43XxDqV
E5VqyUUtnGc6QkTclyWTY1OK87c4fvL/lIb+CpsI4LT1MqXw04UmwfFfLAVHzQeO
Q3UhgPl+jUXaq3HcSMH2mruSOUQELbHirM/yxWL5rpufd0afT9WYh8lZLIonfc0r
NDqFIjm+Tl6pQBMvApiXXTXtHTYp5yIvWICQsbwOXa167REQoxmd1dmYPhkY0Xut
ZPAy7k24gcm8upN4PrSoyRnMEIqUIHrulChOa4/z27+BZ1XDzbN5iIH/f2YfTDb3
YL5jng7RzcbdGO/UEetbq8BGBMo9u8Y939GiKfN0QaDbWc5JnU9+OHrIcHa02tcO
CPLgLdbRMjYCzjfoDHRQrfgZQOH3DtbdS32H86Yr9+EuVwoYYCFCJA7vgTdr6qjd
3tAvfiVG0J/pSDMTezxiENPiy0n8bLFvnOWdi+wgtOlOZsGGyQ8vw/J+Z6ZAH2Ok
Rs/u+kgYTm0878eEZyvIZ1kI3Yb+qW94RzZodjQJM+jgwKExqUNAnGJiv+ZrhWc1
6TTtcdbhQeVCsxDGVPmIU5uj2k8+Q18FWywKnvwv0UZ4hZl3rQxmCASz33IKovZv
9CUd3jE6e9p1EBaiqI/GuVzy7LZemENTesG0zWhVf28D4VWhJToafoXVuZm6fpWl
vO9XBVs4Jp3lo76Jt6ivbivzL9d2kG8OjzgyPxjzfUDkhPaRSuVW9CBLzZ+QMMzX
0+sxzzCwiStxURmg2ZbLXmU3dSA/elRL37eP3WAwQlEkwNqtX73Q5gEguasky077
QiRe1E7Y+BsgMcMcc9RR0fpAnIY+0WyZL2/NM18gUlegwOIRNUUMlqp5FoxtSCRG
Kh9Byc3kXjRp96qzLB8LSjFh72KRKaN96wZzx2Fh0Vb9d7kkH+iUyiLT3BGmsAh3
QDLJVdy12KBiILdraqLqiCgD28h4qCLrm53FbGdz5WIiIRSnNDIxOC5sVU164tJa
MzaXrNKZeoC9512UBHLr8TzajFQvF4hr6OEgu0ckQI/+5ds5QzkSXqzb3VaSlQbz
HBQWwohDEbbLs3YXolt0VRnVbq3VEcc3abJYxBLMxkNuJSgdZ8VpsekTlKYND6NC
LdKJTmNdxqgHk4d6TD7H3Z+C3/d1dtTpisL3wzmsJXcBztolytamMdJwJlMnS3Av
6RgK9JTRreYinXpMGb+jAbrcX9ZXXZmsKcsQNkq9eoro+Vv+AzFXepbHW5e1pJTY
7WzcuiuiBshSZNYtCcXcFTmWDUdCQ5/1p1FKxiUfMLR8FrMo9FWW8hMpACxVNKyJ
cGQln+lrqGm6Aj1d972TCAYffqKcOFdM+BCAeJzpfOYN5NkesFNkAwkqRmvBsf4I
Ot97dXxtJ0WTI7+QGJP5gU/zdI/tqp+suSUpWhkd+fH8ZajUvnw3pYZaCCct+gvb
jl8Cp0zI81JIJadzLp04UM8eyEH3WVUX8HwQ2/9p9w+LCtehk5F4HOj+qjRYNVoX
+c2x3YyBodDIDcDSluGT0noIYSVjVnus/SzsXwtHjED4s5aGM0UTHgoUyvZ8FRyh
bUJMDXgZTjWyHx9KVT/TYviAslqmwwNhCkFMdqZduqksWw9J6Jjlq4g3CVEDtyrY
MPG4fffB2jzUOSalyD/A1JQUA/fdvG7QbAVPbtwjujFUo8Kzj/CIE4i1F9GM3plJ
p4STTVvRrla4pYzXZGSt3SR6Rjj9plORq5F3YJry2QjUXsHA1BVQmiHpZmaTR+0O
8IoMowuP3XbJDsIc+cu8IJCj2RA6msRQ6wGn+pTRAqUmDgBbcUlL243BBRP7q75N
kx5D5sp2RJyzcZAdC098HA87PKEAlTg5g1OB96sydmT7BZ19txyQwV2aQPqlN6QL
GabH0UIwm/W5hefcAbFpxEXzORxORwIDh1NfxMON/2qHOs2sWTzKSbfRn6NSEOru
pBvDNDxvh/hY+q9+sJjYS0o9B0uCMuLepGe6FoyAz6a1ppPYpKqgMGDdZkmbDD/A
+s8G0+paw4qRNCcMVNBaSpzH9324Z2JszTynTufHH7Y5hq4fmc0QCG751NdClGBy
gSLmGe8YoZSSzjqh3ta8NYg4dE9im57JNjXhFSSEvjUJ7ThDeXp6aVhz3F5rI3Vt
E4mb+J7PMbjaebkpE5OtcpnaftyU7vUZuLSYJawvA2bt06M0Q28w4jj+ykwj2tdH
kENOHyKskwf+D3MqJQC9Uz3Ox+aC9E+rc4fvFItDiVjVIaxRZcYdCOIBij6f9+Cv
M1/GoJbPsnWYK/1hTYix6I1/qVXvbECbPNy6pJtL/JfrZmYem8MSoM/WJxEd91uX
iTSIli+m3Y5MMLLbuRe3dQqfAUf4TnCAq8FBvbeatPjO7p2AohCdSruZfv6bEGa6
3zNGik/MiPbhDlcY9ZwTmxVSfaGPOq3iH5fgkmYUyoM+ThVpOBJ2uZqikDBiZLzC
yWFRzQiYFW60W1w2jtZksS+ms6pzbaDIUWSbP5YVgfsX+GuanOwhRUDLE+yD24T9
IXHNUbuxucpipCG/6cBH90TV431/g4YaTy6kTnQ41bl0edRErfHNi20aM5Q4eigS
4zGRAvv5ZgkRXFR2NtS3Ak9uic2XlzL2slRlRrPmROVHUhbiDeFeoS9wkCQkblA8
9DApdez3jG9WeuVrJZQj8C/I+ZSR22Y+UbYN/eO5p2DoVKzCWYfafJgP1tEKGiSr
kY8l21zP9h3GlE2795brhpz5X5HC8pP3L17/AWk3nByx7LdXjJrdQRAYIQ45hppE
q+5h8dL/NbsSp815vztSzh8gl+J7gxYIxaD6uGh6tMVlPw2+iRDYzFgbXxA6eizW
xumKF9vdnYII1FFAi89xbaXRd/Ce8dXIfbgbeNw67GDaS6Kx8vPohTl2Jr7klWKG
iZ3B//Xg9LKatIao7MJ4rQqql3cMJcnbbSP+LUiUirxQzxQKftquGd+ct9JHmBOj
8WZWkerp78eymR7IreCcJnplYV6umcui1Z/fItwdIrRLx+VVZn9XmMKZesZDRymU
BJ3XXbIMF82TAIAPNQ/DbIBTFVssfI4ccaiYWAxCF+CmWXbKHVTh0yhRdqAUfmBQ
MhYItRJC96b37B43aE7cNJpdlP8hh5hwDThaP5PrK+HRPgj2xKdU7Peb9Yxi2dNA
GxJtiON8cxKpWDGcwnX1zFoq2mCIEolVOP9QdVrL+BCq8MdE9PS/UHVI9MKUg2wg
WUpPMiCobzQlODIko0kDzU6ONAmISAjQF3RRD7YaOmBUydG/v/bGueNkPTxClXpu
KDOQZSaYAA47eML4B1I6RcrRGOGg6U8bt7LXUATesZYG5w3J9g9t7vDJru1J1ylY
DiVWR4vJMvLXRx5H3rYYLFX4h8k7Vblqmg5wY8JIm1063/nOVYo3Qwc+E2MfpcVI
BP4cFAAi2U40K5G3mqBhL5AB0mhcIlamESHL6DxbQqQPFHODx/IbRm5pj3vGJq4k
QMlvcGr8oU9AaRB574oQ6szfwlB2Pxkq4RP7FG/XBw1EwN8Hv953njOjIM6sOhFV
gEw+osDTSuTrQSP1kIFbIl/4KhDCCZs5K3R6MRltI/W7veuTXQeu0ZxmmEfYUq67
bRDlyKLbp+lAMlGN68KmG7/cRqoea3VYixyR9Qfj+6zuHvaWozZJDHCdG9paCVm+
Z68DzcX9B/Vnfvk9oecUpYILx3Q09Qbf/9ow9TAr5sgS0tDqIlgZNrSjcfMttAoS
RVGg3eLdPuXA8AgfirQpbA4APZiixfbhkYQodhRhBQDKuD4j54VwMFBqjNc3PAf0
rk8bUSC0LvKDqIo4fwoTzt5QCsbXmBxJ8x1H6lH0xt140caFBo+hdjsh0ZVLQJvP
OGdGw9vnbnRtWPrZN2BvLSst5N22xDcHGu9Zx7G9lDfzpLdF17pBGacNIWmKLiVE
XPKtl/jpkmNjLSW/9Mg0o96LUO/qUlgAiLz4E3uXxU/j/LtXhDIGS+nfmzK9njoO
Or8d1iE0fckbv0CUZud4b2c70hsoNDE1RlIAJIUswsnlgCmGa9fITYqvk5qkJoAN
i7EV3sc19eQIWFtsTx/AryeCOIzwTrX2gaKM1X3+PmzJpmOM9BXORHfDuq6KMBb5
QgoVzYZCW2jex1xcbzgfD3l2BiPWEQNUpCjaF4Nba0SqW+l2nbE9XSVV7bcBQURd
GZuqfHlW01qyPZpiAo+RNYzylqx/84z7MODuSqLXAH5/Rx+WCjIDCHWYAKC+i96t
kBDttatl8BTyc1QgOf+Sv4Rsajgc7GAuhig4jX9VgZG3MgtqqgRsxaRMmirAjhWa
nsKpQre2EIE8riLxTTyRHOlj7oA19otFt6ALGzIfyL8PRvQN+71dj6MUzamg6NEN
HUe/uWq0xLzXCIxjJEvL9FE3E5uI80VITthRm8EUt972oM33PRoY4XUvTwQAkVKg
XZbTsP+HHHm9uNhxNSxprgxkvWVO6FPGAOctbAA6rnxBZ+/IVXWS2DgOYhzlU9S/
ZErwdGcEeRwyQNTKF3CY6j4imsxmI650bL4YwzjnBDyxpoumhZkVAtpVpfVEzwqI
iMgKvd9CmajU1Em20Keur6TsQCfVm3cO7uYKI3C7IBtx/fXBsw47JgCZQdTGqUAe
6E4fp/1u5kdJUTlP4sOynaitB3P4Qk0rMbU8SYMCihrBBLOxBQJthnUaRcqRkGa6
qqVbmJmagqhHKHMQplGUObYBjE22cx8g0zqUclIAqRtoYrtxVHgwPEYZ0FBZp7H3
KGJCGG06DU8+NAYXQOkAOLF6wq2dXEenpfkL+fqkiqCzIBhbWNVzyt0I+1fxCOTI
WCKuuB/qKdObTIcNUL0PmHfEVuztjQuR6weRnms1EvlVoSXEk1MkOYr7+NHtLyAi
K+JweIs2K6lBAnjmIAbbczd2MOO6JhxPSJGaidnxIJXLNcW5jWddmY9x34veccu0
bpnbTCtQMsCGEyzJa/rf2MpA5YNw8V0PwliyKZ6zng8c4tcX4ARxvhz7jBIccygy
rloBMmxSOEBnk9e6yIJkx1V2oTR3P3MteuJ9idWCDT/q5vSxuVjjUCp1+H2aZjOq
wUo2tyQNfX2ew6nfb76VcaAdiqbAW77kj8memeiTLbr8fLHpFCAAwpK6hJZFupAd
9ahrz5R2yzu8akHob0QCezsL2PC+cMp6fW7/5+jx4XzMUihFuzstfZ9LPpA+jXYq
EPG/J9xgfnGuFYXxR5d2zj88DGrQ224kmH7aPx2rRLvukoOMnCHbS1l55QT7Rc0S
4PEXHntypk5IetfHLIARobwqVnNWowaxck5dCJFDsC19rjuDKMEA/YHbiN52ZFXU
GBp6ihta6bKs6x58kIqKegMBaUjBcPwbqAC3t0+kEDkW4wy+hutOd4H4nr4xpsKk
DUqB+fcI5PlDNCaEXQg4vh1z/4qlYXKVkGNgjBX48n4yEDiMBeOmh4JnY1CJreFG
aw/9yBcEyftRsmQc0XUG7R9KJ5hknrKFU9+wq4+KmoqBhAm+KRvuFIKkdHE4GFa4
u0+redWiGSUfhLM91oMewfkpA13CZ/ehi2YUdp6ffJNTtQLgy9SIho91pX/GSWMK
ar/N6Xwwjs8qZpaMUhuabOVdc2Bww+zJpRzCj8RhA2Wek0rED2+vmRby3JMZfb4C
HW7YKP/lSSNxPzf6um7/nDrgLhRboFJ6igQKRZAzrR/oFqay0SPQ5M89VTcIxsLZ
ibWxARAmFqla8rlNeugESnq8l9uY2q45TbFkcZmBTDKeRFi0EbTlJPMbQl3XVJrs
HZyjAL7df11hQDUWAXcQlBIpenA4m5AkX2kh1SdupLgbiFQZOXH/kJxp52uwsF03
IQ2bt41H8wh53Hp1OltHvbyQjG6NVikHFNQV83az986pSmHT+TXC12qR2lJGFWkW
V6NUywp+cHeC0auRAZFaoT/NBroENOwA1/k5TTbapyunLWHD8Jk/v4oF4NtfetjO
Mal7yZ81tcs0cf0wNvOUjL5d+063vD/gPW1OX7B2LhTHkD3Ubxv6bRt/aZvyoeEh
i5cDjOa1JMm+d4RuYGvdBTX9Fsr0UciSlaT3/X269cwlWbOtE0sqYqxJXiK1eN7B
RA+llxBUhnpuxc4hdEPr87OYXuQdyQDo3LET1IgnwpGIptr6h0kK1267ZpRRtnYk
4WBdug5kfMsW54XzKLRwLXVcA7NuH+1B5YnjLSsihtXt9HtWwaylDWjdj5smzAWU
zyndOdgrvzRc+bIs2V6CRvMeNP3NCNOdmzNq2V5tJh8/mbnTwpSjwA2iVLVlyZza
aS8/HO835HCDug/DmvOVjHS90vLvsy4jax0bmI9ozelO6Z4TwTkXSJvfTld+Gmfy
tsfcovcUWOCKQ80QSvohKbyrqHmHr0MnJq2OE5kLnWj/pcn/PR/8a8qctAkGez+Q
s2FNl4af2yPsj2eGo4o0r7hWbP3NlhN54ncjG6PsEHwTOF68ZF2ELzgDdBL57Jx3
WDhcVLE3yRACRqGrJYLrplyk7oso6HIP3OzGUlU/ThCqxprxF8P8C8WJ4jMPFzaR
dsb0TVgkLpaycGksPaq+CUX0PK3ZkxVbEXtXfFiOZoQvCnAKI3AytG11hzgJ1AAI
oR9snXdYEu5V7o0vdApdIyrSewk3sUr2Pk5oTCR3ZY8DlBwnMDFBgRKlb36w7eRo
f7n6TWTM58632qjL7Q8UewOGDnNbfSBG3ELdPGW1eagPFzFm2c79yNcyucvmCeWI
TQr468IKuKXdnCbcMmnMksnaXw+JcNqFYeg8/QX3HU7SXU9siUvwVZYZIXdlrldB
3EuAX0nE7EuQ/z0qxveyJfQnHv4KVzHnHhfY4TECR0ikxmPHkhUyC8zlx8tK2v9B
ii2Qc7Xi6+2I4mlBjKR56qrw8y5NPRnG6sePr9liZdyqT2aQAFbizLuTqh0ekJ0h
QflsY5q5Nd6+EeBrCKIzGkYHxE0fM7pudeVzr6uhLexEZtYPImRQVDSbPCMSVWWm
FNUZfYl1H+lmlHy2hB6WKGGO4aFOPA350yIJU+Hff/xOL4DDOZIqGP+RinwcR1FJ
xpSzRTk5XjlpSX+K0ngxj33POFmN66CniNK+57Fq497+ZzQogtHzXPA6QQZd1i9B
kU4xMaZpAGza3p54v5TQMrhctFfGnYzDZsuJG6+I6frUpjsBLO90bx0TfP9TELtw
zFyrij6+jvoKCC9wEkQum58MBTT1Ajgkg8rPAFu/F5/ffvhuAOM/fWo0ytRY6wAl
qxHAj1BZlE3/y6F1uZPLkiNW+7U3g7n51+Kx1qjXsvSzKMQqLXGEIPPgm7AFm/v9
zMA+Yss5D+OEwePVTX0DAm3EKoGsLSUvA9eKTLFvcDefqhwbo+6PoKgRSPCveIyj
G5A6EznKNj1FAojwHx1rTF5V8618QFvv590h1KGvdCJN5pC/RZ3QLApK+TWG84zz
5gXjBS4BGr8meLZS2vZoZLHr+WewVRG7P2Vhv3NRLHzgHYTECmXvr0E9YDp6J5w0
pb0R8w8tL14XLCuepSSTH4yLVu/odSw/T8MyodXjdLmXg4EOB79NJGdzSgPFvL4q
OCfPjRlI34+4tEYn1Mqqcw3crjFdA8AU6zJM9tVBGTVHbqYHrqU8xCYcpwyoPSbk
YTmVyr5xySA/DRP0Od8eoSR1JH5/hTKRzB8XERHulViFgFI8IqKkWjD44o6D+Rcu
snOzNlMGGgv4gFndYfqcFKdXeFEs0jaUwdN1+gtbQLEtzbwQWJ2PTMgnOAMpvuZ6
s5AughEPecwWr+UZSOizzn/6rFESQme2cou18JKR00xLCGo7ndoXiwmeY64ZRmCO
eUIuIEiQnGj476O5C//0EN1yVt1FR/Sf7xd5VvZ1qV8Tg4ZG9i0YRdr/wxVZIch4
12xuNb0b5ioLwMEmaI96Xdij1xJRbuwo1PqmL+RQumi/clwRhNgr4QvyiG1pLh4a
IXzPW6eALkTaCGlnHnh/s71voj0oq4rDbi3ZFRM2KCjsRkZ2/GefBuP2HzHNH8e4
I68Yle+J50wR4pf/IOgMBtwypwzzDR04AMVxrC2tujKxnXEgkKfCYKWWJqj0zZtL
3ts/eIf0Qrz2OeD9z7Al4iSXy85qtMVlQQ8sS5addBQx3Ue5nHKr1UMzNtlcxw/9
7qTVQYBnGp5sS6QWbQZhytuR/TPDNiZvm871gt392KDnhrxp+m+8BPtdi0ZTthPQ
9F/F5b2tlAtSD15idHHnTH/mhxn73I4rIcqNRPww37bgkB+tFWvHOA9dDf/P1rhF
bDdg9nPbNq9ynPOTpsIPGkaKCAMPFQnbmfkdVU/bIN0ossNmdDU+OUmmMenzVnex
uxd6W5lypFSzNGZkflqyzI8mQWS/zUVL3Ul9W3tSDsyV9gttkeAz09jYhevGPnes
Rdi4b5y8kFJ8VfvXijznwNM40IgvdduE6WXXzRWUWFNyN/tcleoXJT/bbC42E5Gh
RdP47gFT5e8njOhN3VYMIyY4ae/JDmE7LEQ6xOtEAe3OAKv3Cur1UNHa9vzi65vo
f4xsmua/HJ5SuUIWeYNd5bw3VPlgK8T4dE/keG+bvbwDVsxWX4s+EJakiu4uRh1d
wNRKdtIiMeGmp4iDXbYQK9KC6RiODXWrkQVw7bM1B1XgFfnnmUv5sTmL7L68Rc3O
EFW9oBqq45svbwj1wrx2tE2/CDKhjWOBSl2hyp9xLDFgH9aaTT84G+0KoVU/bZUE
mpGAcQ36oC4VlAgVWuRp4cSm3jbSDVg5at6RjzW9PPz+5LVDzhZShJwRiKk/tchN
yetlD/IZW/yJ635xQhR+singHI/A8MvkVNkOg5bBCN+4b/g3i0N72s1AuB8F6J9D
QavGmRqrVVbVosN4p5GgJGzLpAYgjwOlhCEH/nOQZDB6PWIvYTmteWxd0ZhlOPF7
BKkygHgmfPWPMv/aoraq6lCE+O3fnIXQczf79GWFqv7uQySeYAHM9uy92B0RbRJ5
4EtiyLvmMHcdw6rY5JNjUuo+Y9sfwocDjLX2ovyFWpeAdiSKwoqikjX95sby4UuQ
kcqG7MEhq32W05GOJEqA1NTV08iG1i5mVxNm4IpTW5wJQrQN1GAYHLFA5s31/E+B
H8CkDEXoAt0untPxkR9SzSbdzAVN9sP8viphLw1R011E6FrH1W1ypS0gK2ix+IF5
MlWdXUJ39eolQnuNCxYPnPcUI4/SxKnJ+K2jMD3jII+1kN6b14020qBWKz96BYs4
GUanOVt8paDnc8PKgNKyTPZvi0oris99M32g6Fjre0O053XbSip+o/oHQwK6X9vQ
J7NVBOEOSf1UkNIi0vEuf5L85O78I3/ra2e8jqb+MYG7zHFWSeW3TrMJzdRKOdik
xEoT8UgtkHSR2m04z7OIIifMxfeoBeGYie5GJTQwHE7MdNlKKJKSWNJRGe/D9OMW
4aMpT4uMigcgi0RvIPkE/vRR1V6ZyXCiBvCQBI9UyLvDz7k/QnMPKOh6uz3s5x7w
Jr3NaVBGMgDaHU5sUlc0F7DHZg9pQbtogwv4bRUM5Awa4KhQOMzlN4j5jv4iIXKZ
AhCCwcxUwqqDSSeWzgsV9c9g8u7TwTpr06UbTJM7l50NxHpor7FU2L7vjFO+/408
5DiB7Np7VdeskhmaTod0I8QWwDnVNgs3qnT5Nu9rXzUwuNoa3qKkGKu8Pn3cEk4n
MbsFhlEexA1ZxPaoOX6Sm3UQDyYZMSUsRuyEWpUoU+XRLEKzJ5rlAJf5jkgBM0PE
RCEx4IFsHVBIjaX9QQaHWF9I1tjWVafeV4I1d/9a102Asr0uW51QmFmrRN8DcAP6
mtg+TN+TvV7laCQQzdkoSkDXYkfmKKVMmDzSInuvty1BFSFW8a4WckVQH0hdtqom
DExol0/wspE9jY5PpbNsSPueTDNtH/TAlrcJ2fPS6iS+e2sSlpZ0cK38oTnUOpGD
1duKLmBH9pIzB2iuoYPw3lsd6BNvO/0PeF174tKe6GrqSEBvLXNuQQN1+0CzxijX
K9sJ31SvmPH0iN5afVZ5cuxwKW2WeCJMJaDBbwRP3TkOLgFz/hTMsU+HSxxHoIeQ
n1IR3JbvbrCEufm3bsh16n2pf+CfTT4gDW+p/cjVCCwtcWvql2sLqLyGzooDIpje
CqvU6L2Sq2j6eZ7jtgA4zVl6EuFgnQeqKHgrkmgn6jpNCOnNEMT7GjSHjZQjuWZh
tZC7urqm4odHXHDy9rRBwaO/JSIYFb1pSuw8a3Tkdob/ue2Hakgmd7hPTxE2/Hxn
KfuNxOkdJ28pqavnE/HoC5StTMmuXn8lq4cTrqpTbzH2OvRzlDv+6YCNUq9hU0Nl
wf1x9Zc6dIe6Fr+GNnH/2ZWPQFsHA64oRsGIHZHXWjqZeuueuOrac1q7Sor67g2b
nJK+EDFp1rFOvqOVXQfaqv9pPl8Hx6ZqICG53CFTM/mW7iNp8ulB9VJxOQnQ4M+s
O/pwBWHPOnZygbznxQJrTzMLdVSzvQ6uylt9wRXv6Lhb7OUBdZXX0cTZdY/neaSf
I58/gh0UX2pcCGo9ZQ42xBDDmWSY96ydrpFPZETu04Fj+EvQGpCEm0mW8eJ2ShHv
jcV18EcTjYJKiM5aaaDKcCRtG+mA+adxt8NetUPcZ6WdoJVbnPeUMYKfMt1ij4GG
yCly169Uh0ZqfekFuN0bHFCGtI3AM80/b0Lu0lkC9aFM6IodNgirnhgf6PRqxfbH
fRUrpsDSmbdOWjYzSwSp1kYpi5KoVQ5zgKzyKm2B0fhbiYp4ZldYYAG45sLyF5o0
4yYu8HP95iuMu7n9a/2lqNLfwwVLM/eqEscRfUo//VDx71cxFqUPq/V879l9KSBc
hS/Rpd6j5mxpdwSpNX3LXYO5Xno2SQnvZT4o+1/hpeuwfBw3pEHWqQfj1o+vBJiV
NS1ltG44OZswbLQ4Uy2ApeBoLW09+d+pCbDppzkAtDqGxh4ECim3t6Csx++P/ciT
wsZMcXOCf5amvkKcyRpBC/6W0u6wWZS8FyM+mdtJqguHSoL6fv0C59lHOp+cU/tt
UCGM24+pPnQfD7WpVKaEGJmt2YaA3V/lodmKTo2tvRh5/xbGxPKHWjWeM5mBUSvM
9ya3TQgHlkpBgcqeZ7j6Rp1Y5e4xHIJyg8HtE4HZesVKIh1VUCCDUlyBLM6daBMl
wzpe9WkP3UwDCvmY1IcsWIorOeOHQ6LPXyEUqHllkwTtJ87tPdVdi7z5zXiVQOmx
pKkYleNRKtj2NqjN4mqiCTLQb9ymjAyRzrufbpBLDiWnOY5T7tz01MXJOtGdRk9c
dcUDt1cstjKota4yw5ngKuXfjixFYjfEIPt8MheUUsapvsgtcaNc59zQTVKG/iqq
74byNUdd2uHNeuVEQYf3qrxK5qBPUqq62crhj1CaSsmmIUwYhdpj0YRiY89ZXPq8
/7TtHA2FJa05TPkhq6K23TS6iwhxa88UsYhpSZQgjZ1DyadxFdOulbqc4NywiXWe
Urz2rIC23sKE4xXufAOPcN9Mxoc/gGmr8Kb9K7MDL5Yy+Lm+Vofn11rzPxlxsqWI
K/MY6Mp9SQY/2lAI26wuVdk8cw/3bYu5zAeopGFEitrC4TYl6uZAq9oRI+v9VtKS
E/6JIceoJI3wDyevdqZqtZDcSv4q8gL+Ym0eEYigZFsCfmsuBEiGHUjxAEq1SNoM
9xEpijYQHmcdgkOj+ot2hs3XZqfLSoPQ57Om+sJ2UGh81+betvNRC06b2RzPzzoS
cgnWt2ObLTjHfyQAoQyQ5h14juHK7rdegnHEZGyX+c1ww3qgkRgncwQklO2tmOWn
dw8JmhHuoComlB3CfJQj/lesoj2RVOArfkMSaSn5bWr6H/zwqR2blcnpG6N966ji
275ryg0/JkO+ugnZa3xTRbHEUw9IXEHXmqJJSKJj/SYw2PW7A6LTYvdUohHi7hKp
a7bEyvh5sk4KAi635wZS2BdI+UrDV/zUcBYF4qYm5mNBccATAXX4soUAYO6afY9A
eYsAvG3fkZIDL+1v4k3iUlS/H5cyrr6GzVWZRlyBA8Vpz0LxP0vigw2a4Uy5pwhd
3k5tyXmR2VqlBLml3vdlaLQP7sFIYHIr5jAbaBNxVF1JySAQgJLWGCXRJlRbcziz
yBRvA+dj/KyaX6xVBUdJfH7Fmr36QjUOzGPNgpLrtu0JtjYt6vTWcwreJYnaizQb
cg88YfAM37W3mdJGkOhFx4t8il36w2cpJ3C8wTARIL4bn5MNHA1XDJPpVvoHItJ7
k7Uyv9vt+6jTIOtNdtbPAAZbbV62clk4iIWYezz6I4yLUm0zSMbyfcWB3dmhpfsU
HQ30Nx0z90nRkMPqEBhOJ0SN+MlZbNrEm3sF5u/BUCnTpNftE/QzmYFHWMitCCtZ
jhqQAZaMRbmMMJjwdcpN9lD03B6RQ06f5x7p90rENi8oamnbPRjbY94JVGb8T9Fn
B/Z12FLLNsOdrlXDk5S44MaM9Fpz47rRV12QHmdO/QuO8n3FvrhR4ZQM/PSQIgnk
0PknDK3dhmRXXM5dtIgOVEVuZv/rz4VtSu5w4c/LDUPsg/+ctN7Kz/XQbBeSfn+i
x0MASkfMcGoKFvydJN/JDi98Fdcns0xstW0/ogiJtYwoHk/I/JcMeVREKzb7dPqW
uA050HJkKnkeQpm49Xo14+BTkNZ1smk6vLwcd0ZFrl16mGLEgSDZkqNEYwvodZ2/
HcOfQ34oxkHOluZixMQpVFIoSV+mpbyPMNrZxbDFOxNAik7EwhiyNSG8d0ciDjAi
SQ3Qw/d88QJMx5dRoclSA5Tgizidje8Izbxzy9/0LweSki94GgngOoHCYrVcCo4I
D1vYtsp0O2sbrMx9M0/sY5tp3QyAm8YEJ19uvY+ZctvzIQWiUAzYsZvBvo6Opvbf
lIoDRUhtmrvGdBIUX4U8BHhRWYpGl+8Ky0fkV3Mp3fuIk4DZuSn5k13HBhj4GH1t
GaFN39mAdGUxYu9xuHoUhGMVP4U7lP7Gzgo2yyPnq6GATCnZ01EpndY0SEwe8Rdf
amd6rJC8rAt9EdIS5qo6IBGugghlLwZllh/V1Utfa/Rlyxuzvw4KZwF+CZLisQWH
NPCHOVbFgB12V23k0qIcHqhI1XbYknIydIcO/WE96JNMLtdATs1HQm1OS/NIDmyj
dUt65cbHoBr207Ajr1Uqbg7i4EcHt+dPISi1otGDW8MZ1p3QbmWauPhDpri32Ahw
T3b27+WR3QeKWoVwX5Tvm4WzK9/id+vPVgYsKhAaY5E9TFNSNicdxlk6I/bA4PXg
Ci/wXrOixQiH1nf+sVUUQRvHvHyaY8/o2+gBepYrXw36R6ZlNhIjdhtSY3sQgRXq
MS1wwxdJqzIJ07Jc18hd279jUqXcfwA/PICsGPkURFubFCS1e+v4QcJmCFbDI6sT
D6jq0MpGV20SBWKvPOpCIQDoBshfbC2/yQUKEI2/hsXjzXhU+GAyAOJ4RNywixiO
NjNpwZb1gFr45qyqKGU9GoAheLfLxOGgF5xn/AG795DfVWKy16ILnZrhwLWLqXa7
B73cQP5ERTi+ZU8MXcbG3qUd7x4kdAPz/wRh7HXkgyfMyAiwCj/F9LngNIwOHkmU
OCedd2V/KCuGS45IlHTKSKItaljLkHjkhY6QVV5/A+1WwKd1AdRmIoppjcVg/BBQ
zIX1f/ZnafaUZKwa4X3av+qiRY8/NtzALkcVTssNffsirGi26UmjRrk0AxKTmZdM
c1Syhir4kKyt4oKieXfICFbLMwrVz90wF6QyWT7zAgifr6bLmJoqZpJMogemwocp
sImoBmlukPi8qLfUSD0BXWxgrOlJ1G/C5vrXSUFbs+mH96Bp1vAohchWBaSKv5mO
Ftm5/JwL+yVc+ozSyP7ERUlBQlfshoHzqCN28BHKBDgU7j9FTpVBOkA1hPEgv9Qh
Jo9ZqZTma/R4b0WKjdM9juRI6IY6wvpH/PxLmhd7CAIe1gGTh5YsdzLTjx/Hbn1d
Wn3PSC8yBwm0jl/fUQW+MN303VsEjngypfd+JPXLGUQS6TerdkrpZvJJi/z8xdfi
fvdIhqTMyZDXIqPgoXsfZykiJOsViU8crEWomhonIJ9tiLzh7/OKvzJk2X/4wwij
xfl4syNgbzcqeYKjo3tDtNpjNaBpUIqekP3OvBG6HEtU3Nj4MoUwQDKXaL8NkIVc
Z8Ai9n/6tmyM7bd6c+4YfJLjPxrtSUTFtZpQeMTl/MqsE8iWxN2zty86lVTyRu5r
SPq1ohzZJczZ0bhzHR5nu6YN4Ybf/CArnsNkj1Q1YvcK5j+JP9zCZm4k6Tnjcj8j
K88puxYRZtLdTPNonSjWzjW5DFzaDO+QNtjZswnGh0HY30P5zB784IN/j1LBtA2X
TgsIBCIwKBkYFn8nZwvcVBwukWm5ph8PSOs6cOfToQjYDztmiOKv4cLN2olyR5P4
oA5Y6nz9t8NxSIYVzqybk2tx96iDYGCo9eneHNSllVmeJ00VCs5ivWc5PY1ZpRj3
OM11Oxi+hBt4OV99R+PMxadaWiAsb0yHFWg5nkGAv89r3PoR4QU65uJUWdz8l0A7
eIjb4hhVhnFf6CUSv6RCR2cLz1xVaR/wDzmxAU1SZWdIZ5BCkoLjtCK1m/Z+xoCT
ak+ZhA5X4OAhcqUFVMwdyG1GfGad7LgkKtgNhzOdYFKNlNkqrIYRXZ+L9T3pKaaP
vbGMFwEzSEUme/SixuiHXQ03c4b1YbPeLu5mhbO3fgSYgfCSzMU1Vs1xTe4GqEuT
L3evg0Y42VUSD9HpVm3+Uhj555CDptJPpsQAPihAYY7gZsL76bY2/yWTp23VrF/1
0OcKxRB8vOIWmDOZ8jmko9SqsEKzwDVWr+KhEkFJ6XrkhpK1x5PWfcYYyBhQEk2N
yFpqMOXfvO/Ki0DXYe6lT7ViI1Y9wYhZ2HXM8dlsgJQ43tgcO5AaWlqSxzywsNFC
f6tIHbtXiHONP59wSpZlsuDBxQfvibT8PgzqBcPp/IQpLdCZlkoq3+LMFOC9+U8F
yfhZvr4np3ADreyK9XwpgJIobyncPaFWu3XzjVSxoEUisZswXtIwC21ILq9Fvqbp
wO3aFdXdYHZ7InXt1G8Gf5ifU5sqb51t3LLrCksgavTEWoj4/tr/ZQhURj7hNris
H47hpbag1mdRZke9ug8qq9EiQmf6qJIRrGTJ/2DZueJiV4suXVb0DZ8ubob98hK8
1glqukcd57BTr2LGkyc7vj5grn3Aur6vJtCwXu3q1+vReb6lp7gw9qr2vv0hXYdc
jvCsF2KV1H/n3j1wW6aR4mqcQolIyvV60r1+K/TqFpFZbu7vp4UMSSEexlQEcPz7
tXCeEKlbsIMO0mWWTUJLC7kT/hWp0Puwz2awY+6k1A9Yj7hzSQwnbTqHp91nIHRq
6EIT+cX8Va71dPU4AdmI39PGIZA30m1oDnBql51H2q/bI72C3avZvQELtRAJlOc7
miJ4nTdp7Gwe3DvPyRO3Ee7iSU+Bsko0vYc+BnJg+myDl7mGbEpatgAt6HHZbwVQ
a4G1XDb0MlztaONFQRZxQcUsx72QABh0eCNV+NoE60WBOsIi6r9uzrnHvKULXBku
4WHE+PSzIvosJdWAusYxg3BNnBl6j/Rz8B0kMdujgnRTLJZ3yqiphZGho2l+bey7
1ULdKbMYPRjwq4gQn39FzY30GpSlmm2Qb6BDw4soISBWZmqi7FzZK534LF9o6zwe
uLjxWe24mHiZIDg0hO8J3UBbfxMIYIPFXmoFLehvmmziU8kEuxrv2SC3jDdCBG+F
KlkX0qOXUE8SOO8IQ2odpjoxtgAP2HbNPaMVCyMdmwtXV33251d6pewoZYaKzcEu
y0MRsS/43ETReWYWvVn6N4S7DBSV9M9Wh+s/n44mhZSQYNjI77wtuJZmQQXMP10o
AzYaEdQ1OIBch31HiRTfXbsT6E2p2B6kSC/ABIEvkdPrUGQtkXBn/poWq/4kWAnh
zZoHNvxGDG0PiIcaoWZXdyiqUjhfZGEugMsvmBp1QkAeWsU5BDCCVtLZV067hb0K
+UruCSfv/x7kwWWu5zZbJpYevcb60BBJrzELKx4ZY2UW+9YnLTkmlmsIoaLoePhK
7MNGJuEQxVzATeu54ngxD3iBe85xyI/RSE3zEUNZwhngkvk9uV7I0nIT5aEmkvW6
vydlI8hifn+eJRpmFs0WbVTf8PLPVpUOFplE+jQoDj/TJ84Qps74p2wjdfTXa6mo
k+OTc2s9W6cHR6M0L27FR+QfrwwNR4A7U9kqwaSG5viGJsFXEgRpn/XygaIxCfZ8
lAV/vruBqWPuscT3l6AE2hOyf1qKj9W9SkE3BOQB1jUvqC/WXS/9VIahgkIK8wKe
DKwFa4s5W/SG/j0nQMghDPXS7TrLrVUoefl+Lh5giGWfWh7Y25deERPp7o+yFnbO
VHcEAPKRp6GdHPwCK4KoFwvovubQ5Szneqh0FxCKUwagu9qcb+g9M2HwDXTQzJCw
64a2x7HMd2e/bF+hCfNKNNHjMbBd2pSMcp3udgA8rZc/+oYDPRBWRC/zpB0dgQvd
wVtWKoo1hm0aKEDwvvH1PTA/unffCm5w9N1DftiBEFqrIK1CZqTZp1tdyodsEsNj
QnwzyBaBfP0IwElaCyKmubA5ns6mGQ0ubSpdaFux7q13YLdBP9aUqLXQxRmwqO69
L7qAdrJqX9vb8kD/SvLiQp59twbyDYHzcVD3h2Q5ghtkscaRXYYoy4G1tCfqbJGD
m4IUaKMKkv0EHlQG9plYDey+nvpjSs+ZSPd+Y/hqEEv4DwiofB0Ql1UKJRvC4kVm
H1LnF6MMZsDHZIbPaipoJce6HEdxSXau14Us+dE0ezqCJwsL0IGQhHjt5Zhy/Tlc
vtLhIE+BWskK8QsOnFS88rUy8eGeX1fSeQW7j3VlZfA2+oJFEih2lSkB91muEfAP
dxoqvuIK01Padneo4qRPTLsFgNqHp27SYmiLxV+sbHW6sLcTaLcI0nvcmWHmSlzK
yoABBPQjBIEQ99hkjdhbgYkot7SPnFYX/d1Y6uXtYH/29cU2irLVWyfPdxikJfOs
ZWvSpuQfLh3A1D7LawPjuZHnflTQm9s8I1L/5yuo6UJGwmw8iHahbPb2vsvjuf+T
xT13R9JZ8uoindYzrdtjLXuLA3qownAhHGGWGJLyYdxkyGt+aaXxDmklRM5hJA51
cO4WU9yODfVUwEU3j9TmRvJC+PIMmTTTk3iBEvahfeMrG8F8zKN569jokUeMeQU1
qBQwpA5Bqct61WTE3Spf3AT5V2oZarH+WMwnrngi8g8D6HnQ7Pjpx08nhTHQEvd6
MH0EB8ttd1bPruOsr0+XKQnwztzpwa8Rg+iEk6nB+0TcIUNBwZTSuCcB4/62Hi2v
DSYdAWnXxnqy3HPrd6Ta5JFqMnos519DX3hS1dVc8i5Rh4S+/E7NDbYQfwC0LZ3J
jruvezcc2XiVmNyZTRod1pt21aMwTfDlt0RobLD0Ab+DRaM1axw6MiA+wtej6ClG
uq9kaAQew8+iJSYcM0p8dUMcNWqP8i75i0MUwMHzpy8aMxUmFKJ6dP8hRaraRSgP
cACiifnkg8erx1HihGHzn6lbwjT/PN1qn4Pp+d9OuGgmwU+RdvRPNI8JUM+r1Bok
/RAIrYO/zJHLluoKUj41iWkYYtnZ5Pj7qCv9ZgtSOEjmyxjE7zpE8yPItDrEbrYP
/crPfpnMyWeOFBZ5JvalAgUdaEQ+EmOXzM4LTrwPlbQpaLLQDbRu0FSJ/LOvm//2
6eThNSVdlQ7cqXG9oVg92ktF0JJ7K1ooNRvZ8K8o900gu3/jNUF8pP2q3hohyfDq
jZ4jM6OZE44aUkeUm3Z3he7OoCTM5iPugroGQS2WsksdnJCpH0H5LJx55j5e0fzb
0eJstgP8h5VVnyufoWbJ9kv3kd27frMxVIbuI6BR1eoaZhMkhDKIs34lO9r31S/Q
lKeDz8B8Un/Dwuvg5arFOufUs3OpFzhxSQ4H3fnrGuNY9ZyWyOufT8IIIArZl2Xp
SkxfwDeXpOgl2QvYwuLy3cMxdDQCqC1FPcRbJJTeXgWRLykZ14XzaAv4Mu1D3QN2
eDBlWvFwfQnWzkd8owZBpBJaOZX41wmOiImWMwPaawT/zLrNZBXSsfyt6FW5Pfwj
s/jDHX50KdZEma8nUH3sy3DkbBoGSIAKiVyIbL1mGf6rwSAQyHj0s67CUljzFYoa
slHqcXd1lnqfQbJbUThdRg1T2VlC9gGsXh5c1fNlnIYtcFuoa/WEoFQ7KPitolIb
sne0mG7FaN24CL+OM3BvxoFDsx+6Ruv4NJKZQf21WGdwqMsvMeByORIJe9njCkCh
JAKgigDwDYV3hcF23Qj1C0hEdH9R9ThpMx1KxUJ1RJDHcDID6A2x7kEByzFqWxq4
MO4OBhZBZ4w/GPInnHTwkJVBc2bjktUXvvljqryuaGJouvvhn98EOnq/zM+kmNU1
p3sKggdkVAa9oz63rzWXE6XsRNdsdCtarcTrxWK+lKePpg2GpEZSAcfwsoLoyxYr
dFEgsioejcD0YeluhEUZiDCvENBYLii7R/VzsFAQfYReV9SEDwufmIc2qGNr6bcT
78B+vffusIvKrglDm0b8VtGCMKA5Tv13E8pCknHJ+mNktC6FsWE9rRm3Gc8LaPX7
hVknxBQL+UxzUqYQhcakuhbfGz8qbTiZFD2uD7VgsuXvLebpqC9S3eaNgfKSgEXj
iah6Gp/LOFsYXxTunfQi0cOZYmnYffCPRzxAxllUPq7G2CvlOROiF5SSsOxXHJG2
k4gTh/ijESE2dNAilvJe3JxCTBrrcHgITaqNxzfjolj5JrtXEiCi1nI0WNADbyVS
hmqrXExZBjKmYosZmFyNQNPonTrSglodIGISgnfz+eR59daHf/HrfkJ084MqtP9u
HBRFYXbQOnzUgxBWWubFavaagjoJoQeByOiuKxG8T2BuIq7XBFZblGSqLA50SSk+
hEUrF7QPi9Fpv+ry4/J91dp4v4C8MCVFh83lP2m9z3Ur5qFH0halz2PMyHbaQbXW
FzMRiLKR1epSaVIS8umCXHR/0+lGm2UVBnh7aLoGnjkCHKGP/1TJhBnZWQulKlx7
80IBCDKrThQbhjMSCWfhZHWNnd/wEd0t0u3gGvugt2/W9plZ837E4+Bcm6iaj3nD
HGVEvFVaXzaTKsJ9I75NdMizNei1rMUnQVjQuKsA9UkgpIMYkZX4BF38kJ77ETwy
iwDes0RALMUjU7iOPsMf3dOy0rkreunF7o5QR12izlbmTSAJe3MBJR/7GacRJ+sR
20CrysvhKD1Ic4ONX21kZn+aQCmtZl7JGsEW6e+fIKDj8dFsW72bWHziT8cLukGu
I4fceE3uwY08LfvrqGecZc1NkLzHuoAF+5lLgpW626IE/xChLBGzxgUR4xzCWpnk
y8nOzOFFemt6dBc0W9kORjStnIu71KmKes5SxNleWPOZEOtKyYvGusRs6ofXLPJx
vRNDJC+i9ZIzozgL1w/x4k7jf/QlaVIRDYk/GsBLg3bYOGI7ic7DqAL+P6QvizFo
u+L+dvSM/zweKdA4VvNdJD4nmbP8Qj0hu8vyDG17rqg0F8WnrxhWUSMH1jrpWgCF
rLOEufelQU4rFkJ8Lv7r08zwGE7W6J66nv2JNwOeschH08goI12bowTqINR21l4q
c6bdPBjFN/r84r+VpuAAqxsuO36VUL1hZ+12vkHKoiHRo4p0EnxvfSxtn6/vzFtN
tAdfVReVeXtWtkPD+AfC2ynKQtnhIEwI8Cxk/yfY02bXkMwYhYIbaKQ+ngUOgw++
e80dLz4kLwL5sVylazO4wUxAYX5NBUr/vVrLArLx5O7brEHiZFO/5gXniDJUtKwP
5O6A+lEXIPPJo0rNK9QnzVSsB82j1RZeRxgsSaDaU2oqjSgQyNNRlvtW35+PcdEQ
OyCu3KQ6EimxTAhS/6IQ+pasJCKkIg87K9PwtwcQknVQJi51i7srL3wxzRg2/w8l
lnEBT2qQOVffnFe1ueOt0ebGvotp5ZGzzKyQ/V1UQ3r/NWuiBBDUb0xpTE65J1/+
LVTUml5TNb+jqA8gMoWSOybB4MF2Tg8ivRKG5fxWL1A/wcFZUVviZ8V2krpCLl9e
GlPbUxLUJDJQL2p3rX+g9i3oCb82kCVSX/hXURpNfdsDPLUjA0V1JGOq0EGcjQmG
x4PqTOcpiPM3pyeZGdisb16CA70asdkVVTMo9cdyjPev70GOmMMf8+OgYFUtNTLe
Tt8DUIGrfVDP1sQvI3WfGl+eAMHaVHwBHn3qTD3j4nGFoOYJ/0JsTQSQs5LJVsQc
ORX4JG42ZiWnjSsUW8NiNyJEcQEl0f0awAvPeA1Nyehp7hBrHfyFF4t9BWkZLbpA
aVStmiF2sEfW49HmFLYfP6BS6UMnyKCMZSyysg9ix1PCeDhaiCUDJwYEABtiKPLk
g+sa9bqtFvCBVrqIWiG3oBgHqwswIPP48+G6ziYz+susf1qC3DyOULSbrb9bYGwh
kxFZYfaPaQilz+O0AI4KjbUgZvNuLQB0eT6Kd0JEbsq5Gm3VmyxkQZ2pWCDSzzzF
nAIoKyuCpssg0nDYuCO5d9LClLU8ac3kVLRP43Ef/x4FxJZWMKOC+82JqtJ/1ZJK
XWN7OLJs6KHJ92XxdYKuhQOWoTRPUsxySPNt237yOtbSas2M9JQ+45TQChq7b4Si
djATJ1RccagWOYzUHWkFkchA+Q07U4LOcU/S0ruyGn48JCs0TXOb9HZ8Fe2bWEt6
KrQVTv4ZA6KKKV5JiQur7+Q1Wc67PYEX5TKCwqAATrHyw4iQ61XS1ZW5+M/Ab6j0
7HbpQ6MNzlp8XTLUpVnkF2N7PwzXZNH5HcBCOAKkY491lXnCIejhE/cPd3T2uH9r
5Z1Ilmqz8Mn4n2vTfAEoNKuUnnHXFiO3blTIrqvBvcWOFw+nFYzeybKshDcjS7L/
ILjszJFzb5aiIjq9lEuEw9LbWgTCwdQ1Tb7NBmUyTldzumx1Q2TlLwJkAxUKWML/
PYtQYkIqN18R0rSjFLa9p04rnwVVXIHW48HDAf442zPPEgBGV6ZNhiiczYqvLVJs
rrzmEcjjVAvD7GKXSdzg20fm8KJdCR9hkAYbeupfVDQLATRIsf5MAyEkHfOp38/v
ObktOdJiwNbrFFyHkOfFhO2YjE6/xRdrtA7d4smW0NRSrWjtpdAGXpiy+xmSMMT+
qWVh/5pXtbWBSCyGknPRr9Aj4tbYPvLXoLVrb3rcUi/oSpMiwYopnlszlmVWLttp
8WT2xNPdShAhC9dDXT2heQJJWamPe7En/4HvM33iwpZ30BmIckw6x2lXTXP3FYhU
7T1MEBHY2TIGHJYODfVM7cov7AJG/j6VcCliZE4K3l4tw0oEtQnaHPmIs66y2pHD
mMdWGZC4xwmMb3+mDivcY108PQ5wrYFmUOLcm4UI5kc9n2+jwZsVWP21BuiWOYhm
e+8AiQSQO3V0mz5eCZALh+QEx9HuXrCj/xybh+HxpbtXzET1f+eZ/ZWTXPsiV5mX
KRqRH8Dz87js0sYrB52UNf9M17prbeUqobiIZB4a5JDxp1ZUC8p40zUjhokyBNKv
NrxyGCfky9Pd+fB08zAsAHeEtv9GdIQoWgSelZV5hkVVQnTv3Uj0RD81TL9XAfsN
xpJrTZl22JH6jvFM/E8LXLMTkSw7ayJNmMuPMeKckNW+GmGNiPC/TdhNEcRajAxj
0mcjJVuNxpP8lhwtWRRZb2QnzjiY25uVVI3HMC0iZaD9Wx24AtCg3t9pjzp6uqt/
cwki2Dutp4Z2U2icqDwj4W+J3mHwlfSvFEqt7THN70sueYGw3kFVfvS5pELlW/xf
T14a5jd9PxFE/PW4xviW7rtzb/k65pxM2VtojSnpXSR6IGE1Sutg46huq45litfb
lxASxUJNUBlQVarSrYeRRINU7BMMYQM0alhMFWo3OFNIKvWRKtGQ3bdB6GXjzK7E
nyzMxptI1I3tMtR0Et+2JUKtuys0aSSViJnlPhZ3dtn4KDwKP3nB3VhGYUMm6Qm0
36Fqp8azWAfSGcH1vEU93Qki9FvTppngNr+yDFBNWARDuJNSoUj4565sbad4NBWl
qahy0lMLxJ1wgFm4yFpv6z03bJ/pT7LHWioKpTiBlo1Lxr9cXZ3lu612meqmWJ4O
8bMAol4NOaKEq8d1ixkz/u6eXouOxZf/Or7Od6Z/LwfsXIyb/+q3eUQd3DVCZxid
JiOReIj071j66H0NPdZkjt7Og5Ui6vzlkTK9MI6hyPWs9KhB/IcKJbx/de8Rl+Qt
10ToRitywpzNzIwBT/ny4NioGSZXC/72Mu6NaHGQmNSjigMQjMfqLWYg92j7nOnj
ZLpQ+sVU5cPujcDH6ywSg1A9RiGETHtskv1ZTfm9v/CVMZsTv4j2NJ07Rq0OGiAl
gZIUJHOp5xCH4JbKlALX2taOFAPUBUoZ3JCKKbbg/5dI625i+Ttt9OJ+SK3zr87l
W8tVINTq9k3UDwK5cK6GH01azbm71MPs1mTB/kduQPKJRx1aAL1Y9CvMC/OPlk1h
4xqU5i4WIkPi/l8CTXUgvu4m6MKlmPpwOK8NH0UaoN8tGhBea6Z/g0ZOpAQ/tWbp
euRqy6cgqVxSoAJDTZMQOt2aiO+fHJIZh8n9YP9lFkbgl2PmzJ0W7kKSWty6ZIY4
gfnveMtZCDXIpQHoUmndtPwVPrPKh8P5JAofrNyp3Q4ICH0Izc/rFnMctRA3Z+1j
YaIzEUOKGObBL2yhBLWt5HvRH4A5Oad1hfgq9+lWPuQpa+ZplXkM9UaG7agWapu7
rQM2rvfP08un0RPnxOFxa5nJ/RpwiRbjTvC9k8DS/eTvcfkKpFxknAZuiNMM2nej
Z593YnMT5sPxmQKcIZyvCfw7vcIYOkAUJVWYsfIZC67HTCDNKlGwgyApUnvKWMNQ
Q2M8MD0MhSw0BKTN926h78ZD8QwdTceJSqGXsxdxw4LTIetyL0brHO+e6JJKizsW
e3aWj558uQ34jbCCGrrI+y25gXMkZmE5YtLWsnzxnSSucsGhho5GHAVXqokPkrbh
jRjdSfA5AiL+D55EtcbI/V4YRlopPMzlbeiKt0m+EdvQ2NCYO3PmaOoo5KGTxEgj
M9QovuP8HHO8r8PfNw09hNfCr2tbPBEsU75cgxA9X6RYpT9VeTXUlC2zjWnNGkrP
Oh6eAKI811FT/PDBxA5N9S7Pp8wI80cEeptRe1sY/C74kJvAcUHm4yydsWTmxe4X
l5xrRA75cfgeRfIDguzbCZgksUhPoFDydLC6ZmZRQCxAN4QbCYuoq2VRFwstwZnb
B409kls16yFhBhhqbrd/W7rl+FEs7hX2eoGiyNq2dHibTttKdLd6uEEXEBflRDIc
tt9aSulf5/QJ9KHkc/LZLOw6pZy5yXqJhMvMmgEe0Joy8Zfd0dFvnD4bRjE3R+yo
Drm9gEd/1UgUAKIC6l92Vu4sMsQj8sq78+799qSQ1Sn7oUryGSim2MhfePO/YECF
HqyjV2Oem/DeL5d34BOrWWDsJ6SKLm39GrqJKC3yMYEHLlh+uH5Gb3JvLpIpZKtt
eNwkjLGiemuZkSwC+MGsqAOOy442u6BVflDzmJIG9VbyQVlYt/elKrBCMji7xDK2
zFH6wy8Eor9eI9nbyG1K8u9mocUQyDaPxS0O2fKS6L5BFWfYtyayzUscB7ORppOi
DcRr3Udyt70ZbeS/GvWtKZJBQaS69/EC9paJ71ok7WiryQVVXTwsbYtp390UpdzB
t62jxG6JLQh6uMLbqJFie3L3Q0HJjEDVW1Jmark+99m9fcAaL/hzknS37eBc7Wgc
S+JctYi2BtzqxKpJECze/jCzmE6g1/9h7RKHSFTwr+ZMmpVx9odl7pCyQ8aMRIG9
VkexxFq0nabYxPbXwGh77IO43MwPeI44m6HjkrFtcHqYjI6z8UBkV/reqKqf9Xl6
jBWRd70JY5gKV3HSmfajz8qJMeG7K8aM10n4Fw2Y2z/UeExkMv4p+FV3aDD2iKDN
22dC0OMQkDS3UX0R8nJIJPOrekAU6x5HNynqCywnwO2C2pB6ubIo25qGgr97QZVN
7Agw4UnWj0MSfwx5KfHXmtdwyepnLfPOIJgysn5u5Tq3LnaCNxT3cAdeUkov9nME
bGMgUbx5xC95fxb92WTSQ8TrOKeWow5oC83t3/zgmomAMgABfyQtoYNNOIdnw/kf
pB0tQRskjPESTbVPiQdWfyFX1y3U3i+k45DNrLFKGKLOXkICQnqbovPmDjGdcaXj
CBUZmSkBV7GlzgnidWhYfyFjJAgRGcFm/gDAjFNwieD0OtXmDoTbq8M1+ErEgccx
biwgKcVi4Tf+IhUa40eBWoWwMLNIOaklvTnQxujFP7ETWtr9cxQZiT9OiM23W87S
ezffdfflnK3OKVrIydjixSlUdA7fRxugw+nCVIuA7FQyo4jCH/lR9P0E6UduNXdb
NZvLmp5hNGI/YOLcfmJF342w/2KI0Qfx07GbZcfdrf4lgSqBESmiZsvaqK/4tgqp
33B/XjcUTm2nBp/Wpn7v0mvGheNpoSfP1GxlXU/2EXx2NrDHJ3YTysuQKxgKT92R
3eAmqb0LU3bSpzosGv0k1QMKdY3IkL0NUDYShufNphKfaXniV8KdWznzqZp3Dye8
LWQ3FRqRelqm6XQEdQbXPt2X27YWH9cJYnImt6oxNzKTDhcPYz9czXH3izt+JoaQ
qYU16o474tTufx4bCLUm22NfKF0UTxL2H2OqpG3JpmZ9EcxqHsc9toBf6oFT1UL6
Pq5GR+PKGlUjigbIcoZd0bXsQq+Sy6XGzsInY8jD6wx5evwzDBlhddx9Wu347+JQ
1ccdov03M2YBChBtMMmuDW7TFkypIxVwRphKQpglQxL226jiQYn6gC6Z9WkmqUWM
PtSsBD3nL2IilQMumVwI48nHAOnqWGo3GdnXEnIV982jqZz+5rNqFPDI05+ULssk
VFfKVot2YcPiB7ySXWQFqpQYXkuevLgA+xP9s54b3YcUONOI8sHN/3YVgvcHFagy
dCaEF4HMAL6GBispU238Am7walNR4vQUaebwWbaw9INtYc+cijYxV0/A9xsSSj+t
ARmzqWHWvrQdH+zh++y819P1CY2SgxCEQvD2rub6B/i+hv8Cbi0McoaCKbLtALLc
XShUXN5jt4SSkUABsLfEKcKvEEPgSpiyqiQ7TiLJO+MqcgOVYojFIzaOZJP9+y2k
Tz2cTt2TEHkn51t3lJjQdyc/ENOb6nUrG/KLu8vNa5H7r7wGLDHk8dNJDTKEq3BD
fgRZcvgdJAP/SgjAEvVhwwioghe2/AWu+axu8kaZaCY9cnbvhI1TqFGscJYf97m3
LBT/v51TlxZR9r6ttuJsudb9u+ZuXDT7a8Hg9NxDfmqU4S4Aj2LBpUnZymzI0T0h
FNJ6TW+//rOfAvmnDNQik9mt5tPyU0ADOvsTpy0aM9biqampENzsfHwf979OM42F
cHLB6vW/ktiTR/mrLoJyFzxoJ8gHBbDlrZkbgq+VBcQmb7IKl2Ke9V4TEARjYzc7
l2Y3biQnGjZFuA8LcWGJJA/X9WrYfkr/0O5lPQIW+5mtXliJLfl2QtnGJte0K6bR
SXsAT51f8TPGFV7dzuEv4gxpJbkbSeukc/1Wf344ov2aZTvYRz30TBKutdOamXS7
OGyL0HXmWrkZITuX8d9nMfQkHHFS4KACERfQur1F6R1t72wcfqGi/ivIPcaMcHYM
r3yq286d2nuZgp00VemUAEGSreTwIjxUqqPTi+peFC6S7E0NLYHEYFoR20U6GA4y
uSE4GFowz773nwIQtg02HPrV8G84ZxqQjMJaoguYUGB8eXNfQSMAMCSVMiZmD/A6
1stguzDCfEaElU690M1KpLotjSyD1ScJPrvUOeF0iZDb7SwKZfkQCycbZ6oabc95
KOK9lZ3wXsBD0RE5fIXNq+w9ydLk/XVfaqbdYcm8SClZJBTPxUBbLSelp81tzxEE
hhWhgQBNu3yJLkTNFDY8BdlMVMN926jlx3KRQ0CFPZj8Z7KI3wREXy4QDs1gvwX4
/A8Gu8qsTkVOcouipzyzNNbWiL8elwfsb9LRmbNN74yuAk3zRdX7GkhbUX3mKvf1
P96L3Z9O8nB+DGHzBzACOewIt3yj9rLSJwQFPKtxaG6fBwtDY9ZD3nPoPNlFXqAL
wMF7wHTH15Fb9BPlkHXUHf8ivDqZZwNhEwMfxLU46sB7f7vOv6t7qvKj4gCIOD42
L8mni9L0c8Y5HwLSmSYklW792tP6KM8XMgdatbKjrDnuySqgbYTVn6b+1sznEapS
NFD360NinKVEAR85im41YY3btc9INYOO+WObQaAgGt2+M9Wn4817uKAPWXAu/rRt
Nmakt+sZJk6RhqNHezQ/gebEEa+PZ0F60eptvJoZezxJ9lWQovbhqq05KcIbI6A+
YW3FPGMplYij3SOCp/TUaJDTngc+Y4i200isbEmv+27PToBlcND65hmpGxKKTrGn
R/ki+xDqaMrRsDKuwWajA32+aWs8GBgNzDYWauz9LMdXCxg/+D7ZJ3YJUUr32Nx1
f2hpgfzpMkEPRepNiN4R2lxKVN7brjInCMcKdCXOzG2qwhsoqw10b7zefp1AES1Z
pEIbTJXQcTtp7dldjhE3JtKuxa330gBR1Oi9nxorOXQUf6lAhPPqLe4GqZH/SHot
AMvHnsp4AN2hl7vWNRW/HcQ+2GpMlx6ZYIOEJ66/IN4xSz4CsZZy6fKHKMpqEgCA
+bXfFTRY20IXfSKnR1KEDQQArQ+Csk9Z8unrHWnVScW3zDM+/jTjWHHGcaqYnVHj
BHsb+YEWRm/BuSAA3jVdVh/unKtCKIb+BdEdnNj3k9yKtQKhO0tAuLkhd/oEPQd4
bnpugevhmRKWIutbsGfEge58fuwlwNydqTv3fp9gcp7OAu7RttLJyqRnytaV6auz
3etG0jDGpPd5Nq6d9JdFnFWo4EYVIQWGqauVV+BErKMdULaRqlcCFd1PD+/Swp18
Zc9EzTry592j0n4L1XT4u/RuNie22eb0zZDL6fILecFWVfmLFC50jXPZoP/jqv0h
k8gAOtnfRcW+N+IzSX6AabVlmCKbV1pk+eOdD2D6zVuZq1mFEtEb6ygHILqNJJN3
Fougyn9cuG7eN/qSTn5p4d5botTj7folUx56AA67Ya6XYj56tSBoi7kqR+wDLaBu
9EvCrY+7Pt9HtJUoEC7z2M1sfRAuxZzOMy40RFJclk6qRG3pi7VIedaUgGoxoOO2
O+PISovZluzaQ8tUXXNszpPaNv2K7FKHB8K2legZnXoN8ztnWFrPYVKr223CmQeY
16ysHcluJ7Lq0d3ccwj4RBGu+A9skKRnYS/O5CpY0BqCa6bksBTtayPBzR4D50Jj
/nB6vCO9oAC2cj8mX/5LPosFNUuLB/rkZt5bFpEoa/M8OBJ1yDPZubPGpVDi1WNE
BKEPneQ2Hjg63tUWAuY4Ey5SMRrnsxpsMj/tk3fWr50jNTg/WTae8j7Fc9DYjfD2
VJIKwby+lAH4nrLvltrO9PbdPidn3Zf20zKa/Vfrqw7ndHVp9bkf/vyTiXT8tgKY
cJSd/OfU0U6i/uKaPEGpabPGdDfh998Acr0vZCOOSHeUV6p+pwc8J++ORk+KAZZf
sIX1JLjtBbwfqm+n8dLqopD8sYxL3AATAikM3DCKT21FjHGN3OwmfN+KAQpB4X2J
6CRsXAC6rxgAkytqTLp4LvK1qJoEaLwuojfWKuEjQ24mI0RCxUzWjF3WnI36XG9j
JzZabd9sfquexkTvkBoYPs0V64YTN+v8oSTkV9U85qdRvZJ8vBHjjvU/9jdKiJ+m
Up7pKvf5wyEhzAgM3+lfRPBQ8rpc7qWj112dipGhH+64KyCTfxrKqkHCm5dcNjaS
B4oKOHyPrlQeGpoIQ9HHNK1SIpcJlF2gTsb+0mmJajYck+RK68nPpDphFdWt14yr
ep47Wwo+gODXlXUPLnh9toZCSF85hvheEt2uxHwTgWsGSEPPSyNApPEvs57oQnYR
ryW+zrWXEvAIGGSd4wy2+TcUj8cvZQsL57U0BheHq5pwIsYfzSzJ8MiunHyXXsc1
rcmhs81IVSlnjgqIGNl15pj0X1DN2WRmIgV6RqLvEQvix6gT1L6sy4XGYOvv2Lic
G8+BqG1+S6LFc6z5IK424QMBmnQYJeHA8YIP1GUjT5r7OjayAnBC/6vPMYi7tXpA
QJJaQDa6/O2BZ87aZmT887VN1dfxxVm+wFa9jDz9XQV3Ih/NL7l/ps1WrDK12Dsk
2OZdlKaWvzrmxEhOdLm+2CKWmcVysx9i6kYELR5TIbI7EZlSV0ZJNbHLc0OGC9RC
CGfGo4kdAV7XvL027wGt3D36q7cKsHoeIhkDKO85o/rmo8sTKWXqndzieUepyNDg
U46TnlgJNIq7Gomxi54JbyGzoRTHdq6Kpa5URwbWb6/enR7RefgnQLlYOg9bg5IF
QoP+2Ugh9KYdsFqNTohxIPxihidgQg456TgCvI2YBJGtbwhbULOJEugUdqf5IOz5
niybPzFUUSzoieYqEQUYQXIyAA1Wj/zHrwV6ot29VGE4DaAv3Pkxwae2Bs9XMX6M
GxlEvQea1hrsWiOimVn7WhkpSlLdsGERV0uMFrMsFsVWn1F1ONf9JQ0hw8DqEMED
VVhbBo74viEtYmInxCgNp+ObCJDfM+rBcohfXKMFSCVj9bnfvQA0BUZezgEbpj5C
mGzKQuPyFY+b0cTIqAUEuz1ohWxNXyfKwLwzrEDf0KgRudQPDSnFzeULZ50CxwhV
+Uj3GkyeFoziBlA7sWiPDsrZBlD1iBAvJHpCRTIBAj1WVAZHYyJBBeN9lQjwAA0X
Wcv/kZnN9+fkrwDX3QDN/pptsb5pEkfZ4DoWArALSYzcvENAXMOkiZzGwtOw0kHP
xvwEenA+PZC7UXqhgGoBWFS59zaBXQD8hXf/7Mjns99GZCTa3LJFvp/7NzHx4cgH
BrV1qwd705XyJRVy51FcDAPmmV5Od9u2yjMd173tcFSTLHUu65f1eUWVhekAvw3C
MLVM92yUlyd/I38HAAQihQ4qhE31sl42eWOzO79gfRYSV7gOEOQTfD6bmfyKLqDa
gHC1PLiGRwFw7Z4J7p8f8i+e+wuJeIo2PmCYvwxvxvlodWO+lq2nDnPWXtIOLCKg
WSgreD9EWh0x8A/4dpFWVUuTSRzx5eJaa/vzZWwhAb7SIgaRGFbQwSQcGbXsqaNC
nrqpPmA9Pggo5ByS4A9E2/u4rnscmmcNxWKQ1TMcSb9M04fyyZevoOP0U8Y78HW6
GaMPFd8n0iDvcKydWbHqh3d5gUl2N9pAj2PZU+ryFkkLK3R20sdlGDbvdmfLJUjg
Z3jdFv/Dqip1wrPi3cyZhXXOP7JOulE8jh2FQ26MKQ5e8KYPejFFVJ0YTVjRG8HA
4Ufr94E5aXpsO3758+p//yc30SphOnB9OPGzeHDbfYO9V7T4zpGhlPgGny0Ct+Ll
FnO1RECadP8vTDxgN227biOT5S5E7uTjEkESJrc0ZvWyecqx332DgBykek7a/4/M
wO8el2NVD+FIQXuwKn7MqqW7MdGl/msCJlC1NusXwl0K9ZQiUCst/qjAsrAcObuc
2VoyJR2wIFTA+1YT7ppfMVvGq0IrHj3YWhhycHz+Q6CLeQY7dBqSEkgku5lrQTnA
f4igE2agUsIfBv36VSwcHtF13ez8KHCjtv8wvaPyoTLGJXE50qH9fG0MtXXQbgoV
nEmupjKLNGEI7en0NiEPK8bo/bgdKJBLEWczgMXlT1LSBlqpElm7nfTwK/Q/gYpf
wdcsRtEMkMunW51h+7mCyn4m5uu3rC8fok9gxovdYcWDSREwtOGxwWzMDLqpaYXZ
/UVs92vRjTw3FerV8f6fAeaoYzH952E9pqx1Isr/UrJBJj0NYN73Zid9CBNdmqK/
/WnFXUERfBR45HFTOe2l/0uwh2aPbB/DQrSR/Xo9Tp3D1lQ9ffxebva4zPqjA76f
odU7YdV0D3UU8lwS1n30veFSwU/4y8sgTlVvhJPe1JeOpAqkWwzsQ+6t+69mGqHP
HhTCgAwQvn0FceYfwfBX6W//KwcXjKewyKfvDRKZvtdvsE7sJJ7Uv57CJOUhJfP4
KUTLbaZ/9BAwxH6qC91wMT52ONCySOPQkciXvC4Moejr0o4cn/SMdTTOkVSYRXsk
XBzJzT+2Fm+ATNTFL/tderkl+X39XsCn7M3Hzx2CLgYxsIOU0YySIWxSoaKkF+B+
j6lkBhelOkikOij6gvGtzWzpJQw6sSsqSSfTWp7Pj4/o0GsWn0AVdQfOXlRHsA1q
Ak675LV8XtWJBxq6FbDK37jf+rIuKsng7TObEITSGwZ20X+yLwt/WqtmJzx0GpIM
1qxD7M5VtRkEB1qxiCST5bGvm5Ibw09jou4fC8rHZbjMCMIGtY5MHkse93U+NiLo
ZcC3iu43kCRwPiyFSJzdLVZ3KIfQkctHMxbzAoTjrYB6NDcZbRdTE08YFMerSnqH
pKWHDb8TKEHibTq3B5+g+GyMJiILWMhy/FMtObzbQMv9DlvyIcaouGopvxz4X1wB
9pNN2RmurYf9L+i7fgs4u0rmmMROKyond5Xez5EBpZ2Ml/Hd86WOxoXIYS+W7j9M
5M4abrRLa7DOBfspdTmcjBStk6FvV6vh9bTTXlq7hStaDWNIqOWl6Y31BK03NE1S
EpOJx3nKfXTICghg8JKeeCjzpQlGtPtjMIpUIFJFSrrVk50EE5qSBfNZzGR5+0Ok
JqJM/6bQvZRKmizZzv+HY0JMaCEukKdnesX9NPAdFBcjeRtiuZbTX7ALD2BJ5zbT
lcUFPx/qffSm/9cYYv4Dy8hsh+eMs6v2gbcGG26jUc0BGaX0uCqMlTYJBqAdWo9h
wDOVEA5CFQsqaT6gRmGE/T91L9fdSV57c5E0GfWECEBkiJTalKX3OaMIIgGrdQHy
YbogdyMe7hMQyB4GtjIAMNWx4X91IrEPI8JP3lygzH3MiffkmCuXypLh8FYA4+uL
NOBZCd8Aew+Du34dfjWXt2m3xIafsv5ROiUODfgWste/7AJwUXeOJ0AmP93NUesg
W/TXB73OvowLZ7GDRtfbHvEqA1UNUQm2CYwddlvYAwOlzeIc+Fcc2bUzxUWzzB0r
hUYF9ezfuPmBs/RPp6LJFWotuwQntmWp5QpkjNbxSkbQMdZsdRvwnCvvu6uEMp0l
OfGFBV1a0Ab6M5OyAchZot8LipA0riDpG+8U0/g3gzEpKrfXfhGgN5fyhPA7OHoa
SqUIA/71PBZQZLvkMa5KoA9fadR8Uf3kyArHu49oXKXn7UC0IeklyFmYSX6yl7up
ZukJaDyMtuXZxn2QXVUlBVSLhjYZ5FOETdMaLuoySaAKu3rLmjP8s3WlFXqCH5Uk
wD202sMEBsaF5KLmAQnONh2hvJA1+wVljntozJgLheqEoGRNaRjnGbTenofOh3wB
lupm/YTBw5kXfh2wj08Fez1r2y2PErYEtzk4BGFE+y/iKfvbcWDOlA/2s+KNBEUM
hD0uieYh6L8bTJeQKmmi2ffr3RWLcQrGmpJcbE6K9q6teFLlNsJ1nxvsGr06lpoY
XSVQof17Q2vMa2tVXwMgQrCRn4R9KQC70ppBIdxlSkiTpZPRYGEgP6gD23Q/ev9i
6dp1N6MZLKrBIpgntHWwQK0KPgs2MdOQHcjiZaQJa36w0N/vJPPwCOXXztzGnN5N
8sag48vODgDEnUzv3tZ97OS3RJsDdCgCOvt/PWYgFDO6xCSdR+vtRvjvUNTJZDvD
nZukqSf9APVr2hUu1D69xgMjPG+uBQLuxjFnIfF6ihIqzFylCGC+ACERG00nItHF
JekQmPV2kyF+zJ7iPfb4+y/hFV1dBMvm2KZXllvexexl7IAh9qKLpLGQkKdxgSF7
TVHIYRGWuUJWsW6lYZsoJa6UQd7JZeHp+PZctYrA1DgFqidPHbbIA5/y4E4DvWXS
U6XmRzpBRuDazAcBai+gc6ubtmMBOefJcNIV5akVX2I7aXV2hJrIWRBgfkFAiIj9
w7+eIxM5oaTEiMlRDJ/0AaZkx8iTm+bVs5Y4sOgRPb5bPxxFHXfHK3X9bA4iD53S
CW4mrLghqyZc27UAr79IH48R6Aju9MKF46UzTML7n66BqlUmOzxJhXQKnGsxIDaf
Rc+DUwZjZ2pFG+FtGPlHkpbbRa71yvsAZpOik1M/aMxCIagV2e9vnLm5w0JFdxOa
ijrS8EkUBuRWVZnnMS4rkyUuoU/Pc6IpzneL8+XkqMBnmUUrq2QhokRrVI1FaWBW
1GDIvLuzDD/IXE5sPTd38JIONAJ9ot9WOveGVb3CugzM7hVsZn9swFTfot3FUxvF
lVLFG2D6mBr4y1jJdl3OXul4aBtODQ3+lFABQYNSYA0ugBeH3qci943rKqbM0LVg
0UcC88jsvFGPrR3u8kfAZBRfEV6ECsDXDC3eYh+yDWhlAlvWAZLEGaNoqO1ew7ZE
rO8gvWacYsVmC9AhIn+MLtTPc8x0+RwpvTADTtjSmaewA1xCPCtD2ugJS7rJcjXU
U4YwYwFjcMXgwrxeM0SbbM3Yx6pWOLOS+GxD+ueM2GUOjNomEek8h4H2fCFx6JD6
qT1t9VhOSpqcGBNW74tD/7QcKTuEEU4L8JleSrx2ddsn8fO3sGwyu1dXaom2yaXy
93m5BD8C4PPWKJpveAvo7v4LBMd3A81uELx3VaaKzQK2g5u+R44e+YDFplvQOobM
L1cndxJxyzOq2kWG1Ya8gY7r+ieosoTrY/lgwU/DhhJuDuxbnDEviRQYKsyF3hRC
Yx0yWt5qP3Ga1jt6HHyWzvMLXU2aoetSRqj8D8CrsyG3UwKDt2H1GIQKLvsuanIz
/b1fVgGIEZ49hs4U+6I2buJmcg2kYH66KrZaopwkvWvtJUAQwvCZ7AOZclEQgh+n
41FjtA4V7Hn06R71sxNJ+UCAZP44ZWwJlojG9rWIGBu0GxwdYVD2oz/+iprRfhyI
tqRkFDH+LKJxZZmFjsEw1mWLPHs5I9unITlHX2NnmAgqD77ZYfryHt5pxtipUsan
P0raZzmns7XII+g2irwRhdHEHprgp3DbxpFuBGzmJvMFVzFjiNoRf7zpfievwWxT
1owQ0jiJFLm4/5FTlwqDKJtsuevkz9a44006DV176drSJJYhyPWfJnMjYMVEs3Vx
Ryw/IW5Hwq+VE0+MO6h3wGEly1PvfIkB9HE+FCjF1OOoKeSEtiU7cuDYYs2T9S/5
3ipJQpQ22DEalg1o/LLfp96McjfDRgMCmIsSgs1dkUo77zEGy4gAmroUMhp6L4Zd
4SNB8h2u3oMQKx7hh9dBzR3AJpjN1pF0M10uN5HcoPsIY8mAZLG7tSXMEwad6Kn6
NJXoy8HLV6LYxhULPI5OZj5ML3oHmLg0Dzhz5ble96wXuDIkTZO5jPfdjFPrQMNV
7MoHJDKJwK1NDemqlRQ9Maj6/Eki7Q4k1uniNExUNGYO5BL+xK8x9AUY3VirsqjS
lcu9oRK0De0cw1zEyfsRT3LqdVBtK/iygn7/lor4K3/E5+5cVxv5FkSgGvrL4P4W
V9kTtrhoRV6Kc1YIhC3Rii7QqWnIpLQ1LMvKqnQ+44I/GwDk3LEtvBk6qIOED3R2
iwsMXkQkttlhoyp8XQOjG+H0vaCGvWyu4RH4jye9egx2pdEq6HfLxqiouLoeX3TE
nxCnE06CvfPL/FoErNNyxxekLoTS8IHz00T/Y9XmX80ocRQNGmPwoOIY7H4lJufV
aLMb1DEVOLyYzEKj6QfvnBT/iRPnQtXoQ8MS2cDUGIdXthjqDf5Jkcl3EjeJjFVx
WoaxL5XiNwJKORlZ55gAePRakYWfx20rjv7PsgBlMeLnpU98hJJbjuBA++hBZGHY
ndZ+4ZkDsN1WavU7vltZviySG2ajgxaDSDY/QmIkSjghNOGUc/t1Z8VtjKYFmYbk
kD6J0nR7EGkTpqdth8gzqvAoG6qjzbLDnr6G5v4E3ufYzG8uFJcI5tdMcZDTvjXh
7hR+Z1pX6d6pvpzU98oWM1xobIa83+VsT8qNwVsrWJ4+kR0xbQkxKQVANZ92U419
oRUjnHyVMheNlAVWfnEKlXWMOK6MyCju0ysAiQ22eDey4c+CgiDVY9KNetshXYtg
BsdIZmbwLLFn4LDnlARyYaOo31Deb3qJaRs3/IMj+DlUqIl9+pKRqKBvcJ4nGuFd
LSRlc4Msd88k/sGwSpzLJ7iEq4bCIHGMc8wfrOIEMazVMreL+/V6IyCiIfgBLtiD
zS2i4lnq5Wk8cV084ZQycwmwq3ZiddRqtaSevRVrg7fCcf38LmsTYTbx0VIqKS2n
uhyKKZJ904J+CCGwsTvgPSr4aOGNk8fcNpSgWLgsYZLmNbPYnQM38wRtsJdgr01F
+ASLvv2TR+bYkJCDiKhNvHp9bFfFRoeRZbfKL6AQB9Ad0yKcY3ibt7bDFFAxZfj4
n7ggyyHj0eHnaXMQd35flTBCiMNsKoWBTr8WNImO9ismiJQRckyb5C3cBfwakOmM
qjDX4qRYok/u1/qq/e8rQO3vY8XoD9HjHFBD1O8dLJAtPEqGp2osbpj6fyupOWpz
epc+D0CLf/mT8rzOLWDqoDiq5EYwI2qGqcu57tDGvK7WvmJguUKfazItLlQerC1L
yZAWxn96F2UAh93Z6Nl4hj7OmoX1GrTG8xFe/9izJWKUAEL9s4wH3SUkMdRKAPn5
fbDi6jbgT/NomHfK0hXvglU//l7Pf+Pwj1K54QXZqoiTGbZ0EZaccHBSMjzy0hr/
xJ1ijkIfFAmvDgmiBl7CSd5TRr9cbyR6tmnzsV8KKwP0Iw6zcVOt3hZ7ET+yJByN
3T4cP3GxRifuzjuc/gW3rrAcoLvRuiiAkGXHbd5jlG5U7C1gJnbuXV7vfSk3UPjD
gTcF6r5Z4yrWT3g81sh8nOdqNWVPuUnElEAiAelEE9+/WdNLQ79j/ZshO519BpLP
4ayinYhb33r4QsT+0mnnNeS7JeKp93sCnqnrpWNfsUXf/tfASitxV9V0MaNbgm2A
LQ7noxwEWcG7/u0ToLArpOa3Swvz4mNucfZ1Ltbawe63Mcio6L1tnu2J/aPPeJKO
rBQ/cM7HNzTnyaV0i+adrXPz8gwBLu5woV4m3OzW9uzOkvSCuGNPzaZFgrl3QcMT
CDb8oUhbMxM8X92tcTaIQ5KXf/cF6Tw1KSYt+34u4n0cpLa6VyAzqeOT9KJm94Mr
9xyp8h9qeEqqAQbk/KsFsPtsifktUF6BEI24W2GBjCBwQFZNuqOlAt0tVJoZ1d/s
VAggiQBQaTTBFmBRn5gBK5k/FLWyLFMzil/sC+TnrL9Vjl9Ysazc6/PMXFrKB4Gd
pcJaXKZqqmNhuGHCKYysYdl4Hmu8K3yoQrYkvwy0VDzx0kpcgktfaq1zYvzucRUU
KNLKhHR+s+JcHr5c9zWtjCfSymbLDB2WlTPlZflfZzCTegj7MJam8+ADTw6iyGp6
PDNWbYT7mJ3GVMFcm2Qg4Z8Rzpyiqk+T+h64GTB20HLNziSmELXMVnDz1HT3WDdU
wPERb3Z5QodST4Wvr943tb93GXcC3rSeRhs6u7KNva5SqXeOeqOJK99hBOkSd0sx
bEgt0EkimqFnIqF83lpdcucZKVznYrH8NmB7Cv09Av30/cMSTxqQRFCqykdjZWAe
xnRQGJJiQuzMxznTYLE1x+TLhbD5W1A4PPY6b5a1MqmMqKoQL0YzomOgYakRqACr
NqdytF1ARuCFnM0i0Ixps6LgWCB9r9xLyJrzwevT8U9rYMTWwpNz9ewcHfMG/tSQ
MWE9oFIY0R7/XNSjNnaztLphHc6IZPoz4sU8lMPMK8yLBQCPHqicV2dTTKe+4EWj
PIzJGlatW+DiLzs46wVxAIoS/GLurvTJQFYTOJXUcviYbFtIiZtH3w9sX/JVyPVc
FVgEGiJDDaHhEGxERFnrFexCv/eM3G+564fE/JqUHGtNuln8tAEJh5rw1OTe/G2L
aaCgmYAmFOLBlLUFUPmOjUwXRts4R1vefOCFgvaYZvGcZmB+SYTXDiroHAdr5vZ+
uxVr8COoSe4sonCWFo/bRcfRPYxbziQVbDlU8FkQo2xouJq+zzOa3vxBxeaPX34D
vUfJ2iYvt4XHdlm2Pk5wIA0Cb+W/B8HzwvmGpmboD9LAOYyBdFt/uVvAROwVVzRF
1eD0BOwVuQZWveAnXD1cA8vyAu0A1SpbegTmforODR38bGpK7DXLmvVYBa6tX5rf
HJmTVhQOwv8/5c5LoT57yqcxTqamh2LlVInY9efLdeMtDXsHtq89QM/+JxN6myph
TMVIyLzhxf7FPGZgXhvQPDfUSxVR/0DiLDvzDovEtLe1U1Y9vkWwfzYf1VuuaIvX
ZZQK65532BKWmzXRf3aJq7Oe/v0W+WxoGi80UCMmkPWbhT15ZVLYO9pFFh9+LLlh
K16QbDb2bUun9MpHxRYwXvNDcrA/W8RsolAPloyNxYGsa/XJBIlva4S11w2RYwOh
zDsbX6yo3Isbwy06HJ3CR6rq1fDZ0yhB6CCev4sqXhEnkZ+K8l6ZUtN7hCOV/BFZ
DaoKpk+IESZIkHl3Aig/wThhMiXJ9xSb/2+lW0Oz7EwTda2nd+Zg3CmORaI8woDx
jXbnqnGUAKO4tPkJWxy0s7u7leZLG/MKqHvrDmPM6xcuK4WHCni7ZTl8WpQjRPnN
zDM+Z3HIWSkuZ9xKrNR3WHMHwiI0xbJnHpiqjGmFXWbx7VYiTgNP0qlzQOzw8ig2
TQi6Ldg3vgVYhstCrCkJDduArIlx5nB6FWsnKhminh7gVJV9skaRprunVsy0tb7N
h6oPv+4UUtFX0+0Bq4+d5I+y7ENsrL3n/JRToulGMQAfQKXp8Nv9TsScLUk6hi+Q
elujjykTsRW/+3gfPE864ClReenRNRTkkog3Po3nYmI6d0Nql86JlPeooJr2Zrm5
45oGvf48L7K4KiAED+DAi7UaWB7PohshbP2SE4sqWIdrQ15d9dRg0oRn8LvBaWuT
W1aPfWim6wq4h38mdXv3ajX5wO3kS8Ewt947yq/gair9qbeC3AgqgO+RN7g7PNKW
lVLy7moE8NSS36mSZZeaz9128V/Gf/f+xsT8cr1ESjp3qYqko16YVJe4p64Km/Dx
/IA5V7+kBj2Uf1oCZMhEOIok+0ETQSS6HcLuxwW1sihI+KVO7hsp1rELS7Bc8QFD
NlvIFwgaU3iPY6pe9FXq7KuVLcHh+P0CvGttt0slgjkdnuj/c0aBXjqJUOHJg9yM
loy+SM8kQWJwIdAKJCdewwMs/dcZ1hyAAeFEWs/buqbhyYLk0FsQ8opwBkp59tbE
TI1cmTRj2dQ0hGpyRlHyPRKT0KpBdHgUdvBEafRAnvugYfCufjSK9GPRldE2qQpp
O15vCdtPbqC4NzssxcWwqjUq+PTjF4qqVGdJozxeknkYBlLhgmUguT7BGSMVtjFH
dc4dd3xUSsbaLfIz+pBE2WFpkoJnKCccc2aDAMUF/Lzkt93+6fpEAMvNc/8zTTBx
EflL43q40wVta6PkBrL4FqSGDMi7Pk7q7h8rVVVq5FrEZxH80RPz8xNRejaZpw+q
4ZdISzciX+4yO9lFUWWckgcfPJAXnNVRqZHxLou9meVn5UVcthKlmQ6am2WI6c5G
DAeP5f25eeAnrtJ8YjFJyczcIkfXrtyNlPzqkgKoDyU6dlk8ZTZ+3wd1n4HCJzkR
k+9nIkg2IfvMEsREvkh5r1GBc41Fm4PDsE+keU7gtlS2c9GvDVB0ncYHxD2o16fB
kHv1sBkMRhHOiBHKADgOrkT1tjuTkj/bHH/XVzz0iqbaBP05bazDeRPwQmv8pHPa
jE/ReXfyU3NT19VSpBUc4f/QzLpHwRNZJmXWAiJSo7dVap98/aF5U7/OdmDLx4ca
VZ4LQw5/oE4/6IOznjJs3IHlHq8VBCCOrmwYInZQSjg079Yqzpcogi133taOnhkN
Ivu5MsswnFFTcLpFyaS0/XWuBFFvS610OoVTsZJB0UW/vt1w+CPhMOfJ+msV3bb/
utvwE59kcfO8mDIwaR0KFkbyy8fBNS7T4Q99OvANVSQb/YF9wkQme2ItvFSvSkhQ
xrMaQoaBurPnqZVtCtxNQ0cSopLi1qttqCZPxt97xcj4XF5HYbU5z6nL43D/EM6M
MPRSS2uiAlqj2aUvShJanS0YvnSrC5j8j1HRx01YFcUyWXQWD1s3P2FXEpNJFrQi
dH1ntd4PB9n2wxidM648FhYHZY+yFr4UXC413YCb/+eaTPEIG9YymqBO8dPYkp85
rx9csiTb3ufNB1Z3OmEfhV0OSFdOj+ahFeU3vOqoldkmEcuK7j5P0IpkFfo3m7cW
o5JNjkZ2iYigzE4ozHWdmhc9Z8Ksb9krmuS2c9yGQ3hyHm1wX2eY7k3JhpmhW/Ui
AwWYErQIFnaLKKdxGmfr8nGVgwnfX3HOJ1VBgo/k6h1SthPp6M1yk75ZP6LCT32m
lHCEgFuvE3t8/wlBJcyIFjebtBc6F3/XuIZgN6Rb9RUE7y8f5Xxx9Cm55HQryLJh
PVrIa+8BS0xOp3AwGi7j1I3AjWuowgZou0/cNmE+vIm3gECBDm83MdAWeD2S46IM
zc6CiODy3g6pXWNB0oSS0okrIqWYKNuqETKK1LoH/PthmNhWgBx3B5HvMqIBLMDd
K5T6lQm7yjZwMjQbGfkwtIPwU/fU1siVPqFFPEe3d2NLPbxu4zFqzhsF6eCHzmzK
KZq+Ksib4vitB/I3pkVisMac5Nu3bC4bj60QJbluGE1QVikbIf9XgwbMtMs1DQoF
DdWMQW/tCszM1wMmvdXbQVM4imybjWBbjJgegWlYGvUbK/5gh9iovjWZIFwTU7zH
PEq8wllNYY5s9jA2RjZ7PsA4rIKzi0So3IIAyH+t35BdeL1rF8TM/GcdtBmmAVgd
rozyiLxI4U0E5Vr1i/IoIwTQedieRYwI+qfTC8IRCoHsOon4fM3qlp4gn58s6hIw
ck7DOWeJRemFwFgKj7xOlFXHTmCkwww3rqdeE6/69Xic3UAlw9A1/QRQQUwKHY30
9B+zp+ahU34so7oC8b58ZrgfwhAWkUPFDICxUMUmgSIGWi+RHB+8nttAuDZiEYEt
di/FwfF8S5MZTuwEv/ivWx4qHReMO8HaC3ydP5XlYPDCernMWyJOmujFJPlicsSw
AZ2BY79OSOd/s8WYN18TNNDmQBOwDrJ9l1tlFqUf9F1tys47IX7vpKzu0d4k3Wgl
cFJ6qmk/DaO+nOHJCUYVs9y3PsVkyU0xvEEtv8HE7Uksow9u+pThZAN7enFvRlVE
X4UM/Aa8QocFRlyD0qfzCUXbRls3r4/ZvqqerFQm1a1mA41qwUdk3mOQxnZ7u0TO
57MtuA0X8Dq7Am2lYM5LBjldMkaYz4hiPHlYJd/eK5dd6vWY+Rn78ztLW4sCLdXL
XatAqpM+5RIN0PKDZ39CLScHzG7lXHt7uKkkcsCJX32Icuqojgsh+QZNMN22We4q
m+KHw3Dprph/oupAJYKYGU9WGDTiOUuoDET9Px/D1nNd2E+KtkIpk2Ig7BsbnIGX
CJdMjoDcoBiqcrk/ncEOcINT4rSBAI1JB4M5LID4puefUF8PJtRmq9sdHcHVFyLY
9OunfV4h+s/QEq52Sr3WK8RA0yhHdxj6ygfNWgYmSHfedv63+S3q73FrDexNYFuT
DqpGiDH8o9OaGQA3UTZL+7g3Scnofw3xx20GdFFGnsnU50fBYi50Rfh073C1PKAf
r1H0eN08xVijitrE71QUbywnncZHEQs+14wky0pINW+dGFacm2Q9wWUf4/Kk3oSt
ih5D01ZIGZK7gDu1gJ5Vq/0ttDD8p8/0ZvGowtcvrzrfBAhlZfgh9O3p80b9Q0Mo
lEcXZnJRyJywKQ51yqunxu6vpTM+fZVapw4rtAt8BmvqUUFMW9/LVUIhG+udJ+Rh
1K7DnU48XAZ3uykTBaxKZYexMcps4Ftf6Eq+5PTdbkMJGrEttpzM+vN4TgaAS91z
AnYJxLifqTAI16cQvk3UhFlQF6qPWiYcd7j6i0XxWsFjMoz3EYPSEBIXg9EVYNc2
YDqQvuNANg/GRg3BWL3vkHPTyBY0A4HSgNwaFixl/RIJQgK1SdYQ+hBeQ2YMvlS/
fQbBdXKwKjKR3wJgCr3uh259EU2LBAvOuosXpkxoVNX7ZHUik+xycSZ5Hck94jbP
+Ergbzv6lVNMN+u6EBMUbl7Hdplv/92Wb24EK+P5tMfNnRYMMhuPX7Cnwb7nGbEK
T4XPq7ladcIWpAcBv+7pkaracq2L5MhS+mM0sjX+YWuvUG5oPxOJ0/b7ggkptP6o
bP0bJLdgv/9U81aTiCYtuajshReVzxwj2yNPXIjhWwXj7X+JVkskPrhYaf/b1ix+
iybtg1tTRfzRn3hgqYNgjZLCVYvzODEDGsu2HWrTOD4BF0uJ1iMYe5Bxe8NF3HxZ
yAhjTmmyqdASwrF+oTpoyGdoQpGq0Dqd2iSqpFP9++dg7y57vi7L+oE8M6EBSBHo
X380M9dxitE3r/IXUmaQOnjZO0U/l+AeK33lk/FdxtHD2uoKAXQZ8tDCGUNQQpLI
3gj9hdPhN1kMz7hbkgfBS10pAsLKElfTIeevpHHrP0ZYjBIqEmULhOcl1t/D0lmW
gAxBcT8C6hbyWz5y7x5AHfeSFqRU3fN9dMn8WAlqzTo4l1sjA36PklUN/wVBW+M+
g1TuJEZh5amlIdI9hsG+9RJK3nmAFCv0JcD9eJAI6CkoTb7gK0+k38ZBOUNsl05G
flzSM70JeqXxfptkcvjgjkyLaCuHeOZrN22CpiyC1ysMybmBgm1nbUgvN1w21g37
hMrHAVZeUBwCRhD8YkMefewNdI7eSkndQjPB3lO9L0sALZIYldG2v1hzNfYL5ehm
6NZtcm+mclscJgnsl9K/+HvX5dLxfvVAt0Q4hraCfBwD5s6+2ybvrJp7mBrnknQl
9RoSInFGSDLzwPvgaap0tljcmG5xh9vZnfWx5cTP3e8gxAUa28M1PZr1ViW+0uDp
ZKScilMq5C8wO5Kpo+lCzHVhG7UTApA6r6CFIfYZ/m6zMls78Ix6j3iOKVogXht3
VGaI1yOMp5GZf/42FG/cA6YVbD7BdmhfZlnkfg4ruonys9D3MGpYwiNTXrxYEzA6
fAZyUXElnnGAfP4FI4Z48H+wqkmIyl2Gw5TtPR4VzsVM1zyWeyGbXM9Fe+nx6SuV
T2fMrrk7UbeNg8nDEQEwYL7tBMhhVvxL+4bWGqAwq2ObxWhXmuZ4/Wloq38Op9+q
Wxqh3JTaH38NlELY3T9RnPgmZaFXo7o5h6ZbGK8BGNkPpE/e7EcJn7BG2g7ZQOOx
Xkm8vr05JwWmeBv0RoR/uExcNsTvtbJqah/4mUSKHh7DEinzFWKfgPrU3RhNUets
aALoAxQEJctIEgRKG0o8Ftzjx/EedLUyfj8pb8876diWcbHLYMps9TYSB+S89F1x
C0IjAV5GMZuDWAnEYasoQGRBTCuvx6gHJi3MgJc1o8U6BvUvc78WDUzY+gDpHggm
pa4O38nDvzlNXRU5PndaPsUYTjS5A5rJALmcYrPWXu+MCbrnVJPlhqc7I4d73Vei
qux0NkUxMw9lG4PRguBTQKIxqGCTb/mvLFl72pWnje7dIl1I2sAIppXHokFHd9Vq
Hvqjca/cRnnMSXeiS/nC5Bgjxf0zctmfJFrnJCBBlVvMciTCaizeRQvMAVWD2SNn
09i2XcihP2Pk5EX73QCNFxwr757QyJh3SjpZArDwLxNWbSFVmWj5PjMMgJnY29g6
BAhfQE2KAIxKGL2GqQk1bqGRJqymu7kJ4Kd1sDMUycfrtWyUZcCafB3BAyOSS5gH
VmJMoAJeG3J5oWqST+THYJlUwrXWuJ1VIr9V7Wua4vXEofyjKR5mKdg7Bf7AYZld
ngl62vjtJXAZIWzlRDHWi7ykXwtctJ6NAYlgLgTu23+ceGeCFRhzqud3m+gmLEYh
5Gv+iJ6kgeSCHHdTjtl4cx3k4luiAksIaMnodGqyWPzsKxXCk+75i66R2yyO7Yoi
i26hFZLEMjpllQJ/Bx8D6hZbe2DLqTUbBUmsIUuCd3NV2WbJ9GHi07glQqeyciuq
emgbhvk2iptnqaQ0fXXZUNsQK1w8s4KF44GhlGmkNpBa+0m97X6442JwxFtp7i05
cadtzPLTZIeWD0igK2Jut5s1e2obgvSaTmmEDP+1eIPf1Nf8+Y/zBzRO7lW413Mg
XBNT3Ulo2ePhYQ+jyyhBTcRYFvDsZ32t3bYdJrhGKHKM2xJXcklfhJb4wysr2J3C
wo6xwNTSPpJUrV9NCo5g+vmsm3Y3nDDG8nMdGIRelXMFSLuto6gp6KplwAq+ubZB
mwRuWvMxGu6SuNvyQaO0QnFJb317cijmlsn+1yxmkcm1k0CGSKwuLgYZgAu71fTD
MuX8Wcx15b/Hi9jCWaHRoatGZ5IkjfDwe/52WOU+WhdLwrTtpLqesXWR9dIG+LZp
4C9fjUc/H1iktByWh49s30OKHEdX/L81dvPMe5x8yEkijARYazVkO7E+qo/81P3E
v11b/9mSqTp/U61eZ6J3sXwIqV+KR4SDHeeY0oQ3as8B3rNegiUha5PH+HYsEl+2
hP+pP7IWlrvuX+oss6yYN4AAPE5DugPLrbgmvtQJwxz6u/A/MvZZK/L82heX6OUR
K/bLyOvywfw/tdQ+AS8A+/ZMBYXHAODheXWjMI26IO8NBzl6xqEokRrh2UC6FhIl
scfmCNs2Sr1SRk7oUJFPLlarMLvIN/SmV6J27wpze0MfX/kPla4gChbyiMohQVIr
n5OaH+pw1815RvKi/CwxdwAXqvNKgQggVpyybJy80hyhjkzEoPxHEj50l2Ou9S8Z
0oC/tNaJYGOGOJNHqwU+TzW+PMAxyipxe9xLa5argOLUa+P3q/GjqHnoEBjO8G3v
vDeqzAclPcx85mT4npkIjHYVD7gHPucfu2c7lNPWKFk49qGXd54B1rLeg2qDfyE0
hmDXGYfn2URADeCPCC5kenmsHSXkmA2sJkM0pYvbezF6l2j2DOMpVIEMfRegCC2d
/0GtyofCf8DHlub38BX1toN9iy42b4Oa5ZK3oocoZpwArLyJBivtupz9sYoonD43
gvwcrqBCEJtmHKLQeiBDgfS/a7cdA+71fdwanQmcYVue5RWU5YZ3aev1N9DEjudy
f55koW9WXLeMiq9zNEOK1SyANyrVrzgJldIvGlPIT5FxWlVOGFDRCyFV/Ga23Rnm
93LKNt/GjhPgnH2O08L0/JkneLxJxO3m6/3malfvAThhHDshyaNSNEvodSeB8O9+
Lqu3GOCweupfhhsCu109LMt9lZM9euYfM94jAnbDbN4D8CIhKdwIXaQhmHTpiNar
kq5/iOFFKXb1emB3RWbi9tADzZgmVnMSD06EBS1IOzaPX/TIQhpv05ppxlTGnJH1
OEAI7En3E8sblX0djNK5X/9DM6094G5PK4aOZL4KhKqiq9tycnJIvyEldc4bwTMJ
Ix+aa3nNIXwD03ylyFR6h3w/00/nDk7T7GjCOul/6oXWbzloEuS04rzKAWhwr6Jl
C6aE0tCyKSq3pkyNlVNMRVhpCLT5MhAtekwKeo39ekU8/4SD1VAE+DOndSoxzz5w
2xtmKlkE4SMeDNeAt+iKuAe0JD/pncOYpugFkF0ynkDBE2/KhvjNO0RxyolDpwR7
33FVwmbVUqZC5XhDPXFpWAqQWTCwLJmp18JG85KaRli2Q2iOabODj1SM/Q5U/2kB
8Rsv+H3xOfddhEt4hRRO3ifVei91nnxFQZPca4LrSng3zgaJti8tAIY6cvXsDMtP
SJfEIAHl3BvrY4pd3q9Nap2AEZcB4CzsRO7VubFyQrX41IqIdxi+rWmmL5R5TjjL
Vkmy5MfykWcclSbBYGwNlZE5Ka+gvgNIFckpPQAaTnAPOjWx/apG9FwZanXZpG6J
UotFtw0xFC/QjvrRpKXG8GDEyG4bfb/dthBgC6bs17VR09x03EQTFyXTvxioISdk
AodIwhJ31DCSE/0S05AYAj9ph9IzO2yxOxaZrM58ZYdnXw61OIXYR0rQKP8LiaM9
HV5Tess7QTu/YwB8mYeCXDGLTccQglvhLeE2J03fIdej/VIj8AhYrRsI8bXztiLC
FImFYeVilPydnL9qW6jyR8eI1LC0Yl0rBWTFsQqGNifn0X7N0PxLJCO2kxR/NDJS
0HxcFCklX6BfZK4LwqBhmca7BUWytd/oTIVY7yEzeTRiCcIb4V42J7XtG+OdJGIi
os5nvXG1qMPG0SB6Lc1SFCdVgiNWumjpk8AYcJAcmrRFIjWenfJ7ikP8NTjtDxhO
SdlA1G6dg4gSfQ4gT+PPLj7yFUWxs0Br1AslK52Fi7l3L+MoXj82smURWeCbycSA
u//K9SSKOOr73n4LtijODZwTyeXOSzqr3JJIJrIjEwcaoj+eR61MoBfRoOzCGtXj
+/rWwNEFGH5GwDIMgelwyCjQzQW1BxQk3ugyP8btWVbTV6i678wIfe8BPsifit+Q
mClDbtHiNMT1xntLRLjCzi8VDn6yubfvmgQFXxfrvDTu9ATIHR6Bi/MkmupVdkpn
oLjaNQDu++rse5JGDr6GuWwrx2/EYs4mvhMLUCPMhVz2Tki2Kh6QTkXFH1ISUcW7
4uqFF8hoONtDZrorQdMCZhdxglHZas5+g0zLJnuTFY65ojK3hE8N5DgwPOsat4Hc
vRniiThDxdIImej82Ia7FYabrDELcUOefAaRwaqrDh7/+xfZcLAzZ3QiXxkdqiz+
eDgnKT1hJXmfEDV3MDVLB/dU8xgtTaeE4H4Hw4Ej2q0wW8Xu5EsrEWg3Qfvidu5R
Qtdq65v0Rg7l8L+MxzeBdjPiJr/GD3oZ/Kl3m3yfb0ozAu6Jg6eiDn7EqQ295anP
kWk97EGhrDmvKShO7czUrE+pFtmQtZD+33lV8+ogN57YSm+F65xwq67OK21Jv14V
UbEiU0sdQ1JwTEBppn0WZiBrkveFpDz8oEq4d1mtac58+TVQULE3g+goIDl8El7i
a+0JkGCR1gL/3xSdVb0ETBFxVCYhIm36VDtFAIlSl6Zxyx44K6rplJpdlYyFBSFF
P0eHQMO/mZxFy26084P0GxbeBBiMkLKKO5iPUNg1BXTnabR+tVy22ljfG/nEPcHl
8U03Rf+9qYcu9N9Gfa8mThb2Kd6oZUBmC90wTUw44boiRCoRExUF3GlEJck/H9NA
jv9/xhOWqlrnSxrmpFgG4cv8MbD8kTHS6Ub3vSA2ZDqOaNvmBvThd8Ffri2zHbqa
KfdrO3RlRs8/xxk7kIsigl24zwphkOjN7Rm+AF9G/9dAqIL/lbKLhutRTKFq0uKE
keiFpBZ1W4vV1gNdxcy/ZMRG0mGU6Sj98M8MDdYAG78oNURZdCRd7Jd4MzGTL1fw
nTySdRrnEE0Kbxwh2YMjSt8e9+9tSiQ6INUFCJXwRknJnWob+wtn3ZBjTKfZBM23
tbLPsqrcENPAB/8AbLiX42aen4fTl/RbyKMviEvEQlI6OIFtUUxYl+uJKHXAJZiA
FHXiQuzAhnMuVruEOFqYjqqnmJN25AkWnN3RM+aPhPhTuUOEYm5mP1EXbcS0bHNs
1gdtzas8S5yr5zQKvdqhHwnYNK4tfwnf/qdFX/EC7i3DHqHRpfrE+1KCcgKIEM9w
VYL6xUwTNzY2RFP9o7CPpHpNoBeyNVjK2OpeM1Zhl/tVCSsMBPtmjK2kjREGyQbY
Zs2ND0wznHtsKdEFeqrB7HMYPUtZFw7+3mL3q4dN1beR4H4akK2yxDKWPYa1sUEC
TPrsWF4rkeDSuE/AhTuuUmDk2n/U1dL2xfwLNW/S3j1XN09WVgX0aVRQybBrbx+m
ZinuA02b2CSZ3ybBZxU+OpNwa9mYA7iT77FtajsSNKUK7BW18euKHkUNxTcPExEh
OGFkkDuYfDOiYIqdu4DMoAMhlUKSCx2UeYZkPCpE558/tsQkAEtStshtqPDkPgIg
iXEZHBIn3gP0B3GXzRcINvHcgjjdWFEwEMb9XBkQWvWAWaGdhKVlxeqVQExiwxAK
9/MSNJF9a+EPS+dpcmoAJBt9wcnW0lyIs5TnwarodDI346l3wwGPLAlFdJdUz8bc
RGuuNr98AuRtLWCNL94LDJv/LuujpomrccIlb9XTjd5Cc/y1K66fnbsvynKjJgnh
ddHlKdaT4l9iCi/K9CX8EiQBayK7pXZi/G4DHnB+SI2Rop9hDZqskbHvlGfScRoQ
Wq/2snBT/azip15ITqGFvQf5RhSmRC4PFBiXq1AVGJgcwyOa9cUGZQtqaYHT6K95
CuU0pK08jIIbhE4v6Zv856JJyZtpOfDdtvXuEegZ/IbfYYOF/p/gKSNnfcu22C74
4+D6QWLLOUN1R4PGjZl2nTlePu8YHmwG30I8mUeJAazjdhOmwqjEs9qHzvKw5YTz
k8oRKhcb6NKMvAIdPEL9PUjfDKSViMNz88Gqb0whlPy3vz8aqs7+3tBExtPjbt/c
ooGDVCikqWaXbEmMrJh9BPvv/XbeNQOuy3mUDEt1Gczc2okv7x80y1i1o4yCSrBI
fmeeKjcvBO4cHxwF7/V7BHlOxxdFJyOLVOJQyeXlZsjDm+gH4QPiS4dqhy3D1/pL
GyKL7nm5yEmyt3cotf7U0/9eH001SgFrnFbq0x10VQ8WK5TbvED0YDeTbyB8rGEn
nUScP1/4ZBc5a7K/bSZfyPKURnfBpcg4ORD4jGL08JQgWSZ7ILWK8osr2ox3d6Ek
kKU7sfLQOd87KqXdd9kuKUe3GD90Gde4Tq2eDMwUdZVjNwvtieJDk+RgHe1DF458
wkee9xCocnssOS8s2J0hw6TwclSb/QScSvDiZiwULuCS0oEsLc4WgUplyOV+AxwM
1lCzHT1LnI6RKVvatC+W1ZPfDL8nEShCF5I0B2ijpTstdveMmh5M79G5n5mhfpDE
kD/uh9rL8AEZCSLsECjOH69mT2Bh7E1uVVmAMHIuH9SWsrrx/EIKRhaPCMKsgrpm
voESiM2tfxuMtn1S6Zx9PgLj53K2wv9L8bdi6sajbp2vu78ViyZ8wlFDxDVQ9flk
p4ksXEUGbxY4EGwyovwqeceaNoakhvXyFyo0bAPizhYD2EQM+uHjWgTAHgc0XKda
Pj/C9+DZxbzSE29bV+uBH6rsAQnBSRekWRQpszBnAtOEE6xBO4Z3lcsWQSg8asPU
WNorDH0U1pYqQIQJCds9tvAEQvL3jcsaYH29u+12yOYN9NvhZeKkpAyIoU0fFOla
PCjlz5YopTbOCxJVyLcMA3Waa6pIAm1wF8m5VcuPKZVBbUbMb0zFks5PYH+6vdVa
cDw19snIZfdRR0xCLIIQa4aRB0I1ZXHzjD0l2L5OrNXXRkeNdj0dB0DHe5gQyisC
c/SXRzGA58KpjhN8lPc2lU7rgJHuTes297Co1gMKr5Rnwj59jK3A2TqKRTkng0r1
7rSXgHF0WpWfJybYGmctHHVAGGwafZJVEiwch7iRi0HPOrQnIYthfKZ7zslL5R+e
4wXVTh3rRM4BpWGrVeZA9I1h186mSPZyoNpfwR5yskKZOMeUPRnsQfbcKMFa+Yzp
xZ35aYCxJX+I39gERzOXRlkkeMAnzXvhRHoKC5lnugLiQ3J1je0iiI07dudsVfw8
NO9KLktTvY5uvuPYlr7jePhD2cCMfK7YbTLDkn+CBsOhAZH4I8nq+x/lE48CyUnk
TPjTXpaH58R8EJd13WqUbR0SpkDo3wYzH4Hbnz0+BRTJ59LooCbA/POiYSfyKmVR
cAsaYG6RY5ETV8Q5kV9KuTcAmugdaCeVUws0mkgywDnfVZD4NfPQj9UPrM0SUJRB
DxEEr6L/PvQabUcO3lYQyRU1p9C9+CUi8JpOpJH/YzTuoK32BmO4KHjwYiDDZ9g+
TXUuzJCy6rR2S/mFQGIG8WbFj1qLBa13jPLviT+4JmiOEwUgxozluAzmodEPPj+0
AI0LMV8Sa7MSk6PjmOOmXsoFQI6Gagopjdje1oAxl/ioHTIe9KrMqE5CzQnHGWTZ
jdq320dkxq2Q4nKitwyVd89fJu1ev/Ev5CnK9V361a/osbzaBlXfsOB8xGnG0Q3h
eRPB+lAoggarj4NputEW9fFl6ZEweKMr++gxlPS4vwrpDrbf8fa8ieWUBSsuWn1/
T6V5YqfkNWEYvfaVhJ7+NEUCyefXJrKjmjNm+9C275TVomkw8bTPO7Q9oV5MWa4+
xdVu+QLW2wbM+9T454YXFdbdrvqApJ/oE7TZyQXeKColpK+QBWLZWa1LUt1mckwi
bSRro+e9ms9A+gNDP4YLV1m9RZRzjkXN6laAl8WDVf/MbjqiDMmKylj2CWqd8oFd
q/ueuTlXA0gTDtt1la6bdn+ExmlGyJYnOQkUv2es3pTRoGpUnLb/pGnov2UDgjF0
NpGcsISuUEU0dzg+0MNECbsNSnjDO04MGtVj7XIJUqEzgYlaIc5/JpCuVekLzf/T
LaENnHnTydqgF5qYQcuYjMTz5pZMMvJFUrR2W4zkl0Sq7Cz9SRoXtJuAANJ42ixf
S+20BkICokWDbkZlcgoou+nS0aU3y30L1rDHPj9WRnIKUVYtHTGh+i/cHG6mKiq+
5dTMnFAnUpUeaK2GsDkIvyhie88rbgUSXFhRXgQ6lKaXOrC3jvH65CTVFInKN5I+
EI9JdWlmhfBhDxVb5ltgPGsa/qmJ0Nb9wJYY/TtgWpqMqpOBf8iShnBAlE6K0dqQ
b3tYTvDX7hslZWc/ZWatPNuh9mAOI3XyM7w3AQVj91Bj97qktbRYLUNOxD4NfM3l
kpN0/2/Zl8nuYVIoEpGsdldNpr/gBDG9IUgXubQpcxgXPAQmYyvZYcJANXhvAGVM
xcE2dSX4B3xAznufD0bsuxcNvHhn4VsakjOPNg6Vz0Rok2R4ayDsMEm6Ms8J2sVy
l402IVlwQ9K38kfivaq3pD84GegaLraCY5rzPnoNrFgJvmC2ytdh7hQCehvX0I+U
U26yeaj6C6B5djhFI1KpxjGK10adMqg+B7G7v86yQ/WDir+LSVravbilHrYYdkl8
tnyYqYq+e6CvmdxkW7p5x0KGzPUs4mRyth6XQQNKNtZ1BzhRO/0JPYjLQAoUju0E
3acK2FhIZCC0vDhpwSwxJOSUwgmxJUrPTUArIwlF9jA3KX5bZSueNZfbSdZJlVWe
0eiAl607K97Oe9t1HPhPjmtbCg/Na0bZ4giFhjzU0luqkQ5JTywlZSifLkXATtg6
QVupQZJmZ1RnmcRGazigojz1WKHfzNXiXMFBBcwny7EdYQiiDfPiLI5wcA27H0xh
G8/pdS8bT2FMVwFkkTqBBWE9byU3cxxCLHlhadO9AIMxftoOxdGEJ4ZwBaMcg51n
BYO4Q4ily/SdgVGJZloT4kakD7GFD+V0DEXlb8bEbAV5kKKL4G+4hczJeTzXJzi8
X8PPMHd+9OaoFeAvXYDCH6kHGas9V78I54rWY+gDK1YJipuMeavMhun3oMeOSCQb
kLeOD8Ms/rYe2BMh7GbuxfZqz6obIs1sReMUt+c/rd/R1U22NWJeLN7el+UG4iV/
dLtGU8dIKM+zCogIrs8853HOpoBCzvKFI8TjqKNr8UoP22hMS3NItTonmicVq6uZ
iTomXSLlaDkTLCx5Pp4Inn/nltmcx85iknvH6ys5LIhrYgKcDj+eVgE5HZF1FR2R
EfMDH3VjGSuSgcYO/xQsgMYjkFH9JxdsIlbNDjJ4RtKi5wZiCJrK+4ctaMJlL9Ar
ZhyurHVQ0ixa0hVn2Z3wYeI/RSV0ZhlfY1uIuKJHhL2rqXKPsaHK2hFL8G++USr1
KV/SCN2dXoTKFKsNCipQNY/pI3bUGbZGjOvAfBkGGYkBR73aRoE+o1hhb/QMinl7
zUC9OFjCpGbthPNud3TpIMhjG1WtKm5seAC0FQHhx8rahrHxW80FdT/v1PkOLrbb
ZyFpScEfaRHRt6p2OCygYYNTG5IHNSgekE227RNbiR0x3SqesD7lHdsjXfduZJAo
GT0knjT6fVeGbWy5+t1/bRnO7NTzDimXCpP1/kJNT+Je1+jPB41q1iOFxcquIz/b
3JhIDFtl+0G+Y6m/B0Cv7jbR0G6l6l3BgFj5G/X1Cay6hn3yOWdhC/isMi/TE9mt
ECZcY2yr5+3F3LZxFu6w/cZ4qF0+pqkl8FZxe4qCy6m8+dq0QNQMnMDCe7N+Wzvy
cmHNqwslMKby4uRKZmzsFWL+ife6kGKbbPj+oohvcmubTVT6FDOcSMLPdOFSzZHT
Z3i+mAPb8Jod3t3FWNDAPQGsWOdot+j9FkUQ6ji3ZryTtjoaClDlhOQXZjdsG/6f
ucC/OUcaaWZ7mNy7VAa+eqyDTSREzj6DYlUiVNPeLY2YpxPKSsFNGjmDmf+nCOMD
h498WoO8ek7mEJjbVchqGkNPFVdGqwVUD9JwWdy6DZFoMzDs4zY1ZXexp4i2+B4i
Ax3sn2Wks2U1O2f65lJJUeP/s4hAX0S5NZkDwNSpZi7ZrmQDubR7wQ/oPnCSPqLg
qlQO7kd/h30ZeYvzltXKJPzFpLtLSugYsJedw1ZkZ03FJ7T5FQPSlyif8ITR+FRr
GKxRzP85AmyUTs5w7r9D3Y0Q4Y4OdZx9aqq5NYWvMjUPLhAvH3rZrn9rPoHVyU5Z
eAFBSJE1vyfs73sBqr/+YyazrMrkbfEVdNEk07kvNvbSWJxM+83/ZverE3nWdBs2
UWzwD1HYEWVElvF6DJSP+4wT9gWPZY9OC/cV0ixcFkXH+Uzovo877QqAB1KxGItE
H4UWfjgdGlK/083SD18r7F5N/fhpV34BKgaDCohIChSj2AvL2Tgi8BDcw/ZhIgN4
Ncmj7IIqw1LV4Nd7OzE52qYWtDDi77P9rXYh09cnL1+tAKntBnVTK8UEcDhnIa3E
XhZaqTaMUBqbZ25EW1I/o7/RxLxbqvQq6TQy4hcP5DwcDfj3iWuEFiyApKqb8Lx7
o3aRbqbDVWwu7PYG0OiwHyErrOlpXUrgznmwDcoHo+J7pC9JkHPc31gIWB/7yPwe
/aRit5CpwZraxrdGqlGDHFXiZ04sVZ3GQ2zOHlesg8OZC+WZ+JTfoHSOYJ5Tki4O
s9n83wM/rBtMkUU4LS6XUU7Lsr0Opj88Xi7TgEW1lWTIRTORumo6GNb2nAo5dsoE
PSssVe7GlBSXo+XJM9ked041ijqeUTBd2D2A1sdyqXm1SOlLjBOE3WYdVSD15XWF
6pEu5EcODU0KRlUvllTLAOvwc5Ew++77bDZ1uUv/3uk95Vj1fSfmd9FvT9KHKUdJ
3iPNBcpy2qVmiBotQ7vnu5Qy5VyoXKx5NOoocu/niznUNViL9jnRWYuVg8OtryNB
U+4jwekJGi9bLPHzifGkgrgJbPidrlfWKLAAsPwCIL6rIOKAkpPK0SVpL2VGIxTo
xc2f3VwqtzIxBsYy01FDviOdQHXgWpvJcQJ1DHbHR18Cw6dy7qFszLqgGE4m6h4E
BnY4TeQpe3S9WjfeGDBdZct4RmmXTK2X6pp1StWwzMZcM1SdHn/uwayLRXfoGSAw
r8LbsGfjoJsVkOUgclAIwrs0gIG0n0/wIjTFE/PBv+zNBPgirE1TiNeIcEGA1129
LL1pHlQ8IMLh5zfqgLJuLEwvLQ2IXrO2uLu6LHjnMFUSOcMloBU0si2IBTYOOSRp
szoXcnDaxyOZxeu8EMPXGOajFPSQWOOb5OYPj7+SvM1JmDtS3SR+hjxUkXla1i+r
UAxfsduw0dultIyoiBek1zEf3oklR4uG0dXxNktvL3BVranA/Suw9u4+1PpQBtAo
Xy3EyCYy4vdCyRaxpxxfXPwg1+yetTHGHTWOxIjOiTBcNrhjwBIkhs10OKABao1T
D0sPBOIJ4jmI0MG+EMprgcJVE18k0LElBLxza5OwLiS0a+1mxHqSt+gqc+jBsvNf
jhq4hMOPcy/SMdoGHduxUxsmC7kvs5hWzCS7OR+q/9o/aFpND9jyUb5E35Kfyrl8
e9cibmg7fo0LliKnvlySZV9VCpPGjGV2y3anzjaav7UUD/vIGP977Lz8/3RAOIkZ
ra5iNQHtu5eqcKz4HAndoNvqHZVRXWllzyXlP0ArErWOnnvdPNS9zupv/lRXbSVB
ohBiDAlYfV1jfttIdJ2BY/QSJo+N3kOZIhNnppJ9Jk450COjKI9l3CGUh/kLVlkN
/+Iy5JX8Rv63JdZFx3fyP7zCnxk4kVyqMvk9nb0QyGD2bcJN6eABMT3s3ku4DnPP
vqP5ojkxNjwSNyJ7iHvFLD/11Kaf3XyA/mhQibBampLy0Sq+teS7XU8VgxSVNbCr
VIt70ESF9hKsYkRj/Maw/9/jaG+4YjCeYs7iUBvX77rsTvnW4QaJqy7q9SH7C1BD
KXg8sYwIPEQqgJ9I0KwYWFAgoZJNZJDkaa7PXgOkOCErR2xG4bXSEmHsH4lqPPfW
ck3AzP/bn99qEubu5MsUt7oE/YrNtih3kWY6zwGxaz2rPayud2s92IULxsLXa5HQ
5TGT49opGHvjS7LqDOx3RTMpOJXOoc9luUIw33fK4rwzbqoeBNmZmXtb5oAtOijr
lK5oaswq9hanx33JDFYZnPzTGx7FlyIK+yaymSvuwS746AIBiAxyH0lKYRXMRNDU
QmZ3L3o7gns2IY44x9Dm9q9ndVnZt60Za7eQ7StrIqz4yw2fLUjnN/oClFj7B99q
6xWgEVLZFbifaEcBwVR/lYh4Lpjrf+Rc+IqnGt8gcedudKGyqVws0SqCXy+Tzhe6
JEcZbP3ktuhwPP4lCSOlCu9HWEg6kwrz5vOti9so07L3aShIgFP3skTF1KZnXJKe
rUsG5L5py+a2qUVTmtFIBMZWObLzrGXcLy0E2FCIZg//8G7Rbr/SCC79joZV/+mQ
Eb4YY4zvX8hFJgRu3NZZ9SpsvVgUQj/ywoI7JubzgI77awAObWIBZC23PM3zbwkL
XwV45k70uMyAI6hskqUV4sE3pFGIalFflRJ5WZi44fprYVLu0ifLdUCR3GClfbfg
vkwMACeGePBIxX4N6T7rYbT8jR3nkpL2tX850OIScm0NfJ9r0z10bWirP1riyzXP
MAtdXcnLF13SPjH1+bywVuZWKUs7FCJ20q0x/oVISc1dwjVlj32mudUyKS0cJfML
X8UAptMe47iQDTWscIe6Z2JuTAS7J5atD08d5UImgr2HaBXVN4qVse1xVD+Z7/JV
Y9o8zTAtKWZLSQ0HzjgrAFdCs3RkmxpZkgickcM7Tt5V7o9R+0aygEClNB7cjIDF
1CIZVClCpyHC2BbGrnw8AgFbiQqky1+mhiZZYd5vgwUO2YL4xcsu1zNQeiKmvOLy
lcGHIXeqkx6xfK6RJ/KMsSAjbJtKxEPhQCz/xgj//24OxQuJTCoRha0lqKeFrzBf
iGxbUThnkD4xBWsYa4QubZCmV9TWRVSYOGkIJ40tYal/lgomtc67YzfLsSkrKC2l
fWNA1vaU+1AOfdh6t5/wQsI+7enEoM5ywdJoA0OR78aC8nSUlvkOgG8a+LyiSOWy
TpDPSpKg8lyYOTKqrwYBixWNkitwZsrqE3kIgmCiN2o2ldt/YBuE1EZAwYDbfSrx
qxK/SJT0uD/gxmfGvwwM4U6cZLr0CL1WUJQmdOAGX6WgjilZ1yrPGoZ0Vswor1j7
AZdKTk8Bvd+PJbkQwq94nb9INc6gxR13eCIi4EYLIqMLwosJ7IfJ9ifJ0L2DD5vm
zHAvJ6jQc5ILd30KHaVPhvJGmjk/zPJmRd50XgWWQhkSNIlPJaxGLOtRSOai7q7m
g/DQ7EBso7MCz6C/D3f3hFPnNMJHVaNHwc9sCiCQGh3wFECZNHWrZXs6rntazgtI
pFvtyWclBpzXn6++SDIj/fV/fkPqryWQvltwbx2Q2EqCrc/iY/UTLGDQT0yl5Vri
2t/88b7ajLx95AAYiss6SEDLGraMl4j0HVjJ3NyfzV9UrLBQ7McclZ0f6RVsAgry
t7tTLdd0lj3u8u/OTPBetbHbHu/AeNK6d64laovQm8xL7jr0wpLSYsOF8Y7Nkvg9
OXNwC2pUNHh7D/tZ1K2FrIGwfTFS7YUuneVNSCw7TGsjka9/RuOTsm8FAEMOPg/c
BLS2YbLYl/C10Q/4RigW+Pf3e3v1y1ZIRHuHszKbsxXKizwAAD+V1ONkBUZDry9d
sTFUgFLNXPlhcpMpKXu4y3St8t1r/VQ3bPUarKhROFbpDLtcerkMRzIza0D/J1BC
1gZAxoCSK9QY7lRxTDcPuh9D7LVjlY8O+W/7rKZQUXpQrDRTnktuKuF+hiEVID0V
TXDrsuRuK2tSKgXr+q8WBLlt1Ju7H2GQaEG0Q64tSY+vJvrghTZEaaaAuETOwm+r
wjRp2aqWynvPuh+fOQLpWq4CteAa2WHvZNDdi2jQJxq0UMuogG2aqi7zWqRZanP7
lBwg20rnz/xjuOa9ugNiBaRXuuekoEfv56Snjdq/SOwzFe9yrFURKBY54F6FyFwo
vF+78WIJ8nnrzKF0wwWfvBqm8b/h5/WjG+GgjM0CmKVRFTdJRcGNmhJ4sN6eXBCW
zPiHlS1e8SDGHRrzqyYBD9Vt2i4U8t+5ja/Nx+NEQE7hRuICr9YiXsTYXcgx3m8U
klhiCykXwRcfutJBFhY39p3sZiIuozn2BCjfUc4ogVV3KY+SiUDWcTW+XR0A6mLS
C2M7NTgStQT7VrwWKyWXEWvWfAiWP0AJ/oaPjUlAdd530Ah2ClNiPGHJmwBkXC9W
NsxB/KoGs2tues5oFbyoxrcgzaC6aOR9Ptuui7tAK6r3LE+IIfh0O5hjKGFJnwTh
FIUlLb97B4ZUrOJaHvL9z9SEJLBDykWI1zyDe2AQbUJaPNGSNBLQfbwD/GlLspyz
4QjcEKVfbDbEUon8Uh5PGhDKLzr2t5bhvefgUYwS1riV+lg3xNEEUzMk+gcZRg0L
rPX39LXWmKNlg2DJQyv81vVKFQfGuZ3kg/ineSPx4WihUe7pFd09xc16p41HEz/s
Fml9Z5itPeFQAxYSILT5fo4Z5MuiX+H6l1EdKOhr36Ovv6gNESoM6FPZWderguJ6
Ulf+16l8grO77F16CKZVVuzoj10nxSQAc+eWS14nQLPHtydbtBnQ7ioEB9JEwWzg
Tcy8Id/Bh2DU6PuMqYUHn+lUa1hqm2gKzHsJUaul/YSE1uw3IejL5a1AYFtdaV7c
jRxmBnOYm5c2l4ZLm/NPqRoDctIO7l4Ynha9hI0Z3pnYcM59oOk8akDSwc6GnbAl
rPoK5FALtDFk23+RdNa9Z3820GNoZvkWI8OLu2ukVhrQdLWHOEMcUlq5Fazj5RYi
3Ks1hVAMifZqiDJp8hqbUbQJ0G3Rgwl2MUvEpI0xRk0X3KcTDNcOts1xQGOadkeO
mZwGRlDurjeVhanwZbMEQfP6z+PBn036Ajf4f7v9POW21sUet2D7I1bLpWobAdQA
JcgzbH1ZA/3XGlSA62UlKeSargwss1h4AIl19byt7MAzDD5k1r1rKmHLo993csbz
atq3zCPoz1wOj9976PJxcl8o8YE9jpG+Bd/ycFEqvifiAFBK7ZgTaT18WetZGO/P
nEpW25xikOUr1jS9xv4rI1AmW/OqmByClOeyaoRZyFAHBjY2eIAOcdLPM/jQzHPZ
Fb99QJfADYXSMx01yVuCXXSjTExQtLt2LFmTJqN+w50D3bZp02qGrlvYKZD0tsHh
2i6p5onuneLAFr+u2ux/T9wuCqLOf3BX7stE10y96dLAyxBqTgp5XYgU9aaKih3e
lNXxLKHMkvD2lkAepvqM7Hy3DXXtfdvjj8zOBYYnm2AXvU05x6dKVVau/h6+ZL2O
ZaIIRfHgcnlGvxqILFfR2zBjoD8M9AbpEnnzZ6FuYU6KbPa+lfpD/J4VniXgRKUB
cA3Vl8t/N7t4jU84uWHMMOBQSQtU+SAE4uPVOMGMvYo7A+UP6owKAy0XqvC3G1P7
OKZ7EwV/OZ6wYpAS2ViCTEM3fbq7lzzWxHQf81EgCzkJiVLda13Shw9m8roTUgX+
2HHnGurovug7X5bLk6b0UyNQ8bBiBjvL5lKBW4SnvNnbvATSxJrE9P0azh607o2D
RTjxgWYn7PfL8wL+igpMqCmD2LaHNuSrfIV+Y1ucaVK3xygle8yTzKlhFc9TRSAd
vnI73AREUydS+wTponlkKRFngTGCeau+hZNYqAuSE/nyf7VsvyrSO/7Mz4mJAnOu
LKFX9CIb6lwpDRvo/IA9t2DtmxXul89BN+W1uSf9wTyWucVfbtLF0xlTKB+yoLlf
MYlsBQqfFlN9PXsxpVgyjT1GcCY7pBznbTVW45gSEmUaN6sZhUEYX9OIUveFtw+8
JrvJp/tiXviSyX0eF7rm85llQRiakLybqO7NS8VkJtLforI52Z47tdgIuyKfascC
91edkvqOpA7uXNVS+sxojxrYMwETUMZfFNs0CmJmIhu8uRtLFYCNXoub+MyS1cJT
DjvnjQq4pNg5snQ8Gb96QZEO7LnhqXCrSMNAC3frMAmqdt04Q7a9PyibCeVttmYL
y/Rjz/Jad9EK57aTTJ2gxzdE13JLtKutHiMuObggTyW0nIYxD+PEAkjGiQ7tSADe
4IQY7TjAnBIhPy0NKKthOQg2J/QZz2iQON7cRvIHcB22+qEZSa5MPvROxG1gX98E
tIPS+jCfwvxK6eDzSIlkA1HstEdOj5ofjjq2hHNS1FqmfsdeQiM0hD2zkxlJMzr0
mFpO9dlFF/c7g5Ur6luE+M9jEiIAEvMMFMy3OikuPogzZp/mEcEgVOkvvekG1A6q
ME4KZZ97WHu4dh4LW3gCR40pMPyUg7as1FEq4TWkVgIMqTS4H295iOTJPdZjwBYt
/xqf18v09G+vv/bk67EZbMtfrfiqyIlUbjIcBY4mGzyWmt5y6DB7QrU1KYtE7URw
N+5MayElXAi54H+kS721kuIxqPVz00fWO9sO45Bf2BcpR1zK6S2bJgKV3F5bavT5
mJ5CNnoZk+qSLB1RD2deA7YYcbjHx/RPq9WCTl0ySKTS2DlTF3Ns1KqouMpR9Pww
G/N0rKB+oUC6hkE5om0MeL2BbynFOXLmiE7FyPcPEIvvx/8m3weWIEk+H7hb74Bl
cnNkcWGP3NBxD6uCdixedhRa3VhqrMYD7GKC3NdxRvJK8B1BU3gYJRxBj4sPY3qK
5J7vGZRB0X1pqfcpPAiUcwrx0IRBmIR8F2QxHKKNBct2ed0dDk3c8Uw1INFQa3bw
7ESklK/xX0YM36XjfwBrxXmlqSWvsLv7YDrRkCm3sRkl8u1UHR8AsDsclmUOxFLy
u/D0hXdfveFg9bZOZW3iNYJn8X6G4TyDYmkKUa+Lug+tIBgLyuOjrg+HynoMJgaT
mzgQkIGuHOqrgocnTbyHm4HNN3QTnLnJdTbtIkxXA2T9o59SH5ZpMeRQOuRbGHji
/S7u5w/rZt6TCJ4pHkZQ8o7F0XYZAzzgcZnGon4h5lf/XupO0Vp9yIvw/X6TgIb0
nYP31bgdDoBPoUV3PTzuxndFzqW3yHZiH8bFvRSQd83oLeQ4nlBjhg5i5ZGWTSzl
6Zb8s8QoNqXHg/b6wHLfUhmRgLsmz+dvF5Tw5NMq11QO1JuF429EvDcGwHtbQI4w
+vO8Emi64x5Oip8ENTUUZaOpxaca91S/pq3dkXtWedlLBPl0at+RB4OV7rPDyeU/
cpdERhFg6aeK3VeErLfClmvT3KxPf7ie1iVNEjuQmXqQKrQfQD51i5jiemNVfcbI
9vR2Arx7c1+0p8f8FfhWZ7mrajc2QzrPPCKmrf5SrakTSbFIATjdn9b6IIjTvMd8
ZsXqkvNlj9bEP/TwfIVaHhI8Q/Mi3MIuAt93iSlyVUjb7uBzgaVmFQS1+Z0Oa6Oz
9VOw0n0C2RGZACwLlI8s0RNbvUMOCCzj/5Um7HhfcuB/7koLlSK3jbxO7Az2s7XN
xr+Bohm18cPRi8VhGgdvVA90YSfX/79Ig0WtU5P8Q0n12o/7TUEwfsrXOywzVIwH
dZvpeMvp5X1jHnbJmGQIPZTGzPC3SBXQmnwC8RIZayTpgkwSv+rJ9YyDFtuZafm4
hCKXH2bS94Y2wIaf9xGsWEWVDwGigcpJtXYt5m5AFBE4SjUyYQAAxooDiN9lfzpZ
g2Xp4DahxIKsaOjL+rYpL3v6KaLrGqvDwvIC03EtpxWevizgSR0z0fKAzMkZiOVS
1faGCkiY+hrM0syifTZ4ZG5CJniVTRSFoKSRQm4++nOmS+gWjZN3rOf9PKVu+aJF
mleFm7F5lG9oU9bM7VjVLxzli0QyOOu+OilDi5MAEarGUC63uYC0ujjumTi/Kcr+
3owXln/OLlegyvrYQmW5rZwpNvRtcv34kcakrQX1YG+TyOaRmULglFxOJsgbW10S
uz3WJmmM24McYK7KDyLN27MDQEgbDIzH+KfL6ixToPY6V3Bz8i3u1tdHx1F+rBgo
72Sn6/UrojoSl3GHOC5jOQ+KWz+wHmJloOO16yIggWf9K445rpyWV78Or9+A1LaO
ESkdO9fu7K0c4UQbK+RWHN0hxsS5C1RPlDZljgrZZq3syf206v6ZThyZWAjM/34M
h9/i5ryzGlLyiCGZy8WIfKeO+IarDri51eDdVxJVWBlp1BWbgj8W8EkCexRIOiQR
7HRiCFxE1E+AcFGmJ4whGWTQ8523GP44Vigv1cRtZ6DjLDaSFJEYUDtRPPR3ti1j
KJJW60AULtUr30CHprKka3FEsmNfYmv5OinrcyN9doxaDeoSM0hVqTNE0fAp2MME
inP8z39QhTx+geADtSdXLU1sD3ft+WCLN+8UoU6IcKqX9rxyr5LIIYddiQppU0Mi
i5YZFM5vGQvG8fazuZ7jO/o6oZ+OgLaMa90A3tsgA3F6pydsCsVZP/hI0bpMqUuE
/bjh4bWr9kqrahWaExTTLnEvh9Jn0m+NSJl25tE2qGIY0VDYzd/f9XgDrq2Xnxjn
LPEBIcznSsjl9QUjmrKS8CzX4TmxPBPn5Sjmg7uZ8xCPRDpIJimG5XTEuU/KpLK5
ULjPDLxu5sXxuYTn4MqpmrptvRSKpbCQNIZ1SPxkFEljRObxdZlY1pzfHopmbgfd
CwM5/tF8FshG9X3OyNKA7FD9GIP/INWNwuG6x0w7zjTf5i/vp2tE5OLX+1rqDoB7
asz64/qGiXohFBFrkSvJgAB4druZTVVZ0CIdMDdpu1OLvhyoCM8AIfADwSZ15nrk
lllItuDnGO+bXoLmaVu2Z+7qZJau8p6Q8JjbfDyyUl+HAsJ9cjDW9sy3iDsDdp8M
+FlX18ok4nu8WL/PRJ4/Ksp9ePhg6IZU5CkGPtrwE9DR8focNO4LZbJT3xO2g+ib
SYH4L/9JjMu4n8Z0j81KOTWeBal9kVBrWlx3loT/VoT8hHdLzM+JYsaJMiOrvhtx
BhtbXceWu0aU5InMCQQb7L+UrlSH5L1zQD/rI2vsJbaFjgUDzEu58Cob8whyYrdX
LI85qH5O5wAT5G6J9/fKxQGeQAZQ9fOTFn1sJ0L6qitPawTNMP7B4Ti8YIZaKYMa
6EnrMiSWw3oNaE08NIfEzDAQmcKZ4BNtONOoAY+T0FCuTxB/i+l3Bspt29jXYKXi
49ziXcvp1jBymCeRuPsogH9SnrQPd7SsmBS991/wg9TD/9FsOrR5Bt4kBWecaNHw
ob/tWr7hr+0NpY8OwytEJRVkNa2GlqibefuHo+0zHu+HhDuxc0wb6Gs+9LmoJdh7
NF+qnL1Jn85SuapbXtABwo9iirLfaJJTYbpc8gHsA2HmZeKTRDuoX8zsE4Vx1/cl
Yolvk9rQhm8ZKynrInw9X6YZ3+JBtTh/4lNWlrvGN6SoxLTG0iJuqz8rxAnO0yT+
vnBp4gwd9FSOZoCkqau/uWEXVvgXic58t6FqHjrVeghIsGLubZXZYyfJkMoiDkaX
bL0gJDpXPw8L58sR343wBElEYkZLDG/ia9+4hLuCWAhhiDbV7lsCbtbRzSz/NASw
G0SBqETvc/+dfVlCQkbr+UlpO9ogUfmRnfaaPN2iGs5vBrUghY8S/rsDgAtzVaXO
WKGRj23SU7KEkggW9q/jXCyBl5X6S/MrrrjAM1ktSO2pIKDf3yrJsXbwvKG5pDtn
O3ckBRud2Jh9sQOfaEAZdXmYUyb8Y5sjgqhhVMgEMxtiL6pFwz10k/NGu/ejFXvk
qdFPC1+Hf8AVblOkte+YCMU3JAfhlXj8ge+FqsxCaU8xKz30AxeiUOb+4v7/EhQm
leJJYgQlBfkKNi1KdyxBJOU+o28MkGGka7QbBszmiZEN+z+fpNnleBFEOVy0khRv
kJ+dvAP/KXJ5XndzOy3104gOBl4HQF8lDMI9kf3ZHTqnlwd5GS4tW4FCXlpwTHy8
zrbMj582hQFIXix25MiVs+nj1f7mmceDApGVKFgBi8h6YyoHq/t6IqUpBOTc8JNT
uogIJUgvas9259Rm6i8CWIGDsVwEdEoyuXQ0q8Vr0WWsVsnKl/kdwbpqV2Gg+7G0
K3ULCSg5pea6Q6Ij37Dmnes3eR+9LQ5l6qbL4EW0KjA9ntSwhwNCm7wm9nSf6HGh
+W+O4j9C9ZdE9cqiTjPvgzXmyLGKvxFDfHVTedcpUg0yFKAMeoP9meJkxRCRb+vS
ITJrfJQqLc5HpDM8heRdemPBzeroMHSt7EU8LvNr3M8acaWWIRvXEUgdV6OLbJvS
3niKJTQYhA1m51KHqzniB0WHgAs02ePGP9r+p/8B6XZgCNZj7v/9McjUBQG18CeE
FUT85d4nexAM5qcNeX6EGThT4ldkyDFmQgs5cT7fO6cIV2OayrzNFo6P96WTtpjO
18rmZD8+uQVmtR2c4Abn+l7150GL9pHVF+yihkRFuDMaYZU0kjdcNZpcdVtW7IGi
K72tv9YNRKlp4rsFLmrGcf2TvaUNY+RhJvm2/SdrFpAWJLgK+dqQpY2W4sqKJKDq
NAqbzmuG5hM5i/3b6Lb4DeFsL2KkZP3swBAoso+2rd2yjBrVwd7+0BtxGVo1Dl3b
k2778m2/rLqMXKqATkvkaE0J7L0ghN7yFALskwtw6r+bosmLTu87z9xEqKJh0/yz
3mTPue/FsRHjNs9bn8g6kfmli9NpBarvAEZbnZcsLnqrzP2XJQw+zYJMGAMEpRqz
F+pEzYsj8j2tfiM7E5/sAGFiU8sb4D/fsbVqFhvbwzpQYGbtEODmvrIdA4RSzm/c
7mAwrT+8jtt/xoPCJtebymTuzLvq53vfQcYUA/4FuMdJ5AZfw0QfezbtTvroI9OS
L7RtbUiyI2P7d1nj7bU93lyfry/wy0UTAFFzFvT1O5vUeA8Yq3hgTb1GhaB4i6Fm
o/510jKY98CRXdYeZ65zgpk+cUX4UWsLnqBMSdejx8PWofzCC3rcgSvj9LoLBVD7
PPBRE5d8VcnWNkNi1UHz2are/MjHteZPZmg3AYM9QWxKjhudhuzblrEMo0qBLHB7
Il0wv5JsZFz0jEXnPtZ9aAfxlhtexxAnevU+5E0Pvigs7yjjZd+eQEOI1q+PDzvM
9quUhGBdId1YsQGQuFLMbwqifwFlxsglNVUwE2mcvYiUVmeq6jKZDEFMRXxlvrX7
upcmG7BI5jpPhtjT3xhAH3n9bduaaoXtDiTq17ZqB6/auCsEcCnQFXCZeXt6mP2x
G1aRZn5VDM/V/n25l361mRecNZSShmWDlfQj6tuOhs12aE2if/dROcjq2TKe7XuI
VIKniWzTgCfKtVFzPyNdNET5kV759aggRvgmcNfjXI0sEOrF/ovFm+bN/W38oW4z
JZFBWfj6rC8iv1u5IrUwjPEMvSGdXJ00zOV/vULHOq6W1lxUo+CapSYbH8RCOS9t
NOv9RcEzq1Q8Sj+qehzPY+vQ7iSkkmt3GOI8pfcfTgbRrAgf21nh4luZ1xi/WqsJ
Yy999dxq2jKOUjXCeqSQwqHYtuh1qnrwtoQ0+RhZNh0cnKma4O0FfijlvMaHz/S3
R6RuMu7j4vRhua3Pp/EddTf/A7ymd06xGOcXee9pE6pGSiBji8SlAk3lCTgBTCUZ
8kbWvzZrYzhon2wggKOY62sWosxLtGvi7JSihShjKUzGAHDCyfrZgFp4KGI4mqoY
0gRPVtAYCx9dCV5gqeqm15d/T8VSQxOUiFuhRey/vAgcXC/xBBg1F9N4d5jowJpR
dX79AGr6RFqZLCJJPr9p/rKRZAsBvatvXVIh9X+8HSRBRpDC0s82GbZWCrLwi1s1
BRMecFsz3hmeQRl2cjDZy/6+HHO7ArQTKwuUxW0hcJGepoiDzB3I3Ex36VjXCDix
tyFZAQpYUA0Oby8e1+aA+bg0CuN3FmLVBqvCZyGf5c1uMZMABhsxNu8CV/1w+Hcz
5Jn9FDYAr/e9RvS/lHYWPrJMF/U2SzZD3ej4XS7JWDcCadnHtlb9hvCzUL+YtaIX
LW2hhIm9xvkCNa0VsaxU6fc2nkSwYMNHg/+CR34upcp/cktidlAU3wvrsf3YL+iE
+phRa0PzoILXMOgnyL6EZ9U/f4ZOeKqxOyBqLamCHqtIY7iOEJmRBf+MBdyRkjb3
x+HtoveC0/9eeNNwDLjpuxFHBNaoniX7z5fGlxIEoFvbN5XoGYSe7AG+0BDKhR/A
3JNhGDp5g7e2Dq9q53JzesMm4UOr2hlB6JMc6Hu7ixppJoa3CR4/MVrSHNlNgYnr
vMD5HrcMxf48z4M2Xh8e9Be9k5onJ7R3rRLR3+ZyZOqDF+607/pxwUdQoLH1OXBW
NDwuUDaboyhTgOt688u8p3ymjN502XFmo7Sny5X3vamLiueBFeQyRPyanxPTICt0
UbRsfR85F+QvRJx6h/xRfV2nFHWxAN1nbtgi4WSDXx6QZ5mZfBEK2OF00ZM12A/m
D33oU8nRkn6dyLdZyFvNbJVR9cluAdaIkyQxXh+U2vBW19e9DKSCACE6rKsMC129
G5jeLE0M0Vd8tNPD1Ar3tzkyVtBqnpIdUmm+UdCVuhOxz+JLMzzsi8wBp80kuYXO
Wwpwv+Q04pEsOB0RrE01nt5jK+NGPOmtYbu4nty62FD7ex7VIRwjDGcutW506oiR
E1OQQCatAVuY0Z8t+Rzqzo6aKjZ9VvsLcnMVOkDM9qS+y2exF1NTAYAWDViHqehn
vGI2mZQunfakSy4NVzKCD9mP7ZJsMDqLSzAxn/6PH8YdJuezcg5UTpnpUhM/B9DU
TXiIApgmRvGzQ9HFMKqLC8k6AsEuTeO6oR7d7uqJYAxVIxY03JoKTgdDiY6VMDTb
yHJSpRxj2LsBVHyCL0zj7vA6xLwDDZ7D4nHkkgHEvIcGuDlvijjl2Sv+QT5wG7Al
b8s9Gt/E9A/hZ9q3/0Sw3VsYGPReMtIIYqbwJjevx179y2lsknspw+mUe4XFjN6i
ABeXAn+rj1hYo44FVZuCANfRCqtPLzsuAxOUvdpxhhstAAqbzk/oIWkBZR7k7eLn
RVkR+W1+yBy7Iz8MwKa23gQE6KZlryR0udS/iLz8pdJgStlXEzmmGaTimWCGjqjc
0FXUPqXU0G/ulpJJRPC5PPi3/+9DNqX0gKgCHksHIZG8ZIa5a8GbyvcQzdmJWaDq
pH4Gw0CVDn8YoNNIs1WOs6N4joqdxkRWzxhGbE+8rZXmyhZBegeC22Vi+NxS7td0
DG54G+pOu7gS2jwpeH/nu6SdMI3S1+JMoVnhYL3ISx4YAEUPyuUuJIS/Viss/qQM
cB6fYjAWgqHLPJqJCXFeNJgBWoqnAD4Gypc5GVEiXhY40i4M05IIJeWYkYBCfDXg
bAnCjxdxz9P1v+GK8+bRO400u4bhvnXJBaSwH9RLFEPLH617O05RyfukvFPWWsNx
PNEUqivIDNCt0uJOagwrFZjI7RZB8SkWLSr0Yy++9yhx6tej5h+naIKJCOUMR9dq
rIVOfcAtyeMXk1Vy0DHpoTkl2CZsYz3yIQmREuw4N5Rg9mtwhKk0oxKtPO4WgTlW
BeX6+5LvdToLZqfPyJJHVhEuICYrwkd4wi2L8UVGmCgKZ2KWVtg7jXNwprgZa95t
ZVHDIZqvgNVEQTFbRDIYPvj7bevkgtsYwvBYwQgaNOA6cz3z4jP+MmxJlpGwQnfL
SLQj6Fpwy/vF/3xjIHRvEPgoZT2HTSFB2o8Sk9hh87xVoxLusFJGwxIRs57QcTaX
KDk6PWsEfA/2WL+5DWvzNVYO8Du2ASfzegZcNFFk9tm4OnLYaPe1Q5Ns/ITa/U81
uWW2ldNxygwz/bNdFvj4L+4SSxBrlKUQNKEAkMxwZXyrs5/6ca1Jxz8+OMLfy+6H
Qx2EsiuOWA4YemYivTn/FqZgo5uBEz6rqEMoIADIyo+IN3Yc5n5KJgNzr3H7STbm
IHaJLuhm1qwojlAwNKk9GvnprpnldXT3Tcj6K94wEWTocp6DIfJSyIjOXsAyOyhP
UuFm12g5jJm56WY/qpVbEfAGRXaozKJuT5+eVcFK/P33U4q1brFLB7MkMa5iuqLM
OU4EQgW8ElKNjsO7lUmsmWnS56yYts483nPUQEU2SsVvPRVlkUyHHtyIQhcoRuDE
IlDhQT5efwdacI2vdHI0n0L4YZG4vZMVZI2RhtZ4wuNRyai8vCr2trLNHnKo+tDk
zI0jxdJVvaAVq2Bq0eM619L6/nLsURZBGTbV8ZNA5AXieZKbO/BEyJP4G7/r6cS+
i1CA+ltMrX4NUjZWZ8WK9oahWrQ1bhh81H5iOGUUVZyKq7xSU0DmCiavPwXOuv6V
e3amjPX2hbTgyaS/65WoqWdzEF7zR+jpgs/ZXrHZ8ucOSXl5Zoo5aQGZy/MHGjcP
1dBaM8ju4R2kgXiBBNcUZq0K/s9y4AjLv7/UwP6cuGqWW3ZrmNaKX28wwbnEGWRN
HUa9Jb5lLqVlJvYSnoD4X0V7iP8K99L8WFWjs3dF9SjSdagtCJ9zW/JnBxE72zzb
XjJPZkuGj2ezMxJJESHCCbkGn/yjz4T4vFAoj1oCWOIzZetBV96fuiDYRzUrxdzB
JzEu2UMdHbK8AOETH6l63DG8hu9DSMV34HokMT+DLEYCaJ8TtNT12LdTu4Sb/J7d
OUAxqEL6uroe2gpQgUzqIcD+QcUFy5O0+6O6CaOJhk+0aETMEZpW5zwKRGsF2HoD
OxHPa37sIWJ67OsbHPNeZwVlh725EKjf01TJb0DSQ9xN38RsyFjz4EA8J8XcFSoi
zEjkMEle0lkokJfCaEtfCtpDSivbLr+XwLWF5t2AH/5PUyAlkk1DPwpPhVBz2qkV
rrQ23CUj4eplpZ487crIiDGeqeDtUmohaQlLPjkcl+xKZMxklouGBvZD755qPLTl
Go1m2pvHMbv1ZlzTv79/mi8PKFIkaZH9R9+SAnKZHxGGPU43gexAAqGc+bPuGYND
YeM5fI0G2E/cKYuTwyWREWKtPpDbIVRPxnsyCgag47F9VDxc0aioi5lwI9xq1ErU
j1npUfFdirtv+rtfHNFxd+wE/1PXGzC/4MAD/Rc/pPmpqtu0O/u22KabGMvHn6hG
/lUQfpVBWtseRzDNLaQbxo6YuCCF0SHLws0yK+5PpVs/i0J3pzxP16C+BNQC72Ka
KBssoMc+Zp+BBQTAz1wG1EnqVr7HsPfbUvCVK0abptWRy1BSjwwKkFUsiVDr3Q33
2I6hvhNGhS8y1nKF4mAWAUwuDYMa5zC7t7UrcGeWntcpr/nho7fqHqgoFtSOn7Rf
w1CKYpy+FG+skfUR6FOzEX0f5oXMNRXOKUiHmv2mLiObORSfEAjCMocn/BRH7jqk
XwtxyD36MC0xDFbXN5SztHrfOdxrjSGK0d+P5aZkC/YhyCe7D1g/aW1BWc/Updxo
B+MveMnyX4Sp9GX0dVnIx9AA/iiUsbQKpbi3iE7ccqqSfPRQvmwe5K6BDAg4Nm1Q
KBb7vfNxaSG4cVOBp6b2I734WbgZGzSKyzumvY7CeP8pqqcKMdjPvT0gIBKYGfGV
wHCiaKRsUq2tmxMLLN3gPlz8zyihg85x+IxEXpIHtZYn4t/nIU+PhkWQh8Cx1KUk
sjxSFy56z38G+oD58adHV+bfSTw2chtv38BpFEF4YHJFZU45tB3am/+w1OMbCkqf
YBoLLsTysi8Bq3Eda/Z0d4f9N7ajOqTwe7zmApMu4Z41iiuCq3BJhZk3bbm+fW/Q
LniG+ZlmQd2mQuSRb3F8OFQW3aKLqBkUEG1MUhmTEb/gJggApX1m2e0LfM1gp9QN
u6vinByh+c79+BLOmR0Vea24DEZMkyz9NO7ey5ZQOurr4EpZPHXVm3J+9LUPej99
rAF7kKU02X2QGyCddhpRfHuFftPvj7LCOliAsdK1w8Xlv8xvpp9Rx/qke2GDiWrA
oazq+ASnqpB6KF9aWFhmgaIeUDrTdCq/Q6A+6d0+hgjaSy2ezrhHuR1MtFRc3fO8
vfs7QX+VN5kMrQL7TGAqn8B7Omal07wyqfG8wU/SfXz1TUsYbuc9XUtxNzmcle+j
5qpTY3xGjCIRY475RoIzGoa/3C4+L4cpiidmnnkc7TY4HZ8xPv+MgKaTD/6y6n5r
eBs7vWuhd5EvxkFfu4OgZIhfwRUGIOhU9pKRzFvcwy+LPHg0mxBKJIJ4KKBE/Tg8
pBoaYko//Hewf2AzBVgVYeYPsAVYqrKf5+Og9HjEpdOIF5sKwmsAaMS59siK5tpa
J02UyjFaG112db6uPU+JTyooHicD/nMzEPRZotEXPt4dytj3S5p1MuCld27KWTWC
kHD8WQFh4eS8UyiBKqp1GJ29miKB1bvXHy1PN1hh7aJE/e3LcqDIWh3oFisrGWbW
vng/6Jgzh7JyaINmh3gP3yVdNTO8sU3NIt+bDAvLQ9nF4l8fkPyPP0XrDpATfSlV
Fxz6fyOlnj35wQ3bXWl405hThKbLWksXvLDilgoA64+i/hx7tjJxevHfkcIMA/VU
zwoS92w+qNGDZbsGOJTbCm0K7Yua6ULnIN9BtOOfSM6ulPAv6Y9BlS4pI6jpVdQv
Ne+tcpy601yjjLxwSv3dhY/0llWnOCPCF26s4FqX33BgN0n08fzZ5hnyqMIIXF2g
nSrLcRO0yIMkIl6ctTfWKLi+nQ3txFX19ZLesrQcBox28uGew7Hs4Rpux9MNyId8
IEPQnykaAClOZEIZb2Btj6hMU0Dt90cl47I3ojhdWNagTHUI2X8AeO7zS8nbMLzD
l9kYdEnDpUxicPj68TRe/en6qiSp5GbstXXemzVj2tbIXMLdFFSOX8hDJqKOH/7Z
78mHWR4YylVQUeLzEMvOMiZCjQG8P7eRp0En5hc17nMKHCb2VtGs4azeF8ZaKmcr
ChYpUD2HNEGLNXus26030iirY+gmq61J8S8UGD/dWRiqIY6eeNkEEZbApV+PfuYA
A5+60hlTcBNK3wjpkUV27NRIcx2/K8p3yi9kQN2/JHxMq7H83HuYI0L8Om8FJAye
JhQhGqs8v6c9eB3E1Z6elJRCKXvz6RHeEWm0hrWinHAPq+jC4TYT5XRm5atb8HBv
N7q6bodE0KmKI9sPSXlitMhBMMSUrB8xehIg7COx2GhgjqabavkqYj7HG9U9NQzu
Ap6dxAoXSusiPXLN/SAfqnhjWYUrbQDA4yu23A8oAbBhqrF/B2Rf2i5q59yx1nKf
KVf7vZ1ANslA8OmPVyvcw6mCjxF0t0LKRiXER8ARLwj2gpKTQ39u9xyahy/1Op31
+jycBifoOoM2nDZOD30OoCu4oNFPbq63IZsCrC0cKofIvOnYcfLxjqGh2jdG0Fus
LnuOUmYw6itbKH+Gg6uGBlZ7M0Wqe3wevNBLzmheKnC1mR5CS8RDLgcwX/trzWzm
ew8Kikv0ri/ZhGhjcLLrSpmDfbDgTKwtvsV2SwENASGVjEOsJ2hwNhZOUPF9lK+0
2tdG3gf3YbcRIndcNxxr7anBIPW4ZGO22kXnOOXcpGLhcQJrZDd2wgA9qfK+aKTv
2RRBCyLQwQP9McbSrtBhhdVv2ocxOJag0dsEON6BSpKp6LTL5i5RvFZhoi6M36ru
OhUSw7vFuy/wufNeTdusPTRJw4bmlO3RBkukSQAJZ0UrswNuzc8p9zl+d1ZuyPMj
IezWaYcqACi+0YYyDbWG35SgbO6xKVyy9YkCQx77og7AdyjecZ4XazS5NlcPAxMp
C1jnFf58S7dkT0LnS7IB6GhH/c/R9iZOaVrNBOVaP5jBiOOyTxwzx4sn6ld7sNSO
Z/4G+42fhiPp/416IvT8ow18I5zgZafBBBSn/CS0iMVqL7sQXMHU9lEhSZuXoDad
aNhS7srhxDI7/q0qPsbuxXBTm02I7bVjN3FPIvPf9OcALK+P8C81h/rJyv31VzFE
aOQMUp/iyZ651hOgPa4NGbf1mCwForBryTzEuNiCM7pR48nv3YPAxHdPAH1e3evE
nbR+pD82zleexZ/Ok2Zka2QFSSrIy9yTvj8hrbCF2nocWF5rsytW20lH59wpWJCK
RH50AfE6raEptmt9og0wlBvcWwLINHw8WSOm4flXdc6r3X+pSbqk/YDWz4502ZVR
+YHJ8Qx6PQ6Kv/ur2Qz4MpPgWail1eA1zpP1tw324oBvfbM7fLJcYsZ9s90C433m
NHQG+uvq5F4pcYqZ83m/qkuuvTuzybJmKt2ILbZsGE7D2esnmYzTNtg4SB7V7NNv
tddbtbR6a5pdJ7xoLgdpXRTjoSj9FE2Oap5jtaLrHDxY8RE9aQJ6B4jtbLHXT25a
oAJhm5DQTlLhMrXksBDGkC2dIAa3t9c43KXn4VmDmwDcdhCxS9jEuh9hecMBvGP4
vDlRD0GUxkTE9nwBgencirVOzlRvSwjrmrW8z6f0vzRWs0z8gOTSu7Ul82La7uD9
t3LFHuJOKg5MkgvFF6oYMFIMm5C0G99Ynl2Bgaw/Mj2/b24oLxuEN/obgONUrC75
FK8h8A7nLaSjAs9ah+DL++KGJX33a26gB9Eysxk1PuA3kkK63JvWzN9Ybuv7LATC
Ya4k67LtE9w2R9OG5nsRmnY1Q1I08m5gdsA944GVC3IuHTnO4MrGKmBtyiC78gko
J+1NNSdq/AmNplimtf0FCGMb/R3+Ec7rBdLF9WhU0ULQLlEGeykKiQHkKNNfTAHD
/oTjNI9uWNxnpPrcCgIlVhixCBsLTRXFyIEFMDjH3jMKzIL9Z0biLnXPbgr/yRuc
5U8ATMN2MQ2N3TKNmLaoCPIFRMcQGeqi8v4n3XcrgB7OmHpxo5trzMJAOnkrEgeC
4My0DZSsKJ9c8gioutFUj9BnWBni9hrGsqTV4JesGjFXIgTA8fgjb31EEGxMHcRN
0Lb7SpA+qEOZ2Xfav4/lc79S0jd/EOFC4N8iIsmKnVG531O2JaDUIQ4HYvFTfu17
Ckg/Ma63ez2tXXwfrjPqVhGpZRtF+u8P8WvvQ20uPU1OjjmJ0Xroiomt7Ehi8vTp
Lodq8twElDNP7niFkkECUY5iaWFURNajdoUN3PC3Y3J7gtbHmB4pg311P0rbIX0S
WCzbb98HoEc0sARxQhrkuddPq1Ex6Z2/HP0yWdFtEeL43govWlG7+FaFdPFS4YYT
+XmsSVmOFcOEe1iTDta+3TzzZR+8GKY0yr365yrGwfI2O08M228Nle/qIR1AMH4g
D4gQVyc8bLkbxaJjXnsqt9YWBd4iPivQamW+WQ292ifLLDUJekV0AsydQ3rz+qTi
0vpLmBI5dBoUAmJ50rVFYESWECScUYzj9iJFfnaUcs9/FKg7izbUfyG8p4ZUzynM
rZk9TdCQ/Gz9CV1ymyuSI0Ikl1KVOKZ7IyQtoS2UY2jHnjyeoEG397lqn+WzY8Nq
6xmmJ5avmM+7YFGtDuZLoIOoqmwI00KX482GKephP+7HDqNfuXWawln0B4cjhZsN
Kl+qDStsvt04FNhZIWLelk+EOIhNUu3feIBeR40GsOgbp7ofi6tPeIHl9icfh3FV
IwYeMj6bP0hWQnNm0vladnSSTEdxi0fqHfGUQqFbybDo8hLRJombn6WNG70iJP5Y
LAorrJgkBDK+dj+YDvgpIkKBvgX259BKfG+7iLrjbt+YkyLqYdV5dCZ9LYsLpVvI
gnf++Bhcqk5wpf+pmY36g7+2vjqM18ccVdVjZIOZht5d+U/rgPy5aUkANS+Nxf3u
g46d90PGkx3GFUeV7WHJr9tQslOVBskxh2xuYrKYjCGg8bl2vXxlMH2squwycaZg
EG4sKNYdb876vVctXPrGTEi0um+1DB85NtRJit77UNEbUe6GMN4VguNfzg8m+XXA
zDNwrP0BJ9+xdsNP+WYHWP182GBaYU+EK6u1ckWyUgFzj8y4sxGrsVkWU+KYSSo1
jsz6MydbKhKFDupMeefz52US0ntVt6FVxmgS9owWXSdUODSlFvJO6fJ1Znqemwui
z4x/4qp5Gf9r5Oi6XDvTTPxaZtiB1wKw863SoZoP4MFTD5TqqTyivZWN1X2BRYFO
ik+Z85D17vsoQO44Zl7qyqoIqOB2UeKz4lrtTyh2SWua+0oI6IxXgClf3fBLJTBY
2RkPTnnMBVn6exY1QY0ac57CJeMN96k36OUvqzCia39SqLEuaMjSYhAtw/YWpwE9
ASG+uY3pf2RqC2nMJzG4QWJnaOP7uioGfSR0jRYtyxp9GtBgeQ6uojpG3IbwHZWm
vhOwNWTd2NwEBYmHnseOcQiL6MuaHUHlxvuDOVfpyXoGpBH3Bh9vUe8j2rNZUdvw
nNRp+GLpT39n80CcDuOeUW2xzxtoQzScau/W9V/Y17ubwitOvfK+OhIxpp5vq+SW
+Ooy/Pxvd+yjYdmp1S7tgK2VvjWsOdimkPGCOThsx4MkO2gUer7UfhCTP1XxmWVe
IWepqM41VCkFj+frtxQqrqbgx93smrelWLs4Mvp+XQwVxD9HuKCisQocYefsL6Rx
tT8GhHDKdyr8S3Sw2EPLJhuIn6OUiCLxZbhfKS7deP0hDI6nRji0+jvrcc1rCuC/
ZAU/I3BdzhKi6D1Sc85dKkjjSkQOLG22SXqWfHkCNI341IyIuDNg0eANJbDnuI6n
M9vaHtTnnZiB0wrNcWIGkPxKdC0/EKP6AyejX1BFyfkLOwyNABU1zBsN0dtqOMuh
Sq593Lj5bhL7OQWyv3Md5U69mrOM5urwe3XE7NXVMu4MiLckwA4byNVAeVKZSn25
HIvjAshGrOPGqk9ITzXVzt+c1BAzRFoEmH8igXRHHpc96wp4JxEnRf+7xGQvr64C
pPloAzpVVm+HjU7u/nsP/HqbWH4x0nREnnHfDlanN9G7GoqiwNXV+mSh1RJFK6AO
F4Fnp+NM/NEoL74U1l6J/BSo4LKC/ioxMFb7h5Frp4sWIXKYfeXj0GbGjPGvSZRu
gckbXxpTuDJoEmjQVlCDAxZT6dfl0ce/tnt5+ytoJQAzvFg0qY178wgbjasT8h4b
3DmiAPM0iIL80jtLAaFJ3vDZ3AikfR2gi0bOz40R0KTck3sFCckrdMYOCjUYk/Mi
DcTGXAtStpKasmXrRSEOsXDle0+slXguV7XpRsKXCvzMaem7hoFBK3Lk+NMQEH0X
pjDJ9LkFS/iYFnTEATXlPELUTNKTMdoX/CDGR1s9exGt45+3ju62LHv7V+AUkM/Z
LZfd/3XX2MwLoE7Rpga6Zr/SgNE4j2bh05YIpZMOj6Y6SWJaGo7KIWwMGCIeMa4g
tlseXSlFZlMS62IvMbUQ+h2ReJ+6eC62qakvAMauPyef/7/bJhrTObKuZ+KxlsQQ
xNqH1pkqrp9M5OF9dXS7x4aAAPQn18KZ32DmZTj4xxRkVoz8+nCZ85vWBEU6SiHa
ai5Icm0zLqH+TQQ/dVW+MbyxDpvBARcDBqrdIClAY14G5LRkFs2BIj88VvjwGh4L
QjXhSFPSZlE4CjrqPGZfaDpLHZ2SURkO0gnOb0rLm90L6U/SwRvkmhoWPUmx8VFQ
0Tk6CR0TeQW4JhKfP8u+H8siMAJDEw9sIRx70ILfc/ef79wA8qgIP5NfAIPuk49g
RNN160Z78hDM+PIPKDVINfW/24EJVAHZYsqol3MkpAQtV8J5fCZzCSLU7sZ9u5w6
/nOGTXCARHiMjO6UL4MFltUzKEz4w9mw7dKAM39LJJOAh0F7JCqxdG37RHSORCkN
Hl9mdy017EKcwwQFRWCRvS5j/mD02aJO4LciKBAzLmcE7qH9JQ3zXjqpZTspPZmt
HmKdlpp1whhQYCM9VmugY91+zxJ1Do4l96HN3m7gS6SACYsvmCRr+g16dMfHsbbA
m4yEgQyBTU5jh/YnJh8EmwP8syAEdnFfLy+Yb1Bm5Ce9BTckljJDJEpyMGAFF0hs
UEhGF5IjGYwKL58KH793GiSD5qRZA+X2sdysROkoGGhweanOjeQVqemZeiPJlJPU
aJHVCEcYy7y/IQm4jVHUe7OEIhDdAaoFcrqnDf9er6LXBEQ4DZY39GQ5/jA6h27B
VAYB5+ZroOProqdsqA/8jbySfVoNG6uqhfiezbafGYGJ0SmWL3g5pMgWX7W49x2R
S6tvn5YU91DitazTmkfJnGSvtrLaOtrQUskQigZUF56AnMwRUP7mDjlF7nZEW3Cb
AE+S9suH5WqL6tZd6IQjfO9cLW8i3tYkjk9u4ABHA28FDvabNhDHFPXtaXf4B2sj
z0i/gR1hR/IMaNJi39Hm5aCa0ewpWNk5D5z21g5tlFiFNUT5/PhDkISBxQae+z44
r9UQgOo1Q4aCyCYoEEE74MX4lsudW7TOO6i05qrwRnvJyk4kCUkyrdG2fRPAcETh
uIjxc0CP+boxt7ubpRzYso8RO5epY8Pm4+AwtmMg1WCET6D911WxFpzyxNJZAoGL
47pMBodq1pNMkaZmNr2gpXANUagIfuBY5hgft6kwquD9HyP8rGhmfE33AwV7GKEZ
GbKCyZT4sSBMSzOUReNEWAyD/UPGLowKWT8JiejD/LEZDAvA6qKZT1IohwJNHGQx
guc7ffJDrOknyY3zdDirnWqGzUNFiedH1KqMVM5IYD2kxi7wBanNjJr2+GBzO2hv
7LSvZ7Rk7+tB5QfetNmw0Aq5zBAKceOLhVL6eMD8lTw6IQ7VUrbGI0AwfiLk0+1G
RG8ZayEz3x+XkqlizSfNE/xHOfAQYeNf09fkxDWC0ip1AJoFOBhXs8SaXqUC68/H
lM8rxMRTP3SWFqirz+j4ejBNL7YzOuHRhZpSsRqbzNLcpfWJbTNGQ0yfIf44fj3e
dxB2haidSxeLu2yllgH6qzT6m7RQbgwN17Ge5csI9liCaOkGjg8JPRZrxKeG22OH
Yt1bIQ7K6jlzTe4cAh1piYYmoEF2jh388bNhaLnvTdJSyp0dPuawj/wQkl+Grn3I
H2wRGBjzG+U1RjLrWVW6N1vtULjRPwTbMG9XxA6DNU29YmGGRwHijl4s8EuaJbyj
u1XBjdcCW2ZKXoEIKZqO2G1coN/CgCqQFAksSc7pRCBqvYW6vqbWIyMbYeYol291
8SLhyQ97nfnZ31uNRJkgtu7IyXO8Kl902n0MRs4b5kNKEJMi2Pb4V777JUi6jlW8
WOm5RtCEGdThZh6xMj4giMUV3Qs/gg3zWRxDeSZPdwi/MoHWAv3s3jFpno9DcY1o
73g+FzCtd+yhnI7cTcQmxnZC+nWvPMNO41Hvn3bBmYe92z9ZDssyEygs6cPrI4Ao
PNTwYFCt2uunYrHYJANHPDhAxpHqp92HCUsDGf5kGBmMJee63ykKAKa86hr9RL5G
nhWSQMrJJFu9+1PwRBc2M1aBhjNosQafRDYRszcLm0AqJZF8gtP0P3bD8S3lDGNt
T9ljtrrBR2xl2J04KhDVETPLAgFQMCiVrtc3rQcP4I7YH0ZYMPZq1ekvWy5G0pBF
q81761koVpVoNwfLEE/7uXgaj1Wn9ZHjnqXSBV/0/b9RxeI3moDQ29Ns2iVYMcZ7
/FZG1iM4W/Esc3pEzC9p/pHaMx63D+toKNRglXPicACpSWbc2WNgY1B7YQGMyk/p
0fHy4FEI2bcs8KaILBICehU8Yw/bS9URjjP6E6QidgDNpZCSl2yBVPdi1KXViA9B
Z8BTDKloEUqPXHjkO4mlqMW+hAvIoh8F2IbQlIRcwV8ANIlrHEDP3DLgVneN3VmJ
DhaH8qsQ7AbDh7r2lCJMgv52lJr1roM/Mjz9MVf+Nrnfq01GmCi7fFwRxyPpI9vA
5pwFLBv35a8BCx6Hvh3jumDeeQwA7ICS2Gr5OmzxYTOn4DpB67aghDotZzL0bU8W
8Gl4QDysFH3ySwfxh2UXkRObypOMWgm8sOR/tteP3LmESl4sA7VP1ET8ryMg9VUF
Git2NIdG4//PwX6KWgoaiykdWgke3+9TyhjHdwRH+pEVUOyjBYxFOTjd7PewcqAz
mcmpTEkn8cbAahodIBaOB5fKVCaOfuizKWvcEiN8oeMLWc51AjH0/K1I5ujGbG7h
hI6HLwTv3xWryLbxJP0Dbm02UBb/zrBvLaRBl8FDHOWz2Y7Dmhq+91dVFnbqPpZD
sQM4A18u6WE8sumER5Hpj8fA7KLBf1HPsNAe7bjief4aEHpmt3XdU6UpjbWVELmL
8eULhbyUXJKQ3zjZAqH2Y/5MLl2d7dq8Bgofp43qsSBqQv+iHHVQiOWQOjG/q/pP
hYHgo3NF4bsal+iG+NzjzZX4eeFV/NpEUwt2nCGlJdwShmzktA2HKzlfNkD7xhlw
d82vKFP7PANuOm2mZaUKAn70P/qijU0A2dfIMBqdH897l2ccHjqBQc9qgNOHY+Ia
MVg3SKsObNJuVAE+IWL6VsSu0fBvZsmY3iLcoKFiZuJTCd2CNs9Ez+k5E7a/ICil
WRehJ8MADYlAbyh3QhDakm/swIDzhqAOObSqgJuA4qbtc8aghRrwYOB+Bk+J/Lq5
CSQJAdw13z5uWPlw1lQdqGywmJRogoiwoz1rO2wbOXFOcye9ziE361hYiqoBs5s3
hqmS/YSatzDN2M+cRhAPWkvdqabO4jFEpwvNNXRwnDA+P5Q+1BZtBKXm/8zE2nXq
mR1gyuSR480euGztuJfxksaTAlQ2vBTL+2AGKt5uLCIUNnpTDVlbEf14czGYPDbM
ZC0nHfRSYn3k0laRba0Jp+GwdYqQNfzveqv+hWi13J1+O8Bo9ZM+WEpKNwF0gKuo
8jKZ7woAp3Ypp2Z16Vv9nxuVA0Ido84CZT8sgprn/BEDl6XJ+FMpqTI5NybbBNiu
hDSzHhHi736FtP1sscwNBmv/G7C4XHQbR28DjK/HBLDNGU4x/4//6nOfx/oyzl4F
8udH7q2DhkpBmstaz59W/bKhhk3bON44DK/UZsW/9yzRdPa4+foFlQyR6yYcm+fR
PHl57t40fG366d855IinYlXvTnndJEi7xVx5p2Cbu5Bit1bz8F7KDauNV2hTDshw
/Ol0HM+Rst1MHjftZQQpT/GS//NEzIuZB5tU0+RTyPbIEKYZr//iu0JMt1FuP8Vv
JwfD51tvV1BhsCkJV3PllPgqKd15JUFK9nx3qkBh2vQs7p2f0Kxlcawle5CtTsMF
KSKDAvEQ7OhQ1FDd6CQWFUWROV/t0lFV1LPz7cfH4wUSvpsNtkRtVJeqfqU0beMD
xS73bDSAcEIduvWp4tP+yPgFXDqN+RaQ4vLjYR0Ux4xX5KA+i0W2n48kpUxLA7yy
t5fgDiTobE8OONTou3XHCThdGvzrCqa+RhBsQjRNhT41+BbUWqF8IsjqOXI7BR+n
edsQfBKGmDVwaIn9Q6QcRhkKFv7SKwS1/9mtB+tDeLGPJKzfkcZ6NJC8L6F2+faM
n/tD71dUQTqcv9LX0idJpV61CZbXBA8rLHJXutmab34Vzi16Y4JfyP7JgvqhFMIt
efOr1/gOoMPUGx7vTn1hhNc2DV7GRRQYaygXWGwCPnc86hjZq2WozFwVmYwvp6+5
kNIroHSwA/Jvv996+Ig9X7VYJzj9GoJKpSXrwZDDVWdd1V5BykreYIQjvsTEP4xP
EU+GxzgFhPP2NF+oWoHnhf6DWJCOYybQRALdAVk90tbVi/ZbEdPCELERkJguzu37
DqBOzMgxveR81F+lMVMrVlEea3oWGAWIJA3iCw75qP7niqqPLK3Qi+/S5DAiit7U
GG9oHC0OZNZ2maFQEIoSwbwFsGtx+FwxW9FT6BSSmeuzHrxfF2pw6RNuG6NE+6jU
VQGd7A+v6QO8Ng4rdu3l9I4CaqlHrcIkRpAEOXn/TuRZKQCtvSWWCIjPaOOMS6OZ
u30X9dzsln9OztTDldkp3nH+K8YMMTUv0VgURPVekE6j5TZvyA5NtoR2mHuCT8dP
p2iSQr8OWEYk56Uy8pn2GHJvpjei1THhXMtES0lt06WPXikb1VweyK0Gt3eaiUH4
2u1VXjNuTmV3apzhLumlQxY15P2iUVtvieZwSOoZrYKn9soELJY1ceB7FfcSkEft
CVnQclEdsxJmjCgv0pXWjCJlAyZyNWoDvK0OQcdS5RZX6WctXjmG6owsNE/PQZIr
hZDkud5SEWh5W59GQkukZcj5yVN8/7+GgtgVIdYGrFhc4cUg2oxwe8qWe3h0/MQn
1yK3DBZYIE5LULjqgU2HN7ieEoG0OBZ+AwjqfbE27bN5lHMC0YLZkdbOjMJ9XXY8
x5izLhdvod6FA3NjUMiEyUPE7qgNlwa1Htt3ppFSz9xAIzlQWOn40MO42p2lzl2M
suphHAl23qUQqdrpEAFQIqaU0MCcFOB3E7AvYKrgMnfCf8G5gelwZ9JXpdsH531g
yKamIh6rFW8g0xivh7rz4AopdT3remHd58+kXGfl+XmPM4G1jziTqWGqcgSMExNB
fMUDAZBPNNqGxVseguXtMM4Hn8ne48qemI7dfgGJJkTg0Wwyw5xPuOyuWofO3TgK
jQxXTOqwvMfIlSVt6usPMrdLIP7af3nwMsa4mrQ8d5eQC6kwkOcX/am7mfCWucMs
hjuXWF4H/EWuMJaT4V0/JpImxXWFVGyxi2zWQK4wSA7sBkfUu0n0JJE1YGFshI9Y
CSJiLTr+JT9WQyNLuVodskaPBJBap/RNcKgY0kWy77Io40NG4iY778SxRnxAmYXk
B+F7dOWcVDhBZuowVc2HWHLNPZpvF05U17TbyMwObrZvQeCoRfcz74Munaz8VvvY
NgehWM70/qTLmpaB2xLw/zzZxA+ahCq3MPKHAanaXW0UsrvOd4XPn//c5o/ePmUQ
KKr6B+aO9CkVi0Cz4tGlkdEpL0O1HcLFu4wpfhNCIu67aW8iV7967WUYWKjwXuVz
RQOAPXKP1TwOspcW2aLoIYMQjAh4LMYpvDci53ADVDm9rGNNSyg1fMq1Dh7jBY/f
6y97/JS/a5JaT3QbeaB6zjGsfEHKBA9p3KQlJLwpuhGpJSo71qXVKp9sHBYgIba1
PqPi/fbdbfCnfH/gZLeFfDnIHfA0MhHyj6aK3nWrMjCKFMd8ANU8JFo421UQoJ1L
rccmrFWtyeeAAocUH9bx/0+guRcjmjO5A2Sggfua/qyMyGVOWujbNqwb3uU7+JD5
xYBrLudX+n66oziiGT4gyNyIhgmIN9h5IpYIBFWBmjcKtrKTC4/AO8g/t3kQ6bSM
feb8evhQyOXFFSOZPacUkLe5zVVjWg+iaGEl2Q4AVSlTJH+D9clICSvotujls8TM
Nhw2CaNLmxi9nb5FUvoSMNm95t66WfqvFWfPTzqtGbiPl+fOp8Tc2UrdXPZxAM74
buC/iu/kKi7vLO4f59P5nyoxRqML4ANF4SjPMETTiE9AkKxDCLgUDnYHGWs2uQq5
tyd0eq4RFiROOKy9XzXa/05dmS+dtSHYKtberlqaI1LjBcZQryq56YBnXBa1Qoxu
t1XZJZulVUjI0cn/Thg/sX10K8LP//iW4H0OXUBm//eHJGg42TC5Em9qsBUY2l3b
9wKDwBe9cRVxnVDJKykQQrBrClFpJR5vSylomzLqZOBc2EXfYgdx/ygl9FQtz+c2
GQKWkOmzPjUu4wk9/0tCIREEoVKAYWEs2tK5jGWMs1EhTF8FoAMW6nPfIGlC3hxH
lWbcQw4kR+SgWe5NFxL8HRaPbjRYX6MvSucXg9J4WxMkwh13U9tx5Dz/FNomD1ve
lv47TcI+KC3RtvpT9dPfZDH4y8PRQdQVEVTfyIOKQX1lFIE8MaIDW4NWb62hex1K
TY7z747i75asUau9GQx5eXaAEyjxCowj1IYJj1duF957HITxT9pjlDVobFYn/I37
iIeofANnUln4qYKir00/+HC5mUBsdCKZu12bxGiVj+C0hqrTHPAQxQ0/vw/MgPYt
aYAz5ilT6pw7M0OQlWzIEeIps6Y75fF98EVH584/16kIVvPDXY3BZLGX6ziTjN/f
lBe01bcWHNG/8SzV9UjoYLTbtXwNOCCtbHqL7HFwC3PNesjEndwoXCXYq2Zxds2e
fKHPSROOFi17xy9UiaIcqU21NecF1nq+Iu++4vHKXwgHULVc0ZlUIM0ABN0TjdOP
sRsxMvGAV4hFb9uq61bwHeVS1pFGdItx5BL9l6FhTzXGn0o3nnas0orvH36TSdid
zoFGG9iexhN1kEZYCPStFVgsIT9eAm+KQUhbn1AiofvUgm7vYgjJjWClTJsIo7Yi
YqTs4OjqMQu9YajYj+GFwYxMO366tPLJjXeXGAJU/hdDywJ1Vfk6XD+vuCXOC0tr
llHoBpz5YX4ScZ7jexUFVDS6A7jjZ88A0lz470hHC9GzGHC21oL3MEEefg6O8mtv
BeW0qsyI74dfgEflrs5w1q4Wti4RjUyxju7KMDu26k1KzPlOuN5wbkNdIkp3gXx3
aucUJ9KNQD6r5+wh9lLIJa/mqDuDlm0vH+ul9I+KS4Gxbp+TT9Qt7GkJ+Oy55wKs
haCkkpNHzPPgBzDwdQPXH/6KqWXr1Cw4UMkYSI6dvXuhhspFWXgDODXR0BV/0eVl
oXvt9l5qG6impwrA49upjM5/bWI8Ixb+jwdDVlay2OD6/DrlG1mrgYkMj7C7UVwg
uiGhXHVSVYARlyncDBpUWB5dEc1fq3p/geK5FYl8vXv5yI0FIx29JdLq+D1doUNZ
rrhzxJMbRiM7daQJsqS9IMgKLVKtgwonqiZzZaQV/0QPDSHgwybtGxhpuZCSgzrj
HfwTOTTguIAUa3kZwgbm0MED4DRw+/5PHvy3ecuLKPHUvoZve51UPwHVGB5k1s0b
CdTCvTsO/g4Rs4lTcxepO9xRIQ+WM5056Qy9v3P3AUeeVZZZf9Bt6cfLiDSNIsCV
+Zdl0gUIxNMBttp/YKMU7u2HCk/c2d3B2ooYDsL49KkJvkJv/4B3HaiY1NSwSh44
fi0r2COQfE8zlCs3GipcunvtFfNDUdUIC7GOXZRBORLGleVy6NQf6JmakVm/sOyO
aSqFJcyhHpB/4/ZpJU4/OErY7Icfh91Mck/oYMryvn4IGjwi/LRstuCEbPnxLMqq
jiKU+f8qWCeHxGblx9CYnyNmL+RnUZTdPER3XgdpLeOq2RctbuTWBrDyS6W2MaXf
Ax8K1o+U1++udyE9FBuhhxiAMUxZrYE7S3wH6zWNaOpkwHmCKgSCFuxHNoMgupNE
W35tDRKzQ4extPscxyev3rnExj75crt5Yq5B4YFI090VgTw/SU04DK3/jtXzuIHn
IVhbvqY4dxq5jlkUM2vrsfDzDaYTxpuz476G8HAwv04ogfEQ+bVf+dFzB4eYGQBX
uAOvPByvLW+3rw4egnBZj6SK6cEOVMIpcS8jre93k0wWxK9g8UXMruV4uLG5GUbB
9OLUdT8yCeIl5WY/moWZkEc3FwK/6/iypPKjBdZy9N9rWYC/9qrbWA04cUNJhInh
nJV3Sf4U0S4InIdgm43w32laDtzgwfGTO1DcGz64cVAypJf+L/LWUNerbEJtnPqj
hM2+w9z4bT2zG8aBzXdfAKK5fDfXqGGXYZEEillq+im2nq78WedMPzkbO/wScu26
8jO8g1ubFOCPzJ6LLiT/4+wiAW53pfCsVNxVmFnIVKPv9qtqpGp7p4XlkdJBILGi
zZcxfpbJu73ivcqyaZbtAsLRHIn+ZQxWf+9anPH2ZF1628CfYJeNhyCyNjfg7WYr
94p/YzaAJZBXtIk8fEIdV64FanhLC7lTPQwp8PaYtUo6pbiS+AV62nReFXkb18xW
dWxvWZgmFeupXGtq0ZA0fPyx/LB8U1KvDj2XbHEnSBdDsxv/ZwwoHRp2B1YKJlW8
vP2ltP3VQo9VslFQd54ZLFVjKRxcesQvPdDVs8YuJPyAn6TioySYSeCLfxfvc7BM
GrR+DHGmtnCoEou9Edbyi44LGWySwl3HiKCkKFnmedOMizpSlHhJp9TnwUv9jAXk
ukqiv4Q6fKyHRjO885vxSTR+V1fAPz+sojhII8ED9tWyYMYX5UPMFHbgFhtNQZT9
FRonCy8HaGSWaHsTa8ABZEOfkLufCNlxMbeAtM0OxqvP0aZktGS3qqdWruGEJfGy
/wA00F9gJQhPWSFNDFdeZglEhjktDo8q1oeMeiMlfug7VeoWpR5Hgc6n1zroym6p
ibcUyE+kdAWEQkOeEj1Nph4NXHR1lRyaQssUm6/i5TgomMifa1DkuZtiMEA4FPzz
gGwaquthDvuzyQCrLdRG3wskLIfEPT1JlcpEW8aXUR1YKFssGEGhpKsZzxhmWACq
lP5nzW4vNLVaqkjLzSfms19LL0Jz4MCyKShzR94/XNpkM4DzE5aU0zKLCtYJ62lR
n7Fewim/PEfX2vlPu+FQPl2HO7uWrrJZsOeuOCJnH4fAAyA+d3am+5Aru1wc8UWl
kt4OJXtE+jq0KZbrMiWhNiIL00tEmi+XQn0mckqUZBHb3XCRRHPuX35LPAB5wWTK
dVg3xcrlLnPIK7UVQj2Li+05hX3HiVS6pNrVkD5C95T4Y5Zb4YrzBDuToIwvx0/z
r5696xnQbl8B5x+8zb1Og5wPQkp7yVk3MuhUIEz0mxTVonwu9zMlpGHEo3WtCCLw
FXhGzk8L7yJ/kNr+q1M8rVF6SP4P9z9oa/pY7QTKG1ABVpqzr1CB8l2YIn0Zlg6H
EuQuBHpIVRkXwWR8IPOMjIL262h4gBrgd5DqmEMa/kVpN2syFzKL+eGKFFZP+r7K
Pp7NvmJxqjUbgF97i3/WUQtS2lqDnKgRN8Yr3cpul4pTrjWdbz08f2Dj2jpqEkqX
di0iwdnAJTaNNADlgvTRFyAIOPOyUYb7VNNjL4WnScswFn98gyIAhhdLDhG3oUh1
hNCpA6mrDvwDYJkQQbXlcWjNCyN4TGEMGxNrLRXRKVAYytQOC/ZxyJ+K0uwOW7uY
ZRkUkxYn785oEHqMGfb50rG+R6DWUh4Uw+x98Vvff5S0UIbq2fZn+EwkzFtg2eoS
s7/aj7eWqJBP/Iwz9bNNIxRY6JjaHmVU4He14DUP9nirfqXmxXeg/trBGdpbG1Aw
NxPe+pp+9J6VeRfxKDYMiwevmwxQ23plxCUNqR0MXFHhDuLRJDhYK7lMjsctQfVH
9s4F8PmYLR0Sf/N3DX+P9xm9/YIE3SriUBstyXWQ/sBCBsYnkXry3J9dki0jhqNu
937aZk/qnpou6UQFyaBJXyi/tpuC+E6lrbpS8u0lP77VHDiwd4S8SGGsp1wVr4yw
TVHADEyzZUumaYnkIuKOn27YKFe2yhkLHit9asO/0/C3mR28T6cuS8gGgKmvI3f2
ODBVB56DpT4NAoFbx4rEEsVU0LAq10zcqmGyyOA1OjM/OKlF9Q3yXmFRY5T9DlRp
VfWGBZVOGEqmkFz9r1YffGvcuJLj7KFCvOPQsLoNtRInjHMkf+QiTuxDRxPM1oCT
Bzcl9c8lJ13Yua8hoCQYXoyv+mbq3GPYElFBJ+lFC6frxD0ZAKyE7xgEgn4iFtfO
QTEe3Z6OKvZDYtthZwnBvmlcST5KZh6gDloncm6qjZH8mN9jinEN7lu48gFeQI1s
Q2yLyNPVqJ2tv00FjibeEksEEYJjQ5AQETrjqADeY9e09BjTIguoGpkfSQooY4JN
Ro4KIiY6RPlKja+x13RqhAISkZGeaLOX+gzi5mqUWUup1Qf5zT7sqySaQT28LWnm
5RdkswtVtogcBKRmbn6sQXwbCsVJ2rieiV0pmN0vS/XyuF4r0rW6SaV2A9RzS+8+
nyc7TVH26OdVZ/eSqU3tkRRPF4iLThPf+/V2F/WSLE5WFvoS+xgCrClWPm2OffGm
n094Afw+vxMmA+uMb+18OcWylveJsgIsXOGNfogMv9pBdEM93Ok79ms4Z8jHp/YM
oyf6vpUk/y/ewFe9DQoi87dPt/lmk/Oabys8wNk21kkglT5XW7OVNZDYqVdSYIiW
fs7aJBWnaljieLaaU4lHy//+EjM2ZauehEK4OyBP3kJM5Ju51xxldvBNfoEzcYXq
wvnvLBkkkYCxPKXEGucyVNRtD2W+eQA7cH+1eERVEI953DhFXCwTOLfOqcMwmUGV
M52FFwVstiEl/8dCjQRqx2dd8i/1z3ORVr8BCTHPacoW7a/KEx6kPfivcOMEH/nw
wqzeggylgZ/yOnETs/aSE0BqDwECfkJ/04WEuoQf18EifpKadACIcFzesj9s41w9
qGTFsDWyXTu4ysSqL5UiCtPJfV6Pu3JkWsjP3bXoPuWBeaaitahIR5vmLeh9sIUr
RmN9Xj//CW7bQxPkMEE87+IHGpCjLJHHfsU2VK3yVNX+Q0p6fEMUYP4fIMIpC5BQ
9h1iAMn9JW3Y2QTza20WvNT7Ps8I0dHDME5SNESRGUMboiOZDXonDuh7bepzU+BC
EV5jX4+bc0++PJ7f+vIKzFKvI2LiKDsBvT0Rph1KEPJ80X3xZ81l9jC3gyIj7ZRr
lnGpX+oae8wAptp1z94HQPPFaRQrGGnKXYD9qyhfV+4UegA1Y7t8IExe+n0TRi+1
r4ZfGS1J4nvaQFHMVv6yrAuht33f+VPHIGJp02QsmA42pAdtFYDM1peoSIQXaQx3
Cdtxsa9kt0gknX2HC15bpTtb/9+VJt+RwVUwIuwdC+AxjcJlD8hlDuE3Ejlc8JWA
mEQyUJyk5wlaC3MZlEDODyZ+Iq9+M+k4KfFcBsq8Lj0ZgdmFb+XtRYPEL+LrzpaM
czjxScvgUj+JI13tD92XlkX+UGsD5FlQeW5a4OTtMHypzWejZXjuMyfTMD46q1rl
eP8Kk1YC+2M+aFS6tRYpEYrrygE5HCMdkg7jFzvvpaFpwxcb5H5d4+fc3mQ56rGd
Xm5GLhQB2TCBDzLAQEi2R7MT5hoccUWJcS8qxnPtlbOqNLZoGB5T+/jcd8d60PE8
at1uV9/3/c8s5hnZc+ZOK/aUzZ107L19gRd/BjSAfqvmrCwp3S0E3tUKlDqmgHI9
AE8B0EEb4Tk8raBS/qQKIYf8SWQrbB0YmXYS5jJJ+t56d/o2irCaDq3sVu/wQX8W
aAsUVohaTWz/PBTqcACKVe7nHfT9gaEWM7HhRMe3nX+hMQ8/Qkw4dDr+L47XGzSh
hkgxOB/n4vp56sOKXkGZgfMx9t/cvC6TjEbt7mKxtY0B8INooEaTk6K3qgajDBkQ
qMSNwsSOY2+XGZzo5r+2EmdC6WMZ4UGGW3s03PcG43NGzMVeMBC+/pavTXHRRUrN
ZcjSnyfbEhDKuXfAgvxyblXVRY+BI+NRjOwm0mXjJpKWoViHV0Z7V3Kj6AlVdntw
+7o6JXhiN76vZISvI2VtwedvkTVOsUlihKluuKZk+Y/SuLXT/YqahrGbqN4PSIpQ
eJvyNDhiWG2lLyJUILBbUGqYVcjPRGnQ9qBhb6Czyn2acmc1coiVBNMwjW2GNNO7
6Jwk2DTYPffvlLTtsP+XrEdpGJ3PGb7ZpfbuvaSnGEf4JaH7QziSMv2z6qjp4Cqy
IW38x7bVOdArh8awlfbzPDgSYQus1vLs0Fmx5baXQhR6X/qw/1i5DBGU44dTWG17
GSAVYDGPehOzTukJlY7Zia4XMelRizPHs8vNPAUJ3z8tGV/SbkydAL7pmaMxbRnD
0zu06fQ1KmeGDE+oxRoyWp3Nw3I0E4F/oo/7YxDiuKE/2KWsR5eMJCF8h79SVgto
XhavvLPqwM4wG1/tyh2B1+EkUwQOv/gaeA/mVzIHgCDC7fDRkJKQFVNjtovaAlIf
8RXpunNSrHhV9DpLXoxzsX+OaLU4ACuo1HMvcP1bJUvnh7fkhRjJwds5eTjePVQX
OSqE+CO0UwE8pKeZsklF0WPS11i99L/a52ZWojTYDC42LITYquxpG5JFy1WcBNhl
RIGUjc3PeRv2L61MdCcYe0OCvbtwrAjUPeT6C1KCaXRoPUoK8mqUud6vCIo3ZEZn
tzhZI8lxGcucazORQy4YKsG8YctSdrCK1aTDMRv6up4qO21QtrE/M8Q7r5DGlD0i
wrrHjKzQVmE6oMDlYgtugSFf/6IqzWJGCfv6edJGjxB+PvugX7laZvS1cAZSakpJ
IBQBCtG44vYWmTyXjXMxdwj08pPwiuLayvAi+29DVPPI+uBKdhKxKvRbIPm9KpT6
7dvYCeB2r9npGJxLG6xWsO/vh923KoXKQp2wjyOBY//ibq4x5XsffRZVQY4a1enr
3F/LBfsrkYhCahuo9aI4hEWjTTqqSRXRaPvqozWODIJyfXRa2YDLRSUM0NzyAYif
NgcR/CwPeozQ+1AAf7FFL3FFX9LMIeuhLpwLvufoS8iPhgeWD9waH9hrkwnq0ecW
VbpNNaSpFFvdoGA+38z9FD4Ziagj2Q9+LGunBJzjA+puqnXa8Gb+slvuNiMJ7QWj
zyLIYUfB+Fg329MNnid4kQi2FQN9LfkmfrLc0/wNGuaNybF0G0x08Rv3Qhhhupvk
Tz5a8EmVyS1ZzhYsUkvigviD8xtNWyX6K/YtgjLD9NFqDX3VE9VEKML8fIzrOxdG
n78GU6jiBLOdu6VTdMOC5y3eFc/XnAitt5IbhptwZEfwZwW4VuL4i0dY1Cky0bWs
QJu74uH4JrLMFiNWV4iMtTMIbWrKGxDtF22L+oZmrmhReyuI33dtpD6BjXVqP2hy
ofwJFFikoNFVupB//QAPzE2LXf5k/rAo+wSRiZbdTdmKWwV315rRJqQZoUBEy4+r
hF/INmo5GPHo1rXcmVmUM2/MRYT+nSNgOiCBXy/QXcIFGkFk+bNbnpLyzPEK31fs
VIhl8ERHg1TzmfUNUA5D2kpJ3pfZXMtpMg/v0Z254BOddZ4UjY39NI+s7xxg95nq
u0x1JSvmlkzm/oi7jzYOUCIqCRouHj928RBYKWMX5elgmsWJm3wOCCtpFo1uhRYf
apKLVq8OVO/KPCyLoO9gP8Cg+VqlE+UtqPjqbWwCy+2tShCkKDoKc+6ZXGUOR1N7
6kK6MoBnolZg8wYkZrKvqpnZbWP5815ZH260NUJ3Uvkxa/Jbn1Je174mh6y6Z9Hp
Lp/SFsPWq77ZfdsDnV9XvsNa/h7AJitcNohefpu+6daKDbn96zgIeIsrJz825dKP
Jc6GR60rC6xuXstbvsIKkid/KMrGj1i62omZ4QaX7craAxti7BgA/vaiL51nCOQR
pjgR7v7VXTxCPVWbvWTIly+GE2mb2e+ur1IqKI8iDPS96Y+YUNc59MNWZCWgNRx/
D1PjyHNSVgrhA3XUeAYa0uGNKKEkcAs1Xh1thEN3IaeA0LDxvGnAHAx6SkazXa2t
ahVSvwFCYWAv1BluU/7a3xnI8WTVllMsm0GzqCYheaTIVNrFHlgdnfw0ZXHXaHDY
g3VBhmImWPEytIBF0Bx8la2WaOkswsA/OYpEfCTzERcgLvLsFOAuqxd6uq/ofiiO
XiptvGkWcbH4tUzPRaAI2fDeZciv4HZ0hiiPLJKCcLYu3hpctwL8AdaUrMyysB4S
vDkw3Bz4GiGKeksejIyuCBQp5nHGsh8We6utaRKSQokX1n4VNRxQI5CWPTjj4bTf
UUJD7bYW8ZfSqXYwUvJYkMDavqjREe3IdfughupkjwJS+TiyTXNqSuy2gvDzHtB8
50bh5r+K6Jx2XokOouL82I8mbM2nXpGy76FEnZOQuF/sDOSVx2pjldf6CLiztpeP
jNr3tquRujnbiAMZWfoCBBMH4Pmjs/Qt94SdPgh3Xupxi2EG4GaaNUFwrjSwDpwG
w/ikpkhjor8TYS4GUQgscGPEliv+EJyOi6/X+kOM2hcS/kx7YXUAVLpAv8OSnQP0
wSYJeOfDJEPertHItYbQxLY1EXWNpud3B6OD6Prkrn/X2doGR5AD9pc8AHpLsf+J
+uyJZX+iiQQ2BRP+mtsw3TAA+TEMghYeyJyDHREmSkVWeVxFQlvxcEPLrAfCfRU5
xqCLmVVNg3FeynvVl/9uARo6l49JBJdHJoHVL7vSnzJSw0ZDlTJ/cQ1R4bKbdrXU
Wowlh0VXIk1f50peq9DHxIltCy/t2jSE8LnT/iBz7XltZxXLcfoerSn1nBhVekPX
QmfOtFxiXeGFpi2G9mNiXEEPPO8hhCJakCncukJZVriFgIJsRjbGAcDcwpBRfceL
4S2ziHNu+SjN4m3nn8g3vF/yXaTEE7d5vtJVgUBJb9wxWx2johW07aqnQCIob7W5
RdcwpqQEW045lzrKUvcCh3stE1t4Nh33g1idU+59g22uq7EgE78q05NOrZ7bLpso
w0mD2VBNSbfV3ai5U1uyyFLNkipG0dFAp0Yfzpner69mcEmo8x22KUR4Gr/am3/O
rH297F5y7lk5fulI26RuL5SvM3RwaAdnc2atG/0j+/0RsVbD4OKU+tsfm2yLAigh
cTLYGRbdZ4fcB7rj3w60wq9LdhYapTJLxdX9ZYbMRokfwOVMwpg5EEgc9hLpyldf
Nsexlx+xbw1FDePulbLVAk42FY9YQeHaOBompvqO2LfOQKgiecKDYnECVdVtwUO9
CVqAGl7LRJIxnjSsv0WHjFIBlSsjsxS8IT60wP5dV5QbffgSlyEFj4Duf08qa4Q9
D7pQwS36l6usCr0axoqacacH2GRhChBR/WB5KD8doMO1FVu0j8XvbjZlM3dOkFEp
+hTy9UDJ/rof3H4wyER+k/OokSqFmNwuesZUs0vhwQi6pdQFUIpVQrwX+WdWyMzE
k2W9c6TU3jZp5TodsU12Kq3feRCxs6RNPpu9A7BkRryOEWbHmmM+X0csoNowsIlH
/5io5k9sAQVxW21pJd6ch35IhFw+40WgbS0yOKm1XTrrqoI9ISN7V1TlpPZk44Vq
OqDtuTeT6JTPEC8RZtnarL/h7NEgd+i7zrh9SIgIEcP2i2Z5lOwbREPxBnLnTgZv
GC2gX9nyYUvk+Qj1LaKFrGFkfngH0Amiqw24zjDGIekXxeZIa3NKa4o8D9mZtl25
rRPFcuZ0tIrtm6xfNTWPeyvwv8nXWmYdlJTr/kmVicOK5dHnWRaOcuv/oGvS3/5y
Z8ONaPTHgby05q+OY9NDRB8XpUfNGggtLId7rCc0YDsAw6MDLzw+dFb5ZBpDOnsp
87Wq5onAXA0FdzAppN7cl2R1L2Z+ts3PS0j5tnuVZSYT2MWvt3y2GxlOBSZnDrzh
G7kafzt57PAe4rSklDW1/zSDavV6JfAm51w9QFLIMuCNNxmiAszBoC9eGbWArEeS
RPVGOrHgCEdI5t37pg7NHCl+miDznMlKA+LOfrXS+PvbEU+YpidU4gq21WliBJF4
1eF2ZA7yRo0Ra4FP4xZt+Z4y4nSusvbxajmO6EqU34QsJf79+UErvjOE6kdKeVE+
+DRRO+IrDzqmVlWc2JpROrFWXXBwAVsbbToeGTPrm18CTgOrlFjW8pIywxl6RWiW
Epvl5FlIrMGI5LRPWlej5tQMJDTuaOcu6uaTjMMA64uSlTCzNGV7RsM4/1PpaODV
9kLZ3429fBAa9zcHCOmUVnl4gnzKsuHsfcmqV83b9MjbriqnWfT0vT50UI5lPun7
R4dUftVoccW3gTdMAi2EvYwIhByzfd7QF4zTHL/KKOq3uRrJ7HLcSsr2OZ5QOma/
eInDVT+joPwzZRb/dmm5U+z/07QdiOV135gfgrDZNv0YXXryj9R/rnvgLjaBosP2
DxmFWyOx2yqhobgpRWvMlL+tRj1oIOckIJSGqlualRGp45wBsNcV/Tml0z5kAyU3
76nZIz6VqRrA1FdSa3ddHj9OBQiqKWlq0fKAweLAVktIsdNNgUxEmt6T2hsYwUST
e6h0Q+/k8q8NhDzHXQcgI/So+HF8E+0EjQg7kpGyb6Ype8wneEcLc55o9nfpU7ZI
+Tmy73MSGvo/9ifD0+CYCqlGg6hDwdJmAwZnZeeakYjyAEJ3KD4CT6NuRgDDGSo+
fXnAxW9ogpvgR8rgUU10NQNx9aOmqJucyCCR9NZvb4M7FFqHVzMmRgcSp0ftAGcy
L6EGqS5Y/tKEMNxL/O1MSBGJ+4FcN76ABvKtmlH5SFPwZSDTmpETUWUzHHVduUeI
3gfQt82aaQDUf4hY84hrTtuG+rAzo9bq0gxYDowffCo3ibTdJoojuTzk3oF9yz1I
uDX8GnO+o0ODeYPOlRV6aEWpWV6nCq30UHMUA+eycuN1maWJcFh3+tbykZW6KhFl
Sv9pAruHGgYzUlAykVDnWPnWBiXVH9lPEGVe46ie1AZIjUDMYGYA7d0xBQ/4Hp+i
Yg0oIVF0MLGmBvoxQ6fQQ6wAnONHka8M3f24nJu0crKXOInrHhBSoHcGUrvvLNmp
NKEtvHeT9wCxXrt8P/OVaz3gdiCWkbW94qdFs60RFJcuPhif3BRuduwweKhi88qZ
NiBfMuBf0wQW28N2RcdrppVPqn8s7lDhzsZ9bGAjhdjZDmZos6fkFjQbSFQ/HzVI
limd3hD72o9o1/QFxbTFMTi4ngKGeO2iG2HDcdwbvQBKpE+0E+UDGkrVx4XlBiEC
QNX9VLM6AZnulmZrLJqdOdGmb9K+EuKxnXpcAJvaz74u0CZ685P6ADV2n4GenWHp
oON4lWWGSHRVPLrAe+RbcYXBlXLminut16sesXdBA/PJIxda1wX0upc1+eX8ys80
OLHo9GXzvpiCj2VSQ3gbypF3WVXQOADvHyN58NEWFEj2hPh1VTDpBA71Jz7OaWPU
XllRdxLE1Vn3hig2gWA/WC8EdNBNPq508dSfIDLeXSb7xSE3dfGaWfj+aOrlB+EU
F1UWVhhUpRqR7+bTMqTcf9TIpvMfKxOSPfPKbSflKffZ5sP8KBYmjm97hUVRGYAU
WGNzF80IBsVbk1sUqAa2RA1so7XiKiMGx4LsXikn6XGU5l5zLODBRZ96U7tfx6fY
tOm86JtlRBluaftzwko3KRjL3y5V+N9YjutFq5gT+5KG7nHBey+xbr1Q3P+6Ovp4
PcoRsC4TQGHkLl48P3nxYeNTjvBvJ+5i+f15mYAGfd01uKVWrhRSo/gXNTs0GC13
6TwAzSZdQWRUYAvZfI7WPCSjP9DY9jzoIOWeRXfQpATKNfABCl+CzpQ6JbxTPTDX
EW0OlP2B1ppnBlq9+mnKWKBjmBC7Ok3c2WqU9FAdE+57PUNfZ3dJ5eQQgMFPfGun
7hkAifMI5syR5tufp4YHxM8WdzJ1InhnZVVR7K8JuE6Jv1LSrTX1zqGyD4ORuggZ
vro5hSiVmcTYQNoZXdK5e8Cvs/b0YG5667HmOb99g+76Ais/l7yLtAHC32aLNMFg
lgJANwcmg1ebnHmSbmy9KPHEQAeEoTmvkKgTUS8IQf6Tz2kzTuvBvrP1r41rD+K4
rvpoRZeMovH+J5Az10GBb/hiDHyJ46UHjoZZUQXw9DKRaluPX/1Gr2AJODFdxLut
Bp8yIZu8WpFY/sJ5AWijaKltzZwuJ5YUzYGVaXWJg7T7+dsPhKbwPsUK3O8ihs+w
yRGJggSM721MEJYqR+zo/kcxS/RCFy3A5sJXEODoKG66OXDUAlHchUx3JHRR6tXa
FRLfVdPCXU1X2L5SMczrFqotRp3Ai071cqcAsMRQAo9Qh80//eLkKJMXhogwdd2q
4pvRkHTBGb+ssCCggM3RS4dSsCToa8BK9nJuN9UDLeMrmUTc51mKzo/Ou1k2h9De
dAue7cDzKzG+XnDfLE+hfZ0pxQon7aGf8ds6nOS5XKS++Lht+DQD/+eEpj5XbVUk
xk0sW7exaevDMyNmFU1BP4c/6Z0I/TOsVKLqCSWoNMFswOX7GBmTGQGuZzoRzy2u
szzn8B91g1riCn55KrzsvRHo9qtfZDsbAiPz2CIYtSf2wjLFyiOI1UjBP2nkXFBB
VjBPVP2r91yccMHPmIu33az3AYztYMqW+kCadxEfpMOnGF2TP4rTvx3qK7/ZxR/b
2aSPjQSgkXreAYs4PXqN4BqTkOsUnJm1Zf/4wqpfGPLm/DfT22BJ+PpZip91rXw4
L158Tg3oLpkbmOnsDhFcFR9n1OPg+K2gPmjGU9VptsNUmz1N+BndUlQyQBqWjMbg
KDR5tQtXJvKvB+Sbdm2qaqmhbG/Z5OrMY2R5TBCOqFRFuXBTMXOmSsKnJy9Pzvft
IHPPvQ07kvqtdyCGD/fRLS7eWq6VXmJId2kJvg7ZUD9EepPxzgxwvCl0yIIs1Ih3
0NBxSFD0YSJdkrtTvL5c0Dk5y9vwQdhx+8s+IPxdcE5jZJq9GX7OqjwkRSCNis9m
1GchEJXdJRnn8AhPu0NylYNzi5BV2zgTm6eO4eoeNGCSBJJXqH9EToFH0xWr2d1K
ZtoaJedAGU++WN1X9fiK32SUxQr8m/YupAzUj7xbMffTQKDkrr45eARewDvfsrm/
4xfWgRGTLzx5P8oewU1Els1D3YXLGAe2xUM4xOfG7VrbSVDJUdmk2sF6lmP1BaLB
cCyVCZ89W3hqxAl0sSMQTPkaNn/525aQDv/gyDcz+ufuPChz8XbHg74e86ySoQvm
DfScmR6B6huQdUM6xOJwE9nCwOoI0XlsbExm0xpO46FaI1GsS1EfYFQiBr59hxz/
B2baP6XT0QcQeUrQ0MTTWiyOykZq2b2hlf+AjG+KmmUzvltRczYIOqW9FHPlit3c
6bkaHG+Jo0V4fu4EHPRfpbj9uzgI+lh7ewiqdGzNGjNzQ3Kyfvs0F8YJb/RYiIGm
yjdW/Sh5aoQkNf74uavEi+U1cJkRpkaPdMWDoQLX1pB5nG7Sk2GCKz4rIM7PU8kK
cnllJjQ1mbYnqqJ30BgtA1W8oCy9nv16IkutQ67wsrtrv344rObuhV/33PcEZrnZ
HGVl/znEuUzZKuybOzW0xXNUF7Pld/Q/rU1pxGmFXRJtOWa8AO57ZrKtUWIbkCsy
yGZYGHzFLDTgy2xuTPh1ltpIsW+UhLXNKQNMmre5RWEV6mPJXaoI99h0z4GiFEpv
os4/moHWVJxUfz1XQrAPAct0tse5MZArsDxSds7XsA89kwJSjjxtCFZt5cfuJn7V
QjGGeMJktx4EODxo74MAvtGdMG+fvLA67Q67/jf0mJLDDdJe1SKpeXfJFhzoFD1W
7hWIaacpaJEJvovgmqNXsXssNSZQOD1L5KC36aeJOn3cXXk0kpEqsrPwRkhY9kKi
yYmI68VsLzKvAUA0EsyKaZgqFvhBNYIfRtsGobktV+BgJOLBfFqztp+wBE1FM27S
CZnqIgwCBTuF6SlUNXxsGAmna2pYPNjMKBLXn/XnCSXxwJ2yopTVjQTRXpSAvzt1
iwsQz1xyVTzufiwk5iCNiHDs4e3WQ4/HhLvtlS5QOGvthpl/C+b+11NRZQifeJL+
uKoHQni/l65Benlb03WtA/FpiVg1liX3HAgm1N67Scgdttu65i61rgWG289/3ZNL
V3Seo8V2ZB3tjkf9vxkVgXVP0Ln547j9S9cmksMzuNZiJ0ISouRpX8wPnxLsFMxz
i0tnGnU8w5eLyVSwYDPzihh0cCmEhRNoCGlMGxsj4s5mSSqjeTJ1V7PqlOAvs7Ao
b9ZnCtMkCogWZssWCAhIOV+zuBl/RVQosczKRyCzCSUpA6p7yumf0eoRsANve4hL
K9j+/xkv7XqyENpnPGSMs9+jJRn6mYfaoqrxKxLodV3oPOjLifCi4MDQwTsezfmp
YLb4C4cuzmPTu6nZxCXvnTBMHvY0o+ewSkdzoeCMUe+RpwHaO6Mty2Gx1bazEuaa
gFQGE9HE22HE8sJ/DpNGEykfCSUQkzjmpj1TdkUhVT8dOCg4INWI0mmtf2b4tNpC
d68DQdmw4uJli/29hSvzLQhq/uyrjyz7LTh0al3cnuHFBBSLszq4SAPc50THnopJ
IErhVhyE4oIoutPbQ1OiZHuJi6ZW+8b1fZ1y+nE9MXP7e3U/+V6uE/WdT8QvQrV2
PbhTLSyhDFLps6der88/nXWYGuTuIUOWhODw/GkgporuM15jSnzUk8DEgJBgj7Hq
Uf6BNMW1e0J2qpmLAuNjuLOKj3+05webv2ZqpJuMO62hPvWwnvIpoYJTIlDQf2Yw
0dRaJuNIHL+qdaNPOBbUfTJ0Y6lnhkle6d5OI+tiZ4fHXq0d0YT23TUrPS+blTn8
bLeMcbl8a4N19xPDxGMgaDhJuW/Eqv9+zbfYohKxIoiXKEIcLEZ1CeTJ2jzZqacT
8Lu5All/qzSlRFkekiWkGxSQkG2wzSSqjG8/kn12Yca/7Bk/FOgePvemh3/5tkkF
2XsL11sjCGL5wE5TiB8C5L4Ov9go0MuCHg5uwq/9OHxrm9NeZJPIIky+EuvYkKTs
qZ4bNllWY/ueGW1DP/TlPSTf3e2alryhvhygS09EjA96fZT0JaEPSCz9gYvfXRRG
dS/yNrxZdbeMG+yiVUATsVZ7qegkaWPnuv87Cvic+JARAc1L+B01U5OHUx0Q72zA
ZhRE618OzOhPUPtaH7O/00Qoe0DtzdErC7yNdRnLqia8nrgYIrKxDsDxb2Yo1b3f
ehelwOYaV1vKYZxyuFG1kZbfwNX7gv8agGdYzLqDZ8uFxKsKLCJsi6rwhX89NCD2
5DZRsfzkT+eMmLnbKx8IXnJ/9YgxA2p6UbfmvhQi84uvUddPdCdmfQX6h0nfqkNP
TOl7FMRLsY64VX+c6WrMSQuE0aQLkr4BWmcpstPby/P5VZYRnXQKpPQXhNNwBG88
OiGvddcZ5jzNTsua9xpH244ZCZ7Hn92DY/PAWOIjzte5ASx6ck4lmURHVfOLVeyz
VJ1GSYweH9Q2Mm5K4so7gk4CXoKKZgkSdlO3yqkKFwesU/s+xF8HP+7KVWSYEf/Q
2IJ6N8jM+e3taUCsWpfGHrOgQU5qFGRftCyrTCH4iUTdZCQvEtwSCqSTR4wkkWt1
yR62ieeJEi7NJ3nvzjwLffak5a+r8u51KUe8jPKJMFy2QUQCkckZrYemLCV+9DNr
4R4xNN6E/OyTYrUAP3X0o/0kCvdSJSwrx2lVikPaqrUOP/SG6Iq8mhf4xm/d16nO
IPpzzQa26GkPdXxqLuKsrgcVGPx1PH31u+3khOZNooV27UTn1DdbCS3g5bflavSV
Wm+5XhFjYcrfQFXhBGHwvBwJ20bsOZKsqsnR2euCOYMg7iU5/PRH3eyrjH6qnRu4
5QaJ5oCDidHxMrSqxAB4cnxVNk5QSgHIbVlSZzO1Mrn+NHi75eFq5EWKq1Jr53Ux
uOqOdWefWMrLdMUHop1lokyw/5qLNAeCtQpfMxcxz2dPpwD9RLjnC+IKG/sUUxwU
D+r3mTmamYsJwDlL/ARY3Erg59d5MBXCUfgsLUc32w8l5bxm48jPGUY/4C9GCTx8
DrJ3Zy5qWpJuV3+ElCOkvvLVSDGv7Q+ndwqm+ewUzIvRPNvL2m8SRJd1NsPSPb/8
Uw9RAgspQIxd2q2e0km2KRQb6CigDSnjP1HPYTCynukyGiO0aLE3wOuHWtRzhBd8
9Eg5ZURnJN/7d0/MDr+Nxf/9YmLP7bsUSRFCPbIaPcO8SaUxSUyRlCFBWOjocLCV
RMKPVl7H3LSMrW3uKNIEhy1uqoiKzgzmjOUvSvq8xSWNHZ/v63t6amYEHSfnNalb
E52PvHONEr9QQ4OuBqpE7Wl0XtFzVyEyiNDVRXOx/+CjbAevz/MSS0tSFQB/zz92
gC+W3MRQknaWbXlvsbTGiGmLw8WAZTpSCy2Q9gEI/63akWFYSQO+DoNTAYP6F7Uh
3BzQst5eoAQFMh8bd9nnaIG0ZjMqX9yLUTG84GBdbE0LV6NHBdze8TBA5JdMzfrq
xHaN+fLIsbgtXFLU5zUVuNMDrqhd8H3pOGjJbEsWf0y43oEbH+kwXkU63ie0wl6L
ekf4p8r82j0ilJaf66cnGninv8DqgCtuq2KsXQ3MRnG7Os76j+eMVGhVVOrC8GQt
e62ttXcwZYA6PLuyARdeNG5Xp2jC46DiVyX0+O5RZgEpe63izrfuGOYth+8E3Jn5
RXtYa7GR7Cu9zhkHgZOylILFrEG3ksRiaE7sCbxH2t8ZEXIRCPx98MwlfPU0p++/
/IqvVBXhq7/pxQgCOwNs/gU00PdVmxfRZZ3KQyv42++kNiJvruHZ6Kch1TX8XQ6b
fFJ9N6sF3TS3fXFG+fYRu6WFW/jo3dDB/Ivu2Brr9np5k6+vv5SAP7m77qWY6WMY
jkHHQljXOyoKFEgvcg6XalqLDNPlS7WVIV5hZO2XB2CECKJzVTjoJwgjh6VES1vE
g+F+Ahb5YvazGUH9A5TVKIVUewPMJlcgIhBWBkAmVdFveQG2dJYfVueA3ygGWgsc
Y3kx2DKT6wZQY+QiXnS66f270wkA0HzTTfuY/7MT5Hu8qNk2+TA/rvMRxd7QG/fd
g850ED82GVy2KaYmpnAgGmEkjCXBQiRrQsOS/NXl5046uWTMjBGWZr9DNUYpiEb6
HQ84Ytl4p8icnBj+gTuyqNjbXG1RBbRFTtUU9lHou4g8yBaCdqKBAyWOw18qRrwd
VF50+T4hCkB+ugFSVAV6Pb0pQ3DGgWKIWZYvBYJQui9J99KEmRs3P30B+7d+7ext
hi6bXFsO76zldkNip6LOcLpva2YC0eavfJR0bSvJ88MhxeQnyL2P1HeCPA/9kdF8
82oPJBCq17+FR6EXaNtIOLruMbzYVrNlWwDPPDivc8D5zptQ98PlN9oZZLdnrqUE
laDTi6rML6RVRg00qcRhEOBIylHwHA8U77314xWWL/lXeA7JQRbauPL0Wpl9IRoz
L+Zm9yk1V9ZQJ7/3unGChrbxa7bMgRyCuGYLyE5GDrRXog83nBmTUGW9M6X+1jP4
sf/caPM1mI45tQtIHnnfkygFjh0OPygOoLsCgfRIBAKEQzT5PsJQAxKwWR1OrDrP
ZWi5P/n9aqBjQj5jI459096MkjFX9VDJN38TOVaBIZoFTGtX8aXmbAXahVkjv+HX
fCMHFTa8e6Mhq455Vrn28+xIAHSqLIsp/poP/Vp9OEkETFOY+lqXsLUVJAz2Lt84
5ramlprQFzjH+tdrbpLYxAmOueGcfnnuMgd9af1wi898can0Da78jst5XfQfUCth
XVpmWXyMxoD8WjxaDc95gZcwwaR1NuaAcN8hZy9vQVKtberXRAil8R15XMNaZO2+
r9BWpDdiTgd8k+xlDTlHAxhoaQ3vjEinkzRJG7zs8d350vVfMhWkFZxaCBISTgyi
4tdSplokFJU3M0NbXYexW1h3LByXmZKEeGRq5kn+hFRo1R9Vjx6Z3Zln2y5Isu2U
Xtb0GT2aKRmfxy/vey35nYUBRpYCSBC+nZCaNCRnrtRv53Velk+1NUClgDitUUQW
Cidi5oqkEZlEMsk1ivpSabOFES2yqsD7bFb7Sr5tvHcN+km3e1rLThBJ+6pvF02T
ZyF9NX2OVhVXR1FpBAlNcZDm4cvtIGVI5BBhYyMEC+YOMGzwwJSp2OAAAl3RPRRR
zNluU/w12HGfa8oByZ/MtPMTn6kVdfBKHpbGXA/F9GOJ9+TiR2qKovQvhQwZY1xJ
lTxVFZmNs7DA4wiqfaF9IhJO/LXpCO9EHAMhlwN69KYOUDfaBhgfiFuIH9ycxv0M
ORkMvXXgrD01A2LXHGE9BA5qPPLD4lfzvKoRTxV+krX+Zj8//Qw6tPBOIWdniXD2
F+nkosP6VB7BuQsWRpsmcmW1W+CYe4rG/UOrg26Zo7UXzzHf4IBiyEs00Y7YyC+1
3XC4jqnWessgnRtFDoxfJAqnvC0DnGAgIpNPYNN3PIxXb1neZOu1kQ8VjdT3wEpf
XDIv0DVX2XNfihzbjh0x8GjnpSsupHOcaegGV9+JY1edZsQatCigX3k8ACFs71DV
j9HqLQCYWoQO6OFUMFw+j0eMzaRHufIv/JD34G2bLc9wW0eguqnu0p4j+UHO6n6x
8oHGIjrXBpqwPcs9mknrdZ+qyF9CPfecD3Go3X8keZ0Rbnm85GUdSi/eGpN7R14p
Q8ooBmAL3ZxvARPwVr2K6RJcR45hRW/Ih0gN1HkZ+2xXDmpdqpPkYyCJE9kczsQS
Zd+U4afD4DHbPQ1LJYcAvrBfD/6uBBAGJ9T/W8DBOXKbVCoy4QIc1O3Uaf40NGfc
xnBl4lVIxb8YIsTgMbjNjNXnboQfrRetKc6OHUkRklrEGGcDdvTzBilwGhPKwwTs
W8AfahbCKruJgGMi1tKMHiTmfvlfJs7//DKS/o84RsgRf2B0xvh5rLZMoXkoG5vX
9Ii0UT6+zqNG0OZkdBILVi5OAhnbhDr4yXDb0M8SYulnD0oImJskNRN93H/o9II1
QTU6wDHQm7c0NJauKyzo+823OgogT+pYic9dVUulvKhNdSPaKaCGagJrGNDul33X
5QFwazoEVgEGYWlVJdYds2QWXoWOUp1FEeAyWsht9OLtHYYc2YE+m44xNvrOKv9H
cD3jf28jmmEw/0WqsMhPT1b2AuNI/NlSbfd1WQQFu7fk4/8oFr3KCrO/R4mBWo7w
OQaAAc91iqUdwRsT0+nIuAKjNkozEWoHZFX28tD994cHWR9MlsdXsHDeETO/49q7
tLg7fKcEcFES2op28E3BQVDW/FVqZrz8gPyloZlz4xQ7v1n7am7hxpo83jPmGLbo
LWdc9YTIw3qyazZTGTl4rCkFdAhuhMenxxUpxhROmwQySOO46U8oBdoq3QinLE35
lkRgYSsImoZAIbKfyf4vEcepHPedNvZdmffoYQWQ3SoICA1Dr2HZQJV7f/cXadiT
nuKXPIBFLoVv2mQVPToCEm3yogQXRV8FJu0byxLyp8YVGs7Z/I3tWivVTGRgDZ5N
XlEgmrr9Vj59NKCU5+Xc24HzaT7tIv6hcfB2tPw7r8XHu248wr9VSQ0gEZdc8P+P
GVynfNTVvJboY96xoPY5ATsyjmxfT9vb3XL/St70yBNN+LjGRwhNdiQP5J81EPhJ
BFDl22tqhR1ssL+DQKGmKprKAE0K3jRj2zwB6gx7RU3NpQI5WBYZWwWleG07wfeu
cGz80DMvE/BCyeEWQ0PJxEqTReat6JXEdPtN7gX69ZQCAS564qbDYgfBlQ0oJsnZ
ZpTHTNyeq5FMCVwfWBMLdrE8QR7bCJi8T3ScOsz6ZLMXNAAVqDm/sJJS6i8oaqrr
Ce/wzxN5WjS1qT5qWwJLuek7SRX2rFvRaPBITrrxLp5LyPKlu9SkMi4pfXok7q+t
2oN3RbL4J6rYlnw54zJs2fITLpDaQyQo88eC1QqirGrlILDefGHJ1bY3I6PUN46f
bElY+CnLA0mpdAvCA67OtzFCEf91pCp/f/cKOXHHbZfsa7MvuNY4DJgaRYje0cm6
b2Dfqw9nhSGjjp1nlp+kDY5LT4zW8CWYWtBKCVsU1+TPfNcSgp3ECXEKk4VJU0dB
fQZ6E8hapDfF4LUk5a9cBX2j5kRDaV8WXEiy6dyYy/JmPbAyAndyTkp0qmyDojhY
eIgeWaQi/eyxXMDHfKzUfWdY4cDwkBTRL//Hx1MGcqMKFx7L4LMnA3vDzcgQlLnm
PwpV2phcwDHx3iQ7ddWNxJMWODJAgD6JxI+pRvioo/FNhO5IegKR6K6hH8S9x6k6
eiElT2nMYpb1vG7jFNtH3StzkcS2mBFucsBZ2A5HGXZ8zdKkm2g8Fuz9TjB3ZgBi
jXdNBffzT//CIfiFtVnfG1RtWv87sCuqnWWlSUxG5ZjMvQF/7BfEvO0whLoW91YT
Qpln2OhdSCl7LwegBWCT3577RbOF2yzQ7G1uErTfwTLq54t9lBD8DQpqGvfmiUie
6qQiSxp6f7FYi7ufXq4pyN7qvH2/WOKJneu13DF+Vt6G8ivGq2wZaCLbWboUnwJ0
GX1qYRDjiORvmB2h3cEaLYp0tY4gaHoTTX6N2+SKzhkfVxUdk45nvgmzIZKhIWNo
0MF7DkiQa3HRg4NswbSGlm1PJZATo7JzFn8j6Xsn3S3lDfKIoK22yykc2cExA2AX
FBnkWBba7NMXwxqcaYFkFHF3y4DJoHjnyJpCZdHjmuNeVQCljb4X2djOoVzZ2fLA
8H0vQ3U8cFaXxO4c5JwF2nwB8HblGeVjUiKyoGPVK5zDc9EsuS+VVUZe1W+JqDrB
IGFxtFXZ0LATwqHSlpHf5AwVK2O0XEiBokJyT2hhU09sHmf6B/rQtbGAUk1RMsHq
qpVYe72jjRDcJMlra8nWsDl8onnMpINUr02pz1NWlTZFIyMLUUX1AHLix63bBQuU
mY0Qov+f3FsldDXIXmtVaMB8WRxb+7y+322/oRQoldNcTz/6N3hTlfaCnEKlsR6w
W/dPeQVfmBdgt/35ezcN5ol31xPoO10+cK5Vo+1Pa8hWHgGXcNqtQsqYzvG6ejLH
YIonMbH+2ftmFpFaPQzjePmEbNAo6Lzhmh1gm7H1luDCwtICRtQ9KcZQeUJsoamF
J3HNOsYEjMDojOJKyGzTIOvqWcxuq4H/uawNd+/M/X22JbUIve/74u8XP988SH80
5jeec1j9OadWbQve1yUcu3j1vRGvURBQ/Q3WbMfd+rJ9g/Pe+XXeP85PuoEgktC9
Yh2OS2/QKy5PStfdiESIC/KNvRIUHWpRIDinI5gYfGaOZnvGqW5a0k37semTmKcD
34Dle/Q3Z7b8BK24hNPrlfU3OduIvE1/WwJFic6fKrWJOXoQgC1RnDc+Yy/bJRcu
L3jEx2dq2URNeCfrbAvMNvX5x0BDksEuNsSCu61YHbcTR8v8w9LzukKKqAy6a/Fa
PL63vIHFwPpLibCyTnfbQfjL8VNbqgV5AHtD46PhekW/82eEfi15Bbr04MwFtJcw
4ecRsxtnAFCFkxUFnZhVtFRpr9rLx68oi/XreYBdoScn0RecXhpxFLYY5cG/3Pc1
rgCe8oQXeJLq/Sc014RPsdjsVLNprGNf01IrFZixyXJNqpPbspq/NtBIxW1d7Hss
0i5Bo5IxliAyRMSDcOiD09Ju654EC3u5UtD0jpWLdbH2VpYuTdCK9Www7bwSUOw2
LDZFx/fBn7ZPKqACQSUoag+0uCISlPemrgatguJf4W0T7TAuvUzRgtS32I2vrZG4
DYy3+Tg4pdJaNvpZrKbxIlXrj3iVBUcgourUlSWCgM5i+bBz4aKwdH76jTs51+GE
gzmpbGy3U+oKHxdOhNTuncYwlrLMp7FTwql0sPG1BMQSG8z46B/U8zCBUqrs4ERj
l3n1CJTcHA00qL9LBrpCW5K2mU5gR64zAmuYqkkCFaOeyptLDrlSuWTbbc+fXgYR
eQHhZBBErdat+UiRBwFelO7JtJ6xDhMnnaTjIzVRb/Ps+p3P75qZbudCYPw8qk2e
LKbn/yrDe2qfrp9DenTv+Vw7DaY/V1IUNKHIci0YjkhuOV4dF9Jm+DCRW2SZtybe
rtDFnAUNfclpgBN3XWK6J1m+CsD+8XgijtV72uh5rGvIx/bCfwY2Z2mInnHTiVXZ
PNV4W3dl3CUu8vys8xtmoyaPZtk86xwBl1AvbRnyOzG076B05OEuhHgCbmFCyVYG
aLXKmjFGK326EiKeGJLCloho9zwLTRhbSSBNvIWFKXcih1S7+eZfQ3FD6/FC+tzC
RnQsqI0vWsQLv21r1OvKiHJp747KLRuMkuzwyv+fEHojUKo0wkfkOq4jQNB3NIfw
EMYMPxuo3jt/i+R0chVmuDhXG49+k4Wnd3y1roCM93KQErFKhgnC3sZkjaO/LjiL
/V/D+wnIb9jEg0tk+QfN/rqYsjQqszu4xUa+AyKzAvYt/ucunm/LoX1tAfYuixqZ
jg64rFlPLFbB/JxfEwA6DZ786RKSStlAoGXrc5pZ50vF5OD4xGzlZUIjnv/yyi2z
j9ufz25kZhKzcsLkMxsOOPycVjE/DXwhWjWHgbIi95ZML3Ou/hEL3k3x23L+Pgzr
10IilpU7ZKbkhpqc0yxAoxI5mvJzDjpIKrs8PQIh0UF+WjAkyz4X3gE2Uc0s812g
9d17Ess30ZNHzfVExAl/L60LCIg1zGTDDdjlkpLA1XSqw956+yom7mRbtd+kVa3N
KYcezLccglGH+Bugx8bnzOz5Ey7E3omfQfVVbxNdTRBZflGwU+hnnappgfmg4oxt
fDhEN/qPk2haZIEq+skiRTfuO1yRReL1D6pbWLXXWeWYp/gujqC8zVRCtzgT+VFB
rvRp+qVjSAHkPSKaw0bMevJrCwW+GvcO4gYT+e5Dc8q6ALBmyvkXE4CagXg/tr4x
RSe/UQYQgHqGSRwTTCyivnU0M6Hvxyh6ICji3GUwZ7H40jiWiwFSluh+74GiQ9ve
bbltWpc/fcMwqOYOwv7ZxinZIEui1uGnHLAX4+3uTuZRMPqso26COmxpkY5eIisY
6ELvXrYAAgTxmNG1S7ZrTgu3ma7kiQfz5bsvMLaYq/28hlDgl9oE71+DWbWDM7QL
HvmzequV9hnsSoM1mKfdTlXlW0r+83gSZy2NX987Y/RVrOyOTfTJ2MvjYgFBwcCW
y1JEgmxOe+FL/MNymNDLnH3HQQZciI2PflpVAH0l3A1nnkmhH/eqRk2GPwF2uj4P
Ih++at8VXZozp9UNBJWdWfAoU/0SN7s+EwgMWnOlJL8WNEjZkrjJ68qkOl0+YxA8
JMonV6BqBYAiA6amOA52uGOVAN7VXmYaIkZsHXpeOE2OpnByr46YnXZS+r5VKh4Y
bQl6CNd3qphXOzv/J7Sel1ON4wznwlyvmk7KsPI4I+65Y0NXfqmyoYeNTinIDUYh
Q7gAh+AocCUGTTUfcXnJijxCy5B/MPzRO8GEwxSxP711/KcILQwexf9GGCCWsYbO
QTZn9GYRQKme1ZypenN6SS1paz+uzdn/4Hq7jzeqCJ2dAP3wJ2WeFoXyVVKhp44y
WnVBUcYTYaEsu5Z0HneGwvXh2EopdH04OYeKtXyntg3xWgNRXk4jhNRpba/LdFmA
9Cr19V4r7jAW7A4+tP6Ev2Zs4xPFU509YLnL3M+W0DJx0Nr32qORjdcoWIIwhH/A
yR1sG8QH9C1WdAY4l68opc4UnWiVOz74llqBI1I5GyKDoAt1aEarQ7ZpcQCJaygj
Oo6wL77sxsN1glgc1KwujMt/xEr8V3tDCeSedQK11mI5NPkRllwAzEEX0S7Fv2p2
ChxaifFyoPRFTFopulqYjMOJUkYiZS+8rTeMpOunx0K92uyDfLnnCOUHzWhO0Vo8
VxJ7tHDQY66uoSHE2MkW3klM/cA9STPdZAwO2rD0nsI/ScCcPN2QXiCoZbJHM0U3
56zi7euQsEo2Dz4SHmCMYad6ZPnkN7DiUZlekgi4FCP/eYT9flYgzeBX0qgtr5bW
4x8VglZAnWpj0bQiF9XLFteS9R2IYTOJxD4WXdvIOA/76kbzYU/jXtxypKLGp9RN
3c1zkwfLFu/P+d/Z8cCSa80QEgtRKwlgc+AEg0SXjYTURpEFfGmCHWG5BHFKYKZc
BHlxViz0T45sOxB4yMSc6+OMLkKiCIx/9yOvQ4IHoYnfiRx3tbvYu6waQXjE3UNR
EYScW7qNrvYXI73MapH1W4u3YmylShNiF6z12I0+zIKskM5MwsWXxyMOxamGYNnV
v2d+S4tVlK6porwhsO/vC/IMiwMZkxVvZB4jOnCJHo0+eNbC0spkevjW1GZxJtux
GBbSrxSba6o5zkuSs6n3aWtZLgwQAq2MuekrDaT08soTJ7BHZb+aDTNkkv0m+Kyk
RjyMdkL093Gybf/0M/CWWHQppPB711sm+9zT0nqSk1aLEDPC5tzpOW6Q/8isMNfu
2ebMA6F/vSyTBSBCemqtpr2QIXRa8EvUVkAXT09ldyO0iVr5zjPR/rSSGiCqH3jr
aM8qn8RGphsriCZvDvUrroW10JkiUpiM20oCK0140eo5Eb+a9QjLvffyLz554S1b
qNunSVxp10wDFF9+Gm0uOpauDq9WchmVzDde8m0QgUx27iozI43n1+POoWXbjsb2
9vDkcxgFbjdxprLzlK6n1+bJHq1Rf3Yg91TgiU4hWGgSR/QqRy4Wn7SXkAYNPsst
djsGprG0072f7lqPcCKiHBSnp8k4yomTEWPd7QcDPJY3ciJLfx3wgu0yJMnmjx8X
UKsP5u4x3QDbrzFuCwZcHjWPADPoLIYqejTRxXSI18EKwlLNh7M+ON0TSBsdr8XY
lOptUcOGnBw/67OeULexCr9Q7ovxkDu5S43Fupxl9TBm0UToGn+71U2oaunwrDdX
bLQIo1RE9n9L8l7OMH4Aq5ba4rudWLj4mkn3nLns1z/C5mRjF95eoZA2cbitgNAr
yuGX3b8+ZXeQ0glb9fmepWupec+pLhx1bxwXIxkjFLKa9EkozD42UEGHbUQCaFG9
1wOcXA6VZXizqdJ6AycBpaVjFOJn/dyFOnvuLt+aJfSR3jdcY8aQtjvdKqu7O1NU
1z9JHACQERLqztleWCQrla3LVQ8z5qcv1wpwqQi7lHEGAuavz0nszia4Q6H+lFVY
hk1dQwYCvwMHZnOWMps5uDQrii3Kssl94z6QjjJTR7RkOqZn3JvDWgMGEL27MRgX
Xn6UQ9mD59bYLenApEiKQTF8LzzuLZIRbWrWT8NJcIRgA6Em7hhqbb30pAavDGD1
rfzRSlqBq1rxyFXfVuRUTvVdoGzk6Tc9Ijw4KyT61QFl0BeO5zuEa14uH97DkH8H
ayLTcV6xHffRf5+W8yG6kZskv5HE6zaQxqQxR8O6+q8kiLgbS/6wJJXOGezPWbOC
BtrzDnBRYzg0dj5s3lSV8JNjgFMvGVr9m4pPkb+HF60u8dJ9yUp3POtv7UZTYovB
Kg65WaCwQoMH7pUGLu/LToNmrhN3GLWmYywkzmM6m3AI6tjs26NtuWyMTtgQEyke
2jwsvCJJrGuYUFV4jHo1V6ytfQ7iIUD3XKYn5qhOlVtkfc6GeoUfyvfDWTkgofWa
2W2nFgJrwZqlVo4ivTQMJ/LKS7Wu2GtMJisFF+aQMGqSGiwdVutcx+HdBkXVbb7k
nvoBy5NYbyMEwdCVyz5z7RDYCivLsQNCVM6I37GsS4u5zn2AdmZ2dJLTVELpTeEY
tgOHTbqESGdvRwAtCBga+neIT0KMtudZ+J1bPbRi0H8yj1x+cMcY8w1Iqle1Tra5
FzUDIauh9hWODGE38/c+A/cEPQCyASJsEqwwNkS4LdvadLwQ1fPPw4eiKPD1wfaE
0p3HyAVo3pE+PgmhgkWMsqVDE5q7C8FDodVPROjrPDYWLBOHp1HHl2RBaTIA+Q4I
8Piqc42HImFZkvR9fpptlZmzzqftPTV3G/675sGbJ2i+C9ZW4/MfU3Glea+jpIA+
bvuANR5KNGpcztF4sVMOIg3oDB9SQ7xaFORQ1KObartUc4BUOWWmAxJxaoJJ8s16
/Wk1AcfLtHXvg9W+XGU81u/XGJZKN3YV1NkxxMZQ8BhclSyeWlSjENLtFuuC6HUZ
eTYChua/s4/+Cl/jkB1TuQ4BGyyKHctyPeeFmm84rkJ4pMWDRzAipf1jdrX5MOkE
ALWLPQS6ebsfQ0p53G+aSh04Q99CdSL74nDTGQxnLBMwwG3n0b0UE0nI3NEVZ9aW
K/r7QBA/dWIQQSdlDy76boCvkSkuFM0Q3Z3x1C+pda1iEIQFCRoLFol4LCcSrnHT
RnlYoJP7rUo08V4WWRB1vC/arjOYFBEi0WTFtgp18ugIzjyhznrVXxyaiGSHCWlx
BvZWsGvxeOtDm72a3TPs8id331uBv5MzWLhRMOlbtpdC+f1rkqa9+MIgL8ug9dm2
BLns30qGtK+5B9VTPoD6QQETf4nga7gZUIuTmCKGwTTEeEoSA3wuog2EHCF3+6y4
dtMGbwK0etoiV1wpBI/k3Cshgr/01/LUPDhFgyfiicYmXAuADlF71Cn3VbNGdulb
10PjrwuriDS4NIE0Ko/R0QmSwCN4ZlzLgOGl4is++WbWrr9PENNCADz001xuVKws
jKJLORE+Dve3u1pmdOnwFyCBIfxgAHaGjAihQOw8SKs1eYy005o8hBBRLvb+Qap8
+WcFZmo3hcdOCayA0oausbs3ue52cIfM98oJ+781WUC9iyqXPpZxC70B8laY73FR
UUxt0UtqHs1l+U7EhW27aX4QqZco6aJ/nYGCzvlXDaUJurak5J0oB6t6rh0Jsgx6
JV+Yn2sVFUuFAVVRX6rTJ15Wx4/3ljsaOXmKnFjVSv66WBt+g87Fl+QsURbf9C+u
F+sQUtKvtdbPzz+EuGM8lqBFA9mk27+v3CljAr3OP/ydOsMoYqTw926rkufQRNXZ
K7e8pSgJ9LDPhzREkUZz7yO0GFt56rZoSWcHf3ohsU4MpH9+p6bYOdQsEK4rQupm
y3rRwancDmI9Nz3DUw+oeJXnQ6WfEa9CtdBIkR9bu7/FzixSd9KPakoENRC4LghG
2jLwupZag1r9LRQ7POsDyMrUujZ7oVCUQ08r11pxrZVvc8C9wh7GCBzKDX3iopTh
9+xqIJMcA2vP11zVhUdObOoq4xYxr0aw+FdhYSYemIfS+4E04/wsvj5+fx+Um/6K
cYNOF2qRYX1kLBHAL4Ft76UsDZgt5w4yyN/fpKo9i57Pqir8pt1ptBdkXaCVjg/8
76bRv48LM3BZj36CcfQkalkHRG02nIxJlVwjGe9ame2fM/10X1EVkc6eJ2j4rRZU
NGDzbzCl2HJOg2xze+cS3ejNwRVPPFPQmTczlfGYuyi1KcgpZjmF41yoIzEPjWjc
Y3xEtGBfHKsr3mliMuKSTC2tw7w+gKikrWUQW6JzO6QZwUfq6LRvC+Wev1NRxl7y
d4m2leduGcGONA9I5vp0DQdy/olwn55EK5B9MGPlpvyXVkgfF8isMSoNj2l1qCgg
7kvm/Pmd2BLtdJeh8W35tBsDD5P7KdN5Y6VwZBAcKmLrPyOZ87owAEHrNK6YCn11
lcWoap7yfKcvsMMYw4YSvMXdVd1wj0ka3zYrWZIlfNjeOtUGTsWhnpLAMP/x74UC
Ar27cqbHBSPOtT+yMYheW2xehdvG/h1Y2ch8xMVtdvxMadtVg773ClxxL7wOsuxX
XmWpRntniTcuDhJ3y8SKk5/kRZOrUWv1tXWv4wD6t9n9urCxjpshYHAld1c9RqPx
C3FRa3E4MaBs+yCPCs2cqxONdy4NUl5ewrGJVsJG32deW2Ls+mfdhtkB/RxgvLjK
JnNG0eKU/Dc5WuXrSOefQLophyg2bE7BGsUsTQqihJTEl7CxpYa0Amzex0S09Rtr
KdhxUz1IvOvZju7MuRpb2rsuxXy0YExiw5rrs9hMvxwMbyxgP0e6aeZO6L/ITcle
mLShAmgXSQ0z7Bt2UWDhzOfBt4Fcl3v+ojuzzlywBCjLb140kBP1ACvuRYr5NH9e
ignp6elp8bPXSctdNvC6l9RvMlnJmZNmwNokfjD4hXy++xE31MdV0CsQs9CHVuS4
6reUCRz7J/22qKwa1pORnDdRsYgpiyef+olqDmoZ8MCFh5+Hz3mWQWPyXhmIGRaD
poEArE8GaB6aIbqPlB//4XyMwLBq9aVHeKTfHCJQgnmJBxFdMMS+syKWKx0PXGSn
cjZB4p8E6mtBtXceocCkMHOSNzJVAaNhWkXimfh9uY9o5rJTWi3wmoOivI+wDLzO
L0/kw87u7nOiuBGVjDFHwEROzVXoWqczf8K7ijcLVBr3B/28ibMN+Xqk8DMsOj34
WQh5pmjkt+yntaRYcfXAnUafmp+Tt/yHzJIpAgXUljIXhNkexxJAVP/AU6BWAs2T
9HqGkThZXYEcJ9m5vrhLwGX93jggxjW1vLspZiJLs2ZQDavhYpTMfCCBne0XFUJT
BtTqN9jgTz8U2OQbyGc7NaLobdN/doJF6s+YzPardPylHcTPTczWETv3zTwHaI1Z
Xs5Di2rWgumyFjgE/SudDkrf14j8MMYLlywczKC1I55dFgCnoVgy++fWerCRsJtp
yZYB5dFkQ6TOa/cTnTXl3cKo7J+OqHUqhJw1CsAKTKzNgkkkiTap5RYzFcrkPAci
A3XJuURSWC/pxzDeQ2R3NIoyqYVFHGB4ypQSnJLLf+G9RJppxcc21e1b5dQHeDWx
ZjeoT8hyfaDEX/0Nv9smdwqj/bxzyRsoL+R1PkgZH7pUzZxnGwPSks2wUUyUXFMN
Fv2ow3UQWDeGe1U/7Lxj+dKxzYLG1b9U9dvXyT+4/MKhuwFq00IRejbK2ZxMhJHF
JgFWjrSb82veUoO/Lpe/NfEFySjB76FweEHc1Xau84zjDeQPFyqEgwZ5ptZHboEi
YsuYDDQqT/gkdj6bjtwdSJd0/nN5hOFhpOisIVhvUs92Gg8D+uGgRN1Ged29OTG1
P2jtI9orgE/q80SJLr8Dn58KJCg2r8NIuRsSwVheQkPefnMhz4QcXvYg5gDGRQCW
tIf3J/+i2KBEfzsVwSIx5sB9QKPyhGb10XDJqxvVz2WzV/wHf6lY7UMlsb2f5crb
7D+m09SHtNAyxCWSN/a2gwABPuqDza9Fqmk8TvvVNu6vhiPTYwfbrw3ukw1CqBon
NyCIfNmEKmu5AYvCmeBpuRVcDy82f2wGywY8nmsD0V9FbGxFOx84Ziwto+kvOKWj
qfXNyEDVHgrx/lCHnNinoUANhIUZsE2YpoVGS5URe1EH9aSMdq9Wo/RvbdWw/drN
brL1rcq7hKBZTpk+URSLHGirEjK0zitwWLe6t++nPmECwo9y78gTfQvNr3iYH/4F
bgi+niGKXhBA5wFBLc/co+cvaQlyLH0TEn/X2top/nkx9GfLUa7oJ91djGJ/xK2y
aK/CqHOUe1vZsncSl189HPXZwd7+5j+VxAuwQDbnYPBXj7ihFS9P1ingx5Onv3Iz
6kRkiANofTniPFyl6Yxnj3y3DP0DDeDYv3rE5fBYSjDNGpy4xWAtJeyCMbDo5aFm
VZxdcrjOz+JygsJ4tX+RQS3DABEcuLOR47JKtG9yuTif2TIThBFzkuB0lqpIRt1y
8x8Jak94UPyPs84jaZvBtKeNCWP3SkLJlXG9Nyr6aPTVa+MQfe0vDFvXoIcCcFo0
yT//KMGYYl9y1H2by9ytcWHXOmD3TZb2vJiE1h8g8nyGjUI1l9YiVL9l+3DCkwUq
5iF4hEB0mMKM1N8faCl6uO4tOXuSoKxeFMlsDSZVan/WTNf89NvFN8he/m0PcsIR
d720QFgXGtFICzviLymaN7H08U3DuMysncBJLv14RcJ/gjIPgaZP6DUSMJqDZ+mx
PWpLdZVh9kDVeLIr2FlU1POa9JDRP7tdBKobbedOILcGIJ8RhaPkRc+2UJSCg1n7
z2X0gMitI+SmWOo93j4YKTP54vMCv9uadmWbqMDuZmNwoGsmOOPsWtzXcFMN0RP+
CBVNBbzeRIO689kn8bNXSMF71mlSVkvD5VN6I87kpknS0MSOioMqyb5DAG8NdIfH
jqDZChzs1+LpJXxdaTBFfvRQWmAd6b8s8ANsd4r6QGjtwZeQZXfa8VVZh7aJMKwA
i0WkWcEYtLv6w/4KK0zMkNFQI1Wb8uu9VQnYafMv6uINsp95I1RFt9cgxYyFMBTj
+23c3SyUktW42L3HIfkahwwyB+9oskrmpI7IZQOCQEd6w4nBWH03DXaSn+y+Fh40
UN1oR61ZFGy2rFYYbtF9MPTbBXp+3L9vDhJkrJ++nkjGIWpOdiSOKufrc+uGiqxn
K3SDCFrJCfNZdiXTL8vOMrVtxSqNu1tHRDKqdS3RgO99X7oN5h2TlPRh92Itq9ad
WvtTq8QAhScGFzqx+NXDdQOmwRVnDl6RZHNSVGOKI3tlg+BzCvSYAzG9nto4Rte+
ADPVLLlRP6YvPn7rh7SBBEA37FTsI4Yup9BzElHanQ401uRmtI+Zl+tYbDajpaia
c1TEDzgfVDVMGYP9QbI7hJNpy1mUAsffdqBTYJXuRQT5lcLgjJSzlsPMqxXnmJE6
gSX5n3FnMmT6EevSl3rNAOFXi8H0dUzOmbuFlr/Z1s440FTSX1vk5rDgXDNoMoud
VKwmykOD0QFEvuhobW6GXE2Qn/8NqX6nUYqB2MC+S4wog8mV/drH40TONIWeBDcX
Ggaj07u8ToNZwWy91xTTDnoEKxBbEd5bl+o+je4+oS+TG78G0LtO1L9WpxAQMWwH
IQO/d4aMSCFwEWGrU+Jh5bY5HYna6aYBUzmDHdQ3THYvZje0sHXrW+t2DPigv+14
ubWas9f7YurUZ/McwTBaUtkS8gq2HEfUHOBgaM41sSFlhEfxItdQBuijZbFLPkNm
9QbdPOb05sb27GAUd9vnOS+nLvzfee7mUXGa5bwPJK6HeXorivZbfLtkaug80KdP
7uHHt88m6k9zRUFaelVaFWEp+vwvS7h5qMWxNdkDAx2bKFoul6eBCIQ//tOVbK3w
s0tSIu2l7mvbS0GhehrtUSlyJmhvNBAcxSRgADmaUC6Gwzid6+xPkIvxPQwb3j7f
d40reznvtY9Kw9kFz713ZVOhnVCjd7ysGG6qzLkNy9P9SGjV4f8sr7jMqox78yp+
xCGgBnOVQBvRwkv2HnQf6XaKeUHYXpCyYRP5E5DbMZ/F+J8IpvXoSIyhjK2RPcwy
Uj4Nrtkw8AVO+fV9304gAGXKHGplCOy3A++k5Sj8JOATySa5Qw0TJeEunLMPq7cI
rPZk6pDT+oWsCoZCmHNG9REOzcePollI1L/4VU9pO0NMKc380SuU7P1tPSuRgjUP
xVLKlICFQWlk041xtECWHV6MM6PtBT0CLYP33JNlS4GgC4Z+1NkaGJswN/KtaIL6
9ox5ol1o4QQHOaxauVfoYPot9zM6p9EuCD4oDiVF1zCUKF/6vI9UoBGebOj8lV/D
cOSStwpx4f46r1FEcjnkwOkx83QqnY7QFoMoJq78VkzZulr/QISlgyopgwcFgE4S
XRGuiyk1Y00Gnnewujj/BxuxM9GyWO53HgMGZsDOOHAy3SMT+SQNsSlqMoz7KCLi
wMKuKDRaR0I3Kl+AdVXC17XDxbI5gHssY+8rvatwTwOwbyTbEd4fhACNn8lf1TtD
3hDanV2NYUfF0c6pYWHvlBenud+G+e5GAFdP63b1kZ0zXAjQ8348wdmSgRxRg0qf
6od88LpqXbSTBr/pmun1UNXqBAnkZi0+WbKMLIHVR+Vnx2a1348NFhmwBuYy7Y15
6ZXe1rLFwHcGDX8iaXU7OayDfMoSzuRGF25dSY3jNoTZxujhUBCv0XXz6FL0vFhh
QILw6NalcQ42IJDJW5N433/qvLX6NaIx3IvzdQzqRh4ZNQMIE1GdeyPKG8csWhlj
pMDOExIh6D04R4+oVIok87RWWrQ4gWvzA02sB3h62KolS9vlBB6mYszqfetRrRNZ
xFbJTy19JBNDLKCRi5Av4gCb+gP3poLPRNJ8Ss8ILlmUzdz6RPRwiEZBRLYf/Rnp
jwow8YVF65933czjEDxUaHLbm9fFLeNA7uzDSSE2YbflWXv87/iqwoqkUP/kmvIX
pDB3DWFtVFGoEvgqOJHXtNscs1Ac5JBqre2YsLyLYJx5JNK46dKkNd2J8JeHsZwu
nIFLE046jEwW2IuEx7j6voMFwlLEPuqxbPKe8cnUU8GS0E3P6SwG6aaCvlvhgA72
Ktplj7lpt9bYCC2zsAB7stHqAT7fhT3xBVijBO9rFkGumEpezMoB0uc0BDsEp44D
ebppazvn5XaGWySvxgKjv0pmeVSj9KhMbVCZDBGTBWeAMTIoRcFdfBsvdPTz5wn+
YEkyXGey25Nk2RCFe139sF/jBSWAg3yhR6nSZ2YpR5mhkz9mKMmyEft3TAa0WW+O
pC0M1z9yYuqKUQy+HaBNpo7M+IFvYhtDZohqU13A2oNXqVC+riLfjjIVq+02nKC0
F2MCyEWJWQdDDnCJHrDsXmVTf+UK3whxxNT1Fv9tzubVdZFhGb0VhegdjkXhzaE3
Ev7sDG0DgehpJDPFhj6itBsyLoct5UthXMGNLt3P+3i9Z8kxsKBi1EqP6atNwOG6
7jG50qhAbAgy9pQvNFgOs5QA7chhu5bMxuUU5vgAEpXVubMnnZWd9vOlbmk8Gzcx
UmUzOq6ET274DaHr+JteAwXXg1TaqfQZGNyUAgEEf7nJPp7pNrU4ejAhTDfEZPOi
3HvWt3cbRM5OJqhVgSBuO+kouJ4xLzqo8XGnU/EUoFOjyx0tZGm1oCScVqwaIvii
B1m+SjhZ0lUIJnds2IG4rG0EDxN8geiYBo15F3zX+D0O0DIIBTRCa5eyB6bwzaL+
mvNCDP4yuifcHg4ANKS5pYtTBJ3CfPnItj7+jljUP5sC06vhr7b8yd5C7g0nE5bW
0ygqfg0L5mP2rLY27ZeWkNN2zzPhJgPyNd00SfWlgxImJwTAOkWdOofQHJE8xwp+
5vtv8GEMVXJrwR6tKwJQ7JrNnI0XPYrIFBzxzhWuU2l4hhp1l4XXmNG5n+e985Hi
NvHtJ7Vxo0rY1k6uAA2V0uoUgf9NLqdOBOLo0pmnUjBJ8KrS90WwuIbmvX95ZTjH
ZVS3WW70owoCXmjNZtwJcLuOWm+MPnQV4WIj8FHaqtO/I5XF8XDDiU5xP8UzN5li
aPgvAsKBHuZyFrlYykglTy9qRxAz/3Xriez0RggSI/k1A6wPuOnGfKMPI2+SnTAY
qC0FAPIcAq35RLbBc5XiSGsGQfZTcsmKCWwg9b9J+5j/RzZZ+9sHmZNnvEthiXCf
lbX7/Z/t4bcSHlKeOt49ahWv5mph+DHJdJsif/6B8xhzfPqZYw8ZLXgIfsDgEiky
lrpswDcuA35LPA61TxPvYL8uxGwlKyAXIRpDL7HotodXbm31koBeJ2QdkMi3zQiP
QrivKCAueeJrjnEiUWuALYIlTfs+l0kOXfxtvyaBRTcRBxfoWFx0R9S/4GSsQFOF
DfzaQ7NrFEzjubrbnmqGCpvXWaGy3/zsAfywKkJzsFpjKgwKKEBkArxPDcvP48SE
lzM9H7Gvv1d933H+6Cd1N47K/8LTb/PKyaCEyYkKzxRk9OQk5J8bL4m95GQN7vAS
+QvhSJB4OQzeXGd1rPYI8PgaZfMEKQg3UPJV1+ZaVbTCZAifFFDZIJDnZe98CCoB
ZcrykRLBYuVaHsQZUyphSTBpSdawgVXglLe7e5SAxpCt8TptpXB8N8D4MP3jPxY0
R03hg1ZsF4QBESeUI4/50VZ7851apGlqkyVmAnjQiTl/7Pg167Ji/oh76Pi3Rnjm
QYjzAj5MRPl4pt5WJI37smZu1udNRYIbOzFziCtFkTgS4L5ehnD1udNahT8eubdz
ReiS8xYyv95ofCmeA4TsB8XmOC9vS6jM18TkK8TMfDXIS1objYxwy2X74FDfECli
EDeeyMrunT6ucBiT7qqU2Dgi83nY9raD3nPzepYkBAPw0jluofn8ef9EqnAKCd33
PEJa24Prdbkn/WyHs3ltMRR8d/ei3lqLosliK26LQKc4usmuxlwhQuMRc3+22yRX
scgytc4kv/n0ehI+bqR9HIrfb1U/2f/2ul3heZfs912BthQBfhxSxfoeqh3p/DlI
PLTK5nOH3IZogi0oazofiy1lG4u7CI8dMNfmzKunhLILEJog8TRQu7/c5Fi8lyZC
r4jET9AK19YqTBvQx1VFjMvpWUxmJcCBHc0mGQeCaEOFmjC0ni/MDBPzI3MA+6Qr
5r6IoanpvbTOsDdfKKY6rUmFkPvcLWI/iY4T8jzmJD7kLuxw0hkHzXifc63/jb9x
0Rd8y5J/wv1Z+/IDcY28mn7ahc/0XVCgkSBMuJCqD7G0iOiVsa64P3x1pTACDJQn
HBG2cI5dlZS+Pf5WzYdvjN03H4VMjToVkvKE3XoWlpvhxuMM6NUfHEI4xM3BSdPM
mOOhyt8FXZcp6Z5bg6iWv5iOyMl+2zweQjdhUtKzrwiRmKIfSHSne7lBxD8khrIr
FMny7E/9ImBaksrrEIe3Edet8J7HKvuctBWn3/SJZalHvVyapUIOK++adRZyMF7L
HbqLzAm9avvSYxuykLBT3yOGWOOd7/ibbPyRuAIYGBYv+Tqh+Q1XaVB9lGPu3CVI
OvzfWNTWtJTcoOEo5Gcc4TrLJwsbRTZxI400CyUtlRjD03h1zDhBYXPh9brOEWSq
TtdgIjv53hDl7vMRpJA2/93Qy/ZQeg/NOJjet2jge5ESXVOPoHcdp1MRZx05PEm9
ZbVvlKf2oHCR79bMq2SdvrTLJXgvQhaX3auZ/tvYQqHUuQrWQGV5XTlp7/9FfHsi
rJMT/tgfi7t84H6gXi95n9T+UkIoB858AnAL1w+q0rVs577jyz2RkWNkOG+yeWm0
7ByE2/wYyVmSTHx1NVBRtNu9X7fID6BX4/gOB4TwOBVDRvAl04RNQaVhnR1gtzlH
8wHwns2zRd8nDLBnBtXcvgYhSaj7wUNW6HFTv9ob+6kV/DBeaPNay3hgXiaFfzo+
RRtocXwt97NEHiL22kXDOshB2H+EWHmu8/ckp5dwIsx+dkUNDsugAQ58GF4zva6J
R87Tk7lQSiPixAVzlRzmpvs1uUOAQJp2H9Y50nAViqpZmAm71oYuezt41kEe6Hrr
AUYZ17Ll2vyWnDnhm9gajDvTV/dI84VRcN/FALOE5HFE+CntIEleSUsphDgIjFHk
H2ajG62tIhMLyfCxZnUCJXOj+ctMphX0IC++7ys/KC07wnoz7OV7pkdCtKgMUGDi
31LrtTtwnfyfvzjqOSv2ZRiuHeJkdVHH+6evlBCOvgaaTCyYMuKmdmA+r2QyIGdw
O66fFhuT0tFYpqoBX5ENuJcEyqOYWWQk0+roM/GrvAsycX0AML+xH6C83huAoBfi
F8dEHHAmX8ryWNbJtS58a6mQDqH3qKDmcCi4+PI9RI+p4SVjiTFWkBB/vm38syIu
vPvwRtiqxhQSZUourznXfJCOK6p73s1w0vEiQE9ZLWH5hAdaBq9uOHg5rp9lbc5k
UNGrpkCTSfRNqVOl93wK79hE1GQjzjvZqTy1MXXg9cZnpB7ADmdB4CKJ2lPCgmVI
52NK2tQN60mX3EW4i+sgdHC3wt7ftaBwlaU+Vy8J4j6yATQC6Im92g/FdNYqbOzI
IEqC/BNLG4XPMWv6PBzKYXBcL3oBMIbljQu/gajKwryTZFOQQrE9g17XMfRf4iGR
R0WWM0vyBNshTwJRWu/lKobNWFdAfsrvplQA9O/JhEHzJVZdZkuKX+AtIrKmWwAg
zZKt8Kn5UNw2LdBet2t20MxrkiuBzYOt01yQmXon2UoXd9jMAuspueugI0vKIa1b
6OdiTWi4mXN3UaHidELFN+q07gtsSQ/gwqGL7LeMn0B07PtmuXQZqpH9waJeGuD+
V7dZAZsegpuot++SHrguscNN/IxHjhnDMLJ84RV1kFwcRyUAE8Aod68pA9rqZO0A
7ZZL2EN+NQcxkhtJae5+v2PcouAaVfVYL52pTX0B6aXdlhtz/NPZQqybXi2kG8Dr
fF1MpXRrdL09yOrMXZgGBi/C0t8XE7u80Z43nHWo3QCHltuJFzOVOAYqiSHCRHVU
dqGXS/gRr4FVeEx1LuB8HNLwSlY5xD1yub25Tm64RhUmBUit1C962kxOFvwEcuIM
FICPXOuL+x79wclyMoZD2b3cA9lAII2LIWwJ0nPcoltJa6ILocQQvtqpBo/HCJ27
2hFNDpAJsp/NgDkafh/TqQsVqb2qLa4pEsoj60Rwgd0+UUBjwjnR2c/WvnsmfsM1
KpgGzOxjRJPxHMn//rhsZnaJ71xf68y0VyT5XHMvqN/m8RJ2WKdlDZBgzyGEIz5i
ztWtEhbaVFn+8I3KandAGJUu66+KQnoaJvm36bY4K3YCqbLYqfu3eBvaCmJhWmpY
1ojBZQ+0twS+h/q5nYsLSX1dOa+dQX6tNJH++UomgGGJrTFYmgCE3kvxwiTGKqAm
ZbdG0dfhduMvt4kDU4AQD5UeUdw96J7HMHrnlsQ8+pUq/SQ7ocnrQ8pEpurbK1KD
dBs+8GX6/N0sz7qC1AkU9sWxjvN15MICxmiZRwbi8vmQCSJoDifo/iOqft+LM8+t
TfOf32p85HeU8zACo60qHxqZkFcEbZTjjA4253cPm/j1qIOQHvq1vH/CyfO6g5HE
ZnTPn5ID3+5RFkAFfp9eqc5OmX+0rCS2JlGDIxrmo23/Fc5b8YoSYTH2YcM/gE5h
Ge++skf2u7ShAWhLfszNX7K4Y3qUWzfGGcLE7g1jdrbO7LIsEPrLgl29O1Am0SNA
mDBU3bfnIg980XqRN+Yi4B+2LNkAX3AtdsUnJX84WQvTw2kE3B4fhm3rdYFDjFUc
9q4zIsTAoMYGTI31VQciF3a88GXNZ4G/pDYsvVRokW090+ByfQs9HaK/TipW0DHk
QD1kq8rzkzRZq2Eat3vTRgfdtzoN5UhQRpiTk/ek5jeaiIF70Rch90ojXD6vIcK4
XWrvdJytDSO8Bwp0jASWJGlGmcd3jWhqvvFpsHX6mOmIGrwSDPMDHrILFt6u3XJh
5oGgtL6SNxbrvPcfcTwGr6hC/xih2Tt9X+bYnYZqRPIFs/kBH6vH4eiAt3ZxJ92L
83t83xp7TSdRqovQ7p8AzoatmLJRNP+H0qL5yUj+k7kWM0EuG7XXZbWEsyB/EbtG
VGXlrOlZ+z4icVptoFHhs/Ij1KmvNdr2whpVgGhv93IlJtqCgSEmeEZQ7HrJHE8Q
lkBIU0FFDRAB/YTLidAR4JPpQXcBNfiOOgR28S5VvRIsA+r9jXPdhmhbqG0Er4YM
/96xm/LKS4JhWS5AzpGpC/92AIxRQZPIMgaDr6lBdCCEJUEOenudUj/oCJJZb1Qb
usjekaz/ZcVb/diVOFGGFccCvimt+sKbmnAeRDYfyxApKFLLKFWf56K2YrHdEGdH
rRhxXnukoABXwNmXEVg8zdaffy3w67xLb9BJ+6EnkjX0LBQGn1KPrzV0AEN84sHT
rrSeTT6jlDECgHXhItGj3Avcn4ARGwNTDUC3bLjznWNpoLLJqBNcYw07XFiCWsOK
eWiJfl0T+dZkmW5PQRawofoXYdSpgZ/vNufuV231DIdqT4WxvfffXqB3/LsJi+wd
fbCZh5wWZEFWdLB5+1Cd+OkkdnqTSnUtzwSnkykBQk3TpxWMDszZbkfsc1xdtFZR
j8P2xn78JjFqnoAiLJfc/7IezAuscL/NpxU3uI2BP8GE5yNWDD5YBl/5n310TCzw
NCFaOu9izMmTW1gjNsAIHJkD4vEKlK+WtfUjUb78r2GzOU6QhOg0+7fMMRp1sejm
nSakb77ud09GDbnTP537LyFKkxdo3DBUheIR5/GDK8dahl3ko778GimzUclNOLmF
pdzg252Ud/ZhzkW6YAZlDBI8s+axrl5/swaeQjy6u7WJntUfv0MsyxuBT9zD0cWO
vVJfPTiicyLPhbzqxa6HskhIHQabk28Cd/NjE3E/tvZIngd9NjZDT+xjpHg+zzPi
jknL5omo+cvyNMwHa3SEWJti4en4NTAdP3+KTKIHzxbk6LfO42+a/cmCUFe3fxCO
2+Kaw4TpdfRYEDlf3PALGYfk2H9SSyqlEC3b5xzMz4qE9EoU5XJRW6+4Ku+c5mO4
jAo6UYIIqBubGdOyKZJWDvsV2vyQke5m/ovaeBaiWSy0R2geYb16AS+ufpbRGxSB
Fr3kZsc3A6xv6BlThjm4wyBWZ4665zwZvxdKvfwuZo2AC9l8ASi4BCrZEDgn/YMf
hsQ20er4NNihqPbbtKc4XUMEYxrnkPWSeYO6vNbU6iDwkC0Bag+4o7l7wFUYue/H
X3G0tHZ/RqZhxznYj5TzNsHiPGDlkNtYTQIm/qqZ7fxCfmntFeY3ohfCd4pDjTve
RqcU8L4bVHGcKgD+paUR7RBaXXKMERJqiB4FRF+6L0rCuMGDdDTty6EW23tfqGIQ
vazIoBQjjEiiG76Xmr6/3VoJw8r/Wccgo4NjP462paqXLBcotHdQz1TRcVk6C085
X+bBXjT1bwiztR6WImFAh7jSO2K9oSAIq9iGrGcz+AP8mbBMkLtc3EdxX1s+z6mf
dD4X5BGYphYYpIFrCgif0eXNru0v/7h74lyvSWIPVHtZWROw1wAdoivcpPvlGEZJ
Hi44PyRnkESXhNLMXRXgNlDeWGwZkapCK55muLSO1Jt063L3iP+ESSfcyFEU+Pc8
vCEZa9eT5V4o/5+Bv/tAPE6P7UM8IlsQecKzRejE9RKkrcEmZlg/keR7ofCPS18J
YeKlPiTl/513aHxjkOhM9kgigQGD9FXeCNC7AHWbDY335s7ytRHs7SVXmbKj0Edp
JHy2yQ2T3fdWRxylRxwuPLkVXmhqNo0Rh4bWOUlgX0QNTXDVEwyPmAz/tCUynuYa
E+e/dwD2f5X7jbtW3PWtjzUdZwhowqM5tu+8XuuBJlYXHjbhSWOTFmiZBlRa5nOg
mbfW4wKr2D4Vay6LGc5eWSxoy4ALFPs0uZRMPkQINFrSBpKvESAYnZw+X5TI7fsy
yyQ3t4EH1wKDXUgzR/3Kwh7DfKnUB6arail1f1gv3lb1yTXtbqIXFTnXMWSGI1xC
D9VUNU+FuGXz3UbKRFbBLy18jj2iK2Vr5gXSjPIOa1U4J7u7bzhheS70ACYS4kJO
LFuTnQ+qFcbcs1wUKJztYMWbW2fRyvccgjTl+db53cMON3wuNRPMwoqKzAhTGkOF
W7ApumRCaqZC/UF7vNPbVVPiLA3HzOK1R7dDz86GiUdf+9lbo+nMh3EFvuTNwooq
rewQ00HEtmIqKk036rx+cQnZH3RV97iqNR2gBZbLtpw4uuwgFWUP8IghXanQCT4L
w+mSOfefa6JUXep3JuCjz9f7CfbwHo93JxgubYl9DU1DlaeKNe+xYDifQvtPCnji
R/6lc+5uEO9YpyUVQ+/Ymr4Ukt4d5NbuP8eB9URbjliRNsHrvUjp/2wJUPvbkPo1
CRiMB6DzHPvI3SzgRbre2YDGG+vKqNrLgbl+Ml7/J6/TkFcMbkpyXn981vzSW4QF
ReoIMjka+XGm3U4QP19/J+8wy7BQ6IgPqAAJe/okLBrgRvVYBDTSKWZHG+73jKxc
dX5qjg8AoJeAmqxJvTTR0Fp+24m6krFOmjDEgKcSb2BbumY69pd6E1a7Q/EFenbN
ELov66L5QTAPG8FsAljlB1TybqiB0FFSP11aC7aI43rxiVl7G0tYfKAni/XfImp7
K68o93ZfsxbZS/cT0uNT6BN0lf7hJr5uN2H7jLk+1y6sRaQ/kL4DZoQ2DYL9S5Oi
1oW4WyP5Uon0lTXzdY2ROaA4pNEp3HQpj1ai19YErysqyeun74NXCBfRX0X3Qf04
qsLhiiApYkhcSOVpsn+I6ZeY0KKR0jA8tWS8UFT44yZ2NIWTCjahGM7+aZ4qK7eg
TdAs9G4GX2V+J5w+ut/4PP5cqS08tCN7fzmKUExXzAKuB8dBLN2Vqg2bv+wL0uDo
U7mWM3aHJm96VKEV6keZh0yoaK8/duLbtI1QmE+x3Hnc54VP7ZHsj7x54DkeOn8U
aQZt8LOCRN27Wh4gH9QsFfVt4bKhdYnQ5darQs6617Gx8VLf954HdbPeyZ19eeAA
uQg8yUCf9LqKxaGdF83A42fcIX2QHX/KF3hK5tZg+Hv495yLzvAaaVk7c1s5vqXt
6StHjhxar3MYPhOrB8U2g9k+OzS9wmd5RW0xbwo+hGbQg6+j6sg9QWV3EptdpOUF
svxM+/khRE0bYSLVqz0CDDwj1NZEA+kWw+My+gekt1YogoIzfbX7Ja9z04nK3m+w
yURMonfJX/ifj/SiyuRR5Yt4Rf+h1/tQPPLTjBx08Ejwds/K3LtYDmsKNF87/XyB
FYQHp6TfcL08StngpmQSbAOEyX1whr3SvrDdQECEznWxcdRf6mE3grCfiR9oizkT
4a4vuYdCSFJbLGD3vk8uWpWDcyFRQffNEdqpRH+ADsHFC5iHZpXcf8B1y2YBXllm
ar87OPxTZ+3uKmD4WjicQ+lhuF9fsglKJrIUXp9RE50Wc8i2PdEjr/WqOtjehA7Q
TjyHw/vH0HtZpmqtG97m8bnWEnyAXqQ/WVpg6xw1yAjcOg6FJ1q2PNcwwVH/TTtG
uCVlvCoqu+A2x+R1H1m74g7JtuFAhwBMBz/TWZfzkA+CTO1/St0DdKlaeCTbSd9m
jNPqPoe7CIB8CcS62QCGndcNwCnWpt50X/WoFHqKrQOQ/Rp5wU3tMV4saS70o4+q
SssYNwjMDCePwaI8a4Awpm5n7Ve2VF6e4qvFkmuFfl4SBoYQitib2WIy3EgraLqh
JU6/Kpgxu1m8VMXKehEbF710XIpjaHKLyZUxCJyXAx4byeYqBRbVDKbexI6f03Zf
gghRctrP/X8Cg4h5vEyNEc4k8llPSAoy0EaYCGpuSzsOEujvKUHMwGLHkiCb2jk4
eK4QCBAfp7INfll2nKFKLs/ACSA5Ik9ZWisWqbLTJiy7r/i40K97gZ9ILz1zq6Op
NuKKLUd5Jc4Iyx8K4UqcqQW122urUEXh8ttyvpPOKc83ecIMX7UzgVw1Jzr7ZeQT
9JiNyr3yC3pESTfGqsWanjbmiebrZcbovnXuEtbBcj5GHaXx1tUrJdFgwaa+O4NS
pVNZhfqug/Vlng++hLYX3imcoXNEtIgRbRajc2Gy/OA3DIej0oDgjgpRQlDN+cK4
ybXiszV/pZ/J+WvH7+cipWfsrBr8NZLGRsvP4Qo8YyvHmVtmimVBAA1t4liL3jo/
Lls66hUUZ8fkDnioE0kD2/zKwLCgkrSEo/JNFIuozFBPvjVSnausRKbvY9z4klQg
uNp0UoSs8YyqxZprFN5D5Hi0aYPHiAChfPkK7UKehGdLuF84usCM0DgPsmOPlmS1
9HVvvo3gsVzDLG6J/h1KxdPGSUOxEhjKlyRFMmUtmNeAEa3aJGmS5KGyLIS6JiX4
GkWrOAbymYmrOLHCwUGJWcFeRM3wdOcs9HK3G/rXx5WQ9DHYt3b86IIl6SbA5ESJ
r9R9+Vw1W1rH+LsvaU20qMRby5jv4G66M8ETHkSS6mAHaRgQFRuTcmX1a7CMUdwL
SuL5yJj4OM1YKuZ4+w/m3y6qv6Hl1iUvXKZKY7UHofriQFqaTqgMw6Yl0jYlSRWa
pgclGDKWPIG5HSocvLQcc6cV2MZxwclurYeo0iLZ4cQTlurK1CtapHGYbHsnRCWD
4AWcEuKn/dcQI6fm0BIAJvVm/chR9AKOMfb7APDl+Ed1ugaiROWss2cc8MS+oM48
UB4xkaoess/CeBCg4I1BJDl91elbWNM/4sxOpI0go+2LIWb8lV82aLqi1KICcSdL
S3uEO3VV8Jfr+8goe9xSyYLHbK809G5+51JGKV+yd575hENMymMp/JBsqvZlFjZf
RZHRgPGKkbDBwtWhh9Ksp7jfHJXiW9ByU/lbml4gLdCswU4uq6u3C1If/EiRHs4O
M4GzmPFi0a1PYxtsFFlTtKE4yMx6LInS+G/WSFBgX1+5QOXcZYaohp2XcVph02sh
mDVFlwVSsKe1j0dkQSqRx1L7Gko8q3SJmJX4hxjPmqY039uYlxiRGMAgQCAd7n08
Me85xVr9KUJWs1B030m1X1djCk+LexI44hO2NXVirsNamXbroiQUPkafOIJt6M32
Dmhg67QFhy7M62X/GKt1G/l0PfISvhhJVoRyltYPeZ9eNDj+/UbPioyqdeEsBNfh
4Hq7TsUm6WesiPPW/FYycWdEgQRzBKPYgHQnCteawxhbxJqSTIdwMb3D50yZLjRH
dd3r4InM0FSD4PA8RDDqy1uWOAgGX73jBBWkWDHvba5pMMHqg9Bv7W2+vuJnU4TW
svAFM5izs9KUfoOfuRHrQDDP8KgpVNVEtmaxvrJmE/jrHiNWzIFngh+CxZokHjMv
yh9KYJVXHiOtCbNwrTdtVMxwd+imPtsMVtXEbmB5+5ikjMJgzCBSK0hNufN3xC+A
Exs2bmn+zjpXib/u/DfwAzFYwqjSSps5lPouqi8uoH31aqVqfWvAyPg53PxLd0PC
i67BJn8BIH3B291fO9xWEWY44bE7GNjZVYAmrEeVCvAoKs+NMVuYL0vH5NG+5/vg
uLhroTbL40fUdHXucHQU3f7c7NZnp/upnGCXz0jqFjN6wrUxkbQ/Gekszl7x7XZs
/aS/mekap0FT4Q0tyHnE3fey2nNW5z49FHB8/9OVfw6tLAUJUiqB/EU1FqZ7DEPB
CnjaNzMKH/5MDY4GXVEmtMtGO5kakIuQWjMav3Q4kKiR704gUn/lbezZ6S0odsxi
lzDM/82bt7w7pJ3HmK9wPLbcfICXrDxWbaFtcfrHOvDVESJr2KaK9/fDT+k7WPt3
AlZsCmkEIQC1WwzYHrZKe7xW0Uktq2QKfLlgK9p+eHYtGhz9EuH76uNxiKpcdvVU
6NUGZkYXwgqnwfwiIHXgG70q2+L/WLtmHVXkXz7DV3q2GLtjvwnDDPjRkBwvOX93
cUhY6Hrawtcpcf4uMB1D1BwZiblrdD3VhO//6DnlNlRNXglmWF006usSNDVpmNi7
/WPGYJ2vdIneyNuSkTxpHukq5Xrs5Cq9pOanBv49MShi0ZERcDHAfI6TJ/zQvAB/
6S1lyK04IMEFFY2mqpm1B0S/z2HyoLLahHLtlGskr++fY3Mri3E2+nmBxpUyefQH
FPv52cWhuujoI6b2UuqUdP/j3T2uxHaPOTn7qj8FXtU3+GFE/Mgi3x/BPQP2QNI4
IxCFkwtd3HvPXnScCyf1+5NnSozH0jqjjFd3NHZ+XYfB8jOAcN0fcc0Ir1Ytz3GS
UiFF4xnsYAqiTNnDCVMaTCbYhj7e3KjmU4T28qOkBwDvrJwYbngCW1GJnw2FaqWB
F/7CtapQNujTofWjwpQMpiZsTcz5xrJDINrm1S9q6x+cqOSwk/j7VWW5hHRYWf1F
fV83KmNevqoHDjCO4ngnAftnsdhHXeNviY9qytLT47G+D4d04riP9WTuLxpvFG7C
Hz+z+qJms3RWazbQ1zMuzx1jeryyeZsaDNh3U8vRObDFLc9XmA2uWYm4T/yMRedr
hkgle6dA3YKz7Xc+7kOjXjvOhRJK1vlIAw67zQys71+KvoY4ZWieE8usb1PINqwP
66SZh5WlSw+7ovoMgcYPcjYJZ8J+EPbLM1/WcqKbPvORelJCXoadKpBj9ox26cGz
H/+oZ6AI/1T9sCxhbSYAvReq7XbXtp3GjJwxz8F8b2kNf7eHYNRdbEAQ470Se1YB
KxD9gn5v/4dNNa4GT4rTuJT1m15bbZa7vpmu32q65LP4sx68L/ZS29sMzrqpYHy5
P0gjfSGeKijz+7RdMT+oQ/uoS3FIo6FzMjnxOcgv9UyD+fekQl03qS9p9MMjoAbp
r5UtAoEYWipqQ/BYLVkuceEhZ4QuzIwff9qt5UACBiFKr721NmhSVAayealBBCKE
M/FPK8/izm1pE7bjhZeZulkvK3HjZKXhY9ORiLc3uPQq1EAnIA2E4jNhVTOAYf6u
ntA7u2OLyOpSsWrRTuXsAl+tl1ijwQSxep0qKRnJUA8ovWGFjJK8/iDYtRrgmEtd
ORjwHZHPUxCk6DmzweKqsJQ4D8KrSh/I/b6LrR2xK/ZsYDz9gUfqrhDS9HMknnLe
JGFSKYkSRUj8Hrqv4oW+OXXRRmb4svR6jREwLqBhsRjPWxrxUgbdfCb4DSego0pJ
Hb5Jv4Iuh8wwSeDQqsqZ7JSCubdDD7FUoChF48Q2FrAx9VRbeDi6/+Ep8zNlp2Yr
HOk4sYK8zZRi5Uw1azCuske/+BeGS7yIEU2x5bcJ5/gk/daHiOp6hXw1BTfKnPww
fMbhOb0ZAMGxssraM2s3MQmFq5WVoXyxIqY7g7hqrUH236DZN7w17i/CVhzt7ibJ
1xgJ6HBEnIyEQnvAzfMc2zMm6/9QcMsjSIjGgMeCNzHf02GzEApNhCbAmW6DZnip
7Gncdn3KEDM76baADYJj3eseUqZICwUrn9VtSW4+BHmZeSeI4KaQ1eTVCFaQsy6h
qJ6dWeHl1ndgWRYSACcZeMAhZrBITaftKfboicFfOFUMPAAhPJcfeIgI7L/BysBe
IkP/JurRanKJRN1lg7XA/NiWq1ogYxKF62BMs6qW859Sb1lHbb+TMhlNvK+y1tQG
yvqhCAhIC+VIAKMb1Id19ZHQvNdZDttWq0N/DVyW6HWCdYqQeasdbJT5Wg2lxIkZ
PA+bOtt75MOq9oZeUsiJxUIAQnNhaSXPfL24mr4Dtyt+hyxS2Gg64t/r6Z4j3pVN
wXVW3Sv6u8AcmPRNxwZbM/iH8lIORPwzlKWw0jFDvLZBy4siYSanIVzMYUgtiogB
lVEzgmOO0FdKzsMh9L8mmAwduMIgn1dgoTRSEq0ztGJqHYO2wJZE0FA6qK9TIgLD
i8BEUCAhJnSeWgr1PhBtTaJfsdVR2tHkiPxrFTX7oLEwd+HlM+CFIpvIYxzBB6na
CCdbJm68r05dX9IxbnAnlLa764y+viZSxUAW4BBkiq00tuAeVXOELt3zCojfR4Yy
0vNO2tj7RgsHCZhYn3jLmkso+Ans4YgYZMuETlhavQ4NrGO1sR6VUcuo1M/byqhz
ZwY4PRDyCky+jsI9PkubNY/YfKo7NOz6RRvVX0ebwiAcOWywxFGtxxdM+zh2A2c9
SwUTYyBXDDgaJtnccQ99P6/PIu3YcFJ+cv3+MyNpAn06w1QUSWyKHW2VPO4gjTz1
goIbyhNAwy3yKvPeLHdQI2IiHqexYlvl8MeDWKEraivucVOBYurcSjxRbn3bqpp3
K2pX4kxWAE1cyYHHXC6z9nWrPPsQMtbfKz3xXSfUMN4E3xhdamrbtINmKsuApasc
9gOV/6ioHgfrc8Mu/klHb9G16I3mndptzlCTp51GU1cqTrU5lAxAttJ7m0BjjhDC
VmbDfsEuY5ofKv/84Off3SlNNOTXBtlnzGXrmCNYJy8THcJ3BgSff5SXTU7N5PGV
jHvzMQppqy44i29+GQ4GzQGyRIyvmWSjkLLF14BqW0payuBwZVKkyGELBkUHWT+Z
v31MGfF7zoQmKJMsvNgYDjTOWolUcoB2rrmZW5Nei4aiK6mmqpRhdR9XIwb2hLqF
SuOfByVwHbFOrW/sslU4QG1j2JP4GSwoirKs1mYwjEOPAp+IAhFg1oTBkdw6LVra
ymiVGpcSyj/voQruLWHVkJwhqePMQEpxhLelddodqz/feWXDz2MYCP/PauqbVulr
eccgQPxvE5VMRArlnzFIobl0eKLE726tUtgZr9jSN1InqEnJokAkbkdYqVfIJVHM
t7CELd/CaQD4r2BQ7+wzfk0E1Zz7gRhmPmYh7jwsAKGZQWGmMNUxSRfCFRmB6p7I
J0958WIAsMxCOy7VPXM4OADyRAnnJQQEgg49IZ7CFoE2eIqN+wtKAOF3jDyQOAZX
pcmYJdb9fMre0vDq+Jr4eruaiRZ4QJvk+tonqad9HokyOrKEdytJZsrUlWgNjetQ
gPQb5abIOm6NGWGoWZqJGzeEb+gy8R8tQI2gnTIUfigwlERMIqNgfsEH02XefOgR
u5iWJA7DQELhhdwcqrTjOFllHfbiAy/By6kJYaUaDraHT71c2rjPpVjKw9cL75t3
lqp/QqA3Uc33ngP31ck39TxRruXUbgJmPua6r2koQewBXCP1QaPJBvlXVl+moQfn
18zWwN7xK+UIXG93dAQ7o30d0Kyxs1nCGGMEwQDRiUPQMhimdVlHd6Bz9WNZfTBK
FLCHXhY0FVLVZj2wagsyQsb/TvTvzPuEcUQhtUBqvFMwnACwrLuajM0vyZNkAfkP
213OVbxdWuFKq/aZzPdmK7ys95HG1GuMmSWhVEsGfNupnvUF5K2MaE9NhnxXEes8
Y+p0JSLZGXCl2JvRNELBveUCa+wuJBs+CQcnmOcSCYZfW9ce5W6WUzpD7AMgQask
Oki/Sm39ZTqJ6xENlPzw1FHuzjv8TmCd2XXDNuVq/QiV6jxXE6c5yLs2wCg1bZBA
lEHf+ddhMaOcybSnBcSgO9ZoG40s2ieBMbi4ajkXoD+zT2oj7sO+mh2jtyJCAoiY
ri+oQAUrWZhWjSHxT/x9OpkvqG3ACVQC8cahAvUIlwWedx7Fwr73rfXqkLLYSVrW
FZwpR5cvzXWWBe+UFLLYY+AoSA+HOuMv8G5L+0wxfIuDYV39ZBNB0p5GjiTT50Cs
o4obCGIFhblJeYPMAD1y1DK433zaLCKoC/sv4C4MaS2y0JczHnHLXNHIKCaEbxcD
Yb3C37Rr4Cn6nd4bF71IPas5bWovfKigAE5rxEpqm18LXJXGvwQcEVCgUl5cugCQ
0q0f4rn5jfa2hnJBt8vLXf7bj+Mz0A2mhFnPZJ1HMIfwj0qXnbke+x16cMkbdDNn
x/CSrOrqXFCo3BVBfnhhcaNcjApP2jJijed4y1kl9GRxQbCEYwvWl6D7AtgTEf8j
BLsoDK1Sv0V5XXV0dHX4VrLSb/BPHuIR2SgnRR2RPMvgrWs6WnJA3t/FQrvgZJ9l
7E0D0q6xPs+74MSgZDPVUqxBg7bNBcpqB0NHNhtsF//Xf4MwGdJIq2xRM0FjjzQ3
UT4x3XEZTmWBG850Olbf2CYjZnSlKFTigQlNdlsFmttOpjk0REzaBbH21GNJv/3s
ipr1jV42taPPh31KicRciO7yuObfDpUzqssOW2lcea/XyR3vU3ULZ069RIKSARgU
5bFrPABgtgdHpbesvX/tNuY2yfyrpBDpHVQB/THdRyzlodQ4xeSRDfTmA3aFUBxJ
I4V4GDnD7ZmbJ/h/dY5XxZpWTpfO5dyFErmHFl78WLU8E4sLNBlB+AIqPjcydyfU
52MblPv873lh/6tg9MciwhM1CrtBE2qtDGHgo9Kdt19CdFT3RjhQ2gBUrPStNYgk
Mbnv55vP4BIw8id2N+MDMxru3sO7eTqqzzCP/HYk2UUUOuFqJWejBaxVCeM73IqK
VrApNyemH4HuI9e1t/wvZ2b5LY55FX431x+yAQY+ZCSfvZh+KLw3yhpd0M34Al//
LC1oeYmWEL1a+nFvoBYMbq8g229QVWRV6wu1gvvW2zLQT2qSiM/pimrDMTs/BnRq
VdJHc7KA+Wsakm1t9RGOwXas82ViZ4QA5nMd3UKc86oJWM402ukIdwsY4B5YJJjL
rmu2RXFqRDQ1S0bvD2enevhLRZnk30ISW7FbdlZqASP/vFkQCzXYv2nAfuAE6l5V
agdS3xb1lCin5nXhEcpJNMWEWC2LqcVRQBZ6OGkxw3z4587JPAGh97CKUvG4HecQ
YReRZpyM5sPJof7CQvccRnnVCX0OdBJp1V2jzFahv17FY4t4LW61ZTds8JVfHMxD
Ac6IEl5q7J2RpUJnT3+5qwGMsTAY2cwLzyXVnF3WPeBgKG1HmmTOiectqFxE8w1S
E9LglLkoTcVAWUk98oqKMkRzathO7BE3Q/Epfs6T7ndicpMrJLIPL9AhsiAXVkeo
WwLsPQyPSZRyWN/Itp65OIcNpyJzl3ec1Ij+wTuEgSEuvYarNqsoyOHABHKdPH1c
kOAga1E8X4QuaDH/XQmrofxTGL/xWBS3kSWwa+vbZCDnyWaeOZoGPTXiEReJKr88
pz5t6UQKO8t8cWNtyrmG+9P0GhWIyCe50G0hspfu94YOrxvNZONLPETXKtOjZqYL
uT0wBpr8RrzsP0fo3cB3tss577dyCKfVb/IAmjpuENMU5gfsQEgAUyANZYLe6VEj
K90SuOMKc+G2c+qQ66JXHtZ+CZAGY+xbiDhfnvURChsqBN7GeS/mMpuzCMl72HR7
uoaycto2joqzcau78sXdzo7QK7myBWgrC6uPG+kUoYciikyj8gvBnExaH6ahpnkx
f/dxUqYyMEKZQenDoFcGnCC7LsTpaBKB2jmLGoRnm1xqEM7tVj2UilzIivzYTaiS
wlkifXXGCTE/P6V/bayraJTRGSm+q5lj0H9AxzXIOrtzjUo6RyS/G/LrdE5zCPfZ
yAOm4pKZWsgMECvXyoCPz8dUqgPl5ZwdPDlQ6f6nUomN9R6duSfSxMOnOf75X/yZ
ZywYU/2RFQK6263keyLqM8DTifAEgQC6LCIZdjCoFg89A3zOBBUwKGtG7C2mX5uA
Gy+r8GoTwio7zc670eBE/ydLapZgppqVWtxo3aD2mvaVHYGIA9QqGmQ9SqeTGo7I
Tb6EUCyPx3vPE4G6yHRwNCUQJekO1KuNClfT/mYTeWaLlxaxFf8Ezkvh6HCby49S
AE4Dr15sjiOUkXc6mDCT9eoYVO/XJnwzPYIEqF6DyJiTNCkgEIMcixTujVdW8I2J
ih/fhYfvTN882q7EgLt89Vivrb91P0/v8RgFvPme0FtTRTm5jiqgVHYoWeMcRoZ9
TpsxWh7F/N5ebV/PawIniBnH8H/uMKUc2vBA4gWx94VghwSDxZrSqEPUwnO6HEuN
Tncjq1HBgNumAVqL3naWFeTI6mvNMfjKWfGT07VI66Qj3kAq6rV84uegYhZoLWH9
OyxgBK6zcaHkYIyxa8SMg49lzeLcrvD0ZBcEYsYzFC+B0DuxPYHo52n5+8hYvIlJ
DsKS4cqClZMLNTMrZXTIhSoFu141/aaW+lzW5y+ABZAGEyMl5XVRPh9qgoQSip8K
pRCy9jaggJLdnlGA+YtjY7pF9ASkKsYU03hhEAXMtTy32bmjeIdIhOu7/WAbyH09
PjmVdZ5sba7Jt0DtRmDMBS/rBQGccdELzu3E3KRoF9+efMivrd4KZjeJQmSStYKP
IPilPuxHifeVWpqSsq387SUDbl+1XeDdUSvXIG3ZwIW1TC/ywtWlv4ee+Zww9ekc
INxbX7Yjhxeg5sAkgpqPOCCtL8Q7e+XY9Jfhp14pPWhkq8LkaF6i4e4WeBPukOhf
ib5jRKG83EtNUbv9ZzAkfM/fxr3OMmfI6n4F9JnpqJHTaVT2ZYGNe3Vh/hzVKZFr
Q8HlBIr1eUY83VZcgvfAz5Dj9h8qO20lNFblRjvIDJ61f9HLMa6iGJtm0V4KItLZ
pUnmW/bVeuS4nmdHejf8T4rrEI4qMZMy7LPPOgjfHOO9AVscS6ZYu1ZL8SZlUkfp
GjpN3Q+qyAMReh0PtJoFKj6yB/tLmW89rmNRThnLljJvVNmw0zy4UcCh2RzQxdgj
86fyaAjiZ8SABv2r3Zua/+DGwdV8d1y7PUnFv3xrVAG9kZVvoCGlJ25HCN+zHlwx
o4vnNwH9xFDfNP690QooaRGVKCqTQycvt+yyuGn7ajBgNWNXsEzxJFjClrHDp9kR
B42VOH0NdJSFA1IevdNG2get32LRF/iKgnL+xX4LOzL0+jpsPx/bl+FqgsqcWMxY
IVtyQ4Gk+Yu3lRMNsdHfqvr0otEvYvvGw+F13whcCvAWcogfW78s1EAnglljaxe8
ebHyXbpzEz2ESFDfy5plBkGC7eJhlNnZqwfDtnEVuvjCV9Go9ZT5f8oG9uwAmOGC
BHVcajVtKn7YNdYoURYb4W9+K/vle4MLKX43Sp5iKkVg8Krp+jhWE9u41WEk7f7H
a/bV66cT56cQgywuCkxfSP7q/kLv9bYrESF5MB5XqEtZ/AjkYbirZRblhk5Ui4Ui
gbZWSEG5AeezgsomudH+gi0t5/BJZ24Nfmk/Xm9oSNI9e+GLaM+6lDeKf+Xdw//z
h1+4Smyq/h6x4wVDp2FRKw/J+hzbWCQznZ9149brPt3zlKZ6tBU2ZcPJHCuGfkho
ml/9Om2hp5mcaxO1yHSgnxLpBGMKc2mEXnz8PJRQuex9ordXPZaOGEFEdwTzz35j
UyNcUR/SoxEzJCptdrT0I15bdmyNwPgwTiPU6SjEfGLLOcCK/Ujxhe/VIx9lZuoE
aDqVmoboAAxXCdWqS7tXoAnzmBmuxU+lUtsSH1CHxs1n83Wv7aAzV5FZlv3D3U67
PpIW+3q/mVdnTtEbf/JmqCr7C3wXfAt8vjE/5Q6o6pa6O5MrZsNZiGICf5hPuygq
yq30A/2ivvwCGNSQDz0RADpYMPQRWgbkzT5mdx6i9Asg/9uaI2ZOQEfKBLgIaN2M
zSGKzYpws1LBzAPXv6dX+ixY9w6n6Y9zLTqhc8xSuoDSMTaDytR8rZSlmKlDtUCt
T0qQA86Npn5tuYqDC8DBEpnTrucB3nfxzUk/sQNtqPTeK1DWSnWe1yZkXCwTLLSw
0mSQ+FFxM8WUxZCzbGYLA1cc73lZL3mkyBvxSe5G6nEe3eUPl8jSQ4VlxiwP5q4r
nJST3Ygb0+g3NMUHUluOC6RX5CQqEhibx0rfRKLhMSGwDfDxJYmzzgralIhmRr5k
r+6UDP6+oZScp1e1t2k8528gxcTyXvEoU3hXCkizpAnjSXAjWbgUYW/tilWyLSYU
oBWSPEuanrAw+nyhdGiLduZgsRi8t5ZBdtBX1R4LZvIhzbaWOw1g1dJo7SPOehjz
iWYRrLBuFRXCJcyou/vA2v/2ADndmbeLwvjbI98L+s8sMnEnqBve4L8sSckYF3zi
+ONS6a2ieMn3lxfLrPggVyUXNnwBkCxuY9y03QNGxkYEtKkRn6opZrpiaVRmosyJ
D7wzU6KxY7VBSSBwLqh0pympQylixa/gK2+5GE2Dfp4ilBmaQ4ZTSNkxvuDij3T1
1sGFzACs56yJr30FObOLRaOe6TwjkiLEhoEYOMleWFQQScECQJPwGcAv7FObY0o3
oUyLsO57W5kKrOszodf8+1TRoKOsK8EpjBdFRxHbRRYbuhMz9JM2HynuF28RWQ2V
q4Al7Y/Xi/uAaeYj5X1XZASP/a9NJE80thBT912KBfJh+4mzK1pF8g9gcTzZpXZM
/aCgNeqnQkTkIShpUdabnoo24RBOHej46FsKnGW8uEVFVbHU4MqmEbLfB//+z1A9
V0luSvmgNZA8iM4nrS8u52D5qrIZ5wIuuHP/GZAJ63QEhw4emFM55lBC8ac4w+qO
SRSkulj7Dz9/Lw/kJF5Ny7M9VX+J+XbfxErTrLw38sds2PL2vMRJU5NxRe+PmqdY
TJjk1GTO1oYp2nZeukY4Blx2+zaR9GG4VyWjSV88IZZyVX4rvC98TMPqBS9g0C7B
4ndf+V07169twKvg2LRZu22SafIwSkVVNnHdHms83syJbB3EEzpXU1o9P53i0t1b
EcOWkd1zvWHlFbQotZWQOTUX0WEg7bRvkpblhh/Sd/CovvqwldgTIZAEUIhTu+N9
OoaMqprNJgklN8UVjx2CeFfEAjOlIQd4YPB+X7I4iLeUzE0BrN1JhnzjOgT5ma6S
VHEzmz5hzVmFY39CvdF0TEOk0+jJ9BILsw1DE/3qzxgLHazoiL7TjnMw9/FrnlfL
T/FzcYaR0JLHZ4qs/FwyTHQKSToakWq8P7uR75a8A9L/W3gRYpPredgCHWj3U+OY
J8V59w7A7OZcMEqTYpZ9CiBKyL2F10UtQQfKECTvElYEwKW0yaD+shYho27Z0PCp
ZkGHsuhAHZIt6x4cvKYhpZFvzzPHM9weKKt8tC/nRljfd8rBHmxTb3zWpN46twLT
KNkXU1Vh+1cmUTk2eV9zQFRrW/hytk2SNmcesCVHDU1/2HABiuK8zIukEzBfOP/A
3MHZZZjivJQqIOhzpoGBR2Jlwd0tkjn6sJqWO61fQ0ZFVua7l816zwc3bC46hRm0
Zqfw0U2uskrD12LKlLBtFRH5dTSYEfqdcH1qS2DjroQ1tjswnDwSlgVgZxse+lmc
Eg46DgExzmB0GxkpKeaMTb9PmP9In9UbggnIXrdgCBW9XdUa7wyg5m4+gfXL+iqG
NyETXsP+KyWNw7nSDNKZWnoJK/7e8mEgKbxmqkMeAYACUpTOswKzokeqwdvwzvwh
XtcctBdLye/Mj3baoE32fXSFtXk/EoO4dH8zytT6DLlZJkyNuS3sB+TCb3LN1HQF
GAELJxo9IoiU9Z/Mgf8oH2/bHPlsBAhmgLDpJzAJTyU5RGp7Lk+XLZLoLIpPn/Y4
nR2umzk4DraqryY8hkeLpDl4YrWUgfZeXBUZxvAPSwy81GzuBCSDKkV5CmoBz3aS
IwzJ2YAZm9kVAcGDKCoXfj61pGHeFg/6E+UMqQZlobRq1GsJp+cuW6d3aaFma0SJ
JP0IM25Blztx5VpARXN8g3+CdooNhr2LbpuXck1Ti2SctY2KHNnfoRLQna04B5sH
nSm4OMiR+F5RJlRJltyRJKZQDNlVO0ZAg+zC1aifyf2FzCx8U9o3JnjESqlgg8Cb
qPabUT5u06o6j4cl9VMTyLnV9Ry/vHh8H57U8UltTzKl7cAzkj1Osv54MfnRZFr2
h7DedCi8a0YeoxWS90+yXKB9p2I2+sz+VD2z51E3PA/nAQMEdyPuKvqU34ZG5yhI
ZnRUv4gLUCLZK4DNg48yn6lUcuBAAwPbjvaVmiobuZwLAD+a0AwagLK0Llb9+vad
swslqkdHcw88mhpLMiZQFI3uAyMoUhMQe+C3HPKaKaL5t0rfkZXmWmJjHwNq6bMb
441kXeUV7kAKMAuijEE7UymGJUfbGPlZiRexguN3j4v3WEfzqENGTvMvCv+P+UkQ
6m18qql3wucF4nq/txbQPV75+r4spiWQOn9r3LLMOq8bjTzHdcqMXlThpdjIqHgb
Y0Q1xdDtauSD2dzkRT0r1FFYaegdgwmMhpnox3g969rGL1wBp8RAmRJQCpdIQ6ne
WVGx/bYO8YZhLQbKNm96GQA6RXWRg5prGKlvz3bPuV96Tq3z0AnEaDrV95MBCk6e
XgJPlDSZbV30VKDhO1GXCGTvfF1N46ptABd2oeg3GRdErtQfr0M3Mjby/p7zNEdM
Q/uNDxTEc47rj5QViUZLs+jtHkVpCXT9T5sYdKwK3HD5MmhAsTU6Y4t72SsHM/me
M3aX1UXCDMDUKZdWeAwaNkLa02GZQsQe2cc5QxgKcA95jMkxTTM0eJJI4Ttz+jgR
GYZUjUaJIC6jBaU2dNPWgB4CJV5ggma97GnuBnE1eWidxtcXpEu/vzZ+dxf4cUQE
v4z4tzbVFeqFn5WLwBzQ0mUFRce1Rxm/PJmBhbjxj0Pj45HS5L+Evmnk7gwocF4m
pSHAqkmnda+5WDFIKbXnLDeJCDKlHrF9A7Dxvxxs8tF/4Gu85cM4oMo5FvKjo/3o
uMr92i2n5gG1Q+9swT4T4Inevb8A8vKLUkYwqOxsC/omfqSbNRpJG3EkXA0XoHUJ
hSznTvnPIsrPXZnGNVfrtyfnlv1e1C9LzrVXT8g03T9PDnV6BYZGau0uyEaupymf
l0/AG9Z6pKlldfqWhGaIGqUMyrxcvIN+6f6sAWzwXLKa0PsvNdciIB03TZx1x1e/
Kdj9+4rcJe2AGGJdbgNXYgTXd2ndcm3cMQzefXklz2Xs1fU+N5atHB+JFrKS0qKk
ZIamXHqWuMmgpmZms+SM8eNt0jiEslmNFmeZrnwnFkGeuEV3Gj09YnzOVDWFLAUF
pXRtT6gaWBKydiHl6sd58TF8xT4PxdBcCamIjlNvhl5ir7bol2gaFMgCKWGxnvj8
AilK/S4NXNRcIaeyWkR2FyxaJ93VR51M+//8SMrRR2UVJpOBP/goBRazS2D/UrVn
Se/gKhbk56PnP+o8IkTq+NJH2qzpRsMfh5hOkzCHIjlKBYGwtuaCXuSS4C/Xl2CX
gdSF0PjsggiZKomqtBmZhgcqzkflTF1GBXW1nL6hSyai52O11WjHK7yUOBbKa4jh
Pu1thM5kUz6yUCEhE4WGn5iiPS69r4XEpSWZsg6fTvVc8/TZLhnI9MNiczpEBdv6
BtRTic/C/1VYfv72Yetn5u65XFeW5455NXUro99Rxa/e2zK/jv4yN6gE7CAILWx3
P08QkzxGWcTdSow+F+IuytPzjie+/lcyLe3/V7DULpnHwLpyx5aTeHo/SgZLqtVN
zjI3jpj6P/OhiR7x1PIC61cWfa/jsDJnIhiHn96lmjRfzv49D3wAHCg2J+DhbUkI
VryHd+hDu6fnSNF6bPgZgVNJoP0Dqxx4CgdHXEITExCDmT3CsHts0EYNVuD53VLB
3Vp2Pmvgw9UBMzwSTU2CSrE3/kPRMU+WLKPI1eNxl8g00oBcbGwBeABDbcQUyuUE
jzY6DM+L38SFGy8C+HAEyGXZ1CWuFGO2BjgvydfuobymiGmRP/iBVXFOLdbpInGt
GvIdpPfFVGdBbzPe6xFtwxmgRXkDKwjDpbqaA15HRUGufiT8m7ZlJsYuj+OIL2pA
jPBQERyiETyZLAKqtckweokgHVwwq1QX2mmfFZyKA5ua82sKzC/lEJK8cTwqDBIr
s7a4Pu2EeESHvSftp7Lb06PxNUN3Wl9IujEuShKLWjWgF+M3TbKmv0RPLnGw+myr
olxorHQ3ZsHIFd6NQoplb6VTyG62g8MAiDYPbTHbtRNevykmJN4F9rKS5SQoxeOw
JCdIdSWjb31zR0WQyJmHpkqPx395BCA8ehLGLUgGhvHKEBfABk0er+g82ed72F6q
jljywoOLseh4vvhh/3gTe3GKs3nRvCBkfMtn/r/y66eRPGGZ4nEccadWn3Wcoxsn
u+KwqVJKss06LtUG3icEjKQEWFS4AIztQJN7jxuGTOs0J5hzal3oK8O3lAMOnFZ9
u/iqkMBFuDALAtl7C7OfCa3pD+adKZ941ZzE2BRsTswkxiHN8MGz3sYBeu+QG1km
CPM/7hASpTM7vswj8bILbwMp/0OcLm/mbCGaLpiSTq/unb2yqe/eihMh7wp9Agku
902RJWCJ6PZmp0VJ7etkUJtV44aVdO9brYKGE3AmHELay2Fm2TlpmBhTuc6g7/kt
/aPJnG/WJm33YnlcQPuLWMo4v7OS2ZaUscTlj5+Wo3ZtqgXSg4W4mUe0Nwmnj3Fa
Te03ewJScJK27NyBbvm6TOZCaReucRNe5nTXpXbaY/weWbru22IIWlyOgy6BoLtY
1hJ+leuqHGLLYmPyM3A+/wlo0bzjgHImRfZ4mOh0pxmkcZ4+4rQ8u58x0cWuqaxy
FbZoKbLD4BkjJ1eqo1pc5sCw/wrrN8PWRaz9Ydr4qjuLZsvsxHUZ+GGOQpX/+L1o
dLh//OREGHl/0Rw3RMAgW3LGKQeLJH+TYkmP0E2Yh3K4tFI1/9JBgICWifR+50ae
IZ7qYcdJy01NUmlP5OrVLwylJip61Z0YbhTMBsMtndCNFr71kqGmhKV12HlN5Rth
CRqekSkyCUFwRtyLNgh7KYBRe7Szb44LOH3yZxX1qJk2azGRRauhEMdp88Ztwiol
tNLS6/CoHTA6B4JpfLBvGiPXfSSxmG7m/ZrPdmTDpZimRzxEHVmkRvQXCA4ZkPre
20zEe2Yf8YNKhzH/gDjDQxH6lk/3IPfPS8xgW8dVn9v9IiZEnMLHfo4CuGkc3L/N
JhqMZdGyGy4JZXoBDF49g2UI6aeij3XufJFIrCy3b9qhvMY4tOBYmbh+h+CUxfek
X4vnzo1ouqFdwy8ntXg9k+QwZBrv2UPEdIVVhvpUwFsYLaHM58+huVAj9xC6BJ35
TmY4EWWiIwwyk5EuZFOFfjMd7IgR/XDxofYsPumur8rI9obpDLYMNgjNvzkwQPDo
tyMX9Ho1SsI8EF1oXNTKMGBzk/PSwvKjcFlssuOVboVV1K5DXKMaMkWyht81TV1r
8KXcsxHYW2R2oy2N2GOiK0ke1osz7K1Bo4I8V1KIVlgZvVx/TPlNi14oxevq1fuh
vOtyA/Idrs2UHac1e3NOlndARJXF4GKKCdIwp87c5ZYgFjb2NO0dGmf9no/l8UQv
dsk69EH9IQ2B+vkKm3qCRjUABOocGBITuv9aYAKbYenMVeGzvuzdS/HQrvbb28wF
sBxWJdUrPTqiGrWxE9XB9ZBdyI+TvUUgUkzDgOZk+GrHc4kFct778U7etyghBSqt
5IiYP89sXUicyndNhfe/v1M5BG4Hj23h7m6n0bvalyBwKpKknliIR50+iYxcbxcK
7oVRgg5fz5TRPLGduJgThIdis5bVU/A+n//Nv0JFAAdMvgonoDBdCCZDh8uc8ePL
8Uu5S8tZNnbcktPC0ul2kzXAANmDl/Oouep/f1ourN426qHy0DiW1forwVt3khHw
vmgxLnhIWl5f2aJrsnl9EExqA4BfPPTokaMD9FkMMzGb+ZXNdutEm2fYz6j5BMm3
MYLxg5fjJGFsZdPuiZ7Zvmr2AbkdAWiVadKg4KNgP7UU7WxfrmzEfrp2CTA65aev
fwP139o4llLOm/CJ+eEW6/qae17gAuzYBJzYaXnn9KwPoWjFltHK38PwCxc26cDX
Fb4ADwpsWN1xwo4fc9UtXMGAHWah5blt76z0xA3bmoppEpTcnMids/EcGj5B3nVa
ddF8x5GQIE0aV7fpA54g6FokC7c5mt4PllGk4ayFckrMtT48w/O5YsgM5y71LLVd
k8gPG8pYmUfmSY/pXrsur5RybuW5Vkxi+syuRsVD+gsZ17I8zYU1/dLqFTYxc47r
2T4qluTHyUeWZiHzbiWz+L1e4tO4TANPxx0BCfmTAWhe+TTWhMtQkSXcKUXsKhT1
nHA8oq+cwYqgIz19m7LZu0WYUq0K5RQhnc0qoUTUYs0czZUOJRw/iCV8cjJCBU+9
NZ9D0YVDUW5M4gtbmfDcSxXwGsM2+M7jWPJ3J9BkJF9AibUlaZH47W/Aw/Ncg2S4
IVP0/4BxPQWP36/ceFpClIUePOdR6rxa2jPVVvyd4coRg2xVhalYeh9+mZYFNu8Y
lmqTnV3rv7rpSmT8iEtYFPbFgkFQD+kurKNbusqJI0yBH7OrTFTapqbRDoDpwiqW
tDF6BB6+1tQ5qJCUDUpiLVyCJKrpH5dsYEVeoYjZXFn0H8d+TVx7Zz6qYkTZdGPM
fRYxunG9PVKKcIrjbIus3VFQeL0Aar9OlrM7cE8A13c6oMpa+opCNrK5e5Qle0V8
MWevND7v8jEU3rYDx2oEwyVEatbVj6rlpD4f0ravygmcDy96GpU90t9SNwMEsiIw
viZi/u3X/E5swSIZG7h0UWV+wl/8eFHr+LmvCdkZaqtlqvg3gIjWvC0mBUEupT5E
ZbT6MRGJEsGzQS3hClZHiOpaRhhnPz6fffENUWhiSKMjsmYB3bGkB5syIK3+7TvG
KLAlAle38wbAWldjjFbZb4tmodbII0/cMgVMkEiDpaBs6onUSHJCIXYqJpHOuinW
UD/MH0rTZCLeLlaO9d9fglqrEy5duNgl7UWhKEl8enXr++Y/to4ISvEDGWg2x4Sy
Muc26qK1MKsADqb0iw14YhZXNbjmy6eNm5Kef9z2lxlAoaPhxpGrPGSnoB4Hxmzm
omdfPGTMfluvbGY6VS4z9PhKbhbeK7AP3y1ZHCAEUMSopz0U0z++BkTVmjY7/x4y
YzntBuzZOnnlYz4gkxd/bDnNbLqo2rZRofcqW7DrjwFxm+tVpUUlNih305Zp/q46
cYX1WBL12TM+zKmkumZ+a7iWYsu+z5ExtHvE1DZ+JKDMpUVJlqsxdyUpn2SDgqoU
YbG6RJ+q/ooDVgRUJBIiDL6IjsiIc0y8xkCEcYyfUBgJiBZFXW1iq79j7h404Sp2
at1V4MfK2DmS6qfT6TnFUQa4LwzMaq+IQU7GBhiqgSvAeDdTEJ+NjCgUTkJerhtW
iPl7eiPXwVEmTMIkmIxyk5egxt7bl8AECoSexTUXjDA5wSVltTi2ki135dJq8Y6a
LPp5oY823ujzuDzg7dXUKiWtPkbQSGTp8x5sjUlbiiibKi37jFzMuJAQWTt3q0bM
Q71tD3Jl7xvSUz+rOvcT7zpYCc5uUy8gJnJ/8YqwEEcnneoJJaZ8KWt5tRqOTXWM
KnoqNgb4KhWynJvQoQ3TkzH6SXtKgEocx8Ro3xeiKOyMxtvxoVnHLIeFCaZYMARk
tK/jbuvStMCwaofz6fU1BIBEMmJjHiTjhomgOI8LjBKVKnlPJ/dIp6UCeeQlLMaj
UTdAfurtbGxhRzaUmn5mKAhfHHp7er+uJ3ngTWWwDTuvEYg9XXVLjHAxpgLueONl
7KVHy+8CJKhAKymwyNAeGX7JbVtlfNRVqooVTk49XSevjvrmrComXcNq/OsgraRU
G1xbfrmI7PVMabY+nKcaadFW681qusBoNsPws/STqgSQvDWe6jrurkYYo9Abyyj3
IGZmMH/e5y1k5WjX72mwfe8BytgIx9nCGXMse+Zhd1np/ZVAszFeWrrMAygbWuIl
n9bbUw+Y4lpPHfbS8Kk33AJFK1UolVyZ9DGvgzUkbCVjCImO/9gma6/ZqsocaJbd
RqISIojBhyYbad52jpTXCDeq1pusZQ03DcPUV8nfnbxb5yV4PwlWfXI9wMxdVAxn
FLNaPscAdkYIwWe9TQr3A2Jslx8kFHZNFepy8uHp7hJ35H0TvFXrrJDkRy9zgGlE
UVqYBGlm9PY2ZE+1gJzOBi+ZhT6g3Mx57E3nYk4MwuOjVYGoTafqPY4ysfOmtWFr
x6ScO3+d6vsdgO3LJB/3pDcWN+a4UfCOv42Wc3zK+nCyYnr4pmLAUy9VcwNfIBu3
DSb5m8ehm9tpSxZaR6Zp8fY2DhwDMjiSMLyq809TWytPWlz3cZ5MuT92mc0ki6Js
lgose90+IoVjC+3M2H/wkPtu2U8YU7sBGCXxrlKKpZUlcpEsOWrTIMw/Ylqml0+V
WegbdSLx3SCheQECrqCxAaEb59nJkR/4xK289PKPkPPpHvmVO0OW4LzzQcRx2oSa
9QGbH3mfdbmEDJshido5mxpOCS0czRftZ8frHP0jVusioqUiC+eak9R+V1Tp3yya
5sxnZ4gp0bD2m95oj4BX0nnh/3osABSYi/ITP787ErvkQ/Vd+dh36WzbJk/Tu1Ks
4ydOipMYDKUb+BFyoNKQ5zbFve3XCiQ6GEbguZjRu+B+MsURt952xhTF26HwVADw
Fw3h1r513DHZuOLSKaW1QzzfcxsrPlZnFY6Mk0PrS+Q5akVevkdMBUNAkfXtAoT+
ZM/+aQ2gZmgWg0LUzzpgujz+BBpJSrkG/XwJX/tHTV2I1oXdVbjSwdxuIIdHQWjr
fWAPxXyFbewWpwC0IhR33KcsWmiV+iQ4OQVFMdo2iyLfWl2bLef4oHfbYWvR0Q69
IAwc/kfw0+grT2rinpVgJTGinNSFJzpxWuKVn9NkHRfgL5Pn+1/p01/Iv6zW79fL
RbfJoe8hK8kmdKwpQnDOOdHnSHxAESCNPbrsLfx/jKEtN4qhU+Db+jQDpGjchSQy
y5ARtCi5kxegZloKQNfYdH+s10qpxHuzpqsalczrkbPXRml0t6m9vBosRNaHbnmu
fW7DlSl7UV4gA9gbuEOsphARWLTFSn19ukggYWoMTsaZVUWY+RJKS5RBJXV2ia2o
u/J+Fnp7ZowyQxaR4lgZZEMWXI9+T/YDmZWtDJoAsKeIZfEuULgOh4A6WBie7ku7
xM5W7ASMNjzroVgEnbMTMFLTeZq9/ifs5NNDQvFwALuhoJ8nIuO7yfN9sI2d2ziY
8QKQtA51A/t+uf4WyMs1FFKggmA3xgg0WkfkCw+OUwDH55XULogzC6IBiGCtdX3w
ImsF2DhS8QMEscFXQNdUjqBqstl4drLZG0nVwcWUDZ6tciiGaVuC9iHRjcmmCdoQ
Y1I1QAHC/4ggY9b6k1JbWzWqbYZHv0D+zfWqFtHvyiIZVNBdVEpvH/H1qZ1fZzo7
aWjde2v8bLssQ6zeaRXXzyP31RkSdmHVzhDBJpb07f7klXEV0X8/rE5i4cxliKnK
ACVir+/b8GejKGLNxrzdvKse4uM88hqGe9j9cio/UwHqhTXcMKGDlC9D0FA5Lfq4
cACIeA5H6iunJnMGO4MOMa1YDnT8NmphN4lx3g8S4moi6Wrs/5Bd5JrfKv0j8Vhd
UZY/vQmDHnlSX22z7qbn2HzEHfqGV0Y0dT0TNO4apIs7MVBfI/oY7K2tCK1S80Km
lKR85GIDMgdIXFXbtbYF/0qjGC8PVUmcKBoZ9iKxbsHbXfuaVBamyeVNmCj+qNaC
IUSJ+fP0kDH83g7vHnhRxUGtzI5hIfu7n3hRoxag2OtqEYGc9XoyWGRryK/4oqjU
uiOg5nT6oROrQgWJ7gt/sWdxPohTkWT7o8n7OA0ohxnr/Q+Kgg676IacojRa0AK7
JIzLYbV+RT4JTPIawze0BA9Ly34FedAhgbSBL/eiX532+u0ApHqTmBCPcnDFHSc9
zh8jDcDToUFD/55lxlZG41DkVBcfQSJHppDC5SZp9pDRKqrlWiamlfVAY8WIrOlb
nGLfyESgo2E08PMPrvGh+JLQDirGphqcMJRW+CoYQVth31xOrXjRPnerwFtORk9h
HNJJzmgqOpgM4c6wLYmLFKblsYcboqV+FRbSJ+SAjpC6pu2M5uhHZrI+obvK96sX
GakwQejLyBW0J+qrG3h/Et5WjBQjL/+4hvbCQK6ZaMTu5fxMjX5GOQ42tn99SZvh
EIVUbuAK//eYtaUTtwZ1c9fqwXQfLI0GMAW16tJPI4JHfAgQvvfCe+RDffQoHuwq
mCLv1KZf5TIE+zMIjclHoWpn39gV0LjGPOCCnlSvy3UsLJsBDHDkaCzR5IKRvwQb
VE/hIofTZ56P1Vk3dc92+e9+u4s9sLJwFAGQx/H5chwVMvL3TCyfwqZr+7z6yLnL
fRWtDcbfXpvpWBjsrovKlDHZ61g183at0Ezw1t4cG1bccrAs3FzRuvFMgdQmKJkO
Zu9yRZEcz1z0xZ4G/YSKN8bMQ3D1XcfCSGYIJSncdFQa73ctfU+ZRHAatYj/R2Zp
7cIvZoHxwsZPZmd+jXjToLB2C9LTeactY1uGnLjC60ih2TN/iJGuyRuPYXNO0v/l
sv/98jrWfwuHIOxmeohVikd7g44sqUGeVtFhXCeEOHYPGv0Wfnuw6CXzjtvJMH8V
3ZXu9MGo7RptQ6oY/8MEl3mt1gj8fjg4ob1Z6I56YXxqiIH4JM42kZyM1cpMk3eB
A74vEYszDqN77f+cL82/+cYhcqPVH6e4T6TurHtMLsU5IurDbcIHhpcaWzgrNa21
3ydgaXZvttf+9dYhfjLIp4wav1h5tpvm1w24QgYaHaZ8b0fZZZe124JtWRZuQY4U
kRiiDpmAmleu31vTjWv/jqI5R76GLNp1z9j0HtNtYEffOfsUqR5FO5HShZxPyhey
W3nZ5TQt63fDXe38C+v4BFu50nW5UibrfscfBrKmWSERP6gmnNOefdHBMM8yRtIR
BAXqyE3xpe2CdfKctbpk9dhiBevPb0+Vy4SN88mKb+Xu6m9ecFLHgatj4hmEmaXJ
a/NgtaIF8t79ZHBqd0VCFhiFl1CKRkaXnXn8YgpbdhcN65dGg3RALx5KmHHwy94v
I6R40L4YBXd0e5rh9BM7ExF6pcrLsZzBHfTAxu5yTLXqunaRrr0UVSnU8f1GcCEy
dbaj8aswlNWg6J4Dlkaz1pX7KHmRiASbFmFuVdv0ccDge/Tba3tmt7bc1Mu8cgpw
xVC/UVGoxPA56gzaOhuUzFl8e+CD7mmskfSNxtRdBgkqLlQBabnXkSykgd0r8l9b
OAUota9QKI5PV8NdMe/q+hj2764S5FngtRs5L5+8OzRzxFSZM2LWnF+nc4IxBVyO
kmSRoXs2+hAhaUF2C+xW4Wsvp/CuajZU3g3O8PeQP98MiQ4jUqjIfvoR0u3n9XW/
/y7YMz1KwevKQGlABhOf4mSxh46yd4QMiupu/7eZwLqCo4R9z9eccabL+S89hsHG
R4gW2Y2kng83KNujpkR6cy8dq3cqU44rtLy1tBRQF4XxunAqO/NsAtFsb4nYQzqF
aP1NVWwyQb2TIb7Amz9xg20yAwosJHodmW3+18So2zKk+cAmKvMejQL6FgLKvQ6A
o2tX9C9OfUz0qZmWUsmG76NxvUIXaJ0hQnK+UEnnqN9D21zPlguhV/9P7anwFYJy
/1YXUzK4b/NQWB5uzOsEpLhowozFjEj2WKvGpUhKy7+cX8S+kDA9bMm4uzuS7q7/
5C21Bh+ZKw1ZkNe7zQMZHe8HlVrPI2lu6LI4GDosnBmrZbhDwcuMi2leY4GMXIPd
uB3RPMzb5s+R638IfDBZkVFvJyl5IhiSgP9mg82qY7DbJ9KeGg+oWnuTLqJjaj/3
C9qjKkcLlLPk846PBtZwZIepJxPbSn3ioZfo43vLpOyUIa5B3kc1i5mcQhQouYyp
8sqqPGRHmL6W833Xq6M6UgnZbao9r8r6a8EQ+Wt5zXcgDAd02UMkdtaQs30PTfZK
h035a6f58WCU/2SYVej1kKc1aRX6vHHxmx9zGMdoK4h6N3O70ysQ9oDWoWXZUbAw
6sRtsSdEDh4HjXlGlWcZOYcYcFKWB+jP+552F7yqXiTvF+H3hlIQIl8RaXbWzONl
4kKnW0Qx3ZS5TC7Pm6yfOs56tALxPhG/3TlQXj2B7FiYvAD7pp3egHCtx0LLLvS3
/6Dw1hcK64hvwV8OzLcijpAwRs14Jb2psFpuEAg//mLp7PdIyZO86EEtB+Q3Q9WB
DFdp0G+G0ifNhk+LNXw6ScxwFyhdwi8k9UPK2nDTZdZVvH0YNIOJ1YahyQ/v2Ujh
/S+Gu0Kh3Q/aTHmqZr0a9dhWC6r50iUGwwxGTJ0qEoCBFxTgS+it0SSTYbwAO7PV
1YmH70bOlHLcaxRjqck+qinaf8M15EMp1aqg+W8XoXlGvBryAMa5PjqIaDHx4Co+
xQa5KjucrjcYnCA3QdyrrI/QJtHVIDRrS1uX6GIg+Ywk61+1fIoqN1qmLYd10Xak
QaMcmKG8kFLLGruVlMt50C3KNFHfktIRS/xwaVhsIxjXipaZQXK3yDWFluCyZe++
vfoPRbqKg8lPtqms6IW+3j584gYHgMEdwWj4QOyvRI6i4wqjrBPhwrfK1TmLFOIG
OKcZG+5327lYi059Iq6g4GFZHVFVn39NBYtK+OhZVhU53jWsHJ4pb75gvGB9rNHI
DeuWYRzTlTdA7sjwQivPsLwG+Y79aoILJh9QZpWSASE19hwxqTCGR0foj22IoKAe
Bcmh/bna8VLHtysT6oeToZNTHToPL/gCf51+FDTCWX2qXzJBSwCQ3k/EfPEaDDWw
G+JzfjacutrO3uXIfQPmvZVtVwiXHIHLVptjrxVrwsFco5O9VL336Uh2ZyY8bHMf
K5df2mHwcV1KHCTv9FtdwV/QQrmTuzwSmLKZWk6KMUT+c495QRgL4ItYSp6p8SIP
FkuXa7PWGYnyVk7CgJJb1tw85nrn91uNjSphYjyuUhK78ctpaX5lxwk1BGIKlz1O
Kcrp/2s8c3D47OWFCqH0G0cVGKj/DEJnR01Og09/3wzoQ9a7uI16mQ58Dfn7GNlX
YFwtd8NBcBfrZp/N3cDONN4QWCI/nrG2029tkCFqDN5dRgvYAuHugF9Pfwn8+4xF
WMlkUoc4sbsCtqB0Zm0WQBfYw+r7KzOF6KBgiKF0/YOU4bPFA8OFs7dJGnWuMmYM
mV3/hbk9b0NOwgRAshQOSHNy1LZ465QP7zAuLaDcGvJN9fztoYgIOnYQ+e8OugxX
USON7WgXRDCDmJq/oi7W+NZctuLo9oJ2nzp1K4FL6/WL+W5yOIolDS6+Qa2hhXgb
V0Yccsbm/Br+Fr3Uy5idpdcbG4PHF4oM7OCcAlRQBgR/u0DMQhZzkddSu/9KzFSC
HtjseoINIgLcajZ+cfcWZwMWwMDGR0XmsRtFuwirP1w1Ptpm1CcGVObNkd8DW4f/
VxAoVfPvgiIeNN1cw+hPw9/X+z9arwfdZUhcs/3gbZXct2l5O2Nbl4ULWNNvwAXC
/eWh0hgl9+zHAV3xb+s6DjeonYqaF/qjKWEE6U/FEWyzgf/njDvWm22fi9yzCiNl
a/8GaQYQxkfxtbksBP8hXLJOkj4l/M5m1Dg8fcCNmTr0zaXDsLYvprMZOvlkzSeP
bFz8uwIy++cYzd5/WAxcHZfOj6OYY1/FljOAcljzPld7CkiQ8iHYVEuE5Jk1hI0R
cuXEu30okyUAGN/S7KNI+wuO/VhIWt0t47x0wLxEJM/5KFbMJ6+wyTq7Pyiq1P8K
zw921B+1ZNV+CedYT8hCjmNAlDEYYYD/0O9lkE9/S8cHm1WpiFirfKTYr2SmWP83
uszS/NhMA9bBoEAQpS6sUdF6uKCGmaUnC0Fg6sOl/7/vULP2T7kufkpTrcYBaFz8
90smZwZ4jksGoz7wM0ukujqkqQYfIXor7rNVaft/i8oatIAHyENZJfmKJp08uHIl
0oeYDFEb8naHcx0tllGTCVTXWZ6YaH+6i1niB9tYpLhxtvHgVPpWg12NeE6HDTVG
h1ho6DOfNBrTzCa0uHulZdciQ21H8x+FcSs+QQ+nHfMTKoY3A9TCxWO6YKj8WVJf
jwbW6OyYFBqxoDUfyDq7/Uohl2RSsVuY19uGGIaGVODwAyLyLrmZqNCSkGHJSU5A
A38+8/i03WQe7kQnF3I3cyHOLp4Rgj4aISVCdptZSNP8OOZ337HLRaKwb0dTmf/p
Iu+TUGOSBvI0v1cRE7VMzSz9KEuACnbhZSfJqU4Rtb1kZyWoBvkdiq2+4oyg6k9d
AG19AAKgTOTs5WY41zo3IPuhptXNizRtG/TlJbKHhhgvut9Seq9RF2+icn/TaFfs
cFq3N26Q9aDzV2mMYd+MxIfGwjTwa5gcpoHBP5G80j9x3Y1BnsqilQrWs+BVZ7Bq
1nRC/+1ZNv+MytGB2x9MgxFR/11qaw+UslT2l/Ikh7QNcQ2FcPO+bX9c5dCNHd8j
M2UqlcLhDaB0jdSOY/4Ds+TIM2z3gPyd4toXvwW60d0mNgaZz9Ws1xyqbSq2+aew
6IYZ31/Uv5gjI3fRQmLxskYybu7xl9cQC4oQhoRQdoKUNajPKW4OqopubbDnY/cZ
ORhcNT0/KVTMQtG/2ofh7krUz8LLEgfYrLUe/iT/wWplTIuS7JcQvg0UzQGkowIi
vur7Z0V4rbvL77Iuq/C1TOvCw+AOhwCR2hFgBAB+TAiqegVJf3JqwgvmKDKZKMbd
ehFZTNlBuhAQmeoSF+wlewu2NaY8BsmDPiV6lw+9KRj3ReWiu+k51Wseom2VSK25
k3YSh9tP4zibLjJn9oSnW3feKsBspDVkrBhQ7/eMIaidGEcKP1r/IPetfaQLTmbc
z167y1eCYSpr/u4W+3NSz6kft6jl6cpdbiVogHeqcpQuXlAiNiY3sGzaxp6Piutz
3Nf6ULPjei0bIFdy3vUfdFc7UIJC+PnHBdmzKD568jCmADYdmDkDmh8dmMrfZG1B
f2UJ877bthJTymVt4xYgvqAQij4eVNy9nxi16DQmpT6hcXqQf8yDuWu60aHWN8qI
mYXxfZol3NdVzxCGRUASZWydTmrNhprazZcGsQL6j1RARnyknI47/ZG2f9g7040c
97lmnQR0ixiEyVrAsvjQiPKarD7OIKlO/9aHXlSza/LNQenBhyaBUC8kzLKyJmTU
VyqaLNFC6MdBqMTRnRfdt8ukQLZ2Q5rIt8pR0ebE0jv+44XHsiQU8JRMMI5rXW2D
fhY4RyWK7lcTI2lvUzSDgDkTIO7OIjsGJQnOPfYZ64x0amtKup6q9t/fDXHokrkg
+zP6H/LDSo8oqwU3nAvan45Vm+9rspEceVnrhXXS4Srvb6JGN5hCpHVoCwUt2yPe
wU+eRQfQWZ8D1YvgCqfqp5n7X6RIhOAR/BH7pNwNa8C1H0TDorx6twedOsOd7qdZ
oIFdH1BjpOvUaOfZh13hqWxIMBGhi/nht9D5tEvcHP7kKXNuDgLLQAi0G/2LeTe2
G5QdYn9XYuTJ1AaMFLoLL/926Ux0kEC3asab0DgOt57NM9nN+HIIi9OPaWaemTNS
qfDUlmLplCZTKAuZFQbP3XkLaEO05E/p5AfI8/NPJOaj+x5aDD0hWp7LjyzbffBT
/h+Ui/cfym7wppHD1yWfkS7smLIIhaem1w9i9MD0dIAmLccrK5wld0/lB3mID6+y
ZcltkyU7MK3XfTJ22bjMcBuPG/xeBjip28rOE+6WxJcb7zgSKHM+iSpDtlRGQUd3
GBDZETolWsNBE3eq8XM20GqiCj/nuHN4t8HwG1RThEcusVCDCtl11/i7d9f6OGtA
2TxbMLGPxqEQTppKzNgMwACX853uSPyB2xUisKQSaWhpRDNCwSWhqLnJGCI5BQ5D
ncxpFm56CPhepafFmZVet+8vTJkD41iMup52PzgoXzQsd6qtpcjaotbPKYg4FX4t
5HvsD2vaxM35iqN+JqKR5QbqekJnq6Q9XoCZnlCCilyLJLqu+b+raEJDGHptindz
cEykFMuOu4070AGnQOcW2c4lPLmFKDpMgw9qIEDmAR5ElWPsu8JfHeKbgRIYS9U1
J+OPLa4ID1zxUaUNtkfvy/jlrQao+4K0zONQ5IeuD3I3G1nbtLR6nYShXD7EcYtd
kIwbnOVASO9XxfvA7TOdW7v3xpcvTPG28F9eCr9M9dqzL+eZUmkal6M+53h29spm
nURJaRaTwhH4/A/xS8owTq99zEOw5MtgAB6RYCGQ03q1cT0VKBGICTnx5VQ0qKtE
W364vTsPokmsqsFvBU+Nw91esmChrHPhDeneYZ4YV6w/yu/DrTxxKrhSp/fznceV
aadXWhin8Se1fN1/eGP7YIYdpvOYbKx2MUmUBCwsLGfqZAyf3gA+hc8JKrjxvgGH
fPsWgBSwHf1h5XNBdZtxLoM1t90QMfZgqVvNfikbMUEYWjnz6EyjzWykuY5b4MIp
lmbDrBpmGsby9204slIc5uYPAiU29rRWag9XIwpTcX74/IehqhVadKgs3QnsbwXt
9NFej7rHTxMRq3luDBDsGzX77tvUy+HPduu+lAFB8r1pX92I9M7+pHbPc4qD6E7b
ZvGPPrFJJeKW5Ey+QuHMRY0QGjOdbRaw6tz2udHNbsqg3YvXIu0U6/oGTx5LI6qW
dz0yS3Nt82W5D31PC3ZrXJ96JAmapUnMAHalaZ+kwoF3YrVrEiUH0lky31TzhP2F
4Flxn4cuyK2F3FUhauZUUZOs/9B5D62oaTSxIlvoeqLhI18Gk4Sz1vGiPdn8Jmji
l6+ZFmkxSlp6GcbGgquAzQ5vCQCw6DeLtGO0fXLZTiAjxF67dA2QvwS46NMF6xFW
IgFKotlyczdY33diRlx138L4YvQJJpx8/xAX8A/X5260nNAdcWLFOf5i0GgFWyDd
LOpep82z9cmlyBeLz/+EOtVYWdrefGXU9ExpX7xgdveVOs2XU0aXJsPBc5t5I79J
kXR0goXB+LbN+LOehR0WqYBWUNxkWFOeyNy7uvQ1Qez7MwoAg+dm4vzPCy+O0x2U
aEUG32ewro1YRfyId0tWZw7paRQGuMNEKDyTqeEq98unuBOW4wSZfLknlOTErmP2
6gtAQIOPiTsJEpkloDzs2l7YbF4phnZqTZh4H1uYK3E7ZmTsmb8ppr2H9H51Y0NC
MX1DObna2Xy939BD3CZDu4BLTZz6ETcdm6RNxJcnklJBS9mEG8qWnJ6EpsnET9zh
ZsGVE1zEhBkeJGS3X2JV0XJyw0eQ1Bf/z+HYclXP22++dK4mg6A1ga4T8DEiw1yf
1ZGSdy8NHqSYV+lzm+pgtB0d6rPO2HdvS+Xt/TseEXL1O6HaKqFesAFLF+3Rv39f
iv6WA7dSDU9ppe9Z7rIDXNf2Accb+chIC/b/VUDmeCASQHTd88jtCtEQxlRSs9c0
is6hJCBJ09P9QdvDq3CpR967UWusn59Kqx1kvpbSUz9RqKEwRu0STI8/1/7/RrUE
1/ftGjkNK1lhAj1rBbQF/s5VqE9ycHPZmnZcLxfi1bWWdZNlnKqhlpxlEGkcqzW0
LzAbnsQY6utNbqb2YbD1jqGj7+FdYG9iIhnBAcqGJhbydyW/gVZBsMn2WU+jCA65
14sleXGrmBXasQExLH6spb80UMM4zhMI1n04YDEHrKDvrK4aP1Jcf/60wIGo41mu
NuhhS00O1cdo0a/qr2u8Q1SrlNMSvIG7QDzoOkny1wXKTWY1HIS6XWR3HLbgHP9R
jb3CJtUH4nuLpHwN2KAO7QMTHTv/qOVhXcoDv1oIhtxZFZY91wq4uBXsAILG/R1y
NhFbfudcw2JGgTM9KSe6IwSdVnfuTpeWWxCDi02HkYEd4pumFHZQ3DdtPh7BiQj9
TcgHv4eb6+u7ZJDb9OR33mCbKAAQkUgqtZBgW2v1/fBdYyaCUanbJkVsllvfTOLX
BvYev/6UoK4TOgLeoAYIG3hPL+CATsjhhGdxUGjDnXlDg7U81+zMbr+hRHCWZh2Y
+Esl+//pjRXawCXmp9KErjs7EHi+zRmBom12uq2RYtWWRxLx6TK0BsJc9XgSd2e9
LqMRH7c6iPiUzHUgc9Ugfdeg+4sfob+7UeDg2jsfuoBLzXzQWdCMwY8ThIevyze9
7Hb/hT7hAuQjVGUaeTBmxav8e5piW+i089s9qzzOEB4AyHvWeDA2XUWkUzxLny/T
LYhh7FUe0iKcs5pVHl5JgfUJxbzGXIvcPzR45J+Xi2it/P/GstaPLxMUEqRIt9Cp
t+sagPxtQdOySNccTpSR615tGRm9EM96xEtntZDk6GBptxoubf0YJv4bubfOJLQM
5mXkXwMP1EPpy1Gg/2ZQ+MkoENRMhtaQ75c+6iEPgJ6DkdGuQzAHRWMpluWjaF8Y
vZ8QAypVXQ75LWG7NVNAy9RiVBIjKiKlou6pvv8dw9UrxREtU0NJ9mGsarI+Xp14
9QpWliA0qWkgDta7IkbOustw4R9PJ7l3ci10too3PmOys2z1IpPQxXrKCTHa1G/Z
Tg2Ggs/B0CKzpfE/XMNU45w25huJ62xX7zn0lI+sZE9GnDsQIDIm+dpzlB1S+a4Y
ww655Q+t+cgqs8ShBbLZEdGS7P/FngvTUzGNmdygpshnihYPTWVkwitOQQzcxpgF
zYmDejLc1MLRVEtRd+Q1t4izdRsSn8KQ+Ftsgsu+XcioN3HOdBICqBCEdcVvdvae
0B1aFsZcZfO7Wvd03i6WbWzTELGdlF5w5Qwy2RphdvN4a5giAf2iw8CaWNgjzh/v
2Xjkoak8LRzivN/6F4j8psblklP4Gra6WmPyCdXKKVFFyi1nYI+uZXtYSQ6e/W0o
YQDT8b0tEzqTJUwcowG5fYHLGdIgzmoJEfwd8xLnFZdRshIKjK/WK8cPbpNjJEv4
KJct+JtTBPrj7E9T3lsO3cBAxd6CJ8ANHAmUslPM/1gKQAs/vho0GJha2Kt8ZSoJ
rv7N65VuUvN2y8fGQRHyysYwAZmnhw0Z1hA7yDdOThYf1ZVftXTTGvYXdhW+3AiO
r+O2I2o/AzMy3ZUi/rCojADc6LqZn99Dow4ugBB38a3Q0sahJrtVrjnf8gL+1Z/K
b4RevJ0pDxOqq3nqROWF/HuuYFmNnhNtPPGsYbRGzSCVps0ZKYzZlQdSesDrUESP
DZtMYWQyiI8a1E/LNl0wjsZSnirpMjtd0fJXjifPLDGNOqHkRkCz/wlJ4jug4p49
K+1VRHFjph8fEHvew7Xb611ln7m/1a3/REALZvgOeZ73lxX4fc9UAIBsndcYUd6N
La6VMgu5omHrm9tk8dN/ciJXFu9c4ISCVLVtcZcFBBhIZnKVTb97V0heuocPoJHy
OwKFWYKLsTxbuFBhJeZAazgIQsiRXQRqxMx4+gTmoOgRDzAWmf2RUHz/53GAQ/Tl
4YQnAdd+OAVu+KOyZRH+LrdVdPwqZaOBo7tPY1xfOnf3sKmj0pq1ykl/dNEkRerK
hEx7kC9tueEgE3k28XAM6gVEtvYtcTmDOiABOBQWwLJJMj37FxL2GBSymhRJ1wJ4
ATrFCirI3UKrk52EfbgfD9vB8fmcXBwkVZFEs4iGEsKnlPa7NW8F6W8+qGWthqvM
9LWraJQZKG2fnd1iKVEklerTAhpteIp2U8jzu/lHS6/ZY76lSmHD74aK09fPE3Yj
Ax82h6q2PG1tKnJGzd9f0wt/BTVF2FvNrnDyx+keY2GRkuS3qCKJkratcbVPl81l
7Fs5MCbJnkXxEml8RGSlgijTLsAV+5uUgkKivsUJcrOpnYrEV8QGKH6IrKhPPrOY
ev0CDR4SUnm4FayAhRfNDv8zKPz+0xCPqVS+bhx5nZ6Mf66f2QsvCYxAhLl+eOVJ
0rztjxvJaDxW1Fw1qGpMOXQN6XnFerp8eA20dghYzc0/iMLOMnmjZpux8s8Xl6mQ
IBpCVPG17npJjz3fzqXdx5tKHtn2ouqq/8L7Lm4HJ+wngZSokqRCew+lDnnViK9t
NwyASSd+HovkoqsLtOzqyti9cxUkQpWW9gyioySkvuY9N3uu+S7o1Z3w2mIF9Nxf
tpMLlg2Cg7khKcXfm5xkxIyYvqpv8yWoAR/EBM8lrKgJbLqsfl3xnEsvgedGNJV+
bVIyhR+Zii+vEHhafyFNooBSW45IFNThGN1W6UjwQrxurTb0puFLFDugyyYLXcD2
h0SEh8/T5fkS3k1F0hjO+wHUSlj0Qm2YhWg0M9TvxZItyynn19ripfaSKY7DKMwW
FqSEmcW90xkOS5rMdt6onYrD2TPgrtrx8fYmT9y5+GjkOobdVLyLLZvhIFB3lQjo
OHdeQIFFpywFPUYA3EhKKRUo3RFMQPimtPvyV5DqQDlrA1XjbXNVCQzA+wjSb1O5
SqxnMyyoRCVqWGTzZdRdfJklyTwoKjn5ceIQc1G5uPGpahnvStRhk7sCuWyOvwFh
l5RonYSX+dcqhWzF8ewSqgamLLIgqbka9Lzcaa6WLbksmRxlGKLDgFDebe39Ad5T
vf0Lq+EoMS+EXfSFNC1XZU3QUzP2wZEmbqOiSjEgjPB0lHS7z5Eb9/2kxmrg6QkD
1gVfQlkgvgspcgtxhVm14HKqw/O1TRYuofRh5ieC22js03ke7dPeSwjS0NbQzrBQ
pL6OL+D80gCK8KNo7WjxVXtt43Pl5NrNf5K0c5lK1f3/BEZvAUWjaFt9aj60k4ZM
yV7ZOSV4NRMG4IWXcoK9U/EKywj+m9cot7PJ2vbX1gbjxsRgckvBXhuAi0ASXQR9
zBq7FHEQDGxoMI/UqtW5PH1bCB2bmCnzEFAAQeTB51CSR9sHU8lhBBWYh7uGDpyy
FUNFafVMP9g8q9msDCHhrSjyOnTr3nCt1daMbO37acC/cni5fEaazAH/WGQtlMXt
ka0vIU7RvrO+lk6tiEFiRGbvLcItWzGyxFwodEo7GjAo5tWxjbKww1KPklxNLXIU
Lk+hBd8wx6eZU0w/bPPyWlpf3Q7RoRTIoTkmXdchKCLCNra3iJ1Qi9otuzFtZ+CA
n/wbzf/mjE7SrPMOuSsfpzTOZnAq6PxzN+zliFaLIVaB3evHxPB5JjyTtReKjZs4
9zfCv6RTV+h8K6quE7yALsIErF5UVMcK3Y/d0+ddTgp1YWv8qfIGsayeqqXJKMeg
7jiR9wnhKH2X9IGbc0g0ihSLQFt+XXQwyOAsziB4E0GMheExpY8VNz2wqNKWG+N0
q2VLxp7H+m+tXZEkimBcOzutXMDRsCcGQPbd/aQQKdFZ7fEA/gzbdRdizdx/u8+x
RpmYeYx5ZY7ChPBIheDN9RdqJ8kFCnrhOIEWvffWay1SLkZ5Ej6CU3Euh6iDiKb2
tUpnvwvCtz53S8Uk83ljzc5OuPELRg4Tz49DfmXhrpy9KQJ9JzG6Ikxi6LCw6lQP
U6z8l+b21sZhT20xKRzAe8xtfIyCm6a4LkSiRmeakrgrUsI3TPyNEDNBUZeagAOQ
oFZYrpbuWR6pY4ND0L8miIhZsEPSPM6ceIWbz6HAHO9fHfbO6BI8pJlbiQdhapJ+
Reo+rOh/8FtwRsLoDt2paoVutgoiZBwhV6nCJNaG6ms79Zgdxj+lbgB4FANiIa8p
KijPBpA0WB/DQza2wFbkpaMMqTdRSIMP/0oOLfBEyXQwJjBMaKsyB1cbYuRLf4bY
svJoMfn+ZDF+N2SFg3AVo/8F/MHpoAMkFzCRBgMohhUj36y60T/7pj0CGJ2MprbL
MQioTws0SA1DoMus4HJYHODi5HAUl9opsrSTNMwHyxhsUsNE4e1DUvt2DJ9gbVSJ
qsESqSEfVx1G82a7hbMYg72JmiCpdLPPZgOGv0dl+HxVxdpOTHtKTk3+BXbzFh15
zhsKSLjrQ978E3nzoaFE0MapwBX+InGfqsadFr8YwFZRaR+OgFleu+2mBscrjRno
yOgrtG/OBbwke2LnurvlGTncXV9lCHycE28HPZnAri8AuHHXu7RuZNGBkwDquoAf
+6hTBbfBjyS/0hzWpmezgRIctrh03L2AlvC6iK+dwBmmOofv5rn/8EdNUOQXxNTJ
HojztI1QCIn9MQfT6sccE3B+oqTo8D3Olchw6p9upCMhWYKeIIyGuoFdQP6bpQBx
AjHFJVhdnTYMqBX3AhjK4MrgVVq+ZEwZiIbl2CrdBhOxyJcz5jzW42c9bYT5tNpK
5q/MhY2nwLI7NdVOBGfM+Wdw3Ti6xy9gpCN+kCXMYu7yWvzmdYdonbDRUZmzzyXs
Bp9L5Xi4if3WD5HMJi/rkI4KkEAcBETtCqquv1ZIni6rVtVMtRijPw3cNXj0cvyJ
3HRHLfNoX+QnoeDAC9dFlSB0lddC+pGJhwVgfqSeVPc/WL47AgPge/liWKzKkdI5
w9Fzmg5fxjXwfJs+tc4ruUcv/grap3d6JMrtAlvSjQehyF7QoYo7cJ0q3O0ihtzb
4ZMS2V5CQauxGcve6rBdcFytcj1RsLWvTLxy/PCoqyOPeSoeXBCKpRUMJTC8R3rS
ceP9cf14Txj0QGuEknF3WZqKF1mBUx6rDlZpjxzQT6SpIQ3CrMi2CT9ES3tu3Dn1
K9UU2VTKvkKIeFxe2GxVhX8+yLveuQvwSOntQYAAbqzmkELw31UoOcz3UIoiblk7
kvTanb1ItMsJJJuexO9yMd36L4Lc6ZAHoNH8uH2WuVTxl3otkAEAj126p0XOI01i
3RXQdm2KkRJxhBLENwa90PcIvAXnIZC+5Hu+87JpujQrHd4Scv5KY/2Tf2SkbuyP
c0SiAljcBo4mel9hgmq78XcxV5rnLSVo0HiwZYF+XeIleGGEEtK1DKV9h7Qk5lDt
je0xLjLs7mrxAz9+y5N01RXFNulboa8nL3wjepxPazHJEFVSbDVorOAtX/QBZiSK
QZcBmrMKTrvzmebvU59eOwVNBJc8P5zqTkbsQqPZgPuarXi3oOwmwqCKZcwn5CnF
xIEuhi6i3L+FcaYB9kYQ0FAvRIPLCYi1I09h54eGxto8oN2e/6IixwIK8TkxCyxL
ttcPy9C8rGMVRCgGs70ZN4g8E2fwPOI4kZS6Nb81LrfHD9Od5ONNRk5DbkcdsCpI
C2ouDv4nS/2oh0b1k0Wy+9NCYIlWUy1rzHBLFa5e/Y6uUdv3JrPKqZT2Wb4TL7I+
Q2geYRWhELqGVqEgisNNjYEGE/SR9AFickJXMkjHRi3b52q7/MXmVOVPwiwa6Ecc
bqIYMArANB1iFUU3IHZpyQnyTuT+wZ+7pG/N1emc11/pRzzhHQOuK48T0NU/f80L
rXzBJV3Aphg9OTKJAx29qn2Bjm3oztMep0j5UvMvXmtRQEKq7rjvbZuy+CS2N+YI
TWjtwKt2bUGEXJH5AqcDzIipvJslbiFgQ+17IYLVyJuKopB5rp5Kg9n9WeU+CeHc
zXaDMQvtMY02ltkeV15g3aNDG7i618F0xg5J0jD/6mriWBKRQfRl53+av36tEelu
R7HV5uD3PCU7G0UeoJYjKBc1Y3RjqAVjDUQYWy04RKt/YSHbirLbFEliAh2SX8Ss
S3+slfXl3qaI3+cBJk0Vy0nriXvsqOv43MXvQ+KNyV1e4jxeNRWqggJfa/BW7vVL
8bK27Cthkry4Fjo46jtyj8nUNj/MybPzY2cXC9ipOYclnUb7PGrwvuyqjQ9mZfjz
a6CR77ULFBz86Bro+XAyhjm2LbAQgOD+37ob0/3VjzAzbKfwjKRaH47z08/1Puwu
PlldvuoGUQRzT5dT/8lXXhCW9GBcZm1xEq1MMVKROIX3gAmR4algAM8amWYL7oHh
xRJUX+JSfDEGLcMzhNIA3zueTHgHFht9LiGadk3yX/JfwXvihl3/3Qed7Fn6JLAJ
gZGYnRWS/L9BUaAKqeVZWlNZ7WboG/lfbhvC4R8lfNGmK9wUu+oLamELkNhAvC8h
vdW/Adfxqu1iYsu5Vll/qj3RWDmN7S2YofPDtulHtvgDzNaZPrJxrslFcJHP8fAd
ofx3IB96z0GCqjHIGaaDPRGSM9mjKhqMFNOjFrE5cpz9d/kHrnxvxozFC/MB0Bbr
qXCBGkoKkG2T1gByUR+j6CExlES7YcRwIN3XYiPQGaasDYbhGqUoxg+w1w9wLCuO
Bw2tnxPrrZhRfCTqKW/71ThqUmvFu8HmLidUYGX25+UhyhhoNznRZ43aFBZKh26K
p+25o1u3lYpw32Mbdb78jtO0nltRWOQ+L09CwYWXL+zydEmih+OUEnfqKANmwVu4
qZt4crnRHnwXBZiKno7Zfvg0PpkBJtGP5Nr7M3HuKZrQLeO3lKbKxLfQa30HxXw2
f/qFv4xxyQqKF3+o5++nHBwlgKRHAeZ3NNrX5noHkz25kNQvugZX5IOI5idF7a7G
D2ZngHY/ovQCK+Cf38G+9PEyNiYs8Xyfm2Xg56UH5h9g7VbK3CSeXPUxss+ygmu9
bSzYEosQzqA1z44jPwmpxqsZLs47PHVHVbIRMONS9KQQaOIMDW2MaJAtndXH9F4Q
+qcY8qg+Rn1ioXEiym2XkEYF1djhRQKOsAaEUqyUNmFSPBJqKB6gy5Mlp0/VAJml
csjO++wK+IdcuG1s4BGN0F6RdRMWC5fMFggK6wFCHK/ln5g9kQHbVMbSQa9zyrbD
ZYvDY5CBSNScMd2MzOutu6junrj0nFn8ZkSPqlsgyhxtf+VavFF21xNnKiMPu/NI
2G2a65obKg+tY+2RJqsnTLB14ZCpcJkv9YWilAvV6a6J6WoN6tnXQIhDTFY6APam
FGMVEUHhIaI1RPxkP60Mhnchm9qiRq4PmgcOPMU93I7kIX/O5IADqqF0K5TyPmzx
OT7E5U1CMgbR5xuo3WAT/Ostv1URs8Zvszzjvb0ePrSB5W0G6pa9kbZZRzAre45E
ELcJVngHsF8hEolD4IOalP+eLhV1AxQ2N7gzNW1M39P7T8TTN37qr1s9kYO/peOR
GeWDtYWR6hfmDB94hotgb6ZonWaALnD1D9yY2gnPa+oY7wrqWtgGvzyTgKMUlow9
C77jUJaxtOxY39ExKRuaOgNGwJNTGRHfjy16MuJs+WYFK8Cse9vDf9t+6XW9VSgM
ouVkYeJRQ61u4i2qfyUYflDOffCecYWMFPXGB71N1aTsASd50/E6+kFQKjVOmkFs
iMXfpvM0eWh3YxqGrTT+FLnrBKiepJMtDYbIM9G0sS1zt84MHHc6wnWvPLc59kQP
FP8evhtEgD7SQp/ekZ+uXyb1GuOVIUoj4tU3DFl6AVC+2maWHpS8clIjabYbJ2wa
hOX2zXvkgo5XFCHfOfRzO0Qda9fvPgWrXhPeXURuW7h7va5UU8/incear+LTkEAr
g3POPWk5/7+p23t6aNI2SQW3bL+heVpKKklzl3fvKRX1wlledXa7xQnaofVvyEve
FOPs2xK+2NpzS/SvyGBZ5K/LS7t9BdyeoINwRI+T9OLOfAXVtyT6rBw7eRtDQioE
NipEEM1zQxiO1qZAEPlcubVi4ZaXFs/J1oe0EtMf4q4Rh9I9U5tZrAQfXtccdiNt
rjkTM0fI7A/rchMyIQwz8zbMd7Wa2cUdthqLWH7JqlK6hkEIvJeKBYFGFUAVAn3X
NEDyxD9ZHy1kTQ8eBjUKUZiinrq7SUQR7AG9ODYkNN7vMVnmcB+5RmznQKjf62Jj
6U6F/ECXSrmtO0DPBlEVbflOg0vg1Hi7M8pNA+rTOEVcBg2ZIvK4z2JoXq9AEHlN
1eddRx31wVw1woJsfytg8SqwiXwK8t2qbIGEated9mZkVRQgPwQ8KhF7cdelkaNY
iPC9MFnrhEQNRm3UGvXhk/MiCq1AZSf0x/+cTFdOPD4oV0+aE2weGEOBDuO5EXZy
L/fIm3DGLvQ+iSTiq1u8Vn9YrMstmTTYU3C05cRqysSAcOxwt9QghUSOhsT6mBuF
oTP+2YgpZSuacaL0qwE9NTb4R+xeWfrxecEeCHkdWI2ArdsehfmfKv45Lv+9ro6N
ZGLHaT5Uo7639jc58bQ1j+FaWVYL19OEDfEbbyT6oXsQkxhcNx4E7sbvU91jSa3+
Qc71Y2S3SYwCA1yuCf5+6/4E94KhJBMpcDnhkQzem2C+4winfLpkjF6Evquma25i
sC7D3Tq3jIt5UFfSvc4U1O08vNNvMTGHe2uqHF4w1KgtTMx/s/s9jiihuOJGNlEU
zwhSm2hc+W1oF/XnXUrXD7new7NviZzrylbJdDbcsdErsuN1v/nvEaD8jY5RWoP4
OwZKAiQ7s+aq8XJySXfsnIbQdwxkX2VhAtMuMKLfQcW/TRNohDR/+dm7VAeJXxsk
nwKm3tdD2alqkdd+dB5ACnMTCSVoeLug8kC3Km2Psz/cHkL25D3GqHDumwiFdSnm
wy+BLaHvNs8bl7PR+czOjcqDEpCOKnj9q09KBQZtm8YNJ73wfNuyL/Kx5Ksaf0Tn
HpeF/y161BtKKEZpdz00MU/VHIxWSPKCgyYpDnkwyw4TgpOVX1eiYe83JSjjdIB0
JbwA3XTj13mqaR7MY9ErCskeXT8HqGrAn3RxQROaJxjFJnOMAhTOo6rLerMLtvZ1
Nau9tHnQ8HGjulpi5sGBVgyCQ6aFIsirx04K9e0DdeUtUrqU9xcZz5jJMzQ/cHaf
xcfIicsz+ywep4aX5kMj7TtuTsLsGmZxiwCLAh4v6zpy/u4zD0P6yP4b2+unX3X5
l/C1DvF+712n4QW3aK2cM0eFk0ExHtAxsJhGQtMad+YC55WeHuTQtYueDFX58nU7
bwCl7h32BW+tOj8Wbq9DaVojz4zGNwhY0AivoXA9mJLAQuPuAvOvWMIOq94TMOOi
XPedzWLm3PQzYpMGcMWljtLuThBBLrZfpaL5a2F1W0jlQkOC/UK1vwl5H3xKICo5
T2R4t0wFii2u+4hz7kQGZECEsJJahvNYEE0JLRrYFEszqInKPppSJlN0ljy3rVxJ
Lsuf4j1mTnhJcoGjEDfXlAGckMKzj/9SaAhORUeqQAp62bi9n8jsDbJFAniR9C++
zxQ1JK8wTz4Nm0ctffvFFLb/RG7wBny65iWgiNKcG0kQFynjUzzhXyGcVdRJUNLG
8NpnThHXpFmc1aeiR7XudHv6uFKYwMFI0i5qA47Z+jkZ0tZyo2kE7jilcPUZ8sJp
Cdcop/96hUYakGEJn2chXHCrwBRdV0sYy9/3twmEXhXaqZw1uqKN9V7USgI6yF5H
zjTeox/AT4F/draadz7doWVC4jLoUssxM6Eak/uwek8eOxtBMzT4af1LjYxo3uxM
rmsySh244Twvm+uVtUqDtyHuVfqAF1o92fE6La9zS5Wo+R1rz769Ki1bO5x5VUHX
6ClVolVRNGuSVehPmc9lwFXmKl5zOWuanVCskdF5KCn17UPVkAcp8gFLxe2iX3UF
alsUdJ+tCdCkRMZJOAlULDfoKUm4s1zY7vWaTrcKi1xhcETzzDTFh9Ciq7FMd9Po
a4QRqGxLJJytWKsRLK+ezWAfi3/pFK5CAPqk72zQHZHi0irawEjHyhC3sZ2p19jc
byn8Gn/DaEZvrMmS/lg2QOYmpUfZ2M0wRaWrlEYoDOEyIm1cg3LwQDN94VTR8OJb
ZGTiJdaCimdeW/bFp1/aDKdq3lyaPa9n/+ociswE/NH4lsOVY60utDoXxKJ3Eg1c
KMWPk2vrFVtDsQtd7rq0SQ+RC+aK48xLuBROSJ6E+aEG2O9EvRpn6hMMaUvaJK1t
/r0X12hou1/Z5UpkK4SVXGk3ST8phpMXGBg1P25Xbr6QFWrfF12Rmp3+WoFwfz5l
gx37YE1Z+7uNvZZSW3/Uf2HeJ8HmuR8yMGk0AFrfHx3fCuvrKI4Lblg0Z4onzYvQ
r01zAvmVmkQThhJuOJZHwFH5eq//CwwrZpSXXYi7ZXio/3VJ8+dcYMfXic3K1SSt
3xuaTJ8Q6UPR4izvqPWqNk+iPg2b9NchZ0Yuc4saKB1N/gE/vowQCdWgWp8yd1Ud
fWpbh6ElOwvCo1yJwmNE9c8VANxqcFb5HWMsHiY4Semkx617E3A9MV3fv/NWutd0
fZbMHlb+1/QSrYpkUrLOcRJTB0XFYKfZJ/XHXz7SJ6eyUNrSJ7n+xOQuUlpPnbhu
QvKPGNb92N/nnCLHsO1t6bVo0vcR9PfmzbZ/cXRdFBGFm8OFevn4Wva+Mwgadqjy
YwojxQTtbQaBV/VGu1T4Qk7LtOT+4DncxoJZB82YJc6DK2Hxst8GZ5xNrnGbPaHI
/YF/+5ih6gkxWpcljUr+SK2vDeLz/0BC21XkPJ+AITiP+4nFHLq9vVZvfG3DxfUF
xsi5f9nYyLuQKEHD2WsV7/yTle7EFZQiHbdvhIqbeTEvP51mFbnttYarUPWSIAmE
T10a/f5l2FVsj09DZ/PYev9+vP64NQ1F4+/e3K0ffC2pW8loru9lCGAnun4BgMOQ
Tgqg4Rbo2jJC/HWppSEkx6OowshyJVsItKEho+siYM5odPafigBajX6Gr8jYMDGu
7FHCDnngHUFUnTxgpmS8bTPq4RyQBD8JZkOTlG6nA3j+DznIhG5DOBoyGD1drfHJ
Y6ctkdqmOz2gSUlPbyKtJstuqrfHQG82nqtP62NKNNgY11EMP3RMkmkQY6dKByBC
KzkciM8WZRNt0iiu76iMVWLWcSs3wwbPex11riePTDUMydjG6cjXoaOalvUNBCEv
aybKu+UfNH0nrT8V8kInUGPx4R00vPWrkFSI7AWY4tmWQjE9vgYLibQnNj3Q2ETP
QHSMYx2AkTdrRsejyMVHAv4GDrZ/xbbFOjLoiY3+oee86QDcLnRBODAO4pM0rXpV
RTrFvPnM5/mtJWwgsHBwNIZVZJaG0+MLC7KQK+ncnmD31LXGUcykfGybnKOOGHkM
EI//GbwIzwfXjqelSfcK3AyL+NyzRuqtahVgunhe60Y3ZVLqN87AqWHwZ4LiMc53
qIM3J7yxsX1rvU9T1Oa3n5KBkziedecrZ0O19D073y5Q9yu3UqZyhNcFedg5kPX7
0uhv4WwPuggEIDHN8CHDELDvAXf9rT4r1hMatZxCQ0b68wGmASHc1/zQjeDZkwBQ
jeFmBWAdViVfXozNTPc7ubNG33H7nCgwoRsabzGfUD62jHtC2WNtihS/UWLou9yR
m2IodwqJRdXqlOQYCxaJXXjBXoca0MqqczdTP5CQ5YmyU5To0FKbz7F9+WKMVVbY
ZWIH9RIuqbAJ7TI1gNMaYYK4aOMj5MG7T2QX3/zFwuuzLq5UG3212qvUS4asfQsx
THnpi3LkqoFnMxtI6OVLSc+54B1gMDPFgCwdGF88WvvUWfsjbY/pEysnB9ixf1O1
4UsVbN9pxMEF7TKSgHQ6NzLNjp3O+pXOd0kPC8FPj5TLpFveFp+NEpLHBuBOT7iE
lYd+KFDJcTOJ1B93CO1uMdpBbvbbcTuM1eEB1RTkJ+3G6HfnD7nk6mkFEPLixAvN
2MyJ6PMq6mePWkaRM6yTVHqy4F5St81lNMqeGLhZHCNeUAzB1wdMh5AHIOXeMNCA
R8h4vMPrQEgPQ2QIrbqwf3hTLIvX+5iAsuPtrKGeZCGDfi8nbfGmsdxbKKYskUpR
AgmduYpqsYx5TPp07z0TyZsDf0+s7+Dkx48lfaYVe8qW8aQG4GJPUGY9iEp9D8AS
9YhPXNTcnVz2ILAAr3+UqE0vLvUZtEiDHuMXIKuCuPwQ7e64c+V1ulW3be8OP9rC
8Hx0nfWJpRcDpDnqUoI//PRZRGw2uYXYd5OchI7ouavH/FBxp3oDGApgrJ+JTfj0
SQOUTnyygrjDb+nGGbrGb2CUkyyB4pCS6wXTmL6mz/G+GqKrM1HTfYPqNGhCoxlp
rwhxAseIiCALHx9Zmf1+Ckz5atC3KDJahdxwFbFO1u8+yB0/QuDcZJfRc1qqio3h
9PoNGSH0i1hw/hPN6RdZxAVQ9W9ROHVanDd+DdJnIuXdLEVLr0hJtSH28GZc5RvO
VQum8DJ2DX9v85pfMTwBk1BAh2+V7aj9TfQngGl3hWkkFw+lKhj3Hjj9grGXkV/i
AqTsbFJYze1rUDqy37jxmoAhC2UIWffFvT8j0UStY/qyyf5F7fWiKEDDz1sCIgFP
oH5xy79HfZFSbsngMEtq5foHae4N0uGRQdPgWyYmfikATQdabPFBDZzq+mNYc4Eq
OtkiuWqDmPy/TCa1DUjZB70IXdLCWKvrNiLMxtvMgWc2lcaUP9zhnNOLIjIpL3yq
ZbG96Eq9AsGd3OQsHO7S/d6DFkic1YD6YsezQ7bU6BFI2h5vh5U+TdKBK1DIfRcu
W3c1G8zeGflLe52EqRmuPTfnePHIPsPXNIMs5dJB8x+EwpPGTgFXAtbBX94VMOaa
ZX1S4mGe4wPY/3qr1wx7sHoigIE/qRW8zbmzhF+MVew5k92cTWX1n6NuMjuGu4bX
a+4hglIKMRaDoRpfaomVMxVzOz0552tkCFbCJzlo4DFOLutFLkaFkrGi19SM76wC
seDAbqf4APBtbzrApMV8L3ncqizs4kgMoQsQecRWgNfHaMvVgYrwDrKxkF48fGHY
ycdtiHFwQoP0l1d/jQv6OgpI8wMa6Red0k6CljZ+yttx2RDu4cqS1DvvaimPNHRd
VnDXEI41qs6FVvRL9xKtW2dcMVFmnutYYvdBy/CPRpKkQVeOqP/9ESTCK2JLPla4
y1bsp2hWFHZ0sbmpqwHrM5l4lq0gKkPPjbA0CL8hOXO+ZKXzM71Y6g+eJtVOydYJ
pVIDsyC8yCGoUj+kY7Sr1fyc8ndVxrqjRmoBMffIPaJ3jU/sqdZR3DUbaIJKHOi0
26MdOLqghoVTOX2x3BpMalphuuPhpGlxtWDFCdU68ql9HaRstKGmAiztLX8MgRHb
vBpa0+bLtWpAh4xr4VGo4KhUiD4a5657MN8sUlWzpzrOrYjI7UbPBlrKUtI4wT6a
pzsIx6+pmXJbBqL/Vub1qOTJhObb31kGT/RUGl/vNCo8/ftSyftlQZDioiAM9Wq2
Wh0QiCmWhZ7GuQbJMwBWKCZ5j446Keqgkx7M5nbwvFVwZiYGLXgcF+6x+Jign/oN
FgaLc2B12nRW5oGPwiR1iQ3zrLAkz1jq7pQ3MRlLEOXKs6LdJHT6RB/4VWyW8IM8
fg0OPG2PAiCSFHbl8QbUyneZ3pJud6hq5gloF5nmD/o+tzYFg8wxy4Xsu1k1HKGi
nEXGw6+rPY7RGvShzodUWEnEt0LFbvDOQI0OIXtwg+wCSoCjPnqLWV6TCHxDbvD2
qQSKPPWNkSOBIFhTkOPpnZR3839QSMBYBGIE1OzO9sg3R7aqouZwRMdmis8U0mfm
nNKDUNcZ+IeHrn+XO0p3CoHofFwifl14gggQJwA249vFUmPBb0wh2oC5pVcwtzRJ
yDF/2Esecnhm6ONV0gTuUb/tdfdzvFsMQjei3Xe+8zPPp7b4Ep890XtaUOMPI4MJ
J8xkA0UCBH7T/pQs6g/gXU8Osk4hg44A5/mEWlt2FRDtx+6zf1vrgxvjesPMQzMz
WDciuwB1kz5SW6Dqopq/keYTMK1F1nDIxh5hxGb7vCQucr8kwJzEWFs3ryJuw9/C
YRDZO4ZKB9viKVVYhpKXO6VJduXCkEbbUtahq5VXsEeEwqJmc8t8bNIrbqRkn5h0
vvmEd5hpkDeqGtXTDUglwfmXE6mHdXzJKSlMpQDb+EOB2cLEgPnPHsoy3EyugPpn
Mf0Ln8jw68K9MOk5kVTdMdyAL9pdThnM/sLt05SE5CfmW0cVzX8MgJIEBdIbdO0H
niVilvryOKTRqutQ/QHc15uHuGyi2l4yMBMdGEqoULHgxJ5cYnhS41TBvYag5vPD
jPtILkLvawM/e6AtqPUdKMJuX9JNOs3439qbT68GnaU+vQJ7CrTrl1cY96XxvNQf
DXECq2z8jpBOQZYPl2iOE8Z7ATbvr9Y4FjnBDHIkrwp+kbMyDp47TspBz/sFqFqb
6ECrMnAnIx+UrCy77JB6dpY/YvjhkHt1KkRH7xm7XNl4saZ+JycDFuGK0OFu3a5E
OoMxdBmJNSCgEYdiVWVe3xwpghqdSNxhT5jU3sj/t2+fjjRgoPYPjSOvkCsvBdCC
ZIl5RVl9BN3BuhQfcEcJiGg7Li0klqDxQ4emARSNA63e/sDnJ/gYwm4RyJeoNtow
yUuIV0NwXULKTLhAphmLdi8bfLgwgNwfgjjgsIenRmao4SXNMf4Xq441Bq0CtkX9
dTA+xm3N/F3xb0Z9D6cqAIluv/SDk2qAqkwwh4oaORKIxUzKsitXptCrrQZ8lCEU
nrFN87qyPWYbUfkvp7KAteeV4g3t+lwbqaSnYuBxm8d0KksbIE6/8zDOHPPUgNND
VOXxc01TYKc6dVXja5PsYrJu7e733bv7BMqEDtmeFAdyZlKYRSDnvU/R44Rx7SwT
bgxpw0pZ3SUB2grQ3dkzBBwqCSS3wjMyK7xsalHZTFqkS57Y+my0GbLe6L27wLmx
X0fyFO7QIDiXVah21VoGdt8sAJDh5qBsnTOEvBVoA+aTxr5YaLJpmd53cyWMteEd
2ZsuyS1FUHUCFoMqcBgEOyz9O2TGip+T9NX9nJdTq7snoSfY5Yaa5hAM0kR/+KaK
vTxOe4byjB4dsKn+xigU/ifhbT9S57riBMsUHYhCPEuYtmGK/RmOrM8mlRAvsyAA
XwinY1jJOMbJtLn9hVlM7T58aulvUWyfAdogwp1PXBjIExW515qAbFaF7rwGip2p
OUCXGDgqKHtQ+MXlcEMpcuOblTi1jiBmbX2QRUo+lw627Yv94ZOK9YkaEzbNRasm
h/ihdkTz0E4dSzRuxZ+iwoyaidzenfNXsCh43JxPWc7/4ZacD9a3oiKa5r4fDQId
jZrvPxpthkAYmkwLmwjfj+ScrxQr3jwwGPnt3cb7f1W66FdKKjGaW52K/j/DpzCC
Fy+8sVtkDKM0a4psoC2QviZPbs5xfPtUwbGBp/hGndMeVcf116nlS1dcz12hu2xT
NIvrbRjl48oBpcFvitqnKTyU7+wbW8MvPWBmvmfXhICiSDKru2fQQomZ3JIEo7vp
LWxaQSIDneO/mlsVa4DRwqsJbG7plAPgT8jOg+3Nd86/rgqgvb0fub8V7ocvgcTK
ezwF3uCzgHvwnyuoicKILPm3OsDWwfq2o3T5DkTPS3yIAFXPPQ+zhziofQXQUqEs
puhepKRiFAoqIMh2xOaKHF3BTOdk4N+72yG7KY0E/yPbc6sRRqovyWbglSvhpRbS
5r/cAOdwqPoio8iU4z0b8KbGEhbQ6M3eTu11awuLH1GAoYsCaN9sBdvTJeb7WrIr
REGGv1fSm+Lo91i6XJ802sae3F2xTO8K+SYP3j/UNJHFPu7FPjTsnVZVbFvXGkJY
km5tfiCXHhqE6Zf8BDlqq9tEdo5yMesFGxLYkYRQbYcesd7v6GQpJt/bZfMuavoV
1nZwpiWq0F4/UzR9wy7Ho5S7292frA+eZ8JZebcQ3BCAaa+cNZMDOAnMm+GXc++h
7W3g5aTHVP7ky6U4EV+YKTv8o1hvR0NX/YMyak3XZq/hNCPXp/xgDw82Pg4hf174
4M+OGcLsZDnno+tHHgRFmy+2m4WMO/RF86hndogIzNUnS+NQTEj7W/aq0/eXYxhK
1cDDkGwUSxlkQ2k+0lDlTJq//8zC7yH4I6HDuCvGayHmrk7Hdam1t8Aoi1k44VM8
yB8ZPthJ3rWZVXaHx2Ev01V8W6kXHbQqQT/AsqS5/Q+8IQMJjbwOJDJpppR6KV8w
ZgjXI6XO/j5w1KWzk6lLlILhExheqrWaeug5kICF0Yhiohnc/YEsXTyDSq4eIiW+
2fSY5uIx6ZrID34vkS4Q7mfezNu/+ejNxod1svuNNQR2626VR86Y2hFJlYSJ5yrp
Qdeere9IyyWwbjjOTg7/C7uupTccGJTITWABRasLtNXbwP0R/cLGB0BM7tF8QDen
cARGMcdd1XpkipBrkAhGAzuHSJLOdrc4hGK9vwr0ujayzZE0IDooxl1K0jLNYlqp
/41oNOPdejjg2ZXdZprcep+ZwPtxW10WUhSNeCpMvSjjydpiCjoH1b4LFztkob2G
dBLIvVixPZYpv/WY4sCy9h/lFATrrBAH64kBb3Ozj1cWT5qRdTOqCg7V9bdRL6Hk
9ZLBxyVyN0CI5Pam8QTglqQqBVGIB+fu/6i8huYDjL6ntRXIAgPqwGbHTUG8aLvO
5RsrFtnyk6gu69PxJw/9rJCBGTdmpUHZbnPsO4s3tZXD9do+uu+y1akJIrNi3wGx
8HekNtMFoxlhhQ3bYNg43m0rtnlG4VXsYwYSYeCDQtLaF1j8cbFFJZB/p+NDG/Yu
HX6e1fITyz/zAZaTvurHKYJbrdKzPeUok8onLmx+wgUSqylYXADxXuExFDfX6I1a
M6Ab23bDrQkFL6BPR14l4ldHZkj59weL5WaM6F2Bi+e/61qBXdle7lyOZjnDM4Dm
pMDfDRiAQy49Y/74lYG+9wWQTnRhlqJHhRHPVgj7sofFb+s+XkFN+ymU4sT2nky3
L1JPnQKr9RtoFoSXNNsg9XzM0M+W6YLJpUtJLE95EkoJfZ+sKwVlpwjBbxkwXZLr
duQV2wcOLSLPD5/Cx13c5w8qlYIT/aA+JXJZWrdbn2yP2NO2xjKlM8HIHycOaOEU
rGl7+T0jNigJkxvGqDYF/p6mXRR2VKIH/ioaxJGQdKQM+Yro0QAdQXLxNcUZAlhX
zLpTlKs5SkwwFfXkGsUpdf4+b5OdD0VCubuf01tWO+yBktQi4kHpTfts9hfCcG/g
8vCIoaW9sO3r51Y5Y3yMbe+SFGP7cQ6LyqDLlmyO8G6PCieyzYxicwNp6GBcU+vR
AlxEY1FeW6UylQK5onn8Kg0DXT/WXXoQclPNamcl93SYFEGbI1kct2LBoCjJnhPN
1H+Z1eU00bf5xxjDMDoTNIhvbU/hanP5H+ZfFqipGQL8i6NYJ/n/ba3iQDe/AkKB
y9KOAuVqxlhB+IeP6lYtdAotKwHzly1wx9pd/1e1M5cExltq6yeiQTI/uooUULSd
zqkRtyuHH1lCd8xXC65rhpLlgFoIuwD+rCyLu/QQfkJsoo/mEoJB12P1CiFA7EC+
/VA6eHSZvMTrROU1k6fy9UXTAlQT4826Mkk1ADFoHOqkm76lrryc4UQ4uWC+K675
9gNGN5CJBsxdrs+UAe3UWY/yOQhFtEba3sJeta0v3jknT29cv4Xzj7Y29ifnxP4f
3gZFYroCr1549IV1csS5L70WmaS1WaU4ItEiQWwh/o5xv7dwp5u7hSJ0D2L7CdDn
B0soYx399dG+dEEyrgVhYy2L7JTNFvE4+qJSPot7cIt9QkHM94YKF6yC3UXLLHjV
zXWwP3frjtjmfHEZSxaCPRqWWzR86I++Qs3hG1ZCVQKo0chXB+QHc9B+YuXWsN+M
LbXBn27AS0K8Dq/9ItnpFAincVvtOTTT7i7Qbp2TB9VPtrYoQ35cteh5l7cna3+u
5nwaCPwF8uq7SZrLcGW+9j1SWC2V0wiEiN5AJ2fidlKdK51ESbqP9X4chQc7q+/k
MPk/vAallQNjU3lKCR0MVuZ7Mt8o6hmrfNiYxGPv5hzy3kLmoJE5t3Ai37CKj/i9
EIpqtIynSd66kyO5JeKw6zy4G7/u13E7PDknp7TpAMETClDv+ANbis48Dl+lhPBN
ZxUrLDJIkAcFzlZUca5aNLQWduhF9pCcGIwhYoQd8YvhyCl73i1ta94/txx1d7Wn
VRgzxwCZz7TWN5Dp5ovYTryw74LYhCySKj1TDz5TPHrXpemJ+hDuizbfaddfIgX/
LtJga0qLWhdVhtpVb+av1sibSthyRH6Nj90rpJmHUnlSP1N8QZWx9YP4l2roPR9k
kYLenV1J7JR4+jmZi7VlqgxzBc2vVcrIezTy55V4u4TXy7AU7BKrAG7fT7p+QApd
Tsr4oUiKEKWWcY09T2IK/LtC5lR7ciULUeQSFLNeEHRyvwMmNSg3X2jhNHcZIeOq
jHcfcjnIxWyQoWvzcUQOTg5UoCwZClzdZ5vc1lw51dTWFUw7+GkRF5lfeZYZGgIb
LQCGD6PwzXcyNmRIJMz0ouq0/5mWAzMIpjpzADb1czR1XBogifXFM9Vnd2W5jlBa
XWRJHvxpUp6ohUs/wwx+3iULrLRT7F5jCr9wj2auMOGTMxGQJ5stmChXgFAfDPK2
mgI0G4s71heDx8VmnIlPxM0P5EaQAToJJOY7O3pXNxuN5Ysa85+RFhE0mP9kZwL9
oLhin5rh4Xx0ySwDyQ4D2WudoE1+l68C7COZMCj/ttyPySAdMZroLt7dbSS/RAK5
qG3EQ6oNirFglsBq+zKLKlog3wGDdjFqR6G8CNjtjoO5i0SPqjaxwVnWuAzvkQRc
O7JmdWiH04E68nmz1YWSGugjU9Gbgzb79LFsfsLGjfa1w0Zl1+/2GlCymABLGbX9
woNamz8yXdp4fdwD3dqQ1wGP83wjvx9IPcRAOaggrFCTXH3lBFl9rfFA1IB8S/le
9b8qjUMiRuqSR04E5bU1dwsVZSCrV63gDcOqDa9Cb8oagp/jOuCXGKoMFaS59h3/
TSIxQny307/P+XkfRblO6H0hs83wnIynvTs7LGWMrkMGgQrMUTjO0VgHcka0aT4j
cNbkpZor/GjBeZZdb2WO6XiAbvq4blI3SNe2o7bKvzzLMtlziz7E1OYUNhn4nPze
s6sJMyk0xCM1XYx2SeT9yS8aj8mEudIIA3sYr18oVhM8ofqyJaowVBSiXFsn+zIS
X6lhqSVVFmSzK5w6HUnFfc24Oek0fTtpkeycD954MN7dxXl/sJhWzfXLniXrKfTu
sehH6dVvm1qED2hB6bMDSDOOJcviw1tEsA3Y3hI1RK8Zmw80tilIdz3RoaM5YaFs
+a4pH7xoIBITlr6+7U0MJqv+KWyG3YfEb53/FlvuzA6dlLHlT0H6xpF5BERRXLH+
62RxlqfTvO4DHyijm28iPLgGL4QAiZkhLVoAWXCJZSWiVlQrXq2tOTw/Srk0GIKT
XTJgKkNwyPMAovxHr3j/42HY7LmuqV+3br0t8t83EFv8v61oUf95i0NOgeuq4RCi
K+Ivhs+nRVQO4hQ8lfo8rAfHX+qwKAQXGLlK6nhxkarEXHJ489arz31RHJMxbsmN
pLcDuSa7H2VhIpDmW+zKvhQTfxjdnE2PHXKFpkexMmD8932lt1K76o9rE5ZtTkiO
07r3UQXRkffq/S6F/puG9zMje1L0vU/auDsK36x695wS1LsvqF9ORBvSxKcSKomv
h8OD0Mcp6A+N0sWbVqo6fp8lO/Ku1g18Rwcn5ftbjKRtv973iWj+fis+k6VEBhYG
nyQBEsiXyiyVLK62GgVQ5/Q+ue2KAmi8tfLzBpNzCjJx86ATDdwxzy+1mzUsEt+n
BjVKu6yl4CNWY3TMZArSrcEbRv1avU9mspdVg9liu+izfO7XQIGZi7I3AORqQDd0
hiV+Dt4GdNlJeNIfdjIqGY/4O531Ktw82WQkEscHF49oOycEUOqLSxKgOVhhyEWr
5xcV+V+Zd+oQXWvZFik2sCEGsGD7ifNhux1FW/IUmad0NSQyYSUi/UBs2pDaSwhL
q4nf3zLluW1472rGOgZd7oc6Cl/qeL9CoA4lBX+ZuYSRUGcqrW2t2nI4CJaOFEjM
l3tzhA1PqqgGaHPzYgW7fipBiyJKBMLS5Q2JW9b8ETJ+sLMkjq0VNHEWXoV26lAJ
iRksXL66pCX/hWYOw5/T/LlZhrLKNC76hC26/drV9gEq/oyXqXfaY81JmT/Z40qK
dDl7qA6auM6SuQi3xP+pi6HxoWq+kdDL/hBcLMBck30UATOUlJeY3Qzmx5zA0kXN
MCgl924GVMHqOdlThHn03C+EE/Ba/lRe4T2684o8PBkGznhgDLX7jH2wVtvnLaIG
9rY/HuBWaK0SZxqSzAbcFQxnpU5FRu7x0KjD/KKRGIZILPyBR4rHEMmUk/cOWkKN
nnygTCeGB8JG4uDaRvuh71ggnQUjmm25mX8rjv0nR3lhm8XZu5S85UZFGU6BYlgt
xoyV71LWiW/8OHTIPTpJJtONpkZudPbPY78Xkr8JCFTHBVIizWtCiGuK8kIciKtf
zsi9bf1enl0ERsMtKer7TZoBhzKcmwZNCCL14KY7SXGSXWLaMEnFs68t3YDV4H2k
ecL7ecj0V//+kr9B37pShEH3Da8oD9wlFOS2zfUWje0I5yz4bS0VOI3C6UGC3BCG
w+owimcFOmYt6N/z4Ol1vG/ZccUpRlE3uBFx8g/HnP3Wj7bmTvfMdReQ8oX13PLg
f55EPoqoYdtfvTtut05TCpnfWk3p9a91OsZQGmDr4WQc7i2/NZAxy5ZOSGAFIa9E
QeiZn8TSPb+AxNVSwhs8qamnCEImqRA9eSZy9IMTfNpFj08DS7IiIH0O9c+en+B5
O8WSWnObxBJaszJu5AkVhznhLFuQk5W3+QTwQAxnUUQNgHm4K124F2+QQSaDwK66
BXvr4M8xu6z2Y38h+n5O3x30BCtpw7M2OjGds0N8MZ5RtOAlniTjz9v6IRB1weaM
/XThO0MYsxI3ZwoqVeP+9wEy9xatm+jGyS/H3L1lJf0geO2tNpGtSnlqGMuBmn6C
CofKA7Xey9u343FbFf3vnzxPmzyHOt1jmxv3bp0Fd6ehPw7T4rjKr+QMygEo5YQn
DfEJTEVAKUqIJZmbg5T6azuaztva/e+5Dhn5udpDr/bY013t5/zSIuuhWcGCekB+
yk3hJrC691ev2GaXmjh29TdzMtVvm9NKHj1qpCmryf6f2WYIjE8DDCorYHxnr7l/
iovEGrqaNuRTKTmSuW293gR5iAwFhmvvp3JgW6T5futwYyB4hzLz1+aSCQ7jipAK
B6F3un6nc1ZAMgPZh8z7HaM/wPH0BSynXuOmUWrx3g3wyHv0MLVrB7wGJkR0aWPz
1FldM0OaBC7PFHfM5KQcAYcOxaeKVe0wng2hRuLr6wJkU5+s1XVPyN4alwNNdQ+C
ebFgsR3hjb7nJCkOGepnzXsv1JnUwnzc32DO/R9gJNjNdznw/O/4CAqehOyvb7cA
wjW1QVRgrCc5PBKi+tPkj+1jYCo1Aa4p6un/plbjFfi6sMaUfRyUDyvvrPkQm8jG
6gSZl04+5gXZcJyQs6mkBSYNjkT2uVVEi8UeqoVAZQs89qLeVuL1tBWscuQhRloC
EwDM/keVaIdB+PE87V+Qgi/kTFP9VxIwaPY+FcwyxW8p8CHK2nLB2nm3jEkXPIXe
RvNOlMelZAO8WxYnIGLvM/RnK54b17ah/89uvUH+4vllTlEtLu9V5h/B564ky2vT
sI1uDSKLGcEAfhVowwQ+gPifi0EdX8Ujp5bYVCAg3u+GCuA5mSBDjBva300xdGdO
UfP6KsguzQbVezcOITFnOF1S7m7Dfzj+k0xxvAFcR8/szBSQXwQnytN3625WYj/n
RkvHHIq0KHSj8LrFNNCVPuSlKR6Rkc9mvCk/PYYTWNV17HOoZ1i8zdUHgFCwBmb4
vPxNMKyq7OeeCVUG4nZirU7HM3OI/3HlRWXX9WGVGV+vx578jFCO+ZZEO5JFg/F7
klheuKaWYMRplNq59Na5GBezvxV0uiU1BPxAsW6FJaONc8pCU7Bh1Nqojae3dHxS
bi7DdC6YDDRdmEKLWKsbx8rM721tqpVHdhYjGzw0gjIlogyZTZg++MKClRz/NctK
rico/jgwg2NasYV51WbxSq12xQPRUqZ425DUv/vB75GXff2ymX7Sn8tNRUnY8wje
39md1UgKmJYv12c+VHMKIIjYaeWLigU9QKG9wRFlQHL6KvTwbviUXAhxqLiiqSoN
NinanGICU49QDJ5crW2Q5XR0HpCcW7sOg2s9pFjn6NcGESxsCZ5x+oPCKnhSVcZd
rNLGfw0w/pWyMtF9pMicTW5bvNDNU4nMKWSK5G+QbDDJ3w86TtL/CEGY+fAFztca
LeRmEZ+hj/Zg72umlK5n3SPo1LIsQqhNr/ITEV+4y9TUCTUyKwfaog3DHCL/5lmE
mImCxQWH8nHg6cArwALg+34BcAH28hOeWcdplkjDvq+9GoX0DQFyYCAYXJujgfu4
VKfy1rMq++DnnBhssLkdD44/0S6AyGvyZO7vFYZo0In/M0+l2FfJ8tTPbcgWqEsB
4cofhE1ripQnD2gZA6uF8ttPJiGzejzg4xHsia1+TeM+IdEJNwTY2Mxr7eYw5Pp/
sccSe3Pr++Bv589MflSe7PZPuL2uuHnb1FZ2JvxSWU5N1syX2IeUKFauEIQcBKta
+EKSNsCa1Dq9K2mLe0EbZgkdP1BIzBaLFyqLmWMLSWJLttJUbwGvQfBOBNbT66QM
Q6J4M8ZVTqvlKLGFHDDlGNnLcjsa7tVIWPCsC1HenO4/pQwsXjE9ylKmzjhwLZr1
dSIdLTvW01Lku9VKB+TRTBlcP9LbmA/b0ykv+h1PWn4qOxmjEDVmYQXaCKT4BTdc
Pbp3CV2/t9fTVNqyfiEpqVfUhbAy+Xst9GIYlvjBh9F+2eWiMvZJjePZwfP+TbQc
861n9RIB98uGQHsDeSxOPPg9qrlsK3Mg9RotdAP5d38uKF10fgVrjG7FKecm3NW4
euG2N9Cdk+NRTjxP3AqHEYXzQXfmvLa8PQd1+9QuJFQJI2khQvSth+5XlEOjEp+P
PJNQCzssRE4FJsSCIolYEAChtG2YVhPH9mr8ZeHWhCs6VeMGscJYKOV8wrL1M45G
Uz5q1U9CtsqRnnkdSEkBriQjlP9aYKDB5AfWfwQ13nyQNo2ueuzn2B47e7PQvyJk
k445WnduXL9KzT5uU335J96qldyiOdzx5vkSjjjYezB/Y7YvZ0XLFQjm5tidxMMB
9bR4bUjA82InaKcgznP9gcW2rEW7MkJcF7ETV8lNIN+L6fBFNTPgzVhs1cec/KlT
RV925OdE+aIJKCf6lXURHW4Mgjdf7kiC9f/DNvaiuCCPdoNqZYMFKUfxHwgQoXCG
yk4dEuT8HuQilU2a8YWWL8Fvxed2P7cAJJgDLEWbLusVPtDee/aQ92XQHLuEFvzW
2CRo9CYFOvOyI+J6nllhcR9FzQvx83Va/2Z2aR6hHKgRcULqr1HpVp/FXdLGJiVO
fM2gVerakKlxnl4fzMVfwRf6OFDl0jeyDp9PlegQGmqF6wkEE4d9qJH82n91jysW
XRgEFJjQ6fbb5IiAEFScr2fC1Zw3e87zELhYgABqpoPta7/W7QxsCoJOVv2aOQpy
QYbnnVfjRR5Qwg8ob5PyhOO9fVOt96ZsL3XfGsodzoLafZ1ARVnQCveqmH6PXOGm
lH1EAL/wW3iI00bgzxBDY21IDkmMSnWvMvcSjOFMB+MUb3IW+n0IoU7KxwxjcR3O
X7JxDxuz33rxdTmbAXrBZO2WqhtS5yxnVyTs9V2H5sv4eoATookIEROqL4NGWeuS
3hDUuyIbiJiFLBsTVZIRI/NULBHmNw84uDtvICPVDDCTWwWXwZ1Pf210R5bdjKdg
UL0jJ9LHw40URNR2rWDL+sAOlinXixzZCA7BJ196ko5xQqnP5mtvVfXJTuNhfi7l
7GIixJ/VdJ35akVKnMxUsnTI1SAK8qBhfy8sg/arwfIrgR6206M0gwG93yCVviwn
5NYNFSuRFYBYGlsrDDvAShgebTWx+KG8bWwHblSypGhR8f7EE2G31rADKgJpAEo1
rrJEJfc5VhSv25/s0vXCqXzsqGWZw9K26jq8bVhbquSayAEOxOmARIXLt0m8JQbv
A2iTztIxYJXVV0JC7/j3HYBJ5kCWefpQu9uUtxdsvyYvDlyckWFQTrixyK1HN/f8
i1Cw6twa/5UqOEOOMXNHGl/CpzX4KVO8/TrK0zsLkOj76oUM+SxmO+eB9/3LE3JL
5vFCws9YUwlfPg4cwNmWxaCnGx1zfhMD9tQeZhZLCf0TIeTllaaL/lY0kqT2JhPF
suYjLk9ZJjnn7NlxQbnanpB+H3h+DMEnCxjeUztk5526bvBjFNwiMXBa+B5EeoNX
qmGFviiIb2gi9pIoxw4POVa5DPAo7J4poeJ8s6lVmRQdgNrkFulD94bJwlT13wA2
Mv+kaCar/HaFgBTQUT54pGwex1PN9XZ/6nBPKVXKidTHIQBJ/hrOeEiGS7/hNdtl
CxNSROPpkYCCTXbWbs42B5MdTn6ayq9mVmpBMwkzoQxQfFEhfgNUGWTzYQndB2V3
rTSXRrp5/eSg1Zwu0yR+zWrLZ8+1yR4bFLdsUuHd9OFyjM57mqp1VXkqfp55R1lo
Kdmo/oPFMWk5oBtdrt0qQAQmRkp3/F8yA0MA62Xop67sOgwbN6IzD3OtaTwpqbEG
bRJ3kKtEVKbq+3GcaxP7Oir6cvkA0hnl63MUOAQZsNuy406VPqdz47cxFj5axeRh
p6Ta9Od70F+S9nKV+musl4My2LU1tu0+yDZnDNzpedKST1a28dcx3bX/XEbowUIS
GW6fwoDhWoZWcWfVpTKnj4Hx/RI/U8NmekRuhp6L5nZv27djdBDmcFgQdiu5JXJq
xGqk9h1gY+eBnfeN/Wgj+40gHtKQwH9fdSiFupNnAHbemZdm3HSwnKE1Tpo7pOj2
2uvt6qjVwjKul7sS27jzVKNELec9gFYvhh3eQKSqOfpzvAEeJRCg3Pb8yRutTGDC
cQRA0Oz3nG4khB9XF9abbu1w/gbEVbyQeDLDobtIP3Eoc5tCYnECroj1i2sW39em
p/j2kAqOjtnsQGoceiVfP3Yt50ZRD6NGkl/xjVfUrLJ7yZEQTIEV0VHgRz28rZHR
dQGajtzaWJci/7N4ULXX0o/9hKssTnS+wD4YHG6YatLNjD/4DdQ2avKooEmGuNO+
Lz39xi1lgq7s1S72JRc95gqrA24uIipQxOd+HrPbg0k0m+hIiReuXm65uijXDxO5
44AZwuNSyrho/vY6/xVmufSdZrUer7FOxDJzXGeyotsqtCEf1QLNQqi8uWSkGBb6
nQFnENCxxfTzDhImxgD4jilMfDYHy/GAr2Rnw32Baim8Pc5JvSgl6M8lmVQZ4f1t
erbJ5GXtj1GZd9tHa1T43VlxaltdYm0AEVedLxgjzT7qEhnts9LlSSaOwdv2hYxL
aB4QNse+6JcAsEI+Ozpope8j51Q3caCKtjP0WPHo80uxUH4Gf2DR6lPXQBEheSdp
yCqmFmnnfofYaJZ+DVD9DUUG/4houbgCPDnBQbplJXDAW1C1rmPVimjyXGjVH20J
/As0pgZNmlUgVexMw8JeYGGen3lxYrAzqLwlYNIZNruj+aW3TbAeTy/9wrtOHFMF
7Pn6xGoqBNUyJYVwc2oNe6NLP41s2Ky9siTmoKJ8ZMWNeQ/MdkOhKKvPAAgLXdYJ
9lbqIk37Ie07R7HawlOxOCVNe2w0//ggs2Qt3HlDXcHAVaDZ1rFuIT2h7Es8K0Af
o4vDDIvnMZG3cDKafkH9bgiGgaz81prHe69PZ2XsWKm1WvrKmILqIJYpdwYhFaJk
ANwnAIlaRyyKMhXnXzKAIm+AFOxlAOs5N9F0ypmizdU3C1X3ear+DzYmcOjTaGvo
BvXH9RY/Yj2vN71WzqFqXfYNISsW1oZelr/uc6pntPRuCot1PsjRaF6TIPN3P36k
jhKsjWDm6YUetwziAu2c9ySdowOyDVk7C5WDKxjLJl6PwMQLVQ1bDdlvOqLjJRV/
/pUW7Fwk2IpoUg0aqZP/XezL133j98vqfS4kiMqYpIPZqGEExOtJwz8/dRQjpb6b
9jB390X90Afhy2mxdAK4yssfBIcJqwd5mUrobK8FLKFz3tTPfVko/pYvTs6/aSG8
AgqpfHEBxTLEaFfqygGnK9QR6gVNomnvhRIJEiG0USXG9G1oM6fabkkcxP2Rupk+
WTeoMxCR5CBnrNwGdMxp4QSaydq9YUFqXpQbkDaKUZ2HEIrIFU9fA1+Ivcr9AafI
rW09BNTgSuPDp0rNlVhN8lW7CRHxH5/j2kLSXsM8iy+YT5DJZrCoCtBTC4Z0CStH
zAYxOFwQHMTgfOXocqf2qCCfLTN+2SBWWyaBjw7zVeEMtQ3FieXi9pAKwPTJ06gu
P3hWju2WMA+ZBq0F0E7LIdYMvEN1bFW8SiJCRYt5ECJYIp4RBm9IVlEgFaok6g9H
6l2zWjxVnuRieq+dTnycuuKh2GFBcfZWnwja11Ihf/hsRKOs1J22K1C5JdZR2ORW
9ESMcbF+28S6F6s7T4sRRjfWPtLITOU4Xcl/upQLC5nzD+LidEpvuWrmFwxOv5Ee
BflKsYGpQmcGHUm8FaraskX01ZdL3CUOi0zCzdoAJnovuWv52gbIrSWjfUq7ddLv
14VuFOddaMe5sPpucvQDQzoIzpBQUg3xTxt9CCSub94js4o1XvSper+TETdTYvdn
pPWush7elXHxh3Dwqf0y0pkogc8fR8YzVquTc336ElhpQYC6LhlwR4cPi3RAz0zc
KTDgVhILh0XO46FmOH0KwfOZfsCaX9x/npXTJNICVSrQ2ZEEYtip6oO55PUu38qQ
iNnNdzv7I3y9gG0T+3MRWa12VboIJxob8VTRnqp+uqkzl5I3pihxap6ljxEB9nSF
jDa6f7qvb82BeECEqMuyOfbxrskRe8+VkjBfJZ3H9Vautkw7e3I+x4NWwBrcGsx8
FegYnkFO6oYpZtwPFCRhY3/PoKhvYmD5dUdZXI2IYiZFiUhqUrEr4V4WLF05Qb9l
kyqp4HqlUMU9GfwNC+dFS5jolIgjWkhLOvjfNu2gp41REDIlGWXvJp+KdV5horUl
wIbCL6yTcM985fCB7VfFChBDWW4YvGwtM61wmaKRhazfoc6rc6b/qKkfHuZeh21R
4UIIw8mCTq5g74u6xnrp0nzut/LyVTCggsxJqWNTQwvEdSJ5ZOMvzojew+0IRtin
7tWc1482TvBm3fj9uN6gVhyOQJuKk76pfQiMZy4s3w+wipCUZbHPtbhEej3IY/fe
p+qPziEYCWJGfkvh0zUsA4FSX/ASjMnOtDuB37OD/kJxcAvsjIRYKRhxqredI+41
zhA7evw9u1rWn0mEXM5Cj1f9MicQLU4UgNwN3fQwdQ8HKyM0VkBZD+S1rJ16ADhi
eFdWzBlgrQx3IM45RMUqH+sucbDddFwGvEz+7ZXHNCWLob7JVvyha2/rP014k0Ug
aLQ/YXUDGlJ6GbdXF5TZ417wPMQ2x5G8DKUD9GvxQ3GRXvutlwWO7007zH2Yc2JF
Pw+il1iLP5O/PlEWnmiA48/REZ71H+udSaRt0XFMB1kyT+Em5FGlVJm8Z3l8t57p
SRgkDXt0QgCiHNXAqHP/Z+psYqZSYgXQQwVmJ6VkFdWOxbec5kbIyIyY0F6t+6w9
B/XZJG/qhK0SRUZM2Igbk10fZzCUki4yQWvNSdzdliS5SUi/gcBSSmjmyfaj5Eei
4cN2EwqJSxlSk69PnBk8BXcZ1UTuzA2Wyw+OOjwnSdz2klpIGdRh/7yfUHMpvkVb
PxH6MrZ8B+at6A3lgDH/hIPml1btoV62IQbtxbt2muThh00Oea/mkomkatZYnObs
bzPOdV5Ly4/M/TOlJPAkJKIXJAtQs24RMgHGO5RQHL6N4TzI+NesyRogn26QeEvd
R4sKLR9kXBxT4jhGFZogiHBAmsHVOjWaM8LHgDl6g5ec0Rk0xbKCAAwgKFnCfAHs
NZq3oSO2oHyAqRCnxtxQ1l5wiKtsBnokDMethjDZGi3lNzJVwTrgurfPAF/9oQNV
FaLlROez6OVN4LqqwiMWlk6Pzg98Yc96q/35Iq4DEELnPwHWYb2IQoiRNHquI1xW
bgyOaOvfFRWGBnhVYndYWl202L9B09BtEhKuh4pmJfEYht5aR0xMrhGdqeCOW5O6
zi6lMqXUbfPH27WZYKg8gjvSduGD2ecekBN41f5fBbOQx93VJDbkTYOKWg7e9Pif
eatZi5n2ibsiBhYm3mDU/yzmTuXBM5dOaW9X+RXA5QK3YPbxeEaC0SpdkVkEuP6r
qr/WMxA3rdqsy4elsoQm8wGhZavgexBbcNK11BlOpO4QTHOIbdAC4YEypetxW9pi
QYfqX4gFbLng3v3lWudzQvxDYyrxTgPjyIFUpcGJMOQ5oMoGjj/aSJYZGBajQyVA
/ArtG7SAaNd3SfhAgHINAQHCNx94I0TtgrByTBzdoC2hB0Sn0Q5Lh9Rrjn6WlDj7
ir+WzJhuGi4Tn1eAqfJGW7fJU8eoGs9O4kfGfGt7lLmeCiP6ZLcMYh85ctwefQIK
X9Ahpnq2yuG1VHsFJkiD1WIxPH7y+aBN/yqJdpFF6u7m+Cd2B3iQO0QYtDKPXXF5
Z17e4J+DuEXWIiN3OpGlouqU01vxz6E1LkvSizi3dTNhbIvyQ+GTmtR1lsD4Zg9q
2yDzZkImsd7IO0UaJMzlnWza/PKb6LyJ/s0pnprjMleGK53mEoNa+GwzHv5ZYKom
zZ8NCMWWo1k+oMBMOFHZ20AUczlpOo5zB07POa/53s+67cW0slTpsj1qIx2qq0Eu
ygGzbPIXlkFCQ2xStI6YbQa54zW2tvkiFmqUiDpD5AATVFefTUYiLaG0s84fexct
bxSoFfe5wJxDn2awjsHO0RtWobb8ositkZkYn/xB62r11T0+e6FoPuQZ37K4ZUZJ
mciPJR4dp1ZdOauIHOCmlvwo3Ub45sia+CYWEyOfaoe70O6+ICQxhN7OBgrcpY3j
DEfUhpHtA31IIgErFYrWvJbPMp3LPREi7tFdoUP+GjTfGA0p++qi1dqfk8UnSvxu
xw5CAtT8D9m8w9qUD50zB9p0LtkuFkaJkYJ3BtHswkPJUmo0xl47fJMXuE4SF7B+
7nJdK/wSx3fzc6+oisZqTMQecZGx3s988IRcw1ZDQ0nTZPphOUiXklSmw5nyQKwY
un5WxUITDAPHYE+mjD3RXU6ewvG6NLTOLYUBLAOWAVuU6q7NLiR0PHP1Bv9nVGRg
Z2L3zrFcVUkImege09SN2WCcgAXeXDye/508tU6pd4NTaNa4G7P9ApG8OhwZYTg9
3/91xqamT1MZ2VMUpoOLR1KRQ//Mo8a5+yN1byI+xvd9GzqlGCinx5fKtLViqgmn
3bVjAzUv8E56jKPsEIWYe46hIEjp2d42p3ocYOARJGo4Ww1eQeWd7eMVszdcNBVm
WskBIRdJ4A6B4u/aqMIrxTDO0EOJKRBbZXrUR89iB1sYOE3CkpOsMC1j6JO76tmI
t8i6pfc02F1xzSrRLYt6PJI6dXhVPmnz9Ko8auf1drUY7p5XmXXT6U6Lx1EWnumz
RpVbbca/OVFO2/GNciqopYfXvxIhx+NKzU7Q8h7I0en9phdDNp87ThEGJXgIIWr7
uyql8PUqfcVVsdCs/P+lD1yJ9OvZsvWEkenv50HEgk3RqCqeBP3PaMv70RYR9ibL
53N8aXq7Md5w9R32BigsOp54Xet4aAtg7yW0OAQEFbCnQVI4nVVtugf6JcuqaXvW
3aPvGbCPfT4Vt1DTiM2ZsOoSLCHThN4weXr6rtmLGsM5Klm4imkvSEz1Q/rNohkP
MHdTtWtcvjEn3GWEUPzpLvVgLy4SQ/qPttUlEP9ETvAdv9iIKr9UsftgARpcv+3N
JiRPuzm+POP+TCF7CVB7Je65h9PCBI/33q4QjPTljNsJk8bFOpN1Hrm7+xMJ4z9k
foJPkwPpKlxcR/2rcLuCkNV9cAMude2ghNN1RoNlC/cQEDHm/eOnvaf7f2ube9J8
6pHMelbxKqTvkEYa5RUxmCdWwHDjuM+UMwGNuj/uB/+D0v6HpyHlX03oPLFYk2+e
TWu8P9nIVvxpivMqsMaoTSEl+e1QoRovnWIm1NxRHvoIxPyAFwXgiVMhTHlO3/eA
DgHHfI9V9F9nqLNf7lXq4oee7GbbrC7yBDvzLI+n3mddeBONL7RSRMKN2up//9XJ
4Du86QjwLe0jMmL35IyKtnuZ4JTgtICRSVM6XfZaDEiz45WjWk3OV8O/0tO700M7
XOAG9mh1jIj3uXpBmRDWPUF3g3pCrAO2Jf5cEiThcKEbQNkIvIMnaKwK+b4OwH2v
o+N+kIPjfFsS6mrrh7ZSGHePUrpair7fMN/Yp6o4QLJoKZD4S/0HkgxGTbeN/N0s
hUfBXDyuE2B6m5cNo5Q3yOOkad1q9Rz6Ur861Scy1X7tDYQFFC5VUYk9hRrb3dbu
mUNsjuUSC9ubQp9Y0hyazKIv+HhnN7Yhs6suJzBfLAkwzuUkB+udQv+9DwuDBNR3
HtOic+RndV41P6OPRO7wKO9dDVH6Tci0VtL2ZZVxVNvV75esH2g5F7+jZO0bDluI
nKhgOe1FLsW2s/dU0hwtvsNccJZni37q7Znkq1UuQWwn64Ik7PKwTXzNep6lCLh/
Vujqy5F7nXzf+uzwFsgu8/mVTi7bb+s71xzPY8JdDhE+DkDA9n9q50P5nL596uhq
hevtI1o/bcvZ/wTu3Sg6yA3SuImmLXD7IFMN4hj4sbzivoqVFXpYTsV2cbBzd2+L
MZe5+cTO/FaPVFLylmzCoB/EcSFSkynZ/CFiwFUeRAyPQmIxvgdvKJwJapZLX/oZ
UfTWVRaWBpoF6Rp001tNuDoKfYfmP9oWTouWFBMCvgSw1QkkXL1J9ORHVn50vNT4
1hXFoiWI5zTKlHhZYKwmsR+OHAWtIFxZFWhE79ZcdOvj8wQ4N97DR2MwTHa+XHYJ
rUMydZj5sLiQ9luBBsEKMQtoR575kh0x/fWq4MYnSm78R4wHeQQzD8bL8c8tiPas
s1uE0DUc7Wu4BZmBmAKHPNlp5lP7mS7OEiog9U2of/t6EPkpsGVJYwHBqcoGgWam
o/CJFYcZxUSWoTbn6Hd+7olBF8SfsFNghvHCpsQ0yvzh501O/2hh+7E/7tZhmOfn
vLzPiTGLUg3lJATZ7SC9PaRdnGUMgMPLoJTMDdqaofagxVtOONPz9mzHo6jAzRBl
IkHIkHAaycElV3vkTUn4Dp4aPCcsxV5+IIhwDUSjyMr2odfVSnuGGzO4czChaFsg
kqirmw63O9Q00SaPPq26vC/b1vyIg7xvto/afE3W8OrnwB2fHIIfooLQJPvI14LR
I2HrsnzVS+ua3wgEiOtbTT8J90iHq6OxuUAMuNMexaButCagm3dXg+zpxvkVgJDt
KB4Z3rYBrKxW78MIIklWu4j1btn2/xArkYNZKhOmyKYOd7dBMap5NC97zauWTwi9
iM1ydBcBbWbj+EhRwOCZmaiqXLIaEvsLo82vm/skWie4Lf1refsMNpgm2DjvMzn4
P+Ey2vvMb6MF8KX3srwFcziZiKwxk7ATAm0t95Eg//uk55Lo4M0NuOWwIiy1+wNd
hMRWMI/pPmAiYrrzglor/rnbB3vPg8uF4xB8qwqq/1big2m3gseeEmrl4T4tEp5s
+2NzTfxaLzRFdbLUAtPvGcriFE13XZ5Yur3UUOJiq/oOEJbtYN4VwzYueNY529cG
YZrTWTa2gUJ+XRHs9jD88n1J+yUzj4K212JyFzEiQ2P1WHGKNm9IGOZ6ZjGeaUXr
u4JM96pE0l7smqhCSzM3TF6c/xvVt8lM6yhCwZ8xQFV0ygR4rJeV8pWrXSvcDpxS
rmIXOkR15acX2+25HqNaiFzzef9HYE3BS0AMg7UkepIGH2Jc5MwbNuTlOjqD8nDw
6uOG0pjMep2BRY9PaD5mXdA83j0MrUqgPAz+/mtRVxEC2J5yBcSsot92JMklMQHc
h3rM0RiUrSFAG0zXb5222h+exqeUSF5lkP8yAJJLcD5e5vtN+aEDZFYcWgdQwXpq
lluW5H7t6BnRcPW+9p+s7M/oL93HNmB+QWi+xu3cngPAyQL/OhDLc+s8gNJye7ad
mFnOKjOyImqNQ6q82JRrqp63Ze1RZEZw/gM8jIbS2OS8eKrj1IzV6HqefEjGIeFu
ZahWAu+aU0024yJIm801+3qIY+V9kEO3tCa/mN4840PPUoS8ytFab+tToff7RDsW
fJJhUr2LhwBX7VGmnDIQe7WcoQYpqvBwjL6B7I7DU2tYKsZ1l6R3z8btCenwBXnd
sTtoJp9d7JkhTQrhx9nUXG9IWWrgCXc7vDr/ndHk8NiD1GAsDDNd0NiraDTeG6mY
q8jY9fR5REIs08/cOYYnXG9+eOqZSk56rIAfrT+kxhKqvy4HRSCz/WPqDZL4nzrY
cLvFRUpNi0BI1RFuOugrdPrTnqE1kypIMU9D88r8aJh6wLGVRslXq/mGekumjA+L
708GRW+hivpsn38LBZxkXgb6EK1udFCH/vszXFvfaco2lvT/fZw+e7zg9kHSVwKl
C4SAo7/IEHqH2VISGi/gEsJ6glbCHEhtklwnrja4hmSC97yDcFdNu3L9ZlMZ1uZF
69h7qbzB2HHxYUX55G+0m7nN4xL1MObljDFearumE9YPM8dn7o8kBELsaMIAaaZZ
sSR3uwumYZopfU45UwNyPP3l34+AG0MCH2kZLVHKcDTnjlkyHfPcKhj3GbPDiuc/
duW8I6jk+dagee6UexodCKQjc+pQALoOyJt/lONV8oiY1CNNzzw9o23qcgxaen8z
z/3bKff+FuCc93JxPweuimzJpl9+VfBvRUsWZ8cYWRPiNcS++Tuj0hDHkRRwj8jy
RJBowMPfCpocp93+CZVAapO8uTg/+5xXUQsJXXyDE+5G/HKwKyHYnTZM0ldAKheD
rL3r1hahMGo1CUP05L+5QcHAUXa6mUxxlozh1aExmEBAAAkYd+fqB1aGb0+micX5
eVel4pbHYPABdQEmRf561J2jRr9z0iO3frPvKhdPalwJBXkmeK7b+/gVjXfy7m8x
7RXibn1RL3qjoM3OpwT+J73HrL3pHdPUpbEoUUmjojgGq/yoP0j93/mHmGTzVOSU
Mw6GmLb4mKEbUtz2aeRyIatMpX8UXwcURC0BAqNt+FbqXa1kF2oeKBxSMqNMNoor
mAog0xhn0wDiGL86KFQ//Z7PVj8STyckYhVLeMWaLSjYxW8gTquZC0PTEGZFhSuT
JGvCmdpIAqtNjrZO2H/LSwBJ1aeszz1qoqIn0h94CLD0/Mw2/+d8xFIuKYOhfJXp
hYb9s1z/mD8ltjxO6G+5OtHnDvAEczSHVLioblVWsKT8PGtuP85vVKZ4oc6vuTzy
i5ySnZo5Wt1XoYmb23T2zaD4P9+2b1lNqxki2ho4rEC9RWYdTd2Q3M2ojmwbDhOu
6nS4Hq3/lAHxHN/N9jlJJc1CbhASXy6w5Q6OiEoeY0xOiV9kHy3Bgp0XPGiQe+XL
RgaINkMBVlgGe7hkbyO77unNWJqdjJ9PMllhxV+qtPgwR/0ZSgOsU/v4C37lm26F
FjqV6op8wB0Upxpfd0pVgyzZOqRdenihER2P5s7K7j3ZGyzDNAYEf9jTLm/sFFnr
NonTkf7nF+6les92hpa/muRe0c8lxzvto6PVRzwrj77m7LqvA7Zd83gWk+XkZ4ky
R2Jksl+rCdm+Dnrup8m0u7zQRvAuLeYBtozxI50huJZoVGyaZiTuT5ON+R6GAimR
Gzhna566EM51SmAP+qNv89M0f5D18lNecheYH8imYybUlEJZvHh/+RGFEAk9i8Zw
bWSL/ViGx57343gGUHDlXGWEBoFh0emfxZDBgK/H1hbItjGkb6gfXuDg00ROZSWP
oXP6Um9TUGTPdkuNlsgwZJGmWKQ+DWwCg5zXjegPCPWm6I26XCrKFZg1m47cGTvD
84vBIuICK+aAEljXwGaKUK/HnFUW68qiTbmdr8XSZPXDjJTE7wJ41y4RHHgrm3fI
bw8q46PSCYhW68y5pklECoDnPIf8fkjhYjzHuKO8oYfcaaDOwW8EYWiqOTpGgBLS
rTiMSgJncmYWabX33prDxU8QeyXoTV7DRZu+3HB5i1c1R1xOmoO3ZjmAbZFJVocM
vGJdeDVt+0xpxTNQCVtyAPS9y0G67YplBkha8n43Qrhv8VDBP0ei5+74OPN4cchm
VZTXhW8V4cgXOPgybbM8P8byfnp5EpOxUkikNInW6mY7lQDJ5k+/MiAAqK6C3diR
l/xnf7FrzSakr7z1eM+Cb6OLRvYyrLeeabd6FrFgY1mTYy3gxqAm8YXC0n6EDE4K
XKNPyW9qCmwBypuq5W2uEEmaNOCWKVHxDhrGU+dTE3Q9w7sGH6KH/u8tKlsPxQJ/
y93r2m6chgZH3swpkKCuh3Xjs8Gmllzq6A56ZnXtWal+ogmeAeL214oX2dlfiRia
DWLxx8a0XzowHW23q/SWWAPw7c686FLwWFAmfzEnN0zOunFOPlqo7Zjd+nEN/MmN
QRAy/f0rgreoA9fatO4zfBWhCqeup9OQBdo431eqJ+DS3zvR/CW9Q+35V/VRlLjl
Foi7/Kf+QU17syTmtS1BIRAchMwLvPEFktebW9RRaIbSxhMtNA868NSI2Ai6bZvI
8VSr6BhdpB6iAMfbq/YIt/D3mF5/ikvPRprXKdAKSXaAqcBKIjrQwy9jbCh9qjfi
86t1K2JprRxi41Dc/TQGvq7vHYgFq4qiKQVS+x9uwzD90ustr7qZagbktWcIPPdn
bXoFxCL4hzhf6saB2kuXb7mhXTxqwfPntuF3r6rftaj7DNZiuJe1NgwyCLv7+8Qt
qhXxrr9FD1sEHQlm8PaRSUPSx0lrOduRLa8lCfoVbk2fmCtNnaBaP4kaK7p9bIPS
hIfEptWZoo/5vgTmws9Mi81LvrgQTk6+HMWDOUnr0B8buNUb3VD9FarVHzN9Dh3h
x9Ehy+V3ARpqTAlBAYolLeLrfttfXWyHARw2w6QTTg/hfXgaZIqXHx1c0P1JKVi5
nZJGP1aDetjGqB2HA7tcQey+SkIGanIH/56z/vO5zi1arqbQOI/Tf8CkW/yH9Nth
iyXMLpM/zwdYTkWVyYYmObptHqBl8GcUIJopGXqwbA4yvQbf0NvfGbm2QS2AWLGk
2UXbDw4glGY2IOHCzGul3kk5SID1RvjFNd/HYfuBtf4jeCiBdo1fgjXQoxEHBuX8
zcDbXncHLtPcHcCXkEPN+K0sp3NtxebD+MSCGTErc5oRFi6H2iwyydTxZO8ORY4r
3iuAuemvqs2qDN7PUEFrKs7SOd7WQbC5EfrTWDb3Dvm6PzaKW51+nSHBDCGO5b19
JJ7D0rzYdJkseAXsGYz7JtZ/6gfHMxwHGbJhJfLk9GCE/TZCWpR2pv8ujIdZSEeU
4ZJMOwjG3nizZFY5z2pki05hXEwoVepKlU8+M0KIdGcV70qipnpqmP955SU1qUaL
Yj4AQ6rTLo6NdU2IANYQHXfMuv9F1oAyMYC6LuemPGM//xDr5NHzTZy5O6nAqexp
5a3TQXrx/Lt5xJIxBAtpetMxVTR6P60NTiHYnv3vokd99vk+OXvyupn4D7xV5fpG
MzAMt3aQ++etbMaTQ/fJP4xtx5OuQ3Mmu+xbHq8h9lB+2E/SoYNnZCLeql+w1TYw
xLutxPScJK59QBAGM0KvlL0bZ+PHQAsaXORPgxNwdkTOtl+pZFHs1XbP9TR51R2M
QU4a0Aq8WvXJ+YXVe3j4XWY/b2nH0ksXsJyE70os1Duf3lsyXPjoAVYcSgRdEfmz
XIFMCunCOAXu2VHuA/nu3JRM6s50fN4UWRuqvet8GBsIfUFIoziswgoimHL8fPZW
egSA8ujZMUue+gwz6uGaFMtvWQh1gql6yOSiUvlPF0bewOzDMRD8ADizy6MS5Pli
oTckF2pAcIbKxZ8N6Db/8lh9/vIuD5O6Yg7ELMqzIJDbjN0stNhcNVFmblUrXBsn
7tDHDrjp79e5IWlpXP3YAEdKdvJRh7A1h1UDbOJz8bOPE+QaICdVr5UAkuxg/7KZ
8PnoaT9pS0d62BlSlB0SULZLFQb8xsQNjo5C61S9jDOX6w3vbBvSYuP3gMORJZxs
8+U3ldF9HuIBwCr6apuIkunpqgFNevrYs+Gsm0MpuAqoGa/XVeRlR4rMRS4lIzYO
klMp12kbJtmT72BBGOVdou8DEQTuyf72YC54OSDBYEvgUBwa/6d2tklKDGZS6LvO
E7J/phkhAsxulVCv1nRIo1m+JMxJfXmOKUi2aSwHkGAlP0sovW2O9l1uJV8wH/XY
dS1J/Dow7LNwqlBAccDXNbaLGo2Xum9zFC8EZD9g3gD6ZmnhCTmTpeBmBQSbpDcw
eH4bjFlyiedbm79aZrzYhOXVqaTJpI5dbBXAmSIugT/2NbUfAOiES6ClXE0fViXQ
oxnw5YbFbSU0ZCIl2kTyjxyAhS0Q3ojEyVuFpefSNJiO/lx1D4YAA8uOCvE8GhTV
bx5fYZDT31cVvZii6y5mvRgbxm1C+LCqHGolR+jYsCYUjJ01AcuWl5/RugAlX/Nr
drzbevvU0pKl/HD22mfykuR8bQrS9xZ/Ozbfz/vhUxjqdzvGQmgZ2Kv/DpYy5gQP
f26tW4tO0eBwHWXngCgxhqv751gAfdUuc2U8JjCqrI5DzWLbvy5U0OsSJ4awm56U
LdRT8vLrK7OQtwYSiZaqOPN1FNbhA6gf1aH7VQZ1U4rUOmW99lXEexGNuO6jE2fU
+43g/eEpwXEfVknXlyae562rQM2SxEA8A2XvLxtj5K1PCx8wmsyknn71vqmaW06I
ZsYnMXVoG7Unt4bmVd4slXZ4dvLcJC82ipQ601cEVIMlxKukAKzk5GDuF67HW8Pp
Xew+Bm0CN0qPjWD/HjHyRADyuYhP6g/AEzF3k4oYQPMnO1ieCqurZbBcNu3VJnJp
Upf47+7a4sVfBz0r9vBBmFVEAKBLi7doo5DV36A8AYyos02gtBRNeoQWwRic13cZ
YrO6fpddGGJb1knBex2mZFtljqeXTpKFTU2fs11QOpOdHxCCEpUWpHaAgi3UsJpC
yt9lXnrfubA+Q1lCVPQ2M+RS1miJsoNWDEgTUgAMydUNK0edUgCtL6MdbViy5a58
nxgnjKqxxPpWKd7YV9bi6iUC7Exu+MZSyapoA46I4pPPAHKrQVpnJmLaIZptVqox
q1CTmQ3MIYtylZcX8rRW5PTuU2QBc1i3xwF8TRUO/TQrFZJF4e84zIV8O9NGCLC6
tsWSLG3SubOY6rOyVAVjfsArutfWb7d8ZA2sNv6KmQW+RFproyjm/yM6Xa8guPNw
7SUedi7W4Tf1T/j6IzpoXRDk3XcG1fBw/8SLV5VKIjYxPAUmzbVASofFAZjNgM8s
CUFdtz8kSsebSbAMbZ44LUcuynneCabK1n8+SHFf3GoId7Zg1KKHqDwdOMTc2FWa
QmIhpZJus9c8cVo+vLBslsHVf4Cn0gOc0yM4i6q1U9sWcGa1j9F1UzPPZRANO8//
AX0vEtZaoNG7aaeS21nB5J5aIdxyJ1r971mx8fcsVK+d8zCf1p16TczT3v1pnkQ9
+q8PkIyA0h5xb4R3fRzlwSj+ytPAETTa1QEQaQ0XIlL5CR6y4Sa3or8z6i1oornl
7DgFI20zRjSrVE+DsiKjin87doPvX4ONcU/7bEHWWpxFBCC5QR2e8/AeKL010MOz
6u7ItnwrjEb8SR1pe/ft9tgnzF/Rzj8nVpy51GrPrchbwuEMaH1SmzfqjetmGrC2
n86hrpwHvF9i5wO2qf5wsFQdEuDeyaUl6FLUlzkQW7mVgCm5kgq9VBIeBUzb4RwA
3KJuiarVrHlNYVMuYpc5nKJhQW/frSfNQshCS8Zai/QOAqqSnHonnwwo4Oh/IAFg
y0mHrScNn6CF1+2etA5B7ZIXFKrwNcCM866guaA1LDTZNDf3qqMmLbpli9vSC9bk
2QGsxeQfVk6i+gAR6w3TuG8nz46eUKydfKfAJRo09VIjxPDTL6siUoGT6DP/lqNp
q1UCssvr9RZELZU/oCg/G/nCMODyGPpZId/LE9w9l481j5hG3xwX77aBKISzH7bm
w71sn38EP11dFFqoZrh0RCttMO4gdHLHpPo4HIT/xxvCA8gtpQdSlcClf9yW/c5A
o58VEw6EkcPFTX67LqC8gFJopqSjI+FMih5sIdZ6oXcfnF0/D+98V07BrSYSnl10
IOKt/HZePZpwAiE3fsI85T2NYCoyg4tPlRVl6GVxQipUrx7i3EpuvQV3BxPkRZnO
0EdR2Ur3LAQtHVbDoSy8E0IJGG+Pi3/u04Q6Gf1usru/5R2o0l9fmTJaqkbqJnsU
Xao5o/ij9XyLcCREWxOs81qWPt70OeG8LLRMLXatNG79t0GebaZUahAbM/8UbDH8
Vm9oGbl68iwbVDKdcsgROp1JZssAa3Kp3NfaNTO1a3EpEDRnJKslEcwBcu4z0bhe
FVDdK4uz+4N9T3fDPfz3qbASTjuyWnFKA69hGY2026xJRtg1pcd/jGZDZpM8eTo6
xNaXk6tizWK5pGX2r3a+sYGy6cmEv4dIUrFt2qYuGPeO5gaRCUk/4hMuqoCEqEaE
X/bJ+kbmU2ODBPqE1k4yXe7v/IPDuQ1h0GeJn7SbKKuJLGxAG6xueg9xTj+1ddsU
BezOCZrAT0zAfQs1dxXoQKJs+PuV27TO+rqynGVleInrwTUS9tFM7xl3/VpOSlxi
R7HEqUPACbNFUbk9lXEhmkhsarmsCYnSE3vvWErilIlr9mfxwZs6Ex0hlVNNu6Dz
R1LT/aWwXQfkH4rplSQw8gakrl/ftqUhx4ZXFhRlGz+RuQmg7Eq5e+5KAn4wu/OJ
nXIZCIyIqEx5mT/zKRmaHftuFWfuKpjBvbUDR3ja8fnTFZ1VXJY4Za8TasvIwRtD
/2Iw0iviKCtbXWEKQdGJvGvD5N6cuT3s9xMJMeX90ltBTdcWxDP1H18WyRhdwpki
oMT98a2wTWOAzHXeorJjXj2uyVSTDiCmRO88nzDzFOiLh4XzitDXGs5QLiH7fgNe
NOCf35fuMZhyJc2WFHqMKe/iGCLxGvGbBWkV5d/ED4YC41dO5Nvjqj9R13ewo2DO
Pys74ESGmfcZLatH0A54ykqsHvttdPYQu0R7nSUIoNyKGGiUTysz+zGVxi+RUL/8
QrkmOmK79l1sos/i/N+ULV4IwA5oVveMugui4PEVhioaVKpe7s8UvgaWrFhGVkao
5bTT49v1TseUFmi5BXBtuuUzgV7S+lclMA2S9vGvFtpQaO8wA4YPD3Z5GcquGtQ8
5OWvbHv4fuV0wO/5fm7N+b6ZrEYfZNd0y+EL6vJ5+bSTJS5xq3oNqX/q8lAz5AbE
g+zm69hFnRGjVXic76aQ72wUqLemW4QLi5B9+7Hfm9EplVWe7SgYl2XaiQdjJIoL
y030+zga7MUJilpnhi0H+pbmwN+1OZQlM7TJ1puUcXChTars6IJxO7aN6eBkLzBm
ueB6Nr8spNJL6vhfTE/Jf+/sKvfw4Jo2r/c5dPbSGl7n3fpfH+gpex0S1xZZuHvO
v9S8LxBp0BIP4hGKk190J9lin2QgpumVZdH7xhTiCRrMMZGQnXbRTsoMKYz+R/ji
qLKp5cWDAqh0koK6c+fSALvtF9rJTYS2cE+PzYZ51Be4eKkW7JKTh808kARo2UJI
ZErY+FdeKA2rnE8BBD68/X5S4f2LU64QeIoVjoKhh0ojmiMaRBJDXCIKUBnBB3Bd
xs/cqtMrt8gWmUwVciKrOO4X8JAx9sqXZ7YtPJFtVgnesJ2WPmGGUjFf8wTvO6b4
w82wMQqHE1Ip4wqpU5wu9HnmcoQZesDbJUMes4rI+Vo4eltUrqR1rIoeJBZHd36G
9tK2d7cRLiceuW1nOGqd1z9yIxLn892zNqAw98Zx8OS2awkhuDIUc09qzuNN3qh5
pkCWrd/jUvQzALrc1i/l6cT0F5zWPCTCfYrKnu8AjgKPxjoxX1dYkh4Cf0j/MWVA
Q145Evn8bCTOc9ivojM3zmtYb3wNwKnq8PrenE4SDqkHA/Ib3LjdCWbX7QOhuU0P
QzyPu4aNt3CvHxK7BgJYHh+EfSATyr79Bg1IPJeCBp9RYywdQtwYouhan1ONUXL9
JL506w65bMh96MYKq6M/QJDrsHpHm++6S6WV0dGxQLuzTB00zwzb+QbOy+L3DMEA
HHCL1qnKFhmguWutDgnWXRXWHHtYHRg+f/Mt7K80W1obpwGdWiWqWgiKZ7ha8dIZ
KMTFmyz0+4VgDU70+sd/qLXQCWamsCiBsJu1tPBRMVPRAEmTyyLt/zOv/cNcALZS
eIOaYaI8K5BvQsmwZTpFpCZLiEJYyHYYCDheupnCTSenq076irDDshPwdwoFcEam
it1ahnnPLxe55TgDffzRJeIlLvxlNd2/F9DJUNSoXSH5nlcIA8Vthh3wndyn9dJS
lSs/jPWUz245zqiDwYVdsUKFuUXDfkK6glw3g4M59y16apff6d6kLi7aVe9W6X9G
2Y/zd2W1Vim0/CGx0rgVslJEWwOBAGrmhW8Mj9qhLcoMl2HjHYn+wcdBhkvRI4qy
vq7LRRG/jPxf2CrxPv6dcFmhxP5Zf2OFXh+2drQaA/PBbkVPkA2zubdKtp1StE5n
VDtixoAvdzLsEw2ZmdfEi3W/A6a1au0arwqgNPrc2EvZuMia5OXR85LixRZUyFZb
SjMikhZF+tdQkRPVnUK98Jxa7YgOTuupBKUVl7bsG3I5rp04mD8T5RpYwNfxpAs1
QVoLerLIcIXxKDheuv2VGwUPjb61koY49KmD+isR6ukjH80n/dJGs1OA8oG4XSvj
ApWSUbuM3/XjkAjDBvnG9jG4rM6n/wj3figt126LxfdVRBgyW6WFDQAL1zvzKET2
2yxFW5hMYK/x2xM8EeojqH9IY9p142EBePL8IVTB6FIqug3tJLSPkubOm9UIMIhw
PD6ywSwSiCzVAkoKX+otU7RRM8h1GWUO6OC5mzG1CEWLd1YmjtoVACPx3HFxZ7SN
dyxgIKspZIbFOiGyDxWxXwe/mvWDiBBkZunh6YieNWJPPFhQQrSVmFUHOzhnsuTj
wZ8quVizECUfN80xj7c9kJ3D8geurGHyoXPblg5Fk9N08wKTmlnGQX1pTPgD3Qit
/sx3IlcCwwWE5V2BhAR9XS/HNACNXXW8LkY76/EPnWk8SmDLSd2AjKiilVlc5A7e
5+yTh9qjupGMnSnDfewTptvH/tFsBP6vM/wUc9vbPZ38LNH9f4ztPWaQbIH2uYcy
6lhHocYCT2QrW8ceoGLKtY/qE3UTbDYZ3YL5YrsM6AiNt41KbDrE4z33ZjZv8YEL
eBSGS5rZRvdsua9fW85Ko2G02p/HQr2+Lb83sWHjMaxd6CwA5WAFo/ORrnH4BDYE
CVzrNtHzC9ktbqUlJiFa/5cDmivN2qkkP24bakUWFJcHbja41dfwdnu8woB5vRCE
qOwauqv9KYcLVvHm6iE9osfxVrPTYwbIZPEVvRmLgRxopVp/7bAsNWdLHPvt+RMz
HQwjuv3+tJT9lKhKTEH0MwuAX6BpuCSEJQgpNnhtxmJ7c/DEdvSSwYKEkSMXjXbG
6MOe32Ym+Pb+8tVbG0FcxsU+gsNjgQ1bXCNA4HSlDhiVDUhwQKw4cGIkrjievU3X
8usAG+pyezT1n5AW7RDESyIhG4aqjd1B/MGeAXpwuo1Yds67hfnt9RARqtdB7yLi
qJrDepBcsbSf8P5C4g4X4c5YDksy2pnfTiQEa1O19vil3l3M5N6YqlR1ROJgW7aa
L/1kxIdsJoypfb7wANTiVzXVI/t7UA0zN9OXKgCTiMWeHlX0AgvAAW6F1rxPXNz8
eTbv4FvV2CvrHFPdFyYFOyC0SMZCSvah9C/UfCbSgkgQoRzh+ZbOvc+7NVijeQOc
wPxxlvl/KvAeO7yB2JVlefce97lebPdfL6lgr7eyb4q2736oZSPD6AGsdlkuBMCX
MO+tAW95lSWwW2TQ65EgClgH2UF4In/xdb+W8niCrsoVOTo7rs28cdXZZ3Nipls7
ST/7YICm/gVFg2e7Pg7NYZD8qShByUxjvHQemstrTaQq4Bkss4uYBj3iPVB11D0L
WeRVdfSfHouieGXIamVX6hU0G53jyR28ZpbCUw0Y1OzQxBukcfS/5kN0I4czZ+eV
ML0Kv2XKcnzrHI50huMm5E65EG9rr/4hj422MNEZMv7+xHP92Id60kHQKS2BPIwC
7kv8D9ctseFwarZuQDqYekjf1VkMN2deQDvtjtFZh9v5Jfktlx07w4GU8FGiubzQ
j3sfom93yxbBuBceSHOzTM9qxWZdrb87nbzWb7qoEc/Hksim/jiLS5SFCPyuVrVS
CPxpv0Fw/Vs7rcyBHCAx6t4yYyJlh27mIB/bKbOH93o3Go8M8kayhOXFbYDSltqQ
JduVp4y/2+w7nONGs6y5MkcpV75w9Np+k/ezCBZFU3Ff8KWbUtJ72+qd5pKNhCiU
g/YIGOzZCEskFkEPUyei87sWz5RUkpFuc1N0K7pkH1VHHJhqXeF+NJOdvCczTas1
wR3Z8SBvF7R9IQ+rNxmW7Zy9kzGgFwOKNKjWE2LmTm5hUDeRBLDzetwrHnsVlipb
+99qxCZ/BwmbrthSpnyCMtfC3cFx17s7jS7Lj1542AWPLhBKlXm4vjKI5/rfMxxm
B1pYVcCAUCZfYB4VDOcJaBH0WmInkHtnAVSI0MnQPLvoZhbqhfqyu0p5JNnwjO6O
9gLIsiAwcybzy3jLafr4FrQ92gflAPtWaelvD8/X5uyNaHZjfmXH7mEhzoGnwoeM
4Nax8HMtfor/OUvnsTK6ZRKakjBS/AA2tjsIBkfjzxeEG/LaDBK4v+3U3EzIGPdw
x+msHyWIsTlYT+wb3jGAnTbxsMl+fw6Dd5wnrU0E4rpwdikSzgsvOxUMyrVfjDTg
891ax3vBaSSx3Xw7KczlYbT2xGmvFp86+WGpaQe70ZfwQL00Np7OSxD3JaN012tf
cxkPu1IpANb7wgm/GlCRVne2/K0uKlWewSV1BofTmMQJLwpr8Ud9DEUVKaSZeh5/
gFIBtVylDwLrNnfGtG2nNj4zDZYOIt3/Bdw+2oyV51g86tPXrngHaLg9UQIE+njW
8SrNXR1jmPH0f6AioSF9tIdUsVfSs2XWrEE4mmGd3DERy6wRSSPzc6+QtrJN22xi
6JDZ3caagSAVyw9Jz0Sv4B8+Sjq0Mck2BdfQ7nq+aQgyG8OeqYS9SmkHjyW+y8/H
/7KUr9hnvSjnN/+phitFHRWCm0/OVtgelUzZQamZMIx3SaS4TxmTBPoqvYakvVb/
GMYZhGpaFbPPyoyAzmVb+gJJGjMbRbWvZdLmx+s633K02dMi8Cm74/YW77LOqDFb
C2z3gp0j8sf5CVZ/xNo1Me8Fzes0OWGYPWk8VRH7SCGCYv/B53WiBUZq8YI1QAQR
YZh5UfJQ7TO+47Yk3ttfG5jYxKRRoa9mWr4ANtk/J2pc4cjvDzeV9I3bOaraf2I1
MNpgwhFU+dkuvfSEnnhxq9Ei3RTKdl/L6QSq9jdw4ufGxtgzx0MPpsbbkJzwTe/2
I5/IQZs6MoynAKCczoGQTc9qr2kWTRwmhsb5WLW3b9PMQbhrXl6S/VFN6eSTKqCQ
9VEiNXB/jMIx13aaXTpuwEEviQa6lb99BhMyumbosqRgCz7ilZlNIlRz02GNFqks
Tx/xFTccJ0xNyT1YEb+xMY0E3fDYsQYfrIPX6f1lBcTfiSgU14xpQ9YCRXoyAfxi
bGN8Tcht87aVdcaRwLa38JHz5Vn+sbZ4Uap06/ws3U6drYjBe8yDlFE1spm/igRu
THpi+oueoa6Zv9rQIjV8kTByYXHhG74fFSwvf5NwfYC0FotTW2Q0ZdBRi9G2WRGW
4qIZBUFdflUXaerGWfKIlTms3YoK8I3vMjt9SVX84q/V0tITPBcme/MwMv8zF/Wp
szuu0PcKr/J3D7qVM6AQP0nMGNtth8Xok9fgMxCe3N51LVqm8z4UwNQ3boeZitfl
NYDAlRlJ1CknhGr1Mu2oHQZATOQ1Ps/gFA2V/Fr9WJK7uWyxcnl1zdSxwvVpI3KB
k7qzNKmJ3DcHDUGHbxc9suPJZ2YfqDtmdPJGHqWXqQB3buSoEZuRPC26NrcUvv1l
OinLddIZ3gdFfqg2InRqJtvORn5P8F6PEa5SlYK8jZ4DKRwjof7p2faVRMiGTyQy
z9IWOJhKWvnCW5Qs5kBBewrV3Ss7n693+jpDvD+8y3Q+LAwHNymDO+Jn4ON4DB5O
wlaec2ErCADlkUW5HkUy6Bs3v8pONs914Vm1yDjYlnvwgKN625Un8F9EXeBW8/VE
9rwwLAG5++ta1Ha0mFjBSpx8S9xxxI4xhYAfyPeIjxgPEUaTay0l92bmQxu9ZYC4
fvK/skJo95pjTS2E0jqNzGVkDBNJbh21KerG19BJYQgp5Cx71UwKCazlC2ctvI0G
/sGvCMBKWZCt834WWAoMtseBPeITVbFrhmLV/E6UAHCDa5/wbdzP3CB1A7JkTL5I
dbM+CpmNsmwJmlCtaqBsxrWTj3PwoDvYtGAXmLNb1ofu39DNgHX02FX1vxApqa0y
HMEUIFKKWaDf9Dqr7cWkxsu3YPBInUrZ+9rkmKREXUF330AfT6ZMzMhdagrRhcDD
7d5BLR48WHFB4geLwBovSY7gePndNJfTeof0J1VjzaOFadLbGhB9Y91frzBqwxUa
lRxjCF7BZ+IQe+sOm8Vf72NVSOa+hWIiNvcpNp+KDibhVSyyKHFWgBQjRjW3U//q
wbTbweYcytMWRR2vyjPBg3ybFbLg9fu6d0PJVecBD/brF+Pgou2Dg+DMKPA841VG
UvsKA0bf7KblSIksXuDXNw8RGvKrB8TA7Z+rLq745m0gNVnjo27cRsD7LUpqMk0T
rNQz05L1qUlACnWLMynhUrBnrTV0q9Jd5MEA4KHllbDAmdHHdfui2tRHvHkk4qAI
ja8tEDiQhq/xtnBHZkkEB6fGpAY3XWhkNrCfA9Mtqh9zUchxFALjXSe5UzhFG4lT
NbgUOrwHJBCuUlt+KLlVh7z9WkmJmUWSnkk8HMAYOH09k0u4tP9j/MMj+aCqUJx5
beKhLieTq0SY9pEb5psf5mGjUSE6UuZFmVrM3mE55XdIH4AJFh9LjFp5DkUXwf0M
Y9u1mQ95DY9jeit/KsJCdEGOvntxIScfx2JQBGjgqPWXiJ2RriToMvUWwSsMipzc
dm0wq+FLEFCvR7hVq9rJ5ihTxiPnKNv9Bzeh8ZjFp9nae6YnIuVaadDYi+ntTjpd
EIsE7ngYEOSZ28A/rhJNx505ZXfokhVzLJ4frZysi0v1Bz9vmfnwO2e51mpRzPTp
OrpD8DBQl/ATt3EUC20POJqRbqTdBoCCCDOb2Dyyo9Eqw/nc6k6fiiEpHfOUwm98
k6+zIUBT3iTgwTedKcEUirffS+7M1c9B/a3lCZI5WFRVeVUqChXSmgpE1+9NUKf2
y1Dg3KaLlr+oHpfRdC09yZUwc+lKfc1NHkCo42scD2AnjWRliKcpfQxNGbMjeVPZ
UGKxcVC6qCIxWKW1tWEroqd8tFkClSlAZCp4cpF9E5CaQS/S0rkw35Fe4rhYvDL8
FXCPihl60mG0+PrEygPea5xY6BK+tEKyiqLz/F0Nj8/lRrsiA1zhS3m2Y482D6Jf
BxStrlUvwlPQ3WtlKi5V3rUmbwiUWdNBtJ3FMlOlArjft3ieh3QVMQUchXunJfG0
L2bdg4Gi45WWSlycaiqduveh58pPBNkj//sDIpWI80leDyw2bJDSOV1slzVxI6Pf
H2kE+ErjmWgWytQRsKHReuuIyZC3ITDuyscfEq0zuPBcF67jJwIzwOi/H7jipzsb
vBu2TNnb6bBUxFjs2AUrgCveNlYlpS94Ol+Y0ZTvCBfyWXqMNc49+TUTVyGwXHtS
KCO8Lig223GXTPWE4250BeG5Hlj/9UocpI63vQqV2tj23OemSxrBdMUcsHHPLg0v
tNPk0TiqUFNcuz2pdTU8HAdWfhyWuEdkUknR80q/i56cm3FMOn7bF40qeAJ73IvU
84+mgz0ZcN7U2AlwJRXntN8debOHhsT+rCS4R90K/e6LtPTSzb6K3K61lzQXSp6w
puwut0D6V50inoESdZt/e2jYH8p4E4zkVwRdzNDS7nuVsenkVY+9ZQBkDiCWP0vi
7qGHK20Ug7KUyr8P55O5aCQd7ZRYHoeI54lKg25vXsbD4z44BYAO81ivQdBXFEhi
8m9ftEeJV6M0k05NfsEg0co86d5dH+IJFgCFl53aJxAwFJnJzfrzitzHQOtpwc2d
as/+AlZOGAqG16Xe9O9ROjo1DqEVehUJMx1XK3QoagUt+MMx2KW0GvcDSAGHZtLM
SHgt3O0/BloVfTIspAgPryx/rGnEJMFVksj3pG20Dh90tVqNnt5CjS4ocPoeweGj
vGbGAMS3yMxJDG+AoskZZ5inneBay2Rif2vmajpB47KDoVMZkSQNspm13oa8/9mv
zjoMIMnYdI+NJ9FDI2jbJcp9iBqlFgPccDOQtahovUXHA45bpOSsR1Ms0jcwXI1J
lMfWhCmAM56PK2x2lP7pz9i5hINfyZikw49ze+Rp0AIsiPc8s0P7aAunVLrpLZcX
uvm/JnYmUQTiwM7oeNZOpwaKn/Y7Yo6tNmqVISQiYCgVZnjo/endj3H8wisKDzhK
D+7kZ1KUDgb2c4xIaWnYV5IqBOhtddn37bJasW9IdW0yj/js5rc4KE2Yw/5LAG10
1Dw7GAgPXrWpIrWfdJC6kngLvlIBbPVUE3Fnr3xPmibei7uzi02t6Lp5zgDD3WtB
+bakTXC5Z4ZhRwI/ZTBp11R5QLu3m1jYNLpLNeqGj38s1iJPTRabk80Tr1EoISMx
Z02R0JZhZmdCnfjGzM1FeVbbj4CWUd1HLfoppHyq2cPqmOsR6RccU2nykph/HKgR
Ugb3MMKRTVBaCe/E9myzdk4lCGGkDkkzhDz0p0dRH44gORMGzorXeZak4dQFpcMM
KBgcAzocUWCgojHunbM+epN4nhn1wvi80lpwCJmZFV9tePHwtJrT2FjJWn3ObiVI
rSJhm9wtqPAuM3dO/Ub7z+m4t6ujkM1IS9JeALlwCKE5kuLURYHKzm3Uxnt+S2JC
wOC/nP7rYVtTSBV0t3auq8p++lVwtAH6y7FH/RiA+iu1ZxVns7M+9UUCuqaLJ9Fx
V4Tngz1E+f5rlZmcAahTYQBly7BbFQjm/pL87FSla4T/pqHtpb0pgx1L27UPm90s
6Hn7D/zxrnmSr9nJQfTL3Ye1/UoKJJakDsj2aFHaR81d0X8sCGVK+X0Ah+57e4rl
aTvTMUlcxQL/dd2YYZN3Rfc5uP6hB4ltoHTC1SkYY7EwM9TdndvZJtrlc0Naqffe
o+EzhzmTCl0rsIjd8GLSSWPRZL8mWxCiZ1J/h6ia2uvbnH9MdzEzn+EPFpFXPrS4
UMqVDdfDQ4zDipXZGQhrk5Y2XDlT8q9nOxsro0p0UGw2jFdXEyFDN4YoXyNPepIJ
PofsgLRM+nnG9rXdhv+h3s0wj00yUtQk7LQEPoin+JXPoMUiriQsHaB5IOIpOq3U
Nf0p22dNLvsmDGeuba/EQYvWhTiH3ayKNW+2T+LBzNVsyGpHBGObMfUzXTmD7KZZ
6+DsmPW2zQwVwJcELL4/DCX8j5FM3B4uSkd+/ysK7Rf32KE2pWbO75/lAygqUX89
xbP2RqIVHT3IkPwwOpQaaIdKlzqO131sYAV6oK+M7VkM3NGyeUvp7vai60Vxx2b7
47BPSeglmqQd6uuMi0cBWNLEiZ8LZ2kddsGSIGdVhDFPeDOLFJGyi1uhbf34M39v
L2nXs45tvqmZvqrMqF2kIH4PIxADLGrDuPDFM57svefIzbsc5gXroDbmFiSNlGU3
AxDH5Els0IP7dZns/KtbMKaP8LFdL3EVDllX+PE5hIHsXv1hXLE+gcVFVjezRaPv
T4uEW/ooie2Zd89OLoa7f2JS06sYd8xfbdDXJsVIYT0Lh+6673J7h3KpvRyT/Nzm
ZRqeD+9OBCVQpCqRwZbC+mD+snbhV7CUBqx+kZa+/JkX6IAWGrjwvooOtSPFiMPl
bouux9IzulZBUzdWfcCc+7qDLQX+0CjyLBdVzQ1z3HuG4jFJpC5ihdaC0C9hZhwo
t33Tn/ScAAiMXAjEutp078T96zJD5j29MrH1bIk19ZTkwsnabBKfBFpEvMaCHxqY
8/B3IPzc0uAM1BgUyWO2WuTweHzKiCH2pzhF7mgBg8HQ2OGPMmmRFl8WQg2E5Znb
+ft7HnjDZjJ6h6oTLiWhKvCOvY9FH6LwDLUW6gzqG6HTT2YI49pcEAWxByzdypTn
paZPTuju0scQuKTaJcAUqbFvOVG8PBhwGqhGlESebNGtTM5GHoCHM6FJJJSTlePt
WUydmBiwsXZFbt4/+ii+j6WkMV9Xye1kGYxqYsn92TmGMTAzNb2mdIsHvGxD7ltz
1NatUrOjFMQNMKfV3LGY2Z6JOYmWk8AWWNOLHzibaw4P2bjXXJyaY4F7WM50B4nF
8Hl45iotYYjJp2vNIyajfii25NA6RL8AIPdjDAmjHv4bvnhIkZlBHoiQ5qUklSlA
nR30Cm77BjbuAz652NnQwHv1VezHxahTZSkRFqtjNWZGGLPnzo1SOBDooqtZlhMW
r7OIKmI/2HQBET4DGGTw8YTmxLeSJrrOkA3TELdF2jYGTtovswniuWsShhc2V3K8
h64fHscXs/aEzLwtHhr+bhLmURCLIt4DmFkUiwv6sq/3oiAFOuRVMsnDGZiDAUVt
UJzItbLUcv2LczPPI/7xpP5qXoWtSQ28CX+31bbsw91BV2DBlf0f8rOmdeMNjIsF
pnEzGGZGTg04lbfYrGeX3I+zqyj7ge/R4J8b095H1G4TXSR+pF6SbgiyLB0+D/x+
W3Y8phQcFQQ06Wb5ug8lIafw55t1QtT6H/by74MMimvfgZyd7wI33L3aG4VjICUq
klXjmLt3cjrPrXkm76fVacMglReBO8AZi9El1IGdf7fpk4AfJclq25E+4Pixn8ri
camjAJzF/1syy3uLEY0A0X8ZkRdJC9fQPl84sencYxxyZIjA3qtEooVcfM0AJccw
17GHLedpApbnQ6dbxY5UNMpiAGsxIcQ2VvdXAOiRSYECR5bB75bofDOY6VJSIWEi
tSGszfCM9rO/JpaapS+jtxwLwmgY2KMdnZ4UyfkTZlOskqYSSO5PbT9dqJSzx0nu
P2k8GzLe58H1bLLobPYov34wxs98ZAslkW5OZ8kRvRlg0MherskTmf5ZbdUdDQj2
LUmGztX864adZ9+gWaRvpDQhTqGF6JGmR/xdA7SWg3FpTIXTyngpvcL8oCTEhIqt
bWIWSez6BlSKpOo/kvV2fTd4Gq/UElkgWisP/dakLdl6l7BaRVQyiVhRfr4wa06q
YNsoimQuZHB9t3I/vZZot2zZgJVkthgI1cDH2GZKtg3mu8ItshrDlaGcsRxhBidQ
KkTkArCEq+zEhZK3DDyhZwBDs7oCbrABYEFRj9iRnGXfP9NYXTPMTybBO1qFlcvj
4Olz2onYkPdVbalwbdKGHNqYG/371rVtXae151DYrVAvdPQJcyQCKYvNKDQwC2Qi
hjFHs3GJS1sTym1n4VkLBrGFEPccWyyrd6PwJt0u6aOXL8cZrxVuNtKWgZXDY8zY
zQosYNTWNaokDY2p5FNnR8fosB+MFgcasMsqUQCX6WW6UGv98wUYBJXDZOUkw/Ez
uHwg3j5WUbtSlVOp5fPmdZrzgAKKENll5Tv+KqLrGbSbY1dqhp6RA3HsWXoezIVN
I/5uj2n65Bj/beWsYDfRKuiRS5n7R5LVFxMhFDXa+JZSMi4oGcR6ahDyNuFmdtCc
+pXu/yMSm6qNPmBWqYisWxSRod+3Ejr/NdWrwfeiyGRAfO1wiafmRRWFk6ThpiCF
oxIjoJAUGuonEVl/fp4hdinq5Q6mY1XyCYYcAqzJLcivb/xv4LDNYl/vDPHYOWlt
InUbLVGKkSKUhm0oTK8FDVszL2QWgk3dAidgGYkZRFPmKxPIce+k2/3Zb1KU1jtD
vg3UDgkew6UIvb5kfgmXhC/ErNVURoFzaFWUVfoe38tGeRSNvisnyNo9zDBm55xe
FbBdbzHbiU7eclasd6Hry1/TDZLu28H26mpx5JiO4lpC4U4BQnp/nH9s0OyCDu1I
A08tSLXg8Xtvtb5eCpIc9Jek6vLqZsdlq0IW47rin0flNSDKM4uPGzD1Kw6idmQX
H81o0kL2L7u24ko4aoIrCoEeq6U+ziLEasYArbBKo70pU67cirFAhzojNSmGLiJs
U0c9zFbADNQKQVZVFp2Mi0Dr89/jnd5JvazYeQe1TkkdMWf+lQeskrmcFH6/LE0l
VrzhjhUoJAQT8lmN38AA0XhDaN1Ma0SFh6/5ShgVMMY3XFVrD6Je0ypjOUXXOd2M
0dWG5Si4sOEycciZvlzvqd0SpfcpVZIzIsn8PivwsRKLA0qB2hpy5OeBfasOLfdk
bx5+ew10IA4kD0EtLUl6aL2nstNSSnuZn++FDeFADQR3Fypf1A1Q0KyEkyBDTnNh
IYJrbvQSXz8tL0upPspKXN+odom/GMLglj92h0skocGk2a8/suBl72vuXdnCXSy5
NBIiWaRkglgGfO2uRs9QWE6aphTSbMXYg+yD+1U/why/M+NWj4JY/vxWTnNWhOFN
nsSd3M6oJBHyF2Ru4aS5VXHCEhWfjJq7ZzONZUZ/KDt4uJAFMA57KwbU5NOEm7VR
FgoimOqorUYGfTll4GIm3oxryBAURedHxqLyEoWy4oYtzll5W7OZp43Bs6Lw4Qli
ts5sG3Z9q61bCs6y023o5K882aHeUUtYeMp7eGK6AE92WxCocO2ZMCVSdFdCzCqE
8xgl9BLfVAzAoR20XTFsz5DNPp8keHlY+89PqxcJUau0ow51oX82YJ9TnEd+Q7WV
oS3rny8YfxgQWMqWu5glXhdU5BtLy7Ci1W+GgktbEG7uK7gnQlhYUIIzpGAZnhoD
k05g2GIX1bNqVwgn+Iom52id/lj1m9oXCIDW4NBuEoGscSoK0XDnsWzs6wWCLo0B
tAF3zZrUAz632sIJzvWnF5Zwo6Zes+JS/E1A5/0UIU3ZVkJeZainI9bJlIyRbljI
dKKnF8xKOybaq7SRbhOCHfZrZli4SaSLm63+uSn2esoMSV3nzAYmA2d8h93Js97N
2pqT321igEkFlo4G8nI7MhfAoNfwjAGCE/hEZETVj4uASrR9GEr2jdWLK3wrfwrs
7/gcYi4FmLlqki8wMWDRuM32/47c9nAzHQxSNWBqCzLccA4e6sOAcaM5f3tL6C8c
WvCcN9LbPnGb6vSKfW3CbBe8Dfj2Qda43w+3ZtFgtkYFPymIKZ2TIV/Nh+ATs1EY
T76GLDAq0Ggs5NsFxwMrNtAAcXWUWnqHAayKp83NOBs0uUYC1LRMGtF2a90RELy7
dLlFV2LUb0W6vNgho87Addat2ft6lSCyOR4dFpnVjghDVtMHUNFvSqSUdGdPQbBe
HQfR7+HeiBOi+EMddXZ9U2UJ97HVWd459S+vpoWF7KfVg+pqOHTxMPcv6JylRLfN
kPt4zuZkHX/BSfttz/IgqZMTqrAbj7yIkNe0Sa7/bLZI86c3w2PmISfbcVtNRdyw
ysVPeKVnzq4Schl31YELd32iLunIUHaTBo6uRNuFDktg1rpwew+UzwxoQyEqkP47
WdDlLv0vN8aS2j0RdRJ3Qch/vsxj8OwrdCbPWQXecxiSpFYe3PtirXcn5dp82Nyl
kLR/RYMU8V/j11ttianfDNdBDCk94FOAg2d/zrVfZf0SNBX2xwsYX8XmO+Yro+nE
MEkkS+iNYDekpQ0mM1oWeZAJmolkzQmX01frex/uihF16Hb0yv5IcqgoFacWDt/i
W4uKphI42IZo9v+Vz1IyQEq9/qxSM64WBbxz5YidAuFGAyxfWF8ccu1BuYGwkfkV
UUA/4j1S4GmQSZa8O7d4z8aQZiP0PnJ8frjjhjYuoyWPFD0VsGrivqN/MUCjttDq
QYTM6WUoViEdEHDv1BV4kC529QscsbBqd1EDLcmAHi2hydybvep7uAhn9L0GSqFJ
WVXqoJxuxQP82hvNdJKKYytNd/ggkAA8EbzGj5KYvUdFX9GXSFQlEegLBRuTFaFp
JgmAI91N0/HnbzHfDLf/34ApPQXA7rq/PI7AJvzw8Aj5P8Q2xgoEqcXW4hfwkn2F
6Pz8OqJCHK7Tof0Xv6M3UH2hVV2mbbCYwOK7jEik+82iqoC5nO6zUTKYCpFBCcDj
61WDNNLpMogCYS+zfWdD+hQRc9Tnr6sb+Cny2H3p0LjXp25HGGvujY8eByzlx62m
9OKU5zv5zauM9n8AFTccZBp/xyNaZfMvmfbMXltpe+OzbXFaR0+XlHrSfFBZBbQ5
i1wo92sB4hbMnAoQh7yF9BD45Sjle7p0JE65t0Bqj6TPt4TdbnqNim8191gxSf3X
si8LUPI9dvQVbP2PYuFWYEUvO20I9+CRKGdQDgHqgPQ0Tnfcwwbnt3KUPBfLd4SM
YDpcjgFCCTlRCWTWa/u4UljBL6kgYHvLzmx67iI5f3wut/RWaJWSrRfAlRc0D75Y
2zFX7PzvLVU0+UTAo80a/CZVW48LOfKLX+xBGFvS7Lj3ADwrHliM0q9skbMjexa9
l31Pb5dTmpWcnEVejuCIKqv3TiJE8To2x28NXLGzwcB8qT9rHn+jc1fLZd5ri5iA
P6xnXodGUXJYl2cW6J8lmcDeY8eYdh3flh2ga0SBPsK89t6rDt9F37bVkU7pEyHb
QH0VBXymzIEjA5iza44hFoobHLl0jFNjjOCHlEGpC2uuggWOfcjAMoekhjTAdYpO
BF0r77AfFIeKNqPQ89t3vO+MvmBFAQ2w+1uCy/t++8SdBTodzkgqP1oxQsEA5orJ
rSXAkEdNHGQWPGeVCuDOph15dDYCFCcgIxRwogkH3HJnQ/UM+I+a0SOwDl+eWVSM
8i+TKtKvG2URiuNU8Q+NB5FrDSS+e8Fzo20bgplHI+dskhWsX1lKvMUhE6Ag9EU4
eG04VtiYGz6XJ4CMi76Bq76D+F5wYW5zKXmEmTUIyx29wpzIUQ4t5BEiyN887dCX
0vNaQ3uHRaXPYkMr07tQgxMox4EheUhO9qdqvlWKTFB6YXMQ2ZAppv122s8hndq7
4GYyHfe7ISMScYwbyVyFOOme5bx4aB18ya6xKKEAvRNxdkpbZIVBMv963XA9IQr4
Dw3gDg2NWDadlXflbsIxbD7K87kOndb4kkmuv/svux0Tmjb27VuMqE42+STZRsbo
1RUU/njWDusNwKbBuepRkKm7pDOojFT2CY9mp9wR0OkxWmY5aIhv9+5GWXsvrZqN
u95vZkvBjbDUKa1r2Ro1PIWheuy4cjdTgpzqZz60NjZ8O7/KvmWFuP1bWQ+Uvr0/
sfzbJLSz1OPae2B+C5d1duJaQKiixwA8vd4F6dJkfXNBptI/CyBew/0ZjcZBlnZI
W6tMcGArY0Diz2xZ5CvBls5LOeB8XIe/QvwBeu3KT2wlOg1bHCX2KOj7HYnPqMsF
eUMsQMe6fC34bPczQzoGo9Af/m+xJTEs9Al1u6xUVlos8znakDsc5SrlbVFo8a3a
hAxaeTACmd0W8b+E/CZiVNRnGj2GZb7FSNDsErjsNmCEFpZh77WrNpOWElhMLyCD
N0ajkQNT/OIY0Mk8+dVr3aLYuKYZ8TdCoVjf3/j+3LUdWXT341bOCwlu7MnrsB8G
0CA+ydH3pqe8NReuXXh1wGZMYENzMyKxHMkD+9egauXmdUWosGGZKeCX1xXTZIhG
S+6QW1ImuBo1RXnUZBmHse7cVKmozcyWJIZ7LorPzjuTTmpft7SEeyA0aZ1M0r72
0YOs7HgPNdjNoShxrJoVYJYMSZWIfF0ZdOy2KMpgI+mUZgo7j4mc9uiVEWjA71CN
6YM1fW1wzdh7Da173CiX7QpOlcNQnLoQ3WJbnfVbD4yNDiIUSZ7Q5lDkwLIkaSoc
4XyYnnQZOAe8dw19IjEsxzWTsr522p+71c/HFvRZBlZoAmwjSNMARU5TX+LqlXRC
7NFiN4luARs30I92DAmWzi01Pj6CJ9U3gl/7YItKyu55YOtLHlDbzchcfqLJnRb6
QGeqjJ2NRYncwgnggs1hkPIR8CzXAX55EyKGXGf/oLnwWQqrV1CcFhk0xjLWZyfC
Rg1AXhCkt/6YavF3lMT0m3a3S+XJdUdFERNzb3WxcHUQmaTDU+RNUB8332Pt43j+
40zPfov+EIh9x1mHMRr6RAB80cY5l5Q48PYQnsGDRoAVErcOAIS217Gawuj5x7WT
xxbFy6ZBBdjBEYpntZoB4dxyWpvtL6qVma5YKx4aHcKE1w/1GgrvQsW3bhAWtNf9
WYrKuBWPKXKfaPFn7ksO4kzfb7OfwbqjDy1QWhyu0xoof8Zqtp17LzSI//X1O/UJ
kgYyYwTc15MyN9Ni/IZJUAE43xoyXt/kW15acfjwbdx7QQJcK5XLrr5t+hjpzECF
Ftf73M9X4F6iQBMrc07+x/4QVyG4kpVcPJgYAu/Km71KCHvSF+RvX4HHU9P78Rrc
ccxrR8zatjn8kpNhcIvLhJv0iGmtWgOKxa8nP5j7k+46PZ6t4XF5d2RrZyb7UcQI
6oUc2hke+w35DbKchs4nQRVRrvaJfVyBfCKkkdzIn8b2QECPdKq3mBrF3+4PzufM
liesMZjtUo4Pe40fuC7jCxMeQ78VrLlgjmRwTTOkuGKGDU24UKbAD8NlyPRm2Zc2
TlaeMSCpDQeWtVKk8/v+Uv2dVUZxMDceQFGQQVFi/4oUWxKG0/M+8Fw5DerQ0znI
JyzzU6LXe193aqCoIXzSIeRa91bLohs+MJpEDK7y1HasncN2A26AXD3Vdrjrjm/U
9GgwBRNJ6JwGu4FQMpx5zAt2lWUY2p4iu5txD4FQYIrUc0lpLBA/tBLA2LgbRViN
RHTOVT2XmLgeRrVq27D1FnLyfmbBn3aiO32FmgDFEzEvgYPZMKQrOOY0JMgmQWbv
FGxHVcqqbvE9tQ45gnbh4baTo51v6ao/9V2uINTNEgVe8tvncSgBRsxYezF4/hv9
TCOyUfAxgCIwutx39BJp1hNY4VERyPQpYMS2p0hz1weMarFh9btNiqhFvZj2N2/I
AMDL/EKnqq8jH4pgrWmIGvuQtTAymCRtjGFANCbzrcWtJbNFVHRqyINVc0X3O6DS
/DKoXcCaOIi8+zBLtMPzdQAO1HUd/qaPvqGy7nT8YPtXtwAY1ZIMEEDjQYzjm2He
Xh8CElMb6yxA+dhnPsiqEfvcrZrGF1F1VjjW5OmEwWLvkC9IGAx9jBL9HKR+iSd/
nVdwFJARXHhKBMwkVd0+FPJCyrqPQ6TQ47bnkMXbtddVOhCwOldFRNz3M2ZbWusa
wT0oH5d1NEO034BqvGgMg5KSow4EzmMl8Cr0BDB0xYy+Qcn7AiIAWlCP1gDzEDJK
EXRcIBq95CqyM18gO4updTu7pVmrFDgCgDnBrhDMe9IvPJUAaQ3/xnq3Tg/CGmGU
z/MAdJmy0ZgCkrLYq773hhg+VMyeYRYBtKKvd+J8K40B76LCnYsQgIP6V5OYudaJ
uej9l/V5u5u3GKjxFch9f4p/9z0PY6GAyq4VYxTDPEprGKMewxlU8ZaA3kpROKnu
ANL0XRd9AL+bwvhD5bir24Cb36CgvabI5QkE3OcdU9z8E1U0iNxyQIehMr4ZBaks
evzCNXNBLuMiuGVAEyA5nAVaT+Mtw/ZZnlBe9EqKJgrpfM7FEVrwdokCJ4HwsSl5
TtrEdISihqRbH4zyr9S7gQcVSepKe+9hWT2kxHfG1jMpbnf1NonB84M+p8rCj7Dw
HYKr7QLedx93sZW4LObaOvtjitjRsZGNSIo9Tfow3JUytx7UzQDGzI1OwGyUb7Ox
TWBg98I23uemPzkmEzcOYCCO3UKaCePJTDMAe+F7eO6tTnU4p1PHMfTMelgt41fo
Q+/90qCExvt7pTnBVNBh2b6wU3Eo93Y9HBocVFvEHGshBTlSYFs5xqBjD0dBKmsT
sCJp8TP/o3M58KLCnv6HpIJmsT3R8E//qS+IUUmWvl9hZe8t4FBawPcDVtQt78GJ
9HMN3XHfKoT3whmMxDVNTfyMkxJtkWsxCiXoMfl0OBkYU7GgSQJICkloFiVrHszh
OzGgTgcECDkqzkYu9Qo0ZJDUT/T7vfiWIy16r9o8LXuJ3ThbeuRb4aM3gcPC8YjH
ZosPWmfjSjiWmWs8SDPmGUEs/JNc3wIsKIqw5P6gi820ohcLws1EJTeDTOCsIXpo
xa7FUF33d7pkYO5wOFP1ThH0lD8u62vUSgvivrYFYNOMyM44yPyBgRMEV/b/f8eR
An1eTi4imSaUmZIhmlMaK97dspmDFaVDnB4cRVnmvjeMjxHZ6mdcxxdhlbRsLW+6
/ijQsVK9mzVjE0TDZdYLS3790yhLsJQJUaKGs4YqMljLPTYaccVXFceFLqjItV8k
na6MxuDFPvlhKyyZ9fBrhhAvXPGcFOUNvVoeuMcirtFhQenNY80+gbXd7aT+iZir
EoH/0rUB/+JEQ0PyPZCTx25qljwWNyYRlb1gRUqBeTT5ADgxu2I80WF5GdPNvWPW
JID2VAnxLe5O37yVEINIdCuIG3VBcu448kHkOq1Avy9f7Em/aEyJpI0Z9qtlzAof
FgsmxzYpH7YV+a/GScv6F6UIDu6GtcLLbcc/yLo2Dg5Wdqy8qb4wGATXxZSg0zaG
MIadEMBNazmS1OOoAgzJcz92vp0BVsWgqR9IQQR6qd9P4Foi3pNISJbg07XO7vEw
nu8kCiV9McwZ7FZm6WwmCD6ogwygHNcdIEW8qRpjUfzo7T2qItgJt/4TTUJcEl6j
5SZaA09cHjLEdX4EVJfOotPDYPypkFxFqc1Dw8dKtTDGEYJeh7VxzHaPqRsgUqTc
9bqpgtAEJ9gx4uldT0ubJ/E/zn4gLQlZLCh96Q31p8uXxVuWMR/DRsC8OcoutSXQ
gya8T1gyiqeMcacMZJRPWNMUMZpsr5W/oQMiE+NQDaZLOgveH8NoaIrL+BcgRFQq
FdGxaNcJuMtk/DtgGTYmrk/vyobjPVRC9oVtq0syWmk1ZmbZ1kFrFiN0ECOGnOps
O9+RH5rbC6NuqWaqENtSdpUxRmZg+VtaABfzXtKM42FnwfWyQK66JIOW8ZcRk5kT
tT4tWw13LyrS0GFwOnbEAfrB5w3KAGINZyIihuFxEa/XAYxqN2Sx3VtQbf4ksRc6
2Xzq7VC3qWPIQtgfup/O440oIh7vS3qP3upN7X2+rd0ascLCMg77w43/LapXVELv
Q1p0vvNAuHkdUyNjU0Ie1o0/j8sKO2II4W2nWRxJV3DRqccMP1Yr7MmtvxtcQe4+
8ksqpKhPjASuDxUIopRjlGFNf01I38ljKAtGyfoJnpGBuuCJEwtpUuDpfdLZitaU
z58ogqKPtSRg0jksST/XMgAFwNDWkv1Y8vx7ZdS9MTgAjspTxgZj3j13b2NVDTtv
MhoCdIfFCO8vOPOn8d5J/Tu093jLPlYrgQAKOWFd58pGtasWbbUzij75lGjcIzJx
DV+1Z4gwpc9E3LGsIHfknWc8tG5hX+snIt7XBgnwfKc/JU3t0G3owH8n/+2+Yo8I
r940QdkT/WRzojDsmF4eUAwsPuvlI5wmqjkiTocKAMhGM2Eg87Z0VOCsaWaLEANN
FmAN6SfE8BieJT1dwu9uZR8CNV4DjkB/kDJiZkEJ6jGkNALwC7GMHNEzDRpoO2/L
R3sbbId9XDDdotb+OXsT6zzG/dnmal82TDETg/bWdmL0PNbzGbxAmZ6G0ZeHWUEl
WQrYdDLceZo+lyJulR6L8UvYvcaIsQ+QRuXS2fsHs1Di7cckt3ltMRIB3GvPVCi3
bPPEjS0++rlcC1fnXvclMaqN0wz0dXz8Q/EUR3mVqqa8wK23vJAkFJvyLGEXtAm3
5E/L3Z4JX5qkser+D7XG5MJzo4rf6RUuPraxzwtSdOfWgejpcdmpN9GQ7/nbrRR3
6zEkw+CJdymfc0/DvWsqlfZmDaLwCQ0h7GkAp389xq/HOGX71gvmySTEMc+0aGzI
kDyICWG9OrMOAsRf2MTdSaavgSTLDkr/9huoTsob++11yFVkZccgt3A0bEzeW6Xt
WbBNs1u/7/kllfcBQnmjcmgbZ79Rfdw8pkWSkODSzk8bh4Kg5be/v49HyA1AzZxh
QZ9Vgo1dJz29T98HOmXWx1gpRD79vLD2oYQ2ByEaPKO/I3NZ3TpNPQzOySrfLCpX
XwAKFt5FpTJZzAdjtH6aiwKOOoqo+65Dq3gGuVDzyMYPFprZasUX6pBRRtSLu7Dy
3O7dWIY2D2+CeeYaspIHvDGpo5IF4U1p9FI0K944aCpgJdbRgd0v4HfsfxRn/J49
sg39h5NfzUsHXkETDcgUuF7vLaNQmok9sl/W0AW4U4NXxPvERbA1MHdAMSV5uL2i
D0RSvzzIhAtJu3u5F7rgmPZRO7/30XKKcCUjxEWg9zQWdvMjxLM12EfTIbU2DFaW
oeO8ZGeVVT16jRTjzniS8E1BmkUKHVGEB09rlkB9Un3tF7AC1RkjeOCgSJfWpjKc
WjMYeJWXj1dtkz7IGd6z9+FK94njNZGu0P/O9U3E0P+KpbSoS3LgEtZn7I6aTEog
auDcCJUGgb25aNUOrrJNaq8g6EDOK/3EVQXuc/pfVOZ/aOZqugKi2xPCnPBIMYfy
/mXZX1yOFj3xPphiO7QdB2gS/3IjuVh3tM+4xD4hzW/zr6gbjg1u5asE+ssViLfe
gkFhxw8hZ5VIvaiB/xW0F0c8vOkhQS1bb2zhDorpz8DDojMtGipyvG1U1X5wQMPK
b7OJqpqZcyADIkfcLKzTKTfQiZrjoPgVSy7gXXysuCL0G7kNBQB1yMS20J4idzBr
JmfvNn1yqRGU/2KfAuncxN1Q0/QS8qeiOlYoWrm8ihvJe80jMBoONbpfTy5g35+g
OGnqF0r2AyVPiWa+N7fczrD9+dEXXsBnyl1MbH8Sqesx2b9BZNaKSS2fb8TODq5O
oX2CHiWaxD4Xij/+pY7Z/shcTeSLZ/XAL+jaotnRqb2v27HbWgFrl9HFVQKNPq1c
VVfA2hdm8xdGz5gL7gDK5d7X6dB8NpMZ/iq97HCqPt2e8RbX1cQOLtdX35tST18H
1S9rxGz23XfHuE13soykujSVQI75jBHp6D80qE0ucD7P3dHIRBxvmuJp5QlyIvP5
sAhy+tbY9rkwPMPFgbZn+UxvB2JgLX8yvOWfNSlWHifJXrn6Uarlhw+mXfIVkySK
MPIYFknjpG/f2FJy8c77IUqd3zwa7vpsrqi9bBPJWvmXGTzmQK4+bBFVs3vwYaNY
IaGCNZEbACLF616JvaYrOjJKB9eYGRBHf+9r5dZrivWqOtKd06GCF97Xhryhie15
iE1ieCVMWIILsX71jIxhtqxjJlIfgVd4/KpgTmUrKHMvwXmVbeMpAP2v01bdNRs1
MfCgPRap27nlFavfCYtFuKYzNn5cL6gG+t9LlKXqslLZTfPh7U4b3Dgaubj5HyNv
lELJMRUNdqqnnlU+AtvUTmxJcvGhpie1c1ItY2b/hL7pB8DaqgIkLST5/L+XPyDq
ifjTQMIKokrAXGNe/QQlJW7Z/2iAbRAHFjOetXOQ2u8LOATKeC8zkivWo3Oyde5O
GJMDfhTGWL4GBd7wdRFZlGehkq1yxxEtHdfYJCAbsqsYI9lvVx6u4bQC1KCOyaV8
Dpp/oTIUTkGU9fBu/SgBsN7KXSZWNTXTT+BeBTLoRQsv+EUk6xy2SVgS+LPn8VPI
Fz0UCJr5XWkkN677WK3hVNGBe2T5nb/lXC9oUvn5/f3dqoG2+cux+3QLA3cLiS5n
/+1M6kdjlZ2QE+hPa55FIUlEdUB4VsRtHaSnYHeJzNiOtc6VM48YbFvpxZdKtC5A
qcaaDXLZ4F0JbzoLub3v2AQFl+xoCVBsxc/e8nOtOwY+Or0Iaf7N9jhRdfB0rBau
DCQZ4Whvqh7cIdhN5b/VlTWN24KAdDw7S04uyEf7xJNsZ0fyvuo0WFxIDgZ//yxB
YcK+ObZBpr58P4ebi/VByoAAK26+ZjmXfmAh8AEcAee1I9Dt/vE58RVwL3jrftTC
sFsiaKEYtxmrBQwaQ1RCiwDSnGellwjGKa6WWM8QPE1TPJuJy1OhjKtHMGbSvkuW
2rXxMLYmjxlMGLZXMapmJUIMDM6k/VEzXBle0U5GuvK0oILyvdDVPemnIBfYm10m
janUYHTKhqxyga9uHc6zMgdvpdDlJbHJBPHebt91fdLmiR3K/7bkmquJTRz9kgh9
FtL32q9hS6DvqZq00k/xIOsit8xdexDMF9+Rjl2STgE0UFEjRDwlxc66BRvCXsUu
Dd50K2RqwzV3VPqpCR+gQu+Nl4pSz4XAD3+UJ8YAn9iPQ89VNmNKUlRz+nJV26RH
sfNaHzZaado6LIJ5tXBCkDjWQGOjG7bpXwkBDlwjFtnWZG9Gm5f5vGeFS6dCoTue
1tPhsFkbHmf5UrTDkfxDPXuvYDkvL7IinAnk7Tq+Wg1POE9W+CtGz1lg2twYG3N/
2zQg4/lyPqTXS2a9NPL6OsDHovl6epR7+90E3NEdP+A03/pC6qPF96unhRR+qBcS
202917iLkyTtk0BqEnjyvOqmTm+XRrtyTMT4fHhQ8X4d0cnSHE5Bum2ZVipC06dF
XRHKf7jv7s134Ng+N05AiBsg5ynu1KGjJ0tSywYOA+i4ogLSuD1u/W+SCdaZ6PPl
B51V8m/ZZ1kZ+Ju0jTP1PzBvPPTwbDMBMxN40F1rQZzCrHS6z/MrnIX82qPe2j7/
W6D8c4ZepWsynZ0oUAylSXwlqseMFWHEjd+JRAJe2nksA+a7DlH3ane7lGUN0QAM
b8dLA+CEj05AmPf51YF4GUJLplG7WUvUQa1Nk7IhGrrYAf+pM+Hd2r4QGJM7zPSr
+3+uBNid2lbcRGF9YoAJXQ9nwZdTuGzQ85Uxjbf3BXVmNjto4U02UzJB28MbpG0w
6ZumUpze9q+Ti2v+5M4A+TGKBhHRiPl+D/mrL0YgXP06k7xj7tsCjqXC2mgI8xFK
64xcBA7VaMl1wu/K6SGclfFoUsmQUtgqGfR95DqCc/ynYpk3gcT2C1hNQJw9qLLK
Zm+iJi5+qyU1c6WBTVkI1mZRP+/jR4c3CJxxZ5nZKoVX19EAjCVLzHRkLpzXsBsT
gBeOeg/WplN1mXaX7XZAIEvLJbHPfa/vMlzfJEamNCm7ozn/E1f1Z5wF8rPKaBqL
BJ7VGj4J+RCEN8Mofc1URtfPrR9kcFm3nhtlln7ieAGN4VjSrSUTXkTv4OkT7wul
nESAd1Lz8qt+Bjwk6l0LEIfnbOGZFtXnsgWHe8SoIK9dCBMnpnl/mVBgvMFahTJ0
muy1fg2OTPImI+obR3ooGROg1Vu0jFDFa/ghH7LjP31NlNMqWh+Qeay0a/noK+TD
XUdWfWpA+phu7srD6YDm+i8VvDYID2ESKb/Opqg7TXUROfNivG/5qPHZtV0pj9Zd
poX4Y94jg0adY0l4y/IKu7QmpOdcwyNzJinZ6v9BYfjFAACy/Rsgzm8hBtBQ4iZ7
XW52S0pStgzieFi2ODt9/DFCVqKMHg6qspfY7H3S8y27TMzjpudJ1u6XbVHsnwHv
h9k1eg9MAG8gA8KieqxvcJ/+MMrgvVWrS68cgZ2IVGrxmJC9FZ3IAq1muJXETceM
kS+Tdr7SLi35Xf0MAUL026ohcRnC7dkFTXhVlE/cy3bM8JXQKhTQ31rIsc5xHE/u
FV3El6hkhaEZ0/Mu+3B5tJzRfcWWEWGPIQ20hQMDSawL0NjA4qjXmxhKPB16NJWa
U1m+Q2hh8C/nMdFzXgbBLy7j+V4s1YzZP2Rk54//EnLBVW+uQ1FjejG8N1pU6GZG
36lhXXm4BxHAvXMjd8Kzj2v+UDp5a4f6EZ7Ve6OosW0kl7oR3NrKj7Ibhl6PP5Im
QoTaQnY8eFPIcKzOsuSiL+8AMFQE4MiR70KO+O1yMA7bDrQMHxaDPOim43YOcvHX
yeAZ7JWNzQMbOkDEKihONR1bB6myt3fBZkg242VGln9jCgBfg88MhWz6d6/2+9km
rRqJAXjrVp+mV6zo2cMV+MWpi2R7IOjuAgSJYoiik/dXd1YFNa+x1JaneosQWymW
sTDnPsdarS1ud614XDQPUvYOJOc9sHTI2dTPvnJF57qHV/V2/W1iVagJblB7gyFI
AouctK/azvS/pWPCXFU9SJM4MUwYKr5jKhC/EfCAr525ljFV6h859DMxHZZpsPBc
kxVJpdrAsPRy0OCtzOHcgA0wkA3cX1GBDbJFXsSzaUxzNXus6tPzCG4KkGuMvCzW
HZAPZyQbmSXGxby6eEdnBclAnZggFkXg9gsaRq0tFtuIMIwfhJagHeRhyg+TWqYi
TY4PG5E4rZ2/yIptXi/B0Ih23yE43fvnDDvdu6ZUXXkN+5NPM41RiDcZMgRXBDnP
lHEX8uBYGcgeayQfEA56NBAMro1C5bQVEANMZV+4X2PzVrxkpVHqVDoAWAtiFy8k
U6RK0Bd/64zBxiBbLPRLD80XEU1GTzKlNhmQFi3PvsqNIOXfuAHfWYk66rv7AvLl
gzZYVYLbxzTQoyQWH+touBkrrgh+57Z7PYeJSD8OJWn6Pm7MkHsypGjOHf3/GyGH
gDHBciwxylTpfDxc2QswM6hyz3TlJ169SHbumEVTC1zCx6tEVaX1x3baRgJyBdGx
YBO2Azapiy4neMLK6jFh7U3fq0JcbhduDKKoaWI6mAJu5fuyRJ8L9Qpjt0ajCL+e
p/a8aWx8SjqfCvDvorMILScoj+FEHI3OgKPAQdgefQb09F9Rxc6yltW4cy6XvYhF
opge8ladjDOvieRlOQjW17afAdjm3Xc8V5tz4MRqTG7tJaFzxsI6XD6lTbQVzLhz
XuGhR+HNoiVmThPaTzYZICg7N3+ZtlO0DEo9IYELRohJd026ztWNDkCL6jpJme1/
Gts4pVb89NApzV9RDDgKOthpvOTjXe2ITmik5DD1EXwbkb0rWdfeDncaO/0iT5Na
UBMZ2bWkQ1kpa8RA8O1/whOmsWyoX0leT3nWoC74ZZNRWlXq9bep592eU11aLoYE
pBnQBgVfBJW6j9sNgNFtFSZids3//o3STdVKI3EcLoC8Frr0xjdCcQCjFJw9PraL
DnWpCoRm4Jx4LM6hY04lfJfzVF2xoC4WT84IV5jGSetd/nteOeC24CPVN+URg4mr
iDSyohVLpZuXB1VDWCyynUajbViKo//gtUPJhzO1dh6Qbo6QpIEELhAnGrn722Nw
cbA6RbLiknkxhPuLpfxHBLjfLNqtxj58PZNeOBEKKWWnHyabyeiOoSfVcdJBeLmw
8Ze9gH2xXDei9eIW7RUt2Nh+ORk/vFHRYl/J507UuAlFa7uIlmznasr4jL6RG03e
VrvebsfEvJ+i8o3I5p6Ebg7Xi1wvTIE8FK1OwK0ccGaKDuGQHqu6+3l9ebt94G/q
iD6ZVGYYw7H8aPBvNgWlJz5LWs9wDHB0Kixq6LWc1vcjy1SAJW7I+9LsP8iFez1q
Ob87DUHT2UKltTAwCcbmQ76j89z3p8OHxx0Tr+XOYnUy1kdRqeaSDgk1SVTZF+mG
ehP4Bp1LUtRLlqoaBSTBrUid6c6fFR3adwWdkNIDoWjchrpgG5zfPt4uaFZqJHyL
UmcC+5mIb1tZZAzKHxCetxGb7QHFgazatP+3rdi/cXiL7I33VotXU1TWYm+PxM9T
CtlqgmloaIaFL9uAXvb4oHJUhWO93BC5C1QIzpKc0v/Cyb4w2O6e4b9xdqrrzMAN
VEvLYB/itqi0XWQU5ozMy5AByjSRNp/hzLPGGEHBwMqZ/1ZOKGABGq/diDuDrUiD
TMmmXTT/07y5E+SrjkBw3C7C56t0SJrL+d46r1FZgg4iwmii3AqMYWinRSWU4z9M
vsMr/QCA8b+EoQIDyRryuVU23DOMGlVeUUm8PImsHW+BrCvpf93fgGxvcUtdMDjS
zEl3lxp49hLpiUHBMEvwVfx654XImh9lb1j86qSPKJGxnEp1lEzHuTxoMs9TeNy/
dCOxi94DTz1pB+1sxjwrkrp3ZO8A9AhRNcW6FRNBDR2o6ASW+ta1PBYn02AKEJ55
B9Q+Ip0s4LIClfuKpk6r0iveGBrMd9yKdIhUzQ5WPcJmUMsOVGizREZYpDm/sNUL
TSxvPwpUaFEirnYkTZX86XMSl3KO2LNY5yMIp68RSqXAegLJOflNeJm1wY1O4xIE
go6NifwUyix+aKhUXygKFJvk1sE1w5lczuMwyESMgbIkejjEbBz2OEoV4BoenWrq
hbles+BX9s08I8A9z1h5JaVM3iiro9x5OlBa0blGYtdmA1vO6+9RRRPTHamH1/X5
70kYrvnqxfZpMDwVt4XGToaRM4tPBjI/+dy3ul1inaXkwwLSFweGn6iKEaAMpsvD
Za3D5b/is/bJk/XGVLaHtlxCrPWEGKhzjx+IIXvv/aEKgF727+wL1SlWZIzzTHTc
rzoSaZpwaGX+IhERs/6naCXiyK4uR1qkR5j41YDAcgWLojeOG4dfWyc+7yRwpjzo
cBW0BM2WH4Y8yzbTPqLURU9AAPp5Lh7SAuzVVf0OyTrP9KsCZACWB7Ve8rmX11R3
0e4hEQEusjF8V83r1mFDWpf3lWDVMz+iXMivINC8mkBy4yHFY6sbG8NhCaxk2b7Y
Tpw+MF0PJkpn1eqWGxQDHEOZaryZ7+LUbcteDT1B/DceJ3EXe4AjGk1NL82MJlJa
v0JEJHakcQ0Yu0HJ7J6zYNq4zqfybqLOyMFTzINtioIOE7pZtEmxxoVoZ7KFX8va
7J3LFROQ2IWY0TilW/sm+iq69vp14b2Iz1BvZ2SkVilMR8VJJ5PT1Drw7sSmhfp5
jQ7st0AAETkVUP4mHB53vwL/AiYscChuRc7RBzb2VKQrYH5OwVMeIgm+MK/vkS7H
omh+SKOmvdB0oN8j0KwSyi7v7MHQRR5FZzDiTjB1OmkVOQktqUB7ErliuCRuRGtn
jpuCeeDPEAB4dTkG08tQUq+6TQ0iTC96jQeJBNweI8s0OinqTHGKUZHNsztvGsfP
D6DekfKGb6hL55MBa1bvdA/cRlT818XkR3zltznBCoA90WaqmVIAYJ5YEu/6tQoD
GflSg3oj96ydElFUZsVM64FEwojB3dlC9uwdSYmMpFe7Gb/9A18uRk9Or9HGyIYz
PbGhS3o/SDjbfId/D8Vl/LEB4lZXI85bIvQHpUaH4WdMFEdNvobv6y+l8bFduLe5
jhqI6enEeoNaItghp4OytFzdyHVwzXDTZ9mdkI4hBUGuIoO2zXoYyuBnQZffumW4
+P9oMyQveWZ1oibCHEUxwt/on9mm5en7I98i6yUZaPBR+H31NEoYlvUTW1p2RjCb
XZKabg0yUU1zbKMJoYt+hBrCuIz+ScM70ThttyG5RuBMT77jG2VVkzaME+unqAPR
YO2zTbf6tbGE3iSpanPchb2pSW7X6h5X0JxS1UHPzc0XTSvIUsfY1cYi7wQQ5LvT
+p21ZFXwasc24zpPQlebeqs0i7Wrtgad2WIB8SCnHJDGQ256iNkCyOIw0JmmWLQh
EVAWkkyAUXhPXsd3KSt8n4mRJIRKVk47dmh/ZEUwlVSvcQfnicfMGrFnjMEbRjI/
U3hlrGnrsfYenPb5BOoaEz0TOeW5RvmBnFufL54GPDjj8qqdcoeMrjZ1Ujh9C9xF
TSwQh1EOMpCdA+pA2KbKVIC+zoshizj4rdZ7dJbgzTAuyNwrBcktHo2TcHzQkBL5
7kKZeoWyQl9B9v46ibaVQMk5C0hZfJJ5o/edlpT5Y3DDbxz1+4aOR5gOsFQhM0ek
W82y6I52rAzmy0PCUUC7oLd6ENT1qzt8Gn21KskXWmD8psGkEQzB82SVIY7Bt9hz
NSQujit/Pdzl9412tX95Rkr4PxiDDDSNuAv3vAnWZUFOn3C84sYJuWbO2/5+hIuw
X02XDrDnGupgF/aBoAtNFRuhn1///VG1kDSrmdOLHnHReNed2viQl0tgYVi9TJtZ
+rViypMacDUfLjmDP7LaJsyuqePskcJ5X8OqJ7/zgSzVj8wyUdsSFDpEFYzPqbiZ
H8KYE8J698DOQiFS3R1ARVgqrRFFDomjhxFWHfdDBuUI76Sw9BRXkYpvroEO6AdD
1l/jIcV1Yl2xHHAT6V2VuAm+6t2RefBW5YDj8UHaduavCKJ0Iz7KIlYLmMk+sMLP
R0AZ0GgoAm7Fi0Xjw76Ll4rOue7FWxMOkxJt+8JiOKBuGI0K5iYSv3x+ub5uteca
Vri4MkvVGXpE8sZFWhRzaGqAkwbIte8+I5dBgHcNQvABbZn56jRSPAopCXh999oX
I58ixsQkaT3JMiM68Mks/LzfASQmVVWoHDdL2g0ddpdZ3XQG9jQIqZrQfu2RPXR+
bAWo9OuXaTyKcL5f8Afp8fIeKYlNVz3zi2pckpNFqinu+NF6Gvv26IyeT5MOZtUJ
Z0J4C3MzVEJLT7ZOpQShxmo+rxbYXFcW0Fqzm4fEUgbIkqQHbhDlZitOTQZqQwxm
5uaY3159ONuGE4eGTY1qHjp3mKA9O73FvEC+Ab/smuQjcDdZ6tAwKzkXlN+Bx3q9
x1c0QEUdTWEBhwWK4OxQmaOsUX+tJuWNfruiMXOathSF+cxkm/ZiaPdYyEYgt2yB
+h9ENKZpF0XrFpCL0HDuYleR2zcmYpUo91u04I7emRsLizxEHi77mGnmAdCYs+yU
rjKFy6qAzN+k58Gc+hPhOi7Z67CLT1TJ4fFjMwcAh+jrVeXYmZ9HNruV16DgIf5w
4jHlhnSnyYmNcDPpE+U2nbSNCXwDGmv0/gjKW4C2gMYUUPrQQIbxCqW2LNSu72Ph
dBZN7G5sqaJYJxsvbLtVWeHGt5BLytmpCuyEHNiSbzmaub20wdErSxt+DwDPtVtp
Q/5lNA8bznI4YuOxRRpjBvFryNeszND4xHOuX/29YrbrY/VGOzWls08rlRefdopB
fsWxIS8wWpGKgyRIXMi8elIRS+InTyVX8AY8Xy9Zbvn2h6kpke/NNl5PosZuQAkw
1/i1Ve13os2wndAvy171+tGWyN9anYEQV0T86OCcbV6hm7CGtOcS7boku14lQgIX
0QzdXFDJV1h69A4uq0hkkMoNIYS5Kotj3awt6dybC7cz+jDIoEg4zyBmTwCJYTOW
sr2xSKOtUGm90XNszJ7KJwmRsqD36cFSEufkfkzw1GsOvnJqMDdyonAF+nuoqbvC
98n7PeBCdJFDfkC/ve8otBVc8sCr3Ne/DL7pWXLMx/CSGqoTSLeRXC4WxTOE6aqr
RlsJ5LEVlfCOE9o/xeuhyRuehqBKTxnR9KGbpws/KJSZcQtAo1LGzl5p1F3Ev2aW
FkAu/RMcwOtOtK0q6qO5XlSCDF1nWoyXOO2QHl1q1kUd6NQHnbyzoAdqGxwuPMrS
kRhaadwDcSFyj6F0WKrUV7MPLo6ZHcRQeQPNMho7C7QfYsmROID1Hfel46RTCdiJ
R5WTZsuBgavS3F0gKWH/sgDmz7oNp+QCmgf/PqiJZId+GpD8xjK76P/mYpwPkiwq
7L1c/OvIBs8gD4sJYvzKSgP8LK8UxJLEhR8tbTI97EmdvfrmjA1ED1MrPls3/ZrB
IwjIKPBLqTZZI57LQ/ECQQ0iGYsXYSyJxPASw2MiYHy7J6sBrLf2H4uknIp8Shew
hUhuTJYdYAXLCBsAkKJWsorO8kebDvI5i7cQyVnJm/uSUrvJ0jGNlIZtUuX4ylYD
drZwV+nmNeAogqtGgewRzToC/khH2x39u/hpO6VEncQdy/5h1CxY1x1wmcoPlZVj
GNGA+yG8YqUg6+FLJABZuJC0WCKIylJnsnOBmznLy3vCteg70UidNJxMvBYpCfmg
xSZwDio2IzC02uSiREp5+ft/k8civpZqQi1j67bdJ2LoA9qJavI5J73IokGWVnWt
Og9fDGCe6voXnX4fnHrk1JT/8mnpWh+HTRrMGqBCazjUKkDtCcJWhMS7aGSdEHE6
Y1ymnaVjvv8HwSgB2XiG5LERRzXvfIyHL+d4lnuv+o140lDlqgfewAsFURw8Nxdv
RbL1Sqrq2JFV9+uTTnpTt1ItQa6a23JYBdpUEGAawAcAEWokMgzVdcFC1aa3nKkW
hj5w+QPkZ64/YXXahU2LkMxtNdj/g2gwLx/WLhSgvJFShLJaQJ1jBnaepxoVZLtb
TkCYuz0ZiuYjfTAyTf5WgbzaaUsZ8kV7Q+/ffOapHSj4gBYguIeyS88xg2sqLf03
gxYyU4oPvNbRdC6O6wooxICgysHtDN7WDIqnKMahkRAagdPccceKLKmMBGUGyNeD
kMuhwue6H8v/J+95lLvS1MVrr8HS5gMGXbT+STsiPZReZ6ljBcyNu/PmWShrWG9h
OJconAC7uOTSZmeGvQU93m14z6K8mzt74MQDRvMXpVocXzzQ3X9JzhXuxmhDE+6N
JjKzDrmR3SdFa++eMSfBFX8RdIicJ4sZIqSzf7w81D+5fIb3LcVvY2q3/zyDvk7j
sFdoP+76FDruLx9ICHSwWnA38CPLzEq7qVDeYS4zdm+jQC6rhJenjB5dP3/lLryd
ximMBktzy6Bt9puxShNq855WftGgZ9aI9JApl4ryJFxlFe8NCN8QE2h/nuNQ6vIT
ezx9LB/c69jQrzM2vlaio9sGGe9JsQk3eWxtagWri36UdNb1y2qVemfbb9KS2L3G
FC+peZk26nFPfkLGnRMW0DqvsO9WY5TlRfLmvJ4GO0JfAU1F6kS15Pzht23i0iHk
nx6TWhvCHHFJ9i/o678wDu5Egz3vRi5Y8Fzfge4oWAzTq/Jsj1W+9mc6ks/aAhAx
DHfb7KHTNkvm9RRF9glyuvPU0DdJfitCIoXIQcRXeOgYPTy+0P0ScEdOOesq3tlj
yp+uglVo8wJif5wLg6vtTRBVSSoRfQRxCUP06vui7tM9FhWu0EiLGdjmquBVplHx
uPI5utlVuO5v3I00cn8q++uS1JMkyBrok/Qo4/kDMwpOssrIbLpESxBlTuInMZk6
v5EIgxLXcCLfI0klApyYrzlzLFwHXewT2p7MB5ZXHEYpwqhU9jM/vaszaOr3ffWi
Q3/7pRnYLxi2h3K+V+oLf+Q07Z0NDPn2dRXS2+D40rddNUTIAJVZq6ZOSW9/4OTU
1QeVwQSX4aU0uQiDT5g1qayiiJpsZVf6+hx6BNJijuM3iR7Y32YPS1zPsNRwQc5V
nwMeETnb1GgCdvAkbRm0JKZGeHu500SLQmqiMACzTDINFg4wv+Lc0f+X+OdyBAwc
ldzk0LZx6up49Zw6I1hkN4NlhPVMNUlZtsQMJyOs9/Tqt4zPz9I4Z6Ns/izdr3Qd
BNAyHeNKsbo0jwZDiOPyIH6LBaTcq0V1bqngmYqk4N9TBzY+qZ3ySLuHh1Tk5YrB
rSIB5YDmhcctF4tGgV4/OA9CzaKndCiMeFeRfLyPD5fgqfH0Ds1Mwtn1oYDn0xH0
ih1lraCv31JKtS/DeYgIjOZcM+ToS0gkSGyeOFSPXjFbKLnv/De+q3+4duFcK6Tn
ePnIsziy9ohS3N3kL+z5RoZCW+xxkvgo+npuT9MXI51xLF00u6HZo0sYuxiK7cVE
yg9bTDyJQxQMu0093qNZGtto8YUAiK9qxlzCJ8UXVzA2Z+j5GiqRWIre1rYpd2Ob
SzCgzRX1k2sUKTF6jafm8r/0uQEUP1aX98RNZShXDMmkX/IFm+4k6JfQS3jLempP
mQ7i/+bBLDXgdsVfhPFfokHNlHkqIk1PtHIOYC+JKg/B9eEInlUoderwiXx0iu0L
qZyb03om1/Q20mG4wNMR5PC+I5udy52PEY1X7Jgh6omeH6JdSTQ0RuyhbyS+fe7a
Pf+Fvqrl3bPt+UvZNlpXUqZbnuhtwteQYzUhgzavveIyDxtHgtOFUJjb64IwO66G
mglODPfwoXwbADwjZ1boGhzhyjhjUqfUiN4/ojIRLJfbga4cL+e8t9O6F2Ad7w3G
JnsY08JvN0XKUEG7VbhyE0FSBs7MWA2uMVyOE7MUIaHE0/Ic9jbHP/viUP40bZRh
2t80vnRVdc8/7vNkQ0F2R1UcM0sfAilAs1Lv/RDlHF0vXsI9bGVZG2457FzxYlt3
Zzs+jRDwnNsY4cHKvwxS4mQPULU0BeLoDAuZor5u+2pB51n1SjImlaLAiSZpa5t2
5qVkdsPC05p/FaLsbffyohLjvBD1gJ5+MJ/D+wk6u6EBjlUmisfgECWw5CbSJ0da
F17LGeE/F/qrk+sKBPy1pTG7cX3eMqlVnWUxzIIlbNF4mxqkpDa2NotmwFhUp6Na
6k6JwLP4W3hwe52WwFFXHD2KafEVlKhJ1ghFd7m8o1lHw2RGQawYCx/bRBGS5EHb
V3MZ98lBrdRdUSt1Rzu2B0akQp8/NH/pNaGZBM8AqwDqh39SUFoaca/+AHhlyYCD
taoMH6q2hkJVe7ri2NvR6bh2QojpaK2YTcXtvLizcQzXCflzwtSMY2ougGtlim00
kQ0KyJh41BzmKrcmdQxm7CUFZRcojjNxb/sZduVpCVajjQnSipb5FlsWSlUaTPQs
ZVPq1h+scd2KOVALK84Mg1LmAU9sR2PAcNCkNledLvEa0j7iF/nYv1jSitk2rXMv
yMqleGSIJuCWGkVkxYkQaqrWPIl31CvaDXpqP1h3S+3Fnyu+OpMe+zm9EDtuJsJJ
nPxs5s7veEYCKNRCZRAtrSyxyFGiNtB2YWx1MkwOJG3Wgw4jx9NIEMJYFY1YaSu/
ygj+W+A2LgvOKh3zHk+XnI94JK7FWDhDXr3COjnJS/996qhM0RWsoz335vee14ho
ftccP0t2WCemNZWPTO2tnAJHU68TNMi9tZKAugXQ8pP+Pca+TL/n3yoRq6u/NoYS
Idm0pqK4psoE3SZlO9G44gGmTdKkIBj2SI7Sc/sWQkUO/Nm5KBI3VO1rTvw8OmCg
k32Kv+HCWjyqyOpgSVgbh5ifsaL2DCBR0lqiMu6i0Y778QbK/C504HM1FjsAiTrK
sYa+XtQbXoA/sn1Xmh5eH1DxP8R2WsgU7UwtnwsOa8hC2viYtTZ4qB4/+Wq3rUZj
kWr47eVG0tcUoghlXwF3kKMmkIKXkkLuv8IQ+0nu5xqbuDWvkq88IjbVCUidVS1o
FMQE5UlQg2AgxQXUide5cS6Rl3pOdRiDnSW3tvG1/rc+L82VJMWBLAJSNkwJu4cI
nq3moGVk7BxMhttrEntEli/SrZk0oQQl0MpTSQaQXz7Hu2kVoaI7u6snIWoUDP22
tTj39oXP4xg8qzAaQp6ZwrmT/igr+Id8bU7ztVNgcgzvMftzj8W74CpFxcxbAaD0
cgLNO9xZxw7o5pFPw+hi0YTZnOlkyigMt29TAg711LqRIMuaxW/YMb1wUnQQ2yh3
SKA9/Gc7TmJj674oV8IQLTgvmilpRI5QMWbCmsz+STrgxeyFT8zO+U43DjvRWfH0
VtUxNfn7/NtvZos4+Rf+qzSk2tU6xpv+w0y0/JCdjaaL0n7IJ2r/OTgfngbn3Ghu
58d54hbm/AA6SxY3s1iMPnwxKJB2BoAz58Uy335LHGBrha66E/FY8TvlHAZp/yL+
Pc+9puEA8u9K3/ko4DuESAhqCQwD/svHlhJJlyxOiztvuZvDTUsj/NSAgom+DCjT
VUGk3ktYNg78xLAimE+pGa3ANHfTxo31H6icsQsrTozg0PBfUvuD+r9gvzLCn300
idMNxui0++2ZE22oye1hYHJxLVxbpSF1+QnIDoIsax/9NF/PodwvZzKdoyt3Tsi8
+iKmK0u2yWAjQeOtAcrpPlFQnJ/r2qQpq8Y0Kfala5pLFH2N3+tNDqgH9m9ej0SW
F7LH6gaL6ftYivuxQB6wHmJfSGnr9TzSp8k4e+09pOT2/oEQdUFxaxcGJi/ixU//
r/xF2s+T4VHujkifxQpK4CE0SqdHwTkctA9H7QKZqhRgcel9JY21ojzMKSLDNA+D
HjGCoLDN5tml9800hmkX8DwwEhwD7G7m/qBCtRzShZy5VsMMeXvjlBW2jg5tHA9B
loSBghyMKI93ogBBvdRwqIUQVTyaE7UqEIBw12eqoTVwhkEXqfD17uo1xHd3EY25
T9xZYsQJtrU4N/nDFHeFVqEVq6Gm00bkkEyRasnmLBVK5V3kxlBaUfAzYo9gEU/7
bA+JtRK7fMPnXxuL4Q29aPVyFENpgSTBntn9rOIjzjBmovjaYR9a9NMUsq47U/Tt
aebY5T8ie6Fi+zaaUTK5GjY9M1cK3TZNA0NwmKvdKdfHtFF1FibfkxgU6hy6uTM7
wKigxAw/kObnxIKTXKAXMz129H2/mnu0ekf1ZauUJ1eQTWrR7XB7wdexQTY8pb4D
r7V6W/ppMEycdXetJ4BSvm5QQa127ZmENYuwCSmuTTlKR8OJrHV+7WpAyXv9oAy/
/qrpEJ0a4SLq0AZWrxIvYzmk3GZQEmtUCIKvd6rlKZ7SVqOEmnROa/KotuZWachv
3+UruG6deCgJSJVQsI+Yz5srtJ92604n2CmqXms0Ufrz9hcko5tslM+n0+fcCMwD
AIrIsuS1s93qkhvbDEAMU7X7Zkg9G3x8iO2Jg7W9AuiVOkeSQAHEf4zMXQ90ubRh
V3I+/iVR5y+TrETfqaqKMvkUgj6Lu/F4KSkzJ+wHxvDkSwF29pm64+wRU2LzuZy9
2k7EJ3oTvZp/zM2nzOMCT2UiERewz/iNBjO6jiuJQmDQiv9KZJUbjeJhN4lLqM0A
S+t6M+xF86dx4SlbEzcsqklVgv07GF8LBJfaylIhcvS16pe1nMjhXdIUCo+iRE4p
nIQvCx1c6HeemN/Ou2UchjuODS8HoB6xj6U61RwfjiZO3Kj5C7aeXjiBQEYCctxg
0iuCsMay7n2U6XBfanv7h6bPQfsKNjkSs45cjplooq+uWg5NKB6f2wXr7deDzV25
BQb408MDogGesyOMDPpyekvg989/2oiO7xy5MC2yPh6b9kXazs2mct1Vs3q0NiBW
7d6kQZcx4im9J3Y6wdj4Cpy+k2srgReOgNOZyDFdjkK2PQUt7hLR+VDbwud7n040
lrJJpvZ6ehjTfbaS2s60Q+jjnF8he/eb9Tt3jXj6lxf/N3UE2HHmUc8dWKjIpBWG
DGCsgYs/+uGGiO5zOoHOGjfn+grnR33FseFlXMJMVntlzvkbRiMEClbe7pdqCWEv
4gjIVu5OcHWaEZ/CArAOoET8M+ZX8LqIKy5ZBErfknLwzuD+0PNCpm/JLxCibpGz
P6lw0MWRqs+hvltl4Irov4wucEo2JS5jhUMNKrKBCRAHiZFT+oxO4n2QFWGXvVum
3vm4FYEY2FWosc/OIM8uP59rkPdPus2+tlVUGDgnHs1M+Ukgirlv20RrjbO1exXA
Ce03XXa5/EoqRWDWWl/yRUJiXiefBu/dSw7SUe8gVlInAoNMqSFOUKVlkABdGB/O
EnuUJOcJmLNPXKKHRfcgCJOPSI0hZHYZi7IPk++icBFpCTn+VxjptOoYCwK2GOJD
M0CsoG9GxItb9GSVgWbJ4lI4iGfkPNBoEu/wtUm1aKMh2oYRhSMdQ2j6Va6GzDva
gKrGh66kt8YNbuRMJm/MQjjjbajWYdDmfbOVaku0/x0ZBIWalxb6lQU6syfkG0HC
63I7Dl3iAA8lXFpURj1ukKCtVjS86tJYtQYqoCcyeqLXRs77tYZ85u4IoAtnvh2B
dj3IgXXVimAUMB5WDbJmI0nKWsIeqvj9YpCl25Jn3oQf+gRLfmYKEQfVHJmN5rkv
DAApcC0YrZsI5nREpOKowLyUAJS7Qu97HiSkP71tRUL5gZDCw0S9Dzly8+pfUAC+
r0jtXDvHsCC0Bqi3S3Ns0lpenDGVbn7cd1SCNuwQ592lgbO5L7mqJy3r/pQiONE2
9TQdBljhP6isG4H7yhcWSq6K7u5pa2boTKEjytk4vgQVwsUKe9A2N1peXbFYN1cq
uG7xiYWNupv3yFlMqDAIrdBSHMYe/0BMesaED5DN+mypWzhrnGlwsUrY7atYYvih
JkNvCaGVJQDcGA1S6/GL6QFH1jnGcXPVcOqHLCsu9udRleycWlbmyw3cXCfA2jUB
P/73nQvxCtL98Fjki1EupU5zi3Y3dQfqleJI0MsiKbPoXXGTPBOCHkDqBkUbBICg
I6bFAPQ4TyD+5BV1BCJl3ML/F0LkmXBh0c+aJxVV8EX6EC9f9SSfcYgUF1loF4XL
OP2EQH33Tq4TdjfInD2iX2fs/8fuIfuK+yegST588+qShflCnJg6WTfwviryWqil
5fwS1fIhK5j6wqzR29Ne+6vbHyqOicTMERcgYD/ext8DhD63lhVwo3TCr14rcHCa
1CpKuz6UDRzyxfaDh7ElnwuxIa0klQRb8cu6PO57TvbO+xtHTXeeyiTVxWYHjgRK
co250PSK/aLpOrx/HUn4sdlueI11bs7W1keyCCul/a0z9voKnCJGCgH6hsKPibF0
vj9nN+YqJW7OlEuUMHUze9PONFbT1uCGxwYGxQ3vYtQge10kjVXVaFicugUNSTiu
CnhVtuve6VDwUYaZhIWpKOtSvtwJC+zIz1AtBy2c17BhKbxTLccZXweJZFjeB3MU
zguad8J52td7ucllrekizxVseESOb6YCnwHUug8KaJYZgkjaNrQqgY0NmW9tmYzG
BNxYTltYVeZeW5Zy5y80+9ciyAw3pu/L4JJ3RHJhamnnd0UMIuLRCBiyN5e/2DW7
5nhSHjUGCN1DDHqg5qku6H4FHmbCF80aEWtg3cX0EwnMAyR/5x/77O+ljAOVgpHt
jFUWfJJ9iMCwQKinDJE0/FnUy8lu0v7f1jsu3vZ7e34bJL3oIsLtdPUhskF0tmKv
X9GDHNDeEhIh3P2luGn5k+QDAdpy04x07RhkEOAsrpxAwiY6msLJ8+M610tRTF+L
A4l1B9l1LTDiCslutrWtwdUcS82VfShszYYA4LRFZzFaYl8aM2DLkVqGCKKtLszs
dE308eG041ojiWNFPmnODiABCx/lJEpu40ULr9DjJxAExYwKTkPAz1KScIVVoBgR
EgHdpjo7oTIrdrjzcO3i2ZZqLzigTpq1/wYasRwzz7Kt83Q+/N/zY42Ho9rFj1I7
Glw3oYybTZJcuH7fk9aAxu1E8Z8wN8DuRX6LdRvvqSs5ULv6P6wy+0/1lvcE1gAF
waJ6+10APuaqSwhPvb0wZpZoMfcGGzNlJ9ktap2e5I4dFzklRwhqLckN1tHsWp+t
DJuL3ZpaOz9cLR/whkJlYjO5Ju2vkpRgMPvICtatR4cvArtBfrjUxofpDuXsVNLK
B4Gl9Gya7df6P024uz/zT4uSzNyzRCGtSm7tvo11lTHqSeuIdjuAjvvxLeLtIChY
joCbBOUfXf1tnDYWmoTa32AVZuOQfZnT6/hvpeMBzbC2EZCDG1rVdKGDmGo+b7Cx
ZS6DqqysiSBI19OzHJvq3rMhCgPcEF9enWtqUyHM5Y3szVLknkBl1q2uO1JzR6O1
piQWTewjpXZ5tZ5qPec64ndo4+bS3LS9DiDPpBqVRAJGO1tzVpTWkZ6NknTg1jCC
AXT92Xxala2DhlN9QQn6/ACdZICGIKmV4K2RSnxXXc+IqkbhjKEwK+iiswdBufN2
FS5YrWZeWpzrez4UQEkWfPOZk8NwvemGS/7PK4fwhs7LzmGnAWUfx4MVrZZbZ0AM
jjSYNxkA7iQZmuoDGQuWkOrKpoy7oWuynjVX7bEvNnegKKnokSpu/n46DkQzqQlh
rJK5Io4GtPj0gtpvN4qWerQreN771UlGvdZI/cx1x3pqyY4NmQYVVAlPWBv6NO1K
v6FVizfs1Y+Q45TFpWxjcKAFwdRv4/94oNIn59sb2jFCjPey2/AHkivv2PZZSSaR
vBFB5ozEOAINNMMW6n1YNQzl2pEPySBTnI9bBfO/jMrXFlYj88224RjpiTwbhO1M
qrakaVG/4WSLxxHYyzlSH78mtvpnOV8Agzo9ffUBEUwIce5G7BFa6koTXJhMHAaI
k6gaHIfQyHSY+H/ytCUel7s0DVdNv5h7iH8uyRyq2c4hyJQ8VxVMHnEj0xi9R9mK
JTQZpH86Eno3R6dX/LNATh+A01Do9AhCJnF526q+fge2E5tUM5m0MJT7CQXnV1qo
ii32ge1STI34szLB/CvcTWYFDYilWQkf3zT5F270quUHBqAQiR4qV0ECYVEDQz1k
+wgcA+Wi91AegaKsaIkdVREVVrA4IbKkE4YgMCG2M4+e1yq27IGxrhIABGSudvDM
Fu+rEGbKfO1F14Y6k+IWHPwKN9yAYt3/fR2wfIee3okivCtT/SNUkgQmEj+GPCS1
EMswwfN6CsMB85LKTIxC+9C/Q/4zkv7EXUVlXT4A89N2N/nkAMQhM5PimJR2PtWk
XFbUsjOdYOscniD15sK3lwIZEXMxG19gaaAVE4hkzfDn0c6Pg7JiLhSnmZNMGfyj
e5Eoi96KQDRiClZEIZVT0+0sREIsCaEV7HLcTy4KP/nTv8DK7f5HNri4QxKmZRlp
oQq/t0QShkNqcg1WesxwPFLbmz+EdBJgwiJwtBbW1fxQnpJHDixhqwI2Bs7hRXzr
9hoCNl3Ba4ZjOa02qOKozUNYfHZv6j8dyHEwsYw6Iqi8psUaSgtxgYh05Np5kujo
fehC1FWQx3aD0nIctEVZMZoLF6Ntop3nIeApoflLAdmC+vONk+PetVlNHZJ9V0aO
4Q0JaVXY4E0IbQz9VBGP7U8mX+Sq4u4K2PvLwtY1/pDYeube4nl92771Ey0QiPxD
ERDJPl7P7W3nsWzJwcI78GoFZ0Ovlv3CzhXxl62I722I8Lv7ORqWuJVmRFJq0Yvx
ppJVRB0kIttw2sM4zdrDbEyD9KQgf+dv8jO5Nru6rPDQF3HSPtFcV3ts1SAiWvbJ
jaYIPqTGBlJklffAsNgHakou7cbRPKt9hohylKbpdYeZ4bkxiXiOEmAAO75U9UCh
iyDFS62sm6bH3K/HODOfwXum518UbjXbm6KA/s+HRx83DoyHfJiphJ9UIibw7o50
8KsSx/KatB9rmqb5PRB35yyWgcFYJ0+B46LGiwUkpGt28XxGn1TAGWpqibIPDJk+
xEcCYcmRg3w3a3W8tXhZTsMKEtl4668xeb1/nE4+Baa71JLdoqrxqE9q4hQ8T/2W
FFIPTkz7vG+qea2HL40ikmmxCeQ6y+oKZps7pUTwCUq+bGwVkCSD8DcIym0GgOgq
mPmLYFNmN3DrJTFxCbTnnq+P2kZV0CIEAW+Fo7Lin65zLRWOM9ibFWzRm4V2mSOH
Un7wgsjSW4NUtbpmTconEXez/JEEf8oS3R5ufNw1MhiLA4nSBgsUX2MR2LJNlfxY
GtOmI7Jn7zyjv5ZCnJv66/rvsxKyI+EbyFiY14mNItrnZstv+AaYgbgstp1L21iF
MkV5w4/Xw+biKeNXvMgmiai0669btQ9HhNoXkDtWorkjaiQDkjsmRNVNjYgbq8Gu
MXlHuLkvIhnB6oHZjU5PXjfNHXVEsYYO+PfbhlXdNza0rLCINpgLykDMIxnS9Ex/
FaOiQcDTbPa8lOTrqJrIvCZeM1lYKPobmCzDcVSvBN5KClAEFcHBSOTYJ0Zu8vqr
bMtGl/ys5kZsNV6H5yl2FjLtI2aMOsnYJgaFtaJJ3jb9RJ5l6D09UXMXQ13GSRfg
NRjvBRtq4DDPnpfGsufq47ohWXFfzYTzw+z+Fui6BM/QcB5xlNI3GmTzpEjatgsR
JtyK/BSlX625SWH0EKIwYFQVrz+JuD+tbe+2+C4Jft5USuE2ebBEnCANLPRafwh3
kPAuGf2u0S2rrAkpQ4JN/1VYcw0S2x/gbxohfxK0iDTNAHNuk1gy3KPPh+J/RYZw
UXTD4sOxNQPTt5hsPvkdOARuB97ud2QWdMYh8SWDe3vurbDi4YEcjNdOQsk/5gsY
UvD7HxR/kmAfdH/4broT/7X8WZJKTirpGZV4M2fL4PltdQyk1bBlUd9k6tddKm+f
zcnlB5nUy0zhZEEdDS7x3Qr1FSiNLQ3jQ7MyWuhav324UNy/yfnnX1xfqfGR3RDm
UJHq0BBjRCj59dX/LvhdkRU0H3q//guFVqM+s1o1SG7GFOP8skxo3x1s8bHcm0cM
tSczNBHWQsUsMNI6FTvwHpki+qP2RyHHH+NMacbiXuFdsoQ/7gIqaADcNfErLxzc
ZC6DRr59DaGbAWZytHuoJ4ndHOl/G5fUryGqTZpfHe8izhxS+dZeIkeSF6SEfytH
H6fMWDC9abcHE/D43LIuT/XAoxAT037LGqpt1qw4tNU+0WzOx8sqkA8fTF37xbul
K7dSY+4ZuhNCSyJ4qDlryhamxoFpWvRPm/JdWvkdeazY1tKDviNy2MxCnAR3QTNT
2BJj+2drtlhHSoJd3ih6+Ab9oA/DJFwpzBzg3SaJ1tno8kRNFyFmDIwELJiB4V/c
boCAl2ysxp14W9GyXmW3u0rIxj63JhV5k9GOk/3POpEawTA87U9Cca2GSMyUOJcd
7hddGg+ZH2VlVQOJobEmIUImi/aKcZZOC+iHmP03UIvgoQ0X2GGQKzYe1hjd0mF0
reWP6WFI9jiZ/kx1bUrg+uCFieuazJ4AbIpwdv85hu2HJs/dmOkePpUoKrJvJeBP
fsFsbr+vDOq4MWm0oPQ6bhTOcfnfflH5obtwFBHROr7YqUddUbGQl6eddpdMVzJ9
kMluffGv39pfUhODMocOViktIdCJ3uPjoMpWUylu9yb3gzRVDsGs4vPwdf59PxXP
7Gf2LExyQL8RAV4IjqoBN8nKa1Y49SrlDZDFfAcANW9e4+3Vve2fv8Qdkkv+IbX1
B548D3Vdr+8WEyH4uLaoq8hfQMKN0oAw942QEaKGFqUlddWqqt/ng1KFn52z8/OI
AenXdofVOEaBW4CIt14ZGwPCv+V/Tanane7X0py2sY9mjyWBIbry9ctnAPeABGFX
XQbtZ+d7VZPmGfxUt5JEJMo1lAORhmRoqWIWUosEgdGPjiD3zSIVX2w2PQnhZJss
Yu3tSHVH49bPu8PrkzZeY/GSpw0lynw48wVzom+EaITvGKyDo43AB8Id8vJ5eRah
XULKBAoqBb3Sb99HtXNlSFpR5/xVlC6sOF0yJvglyTcff+39Q1n3zCwC5u5dkACX
HdTIr6L2C5gpvkpO8MD5B+6ZwyHd+uZKSS+sI6YKtJubi+FjQf6EyYxDFbYkc5RW
C/rCnc5Obcie4Hs20wCaWo5JzVV0X0YMo3i+22US7WshX38tUcLrEd00Yaj0dQX3
SrgiQOWziqgSXgjDVsUt3dYrjcDLExGlLw2Bme7M/3y/bF27DjSrnOEW48k1uIWA
P88K1knsjCQEmzd2w+sD68+/gT4IX0jvmv0jwPSYVx3Hv+Z1oGEMIcOByGOWao+N
fK032eGbK2YkwjJ0NdoZBXY8WNf/QU7m9zRVSMOm3RrLYmSUUrTKVRhesHcIqBHg
b+6BDcdB9wBDUUs1r43RcKtUCUpwRZQyQK5FodDQvXltCEndwNbIUpJXhHQyxti1
xGWJSXEXf3Ru1RVuWRzGaw2I5yNfU7MaYi4GUAMbUunOncakCm4iOIrJtTDLII7e
WYd7tKuABcz12DMER16Sk1PSsLWb/N/0PcAp4OLONVt2Cfl/0+ppQMrRjuvrCpL/
Lvukvyb8db9OBJ8Fc70GsYHKAKXQ+jC5coUqRm10/RM+JuFDSqJTB1LK5LuqhFpB
w0ppmOvLerElTFj/bc3dIhBfFBPex4IN9OKjP8mFJmwgVpZljXdoIei0HCygKMLU
ywdmExAURRAWmJaTC+CFQas0B7zn3W7RCeT9xmP38yKTUPhHw7d70cfvF6jPavdg
WSOMvb5oU6CIC3tTgRE3U1t/X1gZGFk1cp7CS5LY3ymCOs6UC15Bnm1Ur/pbb1Kg
jBQb2Perf/qlsVpUUR4/puoCfdt3JJBclXQNI3aYGEoHTPHtMPRJxG7bSHZHZj6b
9kq7qcL90tMcTypH7bfN3dkorDQGovtucDysQWbOS7OyyY6un25omGvD52Kev6TY
WonR8zEkHw7tlLAylqchdYl4muZwTh4iAxfmC0aoViJcIwJe3UYzXFBYIR4DuEdv
TzUGhXi3HYXY3jTLbmxTuPuD9d+uY+TM8mNw+H2b8wuTKKGEoadbUKtXeX4zKwdD
yUn28UHbVlT0W0qHtcKdfnf1YqmUHwTIx+aYnAGSpDx3TAmLy8MIg4+ao5+JN4Sa
MMZ3YXGYcqhEUkNIFamxfY4mCwe6JzFcuJQEr+7PGeXCuuUcpk6N2giQKOPPUR5P
EeAJkQe68+4C4ZU9ktlI7oVNzv6r2WeJvj4sHsb9tXiHYDWqaACdnULfkIFpeIgU
Kg354jepWSYiZu4Gg0+PNEYIkdDMWo9nnJitfRiDfgNBNdLCV8HtAi5mVIH/aWxa
BU69Tn1nXl5e/PxkuEH9kFXieu9IkMNivHeZK4lFWkHwJrOHW3vXJHGKvZYV8TOc
66iV4gnbYSLSOIxgVJ9bluaqNwFySofvAZSXhKH7Ip473ES8/MiteUYdPhdMEXtH
oFBAPDZrr6h35YEbtobuWJsRZJkwc1elb+RSE682kyrgLpYsDTsE26HWe0vFwkRD
1NnxALiAMe4RekKQvEloc6xSH/9XLjTl4mikCe8+zOReNFWIg2gWZ2ztbwEQmV86
nTFxzfNdNaFgcsyp2J/liuTHIty2u40D1BV94rfIa9Nvkl2OUsICo7LDxXJJUSIL
i3mTT3931AzUr2O78cTJoWlVRuVQ1vAq36xaU9Z4QHuBadr5L0gF/AFN8i4IhcpW
K96kM9uxkzvb5MWNb52+I4hhA7w53glwDBclivb1IZF3VRUiqxRPl2nCA/4vv7pp
saB2aNOahFeJShsSZ4vJ9rl3XFwZw8stYE6d3GTFBtsmiiBVrf9N55724URwarXe
NwfkCvaHTAO9yKmIQkpR6fKg3QUPj8wfop2E/Ncgf4cP86VqDBQXg8QoethQgfD6
ds1FKcIClzGXGONFcVPvufzclMy2SklBeLx9yxJQjEJoFuTAFqUQkBIWTmfI3IwH
/bxVf5UUUEpq5PrTz7Wu1Bdozkh04zzxBHMWQQeAzPpFD1TWLrGGUZeyTXaWjTez
uC69iU4zS+ccQCU/vocU1gmqf17i8R+8idSTdlovV09q/EKDwBd0Y4vaVeR5UYCa
iBx4DA7CGc+dCxk4LV4tdQjb3mkJ+Fc0vkkWOs6iHm1gTtUPqVUjOedbyAsOyXQ6
0f/qRBMMEivsQTQip2Fa6dBtxxt3JVT/+QFasiscG0k6z/VlnaocG6Zbb61+r/O6
KzevlH9taVoGNRXzYi1/Gz+rIwWG4836d+0MIdpr7uUQHz1qY2rR9p3OuvvWlQCW
EgSUPl38B0X4P5P6ZbULtK5Q95S9cmUOUihUz51qOcxDOIQHI5YLCMqs7VoO3/xY
VT8IHQ8qRRW5bUwjDhaxdhUrQIKN96aR2kdG4LHz99CcUwmbCwE1lXa2yd96seF8
LwbwcQv5a0p7/VgXdlEaF3U7jpWqsqoHh+9bLASr95tQpZ8QA9CB1JoAMSljm7lO
pov98htTbYVUWJkcCiQxA/Nfgz1wNJq6RgmNDADKrCjJAuopIzZzypPnimaARTXp
a7vqP2D2aavDJdrT0uV5pfJlDPyWMGBI2peqykl6GOXPiQD3Y3cXR6kViSmwtwEK
u8FNcaO52PdoTEsytyn9MfnPS0o5G8bijAsAfsoxFeA2jcq9LJBNcoaKQl5p/I5v
DCskxqDet9WOyjw1DPzvaGVyYmOZEm989nf73DeFoWg3yjwZ3H5EPcMd/EFCuji8
i7t+ENVq9JruRWgv41h2Xf0LKfIYkJKe4qtMtcOY45u66qYEiWp6SVkjapT2YXJf
q5aCsgvgtgQWH8cbQPUNm/n1KoYcjRNWhS7FbfRqXW4mSzEDBQ+I1aBtbZbdzCqq
+ZFWW+HVqawMRUkGCf1YxN4NAwe7iFHSq+JbWdwW2ZiDoikUqWrtZcNvhrw7zHOx
yVzTrYlE9nxbNy6QGX5Q7HtL8G2mtXAGUu3uBXeBXkiYSoUz/9OKSwyVzT+SDmxQ
Q2VUnd3+9+P7qo3PlRAcZ87ufOChix8S22UZIDcUbV3g0eljrcDPjQcXmwp3w0M7
bVAxW6OZjyUCpUwSEnBkyURWoKkPNXiDQrql7lF5Pg9bQu2U8jEqlR4N5PprsrH8
SKAVf9c6rY+yL/p9GNqArhdRmCzBReQ11ieDfCRIsACFwpENXr8lO2yzNbjrRPLx
XKtRIQqLxoY4l1TJUn4iLsBUacKzaiGKB5ahB39baI4FlgtokhZKtVi/4colNlmv
plCNIEL8zwUqVUhSiiSsNbQ9aUwXpGESIq3wI2XFNuMRPu5GlLW6Z5MmWJjx0rnl
C3J68HKfem8CdZ0APbsegmGQeBjyoN89xF01bKxQQF3ji4bDg/ToXxktbE0quEML
yZO0jmO0v5fpZWov0RX8joIgGQslKXXhE2e/UPSBLAEOEAFb8wU4eZsJqCkHg36W
ul3Ua5w3PcW6TLrRqoraRoV52+Ua+PAR3PSNNBVUpRYW8q2YZGznglEP26pgOK3w
PL3sOdCcIWB/Me9whF37ZjD8RzwrhVhNa4ibm9ALDGtNkPU0+il5swunVkR7BrFR
7ULNBBpgEYXgyJzS58K14JOuYxYI8kbj3VFkPLRyuHz+nOyqzahcf2S3n05gn/IW
wYryAAm+z/d9GzycxLcbpwg2DyvylLSIQ3ErbFlXz0E77zcL7icmZoO2okpttV6g
+rK2ezj7CIfIq14l5GAuMEOetqxesm+uAJaTie4ud5Gw1EGQaNvhFhjH3eATVkN/
6w4fbzgumIEQ0XbBw/DwlQ2y8ys+w85IoVhGGpC6Vziu+kF6E2Hzzkwa6HJHR/AO
DlvoDO5CJuDy70Nvir/Ju+oN9m5Cr29Aa9yWDIBY2ii83u7DH8eCdHYDojy5qAQx
gPvJDhwXrNNgt+sUYiKGddy6voqkxP5fV8RhCyYfAka4ZdeNBRgd4ipzNjQyJ496
AoGscKFZpOyG6vusB3jqFjcfpAAMsjeAivarJAgfbSsRGq++GNeZNqpNjPShv/qb
eX/1W0pABVME1TCC1fwtk6hFce5DPadIvqhm28cntEhqwWaCIGSKjbVV6JQbgjmJ
10bW1wn5dUpaU/JYnyBsenS/fIgFPKPNO8urFKriU4JRg72gF0icOmz6AHBhuKux
qo0L0QB0poT/XcuJkL+k7CSCdI8BNLg7TX7bSeQkD+SwehQGUdowqIhBAqUqCfoB
waLfZDgCPiQtnYikZxi5E+9IUT1suzs09Dn7hDpGyhR2Qi1HOS/oGwY09KxPRvEB
YHMqHoNe5AJLJQj7lnj7npDzVkozsp1BTGVPackHZArwywz4q7tDPkA9S+++lieX
x3ikOibhcgmFnP/qy3XV+bY9xAFGx6NghGABCFHZ9cP9pnZ0VFHEbqJAPdsHblEG
u6Jo/lH660jv+eiKIDqpCXzua0I4Cg9iic6n88y213l5kCL2Jq8Fv5TsxytOko4f
5/HlXunvNPsw9/TMluOulQX+ZJbvJy81yUOEyE5ykWkZWeU9sKn0QoTQN12eIsZI
ajq0fB/9m6KroyaREHdrbdhZJv6sClCuV8AIslD1MmfDfTeUt8dV6o2UVGK9TZS4
P3eIfgoH7FGqmiANXhKHjC7wF0t74LZuJGY6BGqL1gJRX6ElIi2k1CBrqX4wTGEf
QZ2jVnhRQ3ufHcA7V4j6qz9DQky8W/FCz4A3NPOvRSVRliEXoRpjvrzEP5sP9Hzs
n6FHxvIl+8JY3OVYhs5nL6i67IORTrVoyt8qUdRCj9ByEG+XAz+tB6KfixDRlBbd
OX5YONyJEnC9jH5IIJIdqWF2sADZYddQoXReG3culfo2JedPvRMIsUY4b+nRJcdZ
X0YLxcj2629T09JEkz0XJfJG1smQVfWSNYTSf9gg6VSaqdwd46R/Xx0xmSKVWUpN
qelYIpsXufy1o54WnhoyPZW+iJnhNh41Ug7a7/G0rSb2nylrz/ZxsKkM8yaUVSxV
Y3hUnAthUpMsp1k3x4JOdwGSmhUm9pghtAs82WlXtTLhRahqxCIV5nLgF8Fve5Bl
MVmtto+PC5l7FyCAgmRHVZXPO/P5UToIm8AfGVyT1k7Lt/tydrnX9wecXOAEb5Cy
pbGHCDjynkIWANa1RS62EmBlku/eEiISZ1NIKb4RV25unNpp1nYOI2GY+Y3U1EZu
ftKHTfxL4ZYYjfl0C56fB9p57i3dzrJocDtu3kZwuWKS0TbV3AnxgAevMRPrL4oI
FKGROTB3J7BVRBxwuPgozZd4RM6j/eWGAvV1U6EEUxUjf7JE/nw+wyl09D02d58w
Go8OJGjkVsqdhb7EKTo5Tyd3/rZXqcuEQVdc6yxj/ZxjQDsEL8yFIBL1btwj/wJc
VR7c9C0W7IP2TibkGLQ6us9q7aWrcv+o8JK7Tjhls+IZKIM8kLmo/hzKVd3gIi22
lkcQkzHpwSZOyFynOYFe2UsU93bb5w93xyzrfzue8fzL5KmfRAfS09Rp5q1Lo2lG
8kgcHJ7PTD/O3An5wCc+wMWZ6hsVU7zJtIyQCh3jhW0AlcdDGOkT2cnoTh9bG038
bEWy0Lc4p+s+cXP7LkTZrQyTXtc7hzsNIk0PrxWuKy4vdv2hIf4X8iSH6kC+qxus
OcBEgc6vrX4MUgRShX+cP2udjE35zPpFGnz3XWK6nju+tIdZgVrFUSdIo3zgIgCs
sIW0rJ3OmoPcqsSoRSnhEwv5eqcmPnBIhjOCkczu2d3uJ0IryNlhVdsWtlTi+/HR
GNwebEXdtz6kVGUKP7zocV08eiDOLYqpTEaTuUGVfNyO9cxUw6xPSNdUTijHvHB8
Yc93KZjP8HQ3BjJJbnGZ5P93r/ZkS9yzVrPeKzaXIGBOnjYSictZSGScQTOP2gZE
ltUFnzX4fs7daKE4oskg1xQnPkK2XzZtcL7r0f6lfrNwof+VPJRXZngII5TdIlfJ
ZS/k/uhrgfPcisR70WljnSEQuIX6cdqy1rr4zcMPBdYVyaMy9gMQlx6oObcB+wqY
qifBdw1ftvJVZ/TKZWnfURKd0La1HfiuDfe56/qUIqLjiSvAZjbpSUB08p4fxypf
vrvFDD7MIQjHiJNtOXXCLk4Go/Izw6yHjaBMSInTirI0w548AstzXx5LjHFEHxE6
jCZqjF1BulACE7jR6i3weCvMX4G2nZtSXi6VvpzDhtUa83BjL/CBwcZvgRa7xd83
J0xaHiLwqovMl20YlBYNUcSQlcsSR6uSa/d1ZkXZF8Wzg6YcFNYpg1ZzQj4n0TsI
ahEtkdbNLkSdABYb4MGVMvaEQ/Udi7mJQzVk15PlrYLmmj+25vLB9wyIkvehJ3Fa
ppaDHySkwJTJ4svvT/41IHJ9CRAWKg9LEEfES5NwydGPO2ZMAIV+Jkf5RIb5n6Id
DeXrdgCyHVBas9gqPtm/KJdAbp0RAU8Rx5vq88ee1jX1r+4IpDu8PNI7iQCUFuBU
eVbRAvmBDKeSiDPShcUSFrbRMv2462QglukLnRON7H8vqZayZq4BtkxyaJWTIq5l
1pf314/S3LVJmF6jPqgitfsOgNmYS4HRXZUD92ybpkYh/qcdY9DyLfrXU3fjFY0b
qQpt9V1yD1ekZ/uQYOTfWF1xR34/xamuHBm+jEjprqPdabwHeVXzmp+/47iDnFa8
LoHEW+BzS9bZP7wHjtyieSU9yvP1QL4tfmXM4K2C0fzLHL29RuOJ8GEuA54vKt1K
b3BOe4c4JfwlJufvhorRECM9ugBhMdGC8d/iWWtj35gxChbWUuk6jINmvLmPTBtE
gEfzqWPW/GVkPESQHRLkr7ykRli0O4RZtUkOIwgIH1+HAAyPtDVEuEf+lxdTQ+8C
gvECRqKH0l93cu/5Fqmn4OR8LYRw0xXj1OqJsuOKdGgntU/8I7rjZTe9PSGKkOjN
pvPeSjrXgwlxEV9NEnP1EWR6NAS43m9e01W2SgpZNLQHmreA+rsrVc+AP4Ck1xP2
Dm6Ez19ePtMuYxBGg8AXL7eo+H4BwZOipwNkGX20W69FD49+q6LEePdxj3HVdjeN
0wofWlb+CXKK1HHrz222a0CZa7qJA03UFeKX5k/tRhVB4SyNLtjWPpm9tPQbPaqV
++pS7ZYG5juKra5b8HIPCjTjgldz7T6pUZhykUnFJ4Vb1zHM4tpvSNr876H55hYn
mVknCotrHhn414dxETvO+R9X+tWouJy4sQtBoasgGQ0e/sKJJD96Xo/DKbIWHDRY
OOLeSIQA+5COCEfCjAR8/HtYMLvBE56f+8VVmhM4j+ZHpjNyuazZJbtSiDZgkq1f
xkpM9jPD7PLvkfYWLjYQkiQx5PA32K7XMOLZP2kA131lI3Ecu+TDrlHnBEpn+OLD
r9EYHKXVpzJg+0i3157C3mhd+YritQAIx4vUXcac0sArEZtaJ5UzdpWztCzWmRU2
8GrJu+D2NNa+UK/0XlheBSJAf1a9KyBI9isJoHuc3NcfxiDpGOz2C6xVbIXDzZZc
LkFa727GvP5bruHi4aKLauSxyoRTlzU42P2axfaAiEWJPV0l2lLvc7nzkgy03M++
EFI6nAqDx+TFX50dVw2GpbTO8yIEHqX766CUQe8/MPgvdRmrF2McxNxxupj9FZIh
GNRuxUSDdZlIHWYBcvsEfwMl6tv0hURK7vOqVEyyHhPIU0Zv/VTk1XweQTaF9Z1D
+9ykzKdHnMSAl/cvZxKKS3GR1JTynVUFknhqI+0f0moIpLq7oHF8AtlxJ95DbokL
OV069klSiLQcdXX1kWDa/Q8emQfjazt98IBqkkkGJUoQySMkaPtfB4sdFWj0bB+F
+3DZma7v3Nc/c8ZHvHQ7PsNVlUcqP0dFrpxWI2DRYWzR07yFSfZ8hrVHFzRc2SOw
6H6gv3//ocrLrspKt06/rqZvWdMUxE9Q9Gcgiz0quxqJ6Q7reElko4exZhO6HCg5
RlUY9QyQnLNi8von21TN447/xoY4oyUPGlruCCetnAKZ8WfSOhGn/kH1JkyvJ7PX
6lSRauS9OOh9foGEEFu2t7i4xDo4bDVHEswOhbG1ZFy6GwIChsuiIeto5EhWWeEK
yIjj+FQOWe1EVz97hOqcPEnjCSBEdeMbuQMBYHjDY/XrRUFUEGgQlyp3m0ml8UUe
fCH+OSKiWY9Gnql5K827vAmykr3rwSJOqGnxaXRqiy4r/0bG/jIJvDY4vm8qmEQh
QL2sPLJ0muKUMj6Av8x8TkeSoqdvddvKB6jP45r/dUh8sGj05NhQCAk/+7KaXyQU
1bmGiC7UfzaGx++Lc+R/xh05nesKPDM2yLz42DsS0+OYOq1XWnuorzazE7qvrtlY
AEMPbZSp1QnmqS5t0pzzg2vWLt3M59wl253bkZ2EQ5K3KDOS0ESovxF4rZ9+gaCo
e9ficXsTtfn1IwzWhkx8LN7PwOuNsseH2pVb0tVNhAaRh6aJEvQ+g55GqvuGwohO
9GlQiig9ZRkSw/EHocAwy03rPu9PCoWDalYmsfhQ3jPxm/9Wb7H5jt/NiWfAlvXA
oD9z6VY/wMsydUwE2MQNCp5QrqfrTsAGnnMfHXfk8N0jw5wjG18QVZZYWgtXKe5p
E+GjZSBm2zT+9hNVqXX3RVNrbb+UC6fPrxucFVVL8C7ndn5IA27WWhWHnq/WCk/+
4onHe1I/XDm7HM2Bk0JicOyZkWZC5J/8pY7D6VoObPVkn45cWcqNWtSz2qOcvyeg
BsyZVhzgGybsfxtG+JzCljh7Gf7hEmrVzLbe21mELzfyL8RXZ9FOocPPA48BMbKw
ThLePfVd4bTiqGQNn27I+MhQCTQy/1/W0JP4D4y6NItR9xLn/Tz35IkHegU6hTBo
ilNSOKB/0Jx3+p91Wnt36BdIfE+9uCRFHbNXxHkC9g4oJKxZOqVZdH8Ow5M3Cgxw
CqiW7en1aOJN0ciuHoV4aSFAaavt8K4TOstGcYs/S1TVQUsHURu3by3MVSJuBBUf
5Dtu2VrX7DN6CBV+956/raSK+rPVAea0EOHJH59LNRKe33/9wWILP6jrUTpejJTV
h1GOn0EgFQNYEUN7Bh/0RaFgMc5WUT9ABcoWx+N1XdwOXh1gfAhjljynHRYXMb6m
nHUbvHLo6yjosQ412vvUl9gQelVATiNAHY4k2Hrh9BJ97s3apCAd36oI7aJIg+8n
nbvSNPsD9VDxewbv9+5z7lE3LVNs7uUrpqvNJpRlkcFmPBJ4mhNZLRbqXMaDZZSO
VqHvQjlnLoa1c8tnDiK2VMvkVKkVSjvcjNkC86J3xMS/Md/S8BGHqNqJcN91HXQD
kFiQEcgcdMyjkXla1hSCkQ6cSvNGabprhw0vkjsvuzRNzn0k+Oe8bi9M+0384fk7
QxNkDkbQL4Vr+pBSeXaD7wEo5e4vhmjB02qJEbSvE7T17xL4G/wMALHlLgv5Q+if
0RW7b9J8m9YelVY7ygiPo7YABNJULp/DFqRo0ny1akardOHSldNF90zErAIm56Ro
rnWGGeSBziDYxlDso6bU2Zfg4E056lo9dOCp4k4cQ2Nddldrv+IwI0VvERCrsCMW
7Gg1YLPGRvq0GFgg76BdrFOEUz96/HMkgf6jyVQ6iSt+Gy15X775RvZglL7oJD6C
iIrSjMq4y1jc3sdmSDSL43TSMZx5F5CiSo7tKNBUjIOxe7liErnyn10IVasra2rH
UnNbK4VR4UAmXTjYeo3ykYy344LKb6N8JLhvmbqCsUMEQC227etvt6empEYmwnlE
qRnUyAFldFlXPwqQlJzo0UnY8xFo8OuV9mX9q/utYa29Ux20hQg2TG4REh/JbShW
as9UEazzBUmavQgU9hyHgkQHHsOGz58uwO+gxQiN1GNGL1KZtlw0HD1bvi7mITds
ae+sZkwGqquzX8DIlI68y55eIZdyEZt6+tb8XMo/9r35HnUHJCVsxoNcPdrXEbC0
5JIN3R8d7ZW6XdI7NFKioW31AF+FLu4TdE/Iy6/RCEJOGIkslJPuotSpqrHkGt2Y
F3OYDnM6gJyfCpVVkzxjwNUMNaNRm4umGJAJHWDQyc4B43faBb6QoMJRg7mTRraC
lPSe9gQd9ZHTfSq6pXlKiz2xlVmXVKC7pBIXUwl/iqD9u6wsDQJ5s5uhALiyMHfb
9xTyW3s1hzvfRcNpIRSgXb9l1V27+Exm9vyclActGwcWoywdo6FImY6FYkeiBmHI
WgSMZxZQXmy4lTSU78K5FSAgWgxt95rHesaBEJ9fABLrgrsjX1BBSyhwbCj6+Ke8
dr7uSDq3yB2A83/Jihp1uVU7sB7ukdFyQ14fiOY7s7NZk3Di0LgRj2vZg56wnAgy
ynQb/VFCsA06Kym8B06lDkIunIqyx7GX5F2cIdzAvvX+wfjCAq1eE/qRIybHYsfb
hRMUAjNU6oIQ244FcdNGeWczKpJu3Px97++gGgtvJlZi+WGt2ER8me1NgLwJNCAn
mImLRTgkJjilLwnE25zeMlp0QC//L4Wb6jQKt/JNJC+erdqa0Ith8Y6TmhgXOgep
B3icD8MMvQGXuaO3k19n+zPsDcNWCe7gzlTMbgTY4MAij40y+fyBMktwlAO27wEc
8CQASh9mPfFJHEpCt2+GpGe5N4pRJOjqimBCEZTYMEh32ymHJBgcphK2+2eOuyv8
xzwngTXMautT1zg+4EDIxEBbCHcjub9pQvxPQOradpfPPpmSIkXD69l9Ia9qxwEM
1FTwBs1s/R50qSBE7i3I5JOTb+ku1wjmeX/3oFz8w972ADskgmXVYmCjcyw/FadD
o5iCkQgTo4tBlsLXibHdqhfZXWMVDm0oPClJIwVPdj4jky0W76INZNjTrN6UXhCf
apXXSW4cjLri+K738rd/R1U6YgBiotOMreVW6UeMQarbmuuFAGtugNrGnnBoDnSx
2a2zsY8809mK9hIq5V+JZXk3YpyrDEW3eaJlyowT4+KqmoPl76vVXDt9Hfs+V1jo
T8kZ5SfAYDYT7L2FZHt80EZRpRwkt5jf9ZK6dW45OUqAmylbjZ4uViWqxld7k6qJ
eE6f3TgKCrWtHx405r7zpl3uDcYGOsA2CsCmxM3v9WvL+6oB6iOLs94AQN8MDUeH
DnU77baIAK8qqakaXZaecVOhIX8upOgeleVUuBUi3Nj7h8fmbHfReJ67/MEEWxZC
cHeeHv34uMWUJ9eU71U/X303+zcTAShq2oiGMNBWuGz2F+0CACDuJQq4YPWqApwj
XVRLV4aBls4d3uFMfgduk0QbSS4SyVodS1w6ACagFNT+8svlBtfK6Iyd44N9iBr5
idJYA6gG9dPmh8NzfJgi8eF9f553pnepYwIDy0T2Et9hQYFOhO+dCtthJXlBOoOo
WDrUM4lMBJ5Xb4ENv4T3O/SFnplTk49q4lUxYb9nhADYkjCDkEqkqGNZmlDPXlod
/NfkqbGkA3fwLpYIVxP4ARzbIypiHM0jsgzk0oHjD/LIcl/V8/v8YZvielbHfl/g
YqF79nx6KdepcrAJDQniRCpQ0ckYa80OE2vesYOd3KADt2hlwwCkHekkScZhwigx
vnTpjrQphxVUfYX9JM4em3WMiRomG3jyMxjKW042rLWLETN5nvlxdb6FXaKKDSwD
izoaKarYJvj79cci1YCSTFSHENARc2v2bkjSOxuDNzcAP2+8U5zTJh4GbQuFIWSy
QTCf3LitFbxdkssZ1ZFuF6alTbt1TSl/R+vVgFXgGDSNdSjFykKKyHHVwCQHbwuP
Et0mJIk+neLY2sZda7/xU/BxzADRBc7IjwJOGwm8OjjnBQif4pa6eoq2NfGXmpRi
P2WPDWG7R/zoZcOlxhwow86yqv7wXLHvTJRYglJIH5MmIafmd26L5z7g+5ILc5mW
NHHI8gtuRk+D84hCAprYFYaQ7D9tX95QzCGE3OFCgTov8YglMvhiOQUWzVSgI0EE
hkI5lPT0IOEs2dax5KIFLEcIifQuhmCgQfTvEVeUSBtlz5rbHRrWBvNJWeBt/1hV
+vU9P0XCNAWJk9fCTs8+5RfpdAAIKZ+JhQzeijVwzRSR3vD9+tGz+3sLuja5oyQE
b8X029cnRjt/FFAHaFyhy7+pVqI68NfjfHYBc04JijxZUSunNzsgInHRuaYddaMu
ZFgZIsKT1aXQ/+kNOlVJzCdobIC1IXJ7s0R+OJzwWoc0xDnNFfA11LgQ2if59LSR
fA8vEED4WgyFt9CqKt68iBhisiPhXo5HRrOe+DR38uS5bPAy4eSubIUlY20ZuKCn
2wHuejAlv6Gj27EomwJC2TbSf53nO5aQxNzBsvcFyEcDDdXa7ooC00Wwc7FSR6P9
SdLZ16N6qEK/FUmzAjc5jryokog8tk/aHl2kn5UZWeBWDJASulIJZJRNB5WRMEqD
dR2UH7weBbvpLaTJyRlFXwtZXDk7MXrqs7B22CYtrf2Vp2iUXWHvnd8hwLbQsBZp
XBztpRHpsI/vDY4550WUsSiAIsl9JJ3LC8ZGoo7G/9arxSw+tmGQ6SLK/4VKCh1z
Fx2cQN9AaAivGVMenIBpBYkUCsj3kxGymeFiQnekw77cxIZubbdOvjzx0T2L6e1/
T7HwG7byN8iqdqdytHG+AJANFL6aT1IGqX8fiXAHxEj4MUiJWzMzFaRrv19Dn2Gf
BCeaBaXTQDePqXvxY42UVHgK+F7uBSAIlvlFsUL7FjCDCw8vFfSfV8+m+0qmum9c
0sMZPT/TmzsARH9pKqEIpGeLcMY/yDILHxU83KA+AiO7A7K10O9ZpTmw3pv4Zk3F
meE0IsE7HtzTHtC07oKB4f8J3glUOApst5uS9BaWd1CLUmbWRvgElJGC2SSV5WUZ
iKkoTk95Pl3Iq2nBsMfRJu8DdHCnK3aNOAKYhhAiiIOT3RBHKS83ELR582DVkTOn
5KJZZJP8Y3FKEGK0uMra/FQv5fRoqv1TweL2P0whljzNGdV0xy/PeBFadGMsHvXS
/qumZOQoMmWf0agIAZGWKx1Fh8Ok8q+ENZO7ke1jaBmyJzBBtuFnPgGYWXEbUiS3
+fGMk28Tf65uJansLgHuNhiISDV7WHHmSLEq0V3Aii5Xy2c7B1FLUg64JV2Qb76X
7jdWBS81fgM3ZL0GTSRpzi6Xsw3dgEJw+SCKUvWty+qbtrK3hMO1LO349wIKP9ge
26M25733WSSIODL/gkFMo8OAZGB1OB01TGBLRvHgwq4VqhpNp+VF04VMTr2TWnHz
PDrYkMKCQ7LTYNIFnavTv97DTHLy0NirbKf63RrwTpSjHbQ+NLZm4reXpol0T/P9
R/Tys1A4AZxycOqOglVYk9vtan9eQe0ZCBBjzf/E5tkbgC+WtQ2tZLN9JJdm4V3e
kzIw3sM7gmwOJ5TXiiVYTUcTlhiXtjr/YSeblxgWN7XNXf85NXLHEK1WKhOtTfWY
IwbGvzqwHU5KXojn2C9/TAeICmpsIrTMHhUfMZYWKBVBiNwHyyPw2mqqSikYfHAK
zQWty+ePdzufHReUx0MECIMMxL9NhKck/1//icxXzj2Ge7UWfLXKNcTs93wjKDBF
3HSb2O/7ijqToRY8BVh+pFDUqEOhjlV/3BtJLIj8oSnDHkItL/ZhptkeZpJ110bH
Wp+I55i+21Kjtqe3YCTLzsNDwlE2sJ+I2Mi/Z5JqrzRAQeBe8gPAgRA/58ZW8ANl
AEHiutzBjg2eE3Ls6OFzRFhy1ofvejnBMv9qeA/kZH5apnJH0EQT++TQEnTfjnbA
ao+DFfE4d5AEBosc8HnwFLFPGD/66AJIZ0+e3fd8s5PAihXH2tubKcyy669IcW77
hvd900AClkMXFNsk7elbt2+eTSFYg+0FNiAUK2/+NDQI3XCfHC1lLFvOUy2Kd/gw
odq7ydp54HwfzV2hlAExjE5KRVLz/E/A5VbHowFSi2PY4EGurRC0qm57mo1D/AEB
WHZkes1rNTbCy8EkFZTs4gy2dhCq6JTGHK3kwtB8qUMIq4jNt8QzLQgtZjZqqEYI
Kvh7Mvn7Kemyzvs6NQ4Zq5zsv9Mw9nfEjYyg1O/TWx5PTZJeAkQ6YgbYpk2sP1bA
v0CPG/wm/WJz774bVf0II5eewNEEZayUcJE5tppw0pAFT/+5xMiFJacZDqFm7CG0
rc+K33gz5EeX/sDlh6W3iY08he5AY3wc2h5MMX9LGKtDGROP+Kn8zAq6Ak9tQvqg
xTZwRuaqlkfqX8O5ARf4cYPdT+datA8vBjYgRl8piEaXotKJWSN0CENQ4hf7fgqb
0KEReHucKs3ZrfYO91fA90JfqNys29XgKyVDivD02cE3v6cwAFhgXYLSWtQF04MP
SOJBvitw4O3bCfVG7tk11jN2BHKxd1C2ocL8rSU9v+c8t24t/ZCuY9j+gupTnO6e
u+09eKdZPB5riTw9JWGSiIUI+Fp727B+G6wSrL5CsdCtUw7zH0TjU1bxyWPfEN8D
r1g82YjylrnAWN1VP8hoOld+Mjk8WZuTqHWX1vMM4+/Fydo1ao4Tb+5N8lgclVQ9
ym2Ix1yrpxkUh8yMSNVJeIMeW9+/JKa27+6lsCww/hoaG6JlKsCWy11X/YyibNMv
ZppSqYDpGgWuIyYBGq5MvZpjBl6gWqst57G09a5B+ZYy21ArRAVIJOMp39nRv/ZX
rhsrkA3rOpu5HS9fIVAvCOnIdwh91VWwepx5RoV3bcuWAzUyFpvSUs+pNMdRJiMV
VUn4i5mvVG2LJIM0zTk7rV3iF/zj6vi6ci2AdJsk7kR7PoGET5oNCt6h5Nt6lvbn
31+NLGby1goFCEAGE/4muuvTkbjQg8dUGKvKVoqgFkJ6x+rwNdZCCKisNsiAkYyw
dkshmryhYup4ACvK3P+rM6+zQbXKqsIbLzJC06oyP4TTzxFh3Z/qu7V1X4OP/YCG
rcY9+PGNZPieiCne5LY4J2O/a15oD1uZRUb/uypSSscqDOFyXP3lU8NL1mw/DMgk
A+F0PAgq7kRu6DlZfZOXu7dlhtIelJhavUNgDRIPyhpqCIyGACvp1d9CbiFaccA8
ehFCpXj29AqU2lMWrYo+eWpPNMvGLeUnGwTHRynchZjkkmJaPkMnmK1qqIPIH5Cv
RU9A6BifrxZlZ0fDFcwk+4cboqCPatVods1/LuyRjr6OoR0iLpKe9gwmiO5Tap45
QgfwX1YiRFZliA+60uDHbqhXZWIuCj6l/yYM9mOC71GcQVij6Y9nZ5IhsgIJdRmE
SlqxOcRDFR/C9W0PkIe8xPYZ8Oj9oUPmqNRnoP8VUUTjTFX6jg7ouHfwHTaAiw8w
kQ+cu4M5Rl19NCBzO5wumqSLViF/qvkrAOe9qXLIEEgfLRMCSg7uK9c+FQJO6q+u
Ea/OdE8HanN+GwzBgNgtAwPWmBdbZDsBTfMvTmImJITxrcGbPOBPj079ftvhSqxf
auH2X0i2sxZJ5Yuw4yhjQJW6CR177v0LEpFhR7K7l+o5riAVWqzi8y8/pLRn9eOu
7HVIjp4L/4xZ7U7vTOdWOBNu2ghGpcx+qYy8PvquBVYdq+BywLMwu+qsOaZJ+75m
A6N7OehDfMDjN+VzDo6zs/Ktnjs9kVkiXCWscGLsuU73RJgVrUh7nnYNi+D8vvKL
y06kZHP7WRwUOSCm75P3LXsAlETV6MzW8rNfW+iclBrpebtx5+o8A4AvPP+nYTyH
NJTBd425UiaNA2/5SeBoiiAxkMWLRzqadKGLCyH7RwgHU3jegxdELQo3sCZlt1pr
lkKWEjq+l+P3wTCuB+lTyt7oSfBGSTW39IG/rj+VrFukrZEH6cJEh21qVZqqHo/j
HURTKB9xQWln7fx4nA+TzdXnQ/lfZSzqYnRUH9pLP99iFN8wPxX8y1s5NkA4EZOP
Fdm+L/iB1Rj26JNDgo/SLL3HXl1O5rcOKC9Qg/E8VWyvAwuhyOmND2LwJWNXo8hQ
bknA4gspbi5ZYiSIQLOveqBeoPuqEPpmzvfhaOXN9wadXsBAduIA2145ZDpXbW4P
FHVrmTfPzEnJzhSt3spvFrHZcSPmbVCrEw39xSoPlAh8uWo0PNgZdjasGCcyT8mH
v3SraqZccsCIlcy1EgFqoD7hhvRZSLNq90o3P5KLNUzagyrZU1zPHnCvf/SFTdSr
OMWCVirqBqY9ngvCMV7Vt7ZmI6WEGOuXGttnhxaZOnCyzks7U1Lw25XYTmtvj9d1
lC48i9ypbd+1m7X33k3wHDwIQg6YT5JOgolYNOXTQ0SGmTWVLdHUs40N70K7Mlv4
NrvPGlitCQLDnNeGU0mfd5zwf+Y8/xQnRVQpB8+y/rdlU9e0uulJxzKiL5/HFvU4
FzB+0+uAuoaedredYi5Zc25xZeHDjXQfqP7iuaQ1lT7CJQq4mGvIM/RFmJLy3/Nv
KNd4D9xpL0cGioJmLUdvu85gDzbXdY/I69vZQcl9YejzNIAXdTxo98GczaNyvo7m
AGx3NJQYKG1lniVGhbI9KYdzw4b89jb98Tn/vaS/kTnN5blQGyNUq9Jrb/S37AEY
Lc6OeNLslw/bd2/gvVN4O6GMRrrDxtRaYJG2h7t6pBDnYGYUwlc+YwSpKjI74T7A
PBDoV/OVAaXEgPN0vF5gfadX2iHYUUW+HL+saxzP13lOJIRglDzd8hNIJ8xg7hWd
ky1xwiasEpyDBBq27BN6K2KywezApedXJ0JBjt8L5DfXqcGkTY2eMushXI7HgjFe
Mnw5Yhfs1SQeVdHZ7fCffmIVcbERZS6U4hueiFxVKkxx2YMlkhH3ujjySt5SCftG
k7i/5d3+oKoeOsyVq0gjOwg06qKduVFOlwErf3yg5ymjQ4CgWVNjbe8fKXxFScFX
z24aWGdtaGLobKt5xv1vr0WODSY5a8+sSJw6+tbTs3I+vFejdfHbp6lD5nKSLyWr
rTN4DvT78xIK6DGaJHBJaegRUbwmRinncPc03jc6xLuHH0+r8/YgWYvq/BQSM0Md
Fy+jE10AQrXd/kMq0McH1nc8lKX+vB9bU+ivW403Fj3l0H3nFoqM9OmvjDijrVN7
uWbN+b//1M1J0zQAyh8EgtD6eeszmmyLeOk1ExowzTJGWO5VAnlNQJeNZF5JOp7N
0ufNtwTGDyxQcWMXC+g1brjCIOpS3L2NlrNjKBoAxcOyFaN5xoya9mxT7uKx89UF
cGijRYY1uHKIDTQqBlcCQBJZ6IxDHWGJn69wh2q7yWIkg3DMSQUHDth7kqZAOjoi
a4zUlLP8vKMageqCqdLxzKJAeoRESXsu+UK1WcWALbQzYCPzHbF5QAs6amg7K3Kj
Ej6xrBAA51GhT5+DO7COeQZ6ggXILU+BxadBBoo4qbxFRRRpWDQKqg0gdfTdzt1D
aQh4bBwl6JHnf4spPeIELjkIgRBERBA3/B60HR+VnF5y4qfTyXAGarxAatecnCxf
D5s9yI5MkNcVPFp+oYEyUJGBEymRB2R9Njpic5m287on+zdNVyuKsZHSFwSFDme8
4CGofcoMXjReYPGihIUk82pJpM2U/S+q3LGMdXOp34m/g5XOKRkhZKF6eRpCmJs3
WJqmmGUBuLACrr4ishLdeXXw705iXCr0sbOYjYBuq659bXqQih3c+ak1kY7iflu2
cLnQ9xlrNQwLWXrXj9QaYs47UDApHsugAZ8ZplIwbP4yt7PtQ9wVdwG+2piHqkvy
BG2D8kw7pqOC8D51aPamaOKWUwTcaUD/UaReaubQ+OT49VnDlXSCEBXeO3OcRVtK
L1HXmLBWJzxcaSpgcU34V9/TDyLzzxWJBVVMZmBDKtr5jktTVv2l06dTDIyAJDGW
hqTM02YE5vsGJVrkf/jQk+uTODZu7wiDw7gj+Y1PAwtcGheBT1Ru80wuF12noCxV
D3Tv+lmSQKXtG3/P2Xi5XPoizup9YW8MGv/u7U77qJ+UW5Tr+Mg2g3bgqodr4a3a
3QD+urfpbzRPwrWIBl5Eq5tDTwki3YY0FpmIw+FinK0t4DXgU3/VcWOlN1YZbQai
Ig9hTGztpISGLGmWG9EhHRdgkIcGLXRpE36wXsQXYzcUGHiSHdMLUigV67D8DHSp
tEukU80NwAfFUecOmMZYCONvco41kbz2h3hfT8SNHFfOUk9l2HDWfChJCTtaYp+O
UdKQU5X+1EhSICwY0qCQR9z7CntLMkMzFvk+lpzAPVgRaFLFn2sFqITjm50f6w4n
04O6gSmdISBXPyk6c2MbMTjUzZdK2U3sTHuJK29coUZkQS6LaNJyCtYWnHNnTF6/
zf6EmFURMffd2XCSUIhJN+/FLWzxKDyt+6IsLc935Hm1Hir+EI2vL2XAQ8vIt4lU
kRjvTtF0VpfcOSKEHnEhWZEqY2fX58CGwZJ8qR+qw1DfCFr6VWEUga5t/iVsEqyB
TjtAl3A8rtCE2Hy5qL++XZcl+iKpguoFvOsAz+FyW/nVPpYlWxfqb38HwYqFJGET
B4yGY9QY2gpB1Ni9WbOGtefBVVetmxxXz63ITIYE5/JYJqjkNfxgd/cwpj4K4+kn
v0mpUmh+fFR8CTF7HxQF3Gn7Wtvd/p5DN5IkqBoIYhAoqIjC8o76vjWLS6DyJgPg
ts9MuezRw3pW+WwJgM60UsumxZo+8OISVucO2WhkD27Gx3fzkUNXb2xI6mtlMCbK
CFUnwTQ3wdfxFwdZh+MI5GbeZ3on/HK3RNdYs3gety9sD1Ai30tPabX/PRu3FUv6
3JdjM5YpadGear5j0IxDiH77SCyMYl/xFNIHlNTJ488IiKzPTiGfMjgKrfDwfS6n
WqCandPSYAEurdQf4S5UVD+d9afyuGUvBcGN3DMO8dS3gB1kSBSuAxYC9BueSWyz
/g4LMKIxfgTflbxZHA11oKG/5BFNEuzRMg3MmwKZzF9ycmD8FNd+RRyDm6YQ8laj
+Xqy2Z2rwYyPzVPqIy8W5JeKX/nxvJtCtGg598Ow+t7u5fWWzXd5lyLwr9YNadum
Iyuej6s9wzOUNxp/kECQVSu4FYJuO4t5ecNQR2eD1TrHv+sV1SljCzYOruVMyfRF
MnQZ9TrCfAjfCDqRgbAGm819RGpgmz9BJahhpgxElIqef3fhAfNEa/fPgx97ObXz
Go55uw5g1LwjNbdfkARpVpIk1WxNacseOtOGhwELEepmOExMssQTUiGqFy9zZuNj
/dq482SVRg0/R65wqv+KHOWYSUlMBX2OWdzOQ8i5GMo+PD4MGLLB5ake6NT6IWNQ
ajZg+RxO89Oz+caJJzcz8FtjoQb22HqIW2pGbofuc67jYoh+qhAypBLnVr65yEgw
KtbVuY7bQHaf/T5Oa8sK2EgZpWNF5pCLBbL8oFH/8QcNYUALMB3lNE1dZ42Y5Yzs
WdNf3xLKOdHefuji0+lIbH4r3SNDSRS3voFSXDHD+Is7/xgpIBNDkw1vcK0LE2El
EuwuzfndrRjQaAwpv9NgnCvhzw44xZDH+72gSuOck4DfE+BrVglcteNalA7CynAq
A/9YzLog2N/RLGeILqZREbtNd0kGWuXMmj8luVKqrvaEwg0wCYM5W64l67UEe2dt
1NSTOcihyncHDG4KIcJwkDKOaHYrTwHO01UovULnWn6eZdQ9fLKiQHDF+Sjjx0S0
l6kHBS+fGUpnnlbWYkCGLpBrRKNVSAv4Hpvf2v5csrETzhZ9p4XLICkE1zQddRwB
+RNvRwKqPVxxI4c6yDyFcPTkB/cMbkisIKvK41WDmgar3CztnRtzGVwmaz709Xt7
UP0HgMQyLmhGMbioogNHVfBQKrzg0RVd4FeHyugsCMJUDT4Q6AhznpXX2LHBSmMB
V3p6dYU5fIS0RQLFQGIYba7HLmMlwPG6uNyXX9uR3Li6ZDZI/HaC0ZPk6aoNMbeP
++hdvddKX1bLvnOCVcUcKvljYHLDR9YZca2/ajHiVJkxZ+z6oQku3+Iz6BywMt/n
GegmWUhDgaiPwQ6AM9iOVXgrNIbk+FyHeBRhqTDj1AYwCMsqbKETnCVK07LtZX00
+e3t6/dyL20OP8NFVR0gNifbap2l5NozmzPKAwvv+Il0LWZ978lqohokzaVvP3Cn
FxS60qNR0E9E27AIHfN+LjLmwCs8eUwOI2+8CSqnLNnzQA+IcatEi4vX/hnTwB4N
fwco9VEz2IsDjz1g2MoOrEf4wF+YLKJuUNw02h05SrcKG8Xn0p6MFZLBgSnbVT8z
Ab3l/DurIn6BTLY0LhWuzYVmF7TDUkh7IeUEM2qGEFY/P6Qe54jH7fDYeWUgzLKP
b/1RmZ245Ant3qXqhpDorgmqDq/B2Mv49myP3RhFgeq+ccxQTw2cXdIN4iLyrcBN
c4gTH3k4rwEU/+b28rJ6fgToo/B1hyhM4u+sSl2dlB2OBAFDUcBQXtoiH+rIYrXO
bHQhyv9dwQkyp89RXPvJK5MBs8xDg7NvGTs5WDeFCPxJ64sWognJwsCs/O7HBSzW
Ro6fhF5yEDEOUegW/e6v8jILakWQcNjfzJfV0F0CcpsLQNLdzYjcA0YwdYmYFTVz
MRmrD+gMPw/qtvHfF7k3LyDDtI3yncbC3EKhp6QT/J+ER4IZaC9nSpTp9HayWQwv
Vbh+1aLNuElxWCAyMDdCSJQeR4k9nrCnBh2Wrr1Z34NveCyfyA/WGihPKPo3f5YN
xaGm5pine2x3VJNxZMC96xvJrVYM5KAffkVA9Ofg4Y2KyreUBMhpUX81YqAfygUk
WQS/+AMj7g2Ff/XXuGBOTixrVsbSOSqUP1Ftqut1sqRT087UbRlnpnm2T5qqFkzJ
Cbh3vewwVpB8aNVWKvq/nhE0yHZyfNdCKmjMRmcEsnfAPToFIxaqMOgr5zlg+9ST
AoMp+QFlU0EEbjGc9/gUV/d6NQzMPlehJ48Jclz5D3XhW/AcULXStbNq3lNtSJPL
bFzTodLkqgsxGM4OvltdIJ1+2DsXNdAhEc9SW4oyWmKp/5N5NZ8zwdETsENFRhU+
Po1MRW/3MYytjKsCpGJUdS30BV+9wJrTb1VS40QaVsgsgAgxl7ZfMgencNdPk3RR
wz3nBuxu1fYg5foSE53/ZupXr9EsccG5kAUgCSrkBp+RkOdWm/8Kb0pvwiU2mPwK
6AbVQFb7HjrhW9thBXnXxrrCQFJXXi1NOJxOFtBFGseBi7vMCWvxwkCfs+cbdJrG
8JffrbdrVsmA0NfWXAknMBJdPBy6TLhI06MjBiyTLhUgPP8zymE8Mc+AbNzWF6q0
jEb5goqFNuBuBX7O6XFSy7z6p+R/Ey/IBxroaUzSfmoknVpEZBTBryBvdMc9zA/E
+lI8x8TSFcXuuWS6SCXoJLT/0d6eiv6UUfIKaPWaGBMRCvcqH/7AFT61QcK0VcZG
GNsxobu8RosiSdW5wpN9xZM8nPmQ/jhFMAmK3nkd/PtlPS+JYGy8Gs5mjk0uhKOW
2cLs06CFDiMj0hW0tEdltrvZE2Pe/2bgtOTseLeNo8cJOkV/gBNAm1PPLR2osOHO
ScbMln68oamQeVJqpBzL6Ndiyo7BgtoZRSNKyT9loGa8DDGilU3j4hqBey7PTP7y
QQbqke0ceifrnDJ7bEfQ+dFMHJ25b6mFBQWS7ODDe8B0730LajvZFSFE1qIZvOJ9
PT9nFOe8s0aTdxvyA6EwRcC6p8NVU5p3geH/h1XXZ1h266EiU4FNqmnf90w4K4B/
EvoCALzwwfIuDc4NQ7u8OtRmg6PsrWVaYmBicwiOjJWnqXASpBHh2+asRE5zK8PF
5rth0gQr2lxotOyOYIgw8IJTpD7VA5qEt+qRH80JafBjBLCa6Z+DKxbClWKRfc5T
93r3c3eYCr8vWA7oKdL+xLhx/J94q8QTs4zHV+1oG65Izk4HWB4EA/yeZf2JDYlx
vq2CIbpV+lOQTbGO8aIsnlyWDSL4QePAXAf4dJlfqKb0uC/XAkSEwf1A8d9vYLX9
oyV+bf/iV7wp3HCwDt5sH3pt4r6LDtwBqFI72Pp448WTOPBZZSKwb9oGNc3WoezL
foG0ks784Ltxcm3vh9TPnz7M93z4FzWmqbZr2H2NP5Y9Hya7vTdSd/5OxS7Fyt6N
XgCjfhPdQTyyv6Lj8Tm7HWkmMJDMA88lgiVKHN+PSLktDFTo9xQYWNpzKmF9Ilsm
PBbdYfR5bdcc5vgHUZPARpG80RpOLgrTi5rH3/5jAQty0J6pxvnqaRhJUseapMhc
z51xhv4Lonb5RPNHu2NrINDJV8wfU36m5Gt3a9MgF3+QScmZyMrfiAjk25jmnnDe
mNb1FPHMN+0awM70Q3E1tJj64aXwRFBzvj7W2IsjDDDqDrdSQ1f47bBe+PG+QVmM
it9hC9obHomLcnfuuWMLfr6Zwoaq4Ex4HW2RZVxaVB2TBlmVPkd4cH74q1puRsrP
XX9Y6PfTdIClnptKDgfk+SYAbF5vPHZ3cn/COkTuXK3EO/HwWsV6Ox+7goQyIJRK
ClrgFSASxyTSY2Sz35cmwfFd9jM2W5m6d+2DCuk0xWZSauvdnZ+CL8CTLE3pBPXA
kqSH/j53zNRw38Juxhbplt4pkLvNThTs6IIqsu2VCkQ/e5i67yu61wZJr8gSO8ut
/3ERsI0cyNrKra4J5kCBlzsNuikvGU49ob+AXZVhnzX18jqVOinW4gnB+5Mm8DfT
3cG5NYCU4ui5LGXhFti69s4Pg4CTCpwOa8lfM+bkjBYe1TsrGQGeMFa8s0X6/kQa
LKNeaHZbyRh7uhsMFqIrvwyd4nNcyOZdSDvXc4KoYD0a8kGx0uNeOZOSSlGSOMsa
3CSmnzoWELAz3VkmWCwoOQhVZgQsFlA9CBHbRUgkwx8rHwyq9lp4QNk27pJjd9VO
AUGTJRnsOIgJc+Pb0+JvtKl/Ex/y0FVmon2RrWxV4XyUqVH+/yz85qeLxYIVnq+K
sPuny60S88LWguFyc8Tb6+Hy4Z8zp33Euay/dN1yLEbhC5A9LoFEyR4l150Bgd/T
JpVSCO15BQqJzgRPDK7/HSUvN8hBUuwLgaeCKWZIWLjygtcZ2d7xQ8U2FGXDHVhe
HLbqjZ0Q1ThmoA8FzsxsakDSOWYkwW6J6MBlsSx7NA1ZlBzL0qs24PGPHIYTc9v7
FZ687RQhXdgWTazg3B7ZCBAsx+obLmPq5HIVXPD4Ypns4fli27eErlY29E8fhrq9
v8u7wbMQqm1ha2+NDva4xX7sg0OQENBaF8n7zmHk/b8wZaQdGEvy/4Z+QM1KbAur
iG+qzH++Sh5NWpOiQTMy8WP8zVIUzGx32UDUYxdIN1roNIdfDRa+tKLpZOxoNAuH
Ggl+U/3wW3F3I+ZJ1L1ispowjBmr53J/x5aPpN2WgrUat64UY3gdpNF2B7yxNlna
7HdggvnQcqN7xEUBfw38Nj1T5kMe7feAOIbCVtwqKRa8YIhnzxn15IyaQuqg7YPv
WJKpD9okXa/xJ1saZOo+dYJrsumnhG34yuFAtjM8ZdxQmhH1iDPXWZv9K4urnWcy
ehcLSTxzLClrQS4PYj4GYN3PR1wa0FALp4Kyio52epTqT/wYOKhEArMkS9MUMPS3
nBk0PIX2PYu887quxIvZcaef0oK1pS6Xd7c9USeA8iN75jYTfccJzdgEWfxB2HtO
1r+3pB8XosmGMvj7ymXkHKurjysSjwJPdwuXKx+Jq1xqm8L54aL3pBrlLbe8MyTU
B3ttkwhN7Zfm2J0g+z01gySCZ19agrS3eswZMsAv7HSLMX4M+F/6pW0yHNGYwjNK
mt9SO5x7qp93Q8dOQQ+7KfReKKUpv2n0nSaEQBquhxvlok0yTggAnuxh/ZJH1IJt
Lp/8eu/b0F8UY2cFBnuuiqicz4DHS8GUNp1X9PI7k3F7BOMBsIjhORFzg0uDAjc/
JKpZoxN6QgLCg20wODnQI/XHti5ru2ZPywZr2mpUzZp/w50bYEhDSNCZYYh/ld3k
tTedAEZ4c9pJNCgFeYMbWTUbFiC+MZILuBFifnRuejg9qb7aiJ/s+THQmVr6i3Ka
GaeS9bjJ9slA2/1uxI3ZN4m4MOMSkgk6OD+2ZADkyluEj4dCFpM/mju7Zka9vzlQ
hP9StPhwsxdpJBx5ir2PgWYlHkNBh7VuHYo9yxvyiOs7myf063JZZeDuFYtmXjuv
7kcDcN4Lzv1Cv1tVs3E8jO1bBZ1yP3j3pB19pr7qD0sjZACZijR9+1Zo0BPAXctv
CTl0rPv69IHvqQ+ZsNkL+zkWv3RYzkuB9alTyds9Ye/M7aBxuJlamKlETTpsuTmG
+soeoEMqAuDbabNYEL1JpqP22irn56YIEJzbwkNRahbBQLYXrDtgtVuZHE/4p/ED
0Ws63L1tDniPUVn0abtlQGFbKl1XedV9eaU1nDyKkVm++QngpMaj0amhHyGaORIP
E8VKerITc8VTyHrBG9nqQ/S2IH4RFYJ+uBVhH1S7/QdfI4PpRWlBXIh+VLq+k5TI
AjFGa/8h0xBnSjg5/Eq2YZkCzlwo476gkrJxGuTVBqx33p2Dq/BBaXJmX4qnMDN4
tHHR3HcuRG+5HSd7u165KYvIzKUcy4IQOlKQ97Bwz7RpwoMAEJfgn3jFWMrt+sj8
PlgxdsDNulJ7TUQdgMvCHXTBUk0RQbatHFTP6VGOW01yU1xI8aQQbD74ft3Z1UKn
Hvf6D+pSiznMmlMVvBI1U8qXTE5P3OzlAhP3Blujitd+wIucY9Bz0FoVZe7NQhAA
wVCgV1J+cFu/Grx2OdRengDJLzeod13Yxp1p8VvVIHhuXnpX+wJ3xhUyjVBnntil
q49t+wXhG4YKAkvyLSBxH8NqUIVNySwlF4YDKdLTfUz9HvbypkWAp3bBc1fx7D8M
nliOmrGlOBvbJVSgr33bO0JXytTJGdCym1whB9aCXi0KCNluu5kLkMvBULG5GVy8
QJPWI/T0JeOAMP/DLQiC01Wljp96q6OvVDN0rneEPbCA7aQd5cRsVasXmCDCVZ13
nYiWH2QprTpY/DgcLOKyJk6cwnssPOBTK82/jA5/baz75AfV5RJmXx9t9IUD0ik7
3QAxUhmfmJ2B9QOtwr5j6Ffpr9OpsfdUyD+H1to7syakrnEnMx8WeJbvoKQpBAO6
+6dEGmI61l9icUA5rQYTJgoSfgRWRdE4T34Rsjf6WAvgKrw4viTC3WnhdSLa7NQn
3+4UWqn7+sQdIyO/Quvbjne4s4jIg2gINg9H7MuTaYNyTliDwiYVFuJs87nMgE0n
3Z272U70IfTpwWxANgcXpFiZVXgrHT5oLrDdnNwFFm14xOjWoj5XAUWuGv0AB/ux
OMMGKXLXZOQMX/ZytVHw7+bH7NrpWOJYr431RBH9Y4VHDJ9FjbzMIc4kQQAIn4/H
a50t715TCSsB58u6Q6SNcsHsSMtYOuR3SMDJoCWa0X636HxaXV8IfOqK3VOx3Ifd
hLw1WWbAt7OiHSZPrSRFlzjgzohYGI1hEIcEQ9S98cbeKll5wNl111VhZlmgYcvU
luswFCZCkullNfPocJKLyckLAhL42oMgc1DHmOttLytqHDAyd2czNeA/+8RIydz0
+htwIyl9Ml8lhksa1YbsX4vYy1gEg5LcY04GUXJXmITETwjE0A6van5E1lwPap++
UoenyG2VPTrc4NTr4Kfcjzau7yGAyvqGMY1moRMbJRLoqAjgcaNgC0qxeYau2Wjd
ypSrzjCfDy0rTHvdMtcPKsXnMGscozdqWXPrW01PGIt5sUIddfzLF8SzgfcnDGxi
AbiVSLi2EKgRMRfnomVGcCKrAXGGnL/Glkk6eZgE9RQuaZXy/QHZsFfUZJGeG0iA
vl1MQVIJMoA3ob/7qSyPvfiksyBVLOOclX3h4L6SOE6OBlZ/1sWCuSnHew+SC9uc
YVg+3YimX/rdrm/s8IVoBkD8P55WBxTLpSPHB7peFIBXdjXXvnqCo3/p37fMuiQg
wN2l/jY1rBRuspNnipfxjLlZdVz1auFlwCaPPUDuj+UmNBSl6+c3gDgQQ321mFB2
2JthXTwOLb9XMWG55zEiv2sT/iPeiJeTSrb9SFHCXN3dNLefyYx/v+Nr3VCm67jv
cyuRs8hfu3WLMwPEuw6Kdy3bNmH6lS4RbEGe5JXlbX3M883eKJOCag1LmT5Sg6gd
dumGU2VAih9EMCDsvlrNSlyLHthus1IwhHROW0qmRscyr5f8uxjyIdr4L0crtoi6
ToGEgtKm+A001czGHGfJtdfqOHbnikkpQQNfUsvXdClbTrogO14faFKfYdR2/h3o
2qde8H0woNC77Xg3t3Rqc9gAH+1tObEM6+EByiDqxzQ54cwDWCqDqvTRHTvQuERL
tmJajgbybzGJlD7HgOJpVaZXLjCMOOoNCKGitzNwCivspM2hPytzwTcD/uZQlC3T
KpMXp0tlVZ1sjWHcsFSJYVPXabOogmYydNooILQYBtITwubFk1pD7FSLyyjFRoS/
+zfmRDK8xd29mRif1OeCO2lycAkhpjNU4ax15DErIN2ugZuvv5JR73HsfBNsADAl
pQX/N2KWuD8ALRvbkB+Viy3rrFQ+IS00xnos9AZkgyv2fp+ElnYwXdurDvj7Cizg
rUJPdUQJ2c7uJLd3Br1wUvZL0jHpsniDiX5EANcI+6TyoFK4A21PrGIFUmY+ydSk
HV4GiFOsRwy+Qve6w5VTzVkIwnFjJmVQ75RxymdvtArIdvi6Ub0RASfGSpAGKNca
efVYTp78d4swEQVjK9503VMHguwylr3FD5CF0GTpuaG6PT4tlMTq+TkDOwDIKo5V
NEVnMNheG4jyC6jYD8vq/hd5MVlFHxJfIU3GXJK7r3el4Ldm451Yrrq1SQCWK1FS
4/va73UmIGHO7C5fj5WtdEMi7AnQW4MUg8lYjsIX22nCQEs2ccDwHmMMsshZzka5
NLJvG3EL+jm/yfZALG/qP+mFQWAGqaHmAkKgM0RxFombxOugOTiQQNU/S4JtKZE0
XQ1sZcVcRd++G5RZWzUMNtyVdBGu/Ikl95JxgQwYVVgwJiwy3qDRQqazuiUiqMgG
ZkQNcbC1LrDqUPDNHS1bknZL2NOk39HSTKpZrG0htwzA8nzMw2GSJ6Ub34Kkg7Oz
MNTDQ5Sv4qLgwUD1cN93jnfJvfuCAINslUl01B9KckUaEE1jYwyfAJAsTBMaZ/J+
XWaCxo46AWce6fThMRUwH/1OehWmgtIYLcYKSHz1ps0ccgqAzGSGjmT06Erbn22M
OwHvB8esybUDdfxnSWjkqboTT2WSslXgGSPibGoeGIys7OVZgXlq+xkt9JTjq+RU
GZ0TdtEI1y0/qZ2OIyUUm1Pa8K+u6UIqThNdFCE9d2SNUoV6UZhg3NsJjpxYc9Ii
kC5wMgvhJ3Ds06pf2x2NZFUtXPGdDFgMkIM+i6Sql4zihxvvr0rqw7Us9Ar4Icfj
A/qeDrCH6iHEXdsyjdkQnTh82YIeFaSMqye8Q5qwD584s4nBE1+UgkeUNE3S1mMe
GLBznRhzvo9oAN8myF/ImBldP899niOWt4iA9Uuj/4+Z+ZN/KlJ+9PGACKWbVxQs
P+F5u0zhI3iJeVel0KUZByr/4DiC2YV9Jz8PfOUn6+pDlme4/RYonCujRo+umRcB
xkqCSeIIoOfZE6jowKFprC5/fxb3dRtMCmx2UL8VQW8ODQmXRPy5NVnOofYWljEQ
qNRHNotuSlRvu++/07tMDz1c7gPFgA6gofY9iZoL42C5CvqxRXec7ddy9IDglfTA
lTkxmoTuE/tmKYYCnR541fkuxfpZWZ4bLbaePHnerVAyNxrmA3F3IWKIKpej1foz
MYP/EtW37xSZgdIlIvPY1NLSVZnJbAZgNM5LQ9/tppPAqIRL/LurofGfJW53tfVS
9Db+1WesM2S1cSUKK76QsugQ8B9G/8Q5Nkv+was39hx9nDHXXSlMyXjZwqPN6Zxa
4m2sezo5zdkXyntc3JzI3ZUsXkQMhVXWPZ4Rt6nXbDcfo3vobPHXdxAUUdWtgbCd
CpGNjo/k5NqSSs6FP+PMNJQuHjuRO/B/kYAupKSjpwPLvzfIpXzQ55pgO4BcnKil
qIgIFc0UbQ0fWcRxDKL0Se/L22GvChWhOXZFUudGnhoyGvErGr6ssYUHzRNsFzte
9mtoBBg9HBwO6B3T4Ccki0ki01HeDVy/h7KbJzfhF7GrHIRKJ03/HGhIjZ9ouBfX
TIx3D2m3GkKT601C3JKlesVZlRVqfmYJ7VFBX9X/AzcmMhVlFIqYIQ2E03AoroxQ
hMmliawipTJvHcpdcrLaAE+aYM/idYkpXxk5fSb3T4HiaEIxJBLCWvB2QKwRf6CO
f/+9jqf2ox7UXX5U7jupKfg8Fn6pIGU1vLbpIAGngkYAY9x0rm333PMrfvr9GMwh
8hg5WJ0i5b/PO2yZRllOoFqGhjgoZWCiiuTUoXzmgHLwnxaLjOXgxOF8ExTw5j1u
FKM5CRPFFLBgA4YnVhOP+wQ0yPa5RcoZfxoaQ/g0aQ93ynoNCGrU6fP2lTMp8X9+
jMEJKWzUKjQUHh5x8gb9sFSq39EvIwDVHKero1EPDE/3LPEQAE6D8ePK/bJhcVZ6
YSqPLzjlNfM0yoniUyDF0HNkirs8XJAQwscr3V0azQMuk5O+J/An5EhSbl9hdvfA
63+uUwFYUcK/i/eB299VRYQ0qdclx5K4hIq2GPnl8RSviarefTDcAtepUePkI9P6
TQ0oKw9KrshrtbLaN5mZNJRJJVVteyV2takFFkpTSfHdvy55aczDEGp6tkcZdaZr
rcCLirHl9jFbbwqITMvnpNRszMKIbabEQU9HGfQEE09l/FfoVJy0wK+pFIZkf/sT
0qPjkotWHWur52a5q2eEtk+hveI5Riuv1Jl0sYmnzXMSBY/vk+engZQr47A4QEi4
FZ97M/WnDE0yJHWDPKRobjrcD1zcMgCx5a/4kuhwJLzhiN0BdK3wpHA+txmZoAkC
X27gJ0nzkCzI404YWdO4uwvM0KrKm13Y3dZQlUb/rLmXES8sL/ekhy/YaIgYSiqx
EMQ7oLRaVDXEsIyqweG9mb1cpXEVIlqJ5AxN1KT/fS+6V5ha6VE7MVgYhuHr/blf
I00+xc6ObIeEqz/GH3kfuNGFmGLItYyHSE6FXXfdbS7fza/qqWH+T6sAH1jK9OA0
aqva5Yl4VoAbaKul0KEuK0bAiY+S/QQx5WTRHQdSJ1iEgIWq+iKk7rCKvog6HMxH
O9t4aTvZXF1RPhonnqqFrXWO/hfPlsUIhaq0taETR8CHJOcGVEkK1BXH0HzRMWMc
dJDk3kBeU6n+GrWVONwzCSdUe7W2LgKXTo2azEKQCzrK8t+V0xXHUg3Ea2szYxft
GsTafW4W7EcagLEci+fONw79p8KYAYA7SlTF52pjVqf319+nByYlKVinv8n8djDA
b4NQ9TpRo4jZ1jV/H30smRZeLZ6tooMTGHqCCMo7wsKA82B86ws5yIU/3qykQpKY
mJilXb/vrlYXrjHjlo/4N9ZAUy58Ku1NfQbDYJ+i2UibcBVlnR8XybQBWyjvnais
tIBJ1xyDqrVJ3359YUkF+S8y+N6TaUMOtI8XjtYPpJnp3i5k24ZNad6Wr/7eMHk7
W/bOQORZFKWWmfGPFYLAQj5Lt25d6uK4USoEW4SFrVmNMoZJi3adLCGSz70P6XU7
gjZXJON5lVuqXktmGVZpxOIvOZSJjQ6LMzC+sYVEZI9GFPiMgSsQjWH+TZIck18h
Sn0pGthyl+PotewkdsEeJLCXZgINAdkUKQ8QaKjSO0y3ck9LeKKCRSAysh/eV9WA
J+6xyPPhchkCL0Ccdfu0ZgMpTyPpWYTn3iyP9P/BuaUZj0keiP4y4sJ/tbAFCWPL
rOdvIf35ufxUDoWijUPPoXclBwoMrIZpZvl+Rm/TxOL8F880WkT0ELl0zgK+rRll
I4MFy/3Yr5iRInBrZ7KOMPtpbjQKJCuRoeUYsdOpqUzxU8wnpLvfPuA7UJOWKmQI
nzbSg6+ErIjCvaq3vgb+jJEzSVve2zjlmtWU7uIPntlntpArZ9goWx9k6AHM4K88
hombuD3gFRk2MGOAdczY++IIOoOtDjK0UGpp4e2M7oRg6o3jL0AyNLg0smwu5gPu
cgT+j8Zmuom0y/0M0VEEqmICP2k8l8/oPNSkM8SSRpATBpVk8/FKJDZVto/qdOWY
bNyGWq9ysm98Xfh1nZL9R06CSy9vBPInJacdhjP+ViZ1/XzDDjEys4GhcXaJXZUR
wCEtpH/vCpvTi8X1CxmsW58wlVPPmwyUShaO15VcagCm5b0BMI3gJV44yf6VnF4e
i/rjAv6FVfaMAO9KrMEIOsKfr8rGdTdDhtZA4RDsNss7UNPuhDwlYoPyyltD+p7m
tP0e3vUXAn7OFZBGdmoh2pmzQcZelf/sehtZc67lm9/Le1NymHZkrAQdSmdAHTDW
eR287PfssJS19EI7cf6nS16A/5VTnJxmqUaf/uM9VlDogtJiDUP2xjYLK3YTydxl
V3O6994VkceQXNf9C9N37rdx1TVulJL4sUY/u78HWDIPIbGnqvjWplhIgud/cjXC
p+30ZRTc/9kKz7ZCXK4MRO4LP+88k6Tr5uwistHpLnaIBMyU0TJzFkcpd3NiQX0S
J47pnovAt3Sipt2iRl7iplAM5ResyqfcFvY48OcaQNK32yuKi14yl1GWLz27asdB
1CZpw8Yql4YqTt5B5kx5G+pejHExsCT2BSg4VNDHjV1fWkqrEIxiOWZ6IzD+6fQa
Vr6ha+rrbNeTRjoBjLYgmRh7nK1NxOrP3TPmV1rsmnIiMYs6mL5y12OK5EwwKFUI
w+S/u9MNSBomiHNwwuHtVVVymrLNwSMggLWO+Dq8eskJwYdkzsictlFH1d4Iksuk
/9yOWud94gjoYGj6dh+jA5jBUXzuF82u33zwCk957BYmyBhzG02lVKwWihJ2tmws
RGDrrg7mW6Ii3MyLaxpm1BkxJNYqWXtqnWphgmMlZfeOjVY6BNhN5hQjHN+yunEw
CFw54Hnvo5Kpy9PycqKQ2Go5Wi0Dar0+uTsApoUhcv/s42nouYaWaIxxwFxkkBvZ
MjFa6h6T1tO4ILo8sE83dmVpkEA2UnHS2mE+cWn7YBCaFunGDAvZ9BkaIcEpOnsu
P/1/H74VRcAo1kQl+h0JvGQ3H+58YHNYwFhMoope4LBlg7GL7RAOwz1ZIx2aQ6+x
/Nuvbey9MqcdW+c3+jWoX7Nbj/mPprYYVPwehovWHKqgUkD4Xop9SNLdZ9CMy9mx
MyYTtrBjW+zbzR+rxiRhM3Cs088JrIYWyNRj1MUS9dXScH9gpqUTEwsf7wD41RxD
Quj6DYF9b84WbKsBrvtT7rixyArS/NVh4Wu7+kmuuRHqyyUh3/miBjFjaNv02vR5
OqIDLgn0VsWbV/7R1GsvEpwCRWgTDnWtmKn2HbEWgLaGTfctoMXsdqCEs8XRxI33
3ct6Xxwc83nnEqG7IGDIWy/PZzDeGwfHnMlrJ+6jIQO3Wdt6tDhkinwT9zOauQ7/
KJ9A9fJEVfMagwW891Y58RAbKzyPFY+0vsOTtGXpOTSgMWGPKO8ObpMBZ80N8xr3
IgIqwE1ilYNPQKEG5hCVvTu4Z34LdZVTVRM4ZCWDlfNIp7JYnSHkrZF9pjmKiGk6
Y3NdKzrqpPoy2qUZGf8EYO/c1X2MbqGCXFFoyn5a5CEyzw9QdeuSqVXqyq43WILG
2dD70WO+cya7M6NNBLcy9bjDfa340RZGY3+/aZ3FdAdF+BDl0AIr1KHomvBzlKMv
EPhNtiMulY70zGfrJBkGP5EmkHuU1PFNkEtdLBQEeXfcy5EZfw7Vz4I4P/Pf9TYp
iwpMJ6QJy/GA78wIqhgHZ8bntlGg0TFT7aaNJEL9LlLEV8mf5m0cuOHJcYghfRzg
izwJFu5CNwrFn3Virb9/6ARLBz5AF42FdKQQ10LF7eAuBB7II3Pga2oXRHhNAn2t
D6yfCOorMjofv44u2zqFCD2SZpG+4s6M5TF+I8X5AIUQO9c4/rTk1ezckQbtWJCm
kX123DLfrvA5hEKoNd1eLub4ri3Fzwkzi6eaV9EyedsvnHyhE1BRVjNAHfYmP4ry
9nI/IC3BzGOmwOuWzVU2FsEzsP2W8ALGNi8iK1/sSZH3TuOznErKw9xcEH7rviz6
RaVbA1gwPiv7+sg8IAsRPb4YORGq3IL4nKk4LIuLPdKqr1kma+HiZfD/oPXtDY//
Hw0dZ6eN49H2sufi9Fj6YNU6M/UBSwZXdTViG18N0rtnLACaZcIET6d9EK1x4KL5
klY7EBrAeORmRm8x3IZlIIfmeIETxA71LssRwJKe+SSHbbPgZj5amKxGF7Jb2TQt
iZWrDfalnIvkxa41ZX/oV71T9F+NHZ3//ZeS4ykdC+IjxXpVpjVt9DobUcjGmQPY
EV1R+T7od/vUC5zbUcwhjX9CiQU54FLX1xXfab72LkkWt4BhDXKI0gv9rpMFmZCX
YD3UsBDi+oLYyPC1rtcwlu+qskY10c4P9WOO7B8EhlhRWYHpOF/mQCjmoAQRwOGL
PiuRA4mvfteeAf1+GhwZ+P78ypbr85O8Acx1jmG1jlTmbEa97igHYBQR9abyp7cd
SafYauijsx+XpUamD4KfgA9o/jwNDt8vOC2nWkA+sbbCRDPb3ISnZdVwe3HIy5zo
tPGGoYmDc+fOFf2PtcCzPETjpHYtR2AUJjdoO37BdkO7EB2/FO0gbYp4Bv/s25X5
3kP+QxnnLke0GjC/ey7BcVTvP5wLmde3DBFbCvs9ccqSrs4zT2JHrhBb6Ottpz01
DZSbZYUJTM1Si0porl7ht5G85Y5Y4B+uTyWGUks+hUdhr4BUY4fhcikbhfFDJh9Z
y+L2a9uufEVCpwHyxpcKoy8b8uOM7CS2OPOb8eyZR3IMkEBKYuMxm+ToHJj1ovaW
6LEcEEW9qggFLV6ZPwFsrsg5/8y1ZISb3k3vgUGwZK0so0LNTf+1WqwdVFn2+bp0
OaY2z12EG2DTlH2i9WDK1fMSbaVkP6p63DVgLtmyJirW/X5dRCxF9Vfa9nJod3V/
ONZ+oyAnpJFs8Spgza3SoeVz7swJuS01ElB3tqmVYLm7wMS+Nf3HGcNeBgFQo6oD
/AhyhlPOZG4fXyC8Ah0teZIzSWD70rKvN4ouKt+FIouYORDbVsn0u5dB4J+eInvi
YdEnM+5d0d9JMI1f6eu3hJpX58TN1i1f7aPXfGBHG3WH+U58zp1qWxV9d73TeoyT
ASOqlEIkfzrroFN6AM2J8AieYkjEfUphnBYNkEDfwzkn38iDJmMHLw6JmVwDjyTQ
gF63YvA9WlcaSL7wBvE5I+R0jLNDPSxkjuh6g6foclWiyEEyea2yyj/nd8A7hQYL
/QoEmLCsLmfC5ijEWvslHARg4bglFuDPuYAi6ZRDfQKGHF0sBJh0D19tX9tLGLE0
KPrveX/kPPtFYYuScwkj9Sh8fFhaGpStxGWuh6+rEeGmYlxeGl+wxfCSsQyw3Xu5
aBvO5ciIkYzlSPiBL7EVFeabZkgtjMK5hMJuv5rjMrPNorfkCLEDX4Zj0lMOvhZ/
PSeP7Hbl5Ort0NYTmq3AT8d2prvE0zDmZJk3mVSVgOOsIZ7AxQ+yxE6xhStnrIG5
/cjXlanpk1xjTpDVkMLImYlgOfmCqbQrcECTcsJwppdHElZvnsr3XgaFgaG0dOQz
fkQzWH9bf8t+J+rVlP9S1guri9kCTu946QzoPM+X5E1MttF48Ni8BozGauMWAW6q
CSosjfz0gaX2iTMjDCtmtZNKw53/LI5i4isLb4rQAk2h2VbJ/BnEakN90/l2+mrW
TlaRmHWJLvVpsk8EBxF25Iq3XYuwT5EXwUCY3gt4dqeNeMX25IOcfiZ5hsSXmadB
93XkZTD97o63Sbj0C+HVGbEZQoB05my87vAlhjXty3ef1fJXS9Jelu4TJNBwo+Iz
6G0zFlPH8UCtwLvQvmD9AkdUUL2KqkyJfZAkbLHzk8Ww3nhsU6HOhNrCvJFERvaq
WqYplMCsb9YkZHK5TMQDnzX34ji1EIDm3NUw8M7syGyQp+j+o0Vzoa4zBdU/B6nD
v3UbtTwPvOpACtdPfiH7GXWcI66XgAZ5gexbQVOFOGBqlCTQHzIPLrQvWMU0d5oF
/Y+qReDwVS30+RMFMxSRQQOZOG5TVAPyAGQRfo8K4/9wNM07T3he5AC5YH1La6BX
YbSjzExnT08pW5SZGLtvU/U4q7i+s05/nuE5gWyF7Q8uQEJKFV3VBHjKIzFQXBA+
0xmfBzsuGdKFQofMbvWVUGfkNIbA6IEQiaSUsYpcOAVFJVmnoL1ZcnudIdRpb0uA
70Gg/jfJmJQBkHY7ztYnrg5XpwvNyoYvz89ypyjZGK+f/zlW16U6pzc/oJ08LyZ0
eeTQxBJn8sGWycF5Pk3mMEgiBXrGqvojGectPVtEbD33CPIa4KiXLhXStX7zFVqP
oMt0HLXYU93BCoBCFg5p93+avahjF/omQM7aDjoZ5JzXuZ2H09Ge7QqUjlSgYdAb
DfrgYvOVIaN3yyBzzMCFyCYnd3zlRHBwULgM8tAA9/5vpqNz3I3P7hOKhNtNDrl0
XcTPye9FiWyJBbNHj8vEOwtTPV5SLnGWrj1lXxzbfM8W2FQ1kQYFydVtJhGxSDYb
TUdBqwsLk6NOQRHWYCtgi/+t1pkY0/6KJA2EV0UFNugfJ/cj3i6QAEmRlH2LovEr
42UIM8cHjN4hEa1anNM0ZcOFbuA5ZWYDSc4UxdK1VsXS6EoFtAH0uMO4+rLtabFI
7iiBIx4y71Ecw1JfVz6a+cUf3rCWItU5ppzoPEHztptI2QAHi1ghWxmnPBfiuFp1
VxtU88a+zyEXoRi9ZTp71VLEndgbE0DaTdffi0ZKJxrQX1+g1shmQTcEsgfxecRr
70uozuuTYYMQCn1AVoVo2elSmN8clg2GI3gsoIMLWzObjs1wYmNkvD25fI4RV6Fo
oaiCjWYA3FQt3ZUj410yljOy5D0iNTN/amd01AQQxnw7OAIztX4CF4fRKxqOTGJa
zQ4iQHYioo8lCwOHS30jHBqDqcHM1uPy/wmog1ra5D2Wn6x/fc39HC5eQrVWBTIS
1m1ppcyZZa92/4gEggbICtM70PKXqhEVN1dnaOVrGqMhJ8bdG08SF9Gzrtqs1UhS
8TtHau+FZhPZkdkFZDAlFP+IXQeX6TWOfhgqgwwUwH6ZHKcLi6Abazap79At9c3E
wfy/S3019il5CCcUFWHuP9m3t4bJjBAmIsqXKRvOduyqWSx+68A7ihpiZU61cmKB
CZYJbndrN75JWFE9ezdFFuQSrCOH1nkUdzlgGhpnIUbOv8xSV10WVbVviYKA2xo0
A4qBTAC0loJL7RtTTkoAVBEzyyO4+5TfpAlR71d1ZhV+KF+bo8NZSgJJ83IGswPQ
X23Ql31TzK/UadJKaFdP2/MN4SyycUP+07OjvAIe3al3zPHU0DL1aWXolrRSYVrX
IAL6VAPTwljayT9WKgBFqHRp9c0RnrG09DJbsxENmvgbeV+P55uqBQVUa0PBuJDO
hIyeokhMLNpWHZO04kmA8PHMwdjtgApqI8UtV3LjxH8L+ggYM723SBMcPN+jOJGo
PVoXg/8/hr7X2S4uefuX4zqEv9KairJ4/daLTjVVqNZV8IR1eBZAKt8EIzkPn9GD
6aZdLK653+s8/9r5RIN4qRJvkm47Z10RI1E8Jba3W1zkUtV0JylKc4U8p8ZWQ1a4
3q2dS2zoMwcCjgFylrH6pzbn6kbHnwdkD/xrpifhoKUeG9Kot2uwwRsylFXzTyXc
LloY1chjitJsneNhr0AE2iN2TSjYdbb6uQbgTOwtuM3lKxXYb7CFzbmu0vNBW7XN
V1EKzo8DxiMaNv/Wr/Ae8pPBLTTdAR7SsFfTVU3JiguPPDzX6yEKwDZ/0BAleOZA
ZFwbcQ7xhGdBbSIH6aBPmjid3/FSsO46tfbkhWghXR7oI4gXkF/SzmgIM2BtlSaI
/sLzVzIJP4dKPSe77ZWI2xYQMHX/Kfv7qHDtP9XrPYLgqv5M8DJ5etz7ADWBGBYu
0ecHxWx25s2o70SwinSMleFYwpz68oYJwH5bErlhtYBinExqoZzOrkKDWywCHjwA
50FD8MGl0tbtFcmYJgC4WlVNlCPKg27N+EapjEV9tISAtzFzDgdCZ9LWsPGblKht
eshrylOPCUGJF8PNcJbuUD10aeTl/un/nf4WKmbCWDQq+ojzGEmyBBTgzYWR8IjC
YP9f8yrPA7uruYrJrObl47qHpRdG3aJRWTdXI1FLgQBIBZU5uHP1Uo8FAg942BMG
h6DoyPTxwItyVO/VG5MwvxSWIe5MNJqXpCTbPjdwuuPvmYjO4WNIRPiaV+P7AtAk
oPCer6f/L+mi0OZUaVIXGWJaDiO9sY7QuRrPyGEiHgpO/Awuvc++xWxquNdx+ht6
hk/RrlzGib/QJU+gofp3mXvlDPL9/OyqeTzGCZGe7hpaOkFb+jvCsAh+pli4biQ4
FBhZ0rCj1UeJN6y4ucLTnlYDOedhSiqfiTP4XNtXB18t2wY5Bv+Yx8Q+LYR7nzwJ
qfmWdzIYq9RJ368BpEDTWHRuYc0FsKPZfGm1MZpXKfqmbqjhr1STs1eSM0YPpIfD
ir5U1A32UGRsNwOBkO943MX9+X8syPB9d0+Hn+JzLOgeEFLQAn38fT613h2Fp+vh
cjoVBc+b/HB9EbomsVx/WkydlzuXaBAvugmUiSZ750XGSLGVB4FOSepEYtbnRp3l
RfIDd+hE7tYFMjt0bSDQOuXxGLTlZL8N+2CqTJqrRaM74nZtj6WTF4siCcaocE0q
mCOCi8g5UaoqU67ptUeu/Bl0K0h5Z4+X+uI+WfDARAtPgbNS0RB2fU+UAFZnJdd9
8z19xFd0Nlgj0naIwFqvjzxp/5yy++9hsbvEYCfMxCPeiDjzbhfXadS5jp563D0k
Fb55aRYzXWmJYJJhf9C28hyWVuyqJMDc56RH4/c0tP5vQitRwqNsnQE6WsMOOwVX
ujwrzmMglNdERYWUZUhOnJY5dB2eiweR+/bq96SuvrSSdkZzBdVuxI8EGp2UCT75
Vu/xQl1xygMsW/KIsg06RLnnJFOo4uRaFERf8OecN8krL/GlDZupqpaY2e+GoYdz
5A4Vv4AsTuCJqpqkwSshWeoI3ObaAbza4JPNa+ibQIa0AiCppOqKK/Wf8nyPIoPY
LKhFpapxgHffWZ56nUbpt4Jy2lmcNX8mvN0ZMRuxdNaQSG+UlbV/V8PfL3XIjCbw
7ddK2hOTDCil9yOCeV2pLlXhLdHX2xHHqmLTU+fgN7+iPgXa0NZVOnwDd8KkfmcU
TEgdTFEIVvHmqhaR2Nff8Rx+Ppt/6gpe5IbwJEqWG9UMrwCjMwVv2Qt7hJcV3IWm
zgNq0riIPxgJ1GpPwwkq4F6IEsRazXX/e5k/u9ocj1lsPp9pR8RD3Poo5DlM6CZr
mfTqnx922gqkyb0atob6UL0X39e8ZVxdpCuvE2ymd4mQhtDiWrekpjwxEVierHMT
lsDqI4v7zgPqfGHbNrv68EjylP+gmyZlShEGevytuNYvZQbrQHzgUvrHXrYxlmz5
b2P/s0hy6mih5YRTwvc373pPkTnjYTsAsB7BuYkmFO6c4lLKChfnjaQLUAM+iTgW
ZnHcqk6yD7RqQnBkt6aPi4hgNyKLhVcgUhcj0Gb0YV6F2CL0QNi5zXlTb3KuRlKM
7a01Hn1Khijfk8aAmDvcszvJzYoe9x0IcXCi2Ry/bAVgixLNLkYmRPYk6fIreaMd
y/GDrCNG+Zc1kyXT214Dr/5R3LuBobmmOBIBgfOULNE9ScANAZPWarfoM7TRGU0Y
IXtlEPPo11Splm92GrbHv9ttJZxiOauoZ0ynmxKQQ9yrM67Ia2yfctJNC8v6gAo1
HKlrLCdSAuwyfdVQTeC/fF8Sla9rgxlbC6o3ez+JI2V1/qUOmUb381KmC3xNpKp4
5UeEoOcGail1RZ8SFAVv/+cMLDLDckVJ31Tq6mscTUjET0FGKGOuy37sjGJpFirS
WlajWeLSSWeveQvun5D/sjxghWKLmwJw6nhlBP6C3TA38Z6p7exg9guPioYL+OjZ
BAFVIw4wrQjvr0d41LK7/No63pVt+kQz9dK4rqwYxHSE0bQFbp+I0CfQPU3n6K17
RYJqSSf1r655jbd83YWT35BMG9kyA2WrVzFUNsTUgr/AkIJ4DxUVXpPw3TV8Si2r
BIGe/Mxhvzs7KbVHYjtffUMmpvymi9q4zvyJoo7hmgayqlGcD2RAQaUrxYrgoe3w
VCvNVkCyX84sRwsrVnmm9ncGSIbGRF5PV8wCnnBAOx1h6hH2nbTSDFlv3gCVHtCZ
32r5OcxIsOCJ9xQ+/s1Xh8l8VDYetbh6YdU89uoP1roRe18V0+z4ebRxB4155T5c
HKq4XTYZwYiqAakEAzj7JDfnSfcdRIi+S7d5uRM2aisFUFTU7wwSWnA/8wTyX7Bf
UxMCqB/8y9lWDuogjma6FgX8VUEGOeJWulrPYLUNqEDx1ngprcaSYHxQ4NgCcXco
C7NGXJudt5M8cJJr4Ii5W/HYKrtHzyDuXsNITQcWJxEFlkBGiNcw2UCAf+nPqGiu
UeQWU01SwsVe5MMjweUGSk437XV3Ulle4dQUDc7YOiXcfib3FS3QeaMlWqZMHEgq
9/ySCH8ImnM/HThQOMqqofTmAUNO2Wf3sxdCysU8zEz4Y4Cqcb4j7bY6FO18TrPF
inlu1QquSywOiNC0fcKdFGv5gJZzSZHBEK8z0CHGduQ5ry5jfqL33jgay2/VqQrP
PEpLEH6dIBEsHJ6+M8ygqDV53LC/bV/hvlXLcu4Kmd75c1rFEp7tBi2RpOjyFqIv
3SdOr8TykCqdBdeTuetuENWb7WsVQxmzI77y/oS8HnRFPeo/CdgfYwLlkR+f74Ef
xQE2Fydlk0dwQUVxYxoAyNuFmd9jPdr1qczpDEYmrwqnHAcJdY/w4jTa0I3c8bfX
m8VBQTyqoVMS0fP9e/wyw0mEWVXISlNs3QFDh4p7yyjteJr463Arns7+tyMVYZnW
ll++LXTm9+MvyPyDtboZGoM+sh3aGGqrtps49B2riSSFC7RfAMwX/f2zB8rUUefy
kugONo+KLuHlYoV7oNAsVttSo6imesaBKXHlX9f7IWHI/FrUzEuu5ryC0PYCfUJT
VklSjZkmW7nANlpRuBkQ8nRKvmYKsVbDZQBsH4dMHVshDxaLnVG3bXE5YKL23jFK
P90nh3mmKSeJh5AqFETbLg25Q0Wut+GANAya8QYo9uKHlPjavRdBOr/JvGXVq7mm
xtQGa5xHRGuTRV7b8xBr1YKDXebC6CFaoeYk3XfMIOAo/TxyQmeFOpWyn0PXPSlg
mvODPBa4jSbhCVs+QQErWtry9eaJVoY5ZKHvugbKRx1m5HIsPC96+gtu0u3kNWSG
42+srXInzVINz1jMJhrsW3CtDRn5GP0XY/A2gsjNVXGaVJfBeuNzylDjMzxqR1sF
+gyHLflyK8f9Oo0YFKBu18/6RIUG0FsjCjvz0tSiKTeKHbaMEvSKgv60djXaZf5O
W728seIRqN4V2eHc6XvbGRO3b/2BN6XmcyHCy3IeF/ujWwC8Rbaf04oOxDy8BFgx
fV6etDdfHKJ+Wrh1LvBwApKZd1Qg26jmS3ouquigmdYBALzGaoOmU9W6Dy31TUXR
aAncGVhfaiAavLgdk55ZUf4P043XZwzCmYnF0QSZN947ciqpOWJZYHNNioUhh/rg
ntcVFyokUQx4dXxvjUnhhhmFc8ECejvwkSmUcpSAcg5W4x6eMoEDZxuvTovQ2pkh
U7Rvd/yak9ZBkpMEHUlc3MLPbwM32oLBiQrfi50nbjbjzTewl0pyy6d2MuAHQMOT
n8/n+IK42xagtdVqpE7veYSa3CRbfWwQglWp9YuDWDwJDj8yzXY7J75X9HllVSdX
PGzjkvySaLYHIjpEx+kG6K4+zidxtlQKULrKtlv4YefT2HMhuGd9U8BIp/IfsFmC
fX8Mddsj0allIVyV5Oy6XxJwbEwmWRJiHtzil3CFDdgevIefR6xT+aJeDFE3c7dg
Swxj/dYKiuB2yhSEVciWg5abwnX4eoz23/ICQ4Mc5s+/CeXO+VUtkW8bZT3tH7bv
TMFJzhI8/ZbPtd/2A/BHY1qiRMRPC8mEFy3AGz8kMl/OB5H8PzUIcOFA8sP8a9q1
pWAS/ZG7RapvG+3T2v8ftxxr6+aC5wHoTvEkYXmKPOgdDUrFZaxGdaDV5gAx4SLz
RxHP7F9KK6e1p2tSk4NVo4dD4f9aG5q36v+xbx9VMDG9PxNG8TeA8BuMKBaGoNs1
qrXwKGNZPWDFf0TL039MSEDe7OM/+9yR0FZG0wxh90p8FIfvU3L/XR8gnmECDRUO
hN+xsqzb2ExdTnavvSvRKTTnfRAd124RmcIZhqt0vd1LPTda/7JtwFYweOVK29xt
J2cOdP2c3zoH/WRNA+KelyoKc/sKo7jZDhZ/JJ+IBxQk1N7cBWRO5g+k28StTyMm
xqADf7Do3Td9ycmC8iZoNC8rwN0/S2eXreTxb9uaLV0Ctn31hWGeNOTLW9d/y063
24nPphGYbIAcoz9PIMLydaAkwA9hY6DusYDxaLuv/nPDSKTLL5uam/rTV9y8KBQQ
Yi3vIBJtx2YL9snlwldJgiyxQQfyHeIHy/2cXtcDnieiqpjGYduBYeAFeuPRVw1X
e3UCTozv6Six7Zos3eis3RuVTYt3Kgqso8wLpmo5HvjGzWLEUDU8ZXJvDmeFdU5s
EGkZuu/QOmSfdrv7CHICEqFIW+hCwDx7MWnOBpyVAfSmDRMJRN1W9OGU/tn2Kf0Z
8fD4VsqRFsPGYNWutmL5s5PJ8a7HOAgRRi1KIn1XvA0nBit2QaAUCJ2cGGzjSqOF
H/8ajJ9CvDj9T7RvMiFrAfiSKTWjKYoUNaYdka1Zh1sbP2Rkrjgp4CBj1veNmN95
3xRH0ahAK5UIze1IAVJwIhEhLdmYuVPtdwqVv0gRmrwtYkZcNPZ1JGeu9nlkBXGW
GUljNjK2s0dFYwBGxo7Ylnuk2dzwOQa0L9s7GXBufIxJ4ojMsjzUHqGMUn5wPm7n
RtF8bJoFH2wRuMS4qngNduhz9WXsTPZpLtA+nMG5b4qfzOOIAkHtN7cefU/Gpu/t
MpK4kOyRBYx9Jea26ZUDPiMQdRmX+5FtOa6tvvxLVjsck6itUb0xN5gbtQpDTYjp
KgdCe1Vai7mJivqBhiK4sxlQDdhQKQnT/fqbCQdkDSGHm/dfIs0dJq0NHF9ICGw/
AEM6ERwrqz3voLhYKjBWhRg1jKVyWYeBs83J9LMgv+pbYPJNzCkGI/+CBQy/HwIo
SmnwdqAcvqTxTLu/OtvEuR9H9OdAcAQx9nfknkE9MWPeQb+3C3z4CfuiV1jH5jNv
RyvALWhpWvnBIxW1Sg7yrsFdvLvTKXniCAZGLuQZB3WiE7MftbQ50sd31k99r3lG
nFRrCq5czP8P04k+5ILkBInPI3wZ7VyWVJWnAhlJlOxghGZuqZA4b/hBPwrSZ66t
+hrvA6f0IRzAVG70ZcbokbZf+0XkdQpcT5RZO3e+b5QTXD2kTl+1m6+b4TiS9b+R
ZHHT1pARli9at78f6Ac5cBUdTXApPRaOSTFtkwxImk7ps1lMvBR/mnRro1r1Chjs
h/zzfGH8lsDOeIfCmUBLkDD9RuG6tlUVADVWaKCtxNf0ROgqWuKY8Zs4A6XBW5SQ
Lp9CjnmnwaKCjKddgzB+aOoMbyESnoe8S+jiPvt9etx0TyHRMZ1Qs0xPUYuuHOBs
Kh7WSjU7OxKC4DfkXnfeiqCa2Q3ONkmmpQcAA3rpLZkwutTRdknI6fwJaxCGj1WY
akTQl3XPnWy+tptYWBl9OKYpUwEC2zB3Q5Mto7JRhhjy538Ds3WTZehtGewT0vBb
NVCkroLUd4jeI6k3iPNJomWqmgxSaGvVdnLIfVeFGRDfvGyunNXJMMmX47eRkUVa
kP8J/PyNFoUeH24w6HHLgwBBYcxZBVXOZYW5cKCO9tXsfVAzbdz+cmiV1WjXLS6i
gTPZ+YVUB497a4Sg/EA4DuIzCp3EZ+mlWyf5MzRyoHDh0lXfhP17UYMla8HGY6DW
ojy2nFq6YVOY7TPFcr8ss+4TGZ1kP9wiowCuYhKjCrDic52KvWyA6Uhr6X91Ljqw
+I6+2PvEvaGGosiZ2vxFBeEEc79jCKBXVTXQ9nNCcEP6IVRby6Ok0I3gqTn4QDv+
UWloRcPNV27IL03VsAnZyencKRhfEM+rZ9slKOkjamBF2MbChEQWW0rZPdhO9jxX
LFf8chph5eWOI91IUs2AeXMlNGNWmZ3jxg0vLpNRjThGj7ekepRw597Ww570HmJN
URLrMP+J/Rs8vfpfP4nUXC780GM4QncNOnAkCJ+GD82IXdNWPdouTrFe4MG9tOod
rZtnDvheK53+z5wfo/8iwO6qTLSbvVUsgUj74UM0uoJee67phbKR9rNyfwsAszy4
xHwAZe+S032tyLnx5A5XqtizbT4Xkd+jPzCoikzerselrPAC3zaGQduruSFtFg3Z
xPpE/gwCGSEWuNY0TN/rbaS6J7f4EHHNeidZbaz0Pf0nMsflEiI1d7BZ9dyn490d
sM8gI84kcRHSXjpR+Zs93Q2ZviioGFbgIe/lNDJAhOs+LbyUDbvMbOKbQSp7am+3
gfWgkCEE+1gXZf8ZEyisAWIZ9j9SRBumPo1qS3Aq+oz+eYA9F6LBrGsXlEcQL8aS
jkl8SymDJNQiz9EoI+GHSUsVjkdme46zTXOSz1BEw4IW4yQSoPTPduPOsU9D/ABh
heYM/jbPlSHo1e0MlvwEbjRjnFJVmShJyL4/jPqGpDTU7/ZZsEv1QFpTO+eZxWvl
Q6G3i8XuUJkibGg14T0wCo/OoFKBEWuHfu3bHSU6N74ji4ZriHLgOQPbcIZBAFc/
zjMaG4LjS3xiXHPiOczXx5uA7fJ/ndPaV6J8S9y70xuBd6JCEesCPkG3flCGEqAH
3/AJnRKtNqQ1bbjQ7SQ2ykWBD/reFGaA3ItryKkwGY4NttUI0OYUwhp27uzeEPJd
BLYQ5MRWP2LxSrrhZaJSbKj+nQUi8vrRGJ+N0+5oDC8rYGVyTrD1DHALM4cOSjAO
8iRT+lTjNzQmgiQWJRdu39oBSaHuXV+fnKKdJXSzaB+ioOyYdN9n6dRHdm7MgkCv
IFHIy+Inw7WPMud19bw3Zt+KEZVVi8B5IBYd8l8FSbKCOmmBQe5F7acmzhPB9BKb
OYJIkXznaOsGyqARvIPfPQ84X1w+d0I0N4ScsPbJopZggxZVqmkkmVCyd1f0KSwi
gtx4lqopU005FTAi5CRdTanbtYM5SWip7ZUKMRr8lLjjF0oRKwI/a1GzwU9uBu8b
P/zW+qOPxGpQPtE65hp0VcCCRmCVAutz4X9cCvgnTjSPYT4TxvFcJJrCxlgUKy0o
ENLlQkbYgKaATItqPp3Sg7gPYATK5NQWSQ4gw1SoVTfqfEy+9yQOeRsWcjZgO+Ov
IkSH5ijNUhQJGpq/XOmS7bWDrKnYuoBYIedGKG4Atz6wa0tZ6b8HrR63BqVHvgqk
H4gJo6Qv++cgeBBDlkqp4jktoJ09B0SzKBsZvWXSvwYKnQhKPwFwxqe7KTO9WwT7
WjuKtvV+EkFFfVaN3j50KBT+C9aSXBr3yiYNQaVi1IqGxGvVmGFYXB+dokGQOeqp
0pGtoz4UZc0TSmc8DvvURJtua012kBu2e1J6Qh5gBghq9LWJte0YdwYEaw31TWwp
1g8UsSnfbMwjqHEfVGU45muDvvIQBKSmiX9tv3Abd+8DbEXaJfBAbxmhfnOo65CU
JywZ2mo6M0U7TLDvueaHI7ZMyMJBECzyqBuXWtWwZTMUbBhrb+T5mPb7KTw04bzr
h0kR+qv5DB4N6Blle8x5gBErD8cmu9eE39G9Sx+nKuJOZGYU0cKrvBZAkQu69X3U
Q7xfpPBUD+CvclrSRdVo3ld4iIQcYrNzY+MJbzlvTfLIgAnDtncF87ouU1U0ewpU
S1bNpylc4ZTQtZZgWNi+qpuAtzrmhEFJ64RKCURlpEULwVJcir4dXag394+BE2dV
fqiZKO4S3UulDTiOY+gNGL1mYRHWd/d7TnCzG3wS5pZx7YXj5zt1shDcHqTmpKOc
VydyML77GKslDmDp/BVOBHj6CBFmfZgsJFYcGbdRuDQeE4xuhkayfQldMeoQleMW
uruwLL7UARH3RVlBqbKg/8/nRh8fOHf8t+eHu143TQPOW34Qx5x/NxdsB/tA/vuP
LwVXpl3nDKddcpKsXTltM76svkSuW4VYcEhSdszN5/g3kZAG4ycqAYtmojf6m9dR
pEhPSl1leCBx3mHMs4YVxKdZazPaPYrmmAg1r7KQSHOQZz8Rsn8MiaqToESb4+Wl
WOmMoO4r+MsjJnDEiWFynyITr9AgYu9RPy0Hb4roEZXz5eZLmfv/gqxItHUhIYjT
8exdtGrwksGSrafrewbrpI3YWKFgDxhM34MhRJmRAaL6LPCPBtt/5vme7rxBWEGk
e5QrXdEhZrDX+jFV68DYi/KmfTp1T9GDSfWFnzAvxm1gIccdR/sFd+cVtUfi4rZo
dOrUdcaTj1f27PiU1d8Oe5tjbJbjn79T7Qk9BgHUMWiNycNhdrTXZgv/4gFPyyyV
qud40qeeajneJC3q6Os9Cl5zra1dB6aE+JxD9PPOBbUdHr/nG6v7SKA/ugWNsfAk
7hlB73u5cM20/6CVRuPmOcQL9yH3KNz3hRjBamTKrWp35df+LA20ts3sMpva/A1b
iz/86bBPVEb2eW2MFjkUjTDPXQvY9+p/mNDz5EOD6V3vGJx6XinLEN0tpODPy0dZ
anUg9BOd6u/A9mKiam4QaivaXK5vYvo3qp24AlfR6X03z8+HwFZ3RJSPub7sX53N
QU1hPTCAzWobAAlvp1JYVsAaxsqq3n40bOvSGISfI/InWZjFUVR+nOTzDD+MQZBi
YEKcWEfcy+b90MluIRdULq5xlibdnEsOg9os99uc+CTXxmG2//Z13HcCrPTcCPU9
8iXkaanSnbSjysKElfR/ZK/TMAq6h17oi0CbhWZIlJmDZkuTx5O46EihmfTvqFfX
O/8PGoqgTozlVrWPZfPrPUgoj6CLYzZ+zaq7TiIOHw+n9YdKohRn3eDQsD8dzIJO
z+YRV3RE79lmCdbQQaOaJgp6PbNH43Qu/YrwZoDfkt5wGHexHf2eQ+9OVpFEMfjK
0wd7NWE/QCm14obMsAOSFeHstUpz7UoIvk7498OgzeQi3FrPH4lnE0aWfYASgF+f
3P4kEWdeSrXHsjhKbxoiKsjsmAHABspN4e3KWfBIdeCBL54ZTpVd7v073xgaWErg
pOUApjMkanDx7TLGeQNk9ZxmCD14y9AhKbP1Ov/xVaXZAYI/9YUdQYJCSti77QZk
txOX+6f21BwPltkKqDjaj96Dt63iTnocXI2+D97woi7ovlBJUKWSgjMdKmGD8/g0
fbdICYFlHZOvhxyEfjWIsMoxp+LU06orKJDjmC5llJNhwopwDbFko8PKJ4o2VwCS
cBAC/Q6ue8Kv/pP6Zqr3hazAs7ch/OXrfLs+uCEVXlBcTBKRWyY9V2kslJpTdm5O
GdA3JPGQDzgbPF8YxxqXtXAgvIDN00XjyEMhw7ypSAQaZCBaDTTF9GVZctde5N07
dhDX4aAD/rDnTL3VIQN6k+bS7+1iRIUrbJkSUW5gwTx8IWwAarYbaR1HLRqVarub
Nk8BSKi96mzvAopWF0PL12R4+fzM2omcwK4ociOL1iLuD/yxE/etCRnWaFwZia22
uCcHmrumYbOliF6MH+RfrI0UFwR5UU7o8+9MdUYBgoFqrW8goIWoU8wZ5tasc1I1
msXhHvm9kE63QvPwpiFdfBHh+bizcaHTVG5cTxG7SZK+T1FVwClN3xORtPegm4LL
mL0XO4pMadqMPp2IIKdSB2Gobr0xh92B4ed0A6focOG5D6tHM+MqtxhOtav1bmjd
9WMQf16xVwFsUDlTGudhnvJiVFozrjH9AdeAhWi0yc4XgMXopmgWNmeQ3o3bod/U
DDsCQ+ZSJ5jaHNixeJ8u4hFkuL3Zu1gmYrH38QwF9JtzLvhWs4jPGJ9HO3SXdIRT
1yw/xSdXp2z7Oa62JIHJ8Q4ph2XGqB2319IUDGs8EuHq00KJV8kgJoTqu6hi6UTw
lT7wUbe1LBVhwwp5Lodk9UzDKM4gZBkbkETQ5+QooDIbW4jzKisF8wNSuoy0+lgH
L65XWFWoielzRfKPc1t2GfAA/YxDKoJr2YRo8xr0R3QhnxDgB5Q7WwF2l/trxj7Q
8ApBy3dM3qY1p+6COaUQ1+jqYdSOa6odssqwVNtnlP1CnkB5cT183db0r1qUJp1n
hZCyCkPIOvQgk/qAqBgxE9jnK93jAxULAOROaEojeCTRTUpqVBuz5XRgE8KIZCVs
cIvKdzC7Ijq0+xvwKfxDPpROzIF+E3VCuTem0/fG+ua9/khiL7w6VMFCmOwWVvtT
8ZePb6X8+JAYl8DYDJtThj3Vv9ADJE6tmRlS5KDlFbqgtoahEtBp9E2ASGvxiG/w
ddLsGQoJ2SlmnbIAYJd37wTREOAZO0S5iVAHrUe5bRtCl+8b5abOVYt5ed5eVqjW
Xejoa9DBww1SArUZWevSxQ5JCnv4ozIdgV4a994RPs0YFFntmuAv5iVPF6Y+wQum
udbkSWSwcs4dn8fUL5BsSBt1oCNUO7wOgGsxABLCCw4gixCkzaqoYf7a+snbp5yh
DJVjWy27JKAh9kvg52XSNUAgbH8HWBfbJueRolntvO8SPL7L5Bk1MKYc8tyDWEQo
aAr+4pD7qYsXcudRLaYiI2SfOc+6ikkEVXwhQorFOTLEQIxPb6c7LSqu7WSWTcr7
dl78dRokUETKT4IPqUfLsZaL6JYflm9Pd9I7325+zJ7KEmFBiHGEs22nqBe6jswI
U7RlTKUuQPEL4YgY8yZmb28lKwXz3bg08xYJ31tylPyJXLysfMw5Zmi+CPWbjUA3
X9jm5r2tDsNymE0BFTvFVCis31d5DpgS2RF+2KhFPjxDlUVpnvRw1fKhn6vULgyL
wAxsRE+4EG3mq8WD8r69tMcdQ2tw7ql5v+ZuoClN82AtoJKPNxjJwR6p8t3RSDRo
iD/4yM69qhSpepjfWJMS9Klo1zffc4VACvWTxKonPCUwxGMZeLLTpjuCxZzUFG2G
29AvPa2rZEkQwMrzgzhASffLiTGvM8IPLEx3RmxsxXNnMm5qV07W8IZeFLLi7+W5
3ThsAYp3Evhil4D0LL2SZChaJCdEgv6I3QJjDmCSeawXL3loSsh3X8iLvCdGV5Qc
ow3zAw6Fsm9HPID3126UFf+/r2EjzePHt/w9Aq6cAKA+Dzrj+oLsQK7AzOpAesuG
ru0rlfqYiZ2O3idJqP9kRiJlwdzlpvXDRSCTLRBLdI6gap0Mc6EyFQZ//5/tUpGh
qFtiqyO0HO0uK5/CILhWAA1SBOAN+4Sfu+3kOLVYTErOb6Pl6LQLERSUgkgb7LRU
LPgYsFizy9cc20lyXgp3VguNRTNysn2JAUxBntnyPjMnlXppCFojHoGCy21kVzzF
ue3zOPCbiH2yVZlusr+Pff5Vm9Cdo9juvte8rvlBsEWIIf5nsH9Rrpxn6qQYO+iY
db1KXNgyIhACklLk5BIhhdthEldB0otbznm57myjF0WQY5wgnwlprMw5Cpv1qTrD
WuLIpybHsRZv8l8HHLWo0N2pJjwBo7+8fRZJa6Oh5ph2N02Tz6oPyFSI5mi6p1Nm
QpyGKb5zzkZYYVOkjSLCaXztC2jb2nR9cTuicsIRBW7zs0mlOoyPLd/ChcCJ+kC0
QUauutpcPaW8AlpldbrwIl9UaXzx/4VRso44mevvdGXTAgfdWUz+bzesdPGEBVok
BESsQPblgAdPtAgpE6iRiczsIo3fvbS+YE76FIMr/PTHSbUo0LXWd/jtbtueqWVd
dyouil83ay63vkn8MgYqV+Rp4Ya4Keg/5bumtP/ktTG+VSlh66yzQ6765/hLzT7Z
ESsyPH2yEsVcs4u9jZznx62h9O0gKulxQOuHVGoo10oGX31UBIh+rIQMiMsVRzsr
0pIHanUCUeejHfK9NR/JBGRO6CdclI6zEkrYe1DhamncWZteSef53UbVkqbKKSN3
bHatmHWuC1oY4w791fvixW/Grcn/4KtilOC1FjJEh8yJoeMlpAL1yUUp95iL6GEv
bGHBVBW1akqzJVDpLSAFrVj83a8u4kRg2CXciG5iMMghF9L6JEEp11rDBuyUiSVC
jumiXZhzJJ1tPcDbPV4mkhF8k2/1gPeuPYG36gqphJOm0ttdmxPPpINbg2R99++A
gnhGUa7Za6yffkysz0iszc9CK5z7c4Mln8DYDAnKpL1+UMd8IXizuHraKGICZBKm
FFnt5WNZ+/2CBnR4hL/TL/G83vbkjFvVyr7h+Ji/hv737cVibaLUf8Ay69TVjAre
nkEgbbZ1H/YcDkmJ37xUlxVT1BFy4tB2MYZMHsJehwU94uPe6qeLrGOvhnAqNmFD
3XRGxRB6CYMxtWS+Igdyb0TYohDcNvBDPoDnbsU+8+y5Q7WmIIY1S9DP940pW5T+
4qWTunGgIP80y56c6lsmPVi38sjUgGEh81HxNvQf+4UveQcgtSEIT5GhzdOFIAsM
mPmzMUxibD8rZmG7DRVRIRPNcvpuLkSBJr0uOQ8vWzmioSao084hEe2i1Drmp9rk
woJy1z687zZ9bREgH3wJJsx7K2R+kgZilJj4zo+Gsgtxzwrqgoua0H5ltUqyRcwU
mIdyucuXlzn6Fl8p3669TrgcZKMwBOc6ibaY/3XmHmdcEd4TjZ8eorZbGdpBR5ra
4XyURgbsNFSZM/YTGwHML0rNMQW3uYIPB8BVIm1/JhSy0riL2Tdo7QRBztG3Hrul
7NPHbyefuOAwtXwAx/JzIKp2w00wg5O5ZWOqgJZAiuidsUcHvzqC0+pVexjxs9O4
TikUfNcOxU5RbBBLK86oZ8bfpueRZHUxszaFXEvXlqWhY0wKPIZvuYxdVn75XQPP
sjIxhs8/eTcbtvgG5e+yRHqN/z/8cbrdk0oYWDaetFFSz5912wnhw91VT8Er7VRB
SqK7shfy4zq+ZtGJF6DB6vp0m+PqvIXVnvUQ2gPUmQWhT9bGwJUbhL9Q0vQa7YTh
DpbvCnEENqXo/wK5/tZKiDKAdeQqm+b3zV2poZPJVV7fggsEZsIzXTKcGdA/YOl5
K0lCfLQBBiNr5ZhW6epyT84GIOXPDQ8Wbrbq2QOdKiF54IlsKwKdm4XWcM3lExQk
+/ebdNM6N+YVJ1OlYcAwi5XXJDYVrfv5QJqE1m6RWdW2llnSpRb4eRiu7uKoHuIL
izdHGuPO5tXEMIOb71B5M4KBuBrRMAUhtcTtFaRHKFwL/KLmlb2BwDIPuugI6P4C
46gN2RR9rQ2YS0/Lg/1IQEsRpGZ5tF7hkUDpB9dxLc8lqQKTy57HvYg9r3Go5DAF
Twsr4kZ2bOgmdD+vgV/xFCxbpC3AjU2X2d+K70rduSzW6W8HWGOe2+nkzP/eUsJQ
BZt+dHokhQTr4i4WKmE7lfK/b2mPocgubnqpfWIXdlDyl7e7QFz3nir+rKvzm0i5
6O15l+o/0Z25afD6yVWuRnCBAC7i1LwiSyXdqkfZ2sJyNWylOjx3j4I391AB7YWU
8aGh6pv8zhV4nqXyNkvtMfuK9njMu3J5JW2vTJEfrgn0mE02AdwWTCYRCrkAD1dk
AEVtDxSFpM2R4ViG5bIq0+2TX0hRuRfhWLC+WINdCEsJ1Pyan/jgP+MLDG0bipU0
NZV9gmIU+fb9cYtUk7+0+4qQ6PfmGMPKKEmriqzYyyVFgqz6Rtp90J6gJrX+SaS+
kb5ODkj5awWK7WqpIDQH+Y7va/prD8DIhVztWXMFgcmObDTNJ4qWt08ked0R6CiK
L2TFonFlYgNUw4PuSRXHxeXwHqhMq97Yi0LG921q2oTFWJQXb0Kb2QrQ0yGodSPb
nF0YUp4xjuM4C4M03s+1c5j1jpbUQvS93NUnZOeTD4N+W/aK5iVr5rOMcAn+gPTO
IxYGta9C86ZPzrszBQ/NPgv3m6Lr0DCp3CpVnmLjZ/Dld1BRB0RuUZKWgm/KFNrl
0H7y2DR4wGidKei8CexqgC/xIVAWImfB6yakeg6qxhDB/flPq+JU7405RrM2BeOe
qAY+/cEYUtWlGeQdZJYb2nxFXmn9OqdUYhtr5672nGNcbcMqNSjFKwtUViNuNOlF
uhqy/mM0nEIJ0QN9pQLKXoKPUQHbsdWQw1gt3EjMv5APi/0LIWmHsF9fMtmHRNMT
HRYJAPFsSAadpheYAhvdNbyewTlIDejkqL/mNwFqYfnVvSrTJ3rI12tenlzNTe2y
FdDzlkzcd/co0pzeNFx6Nre98EEVDd3Okq0tS6zzkk2JZQD8myCwFhHD/RkhWQG4
2NC9xOeWj/mo3fIRvetSKQJz/tmF9vcswln1synGkklfVuiAs1+xlmLkLFhwOj9x
qPesezR878Fwvo3t+0bRivfOcxWcj9c7fzrlAA4EkoIxmyBgFrgOYSSr5tAPHpiK
m2w3BcRA207E4GO3P++YZZMXdeX+FqwyRUJ6/ozGz1ldEQVDpIztASuUknTWvkb0
aIJwb4sYiZJWxQKClQNL3IerAX4desHQi6Ml3/Rb/2/BvyWbyteB2OpZI0vk9Tob
5WNChsDgOL/9/qz2QLUXc0CLzvFY6lV7MLymX7jpoxsRY26FfDLQF1SzDdTcQUm9
Q6+4Bt6JAJBkKhH7cJ2GDzXFiwqWfpIZ5PnNatyaApKGZJchSEJqcaWB+GrZ4D5d
wXBLh/ggFyZUzjEKVTx0IHuGFNetoBGKiDwoP7BGn9T5zKTepVMOML+ZWCdZXWm4
q/ANI7xhNNYAqFvqTlunpJlf3tTPjDR/m/ZktymqDLFc2hrcSeBSGxYdRnNoJtfB
vpYkv0FKEpiRTwgt9mIjh+/zWeXV3+ScCrG/Kb3tRgGqrlDsyIkr2JvEYhpiim/z
s+GQVDBfhGtl+zu2KSQlOjGRrIAv1Kc5A1AYLRh5Vqc99LafXcWb6bpegihlI4y3
ZOoh4BFfOExKEBHK1lIh5W9481DXYsR0oNnBGBjQ1vembSCDD7bCgDCOF59G0aVj
InD8s+o4Lz3LuASt+ksdlrUOTO6hneTy/4ZzTwBuUcwAyeb7yt57b9qL66q13Hr/
uOZpyHDabImeqT+bmLGJqq1M+gNpX42BHEM85Ps411o6wps/3AFV3LyE1nl0POXM
fT0l/XQ5V0xAOoOpc61QgvNEZNjQ5oKsDo5a79yH+VkKZABMUDMj3/BgyDnjcntj
HymavC2BNr3ApOVvuhd74KyfKUpdx45yqmnTG7B8y5mp1ysb5o706nVZzdbbAkAC
KV5l9BmC0c/MHb95z0in8R535lkD3buyy47623zcEhrMyo4Pfo1V2JTZQOE3p+Fk
QLxwhMegL+4yz76cl24bEYqGaE+JUhaWH6Pkj7k3xhoEYX1SZa/mrEQR0nZ/oqHt
8mT91JDW41mHG3a46LhZBR1goB/PePvNXp9+f5uQf+zRMOBvyGdFtB+67mVyGLho
5kw3/vjvvA2dHsKiloeBUgSURGEMzEe+QNK4MrW7cfMmusNKi3ifnXNTDGoinEwX
+aRXXtiKHK7+0W8w4Yxwf/zW8DNfav7FLCU8wtMY2ANEFaKyhQ/RmHWkc9i436N9
d4lguf/gpj+epVEwSfn4WwRH62830iCVzZRlCz6vlG3jgWOIgNLmSxxmPeDVfQyR
2x8Df7FGNdLUCuUqgk+W9mm48Mct3rm/D5gWwHSblf5VwgMldB8+iYFPEjLFFpD6
EagTlUTWxKfd+j2C/+dmLsLs+OmIugWga1f0ueuNCrIqz8PNpO1MLTNdvdRCY4E8
leziDO7hL81ZH+occXFFt4toie+OwGLOfLje4eNmckij6e3Ql4WBSm/LkiqLHuCo
g7VoFTAzauS4M8s4tFZM0cnjy4ieotxjDciEfzP2BX8/byfrBSdxR+4/FTUuDpoe
TjqLthmwsAJO5ZG2Zg5OR4LoanjCgXuuyavkXgv6kkZ2DW3DfJyWiIZR8A3t+tup
2257KuxvHu8yX+KJH6ySB5fC4YzSRirF82BTnrrwnAMGsa8N4QUUodLkVsOk9Ks/
iPepwCQ09VhWubh5C2MsphAA0fEH+3MSUKC7N7s7DjCcNEQc5PLBxNhCTrYq0z7+
uPC0BV8LEaw6zjrdw012ugidaNJtOrdVjQqsaUAFSKJXTmRnN9yzYSufEHKY1jhI
Uz/HooFql+mDNu92VG//K/iKv3fHBvxXNz8wBg0z6TAWKkzPD6WMrQthrno8ErYA
OmsmMf7wTa88w/AmYSyl5LcU+z/wWR6n7CqZxfFXExK/OnLYnZzaHdwBlMeUB1uy
HfbLZPwh8MXhVdx3Nu92vSDqqulaDCdT3BpYvyCfQxRgdMbympniyiHQt/k4vA3R
XPkfBQim/HWSbLihgISN7D/i0BIIJw2OiDGAdnEGh83lJisZMGy2eZyciWBaMcxA
3+3ov8P5NzBPJ/Scihd/W/YzyxJe9kRJKHx0onJ0AwCoZYzH6vLXt7M9jfdnpU90
Cc8/ymM+v1pGoUX5mjpqFTpkoBUNr1NqOHhUJCOSzY0JdMovmSjCgtt8a7N6HigS
8Nj++nxKmL1yBLSCHNXUSsvbzPca+Hf0KF/rJ8f2XoN19EfXLYSYaOM9rus1Xpxd
F5dIwUJW9QgfXy2+Hd6Y7E7SeYZqeNxa0FuQaVVrw4BYkLQJ3ITm0gr8yFGQRSeX
nyAIV0GkXryMvY9M2pNmzWCtTW1ATDVZoHQ1Q236jDAW4a2FlgJO9vkk9le34H4x
zkPxL4yyJEDgpj1otQBiZQD3oIz6BkHvl9Z0pxo55nt++ITrJuddvE8toxulCTqM
ErRHy1xosw8rjbgXXKpbjH2CmmDXAeyj0MjS39B+TMorN+hqyfuPONdKZr9T8kIT
ZOZ8BPKyv/75cT7ooZCO/kAesXwB9JX2QJXd8IFVk9B1REum3X3Pk4r2ZTq76fMz
FkZwNZqJJlXNbrXeJLNxAjPqCOQkXCOAq5w9G/YvofHMWLG2OBUMeS6NfJeW5eRK
hxcYJ1ItN3aCui8XfjspBGuEYSJ7jtAQw+grjeBZ2ssTocPglZrHVL0xzTGLAcyk
SUN1DvHIeph/ln+SLk1Ko0Zzz1QM1vPCLYDGaQTYF/y7WCdkBR9wGM4jiYLrGqPB
xbepRWSjkAKPTtPJ8RVaFUaGdxQUW9mx5v/6WMzk5pBgEmhOn7DqDMXiCy8P2oI2
1FhmM1V50vdWkMfJGEvtEGOTFVToczGf5Yn7u4+zOxR6kOZuqurSy6okoct9c/c/
E8NCBXFiWAwV/KjuOPCP5/mWyHeEll4xpEzI/aj4Yr8R4z/sJLsu3Hps6y7bs0tQ
oZAsdJwHE+Ah82BSbuuaaX9nzZj5HCA/z1b+xoNplOKwslPnZrdsOhREIx7Pb7z1
+AC5C9cHMoQqX72ods1b4tUBpnMzFodYsletpvxBX9L13g+/Vb/msEq9QrN9Pa1j
tbPmcVmu283XhZ/ai9yGUJo8az/SeeeZYLLQsEYjE5EvkEFM12lsPVGgnJUpROw0
YqeNWrLAGP7VS6hjJRWzwuqI2A0nNEX//kJ06EHmQLqUnZBIyz3yGsWnjpk/cOMO
UMplTVdHoWdBgOG4yv9WUWrULDDBKp9g2P+aykAF4s3YGbeIo8XFYjzxgpf9dNXb
OVcgFPXB6FGmG3n9cMmEdyebvXqDNCHe6bmRdeiFQiM527ZSyRsUL05+wKNL6E0Y
xQ3q1ldhSGW20yOvQECTtidijJUzx0Kug+kYEp7+KQCcOvsTpYghp6OOU/WPhEA+
SDvqs0BGSjmKJITYje1VDcgih85a6BvrxJMt1cKpJxbrGcrkWIdTmicYUttIpeOE
HxS3CI0BmgqFqJE2ROUjfLVRXG1i9qcH8D1KqRvR3G9Fg991AF9KP5uCbxN8GgQU
sIBda8JTMM6byfQVqL2PoU00rZ1qMXhcf0K3zYLxDqzGmfnWAbeddcxoFTvPzqtl
p7HJVIQWrmklqhv7GnPscujGWFLnCfsZkVYnyd13kAcpLxftnS/FkiY7oXIzPlp1
wQoWT47NnDJpNYK7ApvF6irEny5JYBnEx+54u7vVgpitT2O4TcKlW5CTBPIZDo6F
QtS9zaeKwx9Xa9ynlGjcGHnarPKwWpuQRxy2Ix5Ie31e+6qCwSQoar6GWiTtvuR3
rEBHPtZVLxhUpdwv8P8HdTw6HFSMxN7+iOsR157+9Ka9wVJHxiP/slsv+f1Srogi
at2xwPdW89fB9GQiepkaHYnoNHocNq6eNj1wp5SkopfkwPI2+bRJmfbInNVKGg1r
aLh/SzEj2lp7cJUhZdMwUiUnicO94rNJ0FANrNV/ZuJmv/ZFSdqVh2wNA271/0Le
GNcIu68aw8Iw50kz9NSSxyB3Q3e2DsQ6Tw48bGexSdEpVWCNlq0hK8rrj5m6JLmO
/QZRonEpjXJicLYksfHvHnOgJIRpLB+B6+SgrMl1s2gOoIHWKrWXtTocv2YFdzXL
9VrH0HxuGvSylHVpDYyas9oP+imlcecFKvcBOACYueBDucsHzPJ7WDXqdHZ95/8Q
zwZy6UNqNuxlwkV4fFlqn1EH2MxfdQg+PJPbNTMdrH+IOoME/7Zy3u+PuhB+Cyx9
JxyEWmbKpCYyR4CLMQEM76Iq/+6ZaSGSI9++TQWsMF2YVmOLgOa784f+95b9/TtD
8MCNiwdPQF1lHOBrB/U+il6+QKkSkCpmmVv5jEnffpgJIg85BcPwhbQgf7L8IIMe
lnihFsqfM9zBQxOAt3Lm1gRaoRsmNRjrmgmYyuirScqVsguQJU6xsZTRU5HbpYFy
A+RqHJR6wv1mBYOE7wqhFbM/8xoBa87y2Ura+wpBvBO2dZW/K7wACW2HvdadgFPm
2QNZ2zD9xEqSkLFYUwHFX65ko2zkzk/LO2C1+Gti3xa4It23xoqy10sgoUUaMCDi
3to70kI/tDVtX6YN26Ddm6SJflAguN9jPRNkSZtQFAFJ0sXyxmJG579150GDcJKi
WCzExkMfOd5DbSlCvRC6CovwOf1TWSIZbhvEtKLngOpzBYw05+ZWXnyCTCz6Y0WJ
SQkKHuS7YUCu2866oV1lO6+v/EHHVvQFoT9kKkK2vuFWGUMCsIcpTDobP/+4qua/
zclSbFEk3dn2gAK//j7fbRBgiLFnClQPv1y/ZZ5Dj5snwH2jt/az8oUEe9x9QZs9
CPaFqvJX4h/nHJAjErbblUeGXQ3Qotfu/KTC1ydb8JmgMc8dDc7C/19aUb5eIylm
nF4XE0YW+sZZ7tvxMJytyto/GEdVbGtZL7oAbFbkrsG1czJnUK+N2FmzMlEuG3jQ
gtFa2F2TpD/Lt9C6Lp+a7wTMrebQRDATB1wB0zjJ5T5MFl6oFV+AzRR3jdQxG1LJ
aMeiXmafziqBtdbtd8fcEiFWFAd+6OXAzOTK+UzVx8AiWMR/7IgMGisG+kpCepom
pk7WWA9JM3Adje+fguNWhgx9VCd3zZnl667BHLkYQgkNpQLi6o0IzuR2vQec1fko
BkjcKYf0SLkAS6Dw9bXu4N6qAU1f2RqZJFfoa/KgPTma012n9yr22lLNrhzsBss1
eacUiEOBBup0l0oF36XLRuCoY0zOBndiztAo6xtj/ctgTcGDysIGvQPBOa7v7CHd
+fqEUje+qR3VtnkGFEAbirOrBJA8f4bYkm8eolFER0xafdf2UqNRrrDx0gCdn7hE
uKU86UuIYcULXO8nU4NFHMjQFhkQqxar1NvO040d+9wFBgmQE/EgWyUE+Tpbrwia
3VCpOqX0gaOkunmg2gYVjpM+RHdBRZnwv4xJXjA2T8F/00K1iGItbLUXUY9gD5fP
vPD2S7fedFeDa5CfQXNTepIwQgaHzh2SWWCPk1Su5W4TU7UtaYJUDGSNxeBbjHlh
py3OY4fbAqfKv4HHoAeMOpzG0QCSlPZRysJ8JfltrsMVgl/SJEkQkYwSYXBOoZU/
o2GC8yN7ELwXiFchs+R100HoeE9HCzrynvVJMidpye1pQT7hiCRHBazrOen0i+1A
F8DZXGkx54mJYyqguxIsYKoP5QpUZZwIwW9vHR+gnBhFHGYNJ0FZfCCRfoUuJ/5L
Yy3Oe0Hjtnmu1CCTXOWxoOZ6vu6CVM6V6WTAEE0tDqIX7vtHQGgOVR+d4ydCEXgO
XMegMkibi5rnYCYR975+r1aXzj11XXwabONXX5JhlGa+nA1uFNCZ+jskFJLsSTGq
uiyMwCfJyNrIR1zjEH7YwAlnn2tlBAP+SvZvFh/DSYycRc7Ks5qIepofbXtXeI5v
E83Grc3AU5Z5EJ1Uy2z8h9eqrR05CWa0NaJzzRzZ16H1MrNE7ZCBxd3fqS4Kb7+A
2znybx7vHZ07efTHoq0yaT881ubq/dIdkdgBUVLfEvpQSdcdjU3EUPUqHEeBxvsD
CtQZNKg5LT+HImHj3Vno0ZCxzTu+KAtiANdv3aK8mWv4rqWlvr/OU1qXyub8MLv8
eN0lnNTCQp3hjVu9s1D6F/i4fAdwTJJkcR+Zl8uhP0VZNvWyR55SLC3OEuPjvgG3
G6VU2Ns76PFyQdEMa0Zr0sK0S8QZh4IrSU5IvKDp5zC6vWKGlejw5wn9CwjVBMfH
E3X25GIZDVZchNUx5k2uarX/QhCK9az7VS0ijLI3DnBE2jnaBqe2InAC+fhnGonJ
gMU56zOk0mYmrzqVePCEB9NFbPtosNVjE+Nl6rCCv1SmRg+vlEy8+I43h4obm7Wc
XNqMV9h71LqY2+1Dfgm/waofZKJ7Tqi6/5IO0LjnQG8H4I3xrMkxKpF5YhA7jak/
gBUeL+yI5SpibVFrxYyd+TAPGxnjteBEMtSFFgAFsrUurmDwupVwe9E3cQ6V3utB
X2HLpPhzVrmbe7WJKMANKKAGyigUtpCA1yrvJCBSyxunQ8mQyBVla8H25yPWzgWj
MjtQCcvau0qyURc6G74upY/302blqkOmQLrwTx3MifvKzhWdIxNv72CJfBRXD9RS
xtqnSiBK4cGF+VHEKvM3ochc9OIW6r+jm4HV637IOggjcV8KFFpcEEz13d9hUNq/
SiblbhiBJiGUnActCTCyUzcvRyURxejFdrsyilcS3esmvxKIHQ0QAIoBw7JXGZ3E
vvgGJs3ROn75tTK6mIgebjjDhDwJdRBIfIX5Xb8+wQ4QwtlaWVfA11URw7AHYwkq
RpbVP7I8KdC+fLR7/d6wdKAaBhSUo48K0QcIuUkXwryzNQVGqPgHkRnEHbzwmVdA
ibMPChu65CI3+RtQhNOHsvWavQ62I0FxPZlDYXDzmjyv+6RDYBuwmNLcvEoEzEtd
N/KpcxrDP3x8+DSVuhCEWwO2Ha385AkzEbTh20FpVsnW1EOado+x5Lo6iPpieBiz
mZTll1p9pK+KMkl6D+UAnaGjaH53H9pepxvX4mV5Ys3/PfGqr8pfAd2LfBlyTr0M
u3ID7/kg6LdNHvBUkIK07o7sAknLcJydPnNqZ89JdpuGVbuVnP36n8ON+WPiAcId
hryx8XmRKJSXR/DL3ZZJ0AGtdxfy/n1vCmEyqo+eF2f2ycaD2AvFI9/oo8pMNGk8
XmmMdqrqKw2zWR2YurjOyD5CXDAv6S9P7VxXSk4ZG/OG7yS1heMR1Jm0K4L9yApQ
guqldlkWfZFA8E0cdAlB0Phlrr90WAg9yo8u4c0XrreDjYBTcXhzIN92gD8sGoRk
mTKyVZVO7W4aKszlVUFyDkOQpmbiaszjL8qUglCkLsc9kCK/8Uha31oHmc9i3fi2
h3pmFaaIPDb/DzACexb4F9gXtKU967PvP5a0I34sWUN3MNHG5DdzDpmvhfPD6PaM
dSq5AQLyCmSPOOp/INpIw/iatKAPnJIifar77ZVAvWM3cEnXNV3kyX70W3AKATDU
heqqnStS1NvmAPy8WnFNsVebOXW5M8rhqimxgx2DsO+RbrD0KvWN++RPyOIFhUrg
FJk13yW0OeM+eog7I9mpomSx6pbnaLi7IzFbxW8gQFUyvXzscXpCLVhu4DUq3I8o
3KXDi1ACav9ab1/uBImY+BEOaGCYomUAJwSndpR78BjdwtW1PqUdUPi6OUFfAfTS
n1LJJPqFnBDeO08ASPeLJYYVxkcvH09I3LcBdsrrzR2nEq2naZfBUBww9xl+NOOG
9szMy3sRSJqWgqckeD4iCglV+eGKaHwyr6deCgK5jbcXFwxXG7UbICH+DmAfEwPS
Og5irvPMd5vavsq7CKWuQqvDvhIVaq6YVM64Q1tT2pgdkSwyNRsa/+tHyOdpPWaS
ACBwpZEly2CVrtPUl86exIV6W5EMU/vznnD7kkEpncuskUqo+I+6qvt3SIBZ1V0u
CJa+FFDrzg2avo/Mz+zPMPZNTrfeagG8QUuJq6hRWnpTLMY9tw+SgRb5l5HFBYB5
3S6cT/SsZbbICQrcpjQyCklxjbou2aN/xf+9mQ3960gDzERf3fH2CfxdVkOccHoy
r1mV56gVg0ESzT1bqQcZe/goMg9WuygA32fs3WK+9yuaMuD7aKSbAJHX2pW1JTSu
ufeJTR7NvWyqdIa0kAq56Q2YZS6+hBGOpR0oamWgrTXwJHhO1aHxLs4KdRllsrwO
1D6TkT/zp3NoMjY2qGQDeAc1TAfpbKxtcDA3gU5OPEz5VStEF8Ti7gq9yXSFHcaC
0lC+Qjs1vhgmTHyI/H8Ya04nypcIkv6pKX4++Nx+ZGtehzAHu9BK/9DEUe5gdeEC
PaEEnkGk4yyK+eeq3YME02HiDjJY1baMrsma3QRmTrp7NZLlNZ8ogLp2k0xc4Eu+
yW+5dELIvRwVAxU2UtEAw0VkqAP7Y093qYRKgMBuvS+Hk9n4XBmSWTxf7FwlGZHC
uPKrFKKVxS9kTDKQ79fK5yZlUlEKgbGlV7A1Ea+4Nw7Rg3mIMZ9FirZchEF3BZWp
drOismurLCtildhN5dI7S/rCjuUfHPs2aavnd0YT+dXRr+D1Npu41Sl60BS9CgfQ
6vKhPZ2jSddDoys289+d5Ey0MVpH227ti4hZbL5Fr0XPNrpTh6cGOrGsjxa4nlNi
VWIAEbXrDH6vo1ukiiOgGBGXk2UIOyWMOM0BdoqLQ37jCz3Os9RmtJFUHzUY06lP
jyc7QS4VGzGbRQ/cdObzASl40cuffstjLcGxmUecAJPHIJkJrNVyIGHwPB/7BDvn
x5vcok7kFZGeB+OTgZ8tpBkFRdyQgxznjiPXXK+7kaOMiy3grheOEbD5yIzxfNgJ
Ya82404/L0VuUntMZjXuY+a3oVQCEjmaBD96o63wVVkWZN0hZrIWvu4yVlljORev
+2A9PmlwTR7TCFSXaaYL9C8k6PbHXtAQ5q1ZnrNbxUtQ4LxhR5SOPH+hSm/DsF+h
EQh+a3+7KOAX6OJpgh2yOttOFbricm3wlljd6wELh2RfxdXljQL/d9GVTk3JJFCo
lD75FjmFBxlJhtn5TRDk6Hv5K4k1PNx2/+Fk6HKV0zneJku3afEjBjUEkGUsds4S
tkwus2CKgu2qk/K4Kb6d0NhzcM13vcB34ICn7FZz3sWEAmALt1NNbyfzTperqnT5
Izxkbhrwqh0meE9Kn43bN7iL88iuIEDu7IOASMhqeQPkbpI3jARihjpwZNDnaU83
GlwRvfjFyBrVlP44PZTDw0osrj0FEz8R/Uv1jyki6YiwKousK14l+3KSbKmnhR2a
TtujHwB0vp+ZD5Kbg3nyeBNUet+KuG9jcNuEIxq8j539M5rCxOz9+gyAgb4Svacr
8BDCrdvMBdCvM49RKaTfvxXB2A0p8G2qVKoqy06K8lJAenkvoI4IOeY4WAxLCg2K
1YojFAsBToiYIot0Z1/EjEBgptP4pkR1ftKn17aTH/VCX3GWjClmGdSIqxcqoIDC
xH4/kI/0WjpjA8SIHcwMQqrIQMDmAK4EdLgCOGFlNSOUP2XYgrH4lmmaWBlDP7az
zYn6DmNmsf6C+wkYQr3qsCd3Cmbk8XN5O13FIK+8Ds52PjLJRCY6D1UYgKWAHTnq
ryHRDtRCDbPPP+0Px5RzncK64Rlq9noo2ugxtKFc6UDs4Pgx6kXUg366lyZUBtj8
/sMp5xOYfGbhhv018dBEeNoPTcikkOSU8EyuMKvsUh16nzrZhfID4KfvFLq3uENo
dUmSwGBVAMw0boRsIlYm7hrCUMQE5nHd6XHzVE97WkXR11A6aS/NHWjyxUKx5VqC
xyousDAMbYdiDq+/SBXQ1BZq4rEgScygWF4VaEgr3O/pc3y4sB2FGI4ldq3nvCDO
3KPJAY3C/FjA9TKjk7uSsmAFyE7WBO6LWmoBkzGYMIj7JYWgbSDV3b7eiFnQlBh/
4giZME7EBHU735m7HxEx5nFCOhjeoLSIybInE1AZpw2l5pr/5TuPKWBoRqdEpUiY
pc1zWwLrJ1UuNlljrhcTcfo5YNBNccdcV8eh0+/AwFEQYHkx5S66dVtnGNpFwSTb
sgmUJAtxphFvJFiZsb6mMjN/9OTdxlD2ePVyIj8kt6YybVRoJFgd2YymLHBmL2aL
/N59nXNyTYSfJQAE7uJvywVQwKa08GuOpLiupUHbajJ275KYVQG4YRS+JLR7S5Q8
jELT+/2IDOsDZf8c/btFbj3ls1I6DBGPhdclMHds2fMVdJOkVZmmHA5oEcibcOYn
endpRAofRxhucjHL9CwJRKv5VZ/u1RasZjp2/NFc+cnl0A+CPRQb16aF8CJMT2qL
WzTMGGIRHoRLCHsmfj1BVKG9njrX7gvE5ERT1Qm2JX4bj5Fo7tm4BIXDO0xxewby
szTO4l0PiSkY/UG6t8AEiMIOPCmLT1+dK9oeq8zLVrcWGiIKJS+EXjjyrJsVO7PQ
4vRx3kmg155AT58ws6kLzE4ln5TSRsI6QBZ9KG7eAeTDP9R+jjqvxqTgfq6lJ4K2
Ia6g6zQuDcAU2wxsvZDJlEVU9QlqkksZR3vNDBcYuobH6Tpzw52D8Cj9pQfh7W66
onFZf/3oVQaI4tV8CCZoLvUya50GPq/r/d4c89TMTmsz+b0ghe9xWiXrCdQn71qA
ECZpAkkm+BWaK9gbGglpJwbYMw0MRi8PytYGCNPQeDaQgOKfJQmUV011amGlwrar
UGnCM9us9FZ7c1Drwcs2V7pXsgBWdFoAmKqHNO0pyy9HE8vhpMZiMRQXI6pLPQTM
qcjK3Q4RRywu7qN0KhvpvzEXqtGJymV+XRKZp/atJmMg/xFOsusyJ90IwK/rdWSg
JGOEp86F5n7AwoEL+DgceXh0jhdltYPtO15YWSMvc3/l/DxMfeOCHzFu9tAjXx0V
psNRycJLZErCCQ1NKo9vPXDFqLyqj7rwsrbhTt4tXM4ZLzgQ5DxAUmzUjEFperye
GQlQwLU6OUsLn65ym8iz8doguQeRzFTk/y87rVJzORFlJWkjoYi4DzK24oUvm4ds
v4fVR5Fiqc+wn0hfIxpdUAW8PZA95iQ+szy6sTpAxBuJqy12GbYCSi10hME/vzkE
kePZBI5I71qN3iU+2tNTtAXPuLsyvBrlWi+iniH6Or0G2M89ndW5atg8PL0iMugW
+aDY7o+deJyTn/xn+E3Wf6I/+8IvKZM2Z7coZyTAB98EPSO06wcwK7F7jLN2eeIC
QrVI20Lbw2DQxdpWlGNmYrP4YVg8TFWKFXzUzFQFM8JyLabj/KY2E5u/XZHdP/ao
VfNv5fBAq1sIAlNvfXg4YmYDSfnTNj7n/jruXqzW5QiUZwAaR3yZ+mOI4OI4Haqp
lvyaCRo0mwWeNTgLIDQXwhLPRyw+k+TA2Hi+/hL7Nohftr/S/BwV1RiQHvn+EmVT
LCvaEzf4kJDc4oYrPUXJPqcPKMCihAfnnHynk5bxe4VqOd+nD9RnjxbpcJl/doxp
mdF4d8rD1wt1BHJ79Iwbx8SlNpOnk27NzqBfqK3M91EP9WSH3yG92TMEx4/dZ+vi
0mBSqRCttMg5RYN1lZJsAStEpb7OglkW0mbO15QrpXh2rDVYbWZzr+bp/t/l8vu9
bKl9U4z6T2IIImV7pEiM+SxR/9d2UWKw8y8DV1I7Ws9Ls3l5B5G8Eg6cjrzF5r7G
gigLnko+gSBBaqGkmg6E963JhQlC0GqaQQNjdvubhFm3KNzCZmz3LR75z3Qk2oEZ
mVmLMSIgF/KUeOa8MyOEQUMKhPiTdxwxbPhZUMmnzwgdLLE7ZqLbsi4KbAsgqDrn
PTw892sRmnr3v1wr/tnrl9Cl84DWgB+MH36ysVYAQHARow6Hyh9LdpkmlaUIupeV
DD/jh+iQIJRE6mPV/qqf6SP38HZ7lD6U+cXarKPZzxNs6SSaHOcCFgP8dwgM61Ax
v/R7T0zm8QioTRCtkPTcdosKIUhpJUHt3/6dacQqvvE2r43l3ntAuBV+7JzHP1ZS
HEFgSmwOyFoBQpGWFBmN+ohvabUFRxKgzWCJ83K/VjjQyAUA53gThqHYpkcmoQpB
ESOjJ/22rB0QcEPatEZxRHt+HyXSjjnwqaZNBIz44Uqeogs4i5o+6fRGgJHQrUKP
2FAL1ZmEGHZSOOkmRIKn/UWRNm0ZLZ7MQE59E0pzbdqJTv39H9oqk7+bQZd6WPRQ
/IMtUFAgKnHytLGxennGsfK/l5r50hzQEmkkxwtWKN1/wrqJ8G47txo+7JsXn/Av
YfNtwRH8FS/gyzkfm3qzo/O4H8tSeQrHxtdUtag9HsDO08K+oHguJ5KkeZXdCpT2
Zj6OIWoRAn8VJaJEzT38ZFsFWFIhDmKdGTSy4lr7Etsis18apXavlg8YVmn41TEQ
S/ye9j4Z6MS37vCsS3wzxXVBuUqs+1D31Tg8Twa0/oWeCZ0fG6AshkG3H7kloCLq
VaosvQbQ2OW75/bzm98saNZtpAnumZK4oWGen6SHbi4fgX3NA4qFbTw7n1bwnM54
ylDwUhJgPDbdFfT/gunHUgzLZ36GSsonXlQ8+MtCxQKZI/Qc0c8mxrTOtbP2UuCK
r7Z2hUy53r1qR064RtJR22f+qUlb6Vug78YbDbFPfRuAtxuXsOwNOfNHbR8mq9hP
IYfJuUERnnwisoZsGA26NM4sxZSLanxtTp+tOrhaBSZ4RaLbXWZLegJv6ekDlxuj
PWvvq5P4DouqvdwWlVoLjFvl6AyCqBgw53rsvzLhYRFLr7ldniD0OeNvxhrSLZnf
mmWdfpScuRyZdy4DuaYggw0JCvSJhDTCnOlEMIzFVngk4smyj/HHFncFAPWjHtZJ
M4hIOFDCLVh8zshtwOs5okU8uiJbFJExccBiQ/Oqz0US3591Ems0+jCahO9gfmiN
UQTKb5FSz8iT678OPATuyec9C12w4qX6R6R4AH9Ur2Ws9ULxpnLKPik56p3h1hJe
QnqPv6xtQlNtsMxZhh6cy/sq/ej5sWQnRUIyJyei3ZnaZgvDNKrJWqpEIw9pKYO8
sGTOsg2K4q6JJipZhJMENj3OA64A/0ml2IcaS9MYaKhnICaI4aON9zZXIIH5kG2y
UF4gTESWKWXVVt0K6eiOUj/mtheMQuZmf+CWwifwmlJYiQFgYz0OP70lIkP80TVa
arJntRJRjVxouncHUdZiyufgRnV99GY5+IMtsul+3tELhMezXXV6q6cGLtqqfvdO
/lRpCcnH5Abp/ktBPCwrGIRBbrw1e9lPFI7jCPV8xVJTEHocG+5RUC9+6xC2u45i
ja69kTeHiOKydcsjn63Sm1gn3+xIFRUjmItAqBeNhVmFqqwB4rDO6S9icR11khA0
og9IZ3XGvWzbK7ER3KcF17s29U26jA82a9mJ57a7BybtxG6EkNxFJXcc9nRrmwyJ
qEgdclGz6Vp2Ui4fbp665l9/1a1UmK1B7FSHk0lgkIvYJ8JQba29v8zafSLCJc7c
r6daulO98InvO9w9r7yDv1OfbF1nzmhJ9wLqkK6VCIld44BXBfLHAjfkKAUZ1Q7D
lTGRk+jKSDe8uvo4vYXkaWCwKgIIh/qya7KqSe2JatmuE2BKEuO96Ud4Adr2s3Sv
++RvNzmhGDJIwI7BxeIaeNVB2k2Md/zNjEFDZi0T4iHrrE36PoM92mV/peCGTcVt
P53CUmKztmplw17KWi6NcsGXKFOBol4mNOTSa6lp3DoZyUHrPLbifqYPk/S843fa
bIJr5BHAIStqBp2tRYaMLVgr0tU59gnQED8RSATT5f7PrZ4tjsXIhJsFG+KNvPIk
43gy3N4dO5q21HsATw2cgIcfWakX1RqkOJBTNzlWTKdhUR/c94sFqodRvVbFVAQn
QCsIQQ+GjcfdV2TLGEwVGb+jbqvTldwDfE5lS+q1XCoRKgvl6hfpUgHbIIBDIC6E
byXrjJgDCWaqm6ARyTEWH+WDGMwCzMVvcm2XFr7E97mkNrolTs9d3GEzWD4dzJqZ
4y5vNBrfEkTihyymrg9gpq/+PxfZe7ToUZy/qx4NMm/jyx3t5vgOkpTeHdhR3c9E
RVWpckkUgfTfenANerme0fhMAMjPdFKg+y+Ow54oX3nTPeqIrN2Wo01Y5d5tQfQ+
yL+KVlUXqv2Mc0h8eyWYX3TSKEnEl71Bg9opkOmjl4B/KlQCY0x6p8WM9SxrIEBA
TVCL5aDoW/b5N5r46PIIDQWdChSiCtip583dimsjadZYUP1vxdll9uyVI6m/9tCB
irJ4DeI7XHXRoyTIoNwSENYV4HwCDKsmXvTbpjot1z4zVrKDwU20FkGcs3PLmwzh
3/OWRErGtXSRsZhlwagUYHmT74rh/1WXXly/KEOP9AeekmnDBDGiFxX9Fyx5BF97
jG+sTUuKdboGS3SYF/Of7aKt76e6IzfUxmxt5NVp86CkwhXYU8rcj8WkCnhwQWoy
reOlSDz2wKC2A9JpN0tKOyhUVYeo5LVd5XEdVrlTv08bi2y23s7u11DSfWqQzHSR
bAX0KeHhX910HlGWHxYHN7xhhpmugoSHOxz82+dPJFkqd+QJVMY8eRrihLsBDjjb
Q2Y83jQTgez0wGLInFYqqYCKS7t0J68ELaWobDqvFikSDBuJHhRI92W26k9BADFp
MYJDzBp8ovlJwh0kz7XNqymxb3AXuin1qAeFzQc8fwxLvBxvK17bzPjqe7Y+hC2B
BbSghG8gMPIoNxvTNI+7T5AY66k3Fmj7rgtJJ1mNOroH6QIsDRX/wD+3MbQAfORt
A71YsezTcnTWxKuuB8XfHcUgTlbbmR9qTQIZWbJBr/TYq9lkYOSL/SL+wpAoIxru
RkdejvHGKCTy4GXDJmnafDNsK2E8JpMSgMBxCkIHrdgwGudSZHpg8712IaeAnW0j
uazuapT5LTBTQJL5U8U+TXyFBu18Rjaw3LOxWfjRIOoPR41u++y/1w1U4g+Y76Yj
yoK56BNdnOe08LDuCw8pulNXQciMcVwPcGESoZdpYk2UIj8IlAS/mqIfqqxyTdFk
TNG5JiVY1yaDKs7JnmNMjNpU5AIamMcRNdTwFlE4qToSj8eDgKDWvtVfJ0IdlF1t
RW1DbCWi2j0k4jnv3nnBS0987TgOt838gS/OHBYANsDmnKmZi0KJ9xqRnopoEi9a
tNvyVjYGM1RbGlITJd2H5eF1PPI4vMjarcy/zY6P3h3TaUjaqP/4Kowkaph990WC
Q9ZmiWLmJTBb8btvlbjA3Pb3th81mSiOLR6Xvxsqodl+O4CAVKmK1h2zvs3ML/Xu
xvYO1X650uaMmioIuymPkphScHs4LlniLFKQPGfQQRdQqEwD0Xb6DfPiDkN9CVHj
sUBiY3znXrQuqqnhUHy/RIOQdxwTeQjtGCfVYrMMHGVcif7xm1w4Nl/XnXb3xJrc
nxUy2KeBqSQ/cIK1lVkDq/RY3ZQjeV84radeJVnn4nbph5rfKPKkn3Fu0nhJ4Uv1
zwtjX88Rd3UlfgsCbBroFUbhLICorBnNV2g+IMbov0yNgqHgSFD01I+C2GOwJJL6
WpK71GHFHQB5z2/+NoZXe4lIotNFlJEPKcRG9nXhWy2D9u4szUDSyBwdDi6Xi6L+
27QBAqn57uVcTFD55mcUtQN4Px1t58DeqwH9Ed6fdvqEOQH0n+iPmLZE56QCmhH6
iHkw8Q8Adf7jrsx9OlV8Vt5WBHk/3h2j2jxSX+o2j3NTKafwq8dUvbykEHV7sY2z
5PNAYEI/9qRamjtLVpvvCD5rRtjudcb2HlofhOuh7iTw28a5gGXotv0Q1J351/Nw
qdoYih56VNrkh2l4CKKEpM9An8DdlngShjJ5eeb81RxRpc/Uox2v9nHeQCTFzg5b
Jxa3Ad2sLTR039S9vZQBPEzZe5FS5GBIwy3NqKAEuVji5ZLPWbWmuBHyDFKXIrJD
r2a/kHQWMonb5JFhZXzaw5nCbhN/DSh7luKCA3BIG6GG/PM2FdJ6AiRXmFfo3j5T
E0IljLrZfaX1J09kJ4JuNnO4vXDXO7k1T3E/7uG1BdPwonqIuVW767vEte73rx9t
hsNwmdWFGq+cBQ/M9qFW2NltGmhhISLNIAfdN0hF82SFw8yxc4+FZW0EcgL0DOKo
Ys87XwHWTO6auJCrrmdttazZlaLwkojEpbUqVpH6L79x0mPJtnhcmbjYGg1fMg0f
bc3NfaKBo0oRX1MSZmfWyLZiZu2Jbv1VZMub7v1ugAIs4h0rXKL+Iq57hD2MeEJM
HHYMlGoX/Mv9bB3QFuVHuGYfhsnx0KgKUxLqmzLLGnVFHzWfToaIUooc/pg99tCK
FqkkRB18CQ3gVO7FkHDE59c9wZnBRwyke3STk3BXSU5du7gwD2vKVx96hAJ8Ak9Y
9LiIRi/z52u9e+MhHa2TP49oe3fGyNc7nLfs7tUc6HKrXmITlJEqXuAWhPoK86eZ
LcaHs45yBIkAaRksFobL8a1ZR3FrcUJ4zQL3oP4svyG9wHJW1cQMTPl9qs8Fav3K
tFv4Yji6Wr5DvzMLFLR+9en9wxrPMW1CrLw32nj9SW7AhurYMP5NMInQbjyY4j2/
81Eisyjd9leuJnYWxcMnYGHqZTMjaRRvfkLYLRAaG6aEwNZoUmuzhINU9gPD3MPs
CbZPmamRRcj1hyiwkQnes5KWdvTEw6QRT296CXk1CJfWpX9DYiNa28gOqyGfm47K
PIcHHQXhJlSqZTEJUNEgraalJhggC3YNfbDihoRVj9GUU1K+uR9CkdACpHLX+KZ5
y/fkGwZOjVnpVktkI4PEuiK1Bw5p6kAhqx9gmI1OH+l4Ap1ktZojadTHw7XOpYaK
zf9Zr9S9ByeHeg7wqMjteRDWx2DHWEuUdvnNfoZTZcJvOZtvVTGX4NzcnHytasWL
O8dqvhDYv0c4GnOW9OFwiTbvz9S7suRs9vEvejaNEYzvlNhqpBND4FRelpgSISc9
J0ZmuchfTy9T8h5Zd45WnSxDBPlXYiSmdBH0zM1xVYO7kR0Qark8RDnj1tFN1rYY
ggwL4BcQOPZusGWvdWnewZQw10q5LMkLUGlWXmgLiifPDjVJ2h32Z4HWpH0iWDFR
25aC5zPtwykIHNw1iQwBn8AQpIH/o/LRnlWuinbUYggVJzvTRABNUNRUyM2b3qdo
Uij4Mro8nBPttxxdZ7wMAAB7mssh/flKn7QmF6Jx4g2Ld5CcXmH9QlFbuNvcmHY3
DIsz9vQN3Z9wybgsdWD0sl8tzx+kH2pZbypDf2oQiiZSf5CiBNDYCX007g6s/dHV
C0ZSNnQE2n171cQY48Yow4trjNn21l4Oa/vIjaSAY83ZhLUIhy11TeJfn7DwY0j6
I6wcyDj+m9HFyTBl4rJm2Hd3sv/y0eKxSpRpF257qgjOWt951OfUK2Pjk21vg1G7
4gm1FulOS9bqvOtkKZrBmhxsf0qgkwFdWRKtyDISY+21QZhR04KbgLP2MfOn1kNF
y8uEuZvtXUy2G9UVRkroxXabPtG8Bz21b7tp+KnwfA2UfqkKS2Lv6mH+CmjPWkBO
l5j3FJr+uH6ajgfEutDfVtie7khw8TcVgj5f4gHTSrSTRuiGsRhH+sd4HWHogfJW
zoiN15g6nquPeRg3y03qLNhQ7ciNoWVy5+ldv9ym+eoulHN+fs5DRFqkwfOrbi4n
NP4Xx0OEoNGD8W75C3AzVGGX6I0W0HnGINo0t7q5E4fW2J3FKqp5zVh4ZLb69ZVw
xWWNsUrqs2p0b1lfh1bC39+63GIFzmOq5S/wEsXrDNhM6QXhEkh5xLPgN7XMs7dX
f3zQcjvyB4VpsJflEXwWJ1WmYoNDuB6Eej/S/1U8o7GMFv6hDIaLEipGKwEyk2O4
+nBmg4OzNVJQcqPg5wB3IdA6Aw7ia6wwFJ+WfNdZyfmcdxGMuiVcFWUPTOPgak7P
jpLJzVedjOYkcaUrtZHI7N+cxj50oMvhfalJfdM+5lTnjMHoza6MDSA+IwInTSul
UNNCbepaHbyBvoJSdQ++6lGxUFu+8jclmuUVz8BR07lcauT48FjopB+xnXb/ATqB
pW1HxqBDhBtzC4LNPHiINelS6Q1ZOGc8LSasI7ZVKBH52V90KzTVY1hWG9WDoBe8
FJnGgF0ZcPNJ+5iqqI2RVLKFkZVFPxhzxWbT2xneJmF8Z2LhNUZVSWqUvTDmDlu5
Y0n0D65LtiL8MWHMV7g6HSpQ6RwkObF3c68tKfDYGooWY7iEawijhjkbO+kEn0+w
6QTRwcVB4F006jItkmmceXlU2gvNBLco6D2x+RkisrvUAt+ZZUrWiNDx5eGr99Cb
s2csdStTvci2IZ19dYGs3WiKYFfBpBYq4LASAY5H7r67Itv+0CMOve3sx9gzDIkm
fP7a2NWjk93UY7/+A1ff/S+BeXl6AG7sYZVnCYLehYrWNQNhzkEtrR9JDGLuJACJ
tSytS6ctqZWXlZ3wawGqRaPMZBog5Y/9uLCPDaGThu3lHt/6ibQsl4DVRB2/Ff89
UcUhefQMJ1HhBWP6eQP6RQwyn5a5tDLgD5l3Zr0vNQbhXG3wRGifb4ev/Su5E6MN
YCeZy92G2m2pM8LXqaCq0LG2F7gRu3OdOckMe1uiIu8/EPR4D8vTTKh953Poqaqp
8PG+exodgFISBCAKeRQcOmMSh7YNqwQldxh/sbnzSxEIoE6kD5nivy27MeFGStDJ
lFokMo+3Ui7LzbK8lNcDCDLpwAPJ267og22tO4/l803aW8dSDCVaL0dyETwSjPwz
5BEsv7Xcn7S9HHvGkQr7ZKRG/18Pn9QZp+8lTBTFQ2M5G+Hu2U0jQwUSTRcTxoqc
c65lyual/3teZzcAYctah/iUM76+UKOWdDipHSt2OozQ0Q5cvBZAgmo3Wtv1Psom
Ovnv30hGMGPlJMGbPTi1PwRbNWzZXzGeC3bGcG0uZhjXgRFXvMT1yzhQhVVEDhpc
CCcd94KcPHa7+x3yHf8dBd6EPP+4Gyv+7yILSD8PqcJRzJ9XCePrddaTf1tpaO2M
ODHOUyF5cSu4DFcSHsTqGnoeBHoJVtFOHR9jjPPEcnX/ncSSXKoh4nS+HpuTmpCa
aMeeSmGdzz7DDF4Ycja9PL2FwhA6fc3O0V7gufmymWjsczf35+YW6A4PLaXffyN0
fkqDK6TTGnJt+TvfNuOq3CYuQxtfGSTX13FMRyIhdOD/S12YtBKWnvZUtwuGZsB1
73jSCKAUuXG0kltBhki/mZcn8fEwLswUGz0i2zii5mjYfPCQgkJZ0a6AzeXkycwO
l7TOaVC4IDBc8d+By93qQpceVfUyGdiQx3yZT+ZAdEFxHsE+8QwbfH4rQ1DbKHoe
nhOuDi5xq2ceIG3BN7H3s1ZDpNW6eKiYSfzI8hZZktqQra86YM3Zof0gAezUPzFe
Fw7NPNyl01CNvuBbM7oM4Ap1n+LlhF0KOhsU4Len2WWngguAQTqRyS+Bzp5rqRcI
74GJS4DcUCWYRdRYOrROJmoFYKB2Mb50oogwmv3wWRo3lnyQWaNKADqNaRr4DSG3
rqAFHHkxEZ6ajsKwA47eGRqWnR9dAFa2/kGEkjEMkAbCvKqd59XISw8reYDmzU1/
NA2G469KEn/RS8sXsAyLeFC4yKusHUOoWVxpEHRFEMUL6ZcmloBdsciu39YiDVYN
2RZOObZrHt5Ii26IZpUOHUj3zdgY/uaeuGYeal+aCsUyviBU94joqJK3u00KlPy0
IFxoqsmsv22wl4ZB6hNjYJSM/eh9g24yMdU91Ul93EHxHWjxyWUzJpM8RVIFur9w
fJU1qxoaHUClKQrYjMH8M7WhBDn7G8vdewnjkD9EhRXz7p6rBdCqSp4mOhxmp2iq
tVxiTJIvLBu9xnGPZE4apwc18S8sRcVOmL9ChVhM7t3opzc8zx2/YcK+b3JxdJP7
3S1fYvc9rpJFTfeEVbGnOMb+gzKgeDP6l6WotBUfeatWNUUiKXXdSS7gdwjlzAAk
NqK6Inh94re+7xnFxEcoWT11ijh5tx0EBTqOL8KpMfPYxXAOvbOfxF1AZWIpVx2K
cFJuKLwSV2y+0oKxgTKOkDD7JdWPuL13ZNqDVaeUDjQ/S5BVfl0PRhMUwthWVCKE
255AA5n97U+9f9AUH0GJlxf4rSetK/amOajVraGf9Tnu/ogsgdBu+Qv4XJOB0O6T
K+8XfVbyzdks7eRPJQN04hHz+WYG1ncl/b0uKii6sE+wSBE7C0bhoD48tZ31DukT
0bajwIRAlKrnDM2maXG78G0OaPD0v18hCXe10qVFgOjzzsIj/eNPZhpImtfVremc
9+vqdmXDNQYV9L9J4cBwip0swWLOZStdQ+K7ctCGz8/hjOXL7LjGT8TDsMZsVuKM
aMytmOxXPl6CXcMgr7kvxZDR2TS7vTEM9gXoTHU8OiwjIFRYNfq6u1s5UBoNbs6c
/5gvdIGHpiaX4PqqeaP2pXAYebzakYfEPDdSTtt1ZgRYJSxdj6NIvlCk0azcUuoH
lykzBcQy3yEy/nlRg+6bOb2ipEYn7ViMoXcX24IjEA4On6TJnwWYDx6jT5Zo18yj
l1ouNsZMU8QgMznNhQhE1Ys/5mKndre4B1SBqxszTYqjSVWtGK2ZADDgivBqc4zZ
+1+gtqCepV9vhqOBbNanKQUCQkuD9lsmiUE+uVBXnOIiyP9+WQNVYTXwIofoEyYX
oniFzfg31tc18mJu5tXeHZtWJ6Vr6YXzBvRClKsptUovTpZ63SlX1Y962vfUkLM9
bioAxifcMPGXA31qtfvAevh89aLjbH8pxh4gylOkJnNUYdxJdsUK7z6k2E2icVRD
ohxRCYwg0BuRG7CYCw1xbrCgHvESTkA4c8CoWVsKTQ6aSLQdFY4idPhBrkCb07o0
bIPa7ET+FwdL3exVBjoy2d7Wq3D1CqmfjAycbckLL65T+XV/BARgB2oSyKv911nf
PEEc8bCEI+iPbgzKtgjSqubPstv1IvaLLyhQAVqReYOnP3Ykdx9h7QXbqvPnD9uu
CEJtL53pF+doHjkasSIneYKhojGHpEEMl9PUH+uhak3orHwbwr39WVTCWBr2POOs
lKt7oEMm0rMXinvdgtJiKd62cC/kQrKjiyjTMC0EVylNzFlOnJVcxQ7SOym9lAp2
ta4vUZ6kZClYP1uLPvggef+YMvbn58Tk26WKYwvHH/W8a6Q2oLkRDaP+htfAxaYX
LzuN6H/6koQkU0HIF5vXDOUN4bf0sSlE+HQvwiHMi3OFbXfCiiehA1KlLEPtYwe2
UyhRbZ8U2u0dyKsF+Wh+Mu3mLst1aHRR8SJOzxQ7wy2L5HrRC05g3SrJueqHjxRo
nt/68upWtF6yGzBzv3qaSLYLmIrNrrvLi5Y6xOk5Xs3RZJpbxGdsG9sujOxsfhhO
rIn7Imf2uZ+ZlbZGzJeTVYir5Dz4H6FD7eEWemPvC2a9TotLPv+We3z+PTi+3DuF
kmrT90ns68VcvHFsmKgmvgj9No3zAWve4OcDQHu5QAluDnYSY6w/mpa07QU26GdP
L/tzSpFrARMo1HLsXMs3R5tPifkZ+eNY7xQPc7MguyugdhiUQII89dlceZM3JtKD
NXHnK/GKXzvxn6YQhZ5/AjcqyHpbe3qToC2woVvwuCfA/uI3CFUtt1NEgar2CrRN
R1GNQjXpAiYwfWZYjDggC4BrA3pLLDwJhLJpnROo10YAK9HtwjQGzP8suJh22NkU
DPX/gC346lYb2/SlBTYPpjH1UFXNbMEC9s5Yd1/5lxlsArE1GCHJ+DrFsYwKbLO1
DBUNCtBr012cH1jlc28yRAvSAbppFJXAI5Q3MhxyEX3RmdiN7fEtOBVAnjexgzOv
G2k9TFuVjF8BkXqUwQscplmPasQGoP4+/AlpumZLTsZEqch3zGuF93MpntYNZi1+
RwE28A6kuTcYSql8XkV4fYXe0vjR1+Hj3ATiHjLmD5vnNlTWt85bm9wHqG2uAhXW
mf8Z/BefTGBPm6QheP6cMEShtlVKXP9r6azoFTceNEiAQrcCwqdaCjDGhiIj30Wu
c9216eb4GpW8Th47CTtjuHTuxBH4fbycezPA9JUnG89NpJM913R8bcUhYFKHPhRP
8ktOeMRVTcirGeciWHgnh5lMS6sFWhvXYYmyXdthzsqlVm+s2ztIfIS26pY/hkWR
XYcDVtQgZvgf4TS29pPh9cFVxCvagcpf3rMsd7LZE3YZn1HmxnOEqqsxqp4IcVfB
ik4GNxsEBwyPGSI3+T/85LstPyrLBKs7hVTEF5OQq8I9Fukhs1EwWjpEpFpsYyJi
LMj0vhbV5ufhuGRZin1ZwAO/1KWXvJvYanG7JjCFS/kBZsju6+o0IpHLVJzpG6Dh
y9Aiownei6AFwCjRyGBSczpjRWA59gVsWtJOebeJLoQYCJpCpPMKWZtgaXql+Eus
qTKODTedEwvcNhGTkczbnCV3SYFGznqf5JDkb4pYLAr6DrvflQOd4pdE1dAa/DWt
4hYL3C6GUscEua2GHCc5dCVFyIsNXkCjAz8lnu+6reTTSJjGQYEspHllb9Ogaqzh
zG0zK1SxGNP+RP5seu0BBNUPoVHf/N3H4xuuyg3xqiTNnkA0jFnLNk0QS1AdgWgD
/7CauV/Bk2m1IZJO0CaxmMxsLVZhSPGN0IvRLGd1Qef3a3QjSNTJJ+mFRUtPBKmn
N6bbmWvUJt/qSWyA+HYecA7cdWWoLDNFbHZn4jIOlmACZRQLFfY98DFRpEpP7vaR
q2uOQnciTc4OVqdiiNeHR3qTTOKo8wmArc6SqDIS6bXE1HUbhPYzZlowmnU2v75I
daf/OljBBXm7gbd6FGZwzZDKvc1uF050B+vM59YoKITFvZXdfPVzdAEIezQaOs4G
5vSYtoJN3D7pqc8q61q0/zGRZb8Duu74SGt5eSev/vVa9CB2DTO0BFZRlerMSxp/
Pip+8x677wtxuiwZQkWC29DA9+hDcEQZkFEvCInqF7gCfNaJwkrvM7VOSL8FzO9L
Wvsafv26Uiq+ErH2HDZ+tnZmQL0Vm+DdPw7y39hCI84NgSbiRuD1lTU7SpYXMZGL
ia9jDRWiHdM1pb19Xjnb9GyXeSF/CKyut/BrhE6B5SHKKGyClbUnlL3QEjkcTH3S
NHBnoDjbInKQJGNQlEkOcQkjbdZSYL/MS+V1DSxkt+0nWsikskmhj8dXc1tVxIgG
1jS01B+liR9tWSIbnVmSmEC/pwKj47pwWIRmZ1Hc7Dhu9ZOEWBORVqgZzIVIdyVQ
pGTRLvQBATWe0xW4/vXVPCpJH5swlY4bHTxGpQDEOWcCYZufeW93aKe38p7EDYPr
8D64vRx7KDLgJhOTHO2dbu/KHOuGtzbsQ+BjQS4b21+gaeDwsk2EEorO64bO02kV
iTdIFVmqkcp1ZF4ZZNVtJl7pVso/VNHtSRuVdKeLKJpWBEE9VD437aiLjjFSFIU1
1c7+B6czW/5zCb1yHrBY5S/33hM0sAE4H0a0QwsBon+DbS1D3newlrDYSBkw1VLE
n1QJQngCthYFafHqK3CY1vwVlgi86R9+wggBqpCxnxcduYGJONRJLK180uWv8CHd
B+AxD78Fx7yPNiSocbOq5x43B/qf/gvQ+awgcNFfU/fMjI6wVPUbjsFyImxlwNpt
7/ps7PSVVLIAFEFaU7MYyv9oKOWMQTMJlN2GDOpuuk6mejbapckZmj6PcfcG2NqW
njAzHYyN+fdxSQmNcegnZoc6p3iqEd9c5jMFcMIOq6Eab6gw6+EpAtQHW9vpyZRN
NofRLrBJy4mHViCV37rQekDiH6/g33uSdrYAPV+NfVM8gfgb8NOgmIwDZe2rvxNc
xQgX2b16b6wIxiZOyrDOneHsZtMvTcyzfuY6rUd5jSQjVSWoN2I7qcdWNusFKiAI
k7HfgwVMAPaFMKzmX5DWBI9q8UIgyLHEUdhLTgwPLRtO+RuUY1HPzqS7GL7yNZnL
8iGCDAhDWNuDDWB2+efOG0YSEmv1+EqlyikSzkA4X7AX68nul9J7xx75Ac+0GlB4
RH2v4gIXKK/BGcj85rpC6syfoLdWcFgmkg3jsvARndmSWJNrkoIhxyaLGSOJYqPU
h3hA/rlDo/VKaJN0hz+LX8Ogp/UTXUPXzlSL5rbsegeTH9v3dIsZo3iv3nijwazk
MFJjWNtEEU0djcXUgLY8vvlo3IH7ANMM1F/Ax+ZTA0+eSBJ+E12bMhjN++LUlfzm
x+SGr1ArguLAVE10yPAxSAa8OwCMkHboi0oi1waUMq7aYyLVmeZXdX3ZlDZ/Uzw+
Ly9ZMZzXSvwSA9og/kenWBS7pVlXEeMtsmxfGwlNYxH0GExpAcvqRlkw6l2zDg8D
yMS5uGyIpiRxai1wM/ACZ4GrHg2chQ91bpJzBUT/OTq/cjLZClPx59W2Kv9NS0Sl
t+aYyQfg1Y7lM0ZSf4EbLnYblBRG80815LtO+O2uztub8m+zss7FlXDpVVFtwDU/
GAlAPydHsIZhUPbkqCg0KeZ7LgCwDSiuPFG6FFmgNW369O/ETBkRB/UjoLfG5oW5
e69dIDQTLGcBE9RwBoyiMWlrYnFWd9ntiOIutlSp6Ft4+8an6s8ywjpb3K1vk9A7
NdSsajdEvmm5SOw5ADsUo9FhupgirZ5tHLkzFBSFg6civX2SevkQKwTJhaCkXuBZ
PcafA20kfudcRXhB0073ErFq2Y4vDH32In8SwST9OxPiV3Y3739U5xr6iI9dcHFI
kEsGUP8/ZmiUGDMaNrvYqefjTH3rhQP9QN80qw+OP6FhYK/kdj7wbl8VIXAtSrxi
A29PSecfp28GKi/PaKUD59dwjTTlhfa/elBZXiHUCYLSCQ5OeROjfIZO78MMyVv6
yQuI630zJwMQvUsRlQdn9kxUorS5rKr7ncJ3pmUXm9zGrIUo/NbzPChGggdyHo5n
Brm2lLfAkwbFxw1dqLZ4JLD+dLmayv9Nfr7MwK7Ff+GA5q6nQp5QCkfcsNXVuHNu
SCcWFvKLL42sfTf9fy+bkFKcAItwJ6gv8AcMNq0ltrUtoB3iBQvWdwhBXwM3180m
MnrAoZkVmqFUTCOB2NBNTsGevG3+6STV1XjOh+1TG6pHW1V18uPCam7hvXcpz9r0
ZwbBIfUsB9AX2duvH0UcaHNpR315Yr7Yak+Ot5bado1+MwI6exvgee42MMhiT5V/
MroN+Sv+ObEAIgG1iM62LSsBlgw36KeQ3FiXKCrRZM1s5wPYL4P01HujRJUJbco5
Xwim23z3MYBEhXG/fz4H3/aC/ewEUeLy5qjzX7Uwf1W5iIcTJ9qf5eJ87OQR7w0A
sxQ+2exqPaNnHakktwHgMTIJME4Ow+MQYEBTgszMH15KZJjgvKnwUZv+F+2oPYTW
d5iDvl5IrZSQCNQ9go+Vxt7nbqIY7WT2tdEJmY4nbQ0/JXLdSFxEH4Tu4xoDN622
bGKM7pn872YzTUmz2WTAaV8eddyhg0ay4WS1Ca4CV6bjknggqakdiT64MCH+EHTk
sKD+W6IomSuOy2Q/FLRaw93+ySgdGGJtw7qfb00o3027vxzv9oGJetUew21bdejP
FWMF0qFmymuHU2vCEW9WZ/lmvv+V3fGENIg5lA00HtxfqMAWBAmdqVlk7kPoxEgf
IQsUjkSw23rl6C738jpXG0Ua9LsCewp2pzpd2ffU+W1O62bnZuHrmgHAYB6cpfLj
Klqk7TVvhjdciQ7okLD19WNJP7OTTybOjtbzXZeQR485sArGtO1Ch9AjuJTK4bhe
YDJQnxjGuIKdtzKa27x4zS2QLUCcArGEbl+GEI5OQrSzgBzp6Y9gxCMeeyw1pvIu
kzrAFMmd03S2wf8KhwoyBi1sF8aC/5Ld8rvdZqHyweKzltmRW593jSgQT01Nthz3
jMc4/G0PeHuR8W591pMnEAtt+Ez093Dpd1SZkCGgsItQVJHze9M4fmgd3sCSBeZm
c1GAug6JDMi8aIDz91+LXdBK466i6Nu07kQ/k6TdVnKsB7GJGJWzaa54bztmzCN1
egK6mbjsooxKl/eEgWq5+9qxSctDjXItUXTb2fxpt1UhVBoPdUaSTyBFGowNyfsB
iYBdE9JvkStzxCE9fnQLSLX5Cun+HcpIF4ELm9vkmY+y7+q4QZvG1dNEDP8iwIJr
qdnwmhOs7HYwefgn7bxMvld9uiALaNL6OjEb7w6/SVf/nPRPtHAC3Y7kRVhIm/jX
D2R6VTWYh1ip42DNOuNXqzWnkvwDDk1bmoYQLKstLePLusjBgTbaqy0SFpCFAAQK
qCQllDhC/kTGFQihcaHQgZfUiHPYrEb4OVhqhFA2+AsPBagus0ty80NTT+M4ZfQG
CSzUj8rJdTy/chEqx+N9MyPO7butCe6f1jOZLQ4FuJ5894k8PUdZimhnJcB2wMMi
VDUmCJ6pRhr4oSG1nRfG/LdUWx/bRzsTByhGxN82TqnV3aCxSxytjAtUCyUZ6eJh
ksixi1WT/jJFrQc2sGZnZzQvGMapjKhySRNjnCBaN+wIlT5vQPTC9sSRM+pe343d
b3Gm1Muyw5mjmGY+2nbZT2IOXIuR/5+t42dGHXOC3+vAt31N5TnrLUpm0X8C3nQK
2NO4YKhYA6z5HEm2e3nmkZ2E57vx0jH+YDwN0QYNpQYAKveun1QvQ6wJm09bADgS
YC+B5Jf4/03TRMAV9PEwvQ5+6+7bd+FPm9eXXBJNiNOvVofVY85sIVJ8HU+TahYD
k8lfSFSTvjD5kfR6v+mqjMo8Rs9Eu/QM3EE6jBJ6MqWjDtUQr7671+zhkY65jUsK
aM0DLdYja4BnkM5tfAwp1mnv0pbfDwha1hA3E+bBLPLpXqKf/PviBi8Aae29SfOx
vYD/SRiJLamG/g6JwmeFQOXzs807AHu0fL5GDvO/9tzxMH04sXDiFEKrTVrGuMt9
9a32qirf9PABuXceInvrCl3s+2NrSu94QUoJAkmAib6dfNmWmN9ygEccb9irH832
q1SsnJTt1jABHAHuKZYfMsM7s0nhF9GHriI3g/a+Qjqeg62s0RaH1416/i+NUbDi
iXPwAvBgHMf9pEroqNRjjMOz2jzqiNgVNTlFuDssd+9e04MFMjlvn/ZJBLWPKcMv
PbQ3l61GRa77CPXQ+H6TF7xqyNg9bfCu1ETGJl3hxPco4BywbuN2F2hsQDnNfbZ/
tuy4gAlOiBid+qg5fPNssoXiPnd9yZ6xeTumXGY13v5HtokIw72KLHtcRM1KuCJe
JAB+Soh6tCjPfk8QjgUYqIt8ZL0AVVZYb6xPd7ZyRR83duufa0HlBqG5J1KCo8sg
+SxEh0WZ5rEAMKCtkprRcAZAVvtjcUGmKkgSMnb9jYx2Fx8pXBV7yzO8fmLcC+x0
XDMYJJ6Cn6E0irIomJCMF2DZtow710dSvlLg7Jz07ZfviGmk6xluj/bXmgbzVY4j
9NnRQW0vKgdlbWumzQ8iPFgBSUGDkLfqonlCTqwH+0sjfubkdOidCp9YE/BO3KK9
e/CbVWQbz5J1HG3+PYSvs01rgpI4SiPy/miphCGcJo0WZ8ijZ/48qo81mw8Oz9fS
Ue9cP9HOhSXzseY2D/YieIyrEbIqvUcDsmZTbzDvnhRaYGwSSsmPkQtVA6TUjysT
TEdN8JWetSWwZuxgIBhINLwQkFmNFlignjOyNqKTqIIA82ai+42jDkChLf/ChcP3
hjmfqj/vN/YQbM4dssMsfuuQg7/6T+ooaU6eGKMoRR6x+ZVLFV+bfR2/bBH/4uaK
6NHGZYlXFOnyQ4FWuUpyq74My1+TX3dAu4Ex6QuWyGuJlrLfdR0FcsIBlufU22Ia
qtq23ugK9/nB4/mtqmAnwsLmF1TMX6ydSpKT9lOMIcl+T6Sr3dALP3GgdlrjDyOD
/yfPYchtPI8nWlhoNpBIG3Q/8nmphpYeSDy0bcgzGMIFSHSac9Jz2WxZK7ruc/u1
SxkDtExW4OAKiQG+4lXHRgodpb/ipkdAp7xtFENq7572Brd93FASXzVWVvpKouUc
Nf2MtdWxzFtSW5Z1ru7McbFi20Z57hwXHVR94brDn3S8tExuyMHEn25UIfnirmh/
MEgw9jqQXtJJo65i0s97S1E8aw8kYu+6WS5cTUE+r+6C2k86GjUDab4cg5DoaH+o
fFa/UU96oQtcsCNO5nj5ZrS5tek8ukxltxHTSImOq6lhCEWg+lXgxT5IHG7BzdnZ
HuxXTImidAJW9v4wtJQ3EZH6Y6aaoJC+z3J4jZiGlCe3ZI9lBvFKhBBHGJ7BDDAl
HBgOtXeKQbtZKXr/4sGrgtBOPCjfOznH56sASVQIsxRoSZrqDM4thIsZZhzNyOEi
+pq1+lNrr8rDxSnb4gbo1MVmkfsv6Is+xKaz+L0cQqees/Wns5s5deQClW7WGUUW
ep8MBAcHXvhDtog0tzeM6nOzNpTd7qPscwsY9r6A4ShqDe0M5LyaDBuCcQarSyNU
XieIg6dgwhtKMOMDwKsJfucn9P4A0kyGr0XsjXOsihV03JR4gHYTFmaHPJHQ1Cnm
/dBtvSjEDpDFwG7UGNKmwkOLPRL6XGOyQkD+gwEu55qNdYIcvS0YHSXdQqI8O5yN
xUsqrKuV7TaXEsqpPhAUbvzbau4UmEvwV3U2lGrBv6KnAUPUcSFqAX1+x+4LOJfG
ne+RKf+ChgPDRy/yjAJrg+HTpW1vlmjpbZgUlFNj6wYjW2lWez6Q1JNcFiDJUKVT
tS+N8Vj5k6lR72V4NKAzVBDHF8+NbAZTFKCh1oNAZq+PyBJZ8pM52IM5m9l9qLyS
kqCtOPClCHC+fENxho/9p0ga2IBOwDr8/9tg3WyGJK3Zgt5Q6yge1JwT77K6j+Qg
7hVIyk8UHqbnL0UOFKAA76a9KkL+QPgMpcxaUt0GbrarjQRoE4HXpFhTDEmNHRlE
nhDesyNrGPVhgXoxRqD6OJkXqOdHKrP64RVTS4nMwloBIdMlOkuohpcKSftQwlmv
tZIJWDtICNxe5vmE8p6YXfwEfjPmbsOPAkFgCfYj8I5+N0xxgoGl7Cq/bzxV8Mzr
JSYJ/nAoOPKymJ8E87RRbXrfO2bJ+OzkIoxq+Zc7fyKrPIFA6cJDYUq84dDsqpGE
i6+zTwzzzy22fqQXvLQho7BYhM0yU1MZ4sPMZ3D/SRVeoWgePv5tAEPzI5NMLYF1
cLM8hyhgKc7gMm2uEGVLYS5rCtf5s29xOIOcolj66qRnbECdWF24Psdpnp7wBRW0
Z0Y863Z3sn1luyih9nx+CrWDpzd8Vrh2wfsaeKEdX59rrS+D8VCntgVWJ3nkXv+9
zAo5jTpXB2wq1YN92RfUBvjQ32EiBdpjIBQ5rA7ZYuGv3IMvAOYZ8UN7q72LUXyy
3q9M4+ZA0uIZKifrL6aiG5X3eIap9EDql+dmE7V59m9xKjpOJ9+sGahX1QXM6dcd
dMmG4idty9QNDXhdPkES58rrGO8waZWz1WrGECY+A3Va74jWThjVENv8SKDtH6BO
4qNSQqg4dn1iJ9s4A2cyyHz0mHq3aoQB4r2BXxwLxjNtkGZXCdFnlUkSctkEVfqE
WcsAC4xaPn5hVb1e/d3I/Px23cWwctTR1K442Aen41xMPvH6RIQqXFU8cgqlLObE
7PdNe6FrVPuK7/+K4ja4UVMBztrKEFAjyUNsNln6e27Kxh1UObbkJNUKCsAjyg93
HIWjJqKvZpqOU38aAdLL4lMRQ1cTwtixGOQgP0+FINic7Iz1J1b61Jag6CiCnCm8
W3QmHsiBZYf6iGtjLDV7blsqqN8Z3Dyv67sWg4zQXkvN8jtj7k8Cf7Ajgnl3G0Qm
/r7VRirMlPHq0y197l5FqptXPF3XwUo4ohtnVmZ12C0heaap0EnS2HSuXjTwVoy8
UzCoeukmWy/DjNOmpI21RoznPmQWAfdd7vM3JCL/IEiWGZuCOoIZ/fY21JtMn4s2
UZbCmemiqVUFUTLcDrSdi/eW3gn3a8k+pHXbdb/PokOMdBovI3/wHut5ADvQqAN4
oAbobRuXtJZQ/Shl2FbBzJ+TwHehZJmV3mKPa5RVZJP5iij/J70TNl20uHRPxU6G
l+gjeWJUwyxyblPY4/Zq6tAZXz0VxDSVMPQX4LRJxwxpKu0KLjyne3Yp3hIhPe28
0H85YJ2SYN2ewwGpPY+GHnqXJdnVzBbdvdLWqfsH5CFT9cgyanacWHFRQchRAz6G
MY2n0RbXJbKksJG071dHBc7P65zhahHoYQgrvoBt++5Vy2bQXBTWMAH5u4mJswYL
909jywF30OMIL+6nSZFDboIBLgrJ8I/WOZJzd2k7iq2kQAbgTbD5/9EHN5fH+XAt
7r9oqhDLDARIA4eXzxBpmY+C6+u/dsJXgcYpNBKh65bcNXYqhL5AkRqkYO9qBRrx
rSr7ou5kr1tAa02b9UYt70M3mRoGO2MJn3sIRMIJY+o0MgZFsNkutuD2WtSCM4NN
C9NN9nXe/02Cj+xc3l04w6u+EWltJYslZ6cax3uwdpdzhKWBltZIf1+5KgG2CdCE
6Cj1DoPRC+fi1MhXJ4BXJvufNOQw2frqljG3Vq5+RVFehbl6KUr1rhLhUTThQ5XA
JuXBFMIAIJeAZ1oxhQr5OJcmzgzh5G+cMbkLK2EVY0/czkr8A4I2GTI0jbWwJ57g
7d4Dqe4HbPDAKVBTsVVySWxsOzmzGbW+xVLpDk/zxSdeTVG/yv2KdFnGXSVlLX5X
+YZ46rczngiqlwGV/fYT4MEEkjEk4fXK74m1AvH52BxwPN0pG8KFEpEA+ZykBt2P
d2ht+cFQkgmdhw3wq1wzD3snOxJzZ2Z370KCoID2b5Ko2DsVq5YBoowvySUW2qbJ
yFxuVX7BMZFPsoXvUWElQzR+gVWdicuiRxeUSnPcZAJOVGyIjF8SwD+HEbVQkoC1
AN/COplkakEogzW4Ej3r3nNpk4tJ+7/yVnNPGitfJ/dU4tEfsy2fK73WJZRG1dB+
c2Qyp/je0pBnD3+gzoOZAkPEsT3ewU0oGQ4H+YTdBnzC5KDFgW/yNa5BEVfA0Q8H
5NNZTOFQ1BXjtfuL8Hf7mUsQgMpEgokoexDRzzSb3LVrCveSUeIXZSZgbwlyeR0j
DYirT82NtE49Yr6RfMCWL0zOJuP+sM1721C3jiKjk5SEMIQBBPtl1aOjirHJBYSL
6xr5xwhPYyeOH4YvWq6X6tOl30/GK78Lv93Rv9UbYVbmI3RlBHuD5+F6UjDuHO5a
+GR52leOaz1qkhXq3+Lm0vqSbBzlvJ/QXAKSMeX1sA3yw/6gsu0Tg+aag5yfU3YE
AcnzpNL0dZb3q6CpH3xVD9D6ZS2Q0i23unTSyJN3zEhkcguMElRKGv3d/q+9gqmZ
6w0DY8VuDjIfxmtN4ZnFPWV7zk7ifbhFyOXOzv6746mHz98jApey6aIBmR0ObD2g
w1XtinVmm/A1J+FquKh88rqKWp2Rt3LyVFb1G1faxF7btQk0dXdXemRgsP1avaiY
VA2sQNkZqRI7s7He2EcXj72EXlovWZVWaPN8YPrSL9iCKexAspVsoG3yNKbaYnmn
Sr/ofxxJzYRTHILMfNNE9IaQyV36LAOHExMAO5p2oy1ao0gcFp/HMjpLw8mOnob6
8xiMMUxxNNgCU1N+CK0CVli5M51sclo5a8fBIe5nHIb+ghvUsB3vV6KBkiKQFX/M
4rhD2PF+9wqCksGGeipH2K7PVlbA/H9ERxH4Ufa7kmWY3AJWycrhbirYTAraOUqW
1WzR2+ofbSMMk5TPfCANvP6I9zjBSdyGgZ/M5LMstWxr8VHlB33nidrX98XEXI9w
h+Z+L6UPP4mwjj4M4NIKnIqGVxnY/IhlP4MQORPFBALs581hQCVqg+lFctng/wTZ
qVVLC+dZV555EqovbX/lc6+mYDJ3QXHcnbSMX/TefjZYwlUUoo3TmaP19cmML5IF
9YAWY8U//r+2OGgDav6X7IWw/Oe1XeBq2X1qHt22Kg4R13IgzJqort8ZWZFquT/J
tcpi6Czugl7Gs/f5+yKSEGtpU1K4teGmvCb/CkF1/zftF4wFto99fJ9T7XQoqlXZ
dmLe/oPopJxRZH+BzaRXWsyddDA/6d2B6a2PJ83lFBMduOS14IYoIyJFvcR/h/VJ
XU95XljK22sSPVexzpUclqrBaeK3iFHtWDsxVsRx7SS7CYX67xUMqsB7VV3KARix
sWbgWHCgcJ38qgATjJ3GdVlDIeuuc0ivW4oSjY4b/PLVe+taXXA0oVpKASqXePiU
znZUNsCZq3mf6sjp5qvZpFi2pbq5XSOXi6NbhM3/mBoTKcSBw+NyvwRxv1v1pTH7
hmcVSYGHY6sPjShYYsgjklDGH50etYZetR6ySoVx/H8Jjv3MUbiSPtcPwzKnr/vE
TAFqkCrwXHCqiHETc4kvIedwjrGYOK2UJMMtPBarbofG8T+hqF4UflYeBzmipBP4
VbPzNwUIRlJVgwhI9q38QvX9ACaO+ENRBYIJjd235es0Z2zsDCeZI/bxBZQFtvHa
C9k3kCkK5ct57exX2JVtkOuPfei1YI38iYSjhs3LQInFFt8CaNU2gv5eUwFOTRR6
PIz7kxnEhf5d0Kz7Xr4iWiX5FjGND3uPRnGYcLBu1UbB5eKJjWcSFYSZ1wVPANat
9Jwb9MdVMSPfWnB7BRmx+eiGiTfFjuR6jL0H5TmgdUctTzJqlhOM+ukIY2eqXfBq
vucgDYFzRck+bMqoBT0KGdZgBTqXv8KjgjTBhsd1QFDsF9PEvisnx8juPDFHJYJw
k7P8bIad0MeoWoQrMSZ9JrvK7HOaUOu9pcZkkM+KgAGXfMKbl4uy1+3eIzLocIln
7baOblQJdICtXLlwpogSznTZXlQRFQbEM2BvVTfR3RZKyZb4kTxTZcZ7mGEFjus1
YcJwTpze+lkqOY3Mf1DzoEsv2+rRfmqtPADDGXxEFVi84E8aWoH6CSOm8xQlqjhO
GGAcYZWqCzAduBjZqOK+BXl2JuEWPtnL8DgoJFSGO19SN8Ks7FODZ8GIVMAoe07U
+5MgXs5CQOe5JKDg/K/tZ0I4qvHSGmIsvzKC8NTD/6IyvfS84jkljgBHr0SDkTNa
xdcUBUev10KkiXw0RQEt22xxK58GA8UdKEyHONVSsTr9nWhOhBFXKsaT+wlBx0AR
AZLVwKY4T9/TNlGOggKv/MKP3BQmhn1sIxeqdlHgcRaskfzGfV7UMq54Cvx4at0e
EiAvT9T5x1m9nHKyYR1AEwh53DlJsTVU+Phmm2pTz1p740vlG/NvsAJ6swAqZo/s
UB2wAYM7XiIRe7S4b5yD16VnD4xGNUA2GeWr5Vbopfo18dxmGO9HaPxTJ+cJ44Iu
9yvfHkf2AQJeuJnKDcts14I0NPCgBv7UXHxGUVmAstjtXwixq30DTibA+SxTpaRL
jAD5faBDTEqMor8bN92wohj2A03M9k7pcWFF/uK8ndyjJrLO+K9aJ5+Zi0UrT9Fk
eHDrOCkxvjD41sMPmx3u7duylcckmTPs9xyEbkFWqM7+9RqoNiHUcIc+8TPCIx22
puebyKssQKhGbPNl/jZXrVQ9QKulL3U7dRoLWGKo7+lYHWS6FyoEEpONnVD6Uwsy
NhQV27Prh+U66BDh3B+p9b+d/JeiKdZrOgPPuPhsykvMqsAsgMtqbDbjt2NeeIQK
fdfqBnvQdclENfMY7Q2vcUtbpV7ZWwPPX2BamXRs7hBBp3vWhirr0xG5pDlFQ3Go
NWNsfPK7ehxYjdTat3M7za761YVkrYgt2b/kopchlJGdrxnUOF6yigYGQLxaCtOk
OIIKqw4TgMRjEYbAaDLAS8bvFInNAuuz+Tf4T9HT4rCv+iFsGBXhe08ovlaK/n49
5PnTbOgtprWmpLdkOKBVglsl0eb5fLwzkiY0SEH/9r+VPHkW6i1s8nOldnCYVjoB
Jlg2ocALFYaSHfABtxd8UzoYq4r7jcnan3nqJCX7AMy9Js7hcN4b2d9oP0LbRlpN
bL72EFlnPvxNStU9l5KiTcagaLmA+44m+xJBFbKhClhxp36clD+OqEm4WZz59MSE
scWDBns9npJ/vpTsMhgDGNT/dnAKk9gXbX1B5B+fms54featLPZScKx75HVjKUra
PEzg3i+dxOTkjwhducRJv8vZzwRD18u9FCvPOc1lpo/WW4IPQfjyLqAy+031bWIK
GSQPBHSop/lejbXoVpnGzHCm+k81u5hUXgYIPULuhNcjliJ7dMxKqeo4HXhcMhCa
hv5/yjk9IPaSKMmz23eZyebo/pDX9mCGjH8EU/ZxBQhw3nPW5QiKrZET+cdBonuy
5n2FbkC05jF76EzvIA7NiUYFaeZj/h3rPBfswknX3zMv6skSdf9iq8Yfd7gITGzu
aztTqFtb5XOPlESdZeC0+B8EGoMoPoBRvIQrxEiVcDP13rRbffl4Ge4FXHlSvgP7
15sYEBIFBFVymBch6Ydds8+sVloxZ4tUXax6GTstdwTyIJIA7EuBhB51m5KXuRTm
CjbFewhnVVGdvCmH2dcZs/pz2xSeJjlcs8Cs8O0JhPqPxTn5g/j00ZFwGSpnxjYE
+ZfSxUvHR1ye074ppXj0jrapGJc+NihxddwQJiKpZx/zac5zW2ojfcTaAcVtSTlW
xeD4I7xeVmJqX76rjF8vYnN8ayTCdCbAMaXlqA1XruHiH3l7qbhTT49DogdY0AkJ
sOMZ8So3PLCI7Ri36J/8K4XIyBvELiuS3fSW/KLkz+xCMsiov9uMBDTwhfzEwSc6
yppSnqZ8uovpxqVD7oMHYX8ZLK0eqauFerM6I6ff9o4H612rUTkZDcvStn5b+KyA
UU3gNwUckPjb/dNRdTftlm6kp2eL/nXn0X8myI6IrKCEL5T1K3V/P9xDVgavgFhk
X4hfoWyDrPTc8Qk81R5rtf/o/eQgwah7i7eavukF/rUBTXRhvxl0miGZBgNyxedh
goS1QzP6/xaCGTcia/6UDlMvCCsBvkU0xXM6rNBXw6dCESSly6gozgnYTdYT/NSZ
1S6d1JiZO1uCSIxc2WsGj8nyN1kGk6/g2LjDJRtezTbuK2fLn54Z3ksG8fapP6oU
NrTBa08TSQigK2gkqispUnPSaqIyafuQAdY8Cdeim/BNXjsuCrPniMtaMDvgogV+
2Gu5oMFaT3XjUJdNQMrpw5DocbWzTmOLc5bPMF3ROh0ao7oA6EnoOWP8KV9pg62Y
CDoKAkdQmxSjRKRK4aZ0PfBpzl/FJogx6ptkvqwBCoYPPQGGtCUGOmh0KSnDh+qG
mEXVnoisM3UidmcF1vSE48EY+Or/eh5rjoFIanB0DKINbORkggok7WsRqkrKL6Xv
agQwQE4ccaYk7B75O1s1RWUMQCmjUSe/LpVTIoZ1Pg0Dd/zpusV5VkOrPeCmojrH
wj1ZJ997jkVIRqSkPAjZzPO1e2mGo1C4ggeHjFT80uXHDN6rNr7Xxz/5VceWQebi
FzE9QwjowOAypvoqZu9IDHUU3pp2K1bi4+3SccPUQ94wlakBYkiCnaRXKpNfwaqx
1VDake3YZxlzdir53/yAJ+jsGliOkAFVvxhWCw5LhNILfXCjXkKB1Dc26ESNSb3R
KOEyBp4yxSOfVrHg9oV43R+SxmCxbn/fHQ46T6/GIH/LjvnB/M10JCq2cB9YGpBl
fax4AnV8tgjsVGWXTXEMgeEo6fIgHTv3hhD6EUD9cY/0Navlcm1gHhltjrdHz4gd
cruAHGOMHCSHmOJjVHLWm2KBDTaXdjqDurKlagCo92KMFJB8GZZ4CliNI3uXyL4i
VCjzA8fSEan18LY+7ffQVvaijhjVVRIHHPdTeYcdSlalu/v1Jap8Ixw2e/ZaeB+x
YiXJ4PvdIKZLXQzLsVUO3bN7tv23wtsVRTjRA0lzZLD194CCjpLYcQAJxYFJeosR
YyhCTcRiSkovVvv26Zz1y4PZPaGVXNJmMpcYMz1IIYe/xkGlv3/tkKYgOmWZpDVX
7CM4IfcLG8giP8kZ5rJ6QadjE+Ql6Y/Zk+zHrlrr7Q8Hjtl85D5zZYJ8Mn05lwIU
90nupZbJStCaLQcRj1OWNDb9zmn0omk0vN+ObOt7denmbRM+qwuitzcXiOohHf18
sJLQVM9ZUCRgIr/SCp6Wsp9av8j2YtJMGvabw72U3Fousb/Z4AR2feSJpykKGQHX
04tJ5+lT87BM+79K0ugUpxsI6wzXI6UcsyXwt/A1ztLgXdltQHTs95nWSosBKLvB
rt9JfMJnvku3vyIw7SlIHspy9B3/3LJEkUin1LDnKI8ilAB5qS9AhLh+/Ru9RDB7
UM9T3q6CmT3cmgoHmF5yLiF8zKfEx75JraKl/pTZ8129HevFfewcOT4ZN4xo7+Rc
jPLvjlSlPfoV912dUK8N1l9W2h2PhJr8NpY/DLho05oM0SHpcLM3AdH6lIFsHvfi
VgZjUkQ/Ys9ciZq0oSEzEcuut7kl4JUL4KjUeD6SrKhqb8nGgJhCPOlogfW/LMDq
PYbAMKOCZDG2AmO/rAQEBoBSL/tLfxOHRYHvt3udTpgWouDLH4tINpk/mwLOIkUK
6pyJ668QiUYPKWAAJpSOEc9M0jK5+ktHTC2NIJdjeErxOmbHVkblkqCuFXCYF8OQ
IjEXfK0hc+uoEwxhqoCgdCAnBOjQ1TA3eqUjT4hyQt9BNofR+OsPnpzKDuHfi3RL
Gf8KHjeaEe5r4vVivqwUYWAeExOchsjRllFrKWBmhGSxedGkkgaqozSj3Rnhnehz
ocmSb//vlyNo76wZjZjLZAOR6k524tsSDQp//x9RTEWt3AYTQtvgU6ifWp2B/GaT
ajWHUQaIPzdhmYTqJq8Gky4ZTC0IVNyMGrN4hT3G8mqCZAIb+MbFCiBju3b84rS6
3LCP2Xhr0JnOaXSMP6UlDUEkCcwI2osoMMFbaKOmLa5o0lhnUE9TUF0jnm/nxfeL
wIhik5qekDDHTu1aUqM6FukAa75dHDShUQvXZW1SCBiQnFTbNiYDgKC1lSRQx9xr
duzV8zr/UxsnoWXwiJ3DVQlEJhOvo2svD0FhCRRNhjqcQLK5HT5LuXACwSPmihfr
uCWdr5CvENyf9oUvCatCa2m0SHb2+NRgcVzMkvQPYBiMJDiPbRBh+83I5l1EX/mB
Tz2+8jeYjSg2ra2HI1uU8kQWRGn0p7KWXE2iic/ZsBgFzrPxA3j9v+0pQ9wGcNZx
uMwLLtDPM9+1VPMvHlWfP3czt9LhNQ9nxY5hOaHLo9SEOlqEVD5MSAzPDd/rOXSJ
+gdqloSAuEEDVIX87hXBhIyWrDt2OV7T6G+pVnQvRHHC5SBKVaqsDO3iOs9KEVBT
DYXxQeuO+jTC9yAOFrdgDoveSPs3olo7MOingZ+uJzuXE7EEWjxURDFcA6NL4g9k
GVrcPb2lhRrxv6GKtpLzIesu1XdOJt3fbq1U6gU03Tp0Udgxw3SwfDcBS7eg5NtD
zlAWw0Rm8LsEBpTRRCzjgYO8tq3yJhYME6HS9I3Gm8a0WBfzdhxs7os8TgjrP56X
1u108JK6/sXfLdPIRGV9hGNoHToE5bucTqdSttgnFgSDwbfp01GxrXdnUFj3Avxv
Q9bsJf3XfyPykNMnvB8+rziwdEq+0u9tCU3nBeiZdPLtGBlsxFrE2cyDg1QpUZCV
GjqYIxo2wHJ4ivqPSjLCOQhxDH2hBe62DlxJwlZlhtEj1R3Fw9mu03UwUvVwTdqA
x4PpkzSTN8hsYM2dskjpNPUNJirJ9U0xQvT6dgUVMOl2LiExUdr6ZBX9eS5C9xpN
p0mNQtKMb8O9iSBrpmssQkOD1KgQXT8hWxvb6d8RSGNzLCvyyFS3K9kgbUH7ztZS
V6JZqRSOBtwiIpR1K488lxSF7W5fhkoZqFTY80X/Ymji2YxDIZl6vnGrnux/nA00
z/9TqKxTKo5xlDt8hpcfCFVgxXucn0LCdXJiYuR469ynPOan1zrUCAwZgrOG7w+k
nMETBPy3UEyq1FrgkHWXP9Q2RRZ1ibhoC2MojdsLZ7hOHLdJ9aLJhIp93cNye9ZW
hJLJ93dtiEoPgGTqx59xGzO2Sx7xHlma8XxxkJTi/mnkwvrCaAlqcSyBQgeQLXPe
etRE1cgNjKGGAnZXS9BaThgRR+HAq2SsiTiurfHpjy7zrMge8y9JHogRJBok0vDP
fpKXZkGO4TD2IYHYRHv9YSi84/pgzYK9n+ZBgchou41oR8x9xHrpdzgHKZQW6Vme
dgICHs7YIydcrxgt4r77XqU9mpfAHdV9C8kKm08BfBFCcJbZwJG28W+oqwUmW8dO
l2kySDgvfjsLU4Oglo71ZLqWdqANujGIsYhnW55TDVMwBXv5drIkAWZPuuzKtTg8
v9dBPZbt61elW+ZFagLeLgOU20X2mZfJpgDI2Cr07kOClAsRs6WOgeiig0u5jXUu
JzzPakfkS+Q8fR31M9PNrZyhb8+ASoBVj6K4ZGkm3J0iwezJAtaL66Smu8X/2Bfz
mp9stb677TBSnS8Y56kWkGjKlQxXENZ6Is1smwSJc5lxchYqS2MLX6Xd4lEqd8p2
Vt+kCsOdz/SpJCPYHUEOu9eCv3xORHL1KL9KMTdRfOWOn5qVe5aeQ94c3nubDcOT
v0Tyuc9T/TcpHYaS2s5ImG1Cu8IcTPP4H69sEFB/lxF/FukbE7kr7Az+FEnkNw9j
JgFMD35JqON5rV9BNe9PWNnUEQ/lMZlYla7hpZQFTK/XubbEReRsxZKVcmd/BoRk
deBnZK1Km3uP7O01OgPTc47BKBcc/bge90I/vziMVG4Dby8iFfTKImBrdBTO9n4A
cR4KP48zayh8c0qcACwA8n/xFCQrqfZLi1y11psFBHdAP1E2OBTBrWG+uPxkHRiR
rxILOkR2v6M2AFQutsVGxE3nduk5GkMyWsSrJ3rWwCEjaN/PdEfrFQpSHgfqAb++
kyfFAR7FJH/bFptkj9KeStAbb+dOnXCU4Cxsm3cGrl7iVahc28ZpqH4LMVjKdzFu
i4DeknM1tGhertx/hYjbeGD64BYEuzOkUhGlEo5sXXQ3x8aMdiuOvulbTBCwUJp0
dpKnpsavVbhYJQk8sOnkpM73UA4yTWZZbNlzjCCq7qWJjKPJIbxQHvMMf4+yHGsU
XoQaLR83I0zJE3p+stHh6GeOjlcquFfM5mPAGUXHePX9JyplQBvDsXOc6xjHXZah
t//dCUP5LVeoc1gAjXI61msT4LD6fU/0BjBdfhzn+7FB94Hsy4SQ7vhmcu83jUOZ
iEoDyBosXoHQFB+Gzigc8cPJ9yr5F/c9dg3MXa9YXOG1kqbSwtlJllhYk4kU2UQK
0EVVL4y+oUJkDkgtG2X+IKc3IWBJ8aR4yWk8pNr0YE6dboGy96dHyR3uD11A9JSc
QFZ07HK+wd1Y9cXtoVKg/dasxy0aW6urOFtdVVu0yd/0FRQFdHKoQN9AYQE3DX1E
HTs7mRtIhs0eyHDFNg6BSuPXR7m13A87jO4IbnYq+CB3p0IwdmLL1Ys7Z+VeqkZN
BxervN/ofHh585gln8P+Gw5ZaSCmf6Qrm0V4IcVALLw42GjNuFBJzNjsZJeCXDAa
/k9vLOJAStYhBZYZUU2XpIsJw1OHhx8xMnzi7YeTzrvdefom389v3Y1ByjKIq1MO
mnFpXruXy8gnQwkvjlZJC0e7aMVaVvfTDF4tS/4pn16eUtK4vBx6sZglxRtgyiwn
ykO1lPEv4u9lh4dhZVltcHBYXui5wDKpm5eOyfGcPWT7o5I3KkBtXUG536VzWxLu
4xDsxShaoxWOSgutOymmD2xkit3MirEOqAW0urZP0YSGur4c1jtbOPx9MpckUAIW
NQkkAdH0Gr2WNEv+O+TjnzDK0TsGoy/zTqniIlOn6Qu0X1OMTW557FAYrkgNIbDx
wb5r6EDmR4JUU28gUSB1e6WK8zLgNKqGgXy3vrdtVcD9FKsL2XWDYPk0lFP4RsXc
Tnt3Yo9+31J5lgmCD89O4VPuT4o7mZcD1MZatzMUWXUUKTt0fl4GY5Ae6hWtlir1
JMXNvYuSVfBbI+uJmKP8hklszJtjPQQICwwKf8xbNx30h9x8wF7xdMyZNHWUxyd5
nANWNS7VetN6I3Ns11oUbBTGeucdHSuuzx0dae2m/0873BtpZ07YR8bQ4KzK1SNC
a8EqzNGH1In0SgeRw2EYI+VHMccfcdOBUs4D4+TwLeeGi6lDgVPpVxvtfamJunsF
lmCq+CYgQADC6/2WoSkcf2JMX/zz/TmJO73pDGgXvDP0L2lQs5qX6LZc8giiIQFJ
WcLajl4NNavKTMJjEmI0Vw6BbT1J4Tr5RYKMmXx6tixv+7ogTkwBEEvUn5MillOV
tG3MWmXseN/YVvl5fEi6mRXZ7VzaUoMpRGvy9lAcSPOaPofY/FiDQmDS5l3O9Lqg
cUhhzYyfguNXHjgXks/s+cQKT8XrHftZPa2XgPRaBhFQjPN0n9teDUgpNBRFO5fK
nNUjQc52I0cNwh8/yHaIo92ciRwTEkz6D1pSkFyPXZ95AFoLmKwDJqT9gJIVwZw8
6Ra8dxeyeZRJCbFaaKNfssdeKHZ1dGHoNPm4CHWCenpzkGNaD8X+GQ8/7+GIRA0Y
Da6iG4b02pIR4/GzZjZTWRsFNE0Gl+V8wMNqsn0F+TjhOA2OY8mcPF4fFt964LYi
bAjf7qrjcSVonuHboc/a62WzzRXBgB1W86McnckpM85lVpv2+YCIP7BusaEH+hdH
EVT/SBqo+KSKmgveQKASYCmwTSpveAGIgA+MmUKdnFBbGiQg9S8lw0nvCKIfZmkl
px6M4Pt1IWfji2AvaZy7pLT4czDaZo3K8z3lfujBaT+HLIgqwlgqmM7yssMiT/gq
NGOTxnU6rC3oHRN4y3MSv4eCxHKLixe8kZUGgxsxilSpQKkDaKF8+dSGYXkUvWlC
+H0bjmpEe0TDWWat4TvfaEbDAHFGgVFH5a1Q28PjvYuqhdZ4qMVsH9yb0ScgKoTJ
Og/keNgvqL7em/AHGlR0WVJP81aVOgJFC6faU+3CCO4eemBLOYs5sZH5aJL0tajk
uQJS9r4xfKDHzzINznD+TMwkfXKSpDJ/LhXL1Giv/QS3zzSnfFAWUpOmuEE57UgX
86FE2YxSFdHd3vnC8fr/Ovl16FyAWop/gB3tIaLJiasVJLDJMIFZ29Ns1se1nWIr
xQU7E27m5ftWfvWA+Y/7iB6BRQPog72x2wJP88s83qkM51yXaVqCkiM5aZS7dhPm
yBWGp8sO45FcGVqluOqrm9rSkbnlpjKMY3hafNX5C5/jwDc5yYpWogUw4llUzBjV
N+87gTrfqE6WEaMmzDT5Pq+w7a606PB+y4RtQnofY4ek2D4YqZcv6j/w5NLy2GBq
g0koxrC5aUll3T7EnUPAG6T35l5kqHnYZWbCEysdEpEvHhBjHwlGiYt+XJ1zm4ID
5ah/4E8BC0ZVQVTJF82SoFv9+RhJrMh1VIHFaDGwJt4Pb+Ncn6++Rnkhy28+skOX
Xba3j48XPNdR3ucsxHDrXDiwE3QGL4Al88YPQjv2LfmJ6Lt4SNxh24oEBHoubd0f
E0KUwb4yqlg9R9PkZYPp4nbKpfL4v8OLN9tpuNc7CatNxaZdx7B/9liisA9bVA5n
bp94ValP74aAsOuKnrGEigP8sz7G2czpr6iWuh0UFeOgJtLcjk8QywyR51xxhKbh
Smvk+1mUIydHDjMSGW8vHxM9EVHId5JkxSHuhpFeE1jZIFwrSy9tYcFUzQvvQWf7
RieKRF2bgrsHceXWawVrwvdeZXT6ZG+cw4Kl4Bv4R0MSLeEWu3u9QBjtMNcP2CXN
sqMUjvvxQylU6FTE2ZXwphhJaq0+bEswdvrhkDi5jhY66dTM95uYO8u/6pB0XJzQ
XHccYGajWwovtiQyucl8rKDCI0dAEqqBITisc/S6TfyZUyEB6/5l9r510bkP56Zm
dvftdq2up8wXydKjiJ9htcR/7UKwDHAo3XQhpcn2AjA42YGNSk118T5SuXSwwUIx
PuYReFf1kXKLSwUNTkQ18g8GA3KiWacfhdTFDoBt4wQJroG+UiisA2hLIy3Wuibg
zvAA+1Ps2wYt23qC5kO4BHiD2sONcSuysprnVQZdpYoQ5omLMr+VK6NUZL0VweFa
jKQQ8u7fO6HJka8blnCDUrRGy5pA3YX5uDVGfZaEtXSMSQNcCf+/l4WXCoNdKs9h
h9iOzAj5mz+z33gV2apc+sogAA6RLXDjO6JqOZB4xS9kyE5CGiCk4A32iKL908yQ
Ue8pG/8U5eddRKSghvd9xdaQogs3HAce2Fp2qvvSk/2LwAq0MH4Z2hapEmAllUWH
y5IuiNoEAU8ZicEh0PgwzJILDv36+uHfDVW316oGTyt6n607lbwdeWkC9w0wYQNs
sO9KxD3U3vQUsuZ5+YiW0fXgn8Uj8ThGulkUUwLKluw/mJeo0SjPTbbBi/shCj2s
bltlv5nCZATkfa3taCOXHqhSbWJP1J1sMWZ3AP6CszmZQ0kLc8BRqj/rmDBGyqhV
6hXRFd56iz7aIUzsHEFrFVc5hjtZepJ2f+002CJek+34HJiR/WTb4xdgWvHpUtfh
8KPSuROp2J13bQiqDAbjHQWEWEG4fROoMsMl51cD0gykWThoebNWYgXXHVzhXGqk
X0+qfP/Vl08BjsyVvOHOSWDKKGG5H5QfSsjgdejORezTPfxts10huVHjyQ+a1gLX
hFM95EYmhvYD5JLgMlo1tY/qgSPxyHjwq4XWmkLcTX0tB3czjEeL4S0l3dbvtedc
nLLSSwltIDvga89cFvSrQTZ7O/ofhYwFmolmZwBwt6SkNPv+NWw66U5o5HE0kWIf
JtkpHTyeKOZe9RK4od+ZrK9kP5uCYBD/Oon63TPd/vpYHfEH9CDXBrlrtg2c+xHM
H8ymAmnykoj6aTDIyP4MpOdb8cW/M5dEKbDvK7whHnlHItze8kFvv5EDd3GGmPgn
Yef7CEXyb9WQJeeSL4s0R021+6mK9PwVtY3e3SJMckQhOS3fYajUTdicVc4fnUxI
ALAQAZE+SRgC69c6ka9S7hErlOfWDfnzO0YOemd7Vte+jka2C+aZxhVm8pFS1DL1
qZngCvkDCjqJV8h9ll0ZaswQbAbdYG0q20qkiQ3SilFnFcbsq4600p8D42fvUSgx
6kCQZY5R3OSRkvh/4eMtK4DSfnkUeh8gYkfVwPXwyJd7wcX/pIfS2chhqSm7yhNO
SJgn0u6iwT10/hPpQleEPoiL5/ILQLVHKYvN20qlEpqT/V5wSLJWPkj+S0BbPItX
UNoJcUvjt4IqclH4/tqrKlyIFTL6qYjaw0Vk8/77kINKYN8GbGglwrv6Xg7rItqP
lsDvwv0hKudpZv48yeBt0DllwEOzFu7S9GQXK0fBJIxe7xXw62zZIl+wQgX2fqFI
M3qzWMxtfK7NeE8dZVpvH7uCisuMffW3gCIBJIGJ4v1rCBmfi36hX/1mp8a/s6bF
Z5ZirIILBlIK0UYjYt1IykBzBDwcDlqGKhvhOywX3wZgLwdX8ZAOdtw1EWRDyJri
BJyLe8PfIhqICr3fgGMw6xONBNC5RuvgrPd2iV/K3mO4oXWVviH2o2jVY3aZkQ1n
rCiChTpOHBBeobsFSDIhy/sVhPvdqPerDKpr7dFbop73ojESNDe37JzvbwJbG7bm
uqFtutKHteZLzTu5ceSKKz3lvyP5mDZxIsUSB2WK5DPSpoI5kdxiE8SryG13hYhN
StQ3lBGM9rvqpcN2KbsAphjMZsPU7JlSiyvHFfgbJDvWPUEyPuTplZapp6ep1LuJ
6yipv1Q/mqGVTDjUmk7+ZadK8/EGBWKRZ51Jb/2muQC3tim90LM3tFNuz9gep9ZK
4tQeEF06mzki3ehmGfzi/ThBNXWyK+xWxK0E+y5UzSuQheV2sY1T+uXY0zNlV38m
fl3pPu6igZUXh2x82XWJx0Z+FC9n7OEGpRaKrcwR04KF2HKM2nCbX6ilsCUu4efK
WH/w91bciTVjmeKeJnSZlWHi0UAl7UmGwcihJBZ/MNNe/EZjpnj24ocKqPQ5iMal
jIaSCQ4kgT3p6fK/rYdqfVXkXlGvwim6zJPPJKwy0jA+yLejd+xAwqYFxYiDM1oK
8Op9pEeNcguN4KSrXtxsPX/BD4Wc1tGb3GynNBGeKHJkJYY8h1SJo3B0rlrnT28z
TQlOkDsZ4a9fDEYOwkJd3RDfcYpGhVEeh3tvpmJ6EOjE4b9fL5GBFDJet4Wh9oUs
LMjBFSG/NPJgPTFRZPgIVwqySv4lhUrQ4Cg4ax7SkFihImAvrrqiITlE1jlHWTJ3
TOQmeBYtA5oscd3BlLa7DFk75HmE0jq5rwKB/cHWNXl3MYhmqlM/zYXDxZ7tFY6B
AbcmblSTUthGbUPNg3IJNpZtA8He3E5IcvumfGF+Fz8a/Jz2mGuta0R5V/CB+Pg+
Hd/qaWR1Ou3PuNd9/8nacaIKlXV+/XTrRg6mGQiZZkDzWAJp+a3hBlDXeBj+4WCC
mnhzVm8v/2ch5dsjnVr0Nj+ZMYdx+uauYRho/90CdqlXTkYcykUpx5Ng+fN1mwuE
YYKZjM4SjgaoHx6OK3KOvSjfq6kq8baloZGp7Nr5EpCEfJl2mvCotWd04HIjkXAv
JmBTGRa3A3LCjmscXCSJvlExxNjMDeaHytSsbbiWrvmck/zxgzxr+4Tdn8gnnX6h
zKqqk8W4ZmD65Cm+1uWZlnfLiCIv0hrvKG27Bm5fgOZzgQMK6OVkDLdToI9iOuCb
ot9cDwMG9XmKJhowutUswmfdbhBIfjOQ/gahY23boPNVTFb9HXfu3xzSrUd+LQWc
UKJpyZEYBYHh8+yxllKm3omlgf58nNKWtr6ktAhSxW1ekGM3W9EoEN1UvYWZPy8C
9OTdThRiTJBnIQ/eDPlvHGbISWc6IPFrFcPAlfo8LdB5nIT0Pt5R44iJej+bEXrj
sJiBvGgabL/uIv3mRE3/X8nXzzO7tdDvEYTt0LO/xupbFQiEyFgY4dHz/zvtg8N+
7DtjkmK2jABAfpl5MJU+tiNulaJWI2ibdyE5CisKKNPxPH4VayjPhCQtt7s+Jpz+
ZKR3c62QLrZlD+e71UMNQ9jwMkyf0a4waognBt6xbcxJ0H/S6aPiuGo1j3INDJJT
loUN6pFo/fiB+y1E+E5ixCIgqpfD4WMUQ6QHt/eyBDUrvErTGaT0+MI4uLSU6Sft
Haaa4g7z9qIMcXEnxXD9MNZ67Lt9yhhnT367qHD+2/AGiUtqJ0DyFQJIqhopN28P
JabVUxrS8fb4bsxiQA6WCf8PJLhFTI5mxKviwZtRZZI2FsLDPRCC3eRMDDFQqHdu
mA5OtWRjvhlsPNhtCuyS/+taMSc5LOtVtLK0Z0W8eQ1IUlGUlEwKlOTOand4L7Rd
/UMByuef39hgRB08u//ji0bvYpxZDHRzBfFkdPV4d3EtTLMZ0RGx6DPwjI9tOU9c
o6RqHvB1epuYWsnKof/JmAJ92S1dLxkDFhgArVdq2LYTO8Bj8IJ1ZQLybniwQa8p
lox6yDwHL0QuHaq+Iip2++j6WKswWEx15lTrkRvcoHdCo11ktGmwWKEhd5yrT2la
5PPUJwHqMMkIic/Eo+qQlJ0zSz4IN6PVJqbYCIGWiA41Pu/zsuqWGhZCkKe+EkCQ
cM3y38qLjLueX9UfJM/qs4YJ9ThIpVSSoUNaPMt3SYgS8rQz+eGGLqHkM7DL4yWd
Grba6CdncOve2R8v4sMRy8R2KRbWA+U9N7O9TmC5EN5082MNr87LkbUFhGP7IeQ/
NgxGjlnynZzenyPg1FkhBZ8taL9fn9N7/3Ah6T/PBzjZ7k8zTpKFSxwhxzKnviYK
H3P4R8RoAa2S2qo0HwLfBZjfXAqL3AhLP2LkwrUwCcAiPlU7NmNt/MD+SVv/2IjK
Tz6dCd0aPkpN6RiJsQW17sYFeAbJoB/O64LQRcmGtUYwwaYO78HEfAOYjNvdaEIW
0eXcAPSmVJdkJkjGvUalsa3uLUAiADOvYkQdm9F6TooYm2jd6U0rMs12+ujNUiP+
WS+p/hpyjUq2dmkqNXYZHhI+ququ+81AJwLQFG2rmyxHskNCIXakfFeyFXQArC04
wN8+M1MVdYLCZOBETBqRkx/4n4yCqBmSgXgMTnj2dM/Nq+n9D6/elEVX5bghgD1l
TmYmvkqo5edilEpoFIqYp9rKk5xumrF7xuPnrNiVGKN5fofi9il8d2FNBURLzGNu
FF6u46P4MT+5WCMN6RBhl82LE2WDQMzDyC67uin5UxbsVB+s0j/9HooO+ViYoA6Y
DSMYcUiPA4JHURok4+r6h2gG2+bHI+UyJprmpYQQMwdU/d4Owyj/dUXeSjlokbSQ
4zjif0Ak9unMIRTDqwfpUmRMF5LVHguCylJNWMjuxdMzQ4T8bgnrQbO95x2afgyY
6EPmKtRwHsFLGWwuJL7cW2zVgmEfkv4F2a6BLSUzcXrEGlGQiBh5zdRijSNtCWQu
VnrlhoRwW596HP8VYbuS6mH7bl4Ukv/QaTGPzxnlA7XLnzkm/TAuj/Ar0xTuUOft
rNMynkH8qFB1KLH0lShLBx84DuJemX9+4nd90R9q5oswMsbMHLaIjMpor26pwYGR
uOg/jZt9ewOwqLajgjLZ7N8AlTh/OOQ/G7Uc2YG9Df+BiKiGxE1mJROcY3DJLsKq
M3m2fnDy36YwgUyCRsHm5u4fWqlnJ4j2qg20Q3Ei0jZbkDjUHIwuss/PiBEi7Cix
jIO3ohaNV7Ox4tJDKbjFQwPnTPO7Qb2cwj0NZlRJfbRTWyXOrpGEJ1rrZhdklfBX
E3JOs/3VbbHYEvaFgOWU9ainpQSCjISPUJAH91kQTvMCbRV2BCujFivcirmw4Qp7
uixv9sKGp4+qrC8BxJTdzt8174SM5tYRu/siRp8jrryWdcb8mc4XtYwK8mu4TZRG
HLbp9kpitNHnLVImQVc3PXMCtWgfTDBd3I9dDh9eTcKTf7geFx1xAL46ecmre6o3
6R39uOkmXHBi8e7/GS9W+pNcK5K0bgQvcTPpXhL3GIGqwQfVBChgKxr5n+A0SeVU
UU71yvQXylO2Lh3JUvQFc5VT3BcWlR2jBEI/MgdngYH7n8vQMTIGEgIiNJGrACdK
R2I9oqA+nwTXBX0WBa5zP5aFC1MFVXCtkvLog1TYMBHvs/7S7j5Yu/BM3Ed3Gm7L
1UHA1x+LndN9XjmofZcYve1vJQqup9hposJ+gDHB0N75fbRjHv0Ipe+dAL4ByrGt
nrdP65DiL7+WLStIPQdS5rw2sLuqV9MfOQ7reKtHIi2Wt/iM1/4zFSeLg0vDydnl
cmsfhWKUx/i8BH80ipfYBeqMH8PRg1ExL9G8og8nIql+nsuUdv8kWE3Nk9446f/g
BEk+zFyQ1TPiV5K9AX1OAUD8xrXMU8MlCphP8PgWRzFRKfPeD229Pp6C/yD8+h4E
y1XOG0uAYPUlQOnN00txiDD6WnNvlhn/DoRlrG4ERoYxk9DZ6pIvH3l9EjqBc1Se
0nXpM5o+eMKy4Xm4jjuLxYdElgavkToQUKqgXCFc+Zlwj846vmHfn+/e+y9wpJZ0
72iYiKlftb3Fbb6Mj/88SVn1GgqVlHBtp8lmPOAs2Q98UH4IJ/EvVIt+Krq8XlWG
gsD4KznJWj2vivbfx53JUnr92gYeTf4e4TdO+lBw18mUl10Emt6YzAGOUyzzNzel
VfNRaqf94Sdxalvc4Ntx7/YVDbac16CwkJyj1Kh4cw5kGhlUHBnmZn44QmRxyeYx
oYVrk+NhT/qoh+Oye0wkJ1/Kv8xM8ItrPZysm7+FtGCXlkAOVpTErmOw/nDWeFW0
cGIwJMn5BvTinnNyR51GVI4T+lm9KoupOQXfuw+sOL57Rwi4t2kTIbEkWLTXussR
bG+8DMJhZuf9NIJqFWY5XIklTmk0JuPmIoqnZFP24CH14jKyFnFgnRH9RqsNh2t+
auTnVHqG3xfY8//7MFTfMKEwINxi6mJJcKSjgRg+Sh2+rLFU/LVyV9jgAbvMeoXU
u2XloH9YbKkJI2tcg44djuyQvv1pPpjZI0ulzW8LJUuvqeEGGRs2qLQKgat8V5T5
MtwO4Fj7T3C9DrBeil3HMfG9hSkFl5AiPrV9Cttp0WF4wGuT4MA8MBpYiCUl7mPt
vGxYGdhiK6uLYwZhQemdqiW+b4iBMrQmge8/JmriB9Nyjz/40vDjAZuR7eWvqPi6
eWsPI9+chq2BTXQXAjk++KVz4H8bTt7pbQR2yyE8FEcSTulW4CBgh/4dLGE3A5ME
8/uOOhdjvydfFL3oEwfNraKVjVztb6msZqZO4mbsfPz8g22k5XhKwuEvWINWvAIK
is/ZuUSUsTD0Ob04vVuqykYf6WeaziyiNYDTS0XgEe+Q7Y8sxJIawo5tD7lzmYgL
sUwRznqXrkyprQ+w2bSe5mu1r+K2afX4y68Q/uFNtg4MMZzL58nRAnSlgJMy+Ge9
mB26Z+DTT9ENrd7Ow3heDT8xCf9oXp2//41pQOn+UrQbOmEvmwh7NOEdlg7IVZ63
m0mVfa/RBQL1GQ7pJgHxCgJTq4a/jnrli6lu0/VQCI3VxlvcpgL7F+px+sDLlVIC
7zrc6wukWPYWVFYr1eS0yiH57KJaWi9B4Nk/Z/mtwhwN6fTq5wOjfzn5DDW9Nfu1
CohxkCTDb++Dj0xVTgVugJ/h7e5IAzELLsHnEdFKLcCKFwj3XcoUW9PdA5t2E2KA
KyzvIuhKZKpnpo/pDT4BryFY+4YgF4/AEp8djOYZU7rZipN1oT6WVbF4yvuLY908
fTQO5FV78OEa/GXsZ6JpDFD9F6FsUmdIQTm3066Clp9EYcl+wCS7orN1et9CKWf5
w8IbUMpc8YnfsaVLg6V097bjDNi7mo0xJY7nf8b2eLtgCzQRwc+tO8+ZPzMzhYB0
e1fc2wUz+8ok3PoA+aqXJ9uvqaKhvTBWSyCoTjtmEPIRgs8/tRv3kVYdKiwbXoBS
4saM2kfNWWM4Kz3SFW6lO0VgJJyAOsw//hRUZeCy14eKzP4Qubz/HFKrW8cYLyyx
XrEcL2igrkHuNr5HbwSee2ZP+ZC630LLsKoRfYVfpwhIPOFjBG4Z9KwnQF92l2Ex
rmzEcew03vaGALOauh0+7r2FSruQJ9u9yctOpW+c5NGVkz07+5esdXUoCWKBDKt9
bHRwIeqD/41yp+vABXV9fOfkU1Ck28kse0YFxa7WYvx2FqBoAom7GUkWZzcKdyIw
/zMeEuChV897YKxalvAYdlxebbIYWLBMW2aRKL6IIkrgA6JcnALVj+ZrTQR+8L2U
YYW21NrxA1cJwvhhcWj5hItrZeLBvohQinZCKyKCt+xw1Jx2GA9zRHiq7YuBLqWR
/LutSWc1fR3Sg0lbsvhhNb75g4QTODiAoDTEZ91jcqFohwv2Ir31NE5BePEOnWo8
jBLArVUv2cU0ssEfJ7d9vJBHJZYZ/WaNQv4ywh9VP4xCEG/Xvs0d4pBZK9C2um2O
IfFETxxKWtE0eauPPmrkv9uqeLqxDepmSV9zJEDRVCfx9JnvNZpaMTJc6VX7I/hd
tzmb+b+BfYxC490twGfRWknEPnb64UheBD7sYbdLCu3BFqK8wcRvz9MKpEGUdT26
FW+wvXLnKdGxWreMlaz/u1xr94aLw1ixS9jgE04zDNVyKIKX/E3kBiQFWQhyrwbc
0YakVEJoqq0ixAebxDikn6hN9C+IIfJM+uFoN3n9hgmGEiB4s81xB78++Je4G8v+
OrkwoyPKUMNg0GKezCzS9xUDzAThJFlsch463JicUYPSNTRs6jsaMNWpWK5pghbe
okFm0ueD4sol6nLKnQ/iqnKU5byDA/kUprbbpBlbfR7riLXUxAmoI/S05nB+v6Nm
mqGiVI0O9ZlUQxpl8z+VQ+PRgSQefqUHLleatAa9R2zoqC6iDZH8zdoBdeni5Uv8
apC+d6a0vRSbvjEH+8vwAsh5JzApjb7Ssh15rWae1sm+p5UhOfAWkrOfXeV4R65V
4QDl/9NQIxTx/Yvpfx0BPwN85dbBLSImVIHcporWCocW48vG6axaAWCsxf6cWXUo
ROZ+BL5VZSY8AtuAUM+WQfQ6LO54Tr9KMjCWXPslWpXJRvlQObGiIKx26ICLyhPw
T4ghJNp7RWeYqG5EgBXu6HNaVDZF8XBQ+DOKHweB/8x184vWAOiJKGulRLRkyEwt
CA27r+lE+MNlmyRfGvITTCbPjA8ZJTu3lp5e1Iq4Y9w6oUiH+7xN6Ebrq8j8j6ff
aqfaLkuVR1FBRhzodmevNfls4273qJ1TPknC09o8JiB/pj1Ame8MHQF6f6ryJ6UQ
FJxEAwMChxxWBFOV3cqLWdbocKi12jaj6TkayINWN0/B5txezlEFowVpLJVRxJot
9Y9tBEmsJSOJC2UawIr3Plhl8bKgCwIuWZ3Z1wme7S0RYzcaFfI+dbFHx9f/XMyX
4ODsMH3oMVD9Y+HZAYPBP8LOp4taOGiSmSgo8H3OJy5y6/M3EeNu0bMrmhmjXw1s
Xa4M9INBJbQp9ZYA66GwAoGdjyf+h6w+xQ9v3GlBv54auen9cN4D6ptN5tuGHQ+b
lumzwa8eoGcz4uqWMquPijYo128babNDyAts/o1O3ZioQCjNF097oHJv54min30W
UJXoGTU1+cy0Beu/rU0gEcV6mwGBszuQiSTvqTjO7C1lbAbFqDEB/9ENisRuGMWY
A7cv2vifyJ1QoaSABmhI/ejFmL+ZM6ouYEPym6ESQ1PLMer2Jnm8PPizdE2HWhDW
PkNCr7ysjr7oIZWQzyuFbcvh1jahZxy+ltzJ/sM+0FEkFU5Rpa7+UjPDfqsG9QK+
QGpR8LpeJxps5XzfTBHbQVFqcolKVw480Z+qvU1aECpjn3/5Z2+7HesA82xt/Kzb
u4BaImnQqbqlg5bzcJJU/y5wArTg9CvAxTvytQcizp+unUnfU+1pjPm+1XYl+0nt
4q+JJqwK98enwlbFAWPRk/7lLGPsAoyfP+pynhYl2BEN7F0AHJPEDADkrMaPZe8T
dw46gr6P43/7X5L8+m/WJ/8uvvqOoTL8f0+vHXW4DbC933urbPQGXAcpMw2Iup79
siki8/zPw4qWr7wIfB0rx42rZ0wiAcKI/tzkOOLqW3z8NC28fLobETpmZvvlWJF+
yTcwCm0mpc5KWVfPuvQ089NAbvyNCA5TthXekHd+3OjeQFqeXhXkyti4PHM1kDn6
+qKeZ7FWKvnpZ98bZAIlJUqhh6U/8ZqeexeGRmbU1UTmvCS+Ui5zjba6VESLSD2c
59Fa0Pl1twjcXxmY8DHh4RPPwjUhVN9Gg+hLa/Rym3oj+kkw8GPT9YOPVN7XNrEA
ExH6ijbTMwGfsDCV1Wa9Yqm8J0Y/Zn5WfQVnT+lXy9bTXljvRj8WuKGvQ83WtHUv
9RLTIPrGk8Dpx+jA4rdfvr2vf8Cqtu0qIEQ843qv2RgZTOpvvnVZTT3kx4iC6A4v
RfTbWrwdziv3/CuzLRDclqJZZs+KDHdwOOweR1z7ijuP5Vmjw8mxoll/ZlYNTSfH
0K5yfpACJbKmJ/Fz3B6FN9OdEBANGTz+c+j9INqno33gfyhrNzIEEOrutMaV9Y9N
loJv5EuXKvdfvQc1IhqRYvkAxx2n70CP5wA7GSdwO3XEy6lYh0p3cT/riI8c8XQn
druX5dbe8IX8GQUoYa5gW4pMD8b2PDTtN+ql21dcXkzqImIFnrQl9/uNKtNY20b8
OEKeICd5BoMxtv7cSbvC4hoZi9ld4apiuJYAnu8OyQo+idhpnphzc7kyyaRLxHD9
dlrOjQFOxO1tIWejpSpoATkHZpzIFO8BSvziix0Qo/f1N43CQA4IQEBt/NDXWoOX
kujPF0ggv2oEAhfvdaFkJBGGDd5Cmr3WR6dNLLFjimhPlRoejWS5QHSXypkZLZNT
PreqyD6rEtSKajnbXz4ZzlUHVyGlkFEUqACXIb5E8wyvl6k2QxjiiD4s27OYtGlt
9rv1y+TsNCHE0LgLeUQSIRY2H8IjM7Dzr8X9j67leHLnRIMw3a2kwRxRD2mZsdVd
A/zpHXbYSCH206CbmThdf4XOGzVt3YhpE8Cn2iHr2Fyu8KhG24aHXbVHRb1SBnBA
fERcetm4zHV2aTP2rtIrPl1H+IFzEtinbP/PgZo1Xi3dfXdLY51tzY7BstLst9Mj
R4TEKwQ/oJizgRbs//8SpLPb8l3fPJSm4csxd+HnCiAmglQI29V7ufWGMB9IMK14
IKBUPKloaVkbgg0SMfcW7RyI8DIlDxiBZvjVjNQepoMSqwKaQP55AcGiPnvw+Rl9
Bph32+kYde+wseXNCWzcLA82B/QNf1wNZ/aK5bLXJGs7vJb8BdCMkyADZ6P91lmj
g9y4aQUMtwx8aCENUBbnNhNFwH57bnygOFh/LzoJD/ECEGguUdofA/1i8Pw45BIV
xsoTs9g7vRsjBIrXtFOC7XerAvvgGqPPVefV1gavD19fzIFMXibTuqjdF4mO0W1w
kMey0BIqbEELhsWVOH8sSVdyY+f38ioNapdt9epMD2Lm9B3t7LsRyTVK19mBxCRE
oXi0OmmuPX+39JEj/4t+S+1xoQBbZ+QenxChTMCHT4OXB8cvC7ab7EpnhfcHyFG7
sgrhIGCbAA2gpOfDfkcLk7R8j53+DlXx9f86KQyftajiycAFnFAqjUJ2qPX2BC3u
XnulDyOBrZelAYGyg1KeJbh0i+YVjIgtodQCcR5dIhCuLo/Y5iVZ/tXi6iNYaQ8I
tfpxgEvMbV3SW13rnWCDGLkjtKH9UwAQs/ucA2mpo/hdISRO7go3G4WGs51QdA/y
04jvh1RsR1Fe/Vxszw9Gxvm4zRyP3oHBwrOmNGZWqqV6YVvK+GNKg0wEofCwdgox
FvWJEdrnPYdsttDVKWQxayYR+GDT9NDHHY7oODf0HwAvPLUE2bQuYJ/jnVqeiPbP
sQD+3zgP5QEzyY0y0Apg/4vR2KJUWO6Vd4vjLT5GnANmMF9oluhkw4i2ZHZGTfIB
jywiIx0JnMzexth0XReW7DemVoeaQjPqTdL/G2Y3yuYXEAQsyBtgqSQ8tl6jVZVr
CL2FWMRvlI/hP3J/b0+CCfpcqSz2569JfWD3sYDnF3CO8MDTgjrHiA8oo8TdqIBv
J8UL42JZ8iBoYHjfQd3D43Lg0AeXDk+egDOdL52R/PgybSuh8nOoBfp2CrPUJFoZ
xIA1/1V2r1HPBSrtg1Mar4O3ptU4b5pCGZ1L1UOh/rtNC+5LNthoV2Bm1UkhMAQ2
8Bwa56g2vevH8nbJQeDnwViw/xglQf/i7bh8RcKfxX70tcXKZaqnHYoKaRI04qML
TjQfZ0XGraG0oILzL/Mztd1vt4pQHPpsGvdkBor3Lc/X9OwWzae1GwUA/ZFAuYC5
9zVPl0/wDDgMCp6EQ0LARi7BiUPGTYgVHwOtK1wB56H7H1zVVkbmg5jsSc2Jsk0G
GPnlzkRcf1NRAmgiNtCd1qnLHmkAMcunNwa/qR9bxHxGiSjdnfbc5k7AH4BVmZ9X
U+aMWZUloSei52VJtICOeHM8OoxQQtcBumGlnPdcZ8/xWw1NEVNgR2+BDCQMkM6m
XA4IJJN7AFDa9ixjOwek23wMj3x8dtiweeo7VUjA+gj1+XacPbvxENxAZx+ij+SI
WIjjms720PTS3xNKfjX74LT2rwTSR49qgYco21DJ6k06vbKDLMqlkpWa8lohp9eP
JKwNbvw+5uSxT+q+rtzY84yoS1NNgBA+1EXtqRYpbZwxrwr3t2Mo8rBeuq7srN4I
8E97+Av5XoqzxKjn4w5VdGyS3ZEnw7kj6Cf8OlaN15MYVYDYIW4Oj5XMMVM797/F
mfqBo6HTqW1MooWaYiFDzZBCcUG9hYgU0fe2ku4hhgV1BhmBXa8bY6BdnIpEXpxW
VgwxA4DqV0bc46T9t0/oueae3pXqZ3TfXD2OzDCDNFl5jg706vlhYT3A53tGNM8y
30+UrMlZx+ji6Yq8znxMVjuePSz+sDVl+X3bNK1RQH95EBxCJ7dJDVYwOs9OYMzX
/RSqvlyQyjsmZ+ihA2pRDxWHwNE5Upyv3+xk9yoX8LP6VJ1uInxKa8TQNBg09qzu
gwRm+3ycupw461LWbrzv8nEZEhFl0Jmq9cSYuMFQjXS057hVTSMntoqP7L0l2T4h
fZpY86yEYequt2Ig+AZFcyRMYjarDjA2z8nIo0NcSAJGUrq1+yJ8ciDB0NgQB85h
bV/1Vigd1AbZSbt4c/2ngNaiYIDLdoGMOT4tQknQbrpqBYrXoWVqdkC2PIxRDQiW
gAK4XJHX1KY17AJ6Ixx9vNm3BinoaNa8rCnfkiIRR0quwAB2OUGBsTedAyBNoDDE
mD2azjqI8TpbPA4ePR/159PMAu2Jes8KCsJxaIIlqiWCaDrEO+onPp7Q/gTYh3k1
bzi4nCD4gDGH60JcHyZBribfe9xoqSVRgoDrhuWq7AEn378HfI8kPkzMhmg+lJ6T
rtGkCWTMWOTYYuMFwtbWOcKpJfzEF1JfxG0EPOQAWHegTWnO9OurIVeSGfYrFYvG
GaSExXJtR5RNuRy7ECDjZtbWDZEuizTO0L3l6SHiWeakqOfwORoNvdFo7pO+Thms
KJVQOSLxw9CW8DvIJkqA9HLreed0M3N6TkedM0oRQMM0NnAhd2mf7kQy34TFboBD
+nWNezgZ/sATBFJD6XSqW40ebmpwxkS/D7YlaNxJpc4lvPAWZkb9zjNiuiarEZ0F
21THDTGY+lca/WbSXgqoQkUziunfvPZRwoV6kahKLbgJ/qMTjbPQSOTrHMDJdUPY
g6egrJ4jZexRhJMyVMA/rDBBILdkPyL57niFJIhiaMxlhjtCDDXLWHzm0j4fBKX5
X1QW8AXQCb6QjrFgrJMqEDp8ms0egijEKSor2Po1t4r1RleVICH5IJqk3U/H+VI8
iMPg7RqEMWrTDwPGFVA6MI00PM7jXPFXegxQy6tw6jk915FNopd+boxtiPGUnmpq
1Tb86atUxoHeq5F0LQGzScr3vg60CouuYoN0p+HNW0Chkt7bPSQBA1LPl7LRDiuf
g8Wd8Y1AGdRByWaVXPNeUBw4BHp1CU7c/k8nTig/WXkZhmERM4bkX1IOfMqceG34
1RPNR8gZf9flyLqwlWaZMu3JyhkJ6Ywx6RX2by31ZKtRu22HV/P1hHor866gSJxM
XfldD0nd8v5nUtVZoCIQpRsFOKsa9l77HSLlOUgN/hAUHZjlIeTwN1ArdBHsoezR
raBHMR/bxn0trwU1vgECFDB92a3gneQ7iG6g0GiIc2Ed2VOtFe0KQWX/K6gs11J0
F0P7r3xsc9VZpa6qURT8ttdiRn76+Cnd1fzu/yh00NHi2obhjVtFd7pQbp/CfkQn
PDiSbqS91njOOj7ZwFF7CtdyGjnLHwG6Pmh8tpp+m8chUK9vgDJ7GlbXtJ+emvsY
yOy1Df8bIS0RR0GPatsD+84w6vvgKE2+tyMBLNa0DepxJVWXGfN+pDQoH5wdLo+S
F4txPMgH/Ukro92MdF0Ax7lZIiGrdIKm6VDjhmPGw0HBN2qEEQB1v0Khjj9DR14a
BNLeJ6XhGT06DoB/v3w5WsWEyN7rA0uizJuVc3k5rF8h4bXKcX4J8bP8Q1lsprdb
KCoSp4QyAANehNR/PpGM+TxlTje2YkTEAbxYBrsROaB0VzxkEdorZtq9Nz5gANZ7
7hXYIHhDGiqZ7OpIEJZ99G9WU5Jne1/RfKt9W/yMwJSJyc3zSPrNY4y7rtTlhPNC
3onx8WmaYUoX73294q71UU21CLi4wz4up3EG5FvU6oBkPt2+lB8J8stjZBpcrWM/
uhFiGCq7FBBmmzvibQjsA7QLFe1RFG1dlZAyRrDFT28LHqlZ+2Uxk+funfZEmK5J
P7mhG824I+ZOi/4yyO9Ltm+vZulznDP8OfBbqspoJS+L6eRPDu529+C4wn33zKej
YHIpi9r8HIvkxme+TbOusOA+TABh683oXuRTXJvrw9xqai05ZM8Vv9QUvmyr74uG
7VY0O7FJ8s0fnwb/a4Nl1vRSFvILxBzLukFlzjq/KfwQuWTw3R48cTD3Ct/6mKFL
guub2y4eNvPafas07qsH4r2C8yIeYL94JqMhf5Fh43TgnEXWg111j99ngt+fe7px
s/3rZoRMUjNld3KMZsk1cJzh34wcQLSX2WEy0q74d20H4oVldXtMQwJ6XzCRNO4C
x850sLsOOgdr46GZn42gxNihhvGQ+J6UxP9dpTINSeW7cRo+cl7vQCorfCO9Q0f2
oCfrHEoFkznZPX3y8tvK+ZBIMwNGyjliq1k8gpdgdAr2MOHI5lhz6JKzzFC/BWzL
UwNTEbzeWTjK8KZBBE9v9ABSY/VJb4TUH6qTEZOuASLVIFpIa3UCe9/Wh06a1THb
hW1wTi7OtLG+fNH326ugC1jo79N7iH990P0Khce/S9cu4YAijgD1tPOO2LCMRiKP
QcTw/vDPLIjLZvOfO6w+71CGtZ2PazKSjsYXgkKFHZ4uO6QDmWegN5CB0YdQfhZk
8O4bCv8Za6PtU0gd8dK7SwGL0Sa5XS501frKYt1MahrsMkGDDyK+jmSat17iyHo7
buN/JlcvwrOJeuI47NTMYoXfdjUset6nrJc8MZY4717W85T2KQeSZzZgVqoxA2K3
lxiLnbgPVKVJ7o7ppmNJkVpyEjk5JiMxw9a0VVxy74HFBXXo0aXLmovpy+DcQhx3
9VujQDoQHDe0PBGVHZrTg3RIdkD3uuxrP4367xWlhncA4kHlR/G4aONulcsNPMi2
hxr7crd6edzYCd3o4Bd52FKxR+6bwrx229I7mNXcEbAv+U55G+oFh1lJl5yYaAGn
VQMioqcA71CqyUm1IfnPHyYpRMsTiGOsfL6aojxyVAglVn58uKXA+eRtTzRgwiQy
z1d79fUZlyuEX8rOu/TnP4w6SY1pKTE1svLEfqGeImczzssMMpTq9YPdBxhAgF1A
rv5K5NOz7LHiHjSvIGgwDiXkANkf1rdVbwHyVB8oNMlnUfdH+XNfHh3mvXs1Xx38
5UOE3W4sxNgfOVcckNR2LHIqNWuWY6MsbNb29PCPxroGe0AgD0DDlhw8Y8NfUonO
KIz3w8x/2tzf91NMzeoq3RTeCUT50YKJ14PAttRRYq0VW9RrLus/V3rDHLtqGJXt
HR+FKtlAuXX3vKU02tpnN0eXBG/ObECV5K8BRXR9w4cY6poCCH9Xjcfu5+Bu41YX
TuN+fdLQNmu/02Tm+tAXS1DCiNrTHFBezRkbhwRYLgAaF1ryXQ2jcxc52Lcv3gDN
aIIRNZ8AOA4W1Z35DxSHAP5p3QqjDWfUX6Acwj/bY8iICXUgUkoRdC4mv7/X/FzO
nKvA4G22YZg8iGTYlG7Jrj+2UvsDhYJfhIAulE3MWDw6WuuWrBcyqdr5GdNnMO/v
gwmyfd6UIifcOsGLkAy80d7Bqujw6bqrD37TlJc4QoAHwAP+hNXMns5jfHl9VG/w
I9ZMIfVMkWktDJFQgC9aXNBJk3DlO+7EgqYM1VYPTSjo3o307S8GmMSRYxGkcDUq
ZUOcDcRuu95zovag5icRuYC4pIqhWAD2qCClPxxBa6R1oFj7a6Mb3oT2SNgNpsH8
3UzTmK7MxbQA4Y0eACQD8CVZGxobLVS/CxLTwkI//oUW9GPQJRt0teHW01jjWrod
KpLAnILBxIiKqmtb/hrqW1PWLetWH628vE5Fx/YzgXY8Lxf/BzvpYqIXCR4Q8EV6
u3G3IoC6TA3Gbm57b8ZZhpTwuOTmPWR5wDA0Uz4gTRhsL2G+r4uL4k4Tvztwlv1O
MR5wqbBnLB7xS0r669/6HKkmd3oVwPU4PgObX9xx7v3YTcOxqtamcAGzdORulDHk
d+nhqDdPDYDQcmI0eQnSVzmst8AugOH7ARnYF5JSUb12AMHTL3G6ZYf8ED4p2xkk
jvF060FbYOR2pSuT8tFOzFDfqx0V8rs2q+aAvHNQbylf4l9TwjFfZYVFmyaHj81e
OE65cuOc5XOAd0mqTeLzkP1TzMOp8+GFc1ul68udqs2IVJ7kEphnhN7eC6cSBZ9g
TFzZm07nB8EBrJToFtGNFoidck8wZIGaywiMsZzW6sC3DdO2IFOAdQZspnAtCAp7
HJ8Fk1U18WIrrA19iNR/elqqpwcQOXPZsjKUG5lPK38vye6IZH/d/vkVC6moifGX
jOKpliGewF8/Dv1HOnknH0xN5lQfB86pA+BQREcyGfFlHDblyMXlR7Homw0HRCQ5
zbJX/mpXSM1uC4RHNPPCqTPZ1H3NHD8pL7JRMj/IeNAaWElffnq1ltARt0q5cE5c
60G8f2kvfPjMJRnLeZAg5rA0Q0U77YRE37Mqx4NQZwKkC08brm6N/WSgb8bzQQyf
OpZp2Z2lkp6jhhM4amQkoCKcsG2ioXk+533YHatk8592s1xqvVUJ6cvz+DzxH+ON
HiTIJZPLDOEtua0wUPERhiHuOg1z/xyTC9t1k0Tiyhv/3tSSAszIlMM/sU/RlXE7
2OhO+PKMap3GgRG2upXhH4+12TcL41dmaHHpzFIqoUzFuOMGU2h+gzjIZd5YQphp
9gAf6XqHMiqlRRixYbdB9eP0B8qVp0rlagOmq/h1kehE1lMEOSstK46QnRZ/f/SS
f23fsla3PphtqIl/ILmLwTaqMHYeCp94Xlc8gqMjaEE6eGrmSAyi4ROjIyOL3wXL
5AH3hOcAIfxzmEBcs/z5VZqFfPtgS3RT4gDVlw5VUHRcsTXtZNzFUBIUUx7ctWT/
CZYEqt+chgnM6vbGIkzJLDN/+RcwcENGED528yj7pFsDs3AfZj23RI8DOw7PJLQe
TVcnutj2XnMAb/GOV36FMY4aJI366WGihsSXytLx3gleG55L0aIClkjuSdrjM4fw
Q6uUJ/xoYPpvIZ46dkgbabDEjytwuMLubdW9LaAT5it6h2aDB/j4cW0dAM3zhWiz
Co2LDYBcNbJQVrvmJ4Nm282m3IpuXWNEZ1NOENFX55UF1OYdA1ZK2WsJlXxNyBuQ
1muaPpwHUijE7QmSVglLw/DSwEcCN0IH8nCx6BLix3ky85BrAVWO8Eb3WqflYUGs
EuiQQO6ecTkRt1qfQ+VT5n9WLHfbg78INSirll3FZ0BGFjDlf+0jHmGIqIB4U3vk
FDiKpUt9bqNLaJuMOpyyrwa8NOIeEAd6aSUwvbP/Wg/wZM61lYG9HDcIx4/6eTSZ
TetSYvKUbnUgqI3StAmgf5cFLxXfGH9jx9FzPlWt0bwm8mRb1JOSQW5Kb29nvfBd
w/zrfOoIUa9NtEPH+w5LQuiisF3Q5vJl+Y7kZ8cSKHlm06PPOXURI2MZQ/ZCXMlm
ud58pIwWSn7P2i05pQSaDYUCwzzs9AY0iHeRKimjvavJcXnpKplFmGHtdDCO8uO+
YtjkxlcUOxobPKEkfWlJvaDLAP5pL/tLXHOe1YZQUWo53ZlC83iXOzYza+m3AxZU
fpR3mT3rSuBYTXdiBvzJ0U2d95ZWamjtWVRb8V2T5aI3Q+6s8byCU5J9ARG4UsjJ
ps15GLMdTAecqcLAcigCcpaawSbSh+WMigjeZTyshqYJWQA6VG7E90ylFK2aTcT5
87UucTR/O8AZlCEyXcEUw2w4F/3aDBibW+88JKvWSA4tVin5SgXZBK11/e4rwEn3
se4RGIiTBugHQC6QiCmlPSAKbqpbY8apRWZ+Gx9WKdycHIHR3UbSpKUd4suO6ixd
CLOn/STagsr05zryKiMuBudgqcYvNEvGbjxIvFQGQNK+BLOxlkXEqEF6JPY52JAm
Qe5G/qyraDUnNKl54jcShv5+fwhgMti4SdjYHW3jSld3wMMLE6CzlqlLz9uh153B
qaxmvSh4YMHvM2IWcBELFH30Bgn2l1OVdXzmEFHlvUFTjxgYWRhIxP4MusZkZhzN
ZDiWioTUUi2uAmdbkiJ1llIwIDmfn1Ws2WZXzVqP8TgXxr3rY0W9H4no//mlR9WH
aGjA2Yir5xp4JPHaNx1MUA7dH8DFHlZVrCpFOn20zR08b/zQ/8mAlPevG7cC5DAS
oxgchDuAaTmieCLOrEDg4I4dfQqmkI4NUaCz3PX6eCr4JstPdTQwuC/5OmSvoKeC
cuu6UNOIIj+oWW6E9JsF3JyUWACSl4BQlLEDoazk0uH551G0+N1+e70voJaQf6l7
QvZVXw7Hx3N9KYVmbWlAep5JalOruGy5AAq/o7QW8tRyAwVrbx8co2QU41N83Ofd
FXxhRqz8RogaCICz10hs/+Rx5NKBsBm/b8xxlNrqQaU6AygLvhLGkNrOd1QYp94Y
O/umyS50omwlb5i0eG9wBET4A59nP25yRGeQKJn0ade2gCLIdBRB+CyUd5s5eZfa
/qprBIwRuSFscO8uwPoW2kCyA7UEvnjHiZk1Nh5EY7PJp50ie3i8mnLQv/QaMiEc
5SLrnvMcay0KLQsD6yxacToGH9nezEDMiU5vsOtPmw36ZHDiwA8dSaIORbU1eG1Y
ETB3xY6Oxm9i7zovMNnO0VeeTi9PhpqGQe+4a6LJsX6J+XgQM2+wwJJ+5FlYq4IJ
Apm0LHruuOThcimJ0ZoVsj1BfhBCrYA16KePeBfpJ/MnSxNYg4fnGotOykYkyV1K
5gEs14GPE/DYTY+6e56X/+aLeBp0D0CtosArWBinChWW20iwH0LzyiEIUuHh2Pq2
daxNLyX6FogluJJNL8Se4P09bfV95SrkUAFgySWtQDfZM0e2rWTm4dX76CJ25m3P
S5Mu2sjDEo0wGFFoXXSsrrwCXLWd10Gk9XDLyv6Z/PWGr7tKsMIR43nAW77v2lIm
GO1P5nZCq7gtGexI1cRA96JK7JsYu3cXzzhIKSh7Qu7XWyBl8pip2hmcRQ96/9v3
xtZgkbcB4oEfiJPTxdwjcbsqEn/OYRmdo/T/Z9XZLyfBZJxNh77CepZA/WPP+HR8
Vzl0BWgbUViIouqU2BI0U1WEgHJxYNkoyB8vos/slK3J3Q81NwnKJLjWLwZt49n+
HQ436MU7YJdx1BYGSPU6qjYwi/VWRyL+6IOfNq7ccvl3JZuDZs/bLp/AT+L0wiPH
GishV43xqqF83DZ4KQC/KaKXwq4avrREGw3/NPApAYlH0+KD6/bT8+AFuc/2SQsK
1UIFa1bPO0Zb/Hh1yNaRZTe63mZFGnEOKFYfl6CYM3tpzL9IJ8mh5h+2f/GM97GZ
QoqAdkIJ8Pq+jY1cMb73Z9U8IvIkt1jSFrt2bkGLRwhl3SpT8G4OmcpW42vykR9i
NTBLZfvtLML5brOmOCtuay2qct4AFDgmUafyNF0jxgXdRKW6rZhg32+txBAIs4EY
KGt/EqEyphWuN7yxKyhnGKMlZSXRNI1gJlCUMdxmTeIUklNBixMA6Fjw+Uzuuh7y
z8mGP5o09XjqQQ7k3kH0qsHpQlIrlDze+IiIKj7w1iZ1G/MnP1R3zWV8AcR5hxS9
aJThg80DF5mFFahZtXeneaYRzkiLtEWNyVpuZG30Jg0SpBlvboon0ut43G4VI2nV
i0UCre36NS0AT9Z8Z+UzUOtl9ZeSDv8RATyBlt1Hau0QElVcp0/7e908LcyrTk+B
WB3K7CtmiXESee2Kv+vKj16UNUs4c7cMqAlleXU7tgPWg20hN9bdhVSpZQqtMeS5
iV5B7TrXdW7xQzImnUqH4tBxT/vUeBmFfSA1YAdFaH+73/aOGtJ4GrSDr/6298lt
QIojREH4s5B89J2B1VwOoPg3K2LpUsA1nx9LD+1WMhwbjCl40BAv7gzK9Nx4Pm2k
AYY4DKKN9Q15sgWOPQ0vgQtGSib8Np0xpxK2Bmh4CpngFKc10ljIXX65HzawtVzp
gRDz403gkrMglxFUt+2LnI19EQcVAYxMPlhspj4QQ/ThcqwC90RYZ0PbSoUih4yB
u3kuOlHvWZB5uhHSElOxBTGaVTqadjQf/tzMfo0sEXrOjihabvrAOdDO+l2ahcDG
0KSd3RKABvjeudxkM2juKPhGX+shMvNb6xI4jI1070yHyCTf3CMF345n1jze2EtE
9P+ehJZrXWThI6F9HzyO0bpUvdTXyELoRVCI8PCb5zF0pogpLsJmuvzElcN3U8P4
eRLcOonKL58nkYqw2QCDh9sCqXNmAN6vb/S8a0f/LlSokVNI19UqsjxmA9SXXZ7H
eg3TUvEPh8l8Of7Wo6moyHHba+RO1KBU+WyKIB6GNc9MWuPXbtd8AHhUhHrg/QyU
8w3oPNB9eNUhuLNtR0yL4mWXGMhAsqMPqk/p68tOuTWcH+iBkERORjgl8zCBmVDu
oBG1X7kIVnoI495FnUdfU2d161ZCSRq8l8B88OK0yN1Gtvi2FR/3iKpOKxvLs9cZ
Gu7MgXwkXKYT18QdcSKL3uhi5ywkxsSG6rx6jeKN48rMxJGOcBSljsWLiQ8oNbkZ
NDu5Q3/m+JaTWiC6XhVg49AANpHz2/8QpuXM8UvwNjbPTG63QZY6mCnRxcaC989M
wgBi4aX5YnDrV8G0JUS5YC1tR3IfBhHDbAEB/aXpIebtk4c7YCs0ftGxWioKSeJr
9b4Skxj4cXyFS7Tx0vuBzw1hJL/n95BoyfsLrbd9pLFoTtuDj+NxWblO7A560vSU
EvQ13RvkOdcCQjR6SXbawXPEk53nI90PkXrgqNWCkeNLLOgEnBH/HV1oSKU+6lIW
SB3dsMmPYlUIT3veCy62plO3XFaW2R5+ZsDGf2o2P2bs5joHsKvhvrkNlHUmjY6q
sFuG6BKbe1KoS2yh8wJSTbLRULN1JTnml4QDVBJ62uAm5MnE9tbX9IIiAHABDNkv
K1Qks88YUdPlkjyrCIpOPPUQtupHPrEHyZBVaQ1xEHNYB9PH/KGZckWzJpJQP/e0
K8uWRUEoqA52kxEyVjdzeyZBuGgyEyju7ElI1NDlnhZMTSKFlrcAvXir/poj65/4
8KasvPNkwxZSy0sE255kyfC0ohgLvyPVl342B6YEBO+4KmN0hKj4EhL0RGWbkXTo
iGL4BZ7QXJxnG+cXQ4FkvgurURtstyKKI6v95hXaPOcFs+joXvnkRT/DFH+uld2e
hSei2/9pIW10o09XU+4t4rdEUdD3trvnYyA0warWturpPQTezWjJigufOsr9ZkfG
L7kcqur3nI/0Gj28ISq0DO94l4/9WU+aT1GJPaa4kj5xXM92VRTTf3HCCBJjzing
ynKtxgReCRFrhivY4N0F0PhmYDGu9sa5+4fe5Z4vLmLYlsEFUzixUB22U8aLjwHr
SFK/gKfLrgzhe/45+SiE0e2jOLKqBfbo12BWB0V2wtq1Pw6lXSz8yKcEwIG/Qtis
wSwRJg/jsV4nFb/PK8Fgf+U9TeDpJqgvpzU96lcTRzaeopvWvO2m6NEAdME2VteN
SEPiNylcWUSq2FnZRRJK55i+wMAF9AI5K32pA6zAG+ZwYREwzPTPh5l++2X9lKfJ
30sXxOU3Too6P02FR345PVcHbaLHB+eKKA76pzJFj15m8MtUma8U+R3MhR6vtHLi
pxGfZfhGWZLm/X56XkrRuIeCISbA93m6itO87BCzxybCotY97PJBCdXYUwxJNRkX
0qk8lt1LxAOtGDbHcezQVpxj5xC1+aqR1ZEw3ZhoRvBYcKGQGBEsUbNpKnHiIIa6
UL8BW6xdbGZsYdw3GXm7k319QndF13INqLD9TQ/CscHQXtvx0j/t7sxP4VkgNqtn
yEaQpFw+agJoTL6sEW0FycIiO9b+b7MIk/QKAmPIacCb1PqviEEJlX9HV7wpHuil
3cTRdKGkxmSRpamXPMaYL4ETk+8MlR4TMGu2upzpgz+d3Mgcf00NxKM6Tby9sonJ
DvH/rmE1O7JxTrT09aPMbVsMK+SoeUH4g2GZC6dh7SKIUrEdwveGNUBKWmT6ajat
Rtp/I2sCTf3Eprx1cJ4oTItRTHKEX9E1B06FV8vc4nNTTMLcWiaGqRTWV3V5hB1Z
NuSKKfCbL86U9fohJSUKJtJK07uGzUdyjN8vvcyo5To0Y9opdzKS4Eno1m2T3O/H
lwn8I8cTw/w/oRruRgqBnjOlktRrt1dO4YtfBK3vwTNGJgwwi/Pbql+cXl23ZSP1
tOqwMXXK6pyJQuzyhBrd3NVt0i3QXf4o5drXcOi9CXB+YZncJEu0txvs9oOzv0Qs
+MqVCKI5s4OzHsmyOUE80SYwtkbwKtLpw3FkBwIoWQT8EiSRh7PS1xs2xwnEPWhs
EdN9BaP82OGCcu0fEgpQO+yheiI1U8oqLpqasG0unWKcy9wzphV1OUJPJqW9u1rj
7QNX75PYun+5hZD9WZWxOOG34bzIKOyLHfAqilgtMWXrGR9sXLEjb+VIfba0oB3q
uaplY2ScZb/gKMnrxIjaos+EaxTm6NlzdLwFn60RhL+A2ujqXLcdofBUZaIHncqn
cgj7h89eiedJ32F+weNkfMS9M3MtleFjqTEYyQmWxy/06nTABJRM2JceIKz5Iq/U
5QPG6sH2K0uLkrRw+N/XuZRgB3vlKtg9sc3z6QJWjyl3EPZelgsJdZK9cE07XnvY
UaRJeRKNlY+luBU5u0QxIGjbKDmUZPRPOG7yL4fiGzkd8OWKkroF4WSFw1B4LW3N
GAMwkytIVQTNFNS5gb6ErdycOPQPq56E/DdBpwUMu/tXZJwL2fRMvJWO5d/RW2vb
4yYA3CbdkQ/eEmex63/54QS+OJN5/sMztAQvBqYGqY555ctZdTWvOXMQzTFy44vJ
2x0p8Ovd/hEDe28YJzjo1V80xCIAVkI4ZGtHlokhX1nF502hFchB+5vzeQcocBh4
ZpotCpdsU80F7dfnVuQUlmeLG2GxAtZf6Xs70f9nUNoOy4746StprpyI6QEPgeYb
flg2TSTnxBYkcqBlTimBArQWOiDd/00wDBcyIWXU36vkQW/5rotBGr3pp8LqUzTA
bVwli0j99od7/AR43GbzjdbnakqJhfygZEGf88VZ1nrgM2qsB0GWRy0nIqBqjXxC
XiBMz2/oFZR6gSWJPJM5FhoWTj3vqJSBPsjo/cxNNQ2YAjGl+d7RmJHlXqLaHe8P
uf7W3Mai+q1Zu19rZo3nyFeTEZ/c5aSkEKa6I2LvCxsHBMuGreX9tRwem1ihwEnV
+z975KaFsSYrBSbHspnhwkSTgH8Folrn6vxbWVjXG35lEXoarqQCD3V63TKotUxX
BiGoqmu9IPPI4XK4cmXZGR/WHBiBXADTIv2n5uQKKe4GGBOkaTeZtRY52n6Z/Ena
HoNSW9LjK4ClBMFt/B36c044sAd7Kl5cDbB6Fcb4mGW0wIQngpuI5wYrwH/f2Hqu
W+oyvogXHCmKKXl/oi2vNiOxJd+D/fDIrQoJjGqSJOQiueMZtue6sqE6WXQ9V3UW
k10UZJbzllcByN9QTSziYf/UwZghE36ufs6gYrO4dik5nkS/O93KZ5rNJ/maXVvE
G5SLsSAkymBmz8+8iSGBw4Cm5cmrbvP2FxyMeA/YJREdK4LzjiRI2pknr+j+GGXP
qddke4fAZ6u7ucyKRB5sYlhJn/C3QnnnrMCsHa3l8odjseXrCfqoF2e9+ZnxX7Ha
D35fIbQPNMcdhx4bugjFI9n2VMxYws/roidV+lqrs2MWtrr09KcSpJAiaeybowSC
JuHS9vcyN1wmuoPhHOixmic2+9qUPJpiW0rcdU5zhJ2xUtTbIh/gVFd0jRZ0xFI4
dZkVspqY0hM6A1e70uMh0mulSrzfAKQtcLxVBwkz5BZV54XjIfGP0+x118lrz7zv
39h29doSqZ9UnbOQx1PuGJR/KULILeG8VzxHKadybo4OgqGVKV51F3aUUMtEmENw
T1mOXSsJdHPfcCL0OSmYDgRxr4jFATX4wLmFmFL36ejhutg/Q9R9s6lvJbbfTGCq
2cJ9dn3dlQP4eJfdEYSMuVhzjW4GxXD9K6ZMxjUS/e4iwtVhtnGOZCHVfy+LJ5L8
yeN3491E1nZ07lkc8Pm2zPNVY3tqoOaJ055ys0n/G9l4Yl3r6ZwnNj7sV72ThBnX
sU27EUAAlvMBeA9MGPZWpYQhEeonMWSMHVQ/EVnbV4EpFTtWWVGiJ283mEXO7N22
jykqkw0xk4+RKfiMhV+is4EXRZRhJdlmcsI20JPT+b4g8oecV1ldK3QfOyrnFAia
8WX5BMdOggt+mLVbL2Twsaz5pu+GntyThEWZ5N1i2wsvE8fmEnurOLy3dT3MY+s1
0jdLLniuadimUO3Gna4DUQlCsgLgpDpijPRhDLRxQyK45w3E0u0358HZuVNsoVZO
QLfilqPy68Qh6WjSUAumyPPcQyLay0xpmUPzmHHqaNQzZCHwXi9fjWvkt6GzMV9B
fNph4ZplBpa/ha7KdDXH2Br4wlIhg2xKcIyw63sysl8sJe9GpkgKainCI20BJsiU
gf8oKnURaTCnmM/nBxEtZONRPKTTbD2/qyI0fdgZf5yzamHFOnjYGPnK8IqXaoEH
+C5zwIyvw2wLwKJGbj0LjzSGMvh+vgzhQ+MFC1ZocwRRG/JOMsl+bVUsyc2j96Ki
HBi33glL2YE/Ps4TtJ5/3DB8OjN3Xb35VgZO+PFYDsilL73LVw9G7JoC9DUdWaLc
CqTluueQ/lmyUIyWL6zGct/spwEYmDT14AfKMHBO0fZKPy48bTGfZhauRxdakska
n7KflICO53wiBhp3YdTfGTqI3nSOC9h6CvfAfZZ8lLldtVY0R4EcCI1ctJv7tw2I
TjZ40og63hdQE06wDyimhjeB0gngrxkR7IX26wIsntcdi+0Tp5ZE9t7KOkhOZjgn
UXK4YNquKzrhRRXYL0CvTy/rC1kicEOFXIlDFC+PwTnjBhBI5OC10EmPqqyhjYML
MKO56PtnSQ8MkcOYWPRtnU/Gb5QmVRtKJhwUzqAqU0RxAL9lFHJuaWVn6eEi4s7O
UTGpsW7tY38s93KhXTUQw2/bV/gH8wPi/daWIp9jidmRVf1fkx1I2J+KP8L8mbHZ
IllZQ9XW/+p2n0FWDbILyQmCdKNMwkNT+K9IyfQcefFMTCJkkdtcnCotMgXeeCf2
9rCtwpun+Rm0G27c2PX+DOXsSarVPvTwLu6xw7Cyd7VUxSovSrc7hrc2NHdwKkks
1IHgDZ/Uot+lYL6SCsqiTFeShsLjncBIs++OSl904Q7T3ATJzZeJlTnST7ocL/M3
908VUJYpApJCFY5cDqWKXQUhWocL1EV+Vz6zq2zWS45w1xIHbO3QwH6AL0V3eV5X
tamlzNeY8O0YoLyB6NhLRQg965QnjBPmjJu2dPXIN4ZLnUvhyzLv5qx/hsKKdnjB
EbZgm+tDOenCzl6iR5Tc0lP7ru3fyT3kgfePcleH4WDlG0HPDJx7Rz7bRFSHQ+yb
EmWtMV17qpPeYLWBa2nsKgad89hl2XIqdAl6SRSnAypWzOf+nz26pGYhxYtUwfa7
e5g5LFepNbCSgqjiSyr/7NFJHRM5Atz+vR38bD+bs6rOs80CW2DBBka4o1N0UjU6
ZjiC+IN7P1q4y5+6Npx47oJ/r6WLijvU/ZATZjYgu4CQxiJPZaSKjnTylMx27YtV
AIDk1ohrBqYK59/qX4n4lC5WWERgy5sutUl06gytn3P3zMt5Oe5ISDhoWrENhV6D
7ps5L1OClf9BiXJkX5N0XycKHynBjYOgS3Ob/3y2fSRYl2+9yGaiAh/BzH72kLpw
FvNB+uuOhR8UDYXTq6nBsgJlKa918uaIMKv+JekjND310KS3SVOfLg8tiisNei7/
t0jrsulV1nPnXnM5/9OjLZCN8FStkx1Uh6aZQCpM5tlqQsOU5vfsvX6pLMwcNZr+
cvOiLnNTHJuYr9lCzglM/cJqzXlKt23k23dG9DB+lYgijbKEfnv0/refLhSxkh2k
TBcM24eKQA2pRnl9YSnH2pHoAqUz3g3THk36kSrE6+Zm5mrlLhlvt2IDe2vVr2ze
fnnNq/tMUODBWPEQjDNki8BKudh5TCnSVwfZEYym2LTkaIREsElgf/C6U47S3mEi
5n07eqHsHZ3w89OaP8B6Li/TubkLStOFFFqrunBpwyiLzFepu7QzFIKuKuB3L/Lw
DHo3gcSMdB3alKrH0z5XMvIr/Rs89m3WY+OHMemJFFtm0eij6GZo5EFs/gEEO4ED
IbP4D6qvBi7HgdQLtnENjZ+CeYxzYkwYCIfcg7mE76Uq49UJqU1moxp0X15TzTS9
JvvU+tL3PaWWMvZpNZYTv7+9irvlgCVHyrHSKybutrI1rOalLjSGcmqSgY1Ql0jv
A2fR8YR0Y/kF8xY4uawnPal87ktoAlU9kRfwEkVUWak3PUWybFG8O5PykbKhdOwy
+j9egmNqSHQNIYs9Ke5mLIawz9Kqrw2+hCOnmUSxnZVlcDCcar9tZVPm80o26YVC
XJebZz5r/fpWT1s9kXYweHWTDf8xy/icrv7Y9DZbTAv32lKRr/1oGo/xgXF4dTld
EWPSOCL/ihchPnWHu27mXkx9jRPKD3M3M9N+rRV7bytYWCkxTJ6PR0IFB5SA7arr
DOzSmXn3aSffkEbN3f+2wns+RFJpI8AIUg6oA+Hflp3dFzuJGoWO6Cz4Ybnl+Kc4
TpK5q7ukX7mBR90lTlmDONMoMCykaOuqXVXXE8XYB2BXSUD272FBgB8EwAHcX2PC
/DxpF0MnQ/+PxpydivKwfB7fMFGstC0mwgTrSOQ56/mkX7PkZDU7ZfQIpJ44nEuM
A2Q9p90jN7odhMN2HOU+rC4desGD0ny2DC4qEi84Qgt/dC3N1jqhWxXFOVPAEkQx
NroqNK7BNtNkgO9R406+uSa25LMGS/H0YyGKzbtGfJiiqsbTDrW+LgwVZe9/HS1l
K9gSwKLZ1jEj5Z+pHtLgzV1sgCYxdlmIVQUKEPX/2QADg7SPUZAG7eLNe5EDw/Vn
aZW6tKF6r2luX+RASYD9c1A/taVNTa39ErmfPi1YgRyjBPe1bl34e7vzcj+FgHgU
gLrB0Kv87UvA9/2fMQpuDUQTU6g1cuWVHx/zdZbbzpPx5e8QQ2C8JGf5vTFjRzK3
v3u5NHOB+t0SYeasUCiV0gCRMDkeaZtUXhLySXN5hE+gglJTPPAN2wHPZP26oOcA
8CEG/3qWgyfygJNfcayZlQA6LHrzUhQxqxZV6K0BE/I9mXZOXekgp/K9ADxmBLUa
/cO9l4LgCE3vkLilm3pWAEL9mTHA4g+mxIqCoMBdS6NIyce9oENxeCWLTIOdD72B
97igxlR+8mEfmTdu7PKKumodCjDZ7ESlehpOQ/uaGTtrQYn22I4G11MHkCrHhmlj
Ty1vnporoQd7BBdp70AZQBh+15BQR793CVOt2Wr7FLsahR4z6RtLQ3j1UZKWCFwu
k6g9e0teHIZGOYbPszSzXj6l+qEOFaWsUoqovkjDWND6XtrL8TSL8KoVUZY12t97
B5IAfAAmGB+s4canr48qUXTrQXz+6DbtQNpfIiC19NlW8J6P+kcdUkpLyS+yCnqm
OSF8zDF8KrWrePzUY0l8UVG43ReYuAaAQnhxst7mN4jOA0+mnMUTwn1ztgEL6xsS
IASwLZxYn5N+fhnvrlkxPq7WoMd8NAv11is1Xnz0d1z2o8vsKq0hg9yLnOVVXNzm
HsokQEiMokmh3OS9lovth36eDDrlNsEu4pmWsHeIwEKmfT3dyxuuflHpl9HbJjHN
m2eJLC0AGVbif8dTkX1zTmD/5ZJJkEPNPQxvGGCYeXqwc3+i8dTlk77tvFHgYHz4
VkHH5yNVKyDyXCiWyaE/jA5/lWufX46FuM5ZQcmosa11LI6RCRb5jWT+qa3abNFH
Ey1zwtS6tq24VMjQ8jZYnQrEyDkjRjWbs4opwolmvGZfFOXaGnYgBN38GIUV9rQm
IGgwqyac9lSFw26HTN/XSdyIiAZ++ftmzgQBcVdqq+M6zz8fAJWL3aDvxx5NHLuo
azwHljsQ12a7HaXRWP3rTVNSDRQP+xEPnpV5zAyxvXLb5XuV78aUgrw5T6vmlLFo
z3RH5ADo3xhDS+zR0VeO/0P1doVD4W+Mo/ISJg53hiLs5aiu5DJEl4uyPfVPav77
H/dI7l+kIRY5RKkWuM+EvJqg3Zuze87hguuzYan8b/ANFD+yoQdeyWIDIHXe+BGR
Ub+gGU0vYKA/0BjXR+lrh9tpT7lBwiwdSR9Xj7kAFx7fjwdP6K7UA0uytd3bC9NO
sJWv7UI3pJ4PYTmxIKAPMDgwC2vR7ctmppSR3n17Jd8R9k4QkofvnlL4ChK34MZ4
hRRU++e3Nl0mk8LQl9kuF6TJwZotaC6p9HM24+cnrgAHczbXzHHgFnlLHslIpgGa
3g20EaMaguPaO+Hs/Xja5gsfS2jL1Mx+RC1I/vn2LzdtQUe7GvsgDSzygx6SKy/D
6F4qS8IEkHRoLEHF4VzKso2qbSq9NXqEtxUQVEgU6yx22C+rAvWIwkeVh0GPMwsK
EDftbtCppU0hP7BKQU6Nqpdw4JqxTZ8I+mnCs+tdInsWoPdq4uHybIVmHdWBf2lM
yLp0KFJtG+vNTXepZ51tS7PUi3EREKT5i0XMNgxk9l85YSN8Ehw9GjHsN2FPazyT
GGOjQycYr6ER52/01ew7yD8Ob4At3yE7JxodKp5TgB9AwNwNmKD7s7MBka6rzicr
CxWwFkt0GSFcIZ5nITaY9fc+FvzXCFJA8wxTlb4stJ6mk6gYKIG2l7aYdhlPsWgs
4AqTA+p1gJO21u8+LPLpNyMSWBJfvV1cr0HgS6bkcFTBfXlNkO8Ifer55DwfpXEU
6xFKFe4Rirr8Evfx5vWxwz3mIvB+ixrycqmokGyvwPJ57j2l7H2lw4tLByPyk5mz
ZXIinKQErc7ICXG+at5iPaZ23qFS7HXycQBNcyF6+HiR6lwgj5hAzNwKtQqooJE9
x9HvmK6g1PY6qGaRa3actCZvtDtFRUdMFz80Bv7TO3wNTl0jn3F8fd0hwH8NMm6C
Xq8ja85QfUkDeeXHk97Zpu4bTSDIE9KqzLw/2LKBaltHjwIHLoQWWby7hKIk+SBv
dqQf0w9uTUPxk3loRo9D6tAsillHIn9juJ13G9TxUev0y1ZJ0B+wUB38vlN28Fcl
/S7T/rx5TyWkusdaN/BcOgKh3hOjQsTqNJa2ynhVP4e6YGn3kae16khwC1JvnCvg
Z0nvaSnwjx/GIwJQA5Z6q2g+sPl87I3VYBWtbRZdQJvPLs8igqG4bqkuvoX5Av63
B+3LFqdWMrqTxgFC3nuCyn9wZqn8F3FH3g6j4BRPNHfOfH6dj8LlFlqPAOJgcxUX
bpGFqQdwa/fyYVeNQuV+eD2m3n1wY2rU3OWQQ3RGwz2nf6qbaw3/7Klr5T+Xdzhk
mRSojWtSKTeHzDgzgaCHUbKcS5RSgN/iV9mTpFPJwcOh9o8oJ+dpkpO5GGIczgCj
vErTiNvt+rZ1ofXL2GAPf7qvs9zJ02K4LmmdAT7ekuBNwUp6wPDAN9G1FVCHMxtZ
sUhBu57ms3DklXQNxoCgvmWvuN9kYu1UGxfk5uysRTyyJz6YmP1xPJ8dMqB+ZQry
Tf06Dr0HLwe/q41GqgGDVvR7Qj4+qFdB3V0d96DV7HNjGGRhn5x42+iAJ6kZpsDC
2/aePSKZX+fbQMpsoa5FMJBsAIphcDTtj2gkG1wQb7sQcdct3FKRaGzbZeHEIcZV
yVNHfUP7ofWM73azFTxkciWcJtPYDOGXrDO3GDoN5Lh7LWu70PbCqKxo6KQVGfAI
ZcLavVvqjdCrhdBBIzerTtKaYNfps/C76TFDsV901ExA7Abkjo3hczKosSfCopB3
w2klh8BxzJAzQr8efnT68rYqm1dDEX25jslfb804zoSfGS8FIgBqdM5S7Da9NXkg
FQt9TYu+fQUaD5yv9A3gVDtthfI9yaJvF24g+ZuEBE97XaUrpCPFup7OzIlptRX7
icSv9ydGX7XWomwseMeaKn0SWvbtbr/ZHImyMqEiJJvCSkqsd8tU8BM12X4Tbkq+
A1Pw6gqQ2nKb85WDTFq1cUTLI7AlQuq9Zm2TsQgg040bLXewdiZIFV3aVe68BOfE
+jubPtfMKf5Ozf3Hul0k+wtDtFq4ow4GtgUqrtUKZrtp3dXSrEfLro/HR/5AaP6f
UQTFwgnEYwzfF1/NSzvdab4H2Uf/NgQUvFewKiFrhRSk7dtDUhTqMWCc/kBmDD9o
1xwoioblZZl3Zo/qXefJ2c0Ewmx+r8lVEIlyUmK9FXL0b8DXs2nacvVqB1fJr8VV
4uMhbnrp/EuduTCCfthPYq+JWvWGdksnYeZ9zYYcOl3sH8pxtcEJ3vb5uRBjIbFH
98MKCG4EhNdYCaj9I9M0/fzTEdlmI52B6BT4AwJYBcM7E5F82/22hoEtcpQgu1rt
dP+ergYb3FDBdgVBHJDM4IC5ryHofx8Zpdfaz0j4CZW0t7Q0R39X4S3UyNYqgbd4
AJucACDYuUNAYSgbirG23mism60F8yk0zE4l6VQvgyNcVGr0GCbbVWSBdwzkUyut
0fugTHfgb/3SQ/JDDK754WYk3G09BTYYoXAjnlnIf6z8Te/9IeWaoCPXc6mLncZN
86TI5c9d6ASPubMItatZPjXIXYKFBpwqneRKPbnJDjczzqfbgaDSllXPNcFSJt0c
/RuDenwIX4Qnt32EmMMILaZ4mjD3ptO7LNfOG9YkYmcHZ/eH0ue0aP8sSkRzW8xn
RElwdmjayZ4MFGxa6O571pqHqq0RPUX8od4WfQnHWw1I4IwwHY547F/Y1pBtk2OE
rXaWUWfIi3V5UowafH4XjJwzhFRKq2hMEhfOmRgIQ+PXiiMLIoFXe6wStzLRGjc2
+HPFEagEY4IfEa+iUCWT2I8WRST22erSMkG7Ics1HvsZ4HZawNx4HbuIfariad2T
mCMMiMbGpzM3dQKrEMlljc2P+fJlm/+8NyFGEDxyYy5oxLHH2Gq66yBWAnMgsCn2
ROnokj6tJ7oQVM1uKrnPw4FLArWydWpcoz3GQM1S8HMXU28mUReE2rLV9IhBmVG7
WUWyuh+IiOOrwa7pydUDFgsQongAR3BGr303PeLQWZHWjM1wR8q/fZakmR3xknbt
xhGtNvExGmQeLqmyNUCln/Krddqm6H3l5UL1CEoT+ANdHL2CLYo/UxpWmati9iQT
lcvhhVUzD0p8gsYGhgLNVRyCgzg0gS3BG4vDzYDzinMEEucokykLof7Tp6J2BMOP
a2O3g2ugOzubaLvwIFmS2pLcOs57Dm6YhGjKSH/Aa0MjOr1fzzAh37rmeQkvw+7o
bguCVrc+DzChpmV+xpv8mAERdfLCaIypR8pa/4hJ3jg1+im7cmlzbKBHjcj+SguT
o1pDts5AdzbIdBjQLaiPdc5CCowpqykuuzVXporeZsixQswYeLls9oC9uuF12WN2
WDmk1fTNR0HBwjBeydx7hJQ6BW7pVXVEdJIGcosfPcjMkRyndDP4OXRFBsVbj7k1
R+EeZloGYG6SaQIbzMXyyO5vV84fPA+aZXijeNu7o/7oWydRvXjzbOdaEmJqh/yd
+q4R1OPwPMa3EjHn7+HMKy0Ekr18+ojN89CYUM9utQF5fH2/uooBPCSARNnH4Pmj
72C4YXxzsKQUyOiLjreDbv6GG48w5UygP+lgXLOsHpeKSNCgbarDPQh5WVaGOM8X
8TC1m8p3M7x/+D/CfHJ8P7iCQEqrgkL1GCDA7aaqCuM4p24KGXeR0Dga6q6HwEbP
P0btHgXvgk0OUPnYNZmyy2E4FLheDl3AWiAYgLCxgsYqqT/Z+fGLIarxlApfxxDo
ffcHtzu8F48UbFm5mi6EXDV/EjTe2p/Cu9hWK1rKUJJxHEj2flTGitlUEbYCNved
+5cLKkonAdTjpvGhnbfAEO2lNgTTcdfvsViM9BPm0zChTAokw1QIas/HgG3GPhTU
e/hBMEc9jbfL8qAuMTsuVKEJeFKixQHLzeKjtpmBqS7koQY9NDuUvEgO+45CHvof
kQ3mHudAyXBNYQ2Z593azGsSANc2+6yUC2cR/V8YpQhNhh6YF7tNTIcRrx3TwNAh
QFYs8gFCPrypqhCav6CsnsvkQ/WmQ4sgdGTG/kWvnVbNKAHlGHP/oFCsTgOkdIM+
y2JGePElyStEEmnitSv1am+MTxt0HJG4HHhhAnZ1Jkccq0sfZ2+VWUg7z7WWHKR2
cdhVNeq83steNN2C0kfycOBDbHfv9JE9SuxaGjgf89zu/kkn6mrXqXP4GdLLt2Rw
j6UdT5Vj6PAsGMXBt0fPZBoNVCpkc9zXIvuTwgfwExodG6uRj2WlWeUpJj4t/Pug
j/m8jq0+Ot+jr2TpDyymqahwUgkAS6ZJ2I7XpObZzFySh+StRia2DC/b0bOTS58a
ec9KO6GEt905rwnYaSU2RDYHX2b486rJ5SxBE8ZTc1GhvDPeFBYQUUEN3pZ64Jm/
cZ4c7cwK2fD9YXkKe2Ev0z9G8ItrI8CkTVmRdAs4LEVNcwEVaQCKMPZW/6brJasD
VZ8hqqm0Y4eqF1F2nhp1PmKti4yRKiLO34tGKFfTdMEJ+dyVi3riE5RRfGTJxEMA
BDisPrdMVln3qM4yxPmumagfly1wnaUMoObU4tumSsUnot0Syn1yTGpZo1uqwvTU
tLII6MCxbIcXp8Sb5iqtUrY1tOqjmwCRiZTXFXdBmbfnAl/q5ltJAcp9GuBfoduK
SIlu9fKs0uLOOjtY+yPSBaQf6P8XgEA8eLOtVjkaYLbgSaq5yhv275TVLQZMUKrL
TZQkVw3oPFh3TGCTPdhVVaYnj9+WvzptxMYtOw11HSHdwR2045S7Ia7l47py+dWF
8MmPZBqfHtIgHaPagWcS1D1tDyqbijNeaOS022kgvRjch++gT+q7andalEsQL8Rx
eKqm0ntiM5Cprmkh3lpEe584px6ltd1r1jG4BCC4rhJZNkDn3NhiuxzPHUMoobvi
c2bwlvkWQv2W6byX6+f4rGFEMM+kUeWlqTHcSe+SpfGUrIGqVSztdlxvNm2Su8Xz
z39Yqi7WT3W0MgfyiJVqQuI+ucePEA1pyFId1WdE/DxiCc1ZsDYWXaJ3VArXJKIg
yK+2aoBvTgsQr4wLCX74ymVDSAtjfUFhbzRVhgEEmfYLN0UOJLKcBX4ftd2pcqHO
6obc96Bg3kVzICNE/KDbNRlegxz264FKkPunMk+x1k6CpYRc7BZtPQJ8pse/4tgl
jAmi3ssxHHs1aHgZaa7vf4CB1Zg9wIH0V90fiGsjWjkTMnP908Ks67fYtu6/IDcK
odHY9kisR6Sq1HPwtl7FhHn86e1dRCtofEVXD0UNhqTIAEnMRQMD6MtRscgeS2Al
3tPkOmrsN8xhq5/wMX3wReS/OCkzUpswkujNATDp8LZFrbuku9ocFlox1Bt494wF
TtOon9BsOpzj84rLxtDx+qZWy6j0XO4ELBqtUQNp3VqLAyKnbKngPbFrJRi+njQT
LOnIQt6UMYogPiQXkURqVB1QfPdzGK7+hPv1GPQboswxQzi0enI5Dt6LOq4NyB7p
xOwkI9Je7+Olko866hJ1CITWY3n5aSshw8t8mIdN/LvYNWn341eRNYX7nFNV9x1J
kY1TR9Wl5cxZ4QTcTF4LhyEqAOsVSO4K7cLZUXnEro95obnPGA3M+I7uQc9iIc7q
1d2gI4wLqqTXWt9B7d3QCDNnx/Itdr5ObueU5MY7uy6NSOmg39h8SSFX5kHeMP6K
ZvuDV4rp5tof2p89SIgjoYezwVk9uDUXdfKj6cIFO5oeTV26jvd/TaFuXD7pZDgB
rQKcZ7Wgq9jXBz2Pd46/Ik5sXLEJAcd9TAHkyuMs0m0TZKf6xb6cYsAh1E+XSSKf
a9F5H5pzkahjCJwJ4paWyk82BUdqoRhlY7HLDBHGifVUV2ZnHV8j/r/9XbhzHvyd
EsgFPeUiHkE32m23cPXKfoPXluEwpF3tIgCGOdtKJ6ipI7Ku8h0syGDo2dF9N7vC
D/iTWW5GLNywyhod6dtjcvTG/8oc5JNAxhq7r5fgMLCjv+zrUvOsAHDgUHcXXP52
rhWGVGo9Lw+zklwRW0FnFIVLUdLPKljJFsgwMlnEN/3jWGU29jT2+P2/zKqWTowk
PniYREPAgVF84saSUBgcrIsZHVWLv+fnHbyp3s0UD+VeBOpWCzc9gMokBpfdcYqj
Ep8a6E9D3ynlpVX9OL7YAc6bvCnaPx4NONmvC8Gqm6NRz9T4voMHgm91Q0MpUzWS
B9fUB3twHm0H9Qk4ZFpuDZ296OoPYOcScV1jQp9XLxXK1jHYMUBGyW9rzslcT0+v
QkOEhNHxvUv7HkZp/Sjrfg3c4uNKb6jU622zy5uYUEdtJE9MnUHEmJXaDiNCfSV6
aEJeOEHpg+qivGXXB+j/Lyr9R5Ekpp2/dN/KAIzzn3d4tb7j7YLn7u1bfLT9rdAN
abz/0iGXY4hGTQeWNS/MSnVCIzaB1o6pBM6bViJfOpCSbfDa4AansTApkTSbYJEy
CmCF6c98o7IW1zNQJS1elWptec1lIaKmQMYE9wZ1H5ahgpuPFHx86ZqfDajiJg8Y
vqNigIg7T+gktiLBb/oZxejRjZ757/t7Utrz+r/JahXOIUI8jgV4nPO00TwvJv/V
4l0EvR6CJgoHb1cKgQCsYtWDvHpxfVEryqElnqeh9SzlAtlkJ+zziElDXelDgujp
ks+fpnFswEWhIpIrs9APCd4ydHkjTNkRDHxrgnW4jvGha/y7qKEPu7bPmVVUktBC
gzqrnPqZ/QAYX631ejN0J8VY1weoVJH+oueOqibnFawMFlPQNTgRXY0+9FsVGJsy
Wco3zsws9Cvo9iKUpeBnzEz0tfC2bstCEE7HraqzN+C+3jpCal6uI00rS/mmb0Ci
OsdDa/otAEaJL6FqfE1cVIjUnubR7Ncjpsp+Mqe/CyL70KFegNqe+OJsObdKuZyP
gU5E95pVPig29cTW/ycOfxN5fCF/6BLqEyTmSLx0L5PPE383NAoCSYPlLb3iylWe
uDmpeOmQlkZIq21ymxyZrTPxlv29c5ZfWbBjgUK0JYYpX+s8Uml9xIjMpJGm1X4r
cAKQtOf150MHGyACJNbTTRBcgxmkXOSqKRWhQwe1G49zf+toWe2k5quMFTBzpVBP
XKLYsddIh87y/cERgClOtGBg0zVt/rSu/T231NQ7ys9Qwged6/7tCR18LUDwLdqp
GxFuP4crXLrDg4exfXlJCmqSZJI//uvsPJ6BnYD7sKf0/AuFCgDeqVk/jMQYE91f
C5BJ6SJ6c6i6V1NoS/OB9JU78FkPuUSv+cnrmXJvFHMWh0fC8awrvIOMPU6ckvBO
m1qxlHuE/QOc/xb/NRgHVD3bHe+gS5Q6MXvqhZj55dC417coteVFJewPx4oFVbKg
9qf2qK1IUA3BdUBT+TmUWUq9DlB9+SkbKlQw7sz/THa38EBQ8NXsXkOVXYVpn5pS
sZfRMXV0JdiG7xTr9g990zhF4QiyzuwKbU7wuDJAba/bpnOIXxbBcV5qEZkl4ZQe
0poTPiY0lN/8BE5azhjo8NRhg90ojqzKwj9TCN/76sQ7EmMnhxRxqpuJec8M0csA
1OaypT1n2sF/mjFUnJiL6ikL61CevGekAybuTDvNWHEYmaglk+artH8H1X6ICK7d
zWSlpZZoHZmpE9IRaE7y2DbIwmbvP3lsBYPWgdgz08pvBZgEnyTC5sHmU+QTD3lC
J48r7EPZ6g+CGq2hSGe8a8JtW59Z4e91mV9ZR8C56cLwk3gpoX/WAH5D8PDVXCEc
cS+5zw/+C6h9UpokHIMmT1jo00FVhlfclvjOKCJrjRdKFYlseKtNDfK8K+JYje1D
iD2JyajoH60N130qpTMrCAl0ZcBb5DQBJi3+L/aF+fjILzk9fOibFz+WSCnRn/Do
0Gj/MDghpzCQ8HZH1zVJ8QZyF5j5fT+iR1+t/UtyAFY3sZ5vmi3EWjclazItCAne
/Y49QbJTK2OwOatVrFPgCEr0YoXNgynMKrv11FSR0Q+aWu+AhOaO7wOS2a9Hqd+O
UUKfb6TWa9BPfVdYsFPqHnO+p4zsGqqNSuNLkaFgsrRaVrAX/08xqWCWFkJkZzIa
buoTFcQ5XQ+rjMDL2QhmLyixgR6Y2i8mPrS2Rs1aLPm2q0uz5kT9SNvjNDBTohZp
a/sj4LQCjha3hl7AfAecznqdpWv/8ok2WYCBHI9rgIjuY3CzRhN1kSmNb96ZS7yr
g+sktePLEI/rJMBo7y2jDBB/7wPnaISI2E2T4BcOOmYt+ABP+sh8ffPVAMVEx5wj
Nk03uk+smBWRz9eXPWnHwdgEvZNTqvNnDnVrDaw7hIGb0iML0moZFWLimloVbOjt
2+KiEPNGqp/r/DSEXdDTrkEcTlOGM6ER+e4w/nqs6t238KQF8ZnujNljpH1aTDjM
1kg4c5Dy++1Ng+IWbu3xCXy+8CsAekUs+Sgv/CY42gK5j5Leu2ZCklVajUhxi+cD
LdWrvMgEqphZRETUeww+TCTaAHyYflGJrnVmbbPzaxlny+BQaYEO5fjTsG123v6q
ZDKtzyqY7V3WyYtTPSTcVzgHrQj/fqE+y/jR5jI203cKZouSIt3MyvEElSFXAdyJ
zTW3WMPLWvh5P0ws64nm36fNDq0/V509oTzFd9tR5LvejS0okQaSwc6YxpmjSwh4
O+rheAZiqUimMJf3efvb4dtcctYA9TysaXXKv7+7VCbdaF/YFySMWUoo5ZXwrC9l
eG6TElOTvdqLNzb9DiF0PuBov8TMv6B/VOVJosXN5gSfeEZSCKn5D2BEHfLudoUl
WOsBesBx8kuvT4u6zBAioCnhLmWNiPdZlIPaXFjxMhw/vctvWLCZLphvGtoDKdCV
JhmDfi6mxA9HAM90zGR3VhYONp+XpsaCh4tq6yZgJoxQcX7ZShnEQ3iz9wTZmZfj
FLM3RwBEweAJ+I7L1c+D0PUKrPDJ5V5E5U2zASqOHTq7ug3lH4hjXeFBOXk6X1QC
hG9RLtetYnLe2mVJITnOnrmvc8NbxhqW/pTsA3qYzIak4oe44zLEN4Dq/VwdRXlf
tL0VOsg7oFAnq86WgznXDjsDOay8pXIVTFS5Oq9ea490jXXhuAagk0fo4gwqeEBk
2wl9J94EB7M624nmEEtRDOzLUn4qmnRXddfzhMUEdCxBPQKwB71a2QPxArylY0qM
iea5MIghUTvvciQ365N4o1MeiGAc9a8dBhm5G5cWcGe/uUCHG5y5/+h3WgODIJmN
PNhHgcawNzya56Xo+GgSWvOAsV3V/TGemBBab5KOXc071Xn1bUVNpfTfHJYF0LVq
pgr0SzQNpwClkd080v8lTT7dgN/9UsHBop13ic5BZWMBB3tYTn+7tDsr6Ge435h4
Mcjo7jcUVIqbtC/y37g9q+AX5c1771xqAzozWoZFdzie10K6Wg4SpJwjXXi7Rej7
iOvXiy8SL7a4nPtwWY0gRNeRYNoAxVyvaGRJ1HDwoN6RI3aUnbeHP14XX5CnegGJ
L1uXcU/CfLpw8JfeBTDOzcpE/SHbc6pXm26soATR6WAMSQFynKtCgz8dUgBnQbrb
9egnXBkCB6gQxhgKu772UbYKrEX7ObJPmwjShENOvVDS1HoYzof9SjtGHv96Tixo
5aPVKfHCGwDmYlpDmsbfs2XicyD5TapPBb+LuQWb70wqN0xgCIEiTPfVx3b+//uz
JHPEBK6JBrZ2dBfOeGdVgEY2k5ba2u2lnb4JSn4efTuu0FX+YuDQ+9UNW8yzCplB
aL60ZDpDGgS2L6LAFHsGhdQgK6BpTxZD6My7PmqEBzMZKcs3L1Uyw4cTU3UP3Bie
cy589FeIyBluGmZ09QZzC/Ajosk2DmSDA+nAb1tYSkomsFoRmJSI2tQ2kadWjkez
mIV04pZPrn+BKQtvFHOjkzLlXRe245i45OVQwQX0ayMVKLA7YouOEbbKkaGwds7W
9cWdX88qMgmHHlcZ0ikNeQunCgsuTkN6Jw8lPiqH0La2+LbQrtowk1Zyatx36UR4
JxUrflgoRRgJO169TJMxGqJc3dHFkyPXmvofjCi0+7d6oaM4MWA95izdEss0tgxc
1yl+qPV/XcyvKX+IX4dmpq9/ZPhvzaek9jNyksL03foDBJmblis306B1LRNvT4n9
6W3MH5mrjSoe1t/gWH383GD2Thd41e3JOEM5fApIw0+6bBxc/6MqQH07P70NMBMT
yRwPbuTYBweThgaUqJk5WPznaFkhWaTpHLGHSF8cffbneSAmvmzkd6wEAdsKMlA0
GXucifT0vZWxVjl2yMODKsf3GG696RqAfcoppvktSUwCSewkotT2ZYiKY8pvlFs7
4UWeInLbiMBk33mYAULnp74uHU8h9ixSxb6CGKIfDNsFelQ/1gW8r2++exAv8cOu
9RcRIR1GiwtPlK4gvhd9gYOpBPUgZBvQpSKXwyjVXl4jyzL/cOwrrOCm3w3iuCky
2ByKoJODEX/Iqzzo6/03iaT5s6Bq/iDvEBekvUV9qMYAVIKcccrXznr4VqMesu+q
AWZ3Ottqydn7P7LvBZ65PtLDg4vtEEHJ3puE2yqgPXrodOfGL8H5ojNvcMge5Gvy
aqD3nL5AmSG0HGxGnA/bgPpTXl4mDgUAHVSExe9bVjAKggCZG9qzO2xgulvp+CHV
xZ/FbLL+M6uO0wl/QVMKA2cVJqSFUJ+VjjHXK5FH+0Xj2UJt3Nn2ZLx10/Uw1Tg1
BwJV6Z4ziPK64ZQt+15YafanMjqOFd3rKLuGKTBY8Cl/sgQ4T/7xnK+gY5sFmlWc
ErlzlZpGOK4EYIYk3RDKYZImIlJ+frMQGrCFW6HPMQfU3nQKulVzueQw3ovF04LF
dPyu47KstEz3IWxhkHj3+HNDnfvxqWn+XA9e7qAQbrqSt7vGXLXR0gdR0Ayghz04
0jKDOhfLewlQWZklCyNfe2ZGb37aiJR/ZwDxw6PPU62wyenyBuCQzKaKHqdx/5ri
+2RSKYsqNHLyGP5owgfOx4LldRJ5mN8Orsu9Yx9QHhAXvcycdANI/ktpcFil3fwy
lrjl9YkIqQPrDwPtPdL2l5VTfmqVOCxVq42QbGAnIMhpz8jXe+hIhJNQDvJLc1Hw
dS/rKW8EuAQUhC/mgz8AfdZBssgQQQrv+tTVh8eOq4cj7lYsTM15n97Ix8zITZ0q
Pq+wYAffLURooviW9UinAuRidF4iCg1thAYy1y9suJvDgm2wzgxt8jcKQO2SQ0a4
gv2NSQq3w5NCW0czVLOwgeh6yrH6+TfdGyd3ex7XSESvl3My2ya3dG/UtIacGfJg
gHSeT30t4KM1KYYhDtgG7Sn/EKjfq9h/qtMmmkPYZsfSelgH6TKkqWNVh1Yz8fPG
kinVu5o/YggX51o9DCoEWLa3ANiSfAuA0wXPqWMu+jytBKjnXIE7KTJ3PppeIbao
FlnC6iTzsLqHY1vOgScIF7xlvT6Er/wK4Pl8IqPoFt1PSu4AXuqswnV1b/YaXS+v
iDjLKuXhXtP9wzAOyNykN+lZq9465pDOIlxara4glGfDkS5X/Bv0tDbMQfLBLYN9
AQgK9Dk4L7Au09cEDaLlv7dhcBjQK9m7EiHRm4R5yJGp51qPausOeXlRnfRi2qDH
WJoOL2VKFrqleI58Q1Opd1eVtg/JikT61hRae/PcyOq/64p9LcHNa01BxBx2TbdE
t6fzML5L3wn5eBO7UPPEvY3ROffJ0j+R8QL1sGDNWify2jHZwk0O8slkNYxrgMXD
mgbx9S5117aMPowUoMBIAjEiMXA2/JYrPoWezoxm6/xmMRjHnoDu+q+mEbCfoqOg
bMglIAlU6iQ05wLMYQob7mMkIS8S9I2htTUxIGvjo1DYR+AYpvjP1mVH94ntPx26
ResT3cBWP8FHbwxujAP7JEMKlFC5dSDIGpmtAO7cd0uxNOwbYV4XRb47Zv8kNsFd
wrrUVXrFBxtqdgwmyc3gvgGsR0GLBpaXBc2BUZLm35eaSyOsBCKJ8vBOoIf0HpGm
kjJ5CXixK49HNj6DQSPam1PsDoI5mq6sy2wgpyF6AWoBKaIs6gcR7g0Sk0FFOIFq
Yp4xbHP6Y2yLW8mPzUVX94zeboDlfxtUguipNKcRH3hGG3gnG2Jo7HDDAzKPeANR
K2KguNuyLXVoMfOplDNP0n02NyrA4s+sv1rSu8kmXGPNtlOJuKXJdZ7y6XpkCFV1
lEedKkEWprdpEfRnEt9FWW1Ys0Wrz3ot6rhwsMP7fLp4ixOiUfzLeP4ybq3Dk6Z9
aCvAz9uUe6s/eOx4TuGzqr0oRXJHQUG67gy2toXO6j9R2i/itJQ8/nT7sLHeClXu
3oS8CyC2k81Oo/1jJc8KKBcqgR2a9x+l1bPU4b1jwZYj2yWVUtPYQ4RQGF8CrW7E
pcrkaYoP7ay8u96qp0KVNfxzbZclIBVHml770AJLD5vWf7yBdIyCDXeTVlDwzR32
fgT2O2FoSfhrU8P7j+VxjxLJjNp1rw2M99YAicBWWbvfhEgyZrJAygdjVZzDooRD
NQfWP4mctrjxNi/XKs5JX/xP8t5DX3LDatdW93NSFhU2FUU+b14EqmZMaejOVw/B
SP9ibAdbHFAQsWI1o5Q4U2EbkrSNtsTLrFjpd6tIw0C6/lIC5bHrKfz3zPnPcadT
XMB6VWgUDR4hEq8E7akYPHhts7IoVoCl5IN0jhAE97gc3jN+wVxxcMCb61BWdvlU
WAq+DjVYrMxKAzBkR9zTka1QVzEFo9HSmcPUjJxxJcJgMFdW5bC/a0keUsIPY3eJ
yRdU0p/va3pJYJ6FASFpde/EOc6qrB2b9SWZcLna27LfMKuX/+DcVJ+OSwutN8nc
qeKVFc9AIaRG0uuP69HmvG6CyKNLopoWMAztV5Yh3iMQg+AYapM74Up8x4JIMbse
K59NXZCCCPFy6MdlHPNonqtNYhhH43PM1E4v9fiMxKWQHMOLmbM9vlvKxmNuEeFc
a7o7Vw2UqvzL6R9LG60ZxGD5JGc5T8QH612ajP7PlAnwm+HNue6SDOdvhaQgOfXl
bRaL/iqA2rKaX/p0zd5j/V4Ty21hH6RjNMeHyHdjZ3DIollfEQq7MWZl8Ri4PccM
bV0POQ9hBebDmKYwshq6Soc5CjpqnyQUglSbELjdZQGqsX8pbFQ1L2Km30vejLRp
xsnK7ZtYYNnISIVq2uw5/6EUt3i/gwV8kIUS4DsFjl8KntCKTqRf+BKSWX4QNvHL
Or9PYOweRV1rsq/pmjsHEQl9OfG4Xegk/2l7/AGyUOq92MFYnLUYMXAhDHTwvLBk
QgJIySrhcEesZFYNygUpuwlnrnoIiMNM9wU4nYNTWB27r4rAvvzBfUq11RZaPFc4
z+zAWJs5lp8epGf7asEi/qedS2+DkCjKj0X3T97xfS8aUEdXj269g8oXJZpKBMZW
XVDVLLhoVh1chhJ6+YUIVz6QJKBXAirEgJUOWENSnXdn9KSi63zXrtOjSjpDrdBr
hlwyhx6HmZEjw8YxjXxWaS411raHSzIP4T+ZM1OrKV1xh8qtqWQWs0nzIh4vL3aR
Lyj1r+SdQuktgtzxT1jYNjiWA3wCmapB7VuGn35caE0T+ZofRMZvmlB10uuBFLLr
2lCWI7Se+bWZm2bPFSN6ieB7ekKW3Q0yb79nCmAUWAaY/rJCjcFr1dZcb6HgAQfc
zS9akx2/82+eFOTW2ypJpsZJdWRGgaiYSePE7Pl7UQAyK1Qjjm8b/JkGISKH4UCk
CCJmGHQwvu63ZYq6o+9L0i17pnRhWzgKt4I1qYc7gvuOyrv9VO7HEVlmaib/5HyB
YAD3eaSGyf2RxmzgezpWRNtG3D0xREUJp4KwM+sXR+8qw+ELnD6SU9mGYpH+huF1
n3wnIYtVG6GJH6UpQdewYL9STVeHz31qGnFctzvlX86v1roEfEwqFxdbw3/NilhJ
k+OQ/TqLrOhSapA3dPwCUMMdxoGFdj/EEjLaQnHyl9UeqvvjbXW6+RUr2d7nciZf
vXON1S5BR8KrG4XNMnqNicwBL7w/CI7CjpO6iUCR6UH3CLyYox8F39vrjKI8NQuz
J2hrQlKe6ucZu7iySOVXctl8mmlweFcirPv7OsLjawDb7XLUFyQmlbOz3eClwYsi
ypwXyaroea0AHaeke+dSE8tNy4cWeK2Iil3nAuy0QSHZ87Qzw89xplYgALz09R1k
Y7qNkUovm8ZjWhE8QrJChebFV4aDwtVUNgTk5OP+rRiWtLkCRStD+QJgXXKP6lUp
oSH99DYYEjn2zi4xgKVI0CO6Zy6xuEuG5/HlD2mBZJCoU7CIEiRYCCH9o7R2FkU0
6gCBntaH1uN8JLaB/p8MkmfN+mE683OoZ144yTCvjD2X6Wg8pe0kTjjuFO+NL9o6
hpBdJx9IWirMV0GiGDqKmjntDwsdV4qq5LPiOrl9i4wCTUpuTeZhiQ0h1W5ee9Q/
dDYRajhQfIx8vkASUPMGWYS2D6SWWq0AjSE2dAbw00cwfqiAcewIzTZa3QsRLRC+
fa2DsdZ2rdIL5xVMFwKi06euXTaku881d8rbzpJBL4+192oPifFnMXMuEwTlc6A/
zEoPcJ0ett+EevIY5vL5XfRENkXohlMwEbb7eG68Agog94ViYOxBCpSQY3zO1CV3
aaIjR2vJ0x5OD1/BvacMjhIxM8RIcoUnkMFk4wy0uQ+8WTFiPJEW6hw8h53Y0FOP
QVrZbFFuKN2Pvjn4FOSm+krUEdjWMNJbBlo+wYz98CDQvpVufppnteA324Y+golr
L28reL1/W0WVh5lTbaK/h8s+12NKwRKbVfl7CzC/NSqhuOeKkBu0mEMyxG/1ij9m
IgKoSEzkc2uPfHAUpRWV2/N1YAY7xK0X4wkCJkFP3/1vpKuY+AKOnff4rxEUH43d
ILwcnYPQiAyosp8AfiZwqyUJR8NKWQjI+cq5XNxKjeBCpRTLB+lccXNup/9NWhNQ
Q0Q58GeX1t0TjxEcbi2WVdARJ9njTrHw4VYH5lW6EHS6ltksVJpaWo6JBkrLSK5a
LtNfQ1tQkuHL6Em3ItGaGbtElHUoSFBN+bzOy4kwR8/5nDhYfcX4ErJtIGWiWulN
h5NlmUgO2m8YvfspxhkDzObHSQdHFhrsMuTnXmaCpwqevGDaeQilnFyMhJxc1kR5
+ZIrxUGbNeiK02/JmHp7vBCnDe7rcWeHiBPmgG6PZlHH8aytR6QTiB/s2Yo+mGmC
BccLFyReMgP3VipBVs/NIXDCbeJMN7lRUmhtbycouu+zFkJOJKoAMKe4Jxr5YhAi
vIsRKOwpyjKFKuGSOEtKt8wzybogQyrB3ek/HS5WLXScVtjtyOg1Qssn6UIT3P/i
TYi2Fozi7HaVjgZZGOrHOWVdz8rIKU9VFBEnU7K60bzp6zFx6yIQ5+1zf2jZRpRd
HGeXp6JI0NmZaxmTblDomzykBo62pu4eVq2BpbbCnNjJYD55E5Nl6sYRASsIp+JQ
5x4gxkPCTMRzOyvd4zj5f1KjiljA4ItNTTO1ZsV6fiK/h5swTsy5/703R+9Elj8r
UObGRPjGCAjCLxirWCkfHETHOBUIYxXsYR41gzhZXKA01gO5sdZGfKplPRVRCKR/
aIovDcIVRki/nbpi9WAI+2LYEnCyCGqYy88lbNGYFtceQb02CERtuFGYyqSsp/r2
X7XKxfgsmZSlzXfiUiHrEJNMmrCLR4thMMGTanhYAXYncfrJ+4MoUd0RmdLA+eh5
OXZPDHBAOD8jKW7koaEtZXSalMyehLGFw7HLjI23UhvRbsM1PCL9ACH75TyR19Vn
aqMOcOncqxA4L0CTLJkz0I7ZOK4Ysz4r9kPgchBEtV+sBXStmI9a3w5CxEWCLiJk
SpAt2qAy+ZAKaUvZlm9NJSKiXMO0WgmJx2hBGSmHBEdR527OVvSDelWPx4juXbP+
hIlHFOYFDbrHV8nAI0coLDJj3GgpnP018uXS4kuVpBJoM4HYRcCqqQ9jeXiNRz+Y
dATM2rj9TE9mqPzP/bMP9HUXlebZvLWBYa3POVAZAhZz0EXQJBOPQCtH6Dfl7iyO
9a9b786CHLQmLr2FkhDYYaN7DlMqfj9jwRGBoynyl4sYZSOGe57BS1JX21lCRI4T
4R266C8a/UGdlhkZ7+O0Jj4GNs/UQV8IOiQ8S21LJH+/yzupkleMTNe0KBtKjXMq
5XUB4QSjCHUJAS0KWtrGQmCgKvSST0W/b+It4mYedQSXFzQjGoR1ldogkP2/WOFD
8zas1a8Vne3wEHvzZFPDXUVS9BVZsfZBh6dSy37iCZjUny2ebr9MYigwl19IItBt
Mgc5H7MKKe8Lv2JT2R57zN5fzcdP++knAYKg94gWs7YIeGqkoMx9fOV5SRT+6mnD
2gY+sedG35ksNNf3yAs5gBX0mP9hEYNkARJHDhSyiQyw8AmkV6CICip1os83rbmT
fM5JVvs9MVEkrvm0Y0R5VNvD29W3lil+GxqnQ8eAM9HH7tTR3SslZBKjM9r4bCoa
+R8Hf/GwdAB84mC8Pyttcill99nzZFlpQ0iU5npNyDeNwoaURMOKcvp8GNQkuwqF
lg42hmzzkHdUzsMRc4HuXG2uRkUKYQdd1lakMYMBiU2smVmjD5GrmJ1zdsN/4ZaF
pYXjR8u1GAq0uJZse0j4B3t/r5vl/I9/iFDDRg2aj56HZhesvm5phTo1j3ks3T61
2f/wVeKgL53KTE4KbcmmAjRxklK+Rb9hkRVniN5/LoAIc2y9jA6U5SbsMcW5lOyc
ebBAhsMzKQK/NXz7vCeeaQoCgPUU03J2yQnDXN737f5UQPf8u5J/vuRWY86+uK9e
VB7jEo0ni3fMqqh/AqD/P49U0ZjA4NA7q0umA1DV7/EWctnMiRf7TaTmYSzjT4Oq
r/T5hRsuSar7OQTDB21kP+TarQa5QbKWtS/vboI4+26p49HX1Zo0sSQVj7V+yIfc
wkv3L2lUzPaiq5hfqr8b7BjVfkqqCk/0bPsICSKxKjAYId1zdV4M2P/zvUJ42bMv
RtIozf9UY0ElsGRCtaMwYGoREnYxCBHtnShAWEQ7goupArvVmPOsFT/XfKTYqH2v
3nvGU/82cRCV2XThtd/V66Ll7bNjEuxxlcdU+fD6azC5of5jB2dWp5E1pCQtARkQ
VzI1NoffJWshP7GKid2sDI5mZaNVkytr6b6kdbBlwzW9yUoaHU+BHuV0kFJtEPlC
Urx5rfvlOr2YfBX0qwF+0rSjQsWUJxzrHFyymDR/P9zFDg17RawMhFZtpvhpDLay
MlVLCgJAxggS3Oy/zdvOiFZRV3vNSt48koYtcIdUazvJKIRSyVogwgTNyXgyLLSS
a6f0NVFqABxsalDMjsyyktc8PUYxHN+ZX5kYF2qzGpBnVD0D4EPoyRU4NJe1rhK8
ooud+6di7qXVnd3h++aJZJGlai28Yhd98tSjuG9fVKAEBqbwi/zS0RGm0CTra8/e
EiQOU5Y+EysxYuZYo/XKxcREyT9GGUoYxFCEpb0me5NxrpDMalRbFCQf0x/3QLS0
uY2g//J8+PcnhqOc9nzWCPZ2y8Hjwfm0ZZq/lF+eP0uKhL+uRjUPVJmPXCX5kUHp
mGDpwvLy75tXbqEg09LyyrXdUMcPjQKF3t4TMxqEfHVN2k4HedDiFQ7sTGMrzAje
zXf21MR0OCNcv+oe1CGFSFiBfdXUTpwEfgsdsZvEgvj48SZoec1ilMnoLdHNlqxl
d+NdXLLvXZKvBQoD77Yn8EvqNoQZ8ZLT9svpk+m0ILRLdvL5J3BH1srkAoiTICIR
fURfhsHUyBJtZIHsATECs3kAo33frrVCP2rEn2JZgQ1tXPiGKqzeUssCCscV/S6B
KR8udXOeo+nI51qYE9OMHOnwiJ6q8eQ7fVgdycNWGFD1altC/uKYiDA8H6BYA+3d
Zde38XeSDpTqc2U7uKURBPva78K6P6XkrOF8lbvPhYDoLefS9bbPJ/nh+R7qvv1x
7yxLRg5BGf9rJYVIBbew0SW25ilsxhonEgqhNeM/bZJf7uIUsY2g5f78/LFKx+tS
rGTxz/bLS8GODI/Zq44G2XkDmTfoB9u3jrOTEesPJstxSROHwd4sz/qzGhShBTkR
4A/QHK4dv3a73gxy3r1B2Su8DGcrfWoLlM+w2VBJdqJH0p40pq2WjHUWiE5XrL0L
vV6J1J//Ufw2VmItTSJchKaQLEPAB1W2aiJwad685E8scKosr1sZlot3tFBoXuH8
gh+3vrUUtpdOtRYeYMrZA7r0iuQXwZqJAYtailO64iuMUKgrn/l+ZixNk+apo2yM
/EtTJxcimbXrKnwo5484qkm+KozUWLBzEyna7i3qPPpAs4UYxxPF6mgotR6n3CWI
uKHZd74VvjTBRrXTIQ7GrsvkaZnadmlUrUXxRymUhM+V1xpLdpYrHDoSj5w9ZsAB
xw3RGnRqHd2oYs3GVlz6QKr5MX6CgZaGDgvCjr/utq1xPtC4L+Aw85fNzwT5XXHy
xuFTnlraGcekQxglmo2pHUxW8BTmpjxzu/WiRkMLuS/DWwavfVPo2o7+4ImS50QJ
TqDixkZnwLQe+Z1xzr35/E/l+96W+Wy7sKdIzkcdGAstWICTkYyMAJckNhxiiPVU
nTMNqk0x2TdfLCQLmHw4osJUSuhi2ixxKbwnQQOi0FdAR1XwevxgxAxWN5nSo6pC
8Q+JhFQaNdZfwA3O09MQ5PZNGwzaibxcb1YkM03uFLpB9S2VHa3h5TcmhVOCZGS4
8c2LHc2PbQB+6kYowCLWhlr6oamHE39omaA1K1gAouNWFFvP+G15HL+viWwcTWVR
RrMwQ7X31d0I5eqtkCUow+OSkq122rQhP47lT69XYJcq/426Z8TNjSOPjKtX3Uxo
AiEZY/S8rDoiCkLqSIJuSRPs/6ugKOkl5zka6QvLI/vG3oMLbN3zl3bmZ57rNw2p
mHtUKobKvAGIsZyp3yH+uEMPO4Aa08Liqsp/hMaM9c7aUGSuXtWWf1OHT9RolNfU
aQytkjMKhtTf4MLZ++B24LvBPMs/Rv/iUu6+b/8pnn37RMqJAMKH8SMeuJZGL6op
lZkEzGTgaxjDFEyIibQQKZ2UVb0jmsx2yu9QsKqTrHx+FQj4c2hi65ZddUDBVy/R
zA7dVXaOuu7aVpiRN3CcTJMICPczSDcy0A4z75oQLHKfnsOkr1Z7sddckb6IlEnE
ayrIxig2j70a9nPg4YUY0r6lFAPMMQrxcdWdLrad4B06yNBsthr+T0UnKiNxNP2v
RTl8r/LTeawOxDmw0Q2y4NbtoN5Cd+/2+7od3CR0VkNZbqypPjngfzbtZu0LyGzn
LFmGyKRYBKRg4VwY5OybNQXnyi0e6EFW3A9fQxa9+/+T9tJ6hVPA6g+8TTVe9vzd
NzsL/BixqgK265UMrH5uN28Kb9/ulfwk+4MczGrmPgiJoOBMEIyNY87mgWs18Bq/
rgmJfqvDx2fEJBnfFd+V3lWwrqzTaZSXjzfPSzIbUz6WYhF1juiuQgBZinM2Ik2L
nHPINwAICCQrYKFB0wKFv9jn3pwbmGvxAAnD17dKgCYO1/izeCJR/44GSkrauRgY
fw/3dmQqYNAdkDArNGDFD6pvwDUk4Ck8Qa6yF940beR3ZMCuM37UqTPHptIrPpTj
Msu0p8AqDPksxx/qewfuWwcxCQHaytztNmVTE26Yc5/ZI6v/wWyiaLWC2kuG4Whi
QpEfWf3ajQV4hzdSi9F/iIncS3uN4tcIIAS2dQa1S18pBWI2SCd8r4kjaE3i9Xyg
/zzsp4ULOipIP/PdnTyg2nZYrHRbZzMACIk3HQ14t37otBZdKdshJBC+WSk2vtrW
QpoVtjSOtI+qV/guUG9MQ/ABKKl7LYTbPMSm0S3S1hf9oLG1Nn89/ePITB+sjlbQ
ayYpw0ToUABlPE4llrfppXQFANdxOa5Kkbzyz+iU48nWGKW+Aw6kUQlR4BAJm1Jo
UfCK/yDVRMJOjtw29qcUfF1RPEnQr+kESk4BHEgPnpC5za3HbzFdPrVhIpLs5VwR
ZSxmbX7CqQE3+/uxdZ+H8GdiyGqRBKJ0GYyTUVpFanpmm1e96mhPZbEeMRVhrzrO
Vl2HALI3LsyAYNgQc/eLh9Li4/Ve5BRWpjLMUaAt30InNFYsgsovK2M0Jiag8ySo
Bp5KcTfeL370RI4yehvySfst9Ojmj9/9TXCHK9MZ3gQEo/wHA4LIYm/8bZX9FgzS
7De2Ckqlar2C47L9PaCgE++nuwMuPMq90bCIaNoQGERQb6L1NtRH90upa91mMpTH
5lSb8C7BlEqVuCaDEH/LDYYacrROPbHfwMBDsMvg2hc1oWR09MZKpyMvqvZOEgfi
GDNnXvUPUjcCU/U/fLp4IYFNCkG6XQvbbI8sAIGdBnptVPOyAzzqoYuLw66xSO4O
PQlgkPofnjkoUPn+JLe9sjGCUlw3jWyln94tcaujqae4Gcqpdw+ClrE6LDTaerTi
53fh59IMFGCa8ztx5Fn9JYdH5LWFruq+McPZlBsDnTHmAR7TB4N4iJZixzUCUlQB
1IlAwAl22Rbb9X743u5o3GxgWIXgfyk37laNqN0TZvueEwsCqsNLS9g/zcZJNDiO
04VunNae2A10Qco2955+zRXMBjmzUAInF9JwVGBj1ufd7/SOGLLdEc5ZQHa/kz5b
J3ksAoJSyCtIzTU/2VQe2icnLr3hljL4JjG20+dZruG3i9CQk1rzLbmQ92YVoGgy
6RAcsiNWxEmY409AlNakKBL1oIFjkcpvylbZXsHPXSkuciOdt/0ZJZvDg5vpmkF+
Vp5aXqj6z6uvAbxMLIw8WkzvWZChcWh0Jjjh8SQLfqSQ+gxKEiYVSNYuBrB1I5Vb
IDY0MYBF8oLSxCg2Qd/Y7kwhY+fmRfJ8hwGBPWzjdXvus2UAFxcevH3lMp5VIvAE
V/A665KrYEQxre0rnN7eYXCJNSxFZ4jvD94iQ9N8O+jEukwplIyj/OhjfHobkthY
ax6G/+jjvBTRDFmGhnvGMpC4DS46knyL0LneV4ussabSuTRggVmy/zs2bhSvlJNV
5ZuVrDtADZhnvYzCi4NwJL9sJh8t2It6RH4CXaxjOKejMaiIXIkvjb9ycNVd/Rqj
DE6Q0rDPMK54XKflT4j7jiKM+J3b9gtwlC3mFCVan97gDlEyn38h4QIPaqXsOQQf
3Zn8Z9yhsIiuSJ8TK15u8Es7/c9LduEFxWmdiKruwqQkNdrOCPMny6ATuyWDUF/M
/xOl9l7/vBZkcf4sD9dYbD2WSKQFUjYAGaZL+r2UTHX5W+KvNDpJFSjhbY063oU9
6roy3NVS1Ft1yWsJSdCIaH8rfh/lNieqOv1kvq1A/zRQoZ7w4OP7RDOGGYp08g+Q
FeMhrcWUqrlfXLZdlUsmYjnYpr8n3dZRTcaBTzVBe1tiUTIZzYliJDILnVS69ySa
9I5GRfwXG0H4tKYV+fNcG7VZzopkPvTgwedWcY2z4UOxoam8uTRHzk99AerbL2Wx
Utt5Dg3BjFBMbfh66NpHVQ06KxgvUuBa+f07xsNH3NywzqJNri+C++bcisylEAzJ
qL3sRxwLe5jrTpMx7L2/2nWDXgcVnzJWYyaw6ArLo+6XEo9139ej7OJZ5ctMRyWJ
/o5wgQrG+mtjL+UBFQFoAYx9tryE7V2yKjHGHLdZH2ntOnDELxX40+9TL7cDRX8X
Sryb3yGEJ7ZhWTybYnE0Ct7k4Fi/o4je4SJG9BmPZo27XnjSczw4arHMF7Shxqi0
jEUUzj4LTQANQzE9SlBzY6U9/8T6fyl0VmT2APxD8scPPNvneluBRgzNm+3Iryrt
Kp+SiuzOPrtSndx4BD+Oi1BCTnYOeju+YmYqgXrZOMjsWOkdz/amKINVqTVbpHpV
DcePZKdmiXXSxpxuemhNmrOaPzFA1dqLfq8AXsIbHXJi+SpU9z8lllQeEhIhWzd7
9wDcV8GRDyNwD4VXSbPjTGrNmknL9b3/31tvQ1XTxEIp/qD6hHTWLnDM3Jc5SxLh
u8HKbFMqhAAoS8sdkrfCqLs7O0J3vyte9bib3m2yOUixRaLe7Bf67kqUKbpTaQKv
ORFBPbPK0Tz6ZYmiqnooi5dSrkQrN2LUeSUx9rsce4Q7QEIS2D2M+Eh1AmAC71Ck
DGaniwo6pbfM+pePbf+sDJ0QHLkrks1s66+HXDbPiM0lN1IxXbyQwMQv/EhFzpHd
Tb5O1lVDYfH3GACap7AK8BL7Bq+CIwnp0p9zoCXPGPn0JBy8qwqmMXavr4uCnnoL
UFpnRE/WvKAynbk/hNx0WrFkj447MzZR/4q6jMa95u8i1X0tkxuUTX9UynJ12Ueh
v9vvyd34dQk1xmG1R9siZz/ILFVpM8QVwgF1QyEwWXmzi/gahswCncA+Lrqvw1+y
CmefR4tbuME+oxEnjepv2Ue8t5DrDGG9tnxMj8f8AiymvcFEaveAbw3dlbRVMgg4
QsHPrM/9hi6+lllr3l3hgqBnCE4DAabZMBeFyoXLZyHUfAwv3HP9M/PVKmRpP9Xj
RfYikkNkZFzOLWUqq4hmD/OJoj379CgvODIh20IU7+SUZBsdym2GhuSUn4jl2FKm
g46kIuWNrHiFoEbNqEwxr8VwBy20G7SLBxatzmYTX6E+PPD/Dmldc6fOGRdNl1cF
vDW733Fm2EmxGpaUXlm7jKSYlxoXqc2eysV1Tn1qKqtS3a09AyRxdm2y7ZYDnFme
AZqCn4teU5PWIIimcM/mZBRFDacFuvQwu/lQgv3odACtD5Mi9fDiiwLimuYgJZtL
EgKPdJHmnpoHD1+GHBRzUbZIkeJAtc/Zyr4i7laEv47MLAY4hPRTdgdMsoCuhoC+
4CmNmKP540Bsob0zE1UfhwhKbad6gxzGDNasjEd+9O59UKX7vhnQXle4lh1x2r0w
bbJz11xKLG6CkiVv3Ll6NR6Nha9hb1gEtR76YWTPMlphI1UQbvSTH0xprVvTXX/H
6rOYU8Gvt7taHugl+u0rX1SgBAqzBcZyHCMPHNCESVCJmVTyow7oXdhl/gZcixiq
3hxQ8EFQ1e6Jf4iB7O63AFEkeG2uXiFEFwZ4owecC89e63DXNkB6wrGNoxP+5KAk
hukxkS+k/ACQevcrcjDfIqoGHEYa9FEQE7JIvk7BAWgrmlU3aaZFr8P0rqxG7ech
8VttEdDLO922TdV0c1Tbsuf8+bZS/JTQKbugzESuRroKrRLcXHG7tfvgGUI3GjZs
/tpezRTrHmOBWhmLiT2+Kz2AHSEcDDOdct4q/Zv0F/BNwCin6Whk/gQ5XlqBnBSQ
MNIccHOltIs4KMvgqC1AbS4IEj4XVlIeFQFCMqluSmeYvl/ldMSxXU3DvHIxMBSh
HU4ATHl0/AoM8O4TvG2ljbA5UVrM55nss3P7tBbQH0lK3sQDx20FHyB+S9gkUuqx
9FhusMTF7A3KjU/co6hQRWZ8xcG7oMA5bHOqPnuqH/IaD3K2lQrcU1gW1nkwxozP
vLnMrWgEyNEsvnWqJnTb8Ahclf1FjgrdOpVFvA0FwnpQ6qjDTl+BcktMifUF7suD
V6eetCO01EEJ3euu2hgryJXPYtXZtZCSFkKwmKg+pBx6iXWf59c4m2MzvD8LvNsJ
uGSphAeRpsS233EPGs8JDu9dyILBp+v22iGfNDQX/pDwu44Q2DFZu/MRyeEtHSFj
hCgG6INrsbVDsOeGDBIBFhzA3Hx3XMNM9fXz8lMuF2DTG1s1mKvAWW6lJ+JlXBH3
HhkJUzcvj1K+fP0fsLGI9gXiYuavDVL9m39SjYAtz95ubtIomMOg/XIMbMFZ1Qcw
vUwoab24hrgXmrNTLfhd631O+rWgWcat0yV30wLC57NIHyaPg119Fv02dSPReT1T
Fj9oB6NDKZzDgakgw5ui8nCqTNjHTNPMTsnF0yrB1KFtvCNUB5TFRW1fAu1Dnyr9
hcR6vbiKI09mHPjWF3bgz5vFN3InYMAJIyKJ1izrcLg+bNuiDGwTcxRBq0cQSQyr
l2kk3gkTMyo7DnfIUhDbCXmzDQ2rdob9NmxBLhzXjZIP1Cl1aSrfH60dHNyW1q0N
ywOXhdWO028IGEzQ6AfkTnhCKJwq9h8yeGDLpXPjMCX7/RUtuLHnNIKc/CxD5IDj
9aXcl4jObdyPTsxaOP6XPqRg554zK1JfrLDuZ7Mnt3uuCR/vSDXZXAD4ut7+o+EI
KSs9MYHZJDpPzdrFBTQToNhYFGeHpeiHHy+KnFCZs3CDaPAgalzmqzzmovOqjugD
qkt1lSl3U+vMmZi27cLBnTLHZACVXNHJKyjwDR9tc6I5ccqyu3uzwHwnhDcclo3H
Y5Hr5kPq9Kb34YbA+p6An/AEu5QlaMVZm/rDy378ACLdEhAQt+VYz5khosRxwq33
WAVHN12bow2F9q3EcAzlhyNKr8H6JXWIuEiTJtCGvD1/bP2b6icjfX4VjPpjjgES
H6dBDbbxwLKHt7VZQ9Kdg4rYHMJDOSg/8x9usV+vsy0CLw1/IU6Vbrf87Ahknknn
A0zdHv2rGBBwQhVtFCUAM+L0mMgXEpV//A58uzPYAUCqk2jo327Q3DVz9aZyE3SR
66AER0WzcRNh78imV1uB1BMlHpBUhCpHp/tMsejzOyj4IvN0iSsTlNJ0AILqlKmm
PcLMbbt5Uxzl/QxknTor4eU47U5OiF6QuCr2/HBdl7+8mxey0CLj+aNNq5Hui/0W
mi0YiBO+oJL/+20ACG6hpawN+lFT012sOXTtoz6X0YMEjftpdrhAiStuTkSsWZhL
LL/HKQgeJGmu+ziGwr7W3Q91vQ9evRpd/MV3h7dFPs95wYsqPwuGibc5EVsZkG+P
SPEfdQJiEnRPTiBNKlwyYevBeEHy+FesRuxFk5+gyb3Fpl83HlXEf3g0yXfMvAHI
i7PZWP8kvKPiM6/qge3Jv/qUsJ/VY9yosYEAHzNu8+igPo97KT7Vpy3L/bc+EYA0
1B424SP2Q+PtxVppPQ9qf2GKTXwHhwN9VrlEMpquh6yOkuWjglSphpDDEXIGjprY
BkNzO5kXhY+B6vVabDfL3xkz1uNk0vot39bLWbyxDM7ftzj/wbX9RfdXqk0LAWyc
ePZufamhz933ZC0L+d1N2GeXKrqaADzFd0NT/t5ZigQyYC2rhBXRmrI5CfNwSirF
JXKqB5w8wJlbNlbLgHn2TLHXq3toytoUD4IJVj9AbQVCvM6Q4yTmctfrUjObG5zy
VYVZoASnIXjeufkfRDezgDID4ygunbMYtJqlU9TfpUttzBJY2SEUXsJm6hQOgHvU
QGNqMRRkvcBDWwhTI9AUhGcI7JzTcI/YGliMghpj4mejXZFtBnkoxqvPKzdzbCWJ
yf7hz9USfVgHVVrjsSuUHPY2n91zjhxl9X7M0rR4lEa32qEI2ClM3Ahdmtn5yGRb
U8lU5ZU8/V5jFNqI+KZL50XBmfr/KJX3TAqiZrQHcFDQJVvpU0bh29uCv0WadB8K
O8gtjfhfB6n7zYIZZXEBMpoouJt9Ewc8wJQjHk9+x+e4z6NdPbQJzofQPTpMhGKp
qn2xaJPAL1t3ijv+dGiJRylGVXrog5sVpXav4Ru0kEgGkrwsC2HMN5BSwG6i+I8+
nTBy+LGlDGaE08OV4+V/ws8DGs2urHRObALu8B4Of4L72MM8nkS0A1gNTT+MFwbC
kW2k0IoQnu/WbYxmmrO9gOa5xEnwIQ3kDcsqp8atrxm3zynuUCG9iWQHenKG0+ZG
LCYtXKEGWbZD2QqeN2/xrgvLj1/U2nu+IvF4BLV/9vF2/3kCcaNegQVWAD8aFmjt
cgDusq9CziytqcmGPvUQiYVOpYDW2LBSEEBI1jdN0wmPNcWQDIHzpNtlklcpg03Q
OFH5z8xB+l15soiyEoFDb1LMgv6mT1nWpG0CjNc6YG/qSUVXJD847AbfajLEjae6
Ubm3ooMvh/pkwcWIOcDsE6tMjc8rJj+x4QZ9zG82cDAokZee2vnqMU1omHlVhDh4
FNBG+KIj/QK54uTyDxBilDOJ2IQMXIBqeLwEPE04GUN/N4q/la5rLQoxbWRMco+2
ENs4EHVws10SRnBqO5JrWlrBrTHjGiuz3Sls/V0Nac7Bi7khM4fb8QzxmhQJMdcg
prDY94m88IoHNej1bcMI95ih6SwEyP3j58ZypptIRP98G6FPrbVGmzArz5AKBVq7
+qNk8LKkzD74dbiyY1GD4N1GNCJFwVSSWZ6HL2dseetDjDVdR445oN44JGrWcTf3
rER6hecXiy+7GbDBr5E+nlj4FFda89UWo+KnI1Dy6VeT8RK2iUA4GpmuWHc7sEmy
ZvQqSOMVjBF9G7PfocabIEvXoo/QQUrMyRHK7vhyZU2wIPXQ3KW9s1IC0ngBPtyy
G1JMKIDNsPj9V/k4/rLqzV/Gdlw3vSvlisx72LK/Vz3R03DewXgmGp4QYOUpvpPt
Ol7+vQ//ouq5edNoZ0uPAPRPTm86/F8wA1Xp+uwhp+hPidWDMZlDhxquhPCHqiPd
dM5estpe6Uu7zyngDNFjdRyawE/X8AdeM6vc+EcezPIs16fXsxyBprkAIx20z5gr
hAa6xgnedxFROiaai0uLAgiXvF+nj15C7ZYmN5sdcHO87HXM3P3K/oOrTcKZLG5T
/cMb4JyQj6w3+X3LOn7Ou3uA6wvsrStuJdP4nSIGLLETk3IGw6H/xuIXPPSVDHsZ
HP2WbEuBkEb8KkBLvkvP6ryRPULNY9FLuGOQ7c1vuusgCkvd+KEQ/JdjznA20Kra
Iojdb6wrm4SbxfBFvW5HBKeAmy5MMfEeKKsz1rzO5d2oTYTRe4gnM7lQ6/xPNxjy
3dcCaXk6QRjMyr1UQkv6u4G+X/3JNI8ybnawQ2Ibc75HNssxdOiGdoW4TlndcgJ7
Due9CBW5sReE+J2ohU1gU4Pt0dcMHvlvfGMnT6txgQNkVsGnxwSbAAfg3f3zwTzX
L/UZalv1Dh/7kk2CDl7QO+7ptr62JMd9P4wvrlcMRHo4s6funpMqdM7URu27HH9C
9a91CDjLwAvuqcM6f6fO5oaaSPjoLrisYAzquPt+4dtUArzJV/tE4armlYImqP0B
0d7GL3cbXAq4Yh5swnzS4FkHnwHMwx8Rzf5z3ucG6k3ogMLpVol75F+mGGVkL4Tc
IVyxr9wW1sTxZ6o8L8K+7j0CPjk8asC5Bjfha/ZrM2SpxIyGmS3KMasKbQwswdBZ
bXcagVlV3k1di3qHc0PFtThn8+ujv337q47BhTAtUWqGPNpFg/vrPjp/JlGRpz1U
v7F4P2E7YdELeOVtnus06ujLKYS8aWjUJaB4GVPqXmaXZqvh86fvCp84GyIkzmYg
NBH/tf2QW4hsRntW5TfTsxqgIKODY8SB5EwoYOj1tCgRaqSkktjlw+JI1KubPnnK
p0WDokRDgF86EHYUpBXzBgu8uwXYgM5lGXuCNpB8H0HflNBTO+RwSHd2z+LGsai1
KN0asXhRaU8fHfMpWheW5d/IM3qX8jkA+fwCTJemTbchDA8ZHWldWCMLUbHqyNwe
ADWU4QN6+4aNIT9IvXhvZXFGS6evTMf7BAuo7vUX0yAsOtleJmsS+9ZzSSjlucUz
JYwHzZ+74wEXtEAMRf3TPcLYwyA74PkePJmB/P2wbqRb5lhomMG/9xR0PI4mqotN
Sh6ofzzmh1vb/igMCCKXNRPd09BxxfjumgAaFH20r0ZyMXOG7uOBh+3OTdSSpCPs
8AwoZOPaWHpz+1VRgVk11hp3qK/oMSNnysd68dFxNBevDbo7BwtgLrz5CLim220x
hKTjSswlZlTVCvYRUZKXo2rmBoJk06qejXY5A8WIZgyn5vzVNs03WIXH6ebCS5/S
g4chISvHJ/I5XpBQQ809e1LYLDso4W7duQs04EurzPU9Somi4xe3tNR6A6D3KK/x
tOjVxxUmOvUPRrjPMmeWdzLCdAtqh9V2PwW13H6fQzK2U/4Djp/MGL/WEyf7w8zn
n0+XpifA1LKhGd7KgznOaWyDDP7A8M+hds4SdFi2BHn+YZ1Mjjyq7Tebugn6BtUl
8g+kXhOyYTk5Jf4PwD2nltkNgWLSu1DQvMdwdURs9JZtiV+qtptAbm8xBSBnWn7C
Av9wiuMzE2eivYqBF4Hd2a3uLkoYJC+2wB69QiOdGePlqHsFi9k/BYp672Rpdarz
yqHQW+iHzE1xFZ5KLFmWR9hm4ceGvOXL3J+0nuB1/a+Bf3VgnliD7L+kTNFfLnW4
Rg+Q6NJqCY1OEAE6V0vdCMWzxiM/yievdLpadkqncti8NDiLsrp2GKplgo+q4ZK0
KrfGLhgkbJVD2xEzWyo3UU1HM46BQh/wP0uRe4UYwE27oBtCUgiUIdjewf0iVhW7
sMB8l9v9rImsvj8ZXkrPLf9rshNDKdNZrVKr+rCZKbD2fsPV4I3vTg2QoplanKmu
z17ee7STxYelptsqEboNPTDUaz/wRR7GVwmXd21gmOz+MVufNE0V1+dpmhYw/AX6
4deHH+EragW3W49RxqgZPWiLEpGEGGWNLBmTgh49QBHP7qteg+Aj96IH32F4Xtwg
kTlYnRPlH7s9Bk/eCVKwcbrshcmSkA4SGVtaxHF5IvyVV9/cJa2Ob329gSeKrTuU
lOD/sZw5O4h1wLou5zx4yoY3gL8a+q/v3Q6f/UgAGe670KmtPe6qj7mRltNwB5/U
eETMpqrNa7q++Vr7a+bcjuQaqRxqSnzhnMmMxYNvJAxkZtcVAudl+z6V+hy6GJ15
pQfgTdkGuSytzCR5s7xQDqTccVyNAEV8s6hIKFIr1rMI0QWIarTowAGAE3qM0Qhh
r/go5VqiTSm1zVh5lBJWFk7P23ftaBqTdmjjN71AytRhq8TaoCWvj/jJXRTzaq7L
X50YU8T9mo/MmPeTyYrg98UY/u7TWPl9vRDmv+IHT19hbZ3UJ2AGCf0E3kfgLgD9
twQbAdHEwFAXWuPSMZiQRsJCKwrAscbfzkIrFBdRzlbvqng3abuunBfFGhsb7T2f
lfVFcTcirCwywCzUm/ZcnjDQuFV/YXPX7+JKOAv40L+WJJ8cL4lxdlLjVrI+/lbv
zg/Ig+Xcuinud0THFQSWIUTvvxzGhZRX9vieBUtygVJE+cfvFVB8/bCGYoaJvnTx
HmwWwx8WN1b0OTfWa3DJVd8h/7snYsNug7+z7rI3bniyPCYkTf+JLCTDSAb7dd5C
TiD884ydLPPPbw5q2/mQNVQB2Vjr46NI2hP3xI4lTo6F+x9f+nHNDWYxXBElZUc/
2rxk0wxFf7F1eyIBrSqjPLj/+Y9hJ/cslyri5AD9mVxt7iySGyoGwwhVj29S2dNS
1yufk3ZlyqOlHjCJaqDCKRGdlCcJgRrvqJdkAcg1UKxW7DlP3RXYwlVkoxim2O2A
WDDbK2vsFUWyJE+HleuqoSR5kbwTjWb9+QKVFZ7LPe3V8pJD3U55HA9uWvfgrG20
LWR0HT1ObqFvNXX0aqRgPmaylCqEJqNHl3eYFrppTdj2Dh7PU+c2uFXn4ZxbiQcs
YGvXU5dU1yuVSZI/1NdtlitVt6/t6U2MCWvl4b/+SVK2Ex8pmrWOfkM163TrummS
gRUWjWUf5daccQYm9renjj9/Bu2BeH/fr+6pFCRZLB3A7yIV+D17+8wvu5agpJW5
WU/C1FsuMDjkE81gozjLJbpaVY5gj2A2Y6dBWjWG16SJEcrW9k8bA9Ym+r7P/MgF
nyS/ta1bT/jWjnqnnCggFyaJ0L3UjiIAhuqTZFMZAUwb/MUBK0tGKSsJ1Br4hHU6
IEcrtX+G5zp5Rw9eBk0BG2xt2YZJiRxIaYyv0U/y6BW7Qn1ioCkZTWvsifXfMARv
sGrX5/RdFZzgKwtmZ/1x06vNsOe7VUWK6IgTJGdD9m19TZ/vOv+Q80QbGM+KFSN+
r80qhUmi7iv0qe1ywtfPZhHMuREYB1HZHJoOPGQykWrh2ghHJGcpZwzmIq9JkirH
D3AHXDiLDVglxjMH+ab0H2FsqyMAKKCsZ8s68VEAVh0SyLXti4p0O0hel2fB/bpk
h2JzVajBl/hl76+8epUkH5NpOWQ3I61zCLFX6aj8R6BqxFmrR8UCFN3qf1LPc943
7N7kiEu7Qi2l/z/FAbpxE48bvBXbpRPKsEYw4rJKx1S9djt3YpP0hh3lEab2w5On
dcRfPq2lfL3cgoIl1uCqYiTcCJkcQDlEXq+6sGVbCjHbVgsuk7Y9a9kPlvK1GTSg
rzQmzC+4/TsLeBwFs4pvVkfRveKGg6OL0bkodtgQ2sCDYTZ8oOXfYwB994bJOiOh
om8nNaDHqaHZbaVoSLNgl4m942L+Po/cqbo/iYjpYKU28oLxrDHYK59U7XhOBqCX
pk9gS7h0r/i3imSmuPcHCpdszW/xUmnJiqox+oIBqfTNLsNk8xWuZtgIA2LObBRM
bPv0KroIqctoqsprh8XPekCwow5+VamxLkN2Qd4vxctkC12o1XCeTGDSxQvccnbM
LIDyfXFEzBa8/5khpoT6//ZGKPKWaMPPrlUrQZ7pKdgg7oDsYkTFSlwIYq+/H/r5
FfFJ5qbDrmCKeNyIjcVptiS4rOZrVfhVgDQsc0pIeeuP23rdnan1V7zfO4IjmaRh
wF5Dw0O4fB3DdYpXiUbGvz6HqZF/WR5cTulG7uoTJzkive7EwjOwqU0ob5drkSPe
NdJJa03BalFvtqrfGJQxzr5+hERfBBO9NwWm9arhWGxq6bsdJjtN4zT/yzT4WOq4
aJ2Az0/5O3OU7x0ZUxYS6wjL5/YvbmfcXzjSacSttDJOGQamDjA/z0CU98Ao5nI9
HjgD4hd3482JtV1g6utCfp4uRGysGJczetAhnwnQ0owo5+mQhXFh4zZj6EYTbHaH
HVK6ppnpzE4ZVP8s2q9loo3orMT5vna8nMSyizT2rijcEn+cOui6K7wWr8WiEydf
R7KAvpyE3Ek47Csjpv9J0pQxsYKKG2KqLvmJVGugcDh+IavnGVtbPkH6JcR7w1yV
86Gwss7Yx598E1XuFjz0RdwahPIKkmfds3Aq+BGeh4HMuMpw/v8DRQN+nhylc8D8
12WmT8ZA8tT1NWivrdKy6USaxyDNsbPO42qTN10H4MCQC0NHBqnVprFhqqoJI49+
HoeRShzzDySy0pgMORgvZlhO7sfLTHcKOOlDeDCQneaY+x6yEUlhAnisf+bpQvsD
+k211OnYgWB4RAb6bKH1u44VMtH7EtxqTyH4jDAKjxKkqvU1sJQjXEtYfEqzmAOT
AZDXO94hzhfI0CfIe2nYIjlOdcS00gmj3c9lekRG62Q4o3NdT37UvMIX9P4D2I5k
ZpbYGQdq5oa924AokPnRCPAlqwnGEX0m2vvVw4QQWYArvVAZfaJfdlxSb4X4E4AO
1cSsLKKHThRnzSRmmMxBtGOssNQGCeDCtAXtz3/BYq24bjyunx5wI6Ebt3LTSGCd
ZC1AuJtS0UDf5gdsfrrkTDSBQL1uWb01bnfSdYnWhYN5dcPOu3sB/3MwXv9ctsWa
MFGb0xYM1+KKBOQCr39Cf/3C5FCJIgqUKf4zDsHBIICatudYG7ilAtu0fnWsi3N4
GaPSj/jEneAyX8onwBPB1ZYNgaqJUQo5yfN+WToGcIKa20KqtI4V81IzAr+pTm38
0w8SPKw4sV/BLakvBC7S2ZVkqPg8dQIxbLL6uNeuxo37ipegazdGrfBjcQZ9DbyM
7qgc3/k6suj/cfPIBNyL3Z0G9fSqwNnNtvhR2yXvqbw4XMt3L3E1iHW3JJNqeWKq
AUNCtroqxTdb/g5W6oQ1Hq+I4koNnHGtLEMh5jRy0Ux7L2FbViJQZ2Q/H2YNU1/v
1yjkl4myiK4NZW/jRLcBxfrnadoOHjg5sW6z6+uJCpItmCMxSlPGcArr0W8GhzbY
kVBhCPBarvLjEPvEXv9MbH5CwnVjQI0FQSphiMTsjDXMu7AIEEKHVm4kCZcdiClm
WiOASeS9y01n5DDonW+ip9oRyJijGaN3557wT42InaH+wGlfzFYYFcwy/12rO9ps
e948QpyrzDuaovA71iVWQfmXDy+ToKzID7zdtZXvT8Lxc+E0Z2yJsLluekec6g0v
UKMBweS+98BZZQMiNRHoqnpJXyUbZH2WYOrbVbebjitaHOMEOTYzV92BPZzW4IR6
R1EL8t3DgrJsG93hnFN3iujgdZnq1RXVUVpEH2hv5DS5jakQKKie4giKBXPl2eSU
GydpnPGddjYumSCsakC7OXl11JpvuyhJ/SzVDWYTVl6SQoAlPKE3Hbg3EIFZQ0oW
63Jm8gFDpkrlyhaBjjltmJO+xQPTC2tBkZkyTRxOj4+whzPKYaQCf68WfNcmcC4u
Oipx5C0raXWpjSJ2rBwyUrcNDtIkNyQFvWp438frqfEwJHqx3NgldI7StIgKpX9l
OsE68dMHDlBRU/whtH2II8AMgvfoeaFW7ayq/QGQ4ZJAACNeOdjw03K/SGaB7Ddb
Z36cla/ACHDhBNUyrDtCpdZt8bso9YKUcOP3FKLaPEy/pmliAGCEOsnz81/jxjsa
j6M7oSMfrGWI6WaGQFgVxAxVr6Ptt+JdMkgo8xYwhCmuZrfoEUfWzRB6ZsZopYye
k+ncm7uXHfoWHOeXZSvRn/gtacnDqTHjcKemKbJWGZcLj/IZz2+bmqKtOpdypinv
psp7iEmODggrdXMVqBi2gYFhJlGsZhUoOh6vbCR+ttMsBiq29RxjKCt1icp2szZn
fzV+40N5Pck+5gaW08hkKzKTDNfCDWkVvMCWEwYrOqeLE3+lcGN1Y3NUac78WfBc
wxPRWx6cCnhSeOn8l5jl04gzkufwcbJiLBNnmyAk27lO9WIsr457IYRRYaMUqzyr
A5qcehK8UScr+qk79+eCZGDr7f+K2F4d79oFjiqIpmtAciSGOmaVgLChzuNtb2Zd
At9o26Y9+ut2Gzx9ennNcgZ67SBC5wjWOcIWLdq+sMHpfl8hhqXMRDhVMcSRo/bh
JK2JCHUCYIpNszKmo2z5xQZr7Bg8M9xjAWFkKMnahdqCZ+INqvx4vzaG9P2XfNj4
WKMUouRWo8EcHlqnlktQY5SdnGcshae+JrXq12GhXqVODVPxbKHH5Yr7XmHMExD+
YB1jYbXvgZk8cCJoHoRNuQXVVvcM79ZA3Hd8f9BPGhbDgWg0VVL+37O61My8I0Sa
B0yz22OUNgkNt72DujGiDoMcj9jvgStJGv2epsX3QaQZDKL9OQhKKApRPIQ+LJLf
2hen+4U+DBzCa1dqNvTTmS/ZIvbYVp9D3CA+y/RAGPDuI5l7ct/wBFXsdqFK0o3B
Azv3MLYMqw5l1nHcXNcdS1zGqp2lRMHbuO5aLOxR09PyKqYgRTskuETbSZE5knYX
e8PCcs4ADEPw3x4TqN1UZRtpGeAKN/uHIpUKDlBdWsC14xOiHviPMcZnw/k3Fndj
WwFNyXcmEa0URLiXw1SiU6EtJQTeNpZfFac/umK/WqGEWHcLW1VqOhe9iTpMiOLi
03yv1iZa4b8wyHTc21rmxizGeR0pdOgd8c3jeNps7mqMCnKFi0Mb+fu9bPmoQIzu
Ohw7fQaBCtQrnFpKMhW5kshBZGERcWgAfPug215nlX4JSDFPV6bfcZ5YNpNlVWrc
4hmBVPOJwTPb0W7NH7/oj2VVTwyw6jeiNMQNoVZIOvjLXRhYcw4RxG3bdY7mal+1
fcdjR7LWMeoxbJCDFAHWU9S8hzxCpxgA9l5YDryDgzoXhwNynIdn02ZvjBi5ufnY
P1QgUG8rnV9I78o6BY0yUmr1RJ4U9CaGa1zk/wIC2KsSqnpyaRgyOjdILlehQnIW
gAthqj4iIrek/l6Tk+G9ZDZfDWrhooQGn+XOaT8tY1lbISNJ5n1zjrHvgslydFFK
A2c3fbR3r6EO5kVbvWzYQdhaOMM2Bae9xNiZZjQuzIw8appIuEdWKYeCJFWf1rs9
OXrU/bI3dyqGtgscGdmp+xxw6BbIjDnBUC3ECVfLOPt4nHL5M3qOXwY9lJafMREk
mKtZ8SaBfdl7rtRcsR1m45adkkACiRL6dZPzLmcjFUMHebKGZVhDiX9VJ2Od0SRW
NAZTqwe1vk1MNdMSAIJCDwPr4rHqwe4eKyfs/0Wvz8rVAfYG/oqVyrxt8TGO2dkK
BCLzVvDDgaci28OX0R75uL6Z6n5+LRQ69hihIrgrL9O8enCpZEBigOJBz80NWCL1
x4GBPBFOn4CcRS/3X+TdpOy1ac3JQpdo4g7G6QS3ElGH5aiAxVYbN+DhD7Z5dXt4
U6gWkwXLynyqsuKruCYHr9EOREauFA4Raqumz/DoSVUd0U2MRQZU+fFV+dkwxR33
Rj2iAWzwXtRX1l6/BqqMVNrI5ZHsQTISz/LRKG53o3F6wySJnYs0jNwF3ua1lwDi
ePH/zRtwUtQ92w/rDEIrbni/I1qpHAw+88EUbAPR8qajBIrReyXzeEa/8kjkKcTT
1owNXhcXsKFCt1FPt/Iudo3M3podDBa5/Ik+yzTgCzKHNIhFiVnQiBDX8PgmebAQ
ctKrBLeSj8kgvw/OdI/rgfxcYkGY95l7QUMEjPgJmmtq5v6zwwy0p9TRL6gpxQis
D+ux7zNdDkUJ+fjqBvlPxJDjYZ1S0lHeaxxsqCngQRcJE24MYP6T6IKC6wfc7nOR
n4sbHJebXD+Db/dIDQQCG3YxaMlpaYWPz4AUlgSMx/Izq8a6Kytw93/RV7/PHXHH
jU10YdonOFpEQc+TLaKVyOAkBhpYzxTA8hfSeB7fJlvDuwk1SBDSyvV6jAo1M06h
1D6T2kcFbSwdPJmWAUK+leayJNdFJojw/rrDOWiYJnrTWhspuNkeR/prkuDSZWwN
eRpnEVk6gQUyoLsrut8dwceBl+m1roOpEKn8OYuyUZLSc/JHidNsfXygnK2b5aYp
2Fn8/4IpBQ7NY/3dEdS5Piq3e1cz4KDPOe7g8DfGlGdH2YQ5TdOI6Os55szJr8Sq
CIhr4qEbUW8YjOzz/M38892HhC9hp65PI7bjZSK/nb85kCLoTR1EZErFMPBiMegf
IK9xrN2G1EGlfCJR/mbdY2Zo6N+VpL6b+5rpggII9yG7y06fKDCPtlvxmQZmNU7N
NUzoTDwLPAATkf79TLt74Q+46a45fMgUXl0HBMZ2gXsTOYT/Wn2mn20M4Sm8fwmN
gVeSs04yrCCJlFaMkAwPp4qTOfG1TCH7Ktmu8p0En1QtsNmYM1ZWqLzGyZ1wCGKz
8xHCog9cvsdxshwa1t4Awn4oPWxdTdhD+WFv8rcUWsfm3IpRT69Sz2GMPEN715Y0
n0IuBEEXkfQhIiW/oTqYgkkYjzS1vwNU+P+u4bQvqaoANulkFFymyu8pKcx2AlOS
SMFu4Ur8e7pe722gSBDhGUUyLh5+Qr8loAELKwoNN8gBRVEwAPboYf3etzkC0b6E
9ybuQeRq77VWgDrIWZFXpwbonydWdqOgqIerWHafHj/MxIMGwKgoYFCQEnsX+8/N
r7J07dSAQSJWk2pvTcfdM/R8E0ARRj6plf/il3jvw4S72QLmiLgT8NDn8kM+SeJY
e9pmX83pCPi0jD72FslmVDnVDKR6hVVOD+RYQQP2QrvDPo1nI/kGIUxDXSfnC5TX
8WB/knIty13J72nD5eOEtoWg6T02Th1Ju4wV7CVphzYnIfbk/8KV6k0KIgsDTKgH
p+G8P2S/QBZiRY0jWr7E2XkgV1Re2LgpMxz0L9OTtolT2JsCJXDZvHTMSJwACmgT
58ohHbyLt/Dg/tUL4DCQKFpr/DqCuliTUUgX1GvR/Nc6o+UK81max5VXXcOLka8X
2mQ/vF881ef9dJ3jybIu6FPJAay1m+YlF78ZWcM+hFOTdQmfUHYBVYNkuB2AMzVy
Nv4t/LeXYkfVkUoyE1itWsPhu9z2ofGFFcONvXoeg80Rug0EMmzlJheWX3uJBXti
kRVNl23xK7Z0URqaJgHZt8TwrchYQJLCVJUtqsy+iB/2D2wqIJ0xlSlN5gsz7/4U
ua39sI5OlqApk1zWG0UhEX7VkkVpaEYzECMhT3vzUHmk+VRmCqt0cQIG9YYORsWI
3hIpxqkOvlLnS6G8l4g7Cyr4TjBjtqFGmwiKqIHELMfV4YiVa3FZKtzoiWeocYpK
mYOpzccfhNupsUSzlSMM0ysG79HFaR9LgArFXU/avkKY29tkcFm4IOrSAMkqw9L0
2/8xRnCOp83LtJSb4kAQPIBVMZY0VmDm8NFu9z2ZZJcqppFiGMcQk+ZtKk7vgyDE
iO++YECL4OZJHq+Wsm3T9L9oqCwAMaWPI54t+PDaMFtri8WtKsnEGdfRK7tG0sus
4Si2PJ30xtqi5fHl6bb6rtidH0Y62RK0aWfHU4WEFcevr4+5YXvimQLYCeHVDoh2
QBrWRAEgUSlXMtE44tgRi3ZbnLQAxwDeibGLpsHKPu0c/IABKQTzXjUWJgokbYIr
tX58vYdEPV/UXRW5E8TbEIH1vydtNg4iD/hMfioTCvucILrLE+nBSYo6vXbxJ/jH
WDbGD2Pf6Rn0LZxziXQbkC+9HSlBKALj2q1Bj4rUGOeGnRchD+t+rhj2Vxibll/E
FIet15vr7xkpv8HuXYVv8uL9+BoJjThNDQcuZqkINQqZmpADw6omKdTYJ9eqMl/N
Vkpc+I+VeLhnkE6ic1Svwpmflh92YqC5+5TQoPsROs6QYd/peMb1kVaw0BEJY+fi
UwFo8K0K45KYpwxz8+kSQPyeHFp0xoMgj8IaB4l+X22RyxTSQmpwwOROFNcTdVWL
heIiq74FrInkP6FbsSwh7mUn0WdhjiaDPUtAd9LeRI1RX7eaZrvMDmbWwLQfuph1
YpyTVHJZDOqch1Ci6ET3W17Y5XaHngFIU0M4Gth1ZMVNA+Skr1Mwk5mkCvAXXKGG
BSzN8ptM3CYbE7JxDoQ6dUCRzysbelaGUSRBMz5jxfxR7VWmAI0MuIYksnveMcqz
wm8ePfDFTQPdyyHgm4g/pgZYleFtbm/ZHGTZY++x1ckA2pEY5saIIfxpTUEyNywN
f0T6UVtUZ9ivnpz0IsQd85ZCZ3CoYkD4El1jsxhWa/xdn/MDpDeMmcfjzOiKuI9s
3sv8qJgmjNCrKcoJSof5ApQCnFDZTFiriCaTizACA6zdbonHrt6mJmk60i77tD0W
bnk9ZXfpNdup2WXVLjc6rF0kFC9Gun/TXbLi6ZjFlYWx6dix+tq+DSd17IAc0wzE
tUe6Q0Y354c4u9P1N5+B0qVPm6D2xiBxoP/sqxQd9icTruzTZbS9PkA3Dg2ye6AM
d2Kx0/iJBPYzVg0h9qswhZT/zLRsvhBSJ3URbEbJGWxPuQuxGoPTM0K1uk6FistJ
09f+va/Q5i//lE0YvGpXpHC0NeuzYTvpzwU6sPLPbWigFpbZ0yt0xFEG4GB3Q/oj
+TcNbrRJ+nT9qkKj07Yz1cPf9sfd7/tAuYGiVmysk4rKfqAxYoA6PNVgAFxxxhNt
YjPsg+LahPlcZ4E/qzNeL2S088LekWFjkRPyjqTM5kbOIgXnSdqQNqr7ckYD2SzB
tMuodLzvFS4zaPvdO9vYP+2sUgA0icz5VT3LezJBZfG97v8SdDoaH8+49rrE2iSm
F4rwhXiNXF6Qn9mZH0HFv6/cgGMrwq2k8CrgCRyKkOInbyV+LFG8UIvCktLRe/zH
SvphWDwMyqqqYY0bjkXIG+Caw8Ya8DclaG5Pm8ZwKTlqMNWYk1PnPbSCx5DPJsVx
mM9BqskwuFxSc9tER2LIBO3uFTFj5VvFLsEUxz9UXfNYDRDw+uysGY85c47uV3BU
KNDjJgMWgFSm2O+cXs07KVxvDQ82dXmO1jsxmDS3nM5RmQ7TxVTwFZf4EPvqEWzq
CysQ3yLh0w1b08pNUyQ8RKq3ThszJkSbxlANPZLTX1AxGj3hWbAg04iNb9Oa15Nr
gsqNnLSyF5RznxcrE9P6r5/m9jBp909cMhi4uWvEKamgW6yE7vhONEG/oqTZK+JW
qhhkfVGC5z1MSyfUjLz9KouEfUhVhb6WY22Kr2gW7Kw6387dhC2FygY8Gw9CrcI/
Txk0M8C9KdPDOWkbfOJSeBpP0yFeLtpHV6pNaJozVfSDrKTmJyi4okDAohMHscFF
vItERhHliy9+kqZ+Nq3y4SZztEmuA53c8yCWIk+7GsTwC8keVElYJ3LShjqAs6SB
54hEhndy2EUHkbErRJ6p6e27vxIfz34ui4mKaBKVS89B7qIqW2M4zojvMX8FQcF7
IrDCd+r7yM+8cHnZRWxjEA5uA5WWiICRmcGOsPEa9zCrHUeWLcTRXRXI06x9Wc8x
1Q6rGXoKLMYXToeZRxJXjjWGTCbb2tSBSMGdUbr1uobiQDubAln6iRcoTk3kej4V
pRhAr/2EcHoAI8i5U62iTc9hxtI3EeUhL5nr0HToA1q1qlLjTxDQU+nf2q+ihQc9
H8C6Ti0wAZyroWOQz4jg2eCDouqPAWQevDrJ2zbaHqk408myjj/H7YWcEf+v91pZ
yjbybhaB96FD7o70qlBQKizPtpjSncLGOMnOi6pEn7UzT30TEYqcLx/2O07aCJd9
Q3LrdzhpbmCEmBsoc9pzhPBy4vW3wzwuxjnCoDjkasjueGGGLXDBl15qU94/iD57
V6/mdCmHYE6leG7/30MBD1FVuORqpKCFoIEJbcqWFqvKw2XVEOnZECdb9lWLC0fl
NF38cL7iKd/dP5eVdW4XK6QdkybIN2SFo8f870h1223SuG1MI0VW7CT7CDJTU4ol
V7dxELkYwkmZruTmBJEOXM7ntgUi5GCUOMeI2c57dh+wt9MkO3kJVmE8aWDNDnUs
XYpx0kyaPs0uAiuJjzquvyssAnKT+wPUj8bxPl6wePUPamCA/76l+Z5ebmw23GSe
moXhl2f47Q1pngT+s5KjdhUTuYHaSjlqB/IcXIiKNFg1YIbd4EwhBzkqR8/n6dY5
k4A4nb72T12FusPtuUubg458er7XbCp+rGQD4+vRbhOFudmzN2Lf7s0rj3Y4yrKu
L06awZ9Q5hQLKGYFg1UbZ76sHrytef+ib3jeDBbs5QM/IPBKE/8mWxd5e2FfTiyv
gPwv6mPPkmUUSH9y71pwQbhrJLmClJv9WwfYtv7UvpYLEytzsnLSfgA1wtSLukV5
u9hphiR0hXRNrQxke7wEcJOUB9WxReYtEy2nik2itX2/0u90vnCm1E+eD9nKZx62
jFa66NFcrI4cYLMxH8Yr7cth/wQh+MEQH9RMBmqBsqwAGCJE/ncswkrFoOgX7xyz
9DdlaLzKUSjurlSJXJkbmYkRicwflFATMzH47qaIAt9+i6IqNwrscSjP88Xu0cxD
9anpLg9xUYjvV8/taiTc6hQ75Ubdi/uIrFxL8sVb1xFqptigxgSbqQMCoH+1lY1Q
oyH1EUt8WJF7ULnWTLqSRh93nGYcotheqriL2TKZWTYtf/iHe1VjLbJ9va/Toa11
JHGw24DedChHXco8uoo9p9/7rNTkXBPt7YXvKN1BcBf+AfDF+61yFt7pfZOhbDFq
odoXVUztQXNa2WerwgpCm3b4kZcY1VhQygzjECK931hrX31mGNEXganreokUBc67
27sMM7c7mdoiPf7bVALsDDVb3qNXQJ/ZnkUlcmI4lSMDfG/BLF1eHlX90IHsQFyU
QeTK3+AuXhXPsKJl6ekfuOS14MUt8m+Qx87n2/DmqVts0jszSJiRXpk/awQDeraQ
GD2XxUm5Rzfp5S7jAU141ydcztAifWOQSd5Bk7CE8aL4oRfPWfdSw8Et4XKuPJoX
wBpj8TQwyPt8fFx7E4lt7NEoMJlMZkJY0N70RUpssO3inbPaEp9W8XxoWinXK+Mk
EI8h2jtdr0bsi3U4OvtsY1POfgrd+XCDlAGs6Q2j3LjgKlDD7RdjZHRDAkEldLX3
T/sx7blT/yEpiC0Le2CY7utbQRgYGUo7G+v3UAwME6ULiLktJN43l8XnAoU5BbOB
xoSrGIgRFu2QU2663yawc7M1Zsdte1N7uCLo9WUt9TbHqJhGSBU7qV5o8Zadd1o5
7mwHo6tXSM1hKjuoB9Ag25ICmgzXYCMDE7pVD0E3UnEvUD6oW+bMTClUE07yGxCR
WctJ0StF0ertsfQY/HcF5hajgL5oxzyq3lH0MiUId6NTPzhea0Ybx5C1IRm7YaK3
eFLZxyz8jsiOQRzC9MKZMUQ3AnRgfgKg2SWWTmOoLKNW4+XHVDVsriHyES7selFI
EdZFtYhRfdUk8B2j76pKIab0SggXrVNRNHxg5rCHIx1puz6/Pu5xODxgR3UL2M+V
boV26dqp9aySmTgC6TsQoc9PpeeYPcheGjQFlG7FVNWgkKjGEpWGpzVA13CTv8ek
RjObJjRGu2dJCbeKEib2SV0aWgpYHpe8B0v7Bk3MbnU3+m+TI6OBmXskjbEDZsG3
OOBT86l9yThpu2kMLXMiow55DGWc4mAa2WiCVU+LZznbsFUnppmMpIRYffWNVEXL
jiiKdwk47kOG5eVNLxHwES+9QaRTKNFKuNk77bJEqVYgUFr3Hh7kMl+H8wsUh92h
5KZ+/F5NsVrXpPbsqbanoS/YIlup1YhyW3rxgV4HWgUjk2y6do0MLduNUBncFSY9
Mvi/Y6Gkp/DvPsrtAUe7LDPJ72b62ND0YbRXBZI8Xy6ed3opRGkm5U9JlwJMTPwN
SGTQeYeEJPT2vt6nLKWUVCI6OwlJfASTv4Ic4J2ogVvjJY7R/jwcAdVV71WyvBrX
e2L8HrospXZPZI7pTpf4yJOrnPZGojtnr7rY1MIae8z9dBvokJPmPOjSOkQe3CoH
WBDO4EeJS6LptC4sWHQDKy6Rj1Ov9MKpPyNGgzNnWco8RY7F/FUVitdOLVvphpOz
0rX95XywUVBAt032jsbufVHE+puT1H6cUQdXAZKmcCCl2SKyh9p5cFRXiYFYwFbk
1CN3nGD8cNdv0ryEgbfQ40rj/mMb74NbTP7pnDInIIXRyA2BauhERtA9Z6wfvCuD
b/CzrgtPErtTVaRKvKq/i3pJzh8UBORtPb2CsXy9lEtAuG+G2X2JHyMJB6VcRGx6
N9/gSwtpeyIdPc03lp68tNLe6SRwHCqwc+9K44KAPkvSjx/3tJS8xANesnWopj0Z
UcZrS6h2ouKQcQQFq7hLY1uEyWTsincx7wQXpigTcdRC4V77DrZyeeYoPC8eHZpC
T7GFCCgLhlFyagGkkfnZfzyAMREJRKKg7vJIMz5t7ebpBl3y/PMIfJKtlF8pDGQj
cZp05g4urSRM1xWLGLlN24yfHMu53VPfWXR8s9vTEI8KNPziAUQd1MtPfOnczl9c
kk0ke8FQWOTeZDXVF1naSCbvaDJyM03/0725JunkSXEfkgkDnI3buzI31GmnFwp2
+Wb5mHE3pT4G46hg9wbTxb3yfy4tsNSGDnFFlG4s0vx3ZF5XCqtAjA3yOO09Dz8P
M6B74KQgD0R5VcgZtsUVvAzDh10Yhehk3eHQW8zCCboeE9NmZnQtvy8wH+qwCRZF
Fd7KANI6jbDXsmlIt10Xyzy4GYlW5dPw7f2nT0aV+00sOHRMIXsUK+qgxmFKx8Bp
yVDsN0HPGQMJyzM6mJ4oHIWJVXOn4x5wDiroTPdNQVgItNP6PlfraOCi+bObi8ir
/DnszMCMyQPBpDxrtTc+l61zXeQSDdcVku/CNWHZwMoO15nHMARTMEIpR1EjzA/P
SzDYS725G1hD10g9IK/vnNUz13lUJwikK3sZN1e4mmaEbeG8rKzkMbIp3t8PzRxJ
P2kEhJtC8OezRau/JW6o70E+cURs+TG4MitgKLS0CxHIswHvj8N/L7DeDznqqEMZ
gJcydwBzKhzAws1vRavo9Ab8i3T/RM9eI/UZHkaOBcqnN+urTJ3Zvu4L5gjep2wM
CTzBXlAfXMyKTnu4Bi9AtgoTcZzcaL+d/hknvnpuvfPEjqUN1CAsVhxagXgCFN8n
uccMqb4UkOUwn21iFo9h9bk3rZXZxBhIkCNO5V15aYPAA6sFYpKuGH0vjFvXb9Yu
PNXZLlfCZ2kJyScXTNvXhpGjZRnsbVzCBdStDi5zMlh853vAaTgCcJurgtM+NAIN
8w/dlAVI6YIR/RtKxOVLL80CKxim675+xSPiCUvCEw9UXs2o7De6Pp+nhvdPkxEk
tT0Be99sEqOvjkxoexzY2ecrZMaWzjyt5xJwWT/pcXSEK4Z22qV7XqMY6lDPyNVu
hppSqNMvmKxPR+SI8atvZcdXDN3lfLbmlzMTNe4SROdwYCKwZSBb0TSvgveoci9t
mDDUC++aNAu0ppnCMJkckCR9F6bJjcxz/uBvSXPNU5+sdB7BNbgbGZQwz0AdlpvU
DZBbjAyYhrLlX0+itYyhY8BTKg2s6JTKKV4ewwBn/3bQenMT7bySwpHgQjhOR4Nt
Cc1wWOpI+jsaawzHt0WA/lUPPIybtckBC+HAnn1Hn8UPvcoh+XVgKuf2IGiLfASc
zr9VzTRWEVzVcEqNDc9fajlsi+fcR9Emv2vfMRsJkShiYt8qKtABFblxwkmGmldb
RrcixCxAcSv4zzKdas1wPW1gqKAdktJCeQ+6ZJ1Gbk1NMvepdnHcV0KoEZk1C64n
MSFyJbJxE8zgw9/iG92wqHX3Jwjc8LD4GnhMjZXeYkgQwIbgWiOEtde7/s/ryiwt
dW0N6krxmd2oNHJI5kuvqxanyBwRMmnwQq+e3AuFvOirTobyCVBcGHpjEl5cJbsl
AmL0BJgW3y9nH5MIaafsXjI0tYafA4kYq35R9OBYk/Jbwht94ZTh7u4Ofuw8Khs4
zN/RNgXx9fNoYtRdijBK09YMmg12E712KrCWmHgVsxpE3Mt+2TZXkmFV0ePtc7C5
sMOODi1U1HcX0mzM2B/Xsa70UN5TXcxzL3ww4chSY7I+8zHCYPV3av6q1xDXIdR8
b0TtfOC5hooxwjma4ErV6/VbPhDqiaTwFlquymECJwsW5+jNfWIGy/1dCqBXQ8wt
x8v261gVmTBsugA2LFzi/yHwmY5MaET3R2pt9qrnFAiefne9iNJ//a7TAZ8Kt8ta
r0ZWu6767lkUyMEGwbgkY0djwecEKv0xSVvMUzyDPqmiv2f4fJ5+q0qrHPX5fg/X
C/C4+gukvaXVLuZPmxfjpyQHWxKDuh8xsKo5pf0SCEsaojMY0NpIIohsrjOu0cGv
hmsL3o7P1bj63J/IHP6jgUWZlz3+GvlotCYlg3a18PYcABWlarBa067iVvLf8Eo/
zqyLa0+riAVC+1tImbMqYqGyh2uLZDxDsVOiD9vNpRyrjsxcf0v5QHmDuCS4o7yw
l8DdqE4WSZK2RQ+Z2xGed0bLe2TitoWPREkYlV8b9YajJxLw2XGjzn9IqWs69AAk
32ebLxNTxaGpgRFd/wlSUrFV2LG2wVr3KlVOqEmQQi/yRuLN8JobSz0DE2ehD8HM
S0nNvNBsH4vxjOzgDBU/am5NTiZRlnhUrXSzKncYrzzbRmdvogXRWJGxAIGHahfi
wbkG0Nwv9bJ1/CorBwQY7VycF+kFoh91JsTxdUxQvbE77mZedo1ZYwUMdtfGnbkB
VD8YlqJoLLIymkb3iBekcsbu7t8yXPfVFZZVZJk6pQnxKRtqsmacPsQooUib25jV
Ezr2yF9OsdjbUe55uwH7YYB5dva7Qp9RFVU+sdTnCwcn4R80XIZoAAlPc+20dUAJ
MmjT8oI5ihStIhB5Ezz/eYB7AtIjx768JrwsWNZwwW2bomAFNE/7Dk+N3dEQqqm7
huXYVUu2HgXgLnBvdqTFrs38ktBsk2PoPN2YraQkVomJV1KI9h9QcD1/aubORCFm
n8gZvaFt6hZqLgNm15gRbj1WBxl36n4UxYyKcZ3LYJmXFxree/D7lv+XpDj3ydxC
EU6TqFL3QI5QxTybwMJicoPck1QcuIPbja9+VBcn2GV1ottA+H7Mzu7tcpakv4HZ
iniSvFRGvv2bSQQyXiDYjTgVC5/DieufKihBXKOHt2mPL9nN9sovsCgYe5RSdCMd
5BDLjIwqqA9kh4JLhlJ9QQlcDEhRvZSEHA0jZOoOAi+LZGJxtvgYx/vaRMsCsIYR
1lu6mjDWWwh0YcNQEnkKJg7p99COvw19ShjVfiJ+lKuTVOOfPZNI4zyjEUyAts4N
UBmkUo97KpOZpsJOHtivzeE4aL7j3A0HVoLkUp+ax6VR1jToKJsHWWohF3/7HxN6
ofS4dlA3/trhybi5b8WpF6VjbFd+ifNZ8qExpVatDBsHqhd2yJo9VIxMbSAv2K1p
Z0ExHkDXtxxsKhCEDewLKLyO8S7WlhNTZo+h+8NmpkLn9Gr2/0W+/QqqWF27Eu2s
GYMBWMBNUwpB3FA6ZA/1O800k2Xx/kjUN+/76NxCbohXy3bawdhdLQufAsd7uXR4
ae1EefF5ZB3gpGRhBGwZCLY7h6HmelgvOqJO0Z89QV689evF8XMrQJtSWVThzFRv
QxbxojOm4m8KZywI5R6DZIORYgIgtHwtsxAnw1YL1vOFv4rtaqCFjACGC2QFq1xx
6pTYHNIgW3GcaRK4kVjNYwnzZRBNyXph+EAvx9KgWUgWXQdBVxIHdcLgGIEk+P/+
dNllxwW/1LQFdqXDgggnB8W5Xh1ld5ToEQa3eNgB8GLWV4H4KLiJYePhStmWZcd1
RLEAZBjpxdbZqdHvgF6yZ0dVuiH+WnLU1s7Wlpl93WIIgFYNC06PdI4rqBPbGCja
dBJNhEt/cTf3ln5eQlyy+63qQBdtmeXM9RxwmuYNaGO+svHiu3NFiEChtkPK6t9C
GtY7QI2TTgt1GMAK7zk2Qv0e3VfMet75d2Vnqfw1x6IHitS09MB+JbzPozwPdaE6
7GC3oNfLBgsU+6Ku/669c6AB+hkUTfgbBQr4Q3vXAywe9I3p42vTWK14ig5Jdv+i
jQ2DPiCq35dGkdqcAniOKOIbwfXNobZN+gcEd0mT5sUBey9zifVxMHij3juuWuED
CE2OrVCh87D6rJQ3kW2appFemV9eiIiMw7zLKIHQjNH4yedUKO1Wuap3VY6CTGil
iiwe8veuvPH+q/vjYKbpq50BN3MCfAtXLIptDtjH02DSWMJDLdIsOipOK0HCKlLe
QuE1ycsYlCiWlsSR+l+HSiHH7do0Wk8+qR83A/xJseXPLQ0lUKPbTCjMSUSNIXeQ
wzkvFyR3fF0Rm6B+2JJ6iCOaSz4NuDdHk0GvgoqMvvwkvtUC1uggFnsfq6N5HFCV
GED0dzhdhHDLRH1EqPhmzlhJMvz13+onRP/TO4SA0qVe8gnB0qeFBQLrXMjvcwoi
GMJJ3DohVY3JvtV9+YJBJs0XGUoY4eFhyQ5VmYnxzjeKacQEY1qQ744Xc4NViURk
XNM1xYH0OPSWYzhiSihPNZx/2sV2gZAK8ekUkRKB9fKLxUlyUMRjbqh4gL0GrQ0H
GzHPyFnptgRCOCniJdkEOtssQSAxj2Nq+vLZQ8g2brax2+a07XBMaaRDA71ier/5
VZl6yqJy/Ru641qVG1Dt6ZBRTSJWcUHWoxo12stBDL03CVSRHLJZVa9oPuQp0WRO
lPY78ChPwBat6gT2hFaL0NBRyxeUgaxIAVCYwDnsz9SX4eugx/C1Z9hjrb+DnGZ4
/MsOHDeOL0P1qJLWWsoq/xCsA00klakP21Q2AdhHWSFzMgO473sZRh27rSjePShd
LrNjnuyB2hG1azRBpc9wkfVD0h4qfyyeDMrGfaFf7VYy/98dIacwq2XQvxziNC0V
GP58VjxuM9aGZnz7gNWqteS163AWdiyJdZYCH6kdhS9Bh9bAq9YmfhNYo6F/ED0J
3vcgPes/J0HnU++2fL0LHpddPEijNEEu82+bsqs6pY2ZieFGvLuzVfAJ9GB2NZ/d
9r2KIBiRqC1sBBGGljsOOWS4o1KjkNTa8MojOZUrV9b3zlI1wcmcoxHq0NmylRUZ
2ZcHvNBi6kZ+bGNqh5ddmCvm6BtOaBlJtBe2qfSgP0UE2ZX3UgjVOCUh9XsgqP+t
C3kxUayt23yFHW2wSP/eFSa7LSyQjgoAFv2ur0YAes8vgSMY5xUKMgSWl4aWKz7J
gWkuaK2CGm0WOQkHzPFgBxGSLLvbFlpuPQ20RHPNWLOHyTxFdVEF4wbh2j1/OlhW
Us69PVTUWDx7HEKufbpgTXzw85m1+XPqoO32gdOGNbLE+BmDS0rOQsPHQlR6H5e8
Q/je75p5N4JV6ZwZGs+doSWFC9HzVcWULXzNHNqMRaRd2xaWsAq88BwzVuT6rvuP
rpGaHZMAxan5sw/Lusy0s7lidTG7m3eITw04zd4jKz4cGjU/0en6p34QKlPcRyql
q5GFGLN28nvC0Op4+CoNVcZfUi0rBl4gEDkl/QOaw0DjRB33gQgF9lb1S90+avM8
W5Y9MOPI3s6uhxpdAzuyer6OxfObYdsx96XC14FbPv3cwx1bFA6EwVGgMuDRcEsE
fDye3zThWWVW8RFzbZHUmEejRKi3hRJjoD/q1QN/E47Jyiq9Ur/LKtIlbEMhmwgL
sLZa1CNz83zZYnTUAltXkHRuC5Uvlc/haW05gQ8YwYpnu7eCI/WpBCWq745dqZL9
v5Kkhxrwp81+2K4g11YhWHZYRbUAyWUOS8kUncJUi36UDzoYoCjmRal6UvFWQIkZ
vtn2aD4+sjLhGHlVaD7cbRpKH0VCa8THsZ0qn92QbH0JNXv5j3H5bpCLhK7tXv9a
+hIOWH59UeusPAMgvf7BBZwv+oPKCB6/teJbWOXdKD1Y+a4E1jgmrpwfoV/EjWZr
wUOXOSIvlnJXJaNGNNI6wlj4ukcxlSl0rA+Tr8XraVA4sqQ0vBafK9vQAjDm00Os
kQU20E3+pfbd0LqCFNayXYWgLK+Momvd/8GHzALtO7dJHEBxl6BUX3nynXrOBgBt
FhPC428jXPruRIYN9ig4GodLAM6vdu/spHCOKzaJsdeYx24vgKSFKyBL44pvKiaY
LXG738mCk5GpsiCxbO4cfPfHCUkkVBYVfuUiWv7iHmvgbfSRfIpjh1MZxxaAmZC6
UBf8tNxSDY7GSqSsEf5NbwTdpLLZBJIPbpUHLFBy1daJfYJLjUPNlCS7tdIWzEHt
9RCYeTRCGkVRNd0qD63HBme013kb2znCOvFOvzQXfQ5ezFMZCrdIQvugES4g7AEp
Uc5aSaqkHQsQwHHQDXKKD8t6yILlezbfDSgxXYmPa4YqK6p4BcrB4bJS4ci2TNRw
FAVRN0XBde8jNhyaL9KEexkz6Jw4uRO4O4lHmU+mgXsaVYPAKWYEnvr1yCtYv/Sz
RnJFFQ+xVERO1nuSeg3Lam/7qUN9QYuzlJ32atiBYYa/tUZ3FCYLydBjr/Bfe1Oy
tn8C7QeKsv2l1iNSv80rCqXCVNuHC4NHSaBpinW7WuQXnRVQyUX5/F77O7RVKSYI
zDl6RsMLGgklr2Kfu60Ik3iJS6f92RJw6NAAKK7Vn8HI+EnBI0RmJKglEYRCbJls
Y2ov0QbotIAqHfElgFmwR3tFzdQEdRe52S09tvWqaeJ7NIGuP46Dg88u055aGiZi
QpMm08rNkvrDRTmy6xpkidEdkP4fSeo/Kl74oz0EvBKQ7XCP44tRuuoL2QDdSlQD
Y+uqK5QRSiBvhdBUuz9YxvaPOse+trh8BhLSq/z736mfQBouwKE5OdpjWZ5bRu4g
OrlxUL2Hf/uPvScsGZYT0gPq+CEYT/dx/KE4Y96KtY99T6cai7oABa16sAIYlF2v
j8HRRjeR09V3glymnIYb6xlENBt3AgPuK9MKWSfc22Dr1f+8Wg72ZXjc3RugPLVp
l6Xz6rTY77Asf6BkRQC6HURSLmSkhYAUKfJpWokpzDgEFPA4lYb1Xfs1Qm92bJw1
yHeYeR6x+723PVlePwpvT+k4f59ef7Ai8zTdy2jyjjp54LZn3jdTx8nbC+hcS20S
oVEJAvwNRZsIfeRfeaHRygJxN687tj0lmUyPLAvolKq8E9Uic7wuL48xODBREBlB
/yKr/Fv9fOQ3Ts4Jhl84t2NKoRg2pc7h2LjD7lvMA+xw9I8mYSf8/CzS5nuZVA0d
OgbCVJpBMPxBNsUIgqNkVK/e+I1HGdAA3/TTwmSCwykq2n1HFtDRJOu+KugHhweD
w0JPKs3yMRzYUQ7CYfJ47xYMr3XJ77b9xBbydVHID0WNIuo0Rsso2327jR8rJPcv
/z3eKDCr/XyS5Sekv06skw4+FySdAmK2yNEQbPCTrEPDTajHlicXdQUAf2RTSnO3
haNbVGE61Qa0tkE+ccypKffWOYK9PQ+OeoaxwO2ne2XFQx5iG8WazwCnSV4SVpyT
sf5GA8FBz8BsBOuL0UpFn+3bgxm0xm1JgApfQG9y7a53FOpGGfUKpwS1HPnc89at
xWk4VPlxQ0XWv4d+P95ZGoKKmJQgsBpkNs436wuVqckRz2CRjk3y/cUsNTEgmC0X
jLsfgZOfyJJvPCwmL9x0ZtdBKAr3MxgcUuWTicQ4mM4QTUaurUJRM3c9y9M9Hagy
9gJYaO4ymmi52DJovX/vj4J6/2PwqqKuRA2I6Fo9aoP11lvcNeLJjoyNMPTbjcw5
vt2PRIbtCHEELHT0KefphQNSy0MOJcJw3n+Q8t6sZ26q9KCcQSZtcqeOEX+huw7x
NupzC3kdEN0mvY9hNF57ilB4ltzurQxm0q9Za0gM9JZ0XaaDTf027FlLnZ56ROzR
P3B49PYqckHIZ+nCg3dz67KFvZoFqE1m/wGbsk71By3L0Zq3GRzpL5PvEUB5kfwk
kWYl3jqZ+3mO0YB7H4iawjaXjFGlrDSEx/leUWy32ykGguBAaLZN44GFcGWA0Xjo
hj2GGOq1NvLQP/vR/GTiKlZxO4NFL910y/PmqAB63/f1EUkLoCn2J5JbwPKWaU8O
m9hzONM4EBk/nE+rf16PqgHL7UxIdzzqk/V3pKJgYXPp6zzzRAxg8MQ59ZQyit3r
eEY6es/15+P+e9JndTjoJaDl9O6nqCoFiCVkFo5rRfHdeHx6qp6oEgFPws+gQ4/b
MN7hMbLB79pR7XZmnnACjGFrlJWX5q+q6mbUfEtZLVXoH0aWpme14praELy3EEqJ
rJQmizgZWT/rqGgDnrbZRT7laB0dqZKRJd1c7ZkH5qNsTRKAnuthoQBA17mjBBVF
oEVIOM2KAN0xrn581trA2YRNhKOwVFq3v+jkJqo2tM6dmUBCDBszkooID8HbKOLk
nVzs+EB6kPC/jzVSBiavXfSdzACTc7PT8gxYJ0AyV8Xi24vCsrSnVlAhXkuXqNAp
fpN7M9iwRkL3UgtaUdBqbY7gYN8X9Yapd0p/5iO5reLI/RYRzohdD+X1y2tMmtsc
dZ3O1ncKAJH/+aGoqwMSl/gn9cpYwuw/6n22wNnsQfgOxOt7aHocbLvIKIu/qIex
UTSaQ3DY3iPJcVjoiX7JWjOoNpIDjBEFoktqVEOXAqPvaXXN6d3HnfcXuuoqc3B4
W4lHZgRiB/avl7sAldkhrVusn4GRQhnNTmzIgNu1zuCytFF8U3qmSoy+kG11oIi5
WlwSMfECxC+zz79ADfInN0XmIzG+Lc4fnZWuWnSErAF05Qb6YkSnelvN4gq0+W2y
yamw2DQD1ud2DOWiTpoifZQc9PM1/C1zHh3pWWgegcq5sg9be4hmmNx1S6z17arU
WmgRmoqatBVpTb2lb15Y3WLKQ4KIQM0wwxyvTkxp/oBpxTlOI7zV+QqRONhVJBZv
KDWMMMnXWVibUZNsCyVFfS8H5+KsEkwnaeX/oFx3Bf/u1B0xBmPkwV0t94cnQfTx
3f6meFkopOTNJXXErvyOslvRuGEWsdtulZ+OydIJ/NOLz1A7w32kvgK6qUEnUiSQ
MWa7k281a0ftHTxUp9ne4pyQFX0mf5Qo57kVBvThZd7nm2wGLYyEhnZ2TypC+RgI
Egm2w+cL1QciY/AUaKW6Fbhw0QX2ThpBmOk9Gda6AC6Z5kwjLenpbBw1YEMLGU1Z
sIHIwVeRv+V6vmloe+SeSU0jsC6a1SfGUAzoJPAubRExDWc/ny5Gr64yFdo6NU4z
F4eAWt9lUtPnnQZA9r9aT5kj7mbUEHRIC27Vt6sHKMD70g85O/8/jdiVQ9T3hsLg
46UtVB6HOLuBAIZz4x9Iodm4SYB5kdAQWAS5ixGCsveow2UlpR9qb34NPRdRMDyg
qj9qcv55C1u6Rx3n1N8Hur5rPkcXEnivPmKpGefVt9AJ9KlFsEsMjCRK+kpWW0rp
Eq/g7DNM2DWXp8Ceo7Ftg5o23y5XYCExybheQWch7h+AiU1xPmatNJS5enMJz/UK
llPGjP/Dl1kaNKE4EjbUY5dMHAbmfSpWnN8lxQj17d9QwR4nIkhYyF0nWyGETwE+
h7r/vV1HElX1boCCueU1cz65FOx1uqarm1yhnB6c7Hd33gysNTeYC6L3a2LDn3W3
hRWO3oK37qAh7//viR7TmStlQQ65j4rfUDKvHaFdmqDVP6rXSCuZCFCD+C7AGcdd
ewid0mZeQ2QBZWQFCfle8ZpcqLsP+zFq8K+lcqWy6RHBGFCyBUtx7PRt65FBRbEG
wIdHgT2Iuz76Ba1y5wt5NB77dSGV3wmRgWeIRYdzgayeke8QZ06O8uZKFzgI4AuS
2TNOXeEoLtM4TkLm+IPzHEZyLUWXqYCb7qathKQgB+03GuztrBlqGBRIICYhbn7G
3Ha5SRePClyX6C9s5hZo1GlUMgy7O9wvZnlBIU8GhYfU5dUS1LgRN9Iq2PvOI0+2
3SSeTXjQHYDuyKCMOdQoIB4K71l/8WDzyFl9kjL7Km2KIbIKO5OicCpAkX65Uz5g
OnKqbFSj1wvha+prfS8/hh90jQLu2TEsAmvE2VVmfxMltcOhw1dS7MrpygonmB1G
33jZtieGSwJguHlRqQQanA0G3AUNv7RUwXdraAX2Rpw/ak7X0xdPgRUGn2O5fBXB
1dWM3um7zQRg+lBv/ea4ZWxo2uTnOr/1HU1pe1sOI6LyiUD8wLdJmi06mN/PDbso
O9bfQplPGn05sfct1rkLCRJdKbAUCry4lbLCZLJVYFJ0StUMXhO1CNKIF7Yqzst7
E7p7YrZeCKu7v3p2+PoEtCtcJzaRwmi3Q5dOBVZ2GPO3p7mgDFGpb/2SBiwQR1nG
PMxI/Lvh8cPQNLu5boL81NvEbnbKbv4zdpWPjEvyjOdAgt4J6Xu7qdK7yD2rTtQv
Fvm6L2MFTIPeOXd6pHgBM6Bm3ayo90YmNF17Bc7HbABiFh3MQVAULn2oIi/tFNLG
IOHVY3Mo9wWsLxYstIyduZp9EaQMnokpM4cpy7sSTIPCo+00ssPRtAJuDbCLotbY
TSHvWTD/mtcE96coFldgcmBoY/oVn22+zewUAeWKS+gjosGl+fUkb9WN2qiyHSdV
MVyMlbmoJ3t2IEpsmla2h9DMXIwTY+2RVJw9k+08zPQA7kvFv1i36Rogaxu5VF8l
V/HOe+5E/8JtfzlSquhKLmF0r232xkSR6bZnL+vxwiaembStb2pRLE1UVOf5bW8Y
iehv6B/bTi7fC98uGJ+XY1NSuttHeAoNUkrxvUOuWymHnbAoTnWSaxytqFN5seet
CtBh+97aKo0H88Z6b905V3K7nAcrALf55vtTjfqLS2ynrTmCSzS21Abm/NK1vbBw
eNluxFKAYjHh/+6t+aXZXwlI67q36fNe2FSdyODTuQMsUd9HqGmhegIdO9U0RHww
UXYlZaaQqEXdU+qop2jYyDpD9jBVEkGmMq6BrGVBBQ02NkLGZvWpP/ReLpDiHuMq
setIrblqWv5GXcPE9Pf+e47bMBoZgx8MsC6dKsa4AUMawuHvgW8+8Zq5XxfC1jRa
DEn2UM7N8ETAjcn1ypvMw2onvqzSom4XEf/XbnVL/k8agkotXRSReG1NlSfKgBd/
eLT43iuZdybPyEPKciBwFUTcAVmzAZ12wP1rzicLcJ1gsEeftAktV5I8zd44fdaW
zi783KjARQYARDM606H9knKclh6ftHAcDb9PVLJIqPCNUrzaX2vnexAHMK0cRWMS
fLU4BUGzpJUU9Zxd0uAJn+fjY2HLtP+itBXHqpYlYo7KDfxkqi7Q+oM74vf/wkzy
tODIS8tmOfG0CoemMHwT9ptSv5EFFJGkEJw3Ioqd1oo1NZFvRMlp5OynS9A9Dy0Y
fq7fxYhwL6Jz8WiRyCl6NkOv5ydKknhzhp8zzLF0uKIu+p3hWiyvjTai9od0Bkck
TymaBzqk8xH+927/M7C2SB+Ra8AufyC89R9kLKRVJplu+4QwGQaR+wVM/JBjrHt8
x+eL0bwFa41G4LnVfEUnFOXg4N3e3rvekGHwuPZ6pPLyANy3+glNufoW7we74qBm
r3Fns0Y6Q8uxBgqIlyQ5TahEc0z1cTkOP2DeHjhVRHVKamnnWHMhweUHOBUTf333
wnYudaqLMaVBKNjIZREn8qehcEJJzZ/mRPnM8FIMKyF8kRDS1Bl5PDWGEclrPa/5
Or1hGnZcIuf0+DcbcdmUDtznES+uhUXqBtakRyF8pYrgaglm7OpHskXzvxpxWyct
Uisq8bW7hE6cTjFwyxZZNMRwHKTc+jyCKlYqmm/G0M19rJqYJvaVi9jH212vD/o7
+UR9csKZGp5FJFPV0x/Ey6HEV79zSYFOS3hQhvMh10aPOHeJCJEYtxfkXUt7eWsD
SNi5yhvVZH9AMt3jU0xT+Xn89cMJfM89hV4uNaIP2fKsu69aCzcsUiVcVT477q5P
yPiKcyQLgzUKtsfRbXk2vjD0Qi0y88ITW4VUgfuM73C1BJ2qqD8pR96WazsgCdWE
hllga1G579TvIW71FmFpGK5sO5Ux8qyNCAqZ2qGcrNoeX+TzzUkyWhtIkkNi6wos
P2m+qY6NQE/kmVpai0lGZrom4aB34mMNGOMNgADRsZU3kFDiTq4IC9/5p3jZpwMO
Kp+slF+doi1SWROHKAXPRlkJfb33+U1II86aMpVLl9HDhp+5gzdrMwDuBv8NF9wC
oaJ9jBD5P8NtljgxN7hoTeFWe5+/PmMTWW3eIxC9hbde+TOquKcYTzShaLqKB3/l
M9TpMo225dTiAXc4LFNqOui7a6zFdrRpKsYX711pVZEhdhjUmBGdqDWaZo+OiOhb
WkE9xWJaxptcm0p4rAkgtriuHIbTifWax8bjZx6+58r4wQtNO7cCz4B/3i/KsdKU
yziu3WpvZPSO9pa9FnhQKJQzCsuXOPrGV9XFBM0wvXK1SGiuD62itwDeXby/DaX5
r2ke3neTE1ejHJhzBcQ7jcEEq1T5ybczb/vuzc4kfUwj1E/vYhnxsU/g5ZFb4qo2
FwF6TJhoAijJTlmWKbOh01ImOgrc1wHrTQ1/U04EXBJnIWRv8OX6QFzX855fIroR
HfqDgq2Ww+oIVZ4tWH3a2JGzI9Igrby+kGkvxJNRYcgFbzKuR+AA+M2+Ma3iPNpe
2NZ05XR8zFKupPrcFw3F0FLVOHUPaeivpa2WDl6wEJq+9SjA6yvecAK+rK3lFn+H
83iv4W6+msS8UpvnMevhXSW2jpcObcja2R1zJxFB4+9zF2hbdyzZKpdkA08g/x08
H+blVkTv2ayRyJsXCUpbIK3+d8VgJlIVA9b2WXdCVVdLDWOmrM5ctfef0a56hwrC
c1kbVrFss1M4g2wGL+LZWt1Ww14BLmpjoMpXbi8M8crJ4xlTVORNmZcFbftpSlHR
nsPjtp6s39NOp12zrI7eQzshAUDrkgWkjBXlGAKDykinociOP1aCGTDGtJfSvDEC
E5+SZ7OsnDAgy6sqXi21dFCwSDS8W2sRVj6Sfs36Ix8Zpo2nEYA728g0hltxDhR7
4mKmrGCWsfqIGI3344StUvYQCo729+iEQUfN4H60sVktHXwuF5Yulyv7wdtYSEdu
cgkm+lh7Q+a1x3aOP7WibpYZj/imXAWKjNMb+14Ca+YVP9ZSxtc9QJVofxiF7CaB
HcGHi93nXSgfuagbNhc+2hQFxzLMJXcMC4ADTlCy+wi1XK/t/FaJhuoybCHZwNuK
l18hGHAp7dYocgV3Bgie7sUYm+heOa37ldRwESsX8mCoVQJfq4UdaDtM54j/+wjH
HsOJxPHfjj5vaRQk/ynkRw4NjULL+b9w0wgJ2NRHlFZVQlide/y7ZT1JkkAxSf8r
h1xDnWThtxZl8t0agKONqr+2i+4a9a8oBHH4mqCPTQ1Nu04xSc6RybLqpj3vZDWW
zMgnaIKS7QsPO8vuY+3THQcnUmEu/ghHZioTbuOYEHu9on8cg9ZZOE4BMM0X6B+i
D+ou8hB2cLNoaFIQrF1X8jSaQFHmQi7TbUToAxD6TPJEQ9bLU/i5iXQGpg7/Stm9
oXp4wzABIeqeSwfEb2AMitch8nTl0BhfdsHPPmx/8a0LhqYYPAtzOZcmxodfn0UG
oBYk/6CHShK7EzxXrVHxsK+8FoOxHTHJYPOYzxhYagKkbT+2By275emJ02ji3/tu
xA63C+0pzRq80bmm9uJh+fCQzrOtHyGVUbNImFKDqahFJsk3JPUd44kg+u3wYlKW
P3Fe3lY8hcSDiq3TGCIwPKUm/Wl8laBF10rSiyVjWb7ZQaHb+TDBNENawAx9kheq
658oUXZcgZvzsDBYc497rxQVaDU1JeWtlC0fRaGpgajG6fW+8pR2k3togur/d44/
n+qtDThDhHjrWrDYag9ePZ1W9Zr4uvr9lKbYdTdU9d2gQJBt97VTYH8NwVRiLiov
uiN2MphWcLU5uH6dXAtu+M3XqXSgAQ3fGkArJ+ub1wHiV06GHhXuzpkTMF+YgIgr
FBXXb5RdaKibnYf4yYMNCPQry/o+IKdbjcAefFW9MjVOrUsQ9MQQY21iDKiDxTcK
ln2fAxTtX2lIyr3Yvnfr/Cla1UvP9YSZvqN9TrNzKi9dwwlSBOJINDBzq4l1S/Tv
stHV2vA4Euf1K+rirBHHliQAGbytPSlQ44vQ40sZ2aAmqTYYyzMPrgD9uO3f6bCL
yLVizEe13U2GdncAFzWSgrwa1pWPcaC6rp25I5DjWGOrGO15eDONAjtImOXSk/mR
jkgD0y0Zm2Bo08mtOY0KU3c+iOvo6QbKANSacp5r4xCj6BfZOxBzej2e4o8v4v/y
swzPxmiZSx8ILmY+ep+6ZuSLo5PaCIw9+ErvLavqCljVy3aHXY4DzZf3E5PXAtgO
emDJ7XM0ddVluTf1EkTyilxPRGnXwbl2dHTmvZJnIoVGjYxJ0J4qvBeJ5IwmPpgY
6fFztY3weIToYcUFtvJINKowSmUIMr6nbi08kqWzisyOFngV7LvQzKlkVhpOeQMJ
fNP2eM7QsdB8AnS29Oazt7x6aR0TmoMCBnekLYkKVXfmOoTSRqPxH/gAE1jbSoEL
T3TuUkkScWtFXRvLt1R1eEc1BNLiKAVL/2Vq8I0TiShZDaEFcGb887HHRmJMLoMx
2gAvTZo5i4E2Rc0Ols1llE5u5piuYU5R9NDYinmg4cIkghBD1ezPZp6r4TUiMXCG
b6ocRQXXJ41E/Skh3XOH1nXDnxzaTG0feZz3qqm723tKt3ZQDJMOCw3tB+UBgCCd
xBLB5q/vsVP5dYCCNtXzS0rGyROPa8VE0JIP/Vkq+3M/1kJm+30XLa1GTv24TYeI
re+3E7ZUIvmG3x4tEj5RAV/gdnUqpgKHdqB/LT+4tOVeoNN+nGJyA2rFeiwXZYNN
eVGkzEwGgc3C6Ha3ZDACzt1gCx7/I7GZYa2H/7t50lrOwiKF+CD+4NrdN2PMum9P
f45JAcBUoDaPVG/pzXEaX3nr4qQkQ9VKczo+7odS8j0UUjU6nPKbIIufumwboE2S
xD0VGqCQYtoOaRrsqzDjfILw9ZCNo1u+WiY9XeYA/yarARF6tG2plSWvE1lMnjiL
B9NYJHEFiLVCCvSQkc8biUQE5gHgfYRD9Yf7eEMs9xI20uSE0i4hNDGYoQ6c1Ihs
BeSBsyRh0WfNmM+10PmUV6Ld0k3cuGnASd+S8VXi+CkqIUxQeJcNx2LcZ+d/t5GF
Y6nirrRC81Mk13loYLt8aIuxZNnk6RwSthhU4Vsc0SDuNPePKCDQu+nn8Fh9BijX
HPH5O8GZHPXk7FzuImZFp+8WLS6xpn8Ipxd5aK11WvexwOvDtsr/sntGViGTCzoA
yKiUsFmGbKnY8AaEMZFB8ztfwD/xBW6NqHbx/ros6/7MEMnZLePK6zJCWBal/vfw
Xxc+YmCWCcpxttIjPI2tff7rHMa0TbQktZKmiLxAiz5s82L/+oPqMaoYut7tL/Kt
Y8rv5hOj0q5+nlralRhkRqAUnPQQCI1yYZureJYRzl+xSeYVJApOTPiZ7AnwCuJt
//X+gJv4wh0BGVnfRmwg+LElI0Nb/BDjO/q/UBY0wF3eZGTljUzz0jIUtM4A8DV5
iDl/JW+ZQz+qOlaFDVArzMwaoQ/LZJfcmhi0gyZ6aaOdjYgRUZVS7EPIsjyTITPT
/JnYHQanHYlRvT8sXa+JSxGCiqaGtUhADQ2ZqCqwZyktn5+SmiwRFKPLy0k03nlk
EJo3R3ZGBvWO131OAmgTvaWojGRHwSuULocsZLude0wGTmxpEFdpTjWTqNKnD5cN
ZXOvowma1jPvNa6qCib6yulDfB+SzYzDGQOv7aszV2zeoUqTJLlJErHYrbil6RVn
asYmj05kpPwXAuyTm7sWyoxP3jbne6AJhd6ji38MkUs+CniUetoknTzelz42iOAX
M+LfzpWDNvOVNWGHqDQqRyBL0qYNcYDB62L3Qt/LO0V1CE6YWUU4MmYhtBWcizAB
RI+EU7snGUFCAdyPkbwjuR7ENFYbaE8aHZcL1gOSw3pTv1niPrxxkDe5Mp/lGTQG
XxwCAsZuLPvy23+eNAVBF+4T9ia0UvNG2Tj2tPrOXa9ylbYi7xxbymv9WOqtyiea
Yp2Ab/seu5Px+tzPsrZHITdVhQbUhwZU3pSjGilcmA+Ji+a74FlT6hUc2Jb1v+Ir
1+qeKeYkVb2YSr+ac26DfF7UU2qdbyaNmgBgdb6JO6XEIgiQmA8HJhB3xGpac7rv
zknI55I7FUW9Aidv0YuoJpGjbvpaHWURzZrno/osTkJsFVyd4Sb93fLBT7lCWPsE
LP1uTCOaQK9GO0wawDpNU8id71JRc1yDPlVRh4o3MgHFU4ye+IVHoBI/GT0CFh+j
VWyuYEeMfgLYMSmGExwTvQjlUe8O/+JuubQyeBlp/a2QQ+4A31Scqh18WD/HL+t8
9jHNsv44DG3v73iQPJdZyyEABB/kEQms2Xr5ts1ExDMYMQZ1OIKedU6qhDVP3EqK
jzqgjsCEkLC2tCvFqnSoexuaAz+lTg6maCiX4ue/D75TJTnjD07D+V7GdNE1/B5a
Wpno/kH+kZaC0hhl+hdTadc6NHvn+JQEcd/qC+Ox0fb3A+NTJ5QPxfc2I5iD7Fy5
mQMSeLUxSsj7Lw+nDhOhofiTajOgUrPvBYbIUW7glNlIUQllPhH/70AIOZYcw4jL
M6RwX+OAFj+hECMHcaKTJ/Eb4GjPsNfPV3Lsj7mqJmoDDOOsa98qCT8CQ+6YQB98
42iDWjUhFU05ZGdjqatOP9SpBsoDuSWa8f65GjDA5YJLlWHhQlO39g5VXd05A5zC
/WJggdmGSJpFxT73VuWhY6XbB81vaOrUTXp844zEPaJTrQFAk31Dijo7KnO0O7zf
AoTBbsizQ5BT60hb+47YCwC9C2/U0PnlmpqOj/MnrC32AipS6EK5aeePI3iWycLd
GjJ1c/bLnOaAf4ZLHOwASoBBd7k6gSpTENsLRB0qvlR3hnXa2yTAEzDHuHbfvPM4
eIqforoT2QTKb1VXsSxCo6kMEOHFeWg/pHvVc6GRtUshVGAGNWtarpHp/gqn2uWI
bvj47WV8l9M03thiSrtwvm8IB3wlZLYTLGrxf+PxSgo4nh/jkOb1+yYfyxxLxd5N
HM4Lh34cf60exX469c/MOmYm1RmYrN91jozQFJR44W8nXukWBwoXXMdTiPXjAadu
z4+dEKr6rLz5osfZHygpEPGHfsiJv3FfeH7n2lLfmTeTBIUAXgrsOa5IqULm8JKy
TfYBOoaLoFkrrxDp5fwf3x+LWsm8wT6yDd2bOOGBuGjkX/HTwcRC6YD1YkzoMGxi
TZqDMAfw12vRHGe/54FNHdJPADKG4vJsR5MbYxzIFuB51UmolT3cqtqTpfU0Ldqf
SlT5bbvSVXGUsZyG0bmuSzJo8Vy8V/PBuT9O/YGWIn2DafNeAhKrN0q0KlVTwgVy
Qzgd9Muozc3w49MorJFE9C0hVz1tExLN5stlsViDO4EpR1+yb8fSQSBm9xvnPMK1
CJOleeF3CaGs+U066mDIul/TdiYXrEZqtu0GrqNCRH4dZ8sHLvqeHiUVD1LZx7wE
JQPO5AX+Pd/7ReL/XqfkjNYypoAlFFtNDPRCw6IKeBlM427XRFweY4Cv8aEcbFhJ
d8UJLu+do7mfClYMpdFtsZ24BoHWe97xBkjo81cnt4LA+H2uUILERVZ17u3QSMrq
aDtQ+yPi0qEr1G2BI0ShuW2ZCxYiLMA5CRYHxm1nIaCAvsuJzT6QgjSkqgqJ0JD6
00oB22nBh46EiYDG8IPRSlhlY+u5OvUEr4Te9XrSKAP+7BBxTxc/tM4DWOIQZzOR
Qaitk9deWTTVhctcInnPp9H4VKL4LLbiw+ddXahFwvGP6a5UraeS0C78AEGcVzTF
Ymh/u6EC8n+RsOr3iDhiUcdYfAehBy3DmzLIF87apUg2/n9IzGgRfbFIsbVjPvSW
oTIFUwCEz9j172qi1WAcNkHifgV9k/T1OM1UhPvxnDItjRMZDnqAoTO4g5K6ZXMG
Cmy67dQN8ahA62AcigFqJ6yhfDyglkYBcsSdSBHev9SMkZSURuzyPrnzvC8RdixX
hbJWja5825yw/RPQt1PaPmmrHHT0VDFbECUXF+HGXTqgFwwxoaXUqqbx9IwPzAou
LEpZKLQlZ5gCIznSFb5zYI8ae2RbpGFVmdHdTsHQD8UFRHuay8NDbzLouBDBlKky
XTQRz94ttj0eyRi+xVTR74GhwzHLhcLOsfhXXnlZYXWQvLNOyNVf7RQy547PDPhj
2JPCGjDamBBbo8i8LXmIK7uHb8CeobGr8sEG611FRA7Egw4QkrMXo7KL/WudHcs2
3KjzlchFbnPVtTrvOu1az/2b4xSox4BEKGncJyT3hiP8isqm2gZ4SYQ1HjegoiAG
YWrFdbkCLbmVIMUSFSwwEqa5PUZnQ/kNy5zB/OJWU65YR2x2/eQbAb4OtuUHOfSG
V+khrhRauQ4b5E78v3y8OT1BfQ1LU1QkMR8ZGwVf8tLV6LT6CDriocpqotmafu7J
c8c4YeVJZQ6akHOMt9RbanmOJeC5LL6uup0CK0bIvNQPTZyIdq/Jwk+ncXA8Tm9o
SsOtzxMOjouM81nG+m92SNRMsVT98EMmifbslhC/cvuJn2OfyaqhOFUH007pPPaL
z3c8UUWEtAGvr3Cla02hb2VsPCSXW0HyYYoYa0UAzdTUOMKMAFXbfHwonEkcIDts
zlGGSP6g4jlO9fbZpVLJDJjABBE/RHjIJ73WjroDlaiRYoXqBG0w1TNOcal0G3cf
ucKp7wmgzy2i6eYhHy+jPgoy7UJjeRaTCk7ARq7baAQ7OlrCumzP8b4OQlmRxqID
wLPlftlMNmaAEYuktYjyYMH8Gl+52uHq9PHiXwhHcKCRuI8NfeMDCg2V2jk5LpMp
Y9+R3cngtoMVtaG7JtEMnjdKxkup7bKVm9BSvcKCD6DTp4HIa3iPlWWiZUuq7hoD
nsmVROHU8cPwdlx4ZR3B5tL1XUufjU4X6zEA6FOhOyVoTQAISFMTRRDIlCFZShuj
MixW3U5em6AkedLGzWZrYGTYculavvCUZ4yTS2cAsKzUI9i1z7gTfnjpWmUXoxb2
I2pZTMp68qN5Dst5+Xr6xF0ie9I6N1L47V8ee3XgrNsYLRC50sOBMd/fH7mX+y64
R1FCgTqKPdMIBE8v1qyORioiEpbQj7OIZDTM//dbwcvxAWjG3ZMPhj4YIson8Bng
7KlRek1ME+M0s6QuCD3bjYOe2/0s88o2Nd6s2E9ShsDH2+fanUews42Q4zYTjpN3
MyBECrIXrwSHUZVmUsszsaLbTBrkq83xxP+b2hFHUF+xBMsXFejWDaQw9HKjQb6E
gbH6SFFFrhe8sF9x2yn7nPYp8LztPty4QJIc1jMskSGsPwQFvCUoknRk/jFTbxSU
+Qd3LawhnjDZwRAdziPDuDxZUXNgcmFnOneXEno0ovpV3D8wSDmT8ect2qLr4mFV
1bWoip/X/2fvIBoBGZJ0hvMmToIZMDf5n+fWuTBtQin1ighmPnNeP+BTf/p+ImN/
goF02z3gDtJyM2TuSa5L9yebzljX7wFPeg1kNguYLoti5pOptmJHvJIvJCu0sJAJ
Y9+GkqOWC9zOYRR+RBibx8XyOZPql8xAAbd9NYSVzxieJuHv97QK7H536TFYIBMe
Ox/vDl23o/KCnseeqdsGtl5BQbLprlE54TalL+qsw+Mp7t5uitwDjjDM7JRswjPs
m1me2Tmc1wwf5WhJ4/iX0GPhjyogigXumktqMM4kpgi7whrpuj08cZrHq1SKzhbz
FailRzsgkifSSokB+JjGRoNuwIEZrJOnLaD3uP6/WMNZc7Mv5UjjMvVBldaMUbvZ
r3RrcezpdcD+OuGjTUudp6qUiL1qnkSWnp8FpI1QMKNX5ZtypAjIRmvV/Av2SiVd
OOwloUF7hwUkeY/ZvKH5Rq+w1wg0tDVS/+LGIwCwk/zbAgkpuII0qZE9x9QDThTi
ltTNlVHKD3klB1y/1x73+66NB289H5Ho4fbNbUytu27NT1WnoYWHjpEGrozjrlp9
/O/HWx0/R84SjztowpHANhbEc2dj2IxDre30kTChrGiWXHPBGnnn24ZaPihLn2jO
HCl28TvcHqQ45aiaEcBSabgbfxZDBNX0bP/3Zwu/V2FzFKgkCcxUzTn+RgdrWXDW
THk5i5mnIYverLGSvZmzwJdRw4fOLK5qyU5f9fnhUr+YnsQcDbi974LxlXVEkw0H
NsmfGkYs76JdxdhkgXBHI/t69JaOt1EdXXaz7z1xdWTnG4MGb3aiosijwlTQ220X
+k6tjmU3KoZTceQeyT99CikaRgsivzX684BP+C4yHT2lwfH3UxU2uht4B/iXlqXa
c+ZvwORIaHyl3xKr5H6u5pplCEThSVVOTCPdOiQgcWAapFgHnnGeX35Ad0wj2xgK
mka/HAoq3aaRXlVvlP9q49tHCzGaM2ki30elrR7E4+GZXiVEkNnZDQnyPLBabL3m
0Ciphdxp6z/YEE6gkmY4XQl8yzoCdFfFcchhQKhC8IZqg3N7jtMob9Mt2S5uq0R7
PbKBgpnIPvL38SPHBhoMMymc/e08//IBewB2C54N6zz99Id9qzeDTACB4SasMRf8
zkRLIpUHXJml5tqqrugfb2vhTbJCDvrfhXMz49rSz+YVM9Sxs7Vj2vzwXIEe2RWi
WuWPV3nmULknVqEOd66uLIPd7fdJ46UH99ixjmoU2mqTpCEe5ZeMcH65aHOo270J
C9JToRzkUYFVjGyYLpAAo8r1E5PbAK4VVUFSuVL5I48Zco5XT3zS9m0KSXQHPM0S
DjtEsL2HKvbZZPcJBYbt5JnrBZJA5na+/MpBHcd832WfqdpAaNMSN9J6Gv0Pl4DF
7XdPnfpwUClDs1PcnHHh47OJI4ddm4vyR8BFApkadEXvU0edlb2+e/QZ/LwqKsGV
mp06+D2t1W5oyR8xEfAc7Iax6JSJodj6EUeAm/TOM7tqLEvHFDLq9r+Xshz3Mo27
9WuOICTuGd6wD/mNg+JUxU0gEaceXACPWLqdVlblqn/D4iYNS7aXve333I0uzYW4
aV8wms+y5XwIfeppETUX54umNZNc+wevZXrb3n5b52UOOJlp8wJaAzq+E0+IWwP/
wxUnXO+DiANRyAI39le5GwkZv7Kw1WHZrypd8fVI53Y/7f0lgeu/Z3NnG6jgRKxp
dS0qPMm/5EuRObPUOaseZfnu2gQJ2FhdG8+FlI6kkIUbfYxBiGk5zIyyhjYDBBmP
0iOSxoswfXqaWEi61Y2ylU6EGgUzNuJpt6EwLGl4VrYuwY/KD8ZYIlldXCnRLXJY
9PhUCx3xJtMSwkROYbOOS/Sg7mBjyzZOGYL5D+AiWm+5f9W+MHFyalbvwVhbDloz
uAGvQKwQ5NvT+ivZMMT0Baua3ikyn0YZYMJz5QU3njqN1gCN+CrQsYF9ZeUp5Boe
kk2aknF6ocW0DP/Muc5vVkCAwgeYEu1ksNKAF6565nZXq/PF4PkWM/TtMULKehqR
EZOYW8WvjVoWmhF5L0APj7ssP49b3B5rF6xoSPL0RQJBtM6VAaDKzBUPP/uhgCQ1
XYOWnirJSSNag4xAaZ58exwQMv0PPv5/D+sPcDWK40wvw/+aNbFm8Q4YkJfdkukR
RZTX52F/9b0smdMtiQXaI6fARUb82gCqdIFx3FmbbaHWX8EqhUHO+CurYWdR9fFa
Ax/QjtAaUO+lWjvSt2V8z+BmupQyo5D3Wu1ZADXnzvo8Vs2DXXTF7y2wsiwT2C8q
n2wHgGHOYenL8uQaqBbJDZxoSCsZpv9+bJ4a1PrNSD3pKt3ofvhTH5k+sKsqWgPE
ki/dB+C1ucN4eq/ECGpwUNnbTeeVBZ5sNpBJ3uiBirAZDolQSPyl01O88jfC4G9t
Me32DWi5pkEgj0VMmnTJl/+CVFEskLjg5vCUt5DpyHDm+ZZuE4Iho/1A98UIfz+E
/wpCSEeREU4+gZjEWxfhjVvqOT5vcwEc2hzPpbttYXvGdD1JdLo+6Vsg5vcIsJf4
QzU67MxUoIoHSHZrwLgBVbtNJ8jHl7Zj71hLNBQ+y1PIFlcd6echx5rdcZkv70GP
R5iNic3q/u/8iQSjusAmLSuFMN+uZ37ScntRb+3i41QAvkOqbslD7+R2nfcyWVXb
/hGZPr5FnYQeE40hFBUA/V1Ndh6ssUBgBw16cCT00IN/a12RtBhVxWvA9nwpYUvo
FAOZgdI57Qbkmv2yKOX3hxO+pswaLM5QaQZJo/MfNcGCEvQSGt4ohp/Vy2ukOrFK
kXkhtWg/ItP+agjGWq+98jcJUXSXG37sqjFTU7rerRno82uGw+/dv0P6Uqi9yyen
K0CjS8MR9j1OGaYQGDXhklCEBRF8Ll4arCptbZ7mG73clJOR/sohpyBPmKqOTmV1
GzoE3+O04SSwcKZmvDTmepKqwk8xJxBBKEVMWWhtccHVP3UVSvNSq5O1lP5FF90X
SEw+Qq6AVols/3lIzp0llP67ahGhUh6gpOXLEJZxZ6HbTnJQs/DnGs5Dueo1V5dM
OaRYfsMlwtnNq7hHkczCy8QqrpK3h2UyZRPJOdM6JQF6u4qclEl5V7HHmfBrXJUx
BFN42TN8daNhiIRQry4nN8EZVSn7VrUSMBDS1awbNB50Yt+n1IiPPH0BzwmH6B3Q
3X1Xyk9HcXzQ0clo+ra/s3VJiOPTBSlYH2v5Vvj5wXwG+x4SyZ9Bg9TTzZ2vglUy
+AtNJ8ZEmq1oAOtnmXkpYboDRjVMgogOtHvlVzQ/xpm05Um6HJ45tHNRZ/JYUP2w
ei+mxSd5TUhGur+VkXgFoPXER7tb+uY5RHsr60PKEgI8qpEf7m2YqKUF+bOQ61Gy
n0G2DcUcSeutBP14QiaaRmmGt1LKGQL+NlTGeHEkMP3MVN9D3KmGEJvhZX2Kt6It
+krd1TKpbP786KhdGerhOPBzABxRuhfO3M+yDKXotwah9p46qHH0CJ1ZVEbV6IJI
XjscZa4X7r44oCTvfDx3bTlsstvpfp/S3r7LtjYS4dm/7e6ohfL167QHgOs33BPK
/Z/fbMEKmLYEWXTuIgiTQQJ9mekkZSBKoYftM2WpMnZDI4y8N3CzU4eFuGa2dpKr
nfgQNLwGpzoYyb32f27a/F8vA5pCfr9O5SVQ65kzc5Y+mRuWIdTv3GplBmQWOTuB
uU/gGniMNFy2EJlvncjRjWm5E0GSwzQrFXLtmZxLjOTqfESvOFbyAZANUdfz2zjo
DioHhz+PFN4O2cJK8uq6hNniyl9Al1BmgqF+EjsWSUcxTL1tIctyo67IaIBzgWXF
A8RgasSy7Ddp7D3Df4At/n45DhGdlzoOydw5Q4nch6c4dhqZHkDZsdq6Bs/uohhu
WGlXWzSMQ5miSYyQRSxaqAlkn90vHxmhXQ2017kon2h26evrutBcNs8EPMfwUeKt
/FjMVcTy39ccGIAA8JiwG5MZs4A1PopjVi18fPvv0B32T++L0w/U8EpGu+ZG05H0
8Japt6HHEpf8qXAtna6nQwB6iVfAuGe31xL9qUbpqVLFj7lw98CqQQgi8htorT+k
wrQEkp2afL5WQd7tmvR4ZlbWGKAtAG23CEEc5zSYZfzFp9YOIVZD0kL3ohqA2myH
8abh5CFRYXsUNUwnc/QZP5FEv7dtw8MSin23F9BnlMqf0R+ZBOpFqXbGuzUcSOLA
RDre9yGZVT78cTUWCU6CuBk7+UE+akcVBn0caXhrO0BBUZk/WnGlWMLn+SYcEoiP
JDTVqMKFtjxfdF/itklYVTvD677dQDs+C3JWI/ELllemv6wlUtbQI98k4n/mWCUP
NWc5BKP9DRNV9RpHncjpbCaHR1ldoCwNzMknRr6MAT/lfiqTPqZrLkLUXTLMtNTK
/0HC3SESKdAn6J+Tbp0ZsT3wTyjKYrx3J2v2T0T5Z9mjGepg+2ZYteVoGIf7+6xY
L8LTTdaK1KiRC0t81Xc5Llcf9qJY7bVHTm74MAG56XeRoBTboPYm1jxX8pwIrYtf
qrfLnEb99+ezRwlTWelnBBAQTiuuOnTlyOtWP/GyuCWWgQ8mYSLMl04CyfxRg3Tg
M1sivEs6Zmt7WeLczrfSHFfj1xHywtQ107iVu3qH+kwaXhFkemOfJ6HexdKeso+9
Bg5Hf4s4xFzMraiy1AP0UnadRy0wXA1tDO2OrDWeqXQNnuLzOGrhxoYin5pxihOl
IYtuDii4I2W1YfAJJybJHnSyrA8ngljY2k2LbQrju7KZn+yiWkY+QnC17N33vjSb
JAI5cVgTdcxEPQpH3FyENGEqR1yUqla8LWyQyVD3PAyW9Gif/Gs/ZP5lRSXNHr0u
zgx9Do27ZYTsZGyNIWbixyHi48BMsmoPSltFoepPWUJr+Kio2nP8Ob7teUqqdUaX
3zTVv1qdC0mwYSfM6p8ZXQ89K5yT1V4uK+Es1k6wIXiL6phjquV7cN6SmlgHLgZo
/xxMo5HAH240o+1xl7E+dHTuwv2zdFGlnB37QhxPxPhOK7D0PbS1PbFxeIMb5prP
UMXYcP92up2TroHnYyGYAe1RkV5WnuytHj0Rf25TVo9WEx/wr/wd2w0i0SCryyqV
HuwBJaTlsxAtm3vQXbzvgvPQbFT8oOnMUCIQUJp8mPik0YSzDL6DDViEuQxPQ2IR
LnPP8dKy9+jpIU+KAfvU8I4Xvj0HSzU5AOQWlNkvWSvFzSfueMQ61Ol5+6aA9OZK
c5V8KVjGF/ck5qmbjClJmKipe/0MdAqJ/BaV9/cypdy536ikKQcVKDvsU936/l2v
NbxpS5f/tOyE9f55+uiOjciA9jhdyIIC4Jtpr/1gtjhWdwDPohouveQjkEeEGWgJ
Sj0alLqVp3PxM2D5vhfzBwHbi0t3FJm3DttNBnZ8YME0nOYEJNyUG3YcHgtHIzmt
msY488hEnUg1ZAE+SO3kxrXo9JBvFmTX+n94xcEsue2vhqeIcNTeVpymr+AXXzw0
UkQtWB53aM+0Q2IyQxp1Ey+gsM9qOeKdd3fFuS4Bjlon7p8tay/wv/jk7627zI3f
W97GMV3l3GRAspZHY4M/e1P01gK6MKfOhcrctYif8yzz1T0e7G0qtpPPryXyrgtm
0fadMJQyHMUjWsweBioJi+dv/IavDYE1xBVd0iwwJP2fwSZbhS0XqU8IKfFUcthJ
Ar5jlfkNOOVQTfOi7ZRPCmypub2o7hqzFLQ26QXBCQucERu6Wn8cMza0vzLilWap
H/Cn7ZfBJGSBukj/HVp/2opMwJXus+vtlEBPXhMkpHlvSzwyLda5axYP+Txm/tH+
P7MYNmWeBIV8DlsOXCwcQDzyhNpi6f7b8kvJ5sv3friAVn7evSne94YBhJwN7Ko+
+C2TDDQd043FMJznG5tVKft9juDDfEkwFzDLSVfycZy6FZhf0F8AeSSZ7rAW/gMI
tk8tSBxxSIFYWXzR9Ei2T3gj+UOOjn5Dnz+W4aNaqGdff0DGh6atb1wP6aD/27H5
HCawRqbxK2oEFeGvkfgmiqPxYYuc4xFk/yK1gFKPJJ4eNSTp8HASHSAxmihDO0MK
9egANrl0RNo/+3bkV2AynShO0kZebdsOaztsYV5LdcmRD6oYhlv5/yPHJ3KmvGvq
TEhbsWGWGnAXxkxdfnW3vF67zRLY/SxayNnZZ0FM30TDxKVMoYcEXGAHSrkYHUKI
gMrYzuk5/PTGJA23KlMoJvD7JsGV2HHsbQEGLDY7FMhW5GkdHBK9cWEs9Z+/jedP
LPJj2xOCr9VRQbrmqIXUykjIn1nkyrdppurkjSblhriNhut6UoTz+Cdvn7ThIkY9
+cEF2y9lkJTo0mj+JJy/NUUBfghX4IGSB6NaGudDArbgYWNM8uNp7dWBqsJHU7w1
1BcRZsgXmfuqWJjqqOKZG27K2DqwBYI00RgDpjdiMZ8+QBgWLLPjZKPRj+G7GeRM
Pm9bgFsA7tDD21I4/mHQcqWzIaXX1cv9XNW+D2636KQRUgNIgIGMNicoTVreZqMz
CyPYHbQ7DBvoK8ssRL/4ZxLSNv3nK/AG3chXvqVzJRXF1o0FZ5N/kelNXi9iaaB3
5saQsw9qWD2VL9kRmxruGiTjM7DnO01LoOKhSiuzIysDIfHxm4knscJPQxQ4iA/u
Tll8EJz6FiOODMBHljUnO/82cVslbSTERBtXA4+lSKx7dwKD2dyiKzjp4JkMyPgN
kb8oJ6e01eFYRb+JbP2X5u2ZA3DblOx7gMAJInhw9eXfFPmBJxr9grIr6PRUJjBa
ckOSqgGlt6NCZDBmIhcaWuqi3W+HCBXPK+Hg+forsEOXdyEqgWZVagD+0SMdHEAl
zPETsLQx2VR7+F48UhwTwYWpwqbpb41GmA1EO4zt7BNurMWUcwzSjnOYKD8X4QAJ
NZWi5ke4bPth8DPbK41Tw4C1U1fIUUplgY+/EGFrLiemuV82iP61oBRR+8a0SrcF
ZPLfOTmEMnio5NyIfYdk1FqKGcQDt3cYbR5ZbIEwq7ABbdYFNHIMDjssB07ctSI2
WdtGscTO6PMwtH2TndAykme3VPHM/ADoPBbqrc5BM6V72pJx3nYlsJkGY9bqMkBy
tkFm2uJy6RxuWo5BU/H0gHvIrWO3bQ59/VwM09i33JkZTvfaujN8T7J8/nD0C3hc
eQT38aYsL1ebw4vpvZR4ICHU49+/d5LB5NMeJWQHBzaVVHhyn+VSEwnkjTLBU2L4
xgL6SC1E5qbkrW9hn6P5AgZdi7e5uON79L4HAi1zYWL0BdRkaX7Jhu1AeI1GLrcT
yxf7cMPgxk+XTqqD0I4ZQ9LDqXNMCu7cNN3NSBh+WERgGvsW+wcR+ntCVP3IgGbh
At5beJhfiokQbgzfVdFy6ZM9q7I7DimAegyrpo7Umglj4K5oXD/r6Z88E11OynKx
cNJMvl1W4fwnAkBodWqHlMqtwiN5Mq4R98cO/3WXYWyWFeLj3QUqWcY8cUDlohLP
mlxa941FP7QpRy4bQA/zh/T4MUDx/lbIXou9XxsUY+Sf9NRhjXzsOZLBERyV3M16
dS4I5bacHPuW0HcAlMGoYMbB9FneIDHsg/3dnUZoG2OIoFxyZnpm0DEfyc7VO7Hy
50weehSvHytjkvUsG78j5MjPo/hdZcwyDUf6xc/slWGmK90220kV/WRwNdPmRxqn
91fvjt1Eqy1riODUd/nMxTyrlFUlD8vuGolDTCFpNLKH/O2nQFyAPlUKQn4OUEt3
hmaEwwOzrmiPIf9EaskR05RzrjYf4n9XvKmOTThnv/g99Ex+aGL1pK8W736+u4db
eD9pW/oE6EP/dT17P+1eIOdXSf+HOmfeRRH04vcNgLSD7V8D7pkgLcl/KxfgKRXA
XQWWdwSkwgzxCe4LnJQ3+X8z5yiW50/nt1PyhNL6NjDXbwLAHfWINqjW5A8VILOk
A9LjMcDR695GM6rdlwDaUW2SK2Lq/v5G/BR3HeDLcst0G20YnmFhP0nbvBgeJbae
BB/SDuxr8sIeF5lz0GhxlN+kyOy7UGckRPc5Pn/Yh3VxODm5UlT0WeRAfl1Gt5GX
mtInzHrp1BgQe1cbk8PbqMIW4HP7G3Gc5JF95GMj1dvJW6T2tZyYq9ZONw/OOS5H
Cy+VLZFMWmS45aHyfqRoMtLw/eXpDGx9Gz6lifA5ulSJwsYTfYXErf0cHrUeDP+5
tfvzziAVKC2DJsxPR3ddLTdHgJreEexJlZxNwm28qcYauKJIy3/0+Z+XEobLUjT2
qrYbxWtxImcsq0mypNT7VWKfwvjwgiDbFchNr/k3vBCCQgHa8tUpt5BK9bMkrgRg
f2Gb5Pc4vrI8FnvoujjVE2lxO6NB20/HNHAF6GWqFoH3p2JIKBAXyYOpkPpVgsNs
bv/s18fsmR2PD78F6fS2W3NclejsdBgb0UlehEtflm8R+Oe5Y3WUx+D5nHq42AN6
/TsV39yuYpF/Jxc4QbbUXRQ21iSevMHf+EaJ+smYMRBil8zCO0T06PWCr1chf7ZZ
lDtvphu4IGFQnf+m0oYTc/blB34EFk0OMlbcTS3nj4V+a0rjgPj7llVA7i0SiOQw
z8VbinGJEoJTWHDgx+hj2ZMpyAkMXReHDmGK/5gMqlEIpTQr0GMmr47hPYhRGYh4
CiKK6Z5D4te578vWI3h/wZN/iudoJMDn9IyVGB5b3pRU4ClxkCxEXGqcOnBgJCo9
x/pVxOAXFlLV+7SHhVMgUAZT++qmuHrtDBN71A+F8GV170Ciefe8JvgVrXoLBLo2
ZqlEq/1sZfeGD4KrGJF0ncOXXE2z4i73+HMSrObCdXVeO9QWCWuXGakpBJ7cf7jL
W7ffrFilexgYDkI1SQMhPs6M1ktM4eN+d3rEv/pV5uQG7tJHyvbMkyfeat0LmX3g
2p41Pgs6gjv0VOuyfjLoqN5pwmB5Qj7LwgI7Tg8Sz5OeLFwaP+zjvp7mEuWULD8y
oyCtVhYa5c1MpDFcr3ln7ujvCd7MatUasRYsROI4d10bqKYHiJndnwwwU4hcw7gT
pPYcEuZReH1ugThykWpx6pW/yPatYd8LWmqaNcgZ+9e0GTBUJXKVa9MXbkrABmkO
Ie85HZVHtIkOq7nIczzQ5LEgfHx5WGyRh29Hmmeel/AMEV3EAXchwBfCf9TyvlPE
rbsq/eqcTEoKWSIEFiW4oL7Ae7KmsF8tfrVEg/9dvk2cRY+DVdR77fZ+eM79MSWU
+NdQEydYG7aEKHBicHORvwfb4ClLBBKMrAzncEh6H+GKbOPvxRG7rREjQ/KzHJYV
KTz8gd9DKRlWpBGSTyZ0odB2Ep6Ic+y28oPcJkZ0ELz7IfdXuCGkF0lRE1dReSjd
9O2mva7t3cgglNGQVjqvsEAFNCKappzvNZZur82lkEWyfoT6gzeItg3vTYhpSyqm
ylaSONmKTsJ4ZQgEc55MC3rF6ve8ovFZS3jU36yLt79wFx7IB9S4TK+PGBjCD295
2B3ovyDJcr/qog016o73Rx2JYXhWCdory1LXMV8A55/GSGrWwULb5kVFjsqHxtGm
pYQyvXujJ0rD2xBFl6NpYaI0BymUhNISLm84QnAeG9j1Ou440fhJju6MFTvrca3p
gh5FN1TeWQ9btSOKUA4pxGxMgU649x/Ou3kaiICsI0uXu62Tki2PrC7FQp0Y2ZAX
J6xyquxu1N+i6I1ekvkrOVi+dSu0+PKz90Hw96XFplFkzyirjejdj2qFKk+WAJ5c
vpXxLNTNKxF3MUj0gkKYQeVbvRfEUCoJGBc2iVvX5LEOeqb+9vtc7lXNIDAwPrpV
Iff8wTYi2VtZhqLT+FZ+Ve2uMlUdlhWkjFHVhL33j1dhBD87AYjRVcpY8JwnTkhR
53z7AShMZXX5gIY6Zk8uN7jFX9kOmYFjuEhtt8RI0tXn7NxjR+vlEOG66Bo1yMZv
0t4pHPTF5tjElcE1CZ5t0MQ9q24qafD8v80uJzM/Df5V50tu2/FShgFtwsjdz4Qa
aDrkcj+X2zXhs6zdvenUMpZSrCM+AJN+S3xT3CMgcAP+QeAx81RWeisN0Ujg1Zw0
osqbMwJD1JGL6e3yJpcQRg1qYFow3l298oFlMaWyy7/c4AkJ0X3bf5Yt0FydFtzx
JkH4xH/UuIQFXxYmc9M5HmY7KAzhipIUffWj2RAr4sV5jIaIOsH4s4R1pQtFqIzx
8iY03b0NX8zscHYSh/AntDvnM7FgAlqeDU8NsCBhY8bVpugBLIbDmoFPZgI8eAk0
XPyEp+YjhxRX84SYnULXO9sTsXBJ294t3T2CXNX/LOwSzLwnhAr664pHeLsAykI4
movZ40d7obOLYEK887uOkXKULBaCYfBUTPNyTl0SV1LYm7PYoPFlNbUX1j/+sFgr
dxxPCCcRb7G0DNwjDVQcQ2Tg2ZSMLxAiV24OuOgZw7B8erKoH5wkk4eOJ4SYDZ6j
IZ5aft4R+g4A/cDsaUchffyu4LwLWGq6q1MpkLPVK2CKWoZvwyyzm6n9cHluCuYh
GS4O2SRD03yDzmr3JTsHdwZ3rmyzZzeh8iTIDD0jfGW2cdFuk9rct1ssUfau9i3c
i7QUaKgpCSnGjSOy6Lk+XhZOeGWf+eBuV+iSrWy36BnLk1nr0yO4M5FufJAL8o+5
Mg9tIL8GYPTRXrx6yU9wWzSGr5trXr4M0oETbsqIM34tRyv+IUK2i0LL15ZZ1mOd
4hsrMZoym5Ake9IrWZnjEQ0YF8QKs26eNlxURs5rbYy/w9fsShHm3EnLk9FIUltE
gf9TjoVRoFmnyild0RUUbFy8YvORczXVp2+rk1TVDM5Jv+q0n75ZryE0gZbS0c77
PP6IXOJQk7iYi9/WFHScysHtsNV55pbIkqmarvHtndpTQBcFq4QZdwKUl7pvE26v
dk6awizuly+ppk69vRGYxRcDDx22rRVOzMS3mZ2K0+W0q71lU7xMTFflsMbtUpuc
aU7hpKdNNEhM5oJ+ZseI03Wh8iiYKPtJJKRCoVCmWbJKWw40dAm4m/dL4ra+T/3B
zwtWMQTbIAXI2tIDY1VG1NcnM4BKBx64laj04W7Iym/8L/urSuTacHiKD8/pHPsT
wSocuMCj2BHhnVlCrJNUHC0x9SZGnzwwYf72bDsA7svkXAl7vBH8iS0mBozT+kWM
vlYpBVLPQN8/QXrpdyhSotSP16VTGJdvmOv/tMOmIh+hdoGh4MiL447g/hX07o+F
2lYi1AHPrt1S+FzcTkz0Ulwqjr3qQG0HjND03D+i/Fm1Mdycuy+Wf6EqcTZbT6dx
08nfJMyD5/rgBp3vChYY7czh5MU1YKcVZOjx/pOnpFYxafv5v5Gs30C/q4tU629L
Zv/NJ6hpHl56NC37GolWzjEwdAuMNcjn7036K6BKDJqp3ytqbCUGrbjnO7ma/T/S
U6OOSSr3jWBzda5Jey5CKMwuLDj8Hl+gB60m3jqCHCfqADulbMrQFPn+y7zdn5yo
LHJRjRFE381vpsIt33Je+uUwyWW7aU21R805aJkW/fC6aCNY9vqkbpfQECKw3SNO
S/P5gyVw5WoDdZxbpI7hf5NTFr/Hkh9Gl37ZnumRU0N9QAEtzOCBiZyO/r5nymxO
iHqscBWg8ZKzYRSEMx5E4WBukOL+tPl0EEFrgdzH2Tv4UAZPjlIBm+R+5LRD0t1a
pAevO2PCxQDs/KqDy3HoytyIHQJcW9Jsix2Wyy5PpSirpDomuAG9MjUWrHdLkp1r
QIu1WhWAnvhGQdlwUwEK9V/V47OK6xTlHa5OhRlODzY4Uw+IgRL0iq1gjR+QsP2F
vPZ1lhA0/NKN/WXqTnkZ6QgjHwpiXErhrEKSLDQkTPkS9+xDJD3+QWwiAeT9jZh6
tdSXGqS/GAhP0YN2Ao5L/MeAaNLNaiLTYOnjLoNh6Piyq/UYxmUrLoOiLubD3Acq
T5G3PmRvOTJUsIiA63wg3qFmcwnkJtW/37xUjpV/qtNuHzZvbDLjaMf+Wx8vw0iJ
3m82LEENIixVaTVP4PKmqkCs2ylxKNutqAI2m9BCnC5zcFQuck3Xobr/0EXlV+nt
EeD9duXKGGKmKPSiKL6svly3FMQVG5vWcgKdqlwFhq3GPkCbgjELQUqQCfzUiqIt
9blwNzDL/FByZKlpQvvjCDP9L2umgVXiVE9h+QUerlU+20wxzSWWAeD9vNUjsPnF
z0kNHW5K3IW9D8hZErV5a7JeHXK2FtzJOYb1eQjUKsdvWQV4TdGcg29tY4KpGD/e
5S9UhHj8M6fu7Tlmg84gyPpsMsdfRygAc3rvSnYRIoGxJhSJXPBwy2ydoXB0pQC/
o5xmRdFZPC82mWZ1AM9l43/QkLK3667gO7RYHuieVY1Zmoo/l0/9PlIPIKc8tVAL
EGtZDIRwyLWBljKrCGBguOWt20zQvIQZR5QR+scrP7iMIC6TecLD2CKpGuZ6dl0S
pLdt07NH1K6/CBmGbR82dPH6r5fte2NQFvto2VkqCmNTDt3UbHgMCnXV+eUubL4G
y2b2cdfebB1K+2yLgWiUh2fqes0ANh6B+jecaUZRxvQ4HTf7pohMY5w3M3GbHQx6
DSC1hRoSQUmZMAbVWD9Hkubm4XS6ioPr61r73tvwMao1b3ne2F/miK2wI/cTwn31
iV0//+sLTSt8SeAw04irlx43423POOs023BvkfJ8hv+cYoxeEaYsk39oXeEqOy6T
fi+AkMapOhpO8IRkxQ4rWWRQSvlv14gJNolA+pNhwYe3JsN1YTjUnS4TqiUF+9Kl
pOPhAsu+nXKu9JKyylK5I9q8hrFkftebscBis2DPhPhPf35WyQi52TVzm9yq35ed
bKu362kwmIlBBXSNoa70sxE6wCojrBmLlbUKgFKG2KxgTW8GBFpPog2o+huGkpCe
tW4jEVDLSN4WBBwMw+AObMD7h9j0wx0C6RLiD43R+9ZlqDN6OFy1ivhaHeWCCtjc
C4+bqJOEcLrx+RqfIw+eyUkRmnVmC3xILbfWk7mB4BJinr9MMWdCbRzcqA69xiih
lvlPnJrxFibd+2QaCpS7/jI79b8nscMNuXtwkW/C4nX6jmPFBAIMzW2YqJw21Deb
AOvlh85jInJ2O8MvRI8x9VDQHbTG84iNNQP5z/vL69mgPA1ejC/3ahsk9hU7usP+
Ktrll3RtfJarhp1g4h5R9rmeGa6JKzVX9ffvsVpeQTS4A3+Jbt4JoVDc4tvckPkD
fuCI22LzzFXj3XSF1VKC5VZ8i9nqdisD5y5U9JXJNXAstY2m56bv9rKwwT5XQqaF
jVfb8jrZBX67V6phG2Mq4/+/LvctjKrFHiC+4Kpc26ZOStOvmEcbkBKaBHiayY7Z
1k9AMlbMTEO4Igyn/4SnPCjyragaw4uNE6Z66ZatoZZxGxiKxLje09/m5Bz06pa8
bxJhZ/T6pIEBLHfd/6b8F5UNwyyz5KT4hrtYg4n8r++ALJAaLZ2ojqxxQqhSMXx5
le6xOkp6Zk9yHjcZbKiCY4xHD8ks9TjJCBTpwTeR2RkXjBnWeat/tB60rTn17sGU
JiepddGwXKt/EwYekHYnIFZ4CSA6rxFi/6E/gI1wGQ9CZ53KVK91EgADUV4IWPMK
wUh2G3ZUnQgQnX9hAylEFBJdoS101iv7l/Wn6I6qwjD7B9dQrdtf5fzQI2tJr7JC
SyqZDfs+rzarMOSJSbYGhAQUcCmzfEnISFMmJ5PLMfJcVpLYA7Fno5QA88CPkxBN
hco8Z4cTjPgEMXViktL4B2ZNNEu8jA/POXbgl9Nm81ZQ+pRAX40yFsFBiZq3opEs
Xy+2hC3NwZiv8LU/xqXVklxH1fi3V7YyFFYbxeTYfMMLOMwUds4X/Kvx8NYQH1z/
SJnLd4KC0rDhvBeOIahh+WzhdSnuhmws1fYQQO/Dkq1orgJA61nvmEmv/Ndwa/12
08x1jDMSfY/5+azO1lonRmBr7WXVQOqPsulT/LziLDtH1NfYR9WaKHnKGSHfoVCO
ay3X1Lfbjj59ekFyGf6qKYB/+ARBNi5Ol9TqE3WlFEdSPWufYjP/1JwyRPeEXFo1
BqhUT46UmhBWRLgmBI/lzKCaBrdRAHlODVi58H4+BLaz/UsSXAA7tQw+VIvNw5K6
FzafMn+6GZfQHC8uYzibIanUe3/ukztfj4AQK5WfFGVYjxqXcCYNRIgLcvTt4X7Q
LqN/eBaHdSOuw5xxVJLiKcCYKWFh6ijujk0owViJnZw4ZFGJXStNxMr+5cgHCVl3
QltOpu3tq323IiZqmuFaUKMOW5xZGR5VbPD/jQ1Y1Nx2YHdroi9d23KnVrn983qh
kUZt5fmTl8kfn/NUDSYPk1x55MfvtZu6FfWA0qg3Xb4zQX8HUk+TBvDY3I/5KqAZ
lPZ3rxyHb2YcQ7Ip6aV0dqUqO82l4YXHakSVZPUPXBNaKhKG+nUpm77hEZZWc+nK
3/QyH6YKm1qL9s1WYaw25lHP0nRVMCz9YA4fgt7pecMUivmQOZ625XO82B5mflsi
p2snLWW2M16Sg7f1cxOBQETFnnKE0rWSASzWqHySHz0AzhJmWucPx0VIQ8CsoPZ+
oK/oUI8hD1lRuMkz6djhYHpw+0nRsqhAfiorMNXC0uPNUK0yMYXsPQ1XcETRMhO3
YwFFbHCf5s77NDLvXSA3xcwJQBrr/Ba2YWkWpjj4Oi+m+DvHoxA/n0+9RvrwdsbV
LzbYOmyXTsvVG6WjZyDZV75t4ptVoTS2VjsQ9V4pgFCKSQf9RJ6MO8XbMK8GzX4M
Qs/QbFhD5eysk0w4oQydpX0ODH4jKZsQ+F+8toiHnfZlY1zS2sHKIXms1h7L78Tc
AXi3LUBnHf1JT5c377Kbnp06HHVZaf/DtOqk6yzZ3ugFoyMVKvox+eZnmQL4LL9F
rQExiSMuq6IVpG7RAfndCuNpym0cGdJlvT3VuwOnsN9GvXUsGCl5cOVvUxfHLoUs
wUWf/3CDZgLFlXZrjhgfyNL4hvU3haXiMKslkXIEZ/Ylf1JMfEow+MvkX2Qxp8Iu
DPEyP/7B8dCqWS+t98MvEWLHQVN83OxvKx+ynCMjHbXooToxcyBw9jIem/0oMU8q
kDnnMc9uA/Zk/BN0hxyL/y0Z6EOUrgeGs+1xaheCbo2KU3FzKkCDskqpMbSoBQGP
G2H7CBSF+HCNBwfpekw91tQ0N5hfowxCRaDL7OOHGUdhxqwjzdv3wMWN3Hv5UYDE
t12fz7caFXoJPZOEE4bRGZaILqvnoRgn8beaKN7yUroRq8ET3aJJ6PMuZQu4pgx8
U8X0AmyvQWVGrELmF7REQXtBlLpJRQeTuxpzzkc9bOi4jFFEWrd8SH1tM9nSemeI
8ZHfRwDvgB+2/kr5mSzAZwrsElzsP5JtEIwerRntaQQQwFJo5qU3rd2Uf772nXEt
0aV6D9DsyHwFXbK106OEqJ+1o/6KPfyx1l2ig3MnpfY+iEwVUqOn3FKlTmojFYps
JWw522mLPgiyy43ITfe8+93Rh2ljoBpmvTagLbPZ75HU+fRIRWb1droVd+mgpIsG
+APm6Dw4D8nZZJ29jk7hhZvNCPId/55QmgrPBor3oIOMnr82PfdQ8kS7eiZRmTVX
l2j8nsV0Yy3Ov/aydg8sWQh7+RIJtgUAwBniL7usPRFr9Y3no+oP7lNbknVdZhGE
pY8HrK1k6iX1b8pdmTjA+1E1DnFKdBHAyvSTkx1j8O0efef95r0xxkzfLVpIq6T8
06d7F8oRIRYnqe52w1kGnwI7e6wBGNyoYChx3An0xTCbZvjnCfzqL8gFfxx8/acG
4d+MFj0ADo4ALEA2NqB7E3b/w7QLY4oLTh/GSWlwVMnGWabhmmiBvX4gQ4Pbg/jv
qspMUR7djz4WMuuf08cJ6EPDEeago2d6LnV6D7N0RtYm7uEuWXQ+O50lToilHuHQ
L48DWdd1rfaNoTQi5G5oOSD9BTh0PggE14oJFB/yZKBTcJHvoYPNVtrVTADamcN6
9eCl8+W4a+h4hw728/CW0S3wp/XR9wj7+ROKtf04yDXMRGqWaypBVLovkbLiYJ/Y
5B80MWUtAQuotNXbxk8j0IkkejoZV7DKNryeV02ZPVyxlbwUfLaqKI/kXXNFx13w
oTzc7ajzZDK4rEWnSj417DiNEhWv2IbmBVwCGz0FvZw5CfLZXSXZMsMeaiqSghdB
iVadu1Bl1DZsno9hGW7+3eR9U5A7ZaLlkEnTUYtuWhWFZdE4aoBPyS6fAV2OfuYK
2/MwDHkT2zx2wb30f0rOGL9rQU2xsKn76NPXSUYzS6khs3P/BX5mkp1ZQ5SQB7/N
hhEZnfDpb/R41fPwDDCxLmMLgWkp6I7CqYwqMN9FG95/MSs4VMDpxFkCeBEGhmP5
kduOHsUTJ96Fbwim8OU/fUJpi1Vg220evDPvPcoKDtccbL2yRViWE77bTdXqA2+4
iGBtqcRlqHx+WMXhhuqWLxcxu+EK3x8JnSbFD/adijEnPA6g9lJHkxYvVC9ZGCvg
1dnbqiBcW30u/d8V8Mnk7z6ciOGrwQA9jwB+4LqS2+Rp/3XJmcAIqTG0X+Ok9dia
PIyk19ou7dV+M9ICfvW98RFNnJDTZ0LtOPCSemHoJzTijrlw60KsDcHfvgwNaUQi
IVPZeQHY5fxPjFECe8qGyFSrrmb78Zm0/Dfs4FHs2tf9/mX+jwNU7zI91njyipHf
fuxhNY8M7ZBvI8OuMYsQ43VaOO1mRBng7fm2mwX1K0qFpIxFPtiqC/HeeWloTZ2i
qUuU7ypV/hrJduYWJtZbSl6egVM1+yA7jkuml2RHUhpN5gRoOyiEkERftS2R7GIV
boFKf7MyCEf2ogQzHuR3ZYAoK+oIhQCJ3lcN03ym5zqmGJT4FFfUUknX5ArjxeYJ
3wnDlxVU9w5hATxq7FOZmCRi8JruuCOH4PsFEDwVahlXm83wrWkEIhUWU/DWqWlO
VSFk3nIYO3+4vR4pRJNKC4NPmK2uAFnYNJ4eFigRMc74UvEZkYUiCuGsxYKyIlJN
H8BnE4hezYJHY/JD+hLxE/G6qP5KzP+chqk4Z4GRpgHPW9NEFkbrLX2td0ijavfG
OPBMG5BF3GpyI6JR16TLS72zN6dQQF0+vnnnRsfOsGYbBA8asuKtHQDBZhLxkzL2
ROduWvYDxdVbKBjpql703bo2pUq3UJ9eNgqI5rd/QmZNgYAIh5F8AsCkW7lIssRR
vqW/lPrsFVzSb2DIlb4RNy9h554UDnPNUbT4emVpJaFgwIujpEtpfF+a/HwFDBr4
pfHKhc1wF0t8Uq9bnTcdttwUWLIlkw/Duec3EsW1mhSADlrGb56LmfCCgJx7R5Rv
voHbDvLIS6SUvuHZjipOKxecNN36dbD1VsacQtUKpXHNP/bcmkXD8+2L46ESBUmX
7nCBkK94F1ZKisy9C4ITh7mcQrduawvPJoJK/ZQES2Cyb4wIDqNK8m2kVenX2+Ht
Xa1xtiKTUyzHyYnAM2sxuf6ApI3D4XBax0cA3Fve/Py2l9p5JklmgexCDd+BBCAa
+YAiiF/g+bat9yIbfmgyHy0x6oLoF2NFZvEVr23Gf75SX8SjTOuYiEmdQ0V0y5nt
9n9mCLEFEtjwjQnWIM0TePxbaQpU4GySw75ogGQPg/KwnHb65+HIMKUlrBxqu8qd
c3gfGCDYnc9eHIUxEFwju/DRAtdjvq9/Hif2WGegCJpAT2/H5nxYMkJSQFXCa2lB
bOLGP+O0TWSmgYyf5pSddpwFAUJq+tUADwF6Z/PtffAxuBYoy34pHcHVdftAoCKz
jRImr2YfVtF5SJMyBmcCrbKkV/MsX0HkYKAyHuZb+0V9m1eBkklhjHm7ZW4xP5ok
1d0v18dcv59Ow+1gl7UWqjdXKUq2yzWq00mWfxa3FAj+P+6yhe/ipJAczN3r3Dyh
8EJaLKyhqIKgfXvEaxhQm5JzVhHG7yWXKGAF6d59j5vSlE0hsPD1NgptGSWWEzim
GHCvgc2+HVyZm1+8/BQavUFZg+1CWCdS3eaLV5wjLKvCB/w0HagdUHEk2OIt/YTA
T8JZwH3TBCPPj05usuJnvK+4GUWkxvg/BvGVMPjnHEwCT10fw8QbmPo/8MFlRAtk
ei/9dWml2BLRlQkCUphRC2dlZgi8FbQRIXTtllvi2tvUMRgZ0PimuDO8HOmznj68
S1iBQENXXpKR52gt4iIBLe5ojJ3gQFTBB3zSGWxJ8CVIJqAikTQ3YTY0zAAV0SDq
Hgpqx/3eWjiwNxGagBDgg4q8jIh+lr0BLb968bwoc/jK6obPA+mMnY54r7d2Ge1g
BS+7jDLEj+u8KMY5M4CqsKyjkqysZErtQkmvlcZrOHH/uEafva1pOitkCxVDEQG1
sCjZcNIebfdS/y4wXr/igNI3eyBLH5uv+0V30GX/CGc/tTmjs0j/3LDle6WTN6PR
pv7iAHgEjLEt2wihwYmk/HTXmQMZsL44dDuQMUSK3UUblz62LNMBZYvIuVpO0hnz
SKCF0ynohES+sdEYdA1d83qi8r5cFeULTj6hWvAu5G/LmtwC/XaEDnnnnS9/ZsXx
YNFUs157x21Ll3R3iizic07TH8TpgMWIwApORVRAF1iTrgaQBk7GShwiv4Tvha+5
gY7vgWIKBV9kPnDcd6JcPS1Rv9wNIgx4ZX0ypzr+7ATqMomV8RH0kdLReLnQI1FO
zyXJXm5AeRcpXO/iLErTWmgwUV98+Fp3bZZ17BTEBXN0SBzRh6jtK2EJAmYCFSbB
IqfHlWsFxnivU5acw+ehKtG8myV2wtO1bn0s/fWALiwk9lZU68kbfG87Vlz/8mkP
bMen57D8+HZ6awAxEK9Qa/XzUYZtqP6GtmVQZxFI1JlqIzFZC06VDmhz4uNxEQbo
KEM/EUnC8vN1ZS7zfTgrFMbMnYhUmhUN6dqURXQAqA5QhJSUjpdZBXsZq5LBmUFy
NmG3OyeNchzPvghwP/Mfe4KkzxNBJRmXgVS6T8Fh6+hySYuISgbhr2+t3iPOavLG
o2DbFU4lIwLidc82Sv2n1ZyzlRFEr17dPI/bBEVfIb+zivNLNqNPZPWWg6pqPFkA
LIscDWEfeXqjlRpFgQv6RDwaBA1k/YYyVskG8BKQnWui9KRnYVkB1FPclRf/Z+CO
bYToS/zm/M7UDIAvTTNyLmBbawEQigNL4s35zD8xtQrzIh0stfibgB2mlz09f9SI
s6WDPfN7AP9gaGm/aF43Xy945nDYi3JdicrkN8n7tOKJm45K205yGvAufuD9tk2B
QQcoiZ7s/HAknGJVDdyQUM+QMUpIwCc+mza33cFZ/dBqGWrqfS+IYUJr6AovDg1l
3qeosQzUsMRLzuPdVFSPnyamxwFmGjf5f/W8E50JS7GHr/5flE14s8/OhsWsPW0K
+8aFZW6oDARLyJx1ckoeVS3grtZ3kbjf/wI/YaCcCJy1Z+pf28c32a9gFDSSEW8J
pZ/2+tiKmUqIbvYV13riZcEWHDw3Io5jANq6Ybifj9ph96tIAJod6Me73eYOpImq
MYNZTVsGfs2Ug8Qw/BCy7DOX5HpCLzP+5QnITM+XoAte8n9EFa6fMAzPakCN1w3+
/KI9XfvehVkRc0P2qQOcaytvaIuICB3AnwfGl0m7KAuw6jKUipCuZOXwnDEX7NN3
Ru53moAQvOO3TwPUbGQShmCOSjN8yAs88Y0KTcf7EV7maFuWAZBqd8vyLFqXuoUj
nWrP+b66ev+y03V6DnzyzUUI7YZwjnJyl0d3umxNATpRzasiqCCSFOuhDBNn+MXt
0dMut/dLq0c7VyWHZZ5ZH+X0+pkeQTavkrBYJqOTvoSYlYOjTEkOz28nvwFlqLwW
T1EhDF4X5SfikiXpYX4j9sQzSsaNx2WwvQRSuXjctfsXMr1ub2B/EDjvPwJmQVnj
RP/o4jJwutBRniRVbCOheYrz57Xp+A0cTS95vsTokHiaZi6ZdeZ5Dwv0xFAFPVv1
jrKD3ACvKF8TBBJFsIWUpZShiZtt5Fd9+wHon+oxgDgNXMZVzH6ZGRJxpvixDex4
05FrcVGItSMubUpaYN+0uC6qnMNbzLGqtHGjICyGY5FEcdP3+NNqF1ELt5WCRqYr
l0Af2nqSQkbs3kvCa9zHGO/lVamgb6QSy3D76Icz3H8TnVyvnEK4clDjh7PQRpuu
05qNqByCECxoGdZMhJkmlhhmJNRu+vsnxkUNhEO2eneYDnCRjDm+AiVCncXTYl7P
s7b+PTyVNdQgxJMnYWjAFDuu7caUL4X3p+T7SH+8HEDMQa/Typou/QuEnZOLIoD7
CVbokp9HBkYcxfSH3TkDssam/KKsrJREUmx7CbPDAt3QFlLTGILHkGktj0UxtVT5
t8/UwfKirsReoTkPBwBaQeicMZQL6qvAOFuGTk2RJwQfEURixYoTshlJa1Vkm+jr
M7wCMfcirnubY7Zn7rh1dEuVu88IQ0yLm+VSoT/FxlIojCkkq4fKHlXBZM2jiVOK
TrKUpH/ofiEa6YKGQ8wslpzzIQ28/D9hrIcqLS5GVIz25DJlMNW/KaVjDhSwB7RZ
sEx0g0ua5H2OK1mKqYaDBkndgJeXuTMX+5KxUIqEK7RaQzSM4xRhadcttf7lqv4N
PXysn1G2XlpfNaI1oM0ftOu7oANlf0wJ1GlprDtko0j+LmXh7Au9jfNxUltbqSq8
InjFf4LbHUJfBruExOeOeDwHjoWVaCSjXCq0EPjHIlx170UPXJb/GxMFFapzAzYC
84+QKR3f37q/jigo1GJlZBMQyIka2ljQ24JvIhaNLjQF0xEYNSyW4UF5INBMeaJo
UNmr75M18/7qMC5EmDw5Z5bZaJAgiT19KyOSl6zt4vaAWcDZdx0g5pUhrD2YqvzO
rwwmVw9/d2CXIiI+HvC82cvfRVMuCKVWNEXwZXhC52XDitp+04SMy43ypOnBP899
vM8SV4z2XT68PfIjHYf2rHxjCFeq+PhArHP6DoutLpdFgBDCNFTVslwpeVegQvdI
t7VANQkswomGtwbaALotr0zDfO4W70FXKM296I+rcCoJze6FaY18vSPuaQ8l9VW9
nO+yUNg2hPzJUI9kZ9vUQ8c3a7KgZ/mX0cw5HV7659ZOCGsiugIurlqI6Pfks+r2
9LtYKoSKySe9fc3vgfgzjKXAaS24QwGAn3PSJfqGRtvkIhIsqamQx3KGrL5H6V5Y
y9mqEDb59XvLd6qj4ZxDwvcfWQwvjziGbkliUzMH+C/MdHMUqo+E3ILuA+9ocSbY
l9niCwRQKTQi+IcQ2UfT1cjuYywYAZ5ezH1cnpw+ojqst8nRTgLKXtVCuYJ8Pfpk
MrolAvdW9Ao6fq7zLKnRDdZIwlVUQuY4lwreumFAQVjGZR6V/qKAJmGjEwrUJd+F
M7EyG9M0ue5+K4oWi4QdLZVUrETQeyZa24TbXQ6xR8IrB3ivQ3rz5JA1fC4e3hgm
SHMyeN+NhKs7X8CxK8I+NAVU2rM1KA4pYeEPHVrQsHXK7/tVVmlVhj/3znI6R0nv
d3XtCwgf/jsyilzZsEhIV5Pfg2v73pRul6hKdDXtgj1BnzndQ6jjS0e1ayeOSeH6
SQeQQbt6wIAV7g83mSEx+RAlFAkz9rfAkOdZmoeqOXVcGJoCpHWy/2b0XyMQ2ln2
RNv++XCoB1ZpXg2SCrGZlOJmv6w9xHnmh4OB2u7XLYl2k5kmnL3D2hX11WGqPqv2
Z+6gWEmuZTUUDie2hId26EkSSSOJY0llrM3FgIy/j3mHIp73Ff38oNbmim1f88Yx
1Cv3jzvF+KKjL2f7QjTHKvR4IPEzJYBpqgWn4vENsKTrs8h9wg+LF5zkdqGkhAS9
WdWpQpimGrpVlJ7TvnS0LMDBiv8K+xTln3ZPo645nI50wcxsi2rK6x5bAWAVsckl
1fTBUga4XTkJlQvaVL1HxF+k/M7bLEAP9jOPJvhuUsGmzwwt53gAErVdjjJ9OLln
HaDMva/IMyUSFRPhBd5OeydJ8cVlFDUOEZrtiitNZXEGPtscZdlkVIQSVRv5Lh5c
bhQm51J017iFVlnvJs93CAKAzT+vNkRt/DHyBUsyzFLpb+IksvmYBIeQOKty3uDS
2h87mM3kIQ+7ZoJGZZzTKA6hXNsMC07uE47ov7YRne35VQA8gO5L1h60BR75mmO0
EyE5M3DDGnKeJYYLIjFuNOtrnycpp488gZkodcGKIpUY/zvGY4LkkcGm8xdcYdsN
KL7otwDM8n89CmeOFRxBoASGZzP1aZ49gr/3jt4Cti2CcXcxiZy7G7WTt0YKkA9l
JhbdypdGqogL/9jRnKzGuCYW8yUH5I4KC8njDbzENZgrbouIXCf766tql92k8cfU
wOfMPSEno9vfLxLo4mDkGIjGDJhnsB5MB0l8c7Xle5ip6pqOfW5xvZNT8zbJiDhB
l5boENH1Cjy5y0mtCqi9SDrhJqD/j5FYnuReXSOADSzzmuAWvenyoRWgEhqunnzZ
tDAid7nLWwse4U/+oLAgXeTWvlI25kMGtAfje+7WtgxdKW0e6Fv0+1EWnlWzgK23
YzEUDkkbBEVLrAQVBY1H9No9bYKw9j7k7LhQFSC0+HlfrnTFmGj9gVXdTzUTxIqh
UePW9Ic3+JEMrgPsFgdsUWJzUurrYBVcjPf9htMY5cY9906jW+UaYiOXqgR9yL79
GUiyzVIV0T5b+VBBL00pTmw7FnCwl7MaMCaM+SZ9D0OMpg3EZ6QhIIar0TvTWUCL
NFLwTnGAbdnzL1eNcXglcBlzymhBZSbot3VLehp6oyhtAyjQzazM7ta4zY2aGjTF
qkZ+ucqp6SAL08fMdq5VRK6zmO/6jBWZ5nGdc9HEo07ZIWGx/IFtL98GgeBFr/fb
o0HONf3ZkhJ8xetIHfEXPGzkkjaCJVXR7Axe/2pNJacBeza80SOQE0iZ/IYHz9V9
8D3m82lv8kjjKDwGPUZbGpF8j5byZN/DIzYRduwRn60sRGjoNMK+yfbaMeHm1c9t
7ZrbguZDw2nejuRHbzGSUvzaQRR8M5e12HdIFBVYcsuIbK/oRFqgqYGdbKy3UQqX
DTVgrcBROm4mVBUeZ8DjmlqbibmLBch07SSFQawiQUzABB3s3ib1WaaiBm3ieNNq
qGicrj/aNqYsPUwFe9Nd5l6f86sO5PI/gncy270HQ7ffHmpxJMJJRHFys9cXsuCD
5CIyJXFcoSehSHNY7l/bkiVWS+cmW9bXNIyEWLUud8rPq+oeMlc53nUgpqEBeZuj
bd3Lt+bF08+WXaWb+bgskAUct3KbR1AgjVonyhPxDpPT2k81dE++uWKbQ4YgrHTL
nLTp1yRqDcRv67eNQaZtZF+2Um+GnlCY1NGpDJYpF/9RrhOPKXri92A102+l5bGT
r4ytyKq+fJNF1cxADvPejH47TvXSSDy+673yr+zSBlql4NP1hP50T45UOcO73Xw+
H46ZTDflRV3+hsVceMUxRg/XSvRYl0mt1ro8lk8mQPjMefEhnU7BOJ0WYHmM8T76
jDEUyoiFdoKQ1LrWZ1dPbN/0ZPXuG6rOKXQuPMjIrMtTVjN5K19wB/ZkVr96qhsw
Wj86HMufMvZmmh4sUUWcvER+rFnlSnxz8q48mU3ITw8ypsH8RZ3wzf3G6s6/IiGg
8iLAEkaHCqa5lHGqFaT5nKLQHICkOo4wQs0Ck7XvKqbLeK1Upr/8wpQClh9yVrAy
RrzLEMF1mU4jCY6DyOBRj5PU0J7iggzn9gMQl3bG+WiCdN1ebcTONy+HF3guGVPv
pUwqtjttMBKGJ0pnvlM18h05XTVu7xMWaQ75igY7Rb4fNwITm1/D203G9r4Ok3JC
woUD6K4nyDZb7C+9gAM/LOImFXtZ6UrGWVLIxqcDgqzc78Md8dzOiY5GO1yS5EwD
Ye6xGQuozjqhZru/QoCuYXbQDS26J7WBwmlTTBUtx2J1BJAKXJ93zCn4B4jM3whw
E1RZxa4qxRodx0Odf5PxJLUZZuIl9qjdLkS/kUACWS5R/SmXHNjs49hG20dBc5su
kuVLOTpRJBNBfviDPku9dXnb33s2qcq9P7a2Y8sg3JoQOhAR/lOqri7zkjX04wQM
aFFgyn9hzlTa0LchVfXYAuy8DTv7OsZqpSakFC/PZnwlLoJyeoBcZWyN9Qko2hz+
c/DkgY1ic8g2KG/uZReQ92uuiobvdvt0azytFDcPGgANvbvQVRCCCJut8Nsdhkzi
9R/RmQElebs1w5FUs0v/LLGo9Y/nsr/5/FDIjt1K5GZ4kJqrg5KNwKUiJw75C4rE
PAovjL2Ru2kbq532wVYJNn8Nc7xt77qYfqVvkFm+eCMzsd4hOizkr4h7Q6BfkBfV
oEodUjtMoC8P7RPOgAnMx3Dvh1Jdpzleb4wVex2rwY45M2eFkP3fHIDgTbP2xtNE
eDF/lxHE4ZsBhiCFtgKnTwg8HXVo64IJ2P/iPSc5ERHDy+XehNmsm449Wyib3TdG
V6cDczCkMQS+4rPVGmGBhMOWP3+tNMf8DCW51BiOTbHk9DX7h+A1qQPTyZw5Fuyh
8gsrzC/3TL2OVgU9a/zuoeM7OATfbG5ZiRfaZWcNu52VL8u8DUxOjxYe0G42liNH
8H6KUS6UgxWzj9y8IB01ivNPrgVOTJwxRrq2btqF0AJzgC5nQxacNeOHGnam3GNK
mbXd7XqkcAPfEm4isTk+QWWpiJ7ki62EptXqtGfFy1c2xJJFPpv1wqDmrWZwsedf
ZUikmWMT8a/Nc9dGgzIw1Qf7cM8/WWGhKllic5tTzoNh+vPONvkrapSpJanMRHCh
O6b0Ufkx0s6v/38+QObYR8EtlnJMieMqLKMZEzrjYIt8JvQkYOhd3xxnfsnkkXDs
QGjA/JvyryQJ/wmozkfLwqpb4v7msspIvS6UvzRxqEDjRoNhPXRsd5JMiTqnY0An
J4rFIdMqzMt8F06IYQGYk/cZVy/BtHfdRSmRvy59tO5EKxx0WfsYr1Ej5rayvUuj
JgEjLo/vkve0GWymzrB6Bp+6GWXmhJF1cDI8+lfbKJDYL0HqiKRnTtydsuRocJrB
30R9Fpr5nQrQZwBUD2Vy3zsEv99ZGnWhXlBlwDWfxVM55PTv6yRQuR+09vbo2642
kn2Pomw1kWnF7EgGcRyMHsKm6RfdJNIxgxKvHA7WEe3PeeziLuxsPG+hAm9LzkMb
PxR07Uc6fRzqfWRxaovHyyRjjkD8Ep4F84V4xn852l0OE8mzej4LdIOsrFge7PtA
GBCXpvTA75xjDrAEhXrQijoP0aj1Qo6XvrnO1Dqto7ihbHS3haB0hjoI3FXyPjSK
ZQDXtx0MLcoCOSWYcQdZeuz+AKZlF+wypT/FV0teFkVOXQzzM6xkPcRKW2rS7b+M
P7HL+IRixpEVeg8LNPfDCLpB+/23bbiIjxboWz9wxV2+cP3kefSoKMy1eLtP02Al
+6WLo5EQttdM5T4/FyCxswQAJA6GtdkM4XttpZtKHm3YzbHiw+vZCw+gdvMHtWNv
Ke3b7fawpeu9gTVNeHdjhMNiJYHf4rD3KoT4GaUTN/hHdCqbn6EQSoRoEn5Ckh3j
4gtUrwRFbwlVqGzw8cmwZH2zhHSlephLXMYG2QU1W2WMqVjwSnY6cRRCBN/DSmOC
6+sb7X1x7EvCAHAWVlKKhWTmim8jTUJSyj1UZ3I8B03KB+4uI2AFT5EDsuqRQRz+
j6yhuala8/r9CE9LpevFVT2/DGCR+x52O3T3q8sK0lwL8GA8XrobL9IsJd9nz9Y1
MtTXJ57nZnZVTsLD4T0C0LPyFiw99QTNVRTsP76GxSjacwF1Bn5bewztsdHsOU9T
X1iPk8b64LqHE+mCYHU23np7nKLrOiqqfQRy4wmrWgC/vPf+mtkj8cBrtEA3IaOL
9lz4hietV6RW8AZ70Dnwm3HSwbDv54TgWC/o2+Qy6wr4Ys74HmtS2y4OCzibvs5B
WoWf95K/oJkpUqoKWW9XRyWmFW6UIAYl39ovYYcUHhzMyhH3+F4sJuxqjCWjpi9O
CGZvOAXiIhfpQ7aFVmhp4JdPLTuf0ffXWp+FdYvjRWjkADDD4Eqsib5C7qvYynfS
SOuMMHrPkrGEcYMxXW1x+URenyoBIPYb2ZZ16XhNC1cZhRJWDi0Wq9gpZb1Boop5
H1+W2U3ZBV3MtXE6MXzqJ/VoAph6HAJFwYaRiCfRazRFrxVIMR1raMqJargRonJ4
PmgmWiiGvlpiZgL3W++/mtSv3GPODiMMBFWH5QGgYc66QviRItV8ieecM0rg0kY5
IuYGcgdBfn3WSV5legPMnI/GZtNdjoTDHFzSDE4AT5sC6T6qgpfEi7QKZ59c4NCT
z5qlHzTAepH6Gn5AHOW0yRtIEvdGx8aAAGkS/S9kLlZs6lWZwONFw3kguEJ4M2Qr
4qvecgX4vFoqH3mhNb+bUuBSWCwMsBC0eR/HPuhc0QaUAYwpMd51OQxj76xXrxl4
gmi6oovmvoe1F5DJyYjdIY2AT/yHI7XHVvPRFOWfN5Bm0jeBN4rvDSTHMwTmjuBr
+ly9y/pGV3RsXPAGeUoE3dbdt/73tPZ7vcjM+b6aUBZE3AM8dYkFCEwn9XsovyFF
p1+WsTS9Iy5yQ/F6YlGsrJnJgkXRN63DhC6mjRJJc2n+XLaguN7IyCeIh75d7uXz
+o7MouaHTRfF+x7z6dukr0WZkZCI/1h0asXS6g+xjY5b6LrukH0Pn/nhUHhphQDa
gWxMaCcsQtnBpvQDn6KH0egy0gANbxV+yMGv01AuvjANUZkllgpDS2pcs1ybt8zt
2tbNhhwJGag1ecwIEWP6SUkI5LjBW2AQZHmPUzJ2VCFr1Yp04L1ZAH34bsIb3ZxP
Nv9MhWF5IsK/iEQfgBylb8DZkzQNZr8P3D49sdpbpNzbAgjB7UKQ/QiKX6hCDMy/
NSr2dmOGMdfG/ON52X+lL7juH2AwZWEDILnisENhlmKmyKpUGFx24OoN01R0ShLz
1XhtsTclmyORy3nCYJHYdP+Gi+U+nc/lTWoeHHT5CpN/hoG5bl9Kqa1X4opGir9u
hu0AxgIU72sJOK9jCJzipX/MRDTYd23shR7udWs8QISQ7kHduB70H4tBLV/j4L8r
/QxF2od0g+1awPUTMU/w2JoWPiMvs4NsRuMozjD0/Fx0DcsmlVbiM/I0kuu4m7ur
kKKa2SPQq0h66XolNFBBIjSSEsAN12LnXfjTuOdlH8Ff5NbWKOKadYHS1qrhcfoJ
HG19Uks+IOaQ/puVJ13Ti9vD7t9y+iQX39vAFa5c66y+QEpaX4lmEm+67l9vuWMZ
QL1B1/jgPBazPk+MB1w4LV/5Frks+uq85MHMhVreNt3IHP9ym0QviqE3ygRZuJdU
mxKiLPbF7kJCMVl140IVJ8cU43KXC8mFjIqEhFAbVYDfuNirqGz3DNcTikgu0xf3
A8CsoY96WvITQ/yNNzOJ5UKyN3kdBqoNag4JW4jFUgrxxT6nSDBRbDPBMiFE5GOU
ZLJVojYPMHJRX+x30UvYXNDQjqO1tOPLtYpDWn60LjC9yZpjqT3252AE0ARGWD4c
4xmly77pV45xYlT8D5513DqSlgmkSsp+qQ4lIVhqJ4aggeYJWYDNtfSHY9SuUP6g
KnUEIFyEg5SLIZIWY62bycCj876mx23FQ/eHRVdZDgEeCIaHJQ+xVgO5JR102Oqe
v95XuQEG2KG3ek+XzoLzbawmAi4lpAGe+qq44+2u515VPIqVFpCC2O+akxcc/XVn
s89+RPBvNJetqi65HgkutMIjYNsWs1p8fS7+Gtrz2v63Qi2WxIh+JQfdj0RZu4lX
hx460Ymbf4IHyRpNW0enPXGCtgD+pQ+EQQbc7ktIZZcAR4NEZGNMNorL3MkatBhz
+Rz8rTAVQnIRbXMvUxeus6BFb09jzM3znkRjkwdh9/ibjINwBq7ogE7feGrToCfL
TAgZm+DxmvQ0/+pgi2ibJphUqteeO8dg+/zxhHhv/SyDEQtNk5rA9G8q+F+z1Ke3
uZZi3Ifyzt1uXSZayUr+Mw0plQqIUbksTKU/wwRYIct34diIHujF1hehnAgi2zlx
TheZOVssstFe9tqoMpHaEI8oJTgKmiPQKXkLR+k13FfgtSW4Fcp706uVQzb7sLsI
igJdXKM1IQ1OtIxBe1Or3UeHZKhlg6nN4E37oVYJBa2At8tlWmXs2K3Jyiwn34U0
fukVYolXwnwQbdYcKzAzMhn0TuXmSKmpbmAc2R6j42hMvfNEJhVWyb1lCP5am5xM
5RNNwlM1+BFCFskOTLp4EAXPOKCGp7C+jTCMiFMGgFvFTErlFIY9ufkEkmeHcppU
GN6XGne8DfuzrhV/Rk6VSj6qiqjMP+FwS7RnF1Hr75i1JlBLAx6CGNEZFO6B9i9x
crCzXVbYAHH+wcB8M8CX1B2eSnnAnwkyC6lRu+6vJrXy6g/cS8JXNCkAbjTaGymt
+yhygQdUepjmVXWIiCmLNFDpflivpnnr4KN5PseCYJLA+U4VCjNo65kcYc8afK+c
Wf4hlNUZGVy/9z82YDHnBHZZ7rnll4pTgO0WmFlZdg+ZrHGMp8E2GlP/OvthZk+Q
AOrVRo6czMFMsK/YgA1oyRlS6ZIx28+j/6LNAkkbqxBGUIbRjr+4uSbtDvNRCNDo
4oBFDc4XO2mnjo5MStM9kzYr1EFKFSm7aZ4LT+rfxULUN9E3Y0N5+5bYloqoybx1
zyV4PjdqYYggWzLzJP5n/ATXEKRXyLONKD/1ZgeuXMQ/Fgvpi/sREX1qCbKcP3Ge
6r1UIxEGRDsxrHdjnhiHulZ911K9tjWZTYJxPKRSjQV2V/nkzfwfpCbbfLh7/DpS
9ZP/znRo3+2cOb39MmYLHAZ3V79JcGq5dqfXrdNvZEPRcHlvmc6gmQKtBBU8z3XU
OlXp4JifXqgQqWw4wIEpjLSGmXDEUBMEkz+y6r1XKjsWeiV2Gs3akK3EgUZjH/pt
bHMBv4gK90zAH4dzr1cZDZdfAtzgOn2h04RwQXNALwfEFLVeOForx7yLVIS8SdCD
plsTnaiRSy37fD11ma0TdPjrgRsZwkPPHEBwal/CmTOE/MS53MnpjjnBfMaLH/pu
Pl+VnKhoXBvORjaDz31WhrsNZFv86tXhRyoKLkoezQdx9MvoJkSQFbz+9nhrAxX3
YY03/1MROCwnrXkurxnh8RbMii5B4VRW50QJyHpNl5fe5oPWvWTf1fQ9zGV3++cr
clgPlzNhZmoDDx2PldZLtcpv2/Vqd0RucQUwRHVcMDEznEuOHODGwidUFCvT1Y/n
m0t6ajJIGevty5r96jKixcs2cLuo3HRukLJmJM9OQYgfpwFzwPMw+J8cBe4RUW9t
YXoLr3y7SJH+nWaERt14EVenognnAH3nbPtnAnBuqyGjHqzoS7zQzvkRyYfl9VNv
ItkLh6PXkep840B148FRAPGv5pliwcMnzNnUcwIZKCRz8jQl+MQHXKkUt1XkGCjG
rd7aW8XmwLCDoQe/lN3wAzpcDFx8g33b13k7HuQGVscJdw+k9TyBnUNCcP1C+iuK
qlJaAN3GIcwzfI6iNSu30tKuMzNQWmljOoHzeqkYBKdTSlUOmnGHaHPUzllDBylR
iq1eCgk+0lud0h358bLrZTBHqafWXWip/OlNd217n+S0kTf8FoBQP2/XMKH1NR9M
Y5RrsNersI7FJraNLpKQ+K8BxzUiwYPfqa7vyyiypwuOGKeVqHV/v/vZeJb63N8c
wkfK09DOT1yRQ0w+6lSmiOOmtaMK8jLuwv+7as7ThHkAn9PXLl1VjfRmCm0WrAst
QdS9RGyNNKLMbVXqB6z1MxqywdKyGP1V96bvpA1oyGCpeC/bSYqZz72kyRs59cPt
+6X0EMsp5bRAsNBcOf3SeJsgv744alBRtf5xtTLAMp9hLPvnlvjcRRD+DzQuGQwM
GvrjL7zjNHpSmrsK/km/sctnT0AFiehs86MT/8JrzAbH6ktHa2CzpIyZuv8dM41u
3JTmoWypMvh3lhduKDBNlXbrwx9IjySOVS6t9dyuA4YzNL3iJrkF/bBde8KbOwzF
hRwzSsVLTsSiuu2kLiGUKDmFS4Dn9tJPl6FSnWtZjeNOTJGE3B3u6KCyRejvQL5h
DI/hnNS7wMB6YKvjiMEPThA5H54aGRiD5+4ja2QP7qDAt66bClG+cSULDJlGC3VS
ExGWmuamKD8XbJ84/L4xRV1xfSNZMCCA8bpmRGVDnBQmFWaMTe8A9sda/sukEuHq
hvUu8WRXf9hz1iGuWd43hF0CA3pgmZ35QC2ODPWhgVCSDk+/vwreMxi15HxUY7QM
/TDABh7aPOZI7GuyiiE6WgLFVqGAyHEs7R58mANxdHngAig8yKHGC+gEJI7oTU35
zBsTQE2RBMTZe2FiSxAC26Q+035htaYAJsR36VWtmzN4A+tu44o1m732bwK6R+RR
K2HvKnmqYajKe3yyjWXl/gfbXzQi5GP7DpM1voyE12YruD3neK4LATIDFZCiQ2r8
z+DqQsMj8LmgUzEcwLE4bIedJ3slQDe/rIqU5uJ2pG5lYIxE682PniikSHF7JOYU
eFepSRp2IcUcBMG4CiZyHsHyqqUzcSgxW8ID3MPHy5lmygJaQjxJ7ymwVOhH7qdS
Wl4RD3czwY9tPcciOcQBfe44/psm52r3W/rA8caUWoDuRReGLvvBLn6p1B9M8Iv2
Tp1jtx0w3ponaHp5UK79/C1Ud8V7iQC86ya04Kq59jCUe+a3Jo99xQ6qFjeosimb
Jkd5n07e2yuBxuCDQ7op5qs/634QY2OyLxILbd6abXb2yd0KyDEFWzyi9T3W+5nO
Fs9+YiXkTkFGazRr+rHC5/lXfyJvzALnipFKMh3RTK17R55sO3us1x7XaqvzF2r5
PBPYl0ScmaLY0+wMcUQoTBHEIoqKclf3JVfBEyJQUEVyY9OhdDW+XgLWejkTyV8v
TOK/OZpnCt0FfwCkYwjZ5h7yCa9fiFCUG6nC4WSfmUAuVVKb8r2D8EQ6U8pHzefm
Dvf/m8vl+upCMgGOgyamjHMEQepDtEho9qUVEybVcx9Tn4Mc/AvonCiB+IQ5GO1V
X8bRwDLBLXwa/EbaNwdOOWnphSz3pb1jt1bRtS1CqIzLpAEVPFAu2LDtLvWw08Uu
3PAWc2LIUu24dh8bgcyd6BHrYMfa9bThbVzto+1zsR9OrKIJ3AMfdQ9Qg6YYOVgb
M4jl9iKj65cXeAGgG7ONOc4QYhcrp/3YZS+N6xLOLXTU942SGktLCWrM6O25dYBL
AcqMwA5TtkhVTZYpYPFV1lKzgDhPFGsE++fuF5t0LdX3Io/FIo7ly/8TKWP6zjpJ
fc+BDSoG0yOWtJFm6afN7qO27UMudGMgJsxvfbHkGcNHm8mo/2uuo7I5braVAowP
l9E0P80lW+ymnj14V0N1j21vInBqvNGZayOt192FjKacrx0W9pbFK6NxKdOQAtJv
WITKJqhwOCY1iNwC3QtZXhyqEkJFAdaB+6nByzjFgY/HXLCw6T9SkFsCQbd++n1a
AznJi6NnUmwGcV1t648VMxhaK8Qe1pakbWLFz+1H51/lkHjMMr2Z4A+HMnM8lZvi
JBz3nF6xkPuXTUPBqoLPKqXVO3HJatK5/OoL8UsgO9QHixJLY1waUUXml4THET87
B1gWoZ0IfhIYM6qjKqS8jS0ceRLwI9lXTj0+J/2QvYXXAZrrcgC0uiYgPGuzwbID
ZHdWkp4hFTn+kmrJmBa8Y10itH4Bsyw00a9g4lXewEJ/2cN5GlNOQavU8IfM0SLX
LvJiHzFjwTzfhXAT+ZBUg2pFfsl8T7fWmc41jDabTt57BqI8czXf34zICptaJerl
g/9o5vNBwWhVjpzvNZLcCFed1awhVswj9/9WXGRzI19fgw3WXIuZM+E5P4hfRgKZ
ZNWf2Kzu6J9n1jPhKx/RcSU48GQER4NKX5TN5tvW3QlkQw4P0fKDHw5YBh34TCg5
q3rSrXDysJswsJ0JUvTuEqByjTR+09J2hDKKCeoAsC+zWA5MdUYnMrqpCd9Fj5Lj
t9xcvCooqwmm1IV/ir1tln42399XZ/bbrJ41K5Z6P5Xj4Egofrnv7MFuyPxmPH8/
g5BzWYENgAoyyH1yvkWQq4L9BAbk+O/e4WwzkpdZPorbiNKNZFynz6F58HculC+m
r7h85oDwvAqj2YMM8dyzKZD7mg06f3cQwnfe5QXFsT2sgJg/3GpXL0xQQXV7lREP
ZRWavxYVH74KDrCxqCouf4J4DRNswPBcMMMBC5CDYKQiaMx6ASo7c1V5ffHzitIi
TGUKmBTldzAx0GgmQtHETytdC454Zzu+F37OUDGk0VlvYj8h4A+4o4RP1RNFoHb2
5FtBIn7FCwtgPAwi0m56Ed+cZgJBgMebV6E/kiDUk20t2r/4UHcoOMCUC6UhtGo7
vj31UKbuyC596f3kYv4CRavaAB6M1Z9F+9NhDIHretVl9fGIHamzAXMp8NkeYIN7
PTpzN/Yx9ileczkyrDP5oUcaH+yD/C/xcOfHsHSUrIv9fiNi139RUwi9kk0EtK/e
ugFRi2MR1HQSD7jzlBhdUTE2sG7P3oiaN9SDFaZb8CgxPA3o72tKFgER9bUhMme1
rR7LOzUuwcZMZIHCKzURfQJntmCnurA0eH2n9ry9Ci7zVw009qIytoZNjoXVBoBT
vcm8y4xkGQkal5IfLyfPRhUqb/Ib+R1VIf9Ut38M04OMMi3wSB8PQsd1lLEDKY82
Q0o1+filsyyvFxUYHpgIXu9Z8KKEoJObMZEtMQ1mOjHkSxCm2FQLw3ITYoKHVn+Q
rUXmm4piDP0Eajz98ipAY315gjyr0YKqKcwZv/tqd2EeTg8IYVBVByicHaapjT9a
0AYUJkSYWeY3rcrKnsjh4Rk25z3DqXCigTLzyu9FwHlVJwWJBBCkMb9kJG2hZdNG
OxbkcIMvzqQsf3Kri2x1mXdQksrya1xtr4Q7OBchCJyE7VNDcEj25tCiefWb++Ae
oHncDbeFRBwd+8lH5oE7DoAgUyff0lWCGSY/21riPkqpdpIiNswgVOJQQ6scnUAq
8tJr88xmZ9hA/tuKHgT4skDBXLdXlOK4TG+/h5ks3kQfrwdMa0N1FnJLKYTrVF8v
EJK97tBk8mG1OSPxR+4cPNfkeDJ5VVQV6UIreQWr5YpyaxC5WgvDtWegrls2veXq
lgbcmu7qpKxJv8fGzivAdjhAD9on2Y/qGk8TBVOZ+i1lwe1RLDsXrPKF/Gw02n6r
kYzCeLGaJ7lL4RCx3ESFBK4ekVeFnvcQgiJ75y7+DcF/j2P9K1MY+mKkkSbzXxVi
wWIA94pUhrluB/L9CfmUeqA/KzmuQCxvbXbbiv3cECaYVYaGKobM2LLRsk1ofphi
VFU6/t5+msLJBf8zQ+M0525ZRjqKGZJ+GBaqWKBFXj783yfXMgwOj7g8tqL0KJ0u
o3d9TnVbg/jlLiBJZ8KQEZom9VKUO5b6unKPLaziW19TsXBg7NwknuEiVnkgcYK2
OzgWV1sBlFZBkSqi9cfwBzsSPqa4lghKMDnQZ5JuTOJ+HgvOO5PkNEx4UbI9gWd1
fm4rnnXyyVutT6BE3W4sEElD0yhLOneAA9dqfocgUxsYWcX81Yc8MWry0b728s9M
FgdbIRE6bEVCvVYSV6kExM19UuZu2jAmJAOYr8LXF4QvmE76S0gUcmunX5CMaiMG
4W72xAjLsHRfkXYRPS9Gor5YfwTNpr1pQwl84G9S3U/0fZ3bGofV/qo41eXFfQYU
kn8cNKubCJAs3VJSLUYmm0Okz55HcfAYwZ0Gbpt/wvUYZT0eiMPnJuLK3Kz1YmDK
n7e499mrtSXnr4ufW0V2lc3IK1eHaf1HxRGL5KvljBMX6vkhRrwHd5/ItO76Qdr1
kS02kj1M1GScY9A48zm4SmH9MpQPg6Mmn4pvljt+wzTwFTfUg4AJ41bplZEpsFIX
5PS+rxl+ZGVhFBq+3XX0a/pXqwEXFy1IbXdmhfqnNv1mZE+sllrx/s1dHNtYgLub
rCcXbv8gDM+Ck7dV/0JDfW/koUVWpvJn3b+kUgSrq7Bst/+QTxj3XUpzYMl98Q4A
Q1mZogt3FLFyDvTy+L21y6EvU4lpd2wqYaGVF1kLWVu4QVtbGc88DWckDAKW4aTF
FKuJWAY0t4J/o49kMbgR6rnVIRth8edG4CfaIVpS5KRRX3I1gCgHmQGu/ZZgY6WA
zT0YVogggb8fvq4hRrsmmWCkDxYJSgX+B/mow/FPCaFG0DX1UdK93mgxVmFye2la
6qyGoJdFKc7JLLx9Q2FWumbpGUPDvSRJVRjeS15ziUau22XFyd6T/yL2+qbtViS2
n0Aku6U0GFpmuHGpJ0uTAa9AyB5wpDANP6+OP5yP/c9Yx6R7eEfmCC0Pg1umtVeW
fDChjkPfCZp0MjIzjXnUlKuQXm/3fOaM1sLJVBiuogyWnnqCZGhW9Qsi9Dc9g9XN
TWdcbsXImZ74edvx4VkiqZ0PVDWzLf2URYfuz4ydcXAGokapWctRH/U1PklVGJHY
o8JN1ooI1kidfK9nRdou8bINFOqyCgtmWKzGpTGGRd8Dsww3s6ZhXxxobRRuO152
Bs1/yjd1WVgV9ffpKcvgi0+x/voz6ilPjdBaAOc1t+dzGQpaHk5pOEZaE3wltdDG
gZacv7RBJmMgcLI/Cti4H9rlODTg1dqrClkTxcpWuiTMozENilbdapurqm1SS4We
1NFec1blCzciWAUVZb3YXDNfQ1FuzThrMAQ/NzALu5rgCnnt/Iswr6a9XONqi620
wwK4LexCDqN17SPYfxkrd3KsYhXpgMnyD3aWBNFi2NFnfnOHXUlAF8LwB0TKA07n
5mC0SGkrPeMBBgHdkHw9RLohoU7a4e+GHLyOL/BQdXqHAJubfeBUsT2RdZ/5sFAP
L2AAwWVSunlapUruuPSNQd0sTpRWXJJTjxSsuygw15gEwxBZpuFToK41AOWazZcm
JkLO2rDiEv8ncCk9MKIsp/MWRXfQwYLbbiHB6R5f7EBDWFhNXBrTvxXUy/bP6B9j
C9v1pg4gA0iuVgc8y2AQOgVsIaV2hrAaUzTeNfkvXylszG5sZWfmTFeW1EvrU5xd
KNtNFDCAxP7pnqWcHayPkI1vpfdjXGN/C7S9ANjmjpuFd6GYjDx9BSIKH7Fy5Idg
oqAhmsoxEPZ7w+UFblqqvZ+NfpraO9qwjKP4MdNQaZFRsUi8xv6FDPWmgETT8Ina
NJ+KL+Zs+Jwevb1eGDiofcMMHsNy4OgQmEub1d1rpjFxvf9d5uFO/g6Xm2AwMKQ2
xRH80Uw4f+qqd1Nhzv5zsFcHigBDfH7JDoPhdf6Y5jABupoF8cSYTmRtoMOVFkCG
7zGMbQ7M+rYCWpQKp4TbII/HOG7P7kMG/A1jws2ul+zEpIAhoA2W+TCjqKXvp9G3
PCiRUFsqUQeQ9gmOzA6Wy4QGiE78luN8e8PT/WPF9L8hxe7QLcPT1lTDK5r0EkST
fLD9IfnjzrznNh1/K3bPH68M/0uchAUWH7W7Lg0iCaGoTFLX07o1QLvB7oXfb6jm
e6qOj2AvwcUvILCWROvcWgx1ful1fP+ulaMG0vERAYL886/lONKgrs/1x3FEobCS
TMrHZcne/AqNjT4riw580ojFN79vlitBsTting0OLW/QQsZRcnjG19CbMTEIPAYg
ZPOsXNhBrCHWTer8h0diXSqscUUv/A5zFI3+1trJZ+g7KmMXbllkqxtw5BOeIPzK
WVW4Im87fzACZRDrETeloMh+TaOrzixO6cLW7abYnDJC6S9FNORCzJAgX+6EXC5R
kw1zlD7cGqxbQeg0kG618AFfOV11GLIkn5QEykYCx5MObYIx0/It9htrrkd3ThJQ
IKgu/HkYzBTTnHTlz4osglg+FMMOvKjeF+QWsWDkkEKVHE8lyPBPpJuWoQ5RyfqD
ic4WSMz4Uvj2o8+rv5gFq7PRh0FjJQqVcvh9fHbk3wpvcUIdxy+dOfHVxPGNGulP
5FVyGEKqtyB3fm4Yih/NJrfC2QrR40S7lrUo4kAqO3eI3fIrMJUOHf8xMleSCaQp
SnsQlU0CWUeCQlUyVAKBn+2aGxha5lGK9pS6NXvhsHp5KFCdJ/QJK3Yms3oRP3vF
DYy7DUEbQTOIOMDeHmOJVvYFKToyp8TTfTuV4qu0XlW9riyoAVXSw8pAZb5Achfn
C0QpnHjUemslZf3u0cMAqdkfLNf89CwF8yp44QKtWKnTf/SR8dq0OFvHzjz4UM+8
7pQqHHzZOpf4BBZHZCP/G9M+zcvb71EzpeQpUEOYo92Ems8op0RCWFSDCzZJBags
589nBSpU8ay1zm8b8AT0IBJxWr02qtt4XE6pvZOl9Wb20eMGRgwVgC10Hb/GbYCC
PMkD1CD5Bnve5wJdvDzQonx2UOqFOxXiHFFLiN5fdx6V+6VGb36GvW8ls+vJrYCU
gE8tsAza9WMWDgJOnTXlViyecuXnN1+bFNvnsedoVVCJz3tRmFS1E5oZadrVHSTO
snN9qQtzyPqdJF2h0kLRrKfbKRg9HasYahGrF0XcJl8BQE5x4NuZVSXDnva/GfKS
NrYheRFcfyZimd+F2fihtcMvh4q5HNENZnPAo9ipFhcCq79QVBdmTQ7CuVcORDq1
zHZ7iIoCspGnTg1r6OyP7w3LfSdjkQedL9B0lPUNTpn+zsJLuD1QIXBQVqyY+OJF
dCYtsGF/ECXPxVHWJP05fR/S7Ib49lyNJ0HFiDqzNeDJ3NHLxVgXhfztuKgBR62V
gP0DxeALPP3lPPckF+IwHF5gyGCQ9TDPr3Tptg/gDDISzawWDV0oeX110XPxaMPp
firRHKZspjtBYrFbUDsMvARddi3WcC3J45LUzYN/UNI4LpG2Camu6p2Wwq5eK6zr
WTQj4mB3zqanEHVeJuZuel0/UUad27puODVZXy5aEpyjwE7fTGacZZbBVc11yx2q
bAJ9xtYHRGtboWLDNPRLYvv9QJA7f7qzjHo+1NaAQpRujfSC/OQhkrmMxTrObbNZ
dWkBtIx+Je8ZwSvbPtbpnFPKbj8P6jrTI3MCZsETE80WRO/XZrUCt714ZhUQV4zB
U35Fam/QraKg7BzvFL6glecazAgGfxyiJ6st03bn89rob8eTlM2XsVqsFKM/xrsq
aXOA1YU9wIWEseqVZQ2poO/EuVG6+VpjuAVItTKZ/y7AGv23U22lbEZDfw9PLvsE
sCUv/1dL+iof+OvsZfjlREs7tRKXW6FmW8FYgH6zKRGOlZfS3LNS+6PkfKgFiHXO
uCjS1XWTgEPkconoH8c48PA5JcwqQm/Pkn643h6c2E3aSvj8GsvxKttdzU7E6HSK
5PXJBClDe8DhDDI1Z8uWdSTQMcnnhKtZbx53s7FTHuzlmrMRtGPwQLPj6zAe1PE3
lYUOpNwh+/Y0kOF3B3rmYfL6niJWWqJThdiFEB2SoPuqf6LrLA2fTd9sJis1Auv2
oIz0Jtmr0hK9G36UiC8GhHJW/FeZ//3aP86xmjSV2sDWmiL9PDJ+lT+mIp/fMKju
841Co9zNdrvVuc9aROTkSiTYiQQYbJUtbT4+jFtes6d9G0tkrD7/fpyTHuFKkpzd
qt6VX1yued7USc4aO2s4PjNfbFDfkR8tCimOLI/HO1NbjgxJ4slWeFlyxj+6u45S
gHcfr9gzklUFklB30yeieWyLfRiB5cZ2roHYICIPG9EI8aFEqd2yWZB5J16vzqj9
XPCgWg1AU8fL7exE11mx5vznkCMzrVklCGrUV5bnlFKAzIz8Xx74Co9+q23YLnsz
LxtXxsZfavNkEGV3fkt86+2rWiW+M6OjE1rVNXTGDjdwlN8+NO7/zcuo4lIEEYAF
2C0+kECEqclgvPHumm8BdGQkQ0hsR98tbkDpJUCI4NxQ3MS71brz5P2L9uWRICGG
/9JpYCkcD4PNlik8pMAGvoc2t9QrwGQT9lugf3lDSj0WFZVO4pIxMJZUPWu1U2mf
pLSKsSVAdfpsGY6zsua36WPrb5hygiiKilg/U7ksKJwg2/96iqaTSd7e0WCmSfVQ
wKmy85dzCDa4TlEv9ArHuENiNguar2ZaR8zvku3xoyxY6y5fiUFxFP7xCMc/Evdi
IXrm8LhZ2NdPtN74N1gx3RXHCndqjO2ydTV/tyR/URhUx/fyEUYM/S6xA5IXTHe+
iiWrtH9N2xM9qHLaU/4LzefqE5XcAIVoHOpQTUL0md/CyWnbmnnuoQ94oz+zJFbX
RKfFP8+kHEG3A3FuMg6E7cs/PH53eQhZ3xvUABYnvBBpFq480WYyAOavX9Aeaub9
z1VwTjAtoUWD25cJPsVtEwVOoxsIKXRFhYV+sojUZkAZyAvQCAaM8QztfyBOdRfm
uAxr4l4K3F/n7Eg+sUJjLb4Yh9q3xNtafU1Os3oEzHcWEbK2Ac/2gfv1zt/CfYmX
RqbIdpsRzTUvuABpRYaxmohsHQSiTnMHZXpUjZaHd/kgLq4qYrM3UpuANTua6zdu
h02cCn1UI0Hh4jStNZg33cqczXMnHHpbIL7O9ig/6iqWQRSA5+QRndDQFUzc4Qs/
jljNFCgQ5cUpYL9wk/4nkjZfnDPJMvEGQHbV46yg/Metj1ymBQUuvNczieHvt9c4
63Iqydfu5r5WIDGu4cFq0jG6/2XxROJO7YMNaYzlhhUDN/jc11Y0M79CE6p8FIZU
zW3o6ymDKAXOXU09ARmxL2SJYrpO0AtvDQ6x1PlQibnqFrBaDohptPaqPpjQHd4c
8veLwPHLAdWMCcqIylpvv30bW1dCXIB6FgHRHXrojkITbCqQFK1d9f1ssSgMVH3K
Kcz3HPLOAFNNMnh3ktlEUrnu7Egl8ssy0kYoe6CW2eLfH5AFbbHjJG8WQQyPXGIM
1kjbq0kmyq219bIGaqlu2sqKmj6p1vPlnAYTnnrGtSTYzuUPK7btUFreaYOFRI06
jLJQHPoTjyrwH5LU2EFHO1WSyV9f/Yfw7LInQEwk0nGXtHoA3tdqMtDPYHygHdzj
ypB8jekb6p9m4jTNUH8VRCwwMTwGX2XL0UsmzJ1055IvPd052KTz5j3W+RaRTZDD
gyxTHcLcJPL5wkf7TnW/ByroriMJmteyg7ngF1XtiGMM0sIHmGD6muY+Ugx52qxb
DyYXsliAap/MyDICEIfNEfpNUCSIqF21zqNZ2QunKvfPiNogw9G0lfiCqdRSnHOL
qqaV0ZRB4qFPQP3M7s9XdnZACwCyPUacGzBl9QpOMDg9+gMv51p9GV/6ZmCa/w2T
yANF2mJzUBpZEwEjmcIrRFMkVno5NG+RGV85rlv2wqkEYrjpTyBgs4gxUBvB9RzX
LogxPUm99GCHOYpovVG9L5L+u/t7/ou2//bqdMUFt8k2hqkj60ycGsdp8Xj6Sgq3
XzqPcOeLxyFwnCkL3vJK7e4UU0EpNQXuqYMo8+uX5DBwLykDhI/zVgMM4Dknc4YY
9bSrhLCiiwKybAzUApmmvMxJkv/k13bjziDIJTwdRAs0TAm9sPHsG9EXMYMirvw5
PN+kiJKZSq4jxbDYAGWfR36oj+nZG9+uUtzztM7Vr/eIYgWZ9E2RUSMbHGT0iCWm
D7RVRaH7h1doH2vBxK/Z0LOxKmQ5ObQueB46UbcLH5lFHQyZLMoMkeYOexY/ZB51
bxNw4fLjeLoMCdc1G1AfOcr4Y0OQqSuyo13FlwpUb5/pqFnb445uy9yRAYYkJVAu
egIc/7V+lFtVa3SN6/zLxh7+SvHOM61TLRc368FXKcq0huF90QH4LcYeMeXttPF1
gDpeweSUEsUns3Vn2/tRGhhU+Sma8hM7hO/XS6rdaORBxB2NKNv9eR2yf6gyJofy
f3OToypDhkqR0B3MXUkflFqIyUTt2zDd3jwiIPRxGzjtJcTneSctO3liWmyBjt/T
An3/W+wfRSuSiwWfUAwLjpSqX8fj5kHzQOkdMsp7U89B/7sETZMLIxdtQK5qfMDm
5Ab/G7ZiO5edmwUVRzirgX8SiPsLu1xpmrsu4h6F6TSrmB32WfuWLYJyAO1jR6hz
SCHf+yA25cDS22NwTnMI7t3QQVfbtoC1ISeaVmg97ld5fbTejHjztaTLhd4/WpHV
gAcggolFDyzYkt5pbWj1TBOxb3TMKSfqBGXjPlZVJcEpnYK/f9Z6akWdiUp2g521
dxTdl0WOORE4TvoikhintBTPnnN5/d+47wdByfbfZr2EHo+Xd8xnJ/t5KSpdhtzK
qn5JzWA+8FLQ07moI7n0H1nNKNDEeo4uGZ9cKcWMVYkDpFfTZ2rPQv9bOJXd1LU3
LEt2soBpITMy5RmQ35iuvpKyteFQYn/kYz+riQa3+KGA3W4l1EJcv/JvsOL5Kd0S
yE33LhUFqY87I9GQYKsjA6g4w/uw4pYbB8UMFrMUj98nQDJzcEYrjqb+/O6fL+zz
VHxQzkS4ro4jr/KzYeGkAn2tFTkw3ulXEekVaKc9iqQylNkVyPEmdyLvjcYgFKnk
q4W16QaUbDzzFJxsi3CILPV6TtBgrMf3ULJ9jqwD8UdyzMYHOdV6Psn9HrGaPZEn
A4lcCQ5HpIA+o7g4N5woP/NF2tu48x+bGr2/hz3a/8kMtNb7hLXUtEWCD2J8JQnn
1MFWN039TvWuKtOufDaOEKpqaw2zI+ZxfRerY6MPFYQCgmJFxoEG2upvKNgOn7pK
L1Q9XKJlXu52ziy9oGksfvwmXbYzjZ3XdnIqaTInTCiEzmSqOaVNeHFQrHaI6yT+
1rVq2M7oABjXwjaZC7mbORxV4ghsqFZci6IewtHhzwCb8znWIIfrA4VG8EZGhcYZ
xWeDhKB4dCKmZGN8MdbuT85K9ExotIg0zRpFOTX/sQzayRioqIAtHOCJqOMGJuhL
9GRQSVc+OllxBBfDxa9AJ5+kyQRIHSM9r6Ph3tN9HXmH/t+gTAlZG0xCYSEHg3nM
l2NernHWMTMQUpILJcgpAh6CsYIBIcliBhzyx8NDmVARflrAcRXXXNW685Bdag1N
xFyg0DBHp+PaRlYiDC54G86H9LpNWeRptD3wVIki8CltflbKJN8DWTk/gDhnA27l
71auySE3KbNpyV2Ht10xTFBL2FfCzzF3fjrhmmVIzh5wVDSAtIY/e+bL26Oj9cz8
u2V73FN/+PE2/NLs3alAAcSWCBwyn+nlcodzVaYZtPWCOlzY6FPjTYMWRumES1eV
J/ThCB0mysNFjiuJqK24w1WgSTVvU8b4jqgHFpSazgRLKzawQxTdkSN9SeCRTWGX
taPBlEXkJpd6LcbG4LXdxdYFsnq+uUtsLmLw/tNY2ncyd1IVdyYl7ErwlEzJd+Ri
ZUnpSUS8uIldLr/ZyAqyjoqYc7FkAQFhguVgPQl6NcHHACsf4SOEVWisU4yBnwIJ
hRKy5rc00qNMsZ9ggIG6Tnjo1ojwMmP6aP2ustjfBi1qhqiDLMwSrFxgoaRvR+jm
mr6qMfbyaztmOZysZQq/zkx7V+2UGrI/uT3gpsXcyceCDgRSJQEbWtQ8R/P5lTKC
7F+bAbA7dHXGCT5MpzYd9ILxgQcVOvivXwzSPY0X4IXirstL4jquHZi7E6/PAZ7N
TX7pid/7eu1M51Y8dkEGX6SUoUjTghBxJjeuJ0SrE1uSRF6OfZygYZiTCXtZRA/N
rNguhDsUX2DFtG41nCXPm/fYOss3fP4DQ/DhHRq3QZjRMeXcfyNoz7lM/760Jrsb
/mRD1xw+C6S9D9QZRCOPPfQXjsSf+6JZL6j8AqJiLvyEZyoqv/Rat3V+1DK9d3kN
20rMUeu4nU9s0fM6sJuVyHmkMCw43SX3VKafyX+tdtc46Iamo1HmM/9RRjfF5miS
A3h/lK7HoTiv4dO69JSS19xIOBQqO3bx2xyvIMZ+uPPozuMQYUcfYnvHh0iGFchz
Ujai0CYat8OF6vV/S/lztMOgYb5JjmB8q5RA2Jlqqn0wkWIXQ8bFMiivu7X7d90G
axo+5rQ3+IpXVHv75be4ZfLOh6fn8bGG/LnHIAOq9rShlRn+KG7aaMORnH/FuBR3
sJ15Y/6WesOw8UTywBV9zoQ5SQhs5M+cAKQHjXEf8gC+MWuvc7BOvVo+nPk6t5DN
znc8V8s8HOf8XjmLzUw1ym6DCfsUftEdJhS7UmjKYgGv7fHMHOBlZ19HFydFb5Rs
aSaVQTCpGfzSTM1zGYYQ48m0icOcHAx7yPkPK9hc7X+W7cPrb3G31w7c6+n9ehMQ
qkx0Rjf9o50HBRafJj+OoVUGeQLxGPcLN3uGVR2XhWwYHH3W6KGuvVBaeoZLq1Wj
MqHi71pTIYUyciy8Zwz+1a0wPOmjEagRA/DftYf89W7Pyjbh1uevTW6aOkLFSC2o
OtVMUMEAidSvbWIxTGIB9cNjeMr1x44AzFh0n02l/KApPbDvtH7KMpMIybd0+mOS
+tD15pxZwMkgxcVWFNRqrG9VnVBtG/KtBrQN7xc4LEWeR+pO4ksgSAAEVx4p3PNB
J5Bd+e7RkyYiluT03EIDCYjXP/zoFe7Njk4qSjNHkQw44e7w6Pv7+EWN9gRFNgGt
wQY0Y4meUUJp9vaHE+fFDFLr9ji67vzGlO7qEdPTDPb3hjgok+kBA14vigKj7jZ7
mu1L5NaiyRiDc89B5f3UD5buasYadb6wxH0kKrDyZaHig75YP+qGCJ6oMiXUAw2M
MDaorJTfzK69Ufz/nzn7Hma5eWTCfkKsN8NGc9Z8ReEPmhOPZISWUhaormNNE711
pyxzqmtIqUthb6e8bmLJ1wwf7TbrDC66Uo3ndJ+Q0Oz/0XpJy6bed3RqVzrH9bkI
W9AnCg7GN0HxnlRJHeIW7RzFrBI8Ec0Er800Ev+vL3mm2ANLLhf3c2LLIbUdClR5
Y4u0SQObILNQK/DNuRZewF40E4aSuNKaSBF4mzQxOTQBKvsj3l4h4ULOdbKbzgv5
9cFNuHtjSv9Mv2eAnUGjkVLzbTfZZHx5xMhJQQmqq8JMKrV7q38VDVJA3rJH/cVY
yDD/cDgAnPctCIcFcjDhgEvbWHmhYHhwRQgc/9LVR7tw9rA2R4/HEPuZhJIqVzPe
lOEj4KTQegpBUTqfLLYzqGkW5JU4vQycNq/lt/qFXEb/E1t6AqEXWcQXsyMLSPnp
lMGOFml6eB32gL5fsW6oMeH+Cun4Xg+SQmHcbwTvMiylngdVqXy0EBFxRVibgAJQ
TvUR+Tl7ceHpHD1r17gu1miRMa3fEHhPGsTN3YWeT/2Ox2wm3CEZVpNvUxaELvRM
uo95psxTXociWmktVOQnhmnPJ0v7WF5Bd2+cEI6uDxCpWE8q9oXW9IKNgJn6GKZ6
+syrXFReYp7MbsxO1vTZzDSCDUxPpCfKfyuV40QJdZ20wLR/vOQM1EsjfoKBuURX
CagYqk6RnJVUOvP/2V/e+81NJMqSjW3QEdvQgTTyVeMgAXkwsnq97T1I8CCKJ+aG
+gEOEvLan9V70ZKHGOZ/U0YQy7/52Am5iDVBn/3a1Ic8KholZju+/G6c0e2KGfvp
b1wOMLzqG5RPnc15E9C6zfqASlr3zLzh7vdY+Domu1jpLU8c6T1hbCXyKOpepKN8
cyoxBUh5LKAQmeJqm/sCtl19kc4JfqnljBSWggYFFHOVWqG7lHKAhpPjpJtvcjZb
MDZCHDtsaTpJJ3Ht0bI2F/YR3VK7lbKSKqUpupY0v3ZSaG3a2+YyhYRf6rG4gUjb
IU2eFFlI+PSqMby9HCI55LEwvrdWbVHtrEY05gUe+fyrAeWzThOw2mJARyqds8UE
iniyffELuR3dRtMndm2/cBNm2CBWKIk24uCPVzQAYAa9cDgQ/Uy/zdcwXSnSHiCR
ixnff1Q8Xl0PuvMs+QfKeQJA7BJ7isj2DIKp1ki7fmDcH5PsKBTuZanXyHDbetnt
Fcv143QZJQS084xjRpL7+ThUCxtzT74cVTTFUoo+ZnxE+Ps1wIbNM0qXhqn0m1sh
rqzYR5gW908x1FWymbcU9Pe9KVCoHYbX73jLKBp8AS1pQV9kkaCseaVeOPnSJ576
drdARcE1BE9Z7WMFStG3ml6h1YwIYUTurXTjfL/fyIQPvKoVhsnB+XfbSE8BW2lK
uG9tT802GPk3DrcpBi1JxCOn92n2ama53Kb4wmYLg7eK22ApUsiG7ZLvSty3ztLk
L24VSrBKm+8qjAocdbs2vueJO5ORqUpExnAjJeJn71e/EPD8I1Doz1kJBBLhKgoU
toYoVmcWdUtacyHdTilk7RD3RcDTKqBRVQwvuzheXrblXCECCN4UeethRZmlAec5
Ma7Ics5vG8Rv6PZXITlwnE6FWbEKGzJt6H4pAFMDmr+zUN0lNmMfuLuLQ8besGIJ
aUoclYBmma36DRD2r7QUL0bOVYI3zt/nZ0QqIRNHJeGyX3HkQSvZ7CiCOHpewme6
Plf0qnV/MnesNzWPnHAmkg0P2lzIiymVTW2ixxHzVw7yEludQpXy7QckQlLleREv
zJBvwrcojBvHzyxSHOBL6NzVUM5daATFMMgEccYdMJ5Jv8VvqHa/KrcP1Rny7fC0
4IKhvdIGhyhpMD4oMmqKo2qx3NfREVm0H3jhv3UInkcMVsF/zOqJd0rdyTJm2NZe
Li8bpwOgZ5j6mSLr7i71ffN2bIcj/I3OWhCsoZb74HHOuDLlP5lNAPGtKMT4CpL/
UOSKGWlwZDlkENkD7re2lxkL+1+Zzj1anSorONlw7SMe1euX/wgNPxZ5n3kntGnc
+vkKoyt4SgjuLwMaRwMbmku9qM4SIduGgXXKi06XvTDo2KUvdPJdRn2aIQPMDLLV
RhRAbjclh2fkHXoXp7DJav8y1EmS9+kkn3oY3XmWCbHBrSLFHwSg/n3xMeHTZ3K9
AcacpgeHjepB3DjDEZj8ORSXsOSvSpz3UgpZ6AiONfDws1ddJXiBeXnHlzg2bVPZ
VcAJrWBh93/8qVmBaNz+gE2mnl7TaxJiLzBHsLpCmezQ6ZdUt2CvHPQWsCCVbyIz
ifbe1xphAzm6FcefdtGWhnioDAgxmOJshaOExpqrJxmBiox0HPjxEztY0ZwHLniw
6pLi8NsPgOXCQ6pP5HuKGtz9O1uJVG+VVF/LjxYbQYWmLp1QGKhkmaC7G2VXH+rd
T9HKOk0xFoeZ9hBpjp1WapsB8J4ggHJ36jSqOP8io6XJtb6O/GzvG/kOF6dwyVkQ
uDHhrJsW8FE7LWn+K5/NYtehTYgjry18O+rSdvR49PCTB0TyFSI1xSMLgdRo+Xse
UHYGrAbVYFPlRhpys7rMk8Y1+DOD3D+fXI38AZ4WKXbc01ifZTVIn7vwy4FxKm4s
3iv51B26r9yU2DPScXtZB24VBJJaMto+UGz/5nH72YECTFZWAr/n9z3yIOhKYxnN
6n3q4F/c5IrLPtHCMZD9WdFw76jJr52tZHy4/hfYQUl1iOqCzWd3E/p+k04X9F1A
uWcF3TCmeS8Vzi/mlgJP+FNKxMyKK2ZnHoAXWBpscz7/zJqgWzWS8GKlQaAhBL7g
NzcGr8gYx6/BNK2wFFe9ZlRiNAPjYjmotUW2gzs5oX/WqpCM54pZAf72ftAJuCwA
05Fnd+/6onyB24ipDgVRYZ6F8Ka6omo7b7GNtiQhVqXuYQfX+8y9N6C7w1MjzxQV
m4VK+xTtjywqVYQz8jtJgUKlxp/UYq1lweYCIma3fe4f+VXAtzvKH2pcsak0r7U0
mlk5xoj0JDmgEg36t+DjG+KxPDgT7ZAlY/cKDl4b3IJHj6T1CBDmT/pNfxRbdFdF
iKf1x8beOxpB0FtimF3O3luYWxzDUUDunNNyjZU9EDeB9uL6WZowM6gm75UtTIl8
6CYmcbmv0RxlFV6Fzvyxt1hmXeIk7wWje4XK19lPgwGnBb8DFyLusMsMDyxqB3N2
12Qgq1VBawedY8fmKTzbuR7XBkZopOUhzQpct0kEwYafX6gCkVqEfx5XwN9WpUCZ
fEPxy6Q3JBPkzKVtesHd2o9qSNbfH3P0KpsAMKorqYB6bZVplffqoHEAAAMLH6b1
63CtqWmUP52NIgRckczq476p4IFYxTZlIR/vjSNmcowjlEFecS8Dn54OgUVwaeeJ
c7QoRrFxGxCSU2YPpe/ixbBCDxYBiD9j/nwGQA0isTgKJFckn8KZOJtT/UbbOhJU
6nk9yJJ9PRfuuU3G/ofesT+E8Z0ipdWtuQoXxFWo+9xNWjjTSfMPJK/HO+/r3VK1
Q33Vg8flAkdLa0op7zbBVSyfaWC/PPMF53Bohvc1n83+nSFNxy5Dl73VpZj5/Dct
rDrzg6O4xBPwnD0ZMCBSaxG1bLCO93YXtAeFWz19PNVisBAH68mLbQnLBykEVwDM
jE9kWBHcN/hlkAm/Cg6peUESvFPqcDi80QZEHYIany+7FxcT7djwRtaIZEkJa5ab
0QyeG4ro+yhL5PL/NMdJV6dv5L6CQ7w4aeH0D+sMQZIfZwjb1nGpjP/Qr6+wAqNQ
XrI6yO6u7qIQrYON1IhbpKZZ46uzzOVIcOyjltIlbHc1+stICxKSO3a75m1U9Q+b
eHI/32SRVBmiOCVyq3JoCWI9A84Ijlp8jWgMm/qEV+7SOwLwT6UuqCyRutrBu5qC
Kwup8EwRoE4EZrvrmnyL0+VMFk0dnXyqEpEXFMXjsK5UNpT1PD+4pIqpROeupQiZ
pCs1rx/0h+cW1mXi/pX7sgRnHZQieCUtRicDiBtM0us23PicICSeBiaHSE0mxORf
LrYpjIukg1t+TcsckVqS90aBgZG7babXPE2pWjoiXK3bZcsMSbXUhgfYUwh0jVJf
GAY+NW5qe4byyww9c/bUQpS6/pm/NF27cKE9AenSC9AM+Ugxehfxdls7JPvx6p6S
iKSmn/9rlazx8gaoxDXOhlaC/mMkZ8EjudXO39490Pync6ZZnZeSmmwDIspM36OD
XK2hjNWMun3yAp6TkWgfA9P7/ZtuwQtoH6vXNwEZa5gqRDp/Jbx7XIoj8JUbToKZ
VUo4aDuz/9nJPesQz5a/zGCPYO6wSLDx3b/jSU1anvelc/oaNSWfy1uagJEiirtJ
uMtQJXRkYAFDItXuUR1tApI57bWVKoN9WkxmKWp0rdE0rd6FVUiB7r4pmY0eJoTp
aMCZ1wAXWCZBx9e/7vSsZApJfMVI1/JA6w9O4nBVdFlAH0Gepdv00t9na4HHWQMj
1QdSeEi5aPYyd1vZfN8vVIyPJT8tzLqDKi/SgzW+vpB5y4LwKk3REIcKaP57jIDQ
Io85mWZksgzvw4nlUb0ftVxwEoBmS7673D/WSDA6Uz/K4TWtwnUJ8bIgdbknzWji
G3S7awzVsFNFU8QkvTZqFKIaSFPDW8XITLI5+DF6PIV/oXtZ/q6MfCM9irYPO6YK
g7kGYKr+GWuk0NmAzT5ocyqMzd9a4sXhWtJG3uIqFrHqxNxjTd3XHHlWCkT4BpuY
8KavhRIekap9y9E7dhJW4O8tfOsCAoJsRVkFSwA/6D7o9PDAd6JWElKfbqMs86Yf
xIbsVHirNRPeAHGDfeIE6GiTM1m1HJuVVoGHqXKDqXene6RgHNKvaYu2uL3VioSi
3wCZsDPh3xjEO81WNcsM7WDF01lWFCyJvv4/V5I+oot1u5ElGb9pbFUcpW/kG3H6
jDFgbWB19I6Mhz4oWPMzcbrMg3Sc7pU8DBstaBO1A4t57AykW5OBNksPY8LBdSks
1uktuCJdPpci4FfHvNWlUKIoCUFTi6qQg4hiuwMiF9Map3nqBq1QP3BExq61DecV
RJ521d/53AiRcu8iL3ikDsIuFaXI8VK2GGxMmLuFVjerHeRE08sl/iH9CLw8Mte5
73WBrNyEb7ZWO/s8U/TC0/WI7/s27Aobklu85dsLJwuLCdadPg0QxAS5hUolQS5s
3I43OaCLmhYfud8m0Wp/d7xFwopVaQ+oT71H5FbeLyVILeT9CtdyJ43ktiyLBbm0
pJ34UsLhFjo/p7NDTo1dLKkts8bGLagQF+kideKJCqQhiAVnD6xcsUseTc8h/vCw
F5TM6ZurP9BRFVG5cQnBh9eEKmcs/ICoM7z0bzERc0LxZcm+Vh1fI5jJmQQEONvb
2xsZJ5mVM0mxLZq2iLNucOTggtBKGDigLcuNw7CdPZXWl7C7YmnTjXqeOVMbymn5
F/EmvAB9dxEy/aNJl+yuElMQ6Iqh43BQH6mjscEzN1xWyEdvHeNlinH/7b23YLST
uFUYI9ISeilNYMmmqG7pv6Br9WYH5lXmfYD0LrcW7upVs8+if8s/flotpOzpFU3u
cgAslcSG3c/JOrL+mFNKi8yrUmZsdfhgDPjqKBuU9vyk/M1NTwrI+bjG9T2Npd9s
xVrjzkHAfWAJNDhFe3TnsrEBxfMjpiVq+MKmZk7AjOatcOAjGyK9ZIDMAOuwo2ag
iWILMhttQli2xBrryf6xFVDh/gPNJdnxL1tKBL1wXMRZGMzoV6G67Kze3p45/t+b
Zi43d01FY0D9HZb4+Y07beXEguaELvmk9cr3+2S5FVd/F6QvwwuKXaembElQZm/3
x0JkYBw/4zN8EjdVSyFlZVV03RvsJotLHVsTU1zaHucTsV+5hkca1p3g6PJ8lpHJ
BzpDfOVoy2Att9QgV9T8zazZdfQrIuGWhPiNovwG0uEHCm7YVGWAlu7b6e9TTSOR
nmnNiFdfhk/tv2l3TSw75/tXKiIrA5ZxY0zODh7CWovRibPoJHFL5Yb0lRTUFHNe
uMqeHOb8QLYy6KmSU/tT04W66Ow9Q7ngKJ6wSU5zUB/neXzRTvtciTCQXLCYJre3
91K0+d+JqXmm2HkCjRy0dfsm+djck2jv6rvkq3lKv5Bz1ZeDx8ILvAz9rG+gqsnG
/D5qP9bO4CyfICS2eC1diUO6y/M5sBjku1CheS2IY6WTv35FQHplkN9DpQqHvydQ
fQ+YGCiTABm6zSc2tsseHflGtGiLHPqNxdbU1Pj41JMrDjItpwO8lkpYv1q8MqbW
/CTwfORVZetMDNmxDNFl6E6X4Rr/RDahv2Eb+apixuV3q4mZ3tQzcrFdFFTn4jQx
wMBHaIG/LN0xQK3jBB6ey27QsiIK1KWf/cjoGY1gVaf9t39rZibpAGYr9zdFhD3N
DqmbfbCY/ULgPi+Mey4S2zrYsXtB9TyTtepui28nVLnuWBp78BYIZN7COL8eyQGT
wKSTuzDj99nZrlaTtp+cs0qpRj+lYFNM9FFy8scw/7WKak8+nw3SUcW12GuT0lz9
y0F6jT+2bS/5rh+apEyaQ/ShIK+BaoOvx9ALJzhj1DkjqDae3+Hb3rY61GCnWGZF
l50dpjc3zQgozkqViEiTuM+L/VR3ErIGnTy2yt9qsS8kZai+BAIwZY9/h2WVP+4B
ilwJdGY9bAvkxVkFzyh34O1WXFCUPk8M9oqsCMOU46rerZ0l82XE87CWVRkzBIBv
r3UuHsLgKpwP31Sjhci/K115d5Td5M0fu8K4UxD8x2/pn4e7YGeyzBNCw4gffFWO
OFC3MZjfQrS42OLa6KGzi7of/xH3Woj0mdjCyEDJm8sMnppaKZlJwS3UHquu0ZoG
1CuscOGENPdJCUPk5kjaJmI899Pjxqgt5d1xC3he6xJdB/PLHSWScyuhVefxx4FK
38EUddzBNwq9HjIYtFv/r0QVoaOc27GMdYwNca4QMHMMiBK9SYzP1mMaeX4rtLb2
uWw8hJT/xtJcL9iRmE8x7JHATqBW2OJU9WS7/zrcPaBTq9N+6ddAbc1QPSabkMqP
X8vIy79JtUv9rKXjRUi8s0FgTG7pLXfGe+OeA/jRYXSs69Allf9up4AGOgYgcbJA
yx3BfnyOug0hxikq7fwWtgIlk+N43JjGlZrPtPtyJZ7eOOQ05YLsfAqnPkhOcJOz
vy6jQ1bN61O1Vy322PPYyzIVBQzvdWqcMbHduGuWjsQYd1JT2GCNr+NJPuDk/Faa
wV22xVzfPYOa9QW+2dwQ6crQycBD8uKAojtMXFKUirYxXZFrGw5yEw7mlPMh6ny/
LyRPa3vISylYNC/MVj10G5+nsl9GR504lmbqLa1Yohi/NiVkLs22/TiR8jsHE9JG
YWEkTCxbbwv4MdCQ449Wjx3hYSuNZeHMbFlPqduSSxESQsSD4Sl+wk7vp4o5gyjt
0prpbVLFwvcXg7vSDEx7jbSP968Itao/ni8jUY0M3LvI9wDUksYsiOD6yTh4Z2EL
GJmPTPCpdDbAVLv56ZfCYvpO+l7nDqrDaFBQvVJsQpQwnyPjVviWiNB4ltFb5Txe
XUONlM+HzSoWX3xtjC4cLH6vJjkogRXNawAUszKNEGnowKE9v/5EY+q1r7yMqKfm
ENn+U384rCOERR9n+oaWpiLVIcWVBw6XU46rcI6QsrD6gGZInkGaWxHylHUcX+4d
MXmH1AFKF8d2VMPSNi2UFWBD2SV1Q8yCxVe3xUwTvbvaoWf4J1ZovnTkkGrCnmmP
vwK/sseYnENIfkKtD0rUtPWkeUFEcXMHci61ldbDdfkEq6gaBuW70fRu9ntolhbH
xp9Qn+eDu7xV7RonIqF+SyIh3XRL6TiUE9bySNU0ANBgLPrHLPsUhmNtqci6KbGV
eldRoOZ/AqQ6X1mcEEQob17bIaDg28oDCvlRKUtIjfFdSEohxseDZVHL/goAOQrn
XMtNj1tqOPHuF8FlYUxl34QuqPxDpJ8TF00yERHLl54cYlYqybGIHVkmJLcoIsmA
d1snn+tyMnGMfDdnkpcm07HwrU1Eaz01tg+yMisdrNK97OpnfHkW8wv3u82FQlbR
7r9j94AE8TE9FO7UeztdYKjWLg2lNZY4f1MbzxGmPwf2b1HXQGZZgGs4nZtuhgPZ
qUxdnw6zZRzyndYyfy/0myEnm7tv6xIFiHexYHTwMilmzXOL3nKaGSskflvwraPK
k5NqZLv5O7XbOkrsLdMyMPih7aInJYYKKrctVaB6sewz8lRFv3RRVunDCiSgvBja
pDg7Fd7Q4Swf+mbpY72hNqjWQukDfOHf289F0UzoFl5hsluXHYfQ+mZwMt69mAi9
U2GHdL7JiJkm/Nht1Qyg53UA8vvCCJs3UcdPn1qFfSdwiLv2vMdA7favKPWJOvX+
7l68twXKImuG4cgapbeFdNKnd28NmLRmw6GKwcRVwpWUeAwHY3DON7O+ws7J4BDP
FqjN2NH1SzRiLRTSe/bZSeoO/PzK12QUwkDvfLY04uy6yB5HgTBJs6JJ5OlvtSTf
H3/p+KEh4t/rC6ZaeSqKagGWLPuB6xQ7TwRVY/vq+6y1UF0DQdGPOpX3hXBmyxeW
Jbk2UBUfOSAJvPQVU6F3JP0uOf57CdVTo4po/cYpvQXhiCybIlI1nOoi2ZPF7z7b
Y/nkIvKZUr0lMNtFCngUgIcoj4ohgUiuibXVa7lkbwtSH1K/3R7HmvVsBvrHBQte
/YazkAT36aIEq0FccxcQ5k6di4gwG4NWG/adDBiw0vVz656YvEj9TTRx+JuWr/Nd
AJtrU30hg9e0Ecoa420jhVGIFUShAlsM5BYCwF1CjTXu4fU0w2rddStbnEYENqH0
um8JX4tiK4/dvbz7v75pORXlkJCOocwxaKptU0pXRPEJNXZx/iC1gSMi1wMwmLma
nRbUpD7Rd8h7IZr8aJozX+FJqc/bYrZqbKw6blUkb4jHuM4ckCF+/HGB+VscWvik
prqhE/VpK9/EIPBHgB1p5rZ2erWdtRLJLdgCYg2UtAJNSOEEMl1MfPIenvgSspBt
bA58BgPG02SmEiShiSky5zkzNqxOhVdfiVJXPsjaJhfiE55HtipS8fdpcQJrmdrb
Bbk34mpM1YwIlZAvp5y2SJywQjM7a5Fn4B+wS83iWMDumIL+oYsjezfLLqA2MdDS
Zwazd7kUOjZ5OFzdDIk0+9vcmnenp9QIGsz5sfk1/q1ksayZyrtpnU5hPWijs8FT
gIcwkfqhQqL8A8lQbOA/DaK2pE+bPNO7RBk12tmp3eoaRV+hmaA8YSNOyoiYPqdN
7k3dDwNYTRsFi5ZUxJMS4n1pmMS10Am40SP2sBNPmo4Fn7YZ1xlcbB0cTFrKJ0PN
wbcIbD1RoTp0iHZKPgn+CQp2o+FwvGbMz/l1R8qKjAR6B75ExDF4vJ6cmK0aXeIs
StabDZMAQM9n8DgDppyNHUwcnS9hPMjmjNOpOrwE7BCZu+Hwy79rYLS7sFU5p2l0
ZyI9qcQcdWTN7Kd4DY1ldPkObGgJoXmb/sKsQA7jn+aaDrqwYiGnEbWp9zSHA4EG
NbdYPd6jQTutveIuSBJfvVXlwwdEIIROc5co9NojfkhseBW3Bk/6Er6Q2+VumIYa
CtGdr6TWZgCxd5u47dcHR4faA3StSVWlhnV7VpbjTwlzolhpM9Qk/4AvIl3RCfqv
a+ucg5arJv+GCdZhMdVVDbBIZJ4JuK8Z/9NHerkRCVLnTXtf6Ju5HR7Vv9rUN8U6
XrDbLyryKZVvdNbvJ4eoWwJvp0ACYY6sknWxI16lFp3CJgMWR1o5q6fVxBDgnI00
PW9UmSrZq+JDhKwoq7uGwce1q1QETG7pFZE+jWQ9LEERDt3IHMuZD1heZ0NWUyeh
OhwvopvXJrdnrA4mzAzZHFAuVmL6CHzKt5DcOOXTEC3xV5i5kM8/LkdjvHVOTyCO
PoWO0loeUcy9mgQg6ModkPE8AW+CyuOOmLvkiobmsDXEeDD29QUvxax6RMLHt8cZ
GWArlH+DZc+gNpfJZIL9Na5EUVTuomBY5doEtSnoKHlCeI3ojiTl8HOXu4FS7jng
L9UW50ZyU9HF+cyZ3cBQbEJsaLHXnkH2VChhjIuS/F6ILYD/RAuZbBjv8I6DU1Zb
GaNhIgwsmTB1JDraWA/okkyH1mJPshAIWpfkws2FzhUOEhCVuE6sxBY5d8Xjtr4X
60QIukswbQKDzV8PpUOWmL1yR5cBtTN+ps4AcXx/mtPB0m8o0eeSlQ1NQmibNp/x
Q8iVHpeOQw0Wn7EO+BSB4j/g6oNnMGk/6nZ3mUy1Orm6eKDOnO1+EsjXOrQ7+f2j
GS8xTJDIrnKzzOTgkfKiOJDwjjnJjkfqLkE8P1fFdV0gvH52H8A7mRRKnYnYSRY5
Sb4/Ijt7uVUkg+7dMd9Gwg7O39jjZtxq2jiHku/KdZaDZn0MNnJTuXl74nyQtCW1
e1dq9Xq0AlZN7izQhiRqlp32GtLcs91dJRUOnKWrrCP/2Ibg3yaIXwtsXZHhT7n1
I16St0zZqsboXehUmDsLH59HRh71UT8rVkP1TI1MipmpL4PXB3T1WNRLXUrhvo7S
cRjWe/eePtcC26IZAhpKgaSV9vSp+iwbSuc0HzWDtIHl8jFZ7KV2ZS8KanRX/I6O
Q/2H2Wb2UrBKkqFg6GcQF6vii0pCi2rBOgSnpm0AG5akefdpxci5i/y4NZuaWrZs
3OWn5uK6331M7/dxlb7F/z4r3lHM9AWtbf36ZqoxhzPhgXgQtq5grHWMu+Yipkb9
9S1Mk8X3LLoPLveubXgrlQqOijtzMYqfxIaFms2p4xR9lEe1tiovPNzirIFNAx4c
tdlZSoSYqYu+84qgI5U8J8vW3zgfvwG3vkpcHsxCSYYJn/7XdUTb/4X2761eIlt/
HKSH6b9fZSwKeXN3cgIBLDRJ+LL4rTquGEhCyClYhIaQ0X7sJtgADXXoIO7Sf0J7
ka+SRpXTA33dg1orArb90f2kgESiRi2zT1u+yOnxqlu1qRZzvkYSTWrcP9sKepbF
e4jCHNnrkU7Dq3+uuqR9vzE+4TSJRYI7+RbU0G+n9ad7i+OV/9BghBYu5kjozNap
VnoCEUVKE0t7K4ybgddvq4/1ACG9P9mt8z6A5nKQEhcxb8U6oleNFmtK1dChgvfV
q9iYFTt6gMlITzfCFAArS3wm/b1Vy3mX8KL2VxwOr5zXxbgF/gKUU6GIAivv/Oe8
S05VcpBjfFKF6dAmLmhzs/lN+LIyfJ6yoAeBuywzXtdCIdeaG9OhY0H2Nz8bHgSu
f91uDn+1zED7aY8QXI2usGEe/hKL0MEF+ZsXPGY3M7ghErZwp2rlhcMXtNOvXhPW
E6yU/swYpwz8KKUmQUp3ssDpr7OQhypih4+9Bx9bK/95fKrW+NCJZF4K9IWs4uHh
xa6w7V53wxbbGI3qcfp/qt+6TQQkPLyE3+JO4U0Idz2oInIMhP/cMg+vXU/1Iq/N
thxX+94qAp+7wuuFZzM6vWxnj2qSKBpcLxu2Hv8nTFsNLPFZD3jLJ65dfYcL2DtQ
sGUDVJ/9iV3J7cxd5hf3mLsC1ww4s25cdwI9Nd6auBR98pLKY0n7aOlfPg5Crg6x
ShpNNBu2m6GPtvhgM3BNHVf5lgmhQSsNCRdFKxR7Q6kUx0Z1WTUOpDbQD+WqsH/M
8NjJXIOLpjg4mw+kR4gYsf7DybgRKFzVcjDaLXCwvH5FX6eib3LjL5nllz4JrfAz
8diZNiEWGmyqTxjn5Zt22UXIrlkqdkz2MygOVPCgoPOsjTzgY6zaw3lxJKbWr8N7
E1LPXD7/VrZfrGLDQpahwJuW8cUpfoZI+cm+rgwnb4QMVClAJy1uFVf6T3eUHmQf
xaAJeoi/PnWxz7ZHUkx3IiUmjpEBaoLtJPZf/n3BXlZlmyGWU53CbWiI7j8fqIaQ
YDpguiFBj5ev+YUTDONFaIcFGzbE0nGM0Arxr67BVzOQGtTHsiH4d7bJ75naQg12
A87mColBQprS1oU54JMi7vfRBwkOvrzSEaXfb5aOOQwZ4SaZnHIonQ/QAyZPmN0p
W6P7/HWtKon3LcVDNixe+cl7dPEZZGLbtTnkOqdWOSXrjMnDM1dAo6TBx4Llao22
ZpXe53MIHUBJ1IruYZVJQezSqzwuayEM4/6gmWMSyA3Q0qRO8xlNYXSWci40iTUa
cKTbREz4V3aA4HJj4m+KopiC08pRf+j6hIJAMRqw+UmsCzRjtZjfwoMgZugxYu+6
AEnxVs/Fzdm1kF8nyzOGom6lQdPHiQkNkY9XpWD/cHed/xOmZTIVIe0DJG0l2qF8
zn9OjagLwc2sSaCTaG8qubn1krSEnfZpnxHA6THbnKh5G2aNtPIBlQMdLT8H3WfC
QAQkELhIh0eN/yrSQZyvsRoegX/k0UPoa4Xy4dKWSE88QPzQ5sWKuei0PvcycC5J
6RUKG7V1FKfGkLn9A/bkTsNxh/J2KvGb0qxfWI+da2pOyjiSMusi76Q6d6lSWpBP
4bgEi92meUpYMvZiy0GCyz8jMke6BGLd2Hft+ntQslQPUgd+xtbpw4ZGNAB6XQW1
Bz9XZ1ywUvDuzcd7Jc+YEjs/hfwzCgMJ8JVNH8N9Arp7nJxsayyEOiW0UVSfGPd5
kuF/cW6cIPWdVpKnWIzLO6IZPZM1cXhKsz+gzjYw6jfjLSbm7DStVXAVefOqAZIa
sAgSa2QNvAP5jqDCeKOHlTd++ktvDsCd8NseHA12U7/yI8G36CN8196OmXqtlDQ6
0NHh3aOLYsZHCEPJoyC9NzVtmfG8uoNlmaZO+gX9RJVJjSNXhuQPOFYyEerL2D4D
J7s9FyynbjlREg5NH+PxUh+0p0rqb2uI+QqyTcQteqQ3DGiE5sD2k/2UI/ME0W7c
+93aR3Fqh/b1oESh7I42LjdqvtQfNXbtLDZYxlrvb/RY7W52lNrpWmU+/lyRBoXk
yZWwPJrGQWlMXodL4Lpi5wH5sQk45wTFDRj3Plwf5Y1D0WcM6XOtzRv6Y03x9Qwm
FPjveKYtL9JLixRAb2U4BoqmDL88stUuAC3EA62KZ45gTkjqIKl+D6/G7nYHFC6n
HhhSo4vVgUhH2fT958pcdlIZASjmuvZs/nO3a99hKLwF+ggi4pACbeq4cOFgLnlA
JRA3ZlJwIxds8pJtCotMaq8XkzCvB1UGc5eLo2kOFOEReR1l0YxBEMfIMYO3yrSG
cJPNOBkzJUqUH4vBlV/8eLBo7ZcxIzDK7EdAsqrNKg9QQYEtmbs3o2p56YFPsAgw
qGdwg295YznH8XpJQW/kf4Yj+JiucCBhRQMtshI5xTBd4pyKuS/+iowQODNvPa42
c/fw+2s+8W+IJSSiDRf3aTPlzrsOudl1vrt9gcOsr79CNGAf/5obiQSEtouoJizf
WH0VOJlkXeMkuEDlgMtX45GIJfJmWNZbnm78TI/NcM/hmVL73J0rzqLZDTp48gGO
LSJprOWvMM7wmIGaKdYnkbKKMABvU1vVWfJ/xW6fMY/HAdF901li2MWq/TPF5bWN
clkaMKTxvpFHxO4SJOIlyPC66impdCV7th1FoVwmIB80RMHE+6+QbdK0oW/5NLQt
t2uOHhtGSyr7h+BxxdQ8ooYKoO/tkDMDXKP+4TzuY4qf1pZym7QW5BQC5oYQ8X43
FycQ9ffMtJ3pEjBmnRI0T3Scvuf/DVVXWfZEuhXhtu1KDJSm2r4RGiXBQuoU6XlP
CgbuYbR0LiFgEgwuJh8mNDRLzmWKWzPHIVC+TKPXtPVrvXLFvIvDSkShB/cYXeXF
TLul2bF8KFkeum4yqDDSCCGcxXbHh+XZZ8Ev2ff627gGyRpxbxKWvLVAg/HuYogw
Hmx1W72vGhg2oOorLGc0sCmJZAmRhj9m3/AA0WCfc5U81Vahv6yLVq6qVmSkEKCJ
X09GERFZgTjDUCKynBsGjChiweInsuummpNbAwzrnBzgSzZ3oyhMiyHix7k758+T
W/MNHxz2OBDNLLXV+2iNlkEGSzNAg9M2IuQOPS/FHH8gPMVmvgR6HwOvJvr0FC6N
6CwgePPthqgBHBVzc4TjAYKbXuFJoHQGDQ7tS8nhq9Jz2pYokY1xZ0Pk9qaGZU2G
zglMWiuS8BVQZQ9ktEXXBttQYBeF02Cc/LQ4M6tIrHx9YJRlIqJPDQjzDglXKoTX
9fg6Lr+CEV3qtRzMLqeBZYy9+JGCxl6MjdvxUEO8vwEwQwdBVplnZs3nvnvi2OHv
ToRyxTNUEY4p8hUUwPvJJk2k1Cmo07dimWmG1sy93pO7GG+CKRsADrp1w8qozJaq
FW35Id0wL+32JTXVXm7gfdQfdrt0yHIjxNetEY6qfAa+AdyhqGGoyFc9yx1hO82U
qOD1SR/PQ+WPAksbiWwouA9jWjSJYCTQLd81Ouy1YBKUObXNk5Bls7RXw8Dbj3ua
ve7WrAjpoS9i98DqQNy7u+YAAWFfwlz5ItGaI9JKaNQkwjQ1Tjgwo/2afZ89dT4Y
ZdLQqOGkxbg9CG8/rClMxTQie7DC7qEoTeHk4s7WaET85iLv+tq19onCThFPPnT8
rnW8gDvers0PrYulzGaxwpunriIOtn/usx9ZPsEpfFjb9fiSxP64wQnO0Z8oXiiC
580S5NJ7oFuILdN3lCfe0bZDHKdENf1Jrf0JB+oqpigWpyN2j7wMG5pfd8xDfa03
NIBeKULCMQ94AQxzM6y2UveSt4R0fRAVAdhzD4e199d6WWK3Mo1iS8kVKsWMbZj1
Hj5QJHayxBr4cDSnk4Uiwh/PGJfA3zM+QGZEMy1Sl0NguMl6Jc5yw/+GO/7bbwW+
Wga0V7VcSkCgS4Dy+1HJA63CYxZmqtBtKm8UaPkb8IGxoZo5VkNuzjNWePSOghFT
sXOUkPUCovy6HcjKi2mkZ6sTT3FdyTUhPQjyQYMfP9vievEI4SErsQ6OEa9f/BSA
CiDX2+0/Z+wzI8uwDR2Wu4bKjME+fnTMoCdI+Gp6Nym1rLpy05c6fO1yfjyqo2iq
FGLtbKLMq7aCGu2a1JCLTO4vNOVncRUPtVd0ux7401n4P3kCEL5pFOaP62wwowWW
bIj3keSyjda4tkl0rway8HWt1N+9rdN4ZLuFBhkt5FPHkuu3LaRuA38wZvKpn+ef
1rxq3qXUasfV41h4Jgfz9IgDWqjtJ02/1k+akIsYCdj9fqGU9/HBE+VCGtOudovx
p33mdL3rjhiM07JPfW+a/AyEP0KdMVKr0oyl7TkG2YgOIEvSqGMwokCu/8JdMKBW
WsbsEH36vxu16yy8Y491fo53g/z8gp7HOzzGWDrt6aGrHFOq9uNywDJn3PCFs91p
qR3DizHzYER92n1F7Y28XkZYtpX1us7tnQTJ6EPzdH0/l55+wFWxA0Bf3Z2MmT/z
CXzhCZeQgpjZvL/qXGQUx41cdlpTAVkyvO0ok74V/UK0y58PUxnnBwsfwT+U54KE
+he3Z4ZCLMOuM1rdzmX/nbJY+bYvBU0MkD2dHSZkE2/PdvQNZqN12+8NWZswHj9j
EAwKtQrs5p1vQMcWaDcfbSufRX4vhjMxnVQ9U8F2zuILRvLr6Kxukxq4MGJf3gjy
o03pnSraz2aszWAbo7Q79ZWUPCWwCJLxN/VKJbaYxIlolI2tfW3Y0tB9pm6Qbxpo
6HClc3+5xTvVsdRCs+fEETjIfXTvd/7lBBl49xxq6xPjVSMsFxe57UfJkf53K2Rd
DOePbcXeHYwxZMH0osgAuSbiMWvD1kEMNZy37RMvd15h/1MxlIkzpzt3SbqW15OQ
VUc8OFDGfC4Lkpv7Zg8I+LVjfLbTH9K4sVm+IVcP3ObdUYV6RMebwD/JL102K+/L
l+VlD+PbtKMGltQ7M32z7UK6aK7E9fhQTpMwW1Dg8HcNa7Xw9jxP+BcP0jNoZ8PZ
Z0XUM2qIIZYscsaLgqD9NmLL40CcIhs+rmZf4NZaYmNbavP0W1GmdHOPUj8OtAks
NC40Os3hYwrJMnA3sGo0Wx8oJ7RpkCAwK4D7dyvollj6if6sZQhl/uXKY1CEeu0Z
c+EQPFkdmeaqCOKjCin0NLYX6si/Jfrie9mEgZOE7Q7acSP9JJY5/ESH4qWqqMRE
KSRH9/x7Fav8ikDgxdn+WnAUnajduNh/oqC/eWg7IsUhCK5pe8voplbJH7wxZBxI
VUebM9MxoKA95hKS2Vi0xdMbTg/ERKA+JZempVSdQCpEIvKOTkNyinbSp5Ho1x3K
2qN2wNtPoRzaEoVCGAcJBUyCJ+XdS9RKjeaH/Vun9BPUXj3lGoFsS8UVQnQrrIP9
cFGuLCO1R4Aqs5bs3lCyD9aCOMpwS5jva2IjcUWoh9P8pw37ueBeffF45mB755Fa
DWSnW5A/cx7AysI5K5jEzTOsXe+W+lFTYzRSHHRY8uDyqWhyWSXF+VLr6IIT6eHC
98PTdaiJ8YfFjS6+6J7tyx7+oqRouEUk0QTODM+YbswNet1HBeQETU4QQ2FIrDHo
vdX4rdHJmb3Ogbsuv8K300vpiRuYaFItSvVOG3o7WXXIqj5av8lhfd1WxxD4+6LA
1J4Q30mASF7wWJM4yVa9a6nSXgFly6CW4jSHkWPDNx4rZK9PYGFE1Pj67JJuE55o
PEO3H+pFVV+kCK1Hdojo8/jhpqflb8n8VrHRxYX546PZ4jOl6c2lbWVnysFbmKQ3
B0vc6BdnjmeyobyjbX0a1zeD/W8n1rIrwi72PM2wXnR2Fi/OPvx/G1MKD+okJO9s
xAtvbUGqNxCRuoI9TSA4MkGuugjZwDo44gF0Fw0zqkoF/gRuSLyTD/l/T9anQynd
pBzHti6vFCD5xL7+LCE3Nwn/QvTP4qeE4PdgTLXR7N260BWhq+8D1c8dWg+lIxpw
UN5ITLWjoPyldDtelf4iTkj4K9cSfzaO3DJSXi9OyXOAMW1eQZN4ONnEMcm51ckL
nMitRCAuxijkSS6sq9uNSkijbhgLVgdzw4NtliAd/HJBGzHr0JcughdTyHv4wvcN
CNhQrASVXsf5nqAKjILjPT4glfxVOVRUzzpmxxSxDwD2Ddv6CAOyFyHRBW1EoHLS
OkSe+UcRCdyl8wpLQrdLrToLZBpaAnoVSoJmTAKgcIpovVzpcgrqFx9njmnVXvjO
TxA6mVLzVNvlb+NbNACD/ST3lmPE0/m+01487TxMYc/mpcrV20Bp2GFRYROSMAM3
BaoIboSuhTERGPXuQAYi9dPHLetXzPrnSFdVzhO1SjUNx7N/Oc9YI7Jd7zu+4iLc
xFzAkXoUhcCOk8QJ97fvApLvc3bnVD4bcAahf6BVit1+6vOr+xpVX/KiUXpLWUeM
BHujX0+RLiTfNYZoLh+T4loMGzQBY0DgrrsaAU3zyWJ9CzHkexLb8KD0a8S/ur8p
6BFVr5TtSYHuuW7drc19TaPDl7Sh+9gQY60FGTxwWzW6BInoTO2FXhmOEsQh2I0j
Tl1zYTM57xCO7M/uG4Md6yPWeyRRqwk1Sh6eQICixps4h68uuJWTH/0MgfAPq2e/
ybMp4XsUGGqe0dqsEunN7nZbDVLyStibmC9EbWwCoTSGfNO1jwHu+vkbIOyPq/2/
acNyORBhz/LV3T0lo1He+iDNWZ4ZK8ua8xB37isnwg8d5XIix/Xs8l85rwJOi60Y
OK0SAs73vf1eFPVaaWMZI+9XiIkvCgD2DD15kNxAiG0ziG7Fc3hOZYfViSNQxA5A
33BQc7yuOXYT1TeB89B559fWLzNlkRlFu+96q1uPVoKkYNQvCsS1x1glUDus6gA8
3prwvLVe7mnm2mbW8GWJhCgh6e9TMXySN8fAG0gVNWx36u0IItl0IzMChnxZH5mo
Ck7sloCfonwRGSQhpPuC3Ha/Gj6H3dJdaaF3rnPsnY1IDfTYlyZNw2AW+Njnum8l
usxkio0oKx6RGYFdxZWy2F5/Pl4gHLMVOh/S0TyAgJjppFuuNbd2Y5kATwh5/iLR
tQJtQNitmoSpCQUah2cnoDm83Ls732ENynNCLtNBCtsj3lX0MapbIqHeKT5bjO9T
KJl61qdFzXqVifqzojV/Vkh5WKmS0EQeh5LGZ2CnYi9sZnMCaE5Bblu5h8KL7Jw7
pPDi/Jn41p+/loOeonrY33+1tc3Peq0uxYrvYxYNoRdg3dpFdGjuuSKFjrZIV6UV
lYRUHcwYjOnlyrH4U4vHDT2gOO6demFj3FEs+e2hG2MuKcYKvMbWev9BbocWZNAp
oGin5wR4kgvN8yuTG17/lYkkfqST2iXd9e9hWMh7P8Qze8O+y1N7SBladREYv5q0
oG/2MUfd5FH4V0IblpMVxXcnGBpaxaC1ywilrwElJ6vrVwAYinrwMqW7ZR0zirMp
djc+wq+Lrc8JUUpBhKc8BodirHDWP1TljfUFb0zut926jw5enxtvpRMT6NMeOw+/
pO8u65ttwjNZ6eV2jgQe+sX5qlRzFEBQxi3dFp+IGzkW29NZYA913OpmLOUohK73
5+6IZHDWY5+N7avv3135CE3jxicIaN5XV3l+ipZDsMQOJRiJ3CI658MHBRO1gY5z
bLC7avrk4zc8mCwHr6DCMnp4Iaew0yxzO1qJoYVL6Is/2Ou7Ihp98UW8Y1kt2bvp
pU2mQQOhxD7hWwzoV403A7Tj8pIG4w+JttTbpuLZSRZ0TqFzy510Txek1vL0KYzn
8FHt5cCeRcw6HQ1R7pX++ItStTpiAsj+Mak/JXJ7Dv+nqq7KV3F8SGuJ/fwJLjnw
X5kiDLCDzYy6MyiR7BOxnqZUqlQAv9+nkzySfr5wglK+3xRRL15PRtASxtydzjPE
GvKK9qukGMUlf9u155FAEszm03yfQeNRZSetjVUr6xbmNVtrDOKrk+z8/vM+TSqg
KzEKYgAY2i9Ve3C5V0BN5o9ZmwMvwX4IEFqlyBHF6f02XGDMMfDnQg0F1bdJe7y1
keaZvz4QSsRiguCXJu6pEDPP5rnL4M2yTqMetl9LUjpy11DeYlJicuZw88SS5EKG
lHFWJORFZGjjFOv3WOuEAa5RvTM5lB+0LDikXNLINQ2ZnKZxeypJN2HIVFA934wR
q1CUB8S6OoA3qYjyuq0MEoV0UQeRxe2OJClZAk8gEB5P9l2M8ANLQmdk7/sqKXmo
9fOwvtehBobGTErCM64VhggXh7mEeqex9Pra7U1aqZq07IcBOUnJ82is/23HTaZy
Lk9PPzCbngE7AcqMhtoDGG0qaoz7uDDLqL9b6lBEUQUFAelPPgge+L1Tbr1m7XOg
ftFcL58xVVuJvyMzExPhAMcrLbh9Jrzj/6jzB6NfOdt/KiWfyjFZtG8WXw63iNlB
Fxop3iPJ6NMpuBVgXK9yAU1KPn+kQGWOV+XSqv5t0C8rZxbJ+baWU3iqjKCkj2nq
FTk8JmaJhFi4gJlv6paZsDH72lEw5EsyiJERPJeWpt4QLXAh+mAdaTdfx3xI1+bu
5m8yjfCLtpNI8mq+C/+R0Jq3Yb9PtOVqnbYYSI0h04FUoPdOyLQlXyno6sIDNyKu
mEO4OXY5HU49f/8naB47hPGH6VqUpWwv2bK6XJgzKz/NTluOzSyuGI5CI1dql5ko
zNhuRL652NX5AZokoL3Ym5nLu3Nxn+eMVD7+D3qsoLTv9VhRXCytPHW/AHXo3s8l
5ptG2Aq16NKm4WSMAWWXEMeqsTz5KWifKg8YDIJN5NzjJGO/lUnQYa4JAlC7DFiL
x2+6YGuq5aLp4rbZg154PsmYkerN6XGeYGe0QphuaSQ7txt/rPyO5RLlM0fx4IVX
CggxunZ+p72BTHfnc7Xn16B6agIVvWtO5PPH2LE+4cRyQ7RtBaEffFXs5RSvrzi9
eXf+Nh6mGd/lZ/ACRh1jgrb0RzvOBZHHsUSep6eaCu4m5H1pwVqZNlLeeiMeXUIk
+l+3pOLcazxq9RB3cKIQiB0W0RCkKRNlwZ96ni3Xn//PoGxCDhCXFxJef0tFqNcK
jLJs6M1vhMugG4YKBHtRSmXXXHkv4a/Td0oHKOsNeUnxCBWftjLCGgIOfWU0jcK0
sjr4RXhPXX68HUbVB69sBNkh6EBFHoACHUGGonNOH6oHXDEXau/Fo819FK+P6Xxw
3AX64o9Fy2hS7CUkdVJUVsMCBkYF49xdgxNtom1g1KFRe57wdNB19emR3yJC3cAS
l6d2JylMM+LOztElUuLpzFn/vGTnNS6iR2kSZ6CFD9XCtQbtPO3slWgG1/Qincly
cSVwDb/ix+lzz7FFhyVQdqDZmbWLENRcWV1V5XMG4aAl5qNhhhPsEMYssmnQPa+M
B7muIajF/NmidyRdkTpuhJNiRe7Dzs1M8ZMiTnuwnuXke/tQZso7etkwkTjl59ca
nVT0W3KZMWYlkagqPjD7k/BQlwT47+9t4LyvQC0HPVQA3X9UYu/CORNIPalsTfiE
Y5bfrzWwJeHf3hdAXAwlt5UezzChSN6bnuvonH6EuFf2uUgvmWrwFZHI59kbzTE0
mDiKTgz18iJqyqSRHxLUMfhYGRk8YiQSwmWUFgffkHYIeVKao0Ksb77xnI1G21Tv
cMILBqWlMd96f5vMNFsmLXRzkpsWJ86kbj/Q4KzkgvGKkIrU0mNJlkqK5H2NPMPm
6uD7ghNhhwLByaj1gcaTyF3OwSyCOBQoU5oRJgpHfN/TNJrhRECQlakUeRWfIzF0
QaptnAow9EzKSjyIrlcTbisQre16aVKjOL/cX1DHSnljgRhb2NwTTMxrzTpukZzN
NPAlSgpaCjLPXl+u99ggN+aBVES6LZltcWOu/HXD0y8yzMEVGuYWTrqepfbhZwwe
wbim0C0FRvJJpqxcWpAFEhULkXIiIiU5uo3v1wvxGpTu7i3QH7VCd6xC44u/ixEY
Q8O1yXoY5IhltCByVoopeR7jLo8pMFYVYwFLxZ6T7iHxfDaCEQ31FFtmae7qpBv1
1+Mlden+cowVQiTDiOq9iBKqQ00qjrp4PEPU7lgsiHfnsUCt8OPGPTFMwkfPFsWx
M5BEFzgQ3aaYCYnvbcyIzlVBf5s5woRdl8P+2EGHjXP8P7ti25OfUnJVl0RAYh0K
kk/FvBCl082A304TMbilarlV3OHFnZVWsl1e/1qA9poZ1pntZhoVm8A8ph3QXCHE
UnSD0ZJZaQQuda4LeiL3hDW9zV69HWVrqcBvG9rCyzP6/hn5DHkDsne5gFh65XZg
AtYRq+8+mvb6GqboxqqTW5KhJVTXt3mSIOVJAqRVy7BOBR74JBUq0CIfF3dFH2fF
r2axJ6OtSVd2bwM8lMH2iONDVqajvvhZl03ZUuTBnCIhUhkFM0M3yQ+DBCJYz5Cf
oc2lG8Fp0KBOxsEUCULdyn69n/9cQa5LIleHayv1Tra2ie1+QBfNHCjhef1J8unR
Opq7PoyVjMZ8xKr4mWXElz0pE75VdmTph7fGzxEGAlg23GwAVvd456zYHmy5G6Kr
eKmO6Rxcf/qjcYMkFcd1K0dRzbsYlEkc6kwyUykHtWLtqbxex+npDKAAx5cqn/B5
M7XaId8DSHYGE+6x0DmxniYxhxegidvkXGKaqzLzzCAzZy+avQyifwyMKLppE//x
k3L535KBRLyKyznLmWDMdjfybcMR9MW7k5RqySCAXxH4UHNOVGPGSdrC0O/0LHEA
mAYR4XBsGagmNlT21Z5GFTjq5vDZ50ONO84cdIQHM38mjh689M4lPElXFEL/EY8e
yNqC/bUGjUak3B+D5MJBW7t7aZzLn91x673zZtO2DpVHj/wQnMWnUfA2ClFK2gSh
+B05/Vc9qFWYUfM3Pk6plOJaATRwdRQw5HmYJhul1de0G9FL8txpjbY/1/uJfM6r
b+z7yPffC8D4pUm78+Bk6qY+DlGbLFsdlHMTg1AVnaF8Bkg6yRi9gF0ayhntrmij
eLnUGylPWuwRe8ipj6cPW586O6edexEJ8KoZe1+Oj3zY8tUN93+0RGtlAKEByKDT
K37IUg6D+1FGBWF2EkznXkMae6EnLtvCRhavJ7pRRj0s/UnwIxKs1DRLw1iRS7JU
HnNRoVZx/xm+ghCFOe9uYmLx+ymUs8SUS+UeJISXhwqhWXG1N+FY+PV6M7JkRY+r
apijQwbNxCyaFSpiD1ESdM/e0Njr0J6j3xJdNjf2Mh2UtbkHu1VZOfs8uy1USWAZ
IVdtzTw/DwFwZtNghgeqXPdTKDYjC076vd6Mlk1bAmqAJ9X+zzKWJEk36I7kUkPH
89euxwTa+3deDVVsoXR+IbT93b1rJMQapxOIpos+1K8jkcp+X5BhBO7Le197wEky
kOVGWVRsFI9OXhyu0/kcTo4nYeG6TfFVCUWzaDjlSPF2tjPwZpz9b9sWz8E+6Oyy
apnJe0k0cidENsWWkgEwEUoYJe0yU5+rIpu7lYGlQKSP9XL3Mn7Rz8FtW7O1BuWS
LdwU3eeviQCWQUGQeUl3cGHAWGXYURj4olPSey7tMyvSR+Jckig+gSzAHfQRAcnn
7mF2glYXb2IPdp5GBqVsDNiKALP39vJ70aJDe/EtPmKowDFKphLgEjJAd/fCPRtB
bOiA5nnbXyEnvFhwofpnaY/2fcztOnWBNFeJ8W+NrzW37FnPK6UFgUxj3vJXlqE7
tPSyKJOotVkgK6wFB3Ge6yX8dOP/hwfwSvtJtRldPiDcu3WnSEiFYUwEEZ0KCY2b
Ydtl1CYO5fxRoQgCZSbX5DX3tFObENhl2YEol3OvobNB7IKEQ1ffLbfRt5roRI/f
dzQ3QMWmU9w1J0s4xJCNHWXAXqAs+zmQ5zrheImGn+Ztg3fSXb9rmLFAvqxlNms6
Vp3h0tsTH+zRZ2DexWIF3/ypUTPc1vUlksa7536+hN7mnjmhXn0EaavH+DUHlMHE
rZGCb/r3Yh+x7R7KrJoVKdO4g3M9UIVauJT4V1C9OWVAzePKU+NkXfP4LmL41W0V
qELOy8LTM8bX0TwEzrblO/7KHtdhU5ZWrchxVFupkFEIquYHkOu9dNRwCmmYljt0
vA6OKnMfzyAc/v/O8q1nKlj/u5NQxS7aaKf/5AELfeBNkYkB2RRkgA2F42VttFuK
RtHqtd7UsLnciVqB3iap3bCHvwQmrMVqtk0mKsfcPBiuCcblnQXTCL2C7nR4bslt
kMQzTXCXVbCHpb6zzK4jDZALSp+eYQ+L1nOmfoLBlKY2HlCrPUDPvabckNNrxbx7
tJX7unwL7cjxoFGMGc/0EFrg50EoLMB1hC+bAXmSqkukvRFf25b4+u6uNd0+zwtt
m8x6DmTo60AVfWCXpX0mbcNGqsl90d/RKQOUutVnEynLQ0Fs219EUzJiNcMUEj+u
Olhl7pxOV1z9a27jWm5fsJLOdKxCtDI2gs6tlSSuBx/n85qgr+dAP252x2ASzKDi
X0sUSR+sx9FGHWXVSQO2/zm6WFqbLUNtvW8E6XNGHea3LqIbuofgcNwyrzLHXsZn
AzIl5Dn8JCwoYgXzy1D5fvhOZXh0SOAl3s7al0B10asjqi8TwBIBdScXm7HdfhiP
n2EZS6u4N0q07DtYDrX2gIDaYyQOV7LzcS8//K1CBaHWRaYZITXDAKB/Urnwy9TK
LMLFgz4gXXN28nmFVLW0E62Lk7RcbQCoCHS4tyBIQhGVjlOk5cuMbg/vJ8aiwHFm
yij8eJRmA3n9FGkQPhWaa9wfgkpe1DL/egiKxf12oVea9MskWHs47S6Yg2bOAFfp
jQhAivPyC5CLo8PuIvvPVtvsa45Sd/oZBO2LfQXolFOV9O8SZM5p9YhubVT3rxp6
/6RuI0VGYRImZBuxLx7iqCPnIzXZvC6AUOVexYzwqgEn/Rg5u37FqET4NbPvz0EC
OF/iWAZ3rImpICt8NvJHDv6aUIakt+f/4XgdydQNYVZlOed3/eX6jEE+8k7p1yFQ
z2CsGlY6BpPdV9/wh0qwZfVvMbHtVugolQhLh6J0njiqx0U/4v10pzXm0tnTpAFQ
adgKwefcmqdxgQj61WxKdpgIoLXwroPs4HH2Tyc7b5Lb0L+Njrpi9tF6FTDv+ILU
GzLGguQwivBFjJE3eMTPtx5mu2z1+aBu79kd2LhxhGqKh0l7KTtmhpRYI/w/ynaZ
7s4bjevPBm16683p/ZHMfVMHsmvqRXFuQEcR/yqhD9olUlXOi8LUdW+/nyPyZz7M
+9B3FXOVTs9otkqT1h6u6PvsLY3tkcqpPZ9BFgugsZl7WJlhJZOpCMTulrrBX6qU
dY4BOi2ufqKpPVjeCexNBjf2lnb9H1beNI0Ey2M0t8wkYO/ilYErO0enXIWfC0uk
oAorjH2SD1fnoPj4vltjgQ4HycatS4g5GEtt7CZDfhafhQIj8xrnoQoTP075dgpE
0hTgb149REebcibGhOo92ekeI7SI8kx1FeYtfiR7wPDIM+zNyLLBIL2se+B87vd3
l7FSFOYjPtc5iBytcVvxUvaqbxFCSrqk43AovJSrUzLAccWERixRxfXAWEFHWwRL
YFnFhxEIzwEwcrvLTbRgDmMaAgmdugHDYAB82rdQM5Ik+6ZgiJahMT/5CeQFmaC7
Y24VRVymP0q1JuzaNPns+7SNnRmMzlXZaD0xntbnhMCLinP4o/v8Fj/5pEVGcadk
oy4HyiDpaE8G4ZPW+SXQkXgdJjoSzCKbakICcTSnKhLNmqgyayVwUHF1PKJDqhuP
BD2YzFJuNAopIwS2dew71Rq1roj4S+jwwp3BT2fGfI9qzApv4i7GYdX8SINoXPMZ
q4I6Hqj6Tx4+WdyDWmYcn5nK5xM6ZE+4ye/gqZQTK/i5eOaDNq7jFpPOiOyLXKuF
WuJkc8hguYUzD+GJFmKfy7XELhp9NrM46oWVnGNyRMbKj9arTuKPt3aZ7WKXzahL
+ACmimhrk42OyqCw0uxfGaojKwLShEs3gLYNqBrmpim8NM/5IiaTtvA3rL03thD2
X9jjOy95MAMhY2tUWwwyYJmnEljjoGJ7flS6kkeRrIp4SB0LZbCbu9TkLhnRGJjj
8YvVsqG5jfdgyWW6gAI/eEKyYSG11rqqEdFV/2R+JggFo0V6P3n+YhZiGjlNkV89
s/rFzOLh9qM7YuNuVdI7PM1w0a2EQzYiWN9y15q63ABtIeJrUzZHMYKRqupwxkt5
yfM+7dX2zT3quIQzSpfVb0dpqrrqD3cBI741JIKBU4G2ogeUEfF3fncA6PgTAq3G
c5a8wuWRsHPMHIpwhiH8XepFVRVYVf+gU3Sl2WE7lX1EZdy1KHnCPBNpNBM+MXYS
gEi5M+5EGLdF5VNaHpuc5BrMvbNpuO/1OI5JcsRJ9q9LXur0IzWFsfrAys09WZb0
Pkq58DPVrNzDbEbVzJDJnOGluxVCsLRG70HzDxm8js27CvM3AWydzQo+yBF6GXtw
UsXvlx7IaXjpnqU9hF3dwMxqUpMgrbTxi++9NSxGkjR6UhKc+xxomX/QSau8gS+7
s219mX9cJv2N4Eej6e8R/FxVFtoUmY6tEjctmUMZX9Gdl3pibfi2Z5cMlYVbrzET
6vumYF5CS/FMkffhoAZXr5HuiAEWQmoy1S6hrTo6rZh0HdHJ/AtgUnuDS/rQnjoJ
U2qDVvFw5ba1QIx1b1b3U/8IrLOYleMXcMZzPLYUlfR9FIO+JPdurZDPrum3yYlG
Qrir3RCX4kRJixialo8y78PiuEb3cfx/UbbDU16kVGsAsFTzKOej6pi3Q/pFXz2J
Npa9Y7xrjaB6hCWZJeZlkXu5Le84dVXghahosWCxmsZye+Q9bNmIem7Epr0rJu5d
JYzKrKUmExjoJB1jYxQGgHWE6tzAE7yktuE1ZNY4JdX+HXpZwDPWe87wgHcJSTWo
1aH5/zHe+w9olvifKhS3Mpo7oh2bzpIarGIFFaMHVJJWf7+8ZXMLqTObREww66ht
SyGeufaRkTjiXCTgOXOhHdkhTqvX5s3LQXKWSH/SE6vjRtMZ5FNQ/MMHEg/7ph5b
NyZOsB/39eM8rj7MMlnikvvBg9xbnH68FC3LiQiwY3f/6pb/ItyxW8Ew1TOL24Ys
pi2W+umYHrvlFdCJZmR+Yv1UlwSInHYiLF2DVsctHVzN1WoyuS6snzbKPejmMjjM
d+Pu6RziG9szmDwc6GW4dpOY4XJGeWw7c5C7nUUjOvX0m+uxuPFDuuprgscfpfW5
0bjrE+5PWHPL6JpgG7L1rJlbCMOYMOVSLe1zP4OBixB7+1mDhnMgB5exS66MWm2w
ioOmPOU6FSFwxmKkQ0bM1uVZkYhZ3Auq/M8dO1zxWIWok/iKZo4GTW6p+2ewO0MY
Agb4hzSlPdKq/O9noskGhn7zGHq0i95/CI7REd+EcWCUQ76CJxYpbCAOfpONFnQN
kLe3+2ID7+Hpgeqzqp2M2r75sdrfb5zl6YAlCgqxTBpNNQkCLQvWtAdGt5+XTvsd
eSPM16QXU5xnhGqIZTGOyjhODcCWDzrGMoLsVRFCKB1bUjhTUQ79zGdlueayNF5o
XWgC31823UJ1j+XZz+C8ghT+ED7lep8TKmbzcD05bhmHigBs6zyG2T9fYwSdUDNm
08gKHMTtqfz0pO/iS9mYGLo6mC7EskwQNcWLmX7OViNoYkIRMv2Crt4vA6i5cMk+
yFzb+Aocn7+l5IkyO2fHmSyA05dHcOOCoI2Fp1iC1lt4YEV9XuPpf6eQMawrIGly
gp2806XydgKcHToS1AXa1tnNP7X4z4ZBQ8Hr839JE5RI6u/CJneRyrJYMOQLrfF5
+pzrXTBfXLuaTnVXXKxFwGJ1e0jSqUrGM4scK7bL++12eO4NpPKb4bwnPWuGqhcQ
QSimg0AGH5vAvxGGSUklYftkV1DlT5xNFs3HFSmGY8wU6ydOmp9tq8/rjTeKDfyF
opth5TIqxLvaknpMjf8LE9BRjSgK7mz3TrRs8Dvl6idnj5yVL56QIBm+gJ2j6kWl
iwMPWCtVxlB2Yhbc6VKbSzGrSAljYNOSqVFoDsj/p52bMbFYWPegfv5ithyWrWEA
lPpSiFksYkDG1QgYBHJ/IMl7CO7UAIj2AZMKRBJ9Mq8kgWn+ATRvCJaRWFENtuyS
jxr7dBTuO67sa5l1Fl3aVcrxXnvZVP7tEouO1ISkX9zDyH9QNXiOqKQ661gMcer+
1tZQsXVadT3DiJbVCbur4VZokbg3UzEX0Fj9+7HY4i79R0zm7B2agq9FvI56Fy8v
UzORm3aSvyM2YTzs83uWgr52+4ruGkJYTDujald1T8YctI26K+EojXHj0/YbQ9VM
8orldkT9CFNiRN4mmCpAaIMNipFgoLzEH61F6bhp0uEmdLnIZjyJePXq29QIEJFK
GkE9iBJQkq27z6eLmChGgZG0HNRVcG1es1QBfvDjs5yM+BANv90IrMcIxsufe5JW
Mvj7iu1/n13Pbjf+PV5aZf1UuBU+PPPMyLSJ7JKZD44/V3QlOP5SCWTiR3ZKjpC9
r7iaVT7x5YxYxLr3gJxBIINX4Xsmu9/+VWInWm4PL+FV+aLB7Ozc9Y9SLXUPWPRj
4WU1BryzpC1Fl3DrE0Uk5blTbcuUt6J7xLS2hdr3cR7O4Oi76p74FcFQk6KGZnb8
CCIdx+Ljn3W8EqqMy1PSoOB2GJ5Y0pwXqyL83IJo2SxMyC9RjDUFD/aRQ4Tc1f/d
sNmZE4exp+LU0/fQ1K+oVGNJ+AEtMY0OoezqofmkiQQanD9Wp8HqXjVAszWRWizG
G14lAN6yyuQlj1cf1kNiyO/5SqG6n2cJKrYxzyI6hYda+GU8XoPRYHCpiR+4csUj
480XFTU0UQJJmf3yJGVox/Jx4fFrziG7E9FeehJdF9pXa9vjP6nMxpOTfoUl3o5R
gBwGCQno11m5CLZjcE8mtDKzn/HTi9ulvHaRbHdOjwPwqZ57hJXTEtXhleFLEvsz
jtx75kDANN9iZKPz4bywAKETXrnzTmV+4X2nBBUPD5S0NWMHy/SH28hq1425z/qm
iIUzB80+Kh/OED+dB302WE5RjpYOaxm2RuXVO3Sf4939yDJaR8J1VwHSVe/EnCPs
IuuyYoRL4RqvH6Y69G4juukj/NxdGJHDO04ALxQRaSPSoc3wnYrLZBQnO5+SKwgo
xbSzWLAhcyyLiV07Qdo/JXiEKwE0uPbkPbeS2EBPvbMWhPRFxbJXtCHmgUkJyoXv
Wxjt4TYppyHe6fMuLYJ7x97Fef7xE9t5eVy1lb6ShQG4giIN14rH30pALGWpEPc0
4f1X0zsstEIGahm2ftvr8ZyBFM7I94RTb3fXUzLVAIZM8PwLQikrDfnqWsxia066
Osev52zRRS0u06MjSkRxGNSJY62dNeet+R4cmClMsGcNHZoYiETvdOjUexk2Ya2F
fuJI4YCpf7E8FM/etuL2Hmd63bC6q2Tfm9rDIGZk/Th2q8VdFEgsNHouA/NvVZOy
XyqULFUZ1JwiUIOL1vGA5WCOyCfRJnbU71hUUlPnUFOaw/3UQsWdCjqma4BdOhJL
Li10f1VUtIztfllXONIFeu+BGk3pg7Hvq3CBrLKUolqbgKs3of47w4G/px+eF3do
VcxmwRHj2YTgra1Y3zHXB57F/o+KShfk/J/fRblZHrZRJWSZCUwh+TMsWZfxImE0
YrdT/vbsEgIbLMzgODKtbkfZBkrOFA1TUdwCH+EEszG4wqGOQadBRIF2ZY5kVCLC
Krtq7Skg4GLjLEN2uan4xqJrdUpKX0RfaLbZ8ys9B2GhUElV2w1E7cHrHbTQkM0P
lwWqkAvi6tZ7oshJHIh/CisY0pYMqjg97NYoldKM6INWwyiZt+zrzwn3ck1VCu20
IBVzmSvg2RYlGBrsmUtReWl23rXdswHDYOCSKvJckom/h65AoCHrHT5DGBmuHhiV
eIWM8gXpO+3RpqlOFBQvV8NJ1deS2ucDixQNyciTzyhwwp52x4ufD+8Zmbzouid2
VYE3dqUzg5i7NvlcBUyWXd4/PUCmo4CZx8SuKLq9nDj8Jp+tQw7hwG9ktIisH/Sv
6iJ+B/eNdyJFYiAx7pthe1p5E/77yE4enRqofxG0KHUstNvNu3Y5Wh3r34xCG7dZ
QxlxPOkNZEW55KU5AQblpUnxclmmpxMMAQ+EbCjn96hY1e9av+IpCLZ9sIjWBrMZ
JLEj4LcBvovbddP5mZoR/RebICsXxUzCkDWUaxLJCSo5TTy+Nf/qK/YFiJc8JT1h
kB9doB0KA/4HLnyWEqn34fTuvhYHrJu04YOVSBqTwB/vP7/1Fy5YobHgqSNEvfvB
VRTIy5ebpd/V9AJazkwGfkV5N5xJAf15y/trqHouaWSg0/N0Lkuj9LgLgb6oX7z3
LCbymiVtE8SFNo/630StE0qwfFN9+KjKApiEXJg1dpOq22fZrYy4oIhnNPluPR+K
UgSIsKfvMHmRBNtkUSZLCRKFCIXghg7s1NOtZqATsj2scKDbDusSYLY0+HL2Zy5L
KEYUVlAMKJOettOi3uDJdSlvMn0eX6JnuW/f/SkF3uXBP1S0Wl0gQeXV/+5iCMd5
4RbdwK/9VTgB6QXXa1oFOyg4f2DtAPJCva3qkYLlxND7bF5sVNh11f7YPHTuwVyn
BvjwRT2KOlWdNZumjvukxXaijxWvMapAOlb1tsHMROx56WkTinnvho/S8+3eBcPO
c52Ue3/4uwCR4kU5TNQOjWgjSApkBzwK3NdH0x9I3/3JDCva4yg9wxl5/jkAGcOX
067czfnpA/YTZRfiLFEKv+oN8zyYWlGXlyqcW5C3hj/1bVCrsBJpGWEUD61AIAWo
OCj4yg+5MhR5w9VYvrQwSusqRk1OmwWFIP65eNyDdw59lx6Eqjk+dHM3HCNGzFoJ
/wRTqKyL4lrYjlBSIqD+EbIbFtuzp3ibbVGhgxwi5xquNlHEWDL48RJQx2D50iyy
+ra5XZh/8QbqEsplZspwp5oM96dLEKnLTPAZTAX8j3cyqiiZw0cuBaQpK2xQH1Hd
vA3W/lAR1nBQTgW5dla+FRUOYHuFQ9nE7D2zJbyHBpGIN02SO9FGEItrE5agq4Rb
HCGSpyOZJYm61Vo/LtGHlY6ORZsL+YysP3qgiC/tnO0gcFwI9uiAPUEx6qISWalS
YaxStQI9/1MELGANTIRal4HDvwWBujMal2TUKbX8TA9/Xr6h3fiupNeJIyRViGjd
eKocrDtkjLwA14AyvR3VuXL8nUOeJLgy8RXEBlJ9mNyCUdxpwaAk5DzqMR+1hbL5
waHy2713AGMOkO8Dp/erXVUjY5vbeLNV0e4q4Q9Ow9BgNl95oDmzQvRj2QhtBeus
vlh0h/twbb2GbaBOA6O6yJL+rN8TDxOlyKh3DtR8LppRhEB1/L1shp/LPzHth50R
6jEg6J+7ewRMeqo6mbgXgTU19te5iobEL6u5lNMCtAVY3tPNgo1oxYj10KtMzgTl
zbd8NAFfuU3YPhFaea/JJ6Ukwje9eNBnzApgEyf1mO4bj2tkOYM32h64wSpTKN24
05rsJVyuwZRotTSQpIBMmuujOu49aX0jSPYIV3qrEHn3XhErgkPm/y+9xWDPU/Uz
m7JzNJWMgX+MSk+iP3Lc0tuP/HelgWlnHoYUuNl+EDFustfis695L7Pj/IeWNoFa
ln6g/D57iNPEhnsZlx6+Ritu7RN7A8PHo4A8iSZU2iwLcBYn+mKSDUowzpY2KeLd
9VfsLAQMBzM7ym5haKNBzZVNxhvKOcmdRV3ZGOiIy7YFMSNx35mkLltYOXpgdnyN
rc40S9RM2YjMgDfRJRMyrXdEcijgyngQeD67MdXEm9WsKH4w1cg/VHI/dJzgWf9s
SCysoWibq/n4pez7uAs8fO3SNt4x/GDgfGS29jo5mAKM9PjqBN8Tb8KrkovpXfSu
zYua2CR8AIFtimRMDf/CuhhbIElsewtVSvZPlOsua994FMyDq+1XdtNTPAaei3zM
dZ7DTEy3XnPY0U8yEAK1yN2i2HINjJHZAlvXD9KYQ4QuTbTnmK9qa8EYU6lCxyGG
MvP++ubpg0Q0kD36VNUHDneAg/btvZXHvSE3jeH4q2lZ1kLT/0WpXefbgi7L3AWE
2IEG9U/eEYWioPLEYh0Ia+bfGlU9JnaoCHJQsqHcFGDPFQAswNDhyFHa5ZSsLPZP
hEVfVr1h3KIJhM9jMktr8dn4TMfZnUwv/ZrftxoHTRr7vKSRWyvEWX0OG2XDC3kK
RORkrrSy4Jq0HCGFrDRz3yuraqpikh6IqpmANMUyDgAtczPbrT+lFyktSvBglJDU
PAtRzYm63CzXd13S435+AcatezyVbt9XuEbpiWomiY1GW05D6w78HctQ1788M/iR
rL2DRbqPsvDsyctlMj8PlmObSrpEccXaiZFIfd3Cn+0gtsdipu79ZkjE8Hc9ccO7
uFd7ANso7hgqCFHVwzMx44cyJBosmDucbU1g+1lOVyprxBM1KwUOCSOxRXDR1O9y
X89kMvgYFszFdjtItTJrgZ646ofP5MNfXc1jXIE58Sdy9izLknSWbobCFFotN+X2
QJ0H+XRRH0EG1a5/VJ9jALYzgg5hWXaYu+8u8QIiBBtEXVVFpfO8rm60owwpf5Qe
kpjYzZduP7OAhIhp79h7FaQGhulVVDetuErtovJym7yj5GTDic6fVLPOO0cQrw1S
ogwuF2ZPJEQR3tK10PqKtKNow+GLYKVWGpgBp/CqKaFlpRr+/XKFzrdRGJq32ppY
gxsuY/fTXgfuf6t8VaTiBYT3Jsrw30QPKD0iXaCXwNOiiYyQlGCwog3XwDxZ1FOm
SzBtq0ZLg7r3hcJRWn0vgb35E3tp9kZmKhXkXtr2tKaOG3hgb5iEJpfgM8cHwyme
4HVysJ3J/V4Ypu4ozwuLxeDuZ+OY7Fi3Kg8m9pKHhbG5/Z5tLHy1N8IBNopYBXgB
XKTM8UqU8T8TXj5Iv/+8t4D4lFTpKD/z1MI4KQtLFUfNstRP67lZ9z2g/23cBz8E
GQg59v5cDffzu5NTOVTgfMiO2Lphr03LS/C9woqAUla0yQ0X8acKrxvpKyVHzmpb
iIQjIsDCO1TkGAQVSg4ph3bJlV/uEBNz/xpOVyAvd9ZnFjf0E1KtwtqZzZ75WqYA
eQOwO0qavfgdN3Ev7ZrlDx7tW8eXFmdFooXToMspYmUsQ8JNr4uVV1kgoBiIdat8
mykD0OfdhYhmJHdC7HTxf/+bSBjl2f5JIN2peLe9/AByRuQVFPQKXvC7QpPKJQ9J
hQYtI9XuMq0CN9uClEsmfpl7V8UWtjSH3gQ95H7Gpck0Ba2H77S2iHSCG59LSgnV
blkCEdvmBGbJ1BFAJ1wKXnjHe8pAoshTIF8j3f0G/L0eIWdUiTWadPOq5X1rFLE6
Sblpd7415Q3/m46V2BHmKZ4ObLye8zs+qT3KotMdpoK6fJHVhNARHHXf6IU1MJ0I
P3Z+pOHzW8VPFqwIIhrjbtcRCmmfrYos8IfFdXkAwO4co9LPDKnGqYeZui3JV4yr
g2t7X+jKMME2kHicBCJLhoh35q31z0Wr8iXyEirwtC9FMTH1B+r5PzDJO5nW09b/
OD1QrBHODhDzzOM7vve6vefuhNgRQhK1md9Q0OIQ+lDyvVXFXDj4rQ63THPSi4Iw
GJ3LMGQgkwy2XCnXC55LLbB2kLoj2GVjuUmIdcU7TMPpQz5TbLc4htibeiQm/1ur
333w/AozkazpOteaKDrBkeYLkZBFE4UKFYPvpCEje4sHNiEneaHEymA95S1QTWmt
dFGEuHkDOhDv9VJugQR2x+DNK4yf9JCf4yNfFzdRB7VGunQ+m9xTs0lr/zlPHiyw
B6HFkkNxKYjMD89AB+Glr4GjQjgxYVR17ljMav1Mcsk6ME0dkcxC3IFnixG/meDb
UOs/jSgtbEy0QhY90xtvXv0hlCW7qsfGMXUfSWRzBCBTy4U8cv0jODMfMDP64/Yx
TYnamKoVTep4KNul54Vvdf1aQzSNPevIQQamyy1kl+obZ5Z6kABCgxNupUACvnmC
I+7dBSxKYbfjeCl1g9tWY4iCLqnVXrs+x3ndaR72IVdG5czl57u28iYtD5tYZac3
QBu0oij8U4Y2WsvauQY2cUINdtHrK/cS4Fy5qDcaLYj5Oh9/Isps0B0g2pMkR/Jg
s3i1Wo+7niTJHvWHYf9YKRWOplA7DOzy9IStxKhxHqIU+5BnmNb6Y0RrgUj2nKhL
+7eJo+J0IcAdPJnWnbr4j7Q1gNdc0i2v08JlDqGl4Bg/oUIGMPTL5DyDN1lFos0T
BCcxYkVlUqwlz27zsqWOfnCqTRkY6pwN+IxVudKZyS09sBTy4qRNBj4FW06EP1FR
n41iVgX5ognnQlnYsUL4kiN3H7byFcwBk4WKz5/LaFap4oFyWMuxaMRtCtlUppAT
eOBRc8k3dNLb3NcKmQB9uB4NOVKgeN0iPdj/AdbpENDnGvK/0icM5EkjEmb4OrLp
o9JsViNx7qMd59uFJ9yOYcIdz+39cW039XI7hOGLngWxem8EqkOIgR/F1YAomR5f
V+1+Bp9VKAX9gpP4bhjxxqmlEWKmXZSj2WcMqgUm/43bb6xDbkOzAaavIfkHOCZF
IuX/uUdkdJcamDgLa/jrAwQpGxoL+fnSm1DvwHYWT5N2xIQbKlpmmy2WSjNSguEi
kBwgQUNqM/jrfbqMvTTI23yFGjrl1qsBCrmS8obJ2XbvRnbbgNRYBb+idlRUiVvx
nFliIKtlFT02Qw5KfHxHGPPueAsjupwbXvTsXX6RRxwstvUh+/LH0YUZXvxTAukd
ZIu3Ag7HXvrHawu6eiFbAV+38xo/+4v8O5dCihZSqAkfzuB4EAKk5YfHiZdIGm3w
K8ze4nIvGroqmO3gT46lK58DVbduRK3uDC5K/V0As5SJnHn6A+aVdfUKDcZ92vxR
eFN1daPB/v0KeBHJ1gApY0EcS5cPMhkANiPHT5dMt1Oclg/zFWvl5yEQDQUg7c4t
8btkWHkKDsAeDpNAFaeg/TYm6ugLQcy5QGgiYh7GSX3HhNJ1rRABNjR4AiwBOZta
iHA9+7XqC5ojEJCVclePsiXbjPtNt0tSXXlo5C3slKl7/Qf61RgnsFV3aFbb+yrM
hRAA/xS9T062KUOrTvxTGM5JwKI1ufkvFweCsg0TH6Sp/xAHJY9UhIkE+2/+GSQQ
Opu52qLVTXPeo0KKNY82A2ZYFq1m2T3baVa0Y6ggxsdE9IGTWcexDhlOSEDv6MUX
k0FXETzPybJH7vTxOqegVpNfQx0FRzYHVwqr1eNAZx4GLef1Fl2Z3Kv2wCKnAL3n
Jtxp5cSvnAqVyqb0O5ABirqtO4GxE0Of5ZB68b316KXvcjK8jR6DUQ47YuBqNpAu
m3gGt8OK7gaHLQfR+zLDnJzSwEdTYU21rRbEwIgoI2qlQKzIoYKeHS51sOsFH5Mf
GaBV3daqoCWGfyxH5IUxotKqEz2zKT5A2CunSVAXtjnjhvpjqtnID+inVqsLt/q8
D92170siurHxez29xOweg31jGqd/oX8njMF8U1f/h1ovYD9IPnt6/rCXGcptT5f0
1UzJ4f8wZHdiHfua6Oca4A9/hnk4gMc1PVHiBpO4QRdjwtppVPu3ON+YybojzkUP
UWTfVkaE287Y5/WlVt4jaZFFtE8UAyThdXFNXhUu7ViVC5Vkn/vuFqlCaNFGEnO4
kQ4zOVNHCITl/F4jTgyonJkokpiQKR1OFIE1M04j3Wrlp8w8VkYzlBZG2Jdg3/SV
kgwWABuNc4DFvySCjPz9Axc8nB7X+Dpq841daSmy+niPlmUDKuVPPxqxAxef4tHa
WgC2lpSvQnqOXeW6n3RvwXqtz5YuxQe636zxQvnv4c0010iaCwSuyJJa/2FAWHJJ
NGERfgaiARo9FXJqrZkrBrLzznV7BbiSUWx1r4KKQ1vr5SQkfmyEoCt6O6Ej1g91
cjqK1ckinMpQ+hBWkBMkJOJCMnf2bFf4Gyj+KYr+4s9bU4d0LYgsFJiUQjwS2FMC
8edb1gDGuJGZVy5dL3RwVPF8xWH4VGvCRBTbg8H1iecN4f0xb7M1uCPwLE9HuI1k
NfmPpv3HXGkPDBDF5F3Cpc9EAAzjvRrfEPfVaDKKb9D4N/bhd2ya0s6gcuiKxPIx
P56QfmySm5af0Hae5MhqN5eURUgz7bcIj3TTXRREng7jZVFl45GfL/AHyNxLazN4
N4gb5CZGsMO5+oiqFStJ+jfqZL1hxBgbW4BSIjixAqMtO9t3aMCU860eePGeZAUu
xxu7Xj1paSjl4zLNSIPFCkGTfG3B09OYP0o5YEh7B0JuTqV2iDsF474LFL99cVKw
Nc2tqksdwlmcabYf2XNR/Jccg79wZ9nbefk9/QWHJwJFNwXHf27O8kZP2rrDYuP/
tMoDM2o0pat5INJ8LOdYvMP4KUsVMhDY4oexUzh5DZAvqoSTb3Yt/7J5eGu1epJn
fT3dv1DhHN87imBbxGzfJDAffJaxRxL7O3VGrOCuOZq394SWeScimKhLbqBg73Bc
rjp0DMHxDF0XjYJStivarhuaGBZjiM1TwqdUyO0VLeoNtYaKHootVEo+7OsQ2Nft
weVjeZUK/n62ghE8+8tFmolOUoeH1zZ2EgyAXaGE8l+1LTmE+SvY5xikVO7FFuSv
+vs9VdrzXNxelqh4UhaeNatChqOi2rIkhl0/k0tQ1E+y6l9QWIyqHNcZ7fccSFpt
a8KqZ9AUAc+2VI85QrfoGNnTHBmyVBjiycpdfB4UJ3xABVmUY3w7R5jsb+qYtSB7
Po3nSlDadn9l0yqbB5yARhxxz+KhH6WXe65/dKiosvbam8Df7ga2iyNCoS90V1Qh
jw/mLi+srseERdwTmk6UWzgOfprz8mhdKhN+WlnueMfDrR/Z4UhVgjfbNhoP5pjX
l9Ca0lQFepKZzJVZPyQNO63ZoAGQmEKYu0PE7xV30OK1sNkJfeFlbvZXzMSxLw0K
k3BB7mcer9eMZdwWGrRYrwgStBNDOAV2O7Wnl2ix9LR69eDgDCW3knvnNrKJPin2
2m3GcoG3ZTf9WylDvrAI2YISgbRfqN9b8sFSsxJyemURL+Rl1/3DzsN9hNZYu9Et
zaQ8X9HDB8LsVwrQf6Lj4gwEAP0qWuOI7ZDedHO0oT1bK1sF+MWkHcGPLyuBbcG4
atskm2cZz07cfNJtReKqa2b80m49P5cvn8cLkwgEA4fDIT93KjhIV4+2a0Q1PTed
81Z8+SiVD+AAWliS8M3/ZmKGWB+HSAZaFfkAXgeyRRnx/vDqu+LCLgBdGaM/D6ux
7+z+jrVHmXpNP4Ad92skaQpy31szW5kgsNvkHXETasMyaqYt/x4nDaD1aAu8OOC0
l9t37umOkNzVHKt9Gs2a7u6y1HbQPLpZrnUQVUqQp5aOcZni+Vyw2W6AolfHQk+p
qbiWsFKYm06YJTYwbAmoH4qw60FA0/GcNvMyA2YkidQaHubneP/bGrs2NkS1asWa
QkLkB/6TVyDCI5lMgMcR6urOX9ymz5hdw8BpGBNkrD8uJe75qC1V8o87ygA+KrIa
V2/pk+EomcvlgqR7wkQGASil3n/rcjgYu4mWhF3u0Say/L3+KpXUf/uqBtg6cFWQ
uB+DxK8OGu4wmYQEtue9zABPHGNmkAnKbgQdDZNzzqMx1qT1yYQk9Xji/HN4DDCx
VuAZTbI7G+/liylcJmKHkYuy/+7Xr5qMwblpkjg0Ex+LNcFG3U7VkjWhcH7Tnq5u
Qs60yj1JmPp3MgdMWuOM2Rb5rirEMvI/8eQZMKI2abu++ybqYDxfhSii0nN5hNkS
orOCgPyiOIZrNlMEvSNohU6zAxvAA1gvBx5SsNXwlFzolGAOqL7SltEmn1KoRpKv
sZFYtpuTZrvY7MZ0kf6J3Wm2KbyoIf3rnL8WkZRSH9UBo02H+LUf+6adqRsERUVS
4oICkl8nn9NCthnQAXT4geOQrasN4LeZa+zAECdXYzC1DpcyuPwAVHGeIK9EvPCf
+MEkGTE7pVdmYI5eN0tK/7hanHFrWi5169etN9T55JbDERb9I+trBHpU2iOXPeso
rk2abR2WggugfDrgx0XDN9NZDcnUNbBC3QR5RvxdAl/dZhruqJmuDC2xe3QuGHzC
RTBCrAdm1vXdrxHQqwRKMztKGR1gMpUGjGFJiCCe7C1S/sc7UBmr2lkzJGjrfaZl
Q1KBZ9iRX86yba3sbgvHNRUvnE55XKFnk8xiUHrUEJSjpM17nWBY6D9bRyIi+5sK
4pff0JlPGbxocNKPbtRU8NjoC0x9MQUCnL8SjJa7sk7E1givWLUEVy2P8nCIB7ko
VKQCZM+09CVptLdISvbI9JS3D4yXR10dy0MGUPG2MgviXsQrUfiQchYcJcKs3irf
9IwDfsz3ug39YxnjBGnlxRoEVqWA2pGkud8oE3GZFWU3KIrDiRfJ25QXLFBHjJEi
jhuMrPV8wSInpKNi15TVpo7VyMeA2WEhB8UrJ6La9RfZq3ZM+1W6QqR7xFMnvRwb
8hLS7w/HvQzAmhDHaQaxuxwJfD8mPXAx0UIYMH5HhRsmRn9ZG0MAh6OT6Gq1j2/Y
vR8idv9q0kuI/lopWXzOKyUc2JAGCVGWBqhNtV9v3LCHrZjS1dXfH8frpFh3BeGI
j7GjFa+gFRaWsLa/er/tsqVl9ZhJRZVcy2KQtY55CvWghYhQNsAkONu0XrPE+EUw
oxHt8KPYWUUoqv57v45UWYOjUHCGWklFxEXV52bBjuc7EtgDzT+K3CHfwvvVTMQN
LQbXc0WIrwe9Z933rgYlKNwBuS4HFpQk5rU7Pfbzi9GCb77gQk8hhgpoPfPkHgjg
lld1Q+Yhr2YMedAhe4Ya35/QAjViT9k3BxibKIPl+rHoCwZspxdhWCPMImhOeW/0
12ip+qJ2P+Dla0Xon4ie4H06hl4LqSeAcxUq9K3YLxpNmKn0tBVeu4AUe+/pfUgi
LAfRmbsJskmGyKkYjd+qgecVlKu3nFOJL5bMzhP9d9jskGH+Zl+z3dPSnGQCGS3S
plP0VeOj8gM75N5Ls6IWqOBaGT7RaFJkvxs3vJfiFn9VLYoK/lJTbQFiaG1Y931i
9tD/RimpF+Fj20ynCEnqvXGzzv6xZoTBl+ew+vrY7kD8i/VIFEzZqGYUuDbHbwAV
P5HFD6khUFJaq7tZHvmvDGq4BAmsamxzt21nE1pbMGNlzwCfMyTDBVL8/kqXW3RT
QezWZvUhcF6b2HNbkCSGf/nGV3/mi70+Ew0eztwdSCvrNI6DRAY0zFZIQscUeH57
SXnsi5pYaRj88egLElBDE+Uyy7VpB+wYUNrR5PqycpG7kruC1rguuDL0L/5dDKXM
7p+k98PMzzA4YcUWWtyz/jT4OSxFTV46WKejrRqvYXqdvPo9EHjt7yL08OBLvW7B
r++rKNc7Onjl8hdu6ISh+Acggckx8uV3k/QKwTwM1tSEWPMHSY7y/u6ljSG/0J4l
ATznXS+TyBWrhd63kVeZUiFT3bxKyb6XHCBhTX6FeER5TqwrnmbqbgGtNLHlCJs3
vHAU9GTXhGFgyKKxFKLtTMPBnSmK2USfxoo46AkDljoB9UHQy+TWRHAqsRKCChDB
nDxZ+VY5B7+d5sHtEolrNT6Ykr4FDPiD47hLszbADDA66MYeiQh0xPmv4R8hFy26
FMGU9huSpoVKtY/taxNG4evl3+u3Ar84a/wWwih4LzkJmSo8gBA6Qvq4DBSs4YIn
PdorF4Z2AnxDn5poNR8GDDC0yoY2vRsrJTKlJaIuOVR4lPgJ+XZX3Y/oih6g5We3
ygMWgfzta834V0zpvOA2XUDUeCafagZPibRWhLeWaFR8zGUkCsupaySyy8unzzHB
6bNmqSISWKgnHZ6UKNQFVX4FfFtbw1t2xJGbKYeqZyRORukCZ276ZPGpcQ/a/7mp
GWztb54RVZxjA+4WiVcYrADuaGLmJjztnrVKdbeifyJpRo/RsmLUrbfMwkH6CrEN
mO5kH+I3hYgYIoEgRCrnqFt+hzYFBHt2ChRWQTrur6CUiaDyAuGDKsGAfAIneCGb
z+RSPcrzeaxYnUstBfX6b4o9Bh/FDQSUyl1vhKux4WlyswDAt5U6LVIPBFJucx7C
jsv4RGJ0mRBUdJac0QIG+zqf1W1LzrboHmPbPKXSZyGt0xGPi7eXWzTqlxOkVPAj
5f9isr2GnKH/C+2FQeNs1A3LR2quf4NJmLgnoUTlJl8KGgiS3MBuuzeKY0yZoxki
K7VU3moioHH5kawkYGyWz/Usz1aUZSd59ya+Z+H58zjKXdL6D7xZIXdfP8hlyDVN
4Q9FUIkGlFFmU/R82ytJLoW1Etr+jqhqLM6peW9BiVmEfCfl8+dGYXKOTYlcMk3b
XuVCEMRbThHmLbJRI0JCgq0uRcgxKS6FA9QWCmP/bwE3RGiC5l0fexSBwE0g3GCH
A8J0oWdsCZXwhQNHx9IarGouq1IXbLHCZbG+1z6E3b+x3uOAUlXVtZQUplxffux1
+KH8geuxbjEt1uVLAUWrAYaj6Tag4bEArfkUZtJeKoMAHQyY/nB/r0TT2soj/hBb
bCuGrOygQR+B9KnAsZQELZKZho12DwQENQGfQMZrk6IWqFqH8jaD89G8IRpktRLQ
wwBGxHsEfPqWhfpnEeP+PkTGU8mDwF+BNQqu4szoy1CGzwK/HbT4Au/Dq/AXeCIW
xqbg8jTaPFGrQD9oKNARtiGBkMt7FzOjUL5aiMv9fLEbsnJYngiLwKlY97UPn2nj
RF7sfvAJdYm8Y3Zx28mVqM+LNNYQFfqmD5hyCGdyBxsHjwr0t4Oocm5IhQypDGMT
qY7vSgNFk03XzCTw07iDYRwvJprRe6Tv13BJXRsHF/iHoVWgIbVjH1yRBivVNlJP
s40yNhg3CTLxP4dSNEQSs10KkXMjLzoyZLbhAC+qIw8HCNjnBsCkl5ufhQw6DwE9
d2wJVNLtjGRhFTm9ntEehpTSNl7U5suak9FrSW1EU3ZH6aNrOHLjqdMoZAF3pMM0
drMk9ZGCaNzLsV8lmaAM5OQUkP0cHXfe/KcmKyQRvgDDtVrCylMrmfkB+mp9F4Lg
WbXoZe8HyCbmCwTCdu8mZPeWaDXYyn1fIJblDrc3dOmeaYbyyRd5f66QLqkUJv42
MdPRLr48lSYg/8/xY7nprOc2go1RZnrotc6ZaClEeg5t3RcxZR/hcRTDcHbDEZed
oIlZ7h+tTfbexuEPC5l8wGrMNGRKCkxc7FTnGcClIwtbzfILRiVe/b9CRKoMmgEr
SxLJczH/AtJO5iEF0XUG5C4zxRDvJZ0LwPZEz0LIVmY+v/V7/uR0qQZA9qKbot3N
RnRBNtgEO/OiGFxERSCOSZYHPv6a0vyZNDMlxERSCm+XRb8n/ce2GquDcBddyloQ
myJzQj0xe3YM5FhDs3d/daALxlJPQkjGY2CCcI94sQk877t2FakirWGdyCmFgDp7
WcD68tY3QvVbnHAL6l3WSO4XzVttVVzWa4LBtU3ga4KUDMec52CMnI3JRc8pjjFZ
7mE74PP8ge1+HrKOPQmplrdx6p0xEbkbUvHne7bDAxw4Y9AsLzkIHWbF1BD9E6tq
rbsNoRjXCChmYYF9mj/he3Pe+Y8zuFZ/4zGyJrlfVB/77yBhsuiCFUXhQqo8pPM6
7KNYpAq45GoK3cUQPGZB17/0hSKp03trtYaUAoqRAeWLZuV1nTw4lZSl/coZ1gBq
WqT0IKoM8H16/q/dFp1YXPYrFqCtnsyq0r084uReKwl7UFTbDmac2T2GhhqtChy8
zgSDBmJF8dYt0cUDridmRNaHIQcBxH6vaGjugHJChej0XF032TbORNBQfPjxq3V8
Uss1h2zzqF22fJvUJme2EbJKvVfKfLkJyHkGZB1S7vSkJ2Rda3VKonywHd2/Y0L/
4guBySBQI0tg32wYpdf2gKCHaXqfqMWq7QPGrBr//SHCmHZraDMudOOkOR4e/NS+
MoRj4vktqiziaFfUwuqg+1KmyZcYMz2wcXW7S3mTBM7oARk5QqTpd2kRELDQYd7R
HCLKMDHNbGu/TYS83qdgyheTsBSO4H8sjosH9Cvw8gZ6ixFA1GMEsi0tX8IaCp5u
Jrf8BJZ8dYNXU1abJ0PV3fVRMhUOJ1xev6gexxmFjzXkPTgdB61g0KPI0rpMjnCc
VHeGsrLbwW/Jd6vXqyy7742stPF5GmINEOUimJnS12PBKpPTiXnoHExURnByagYE
/6yrt5A+9LzeT/ncz8fDtvdgL2AWXM5Sp4T87R8Yg+7hkig/CrOqDu0GXSJY36k5
jK303gD73QQ5CYQa9BbvqZGd/VqXp4gl9haoYYUMTp1mSE+mkWmQrCln+dYv6W6i
XZjR3yr5OkJAWb4J50N+u30N64dLDDErV/4G+yMV6tSR1DhuK7fCKYtO96oDPGCc
okuxnfw5P0Brd5ApphtpveishZKm+hakk9Im/R6J7UJTuS4KpcsTJRT9ObrfJL/E
HD7TD+5+oCdg60dl+g7v9iUZmByahVpuUV3fcGXWkZSLWGefMYOudO/BbYji8mmS
VZ47JBfjcXQ9Z7SlTfpmwCpMu7fWbn8zJHNjDRwoOtvr1cfRH/q5tK9nzYKvXr1Q
G2UFVB4evErdrCoonJ9gzcLBeROmROhxjwat/I9gzsLXQIXYrM7Su1yDFsyQU2Mr
XDiM1g3mzqIXWR3GUV+xx+LqYrXPu6ZGqrX6NRhDJ6HNejR5C9/lxo/4yzZ3fapx
TheiRLdYClW2Ekhxi76U9dSHsmlQaYtOloARfsfXDZ8XyOigu3NMONvSay3FhtEB
4kO/rPt9u690shDgv9O3ABIknk2YNbo/aYYD0gFHGzEWt0cAazeDms9iLnjOj5ki
DkRo0XhFIBt2Si2ec1wattU0xbD9IFnfcpPKpsXJcIAFAh4ot6rMeInsWMRB5P6C
ZF96V0njoUv441BbfHKgPTs8sjDYlIN6/0fWT2MmpZ7UYewi9FWdZG4RZigStysq
QBRj09K79rNjLYn3R6U5gom7WSLpXmfhnLLOuE3m9+iaHjdYJ83gB1ED24bP39pX
so70yBtJ9BK9RnqzMyDrYHyOad1kRDYXjMo7SH69J6s6nwJYF/WEfpqBfYTmw0uC
1XJ6n6plygGXP0HShYCO44QVQ4gqofLHADFkULpbyA2dtR/F8SglJDldSmvUGlB9
Oo0hJeoA8PGjZrDAwL22+V6MOHzG3g7KQZitHlBkO/dm/IJEsJvjDaI3qrtlnjUP
nQOSL72SDmDCBSmg/ZM9i6bASeDZCCaYqQyrd6JuR4WwMwkHkj+8ykOQoevAyUoB
dZPM9a6eqO/Q95znqTX2BArB7HgVH10DY+/oLpGEbOhWlb13ZjIePdUJqbBpULYo
fyvlq/2vjxRRZLVU9Y4Mr4oX9k5T2TU8ueF0BfCfUUXEg9N0bXH+kNUhGPszGWBP
6THv8gmHlz7Dj+UFuZqvRoZ8MSw+mdiv8NZQpJOi621/86pYrX19DsPV23BsYVUL
qTiQhE3uCLWWt7QhKVzg3rGMnYAUq1m7dHLLm4UdxcxeowS8ANTaafViDciy/Zhn
jwCBCqZBh76hxdLOqlOqEciEawKbwNadGlM36J2E/1vTUBrfnS4G2wezq4zJR1wZ
5sl1Zqju9sV9iiPsDcEuhQbwEGRynpEhxfN2LcwH3rOl+8OYUA02TCrI1V3jCxAM
nJpg7GkT9q58dHat/e0qhw5ctm78nodSELpoIm+gXIu8VCyKqdQQJLu6PDqzaCgK
n1Q3dDW1eRjXCOp64qDe5+m519EOrcPpt25x2MDFt15y53o18+g9wJmmzkmL/NKs
X/tGto7ST/VkKQk2EUnDK8XjbjI9ANvpyxZ1bDjO7AJGZACnnfAkdWWWmLMpmuob
Buhiw2/AMc1Ab7NkKUbjTwmkgP4mIY12pCbaf3FlGJuHXUMo1dzTpj99vEpIaqik
NOHjxpaKL+IiVy+ugobBnaXesdiaxk0fdk9EMwKDoQdOUqKTRgTF2VxAidqzrTDb
bAJ6VqP5VSYHCJOjDrclhSCP7GUv9rhQl1KNY0R2hzAPAtu/Y3CwAFHrQ0T+1do9
JHjuHQ2wLAySHDib64NVxugQo/GXwXZwPsblsSw86FSu/Mzv8Q3hf3DXKYXC6Enz
5Db9dY+5zXvh29py9V9plKAFjr3nZB8L+ffh+CQx5Z1pa+W08nFhNeCgnSebWVt8
6Vf7lZN4j9MrRw230HxdZqnHWCaVMcsnJ0/TFI+EK71t6rYKa4kCwtQ1N32shiAp
aP6P2xby/8wOd/3IYZ71kxOvUFGZRZg6B/e8tKpfiBtpsQAmYpWieTFR35lD464p
b2X6CtECd/mWUARmA/VBK1NsdxMfyDDKPg4ClJ1YsMA+AysPlsN5Z48v2cl9qzG1
IOfE18TafznU2J/VF9Rmcq9ZH5EJjNkG0zJkUgDzZKgOjmwQecICuUoIoTzxpQEe
unPjvaeKanXri7hbG+soZAOXlyeyuDWHIHokhWSF2KTTuBQhyBEg8Iw46p1UR6Yl
B9kOdbGGhsEXj4tnU8NxKSj3RHGDW2wYoAxrOjbx+Bi+VI05NGoovEbszYC7FKDV
in/xSQbi1UST3iYHsHxOcg+1dNiVJH1NCx20KubYTotU9y/sUbKYHe68/PYGBc8Y
S/H+ngcWTQgJKlEcjgTpbKstcbZi+2czi5or1t9jLzJsls7FQzIjGMt8ZJIVdFg7
zEFXks6Qgy2/rhqXjooEvzyFuE5/r7S0BGeWYdXBdr9FJZksHT8JdSZ/dW4+CYM9
7Z7/WglF4liUrHhFBY9y2T05TBxKQk9ipeygf7/IYlvgava1aDghGpLhxLmEXAOm
Axl15GPCRIJk9zk/kofAcWgKDuRZUmhPkcmlgdV/KsjZ3FdGs7046hdVfECVtIt9
i4H5xD3vVGxMkopF5XgxceBPEcIXMWe60u4+BUDwSNZyLgqmUZcxBN9LcdEGlTfh
5FgVXyLf2mdZrlTB5fQDsjxA3SbMvwOT7DXZvKi3Oct+vmV/EPNF99I+LiKwpsPh
71kw6Dva4cZCA+gHoV10gYKGOn39z7Vi/gLq64j4zQL30W840qqLQl8SYVx6Xc3u
yucnWs0G1vJEhU/R7SrBQzCbN3bww2CfMUgKlfldoSzVUwSQuW0yBuAe7Mc6+15l
RsWZJjYAS9MorVandZlqpFTgRYAIiM+mewFFvgumEuJoBX1ap7/tNsaDheRky5UA
raUk98Hk5Om0t5roFgD4n0wlGPoZSzoj0d9sUpWcpebb1/KDHWG9Z0aoWr/Nm7u0
xShrDtJJjioqEGkvbh61AV2AdEch7vKrRCTw1US0VVVv5N+RUpPRY7rkk4ORJw4O
NDiNN/Md/hxTMuzWCwOEh/Z/bUeC/feHhaVaShmekVm5U78vSetSLgTxFIMgRuFk
UHDylwrXy2glFQ161WfPPAYXv2xwyEoS2bssMDQxS4VZzWb88j1rDkKKACVT3N9p
OYHfT7y0M8b94BRdeupmu8flCi3MgwyqMvb/JKPN7cA74BzzsHGpZ41wTJuhfvgt
1F5xxLu95aSVL2fN8bfpeYhlubYoInamNAwTGcXUPOMss73nRnirG2RWuhGoiXDy
FcZvWH7oHWcZlgC4vx3Dixml46n7so6s2xerNS3SWj53laK5X6aq5/V3ZOHvL6Mw
i802+Kg/+KGCaHrJ9ApwH3AS8R8aGKUIGshuZBf3JZRCn+/d1u7BNWDx64fOTCqd
zyeVS/3sNBCGAh/ltbpkCEyVd8z2KIwa4cYMbq8IVDvZe8+x2oivncY7mZ03yBBO
sU18hot4BSyTVKbtPGWtdp9wNvkHkWQFoagN1M5PhUJKZYymdu1VJIxdoRJtNpFA
ZGOJJr/yYS69kaXbNTSsBAdwoPqgqnmxsg8UHB9Cp03cr4k/9QVuLWO8LD9VqLEn
yO7k7Zfwvn9j7qNP4TPM+EWll1KuxGUHNJI3Al7E0Wc3PRvrflTMJSdaCo8jfQoQ
ztHZt1N3zJwaICY2Kd+DVRwIqeUYiDZDEoDTfX957bVcfCmHt2Q+DK8+8MygqrXj
CLy0S9DJVTLgOkRVeAt9+KPeQ/SsUZIuEjiw7nOzAfDlPVfcDr3ijUeV83ClQJmA
U/DlTMxHftWa2bwxtTMpyj4L2H3x3QY9UlnNdSTd/sKS8DzDDsVNg6wfV1u/K4h/
4RcW08KJERZ80dLQr+1CO44ddrQ2cUqL7GXoVHGbdVche2uwjNKgRmiPx25xUL4u
D3fi/sWmZ8wGEzn8uaeg4kIVyy9KdUlBdy2SL8rQyR2bprYIdjJf50gL83xcHwu5
dYXlPA6+1VBxYNu06DEq5Y0YGhEqfK1X7A7ro5HuoQZCSYxmhvXaepeXlzK1B8w4
EN9gcqwm7kNiSijNVxIzYOr+DUuo5JJydAQ604kEqC8QZPYid4d8tyHuaDuoxIxh
Voqr0xIGUBJd4Cn7Qa9Bf2o+78F1OFKSHv26rCNeYke2iD1b5WMENsfZ5OyZCO9L
tkUzGDHnG/DnoXRIcpCgqpwxkyJsIWmR8i9nw/sRF+Y4iisGVcrracaySXp2DR7s
v8S3b07w2eIzt6A1G2RKTCCpKVJSEZa1uvAh0LjtazHn1WqbTQGY9x0aNj+tJJ02
TJCGvPN9IXbCGS6qaj6NpHMZa3HkIcZ0Zuib4Z/gzP+37ar9WncsYDUczn7YE3Lf
riViLt7TLoQUysFmVaf7o82jSqB7uAaXne1P1e9n8j7Es8b9pQUc2piLFHHTCwF7
TvugX5vwuFPE2CYSuSofuJAUkx6uVrjdTJRdfwx0hx4XLpXYpFbpaEH2odd+BwYh
REGJEGI1wMD2GZKa9Xe5VPKzOoV9EgX6Ln5lVhKYtmV/5pE3BvT1ZPUtQIMvOaXA
JAV19WouseBqLDFzWRtpH4piOaWZcUiFKFEydWVJb+UreIdpFGmiOKg98A9ToDz5
qfc1c01LgM1gi8kRsKCarlSfeQ8kHgG+k1Yu2Fk6/7XLcIfMGdKiDvLzePphP5uW
yv3RotH+/u1yoXZwHijmVoF2DOm66qK68Su7hHmFnzBwkL4wPKhQ57lPXg0EQh82
4M6c8l2u81EV8cGw58zGtv//cIpxXVMZJ3JoI3ISnNw/StL/eE6gTPRblh6Z+m8o
vBjZ2DZCy1Dbz4LXhFVDw8LQsouNk8+1iL0fZTZOHrCP7ke2QOVAEE+jTQIOeypR
XX7MGFbA2IFBwMuzrbbqsDbaQ+2UCt5zlCHlCfsQtWVTqebC8O0huPP5eD/RMvkj
3nwSBafGJFCnOkUBKM4vSSvqDdktjsOdpIe+2hG5Yk52xujZj2M4kR2tLxcxXpCj
NsAdXbV/+zML3jNnlZRWDrE/HtW/Z8VDX3My/rbqX1amvgtpYnR0ya1TT+4U3/gK
qWsnZYCHfX568AR+FvAYltWjhH4BdImQqgFIMkaaS+i+NkPfFhfgRi98yVMOGobg
1dVW8sN8NJZeQJ09w6/KCJ8R2cX+/ZlxEzoPuspglmVs6xoXPbbUGdMpNkbAG5O0
waiggSIwLCuR+6PVeyUB4ogZkuKty9HJzr7FHgMo+QH9jlDFLjlCvwFugBaYYZRH
tP4vdx6iwrKJGkIi7tVAtkl2a2zLypFDhXaOQyFKBZIA/aXnT1wA2VmE2dr70Mzn
PxvKgMRR5vl38MtbJJXonZGw4AXNU9CO2nkBKKwx5sIQm6Cud59qMyZVV+EC43qX
9EnK+gAYw6dG6W9kxuySro2nk2dlRgbeiVeNpxCszJz1jpXk5LdZvzYNBFRiqeYq
HQbFMOWPpoHJ50kFtmJKw1+/RttM+ARrz0PV7LcAdULoSEUAWlU9W8hPiAkatX+a
CHNGH5FXBjlXmVxyL9Bi2RCsZ81/jO3Q8kA0/hJ9jxhOYkcjTc2QwYOvseKcNE9+
sKFgkE6MJZbVFQt7bjdUCLMOV25lelaqpqbKH1SiOS4VlVLHOzz8cXdXTrRk7ySV
PvM0Hkemqk2q/wh5PMEhE89zkHNDsUelPRnQKV5p8n4tnqMDuotdzqYOWIMYxkYc
6c1igkYanJ2mKC3XTdBuC2r3/mZI/A+Ju+Ip+MAh6vu2qN64ZvdKsfMHS3hDGS+p
a4lHs2GuOiGI5lZs/oq9tNkC/1iI8eVFt3/5yN0GpixNqL3HcSQUqfsavV8L9SkJ
GdnvckJAxtN+tR8HY+AjLvaxGuRhF/3Stxykqu9iZIK04RB6Gbp2LPCFYM6DUMg7
cxPsW6xjh8jvXBP7D1wUljwy+bAKDqSOM8Fz+rgGz6YrgvoYJPxt1EippVjnne1D
Uj/jkBO+vgbE82WxmB+W3+XYzXznMaJMXxu2oG5FPWdASq6wGAr8KPV6lf6tMySb
4F2HjBUhRmEtP/Ik+juHP+ZuhPioJXqxh1bR3HCS0vRAredzYjaRFsmtRN8/GZkd
s/UbXj2O1hRZweG0MQrkpdxgX7NHuz9GpWvmnMbulPgQtXA8k2A+tdvVEcClwpbr
3uyDzbBMyiDdrzeBwE4xGg7hOXd0eagGX1uJD4J1AJEUnDvNyY7Mf/LEmQqsnRDg
95fDQ6JFQv42q0OHA++e+mCvx5U5E2PJALhUgtf73Pm1E/2nk6OTp3tZ5F+5emkz
jU/rqAlDHSamf7wnjWFAQsfXuEen/rZ8/5r2wcpIZsYwybnP4vAbN0pZvdzPMMFj
/lKQCM6+XhuEU1LgXf02PZWWSgQZ2ChZ2zcQ9h36b4PhJsZ2/j7IN0tPD54SxGLp
Xgrdo9IqjyBI0q9OLMV5nCmHjIREm9lDCCSbJTFa2GJ2uthUwhXSIZnjOIcMGN6B
ZIt6bETv1xTIO8fTs0wD5oZ6X2wcPqYPv+gNIjJx8raPPAS/gVcfQKGn21RazBXO
ETipNoBtlztmKnXjdWdnVAh/RtIBYrIBF+5CjzdI3CnYEEmPMVlviUicBqOo+b1N
yrZXzeGl3+iY/T7io2t1gzPXa+694XNWdmb+qxJ6gzlRZW5eH/11fuoLbJhojQpa
69EXxz9WBKcZIDNciaqbtgrTc9yX7l7k0Q1HTHjjWI2dKJ24V5GoW6qOdkrodHgm
pBQvMXlWg584+G1TxXzHLaLBF59eBik9T93mTieaoximWKH97ZVYoGmCxuK8o/dT
WOfA5wBWXkyHKhF+sxRPRvugOLru9TSkYS9RjQ1QLfYNZ3MF7gyeK7zkcC8ifkSO
votWP8PsQ/OoB6f5l623M1bqKJpr+patROZXcY4VN1Rspk96ln7h59cZW5vuC0Mv
pafQL9rWlCsbAZB2Qolh3hrugXn0eE0L9pSTbtpuSDgN7B2oZsrJgODXEwkuwGgJ
fi6xLFqR0y5xdZjU6Guf1PsjA73mmPDax1arr9BSD5SA//DQxsRNoxANEacHq2uF
eDCbMQK4S9UpcTasEyS7DnmZ7/vJ++mC9KLaWeGddkBWtrLoLOC9DUDSmSow0Aa/
6Al/htC6t3kyAnNwfvat3COkCIT+OBr9v0/z0jeAgKnq1Kmmp2/Rm66TGV7pfpLj
X5hFlgFiuZ/EIvgHGjVRazJfzY2CWjZZHYtE3QwNqB6nlKoZSdaWhjH5+uSrZPTh
Nwid9Kbzi2YNBC/bJQet2HH/ZkCEOguvwNyZeYDJ5H4WRA6OY+3IYpn0j6MYf0S0
8bUwXSEM7As6ju/brsmyv5an4hz/QB0ehjw4v0UdRc8u0Wy0odeLYz+NpcUgpnw/
cAh8bQ1SUa5LTgfQ5fzQ8k8CtxRFwcxjVDwUSOdM0WjdiVtskB9iVIWdSrqUGi3Z
ZGSpp8XrqKJDnexL07un728FOUOHJotj3visyeEapzEnCkp3Opv2PmppO3PcqNB3
oVlVYddTk0N77SMD83rwKmZESsCHIFextXk7lQHdg+sEpc7wryWFt/AgTuv+qPe2
yc/sLRDyUjj5lppnqyThV84ahXYNoIKX8VQM22z6VrPoY2M4CSltn9dlcDWsBqxL
lHQCwIY6AWXfGxi4JxSDlW9SidbRjz/ssFf+m8FRm4fxnA43kkJaTMr8HRLzS40b
Zil2ySLJcjPPGAAX33A8eZ2Fz9+jewyVHi/m+8NtPEyjgmIgb7tWBHC3dh0oZn0G
qEDCg1a7MgFcmIkZ4stAcugmcxMxL0GuN2FdOuA0rB2VOuzbQrlMxsPjo5Wxn3Tk
zMaTJfSq1q9jY96GrrTM3DA9xcQ4wf0PEhQURl3c651E0j1a9uZFOVGI9YVW5OfU
pnCVlMRRn9n6eQjJgvdeutsb9mwz3GlN7iXI/8PK78V2wrTiHBFNgGRK4uE/Tf06
DC7Zy/QrxrDPuRk+F2s34swPDN0kJ/SktYAs6bft/F7Dw+f64xaDlog80xb+psxh
SxQc+EcO+U8usxmqb3nQJR7sH9dQq89PyqPbYblAsXzDm3T8EgOzh+TKywLNsxc5
zaMbn6husFxCB1S36T9mtN/P/9m90fFTHKjQkbKENsKiFLhvDC7NyXwiD47M0i9c
dssM2vbNCa3mFvZwOQPHL8uJdVl4ejtC2i8udVU1okaRL2sPtpj0PBgIlVdR6y7n
/Llf3MhCEtokz17qop1KggcjjPKkn4ueTpjOJhKSjh5eSwUaqce/jjBeK7OCTMhK
yqeZfyt5Sq92dFIzEG0WiHbx7aCENO2QKjmOTs78O/tx/QgTFrYJbTgqDA/OjZiH
shgkm86Xk9f8nxwMrV0k3ldLOecKzFRZN8bv4bltXyX99ER9pPwinRzUYgdY+FdF
+cZMBxIOM+wkTGF5PY4m8qmkzDGZsjf/v373q0pzi90KRcZN0TPGC6c0IlY8MazM
Lc/vdw8ATfUoK/Hya1C3zogHuCbmF2ECVYfehc/7Cnrx1H+BX4RHp8SsDO4Q6nxW
0zyRZ+S00KOYSpJ9cu505qVKqsoj6wix5bQtwGSXs/BmGT0DZ6Q1E07JtyhAdQd2
N8waXifMXC4kbQNxSNmDtAfFzAFIJcX4cvuao21FqWvdBIzRLIW9twQEquhT7X60
1P859drqUkTS3yuNIvbnCcaJWkqyB9Pmbyb2hFrQjt8U5EocewzxYWGF3sj9LZNU
HGLAcOE8bAMT0DmwEf3M/tOE4kJHsHFCU1sNJEZI6gn1Rs50qN3oQD9RI1tOznUy
U8KtqDCjAD+kOcE9WP8gmCLjldPY6HwRkkUv2XkvmTvOL/EBhhOW5CahV352Uc4m
lXAuoBWADCwN0tU0fNT++cU7ha77USsxVYtLmAkDRlFetBXSDKa+gbI5Mw6e2b3s
8Cur9IpGPOlbCfWbmWA7O9K3MtLPxFfbE/E7mNQi/Uy+Zwvv7OPd9Qx3+eLZEfKB
lkKm8dsWIyQ9V12reZ8sYtWRXVdLn8cDDX7I9PkSx1JBIiSK3G1YKR7U1RMCNUt5
s9Shhujf2W+KH2qXMirzg5xe7+Gh2uud5rFEDRhqBmRbzfwnYqY/iXUSHPekMvnl
yO60i87jVeH+HD0Vf8gMokub0IkaTt8ZPq2pH6MDKyMPUnCl41+RT0kr6XHZslM2
Acxn2CcBJ4EYpttXbciWoi1NznOQoF4wXX4DYjW4O1aycLCG6z9YEYpXUANB6JEY
yewt7nNLoP19SCG+x1m7XMafPB5T2J1PS+f9e4wHWLQdMFHERDRuHzbVeI/IYC9D
xnSrBiXc8n/aqh6njkl66S+oHYKBFWJTZj796n0mfyqBx2qD0fC9gKLgxxw14urU
18mb46WfSC/suJv008kn5S3dKX7M4CDGRDFqhyPGFVaAQpkEy4gBCx3W/8MrcsWb
jDek+QozKPw4Ac9juJ5jUQVUdrCJ6qv4tfnqZ11Z0NQB7E9JHEJ6W2furAn9uDP1
TYfRBpips1fyk+G2EAbCjdk5cV1n4uluTmHuAd3Rv2AjjEGNU8ZBUfh+h0ytAQiC
zwDYFCmkJ5XY6TjBsfVn71UgLkZDeev0rpGU2TO3kc2HReNTunDjumk8s75smct/
VbSV1Umbq1GGX+LCvPpzAGO+hvtZ5SGwDAbhN/irWKYuQgoQCJFCKBA0fmIxmg8j
trwEDuio89ZXwPUKWwpoFYLqTa7hLnBEjhJHZslcLcwDLWaXIGgYYwpcqoE/nZw4
UDgpiWe4M1zWG0xqRsXHmipkcefBVZ588CHvh68VT2T6+H281qpK5uLRSlui95l3
rIYeRTlbHxs86zT9RgXYTmQn4efQlXv3N1L00v9VkxesOvS1iscHtPCUWM9AefOH
AUxrpbDkU6XSctBfVABU5MaD37IFiFVJIBEiUxwh+MK/KCT229Ah1gu7tjyUlmkK
dgwu0OTKG7VTkSk1ouaJQYo1z279vveQ0R2XFhTUA64bWJvC5tddwEqk34gJ6d+v
Zm4+9TZWmq0LkcGM8ASnF9Nm8UdDGr0pNszXpwsR635l4dE2o+wQTH3fEPgFzqFf
PEQYR/og4N4ixJFcx3llDc8cDT5TlcRFOXyg9IsKFVjaqB5NhYt0m1kvbf2/+bXr
LlXSX2rz79d0KK4qX2mj0aJeZaz0Pn8G49IMFS54RU9LxcBzdF4xr2UW0OjwC/xx
JVomyEPi2cFd1glXAo1/15YKWN0We3ZXRDSt5YpyxYyubXjVsPz5GAvJn0HoSRf8
WmCee3NXfdRUCMMyA4ccrE+s662fuBQ50D+k2LIidpY4lQAgLN4I9vfbih4SUbO8
oLE6EEWawvMMe7ENjxyHDVolHxfx4F7XDzg9urtNLA+rdHti6LaLxQpSm33QyGhq
WsJ5PTJfmgNY3oSjJUFH6C2jUTYsZroOutpwo3nas6scyoZwXO9aANZexuNK3HhY
fCWlA1C/DrKyTCuJegiEMuDcoN8eFocH2p4Z6abnpLVNP9bQappTs6aZ34ponjd2
BCv0xxsChAgIXfnBz4gdauiYpA5iddk2cklr1OdBDgvmyQ8CEvoOueYPwTjM+XWX
abtDnuPT7nh2iNRdKX/Do/84YYKnPGYgOx8GhdeJUVbnm+Z41sKJSDJm5wGgy4pu
2FvFLYXOhp0srBlWccKliQw9yDWvnwm7+MSLG10B3lE+ZWa6mDcZ5zb+C1TGK5E9
Crpi1H7WwkrO0tevX2JE2MipEQw0De2zcYjNsqqC8l5YcjlRP8q59i0Tk7h4hKKE
B0QtLqqnm8nRFA+qcjYBJZjubQ7iGUJV/D/w7N1gHBQA5WtgdY9O6ZiYxIW09Kw9
eCw2c0SLuPliVk88V1HW3OBn8cCCayjTukKQrqn6f+doGZuMmRWOXFPeLWA+S7Nn
REe/V4TH92FcIXhyGeEnCz05WsCsXhDhvX7CDRGmrHNbfzwaaAsO7hQoABw4a9jU
/oyMrRuARXoAMPXH6W0vNTTiNiUQ0Y4x4rk2APFafa2QcybKwOqG7PSi4lOMrsQe
hzQbKoF8l+/Ep9UVFRQGjYDtKLeCzbCKfLBRlJurm45DAuv1vyCkE/Wel2HwZ4GZ
+zh5j2SQZs0CubwyY1a50U3+Echvb2HfZUJexnls6uuZLqYbt9kM6KzN3cOiuyrb
Co5vsz4xFEnb5aTj305jstlhGcm9SIDz8826m+WFyyLzEJdMjvi3GVu0TNA8HU4m
xcRZ3jxxJSAa6Z/WCdv12/iWAXfLKb+ICqZ75BLWf+zJjB+F4Lu/1zNaY+e4zUjO
Do6OI+ho0z9cX+Bu78DtQ0+fu6ZUkZ+/i+g1d6Z+SzqYBoURyPpz2saHRMPhAZJu
+3NEdHSV/wUUukAVKiP4mOjqsYz/hxG9wNwocpmXsxrdEdt+hj2adeFlNXC7uw8u
h7RZRyK5iiP5RuHSnLOdWQhwDYm9l7USJv9Qj6HG92PxXp+ulTb8h2nb9caFuTJg
yBQSEHLqTsbwQj0uvocnMb5pcqH1bL4AKCy0b5/wpspNES+qWvMgzkN3/8UGSFdC
AeRNqprXb1IGUl7cOuTlzMnMMRYidtVCUrUINHpccSfHSiigLO+UUK7U9NKrJxoy
P8LrSWRx3U+wdgy/hosmLAk7jndKQSXZf0/hqs25DuM9yLHzldQfuCR9hYcReEym
vidXRQZJSGUsHJAM0MHGNeutm6l8CiU/CnUlt3XIb3KFb2C0dupioqBo509dyrRa
UCQqJ6JPj7HmdpkjESwyBdsc9nuGONiC7d/LPt1PBQkTC2qSNzT+O57D46SkHEug
xOlG6CCck3tAvsG8cPk7tUyEZw9txY8EqVzPNgJKF6EawT2eQAUsU+LhAT0+orOW
kPIOEpw0Kmn+ds5+CHslF9DCIMrYdWjRaf5KtrFZDlcupxLy2/UXLGHR3CHrK6fl
wz8N6nVZDDHdRbQlRLv+niENQ2WiCVo4F7wAEAYmORpZKtEYm4t3Os+dXTbJfXv0
fD8cqBu6wwGlWMGwpdkkjfZILKKVyZQzKwNfBzt9nm5BQRPxcrMJBc4H6ulmHG5G
V6JEKHJvt76vAMUTqO1KqtQXwhl3ImiTGOqJZQagSOltiAUzcTORdnsYngqG7esF
VCmoxgxwd2Sxwm7apiekttBuwIAQosaAYAmSVEHNTBB/2pNNFgypyCTNmwCKxVns
5dnn97WwUHcl8HvGGGXVfVisqSSgdHtF1PH+0cWN2KPOtd5Nij8cW8eEN1kayL3o
LSk6uKpykPoZaXy0jEqAdiRIt9s5HxTTcFym+zBKaaLKWgA3H7hfGyqFFm4GtW8N
GOAEsMMF7O9dKzcKh3Sedymc/9B53JIm35Qg74c/5sSewZRki+455riM0NKmdtl9
SSP49RDUdTfDCMBuZl2FxobMM7Mm9uJFYAQjdMoXBl47ZNVObQtmyzj63nRMVls5
kBCNQwRVEgfUZvOUEp6p1GJIqaZ5VsbjENLj4kEF0gn/oIlsFePh4p7uJANZ33JD
VnSuqBs4Nzm+0IEzjCT0wScBDfJBvZr11kBu6KJqlW2G1E2IRiatEfbmRogWws0w
v7RGDS0KF+ibzglg+qsEIjHUG/ydbuY/JdGBySYcLyRXQFX6PqcTStedWoAUfu+H
cRmeHOMrJdp2UqRvUhPoo7uwhTPWw2547cjTs5aqBJrheCbn4nD0PIjuvbPX2fB9
YQja2UdhpK4T0GrTpGeOo76XcvUP6qUruE1R2Cydw2aAxeukAr4yLzRkPv1N1+p4
eJ7RPT9dVTu9JS5MWA/9z54K199IEq6WotvPCNbhBWwi2o9A8/RL66xSR3ZM9hw1
wJqtdPDy7G1utzSpBTHyf3EAEEianDlfXvgsU+hN1eHOXuMOJhCrVO9Y/hFGKNr8
5gQfluLUtAT3nhH1xsta7CSR0TuW1rZvj8iklohP4NsnDpW4ky9aq2CUS0cMKiRR
wexsyAKKzkkDtxzADItQ2TNkAqqe8eNy+dBTwf0fEG9RtM3thZz3cn39kPtI73Uk
KzKETJSuOJ2+oZh/Acbq+O0G/qAYl/ayBX2hATjY7fSs82En3zwps9iH9VwuF7uP
nftI1MJEK2ZSsdqaSmBR41JLxuRQnvG5G8+JNNhNEtYohivICWE5IrFfXI3VRpCn
Fd1vj9zk9VteSc6xXf0A97SD++Xwes72nk+GXlxbogkfL6DrgMg3fVmH7sK/0/l4
Jdo2PZO5A2gls36rreMswchjva2FEPxGSdpmo00lCjxmg6dmk3/AO2Gv2W2PFpiT
0S+b4P2iRXZdynBptyt4zvSAv1DHsgRobqKx+b/zk2uxm2TRQBFTqiNnY2qC0+Na
l5kPYxY0Za63AZs7thglQODF4G8v0TiII/OUu+Gqr6jCL38fRbJr8mf9KIb5oJ9T
ROeIllcVghmtrijcSmYK/5ucqFTbgYsvNY2eVU4/Jhwj5W+52PlzfTyIT6Bxkeko
txDIYYhvEjtuxyUnQEFtgpQEJcDiT6PDFMTBU6HjSt/4XvszfDNYz9qiw/YeTHqw
gpBGB7WnBf47dVpFvsnWjEyXqvcPb/B7Nduxa5f83cmeptnP93XO/3uM5yeTkSbW
qPbivzPRQI30vSko0SSDVCu3sbjMX+p+EqnL0zFQEUt4sTWexpMu4eGbAS6jZxue
hBB9x05OUgtpsbv5TPjHwGp4lLv8zy+NrN09zR87MFAaCPNk7j1bxu4ENc3Mg2nJ
Jghkv8nARm7JghM4aEhsCV4GQGZ4VSOQVBSqUhwTp9cwwJF5EA6ocjtxsL7p/xSU
V0q7h6ZU5sklTjNQrvAsuf58tWfvEf0ApyK+ZFAz2jPzm1UxbuzLK2CyrmqPA9Da
of4G53ub1oXKmHr52ir6QJ6MFMPBhPTVghbMhXyGHmOPko1KcfKv3dhJEL0zQyOQ
jM49Y287OhMqXuEXlbCs2GAnXBW2LuGih2KTl/b5Xux4Zwa3TcBX91hr5wwmIxXJ
XjC3jxHR3RTcNzcBmh1iriobuYOp75/ZMCxOYTOMDg/fBvCdUBEAtjvumHTio56K
e2ZCZF20nCI6iL7NdFTmIBI1vL9bidrIZNz6Sb8c8gLn331Qc1WJFkVe2KhaeA2f
DWyEBqJ+vjVTDKem5tQcW1ojgkoSfyU6i7EqiVVgjEjJpOH/34xGR/LyC2zxRLda
6Gh9oESWCZU3RWOlvC7yBpnczBd+F0OWhQK2DF6um1oinqRObIp8D6fZnNNndECc
UwaZBcIiu0wJCIcl4VEgYI9eY7ihGo1afPwhiZjHyNRKMEqAuwkox6M/td5OxnBq
EklOU1aQTlCjNlnKcMLyPgIEMWuEuAEhQoMH3t8BTSmIa9h3kq6J/OILYj22gi92
pvPkkKV8kOtst7bjLYhis+cB/DxmDwRS6meyGMACoL+GT41LkSf2NN+dtCBHV8V4
9KNV7ymH6RZTTUI1paBdwnIQiyTPvHcfUHXo6eM161nLG0ZzbkVSYHHIrVo11k5M
zfG3mnl4H5m/eBAhKPMyvF9qmekN6h7Vfws8tWLbR/2ULdSojSrPcwZ9OqJmX7Ic
8iflGBW+vP0LNO+dpc5HfYUHtkuo0HPdmjRMQvapgUQWSRslr5hitnbO/t1cuUEh
8ktDge8nH/OUYy4sagyLWmVkDuIBwlSn8mwhwof1xWlL35ufcj7o9YNBK8cNBQdG
9tzB+8WYnlfOlOhvzZ6Owv5oi8KXIcTYWC2BX3N6PVTID6Ex+asWzYNg+qu6CN+h
75sBb9MzuGdSTFtvlk+m/7dIRj14tYT6+iK10/vVTZ1zFoG1VqNlWVZtF186xUva
BjTsNMQ9VGcNxn2beDdUCkAEZHntgLos8ctnyTvYWTXTzFCWd0KSMpjfge6GxT/C
LgAdS3Wry5QcINhQlImK5o8zQdz1JG2UdxB2sblIbqJs/9OdajAIZaiy4JhXz1t4
X90ctTRmVQwjCWLkfHN6NkhGd2SkDk7Bvyy8s16tSXFcrUvf8if99JzeBh1+gYAv
4puINqpKM+g4ADGQjMJHWYm0LNhuCPlDB/Tx2vvAUQPP6JTCHGdjIn08HPsHktZY
4QYPr7x29ttqsEzqacMSFJxj5vGB55AnNdiRjmBI1CdZNhAuSCWy9HFQv1flJ9E9
DpMn15uBN+W5bcL1k1rQngcH/1TLXiSu7ViKcir/VN4ehEqx1KqJprxHrB0WaEyk
JwQSTfxYTLhMgaFdnsTgm4EBLcOHbWGBgsbRisXf/gNE92Y75xlJ27KCfnfkk2Iz
2aLCu7QfxbOJVEO3gy5QQBtcVLe9/ZoVOgD/mpfKPu4GUFBQ7SrfGtdBld30dF2t
xHnn3NAf2TKpUfM6dN+LO45wxIBWJ6uX+LGvNXWlCn2pH4Q3/DkGSfGWYG7kmDsg
W/ZpdR3yVRbn6ct3KNc5QkH8tY8KP62aC6WiyrGU6n5Nf+jObYuvy9E5HID26cRS
ymFnfJrMFgaJFcQUT5KQ+mVrln5xnZOLGzetvvaVwlZJHhR73uRZbM0oSqqwM/lz
uOKBGyCv7Er8cXH5EC7ZcmL3wPIdO3T4/fNtPR8xd66LOmQSO6MDpAoqSKDgQh5Q
CECtM9c8OXBrb3A/d/JkrSYcbzaZxGSBvsU5LBYUEoqMcn2UPKY/rcziHw4xW82Y
zfup90XrtDaD04vXuSARrv7+sESzIfN05BC0f1bHOU+bbrKyJpwBsXVFA7xjPBCf
WtmQxneA7mxxcUws2gEwWk3gpmrGuh6hVS7cFgsgqwy2Hg2e/oQyDI0RTRyax158
yinsfabA+g0/VYiSaNFjIa+ARVtQGmyYLHKClROZ/8o+7dBd+EAU2LZx2pJoBOGZ
spgi7uZyZv6W0wGd744qob/7AMXTaPnIL4r2v9c4WemlhZajaie4lu6bU4E/uRcl
tuTNfZ+OQQ27zLA6N2KovpoDqaibSxR/SK2A8rSy81bG4fTciS3eVBWeTGq8GXHM
LChADEObtbO3zUN0aDXvnhK0PpQwKfifRvYIUtbKWMNdPMmrCgtshx3JIgU6vlaj
XRfGPakm9siBXZE6+by8HHOgDR/lTIeGvZtToOItWFReAVvHc/VnY1xXRThh/TBp
CGnPL56oQRBykGm3RGGdCXlq3QRMwHucMLfdGfxdcJBfm5LEmyRW9NOXdOL0E+0c
Rhkg21i42kfvE77OmkdKUoWx562XOJlGP3wSgdZG0DgJzrx5LnFb3QmVGyfk+lNh
XNJA+e6xWgwWfeyayhXGvL9wRXFlI6lcgmePUOQroUtYE73kVr8z+A7kYhTlafP9
d+amj08T3RcN9uYHHi17KQVT9s2D0YESY8tabvUMveb4Mdu86Vovt7N3B6Bk54OC
rhAi6kPOH9rQskLA5Zq/D+fM7GY0zEBMk2Rbk5t933uNxLN8Ir2f69Qxs36Hwr3m
Sp6P7E+QnOUSvaKxLI4iUi1lILlVCRRY421HqIVVhQ7FBgUYXuvBmENyv3c3ZNGZ
pdcjh0ru5vOzg9Qd9Nxkeq/tN1vh2z7y8SUMXVvTZ2/PB5HxuaaJcoMFGtoRRHzA
WcQNDQo/ETX9QWTKiUPzB4QjhYK9DzzFhEfNGD6ikS+jQXIfCgTKm9Vho4SfNk9B
A/04ySW82oizKWA2nFXAtR+KXBj8bejxxV5QrsFQ1X8r0ZrpuDbcJGrDLqu0RPZo
SeF09Nw+lOGg/P6d+w+qWIK/qdP8cr4rCwutYBOEXykT820QCTLgZgq1zvI3wyCR
RoH6HrGCn7riOeBiLbdU0rrfxXvffNzX+gIPXZLOFjGmJNJxFq9JqN7+oQ0nNfnr
ijVJ03O4QYB3HdQ0VFl2lPELt2G1DMg4n65hqE3QQZ5JY/LqNfYMgLg9evVOe1hu
39Zdt26GutXYSK00SD6/lIFLmNC5SUYms48eYhpbfmT2woAx4lBJs9IoV1sp2Qpb
YnreLc65F4q+wY3kj+uKIdStxy2Q2Nh4swqlAFzrv8FFJm6vMKA9XXMjtgvbH8VQ
gc1DTH1EzAs6z8WSIHcITYJNgevt5u+KzEpqN/DP3ypP4mPXagIK5Sf++4QkalYv
9xYBmQRLJ9MY62glQBGH9970mEjMBe1kgxyJoJTDxJRrVmPvXy5aWTGnB/fcK1q7
5MjUv5CbvvHXuZbOPlmU3DJSndEF6MdYJM0WMbv8kOF3uA8HWeisv3BJ0FqTuVrQ
be9FUNBpuGyCyTOZjtidN+HcYj8P4LD4GZWiL0Q3cgQbIZyaGSitMuHRVQAR+Gf/
BmndxiwlzZW4+zwW+nEz2XsZ6fdNQmYF7KR99fd42eNtBZT3cPc/drhKHTIejNKf
ZVzKuBYkkk40cZWzllc5ymQr5jVYR1Ed3MAjnuemE7m/xbP4bp+iLy/9Y6Ld1/1E
jv3zFfORSRvdEcjXjj6whdtYkzDQEIX9M7lgyqVQqrfP0zDV0vsxB1FvYJcPuKRX
/cZ9GaMdZNnD14orUDEFl42WMqLTWSUyGqXh8NtzoYda6AdKDu8q62gxUGfDX3uA
VEbBaj75DZ7ykHZCk2lZP+qz5VsoiXAZodfFWwKlDYMRwl/GGtJC76Eump7XJlmT
jn7x8nysz1SjkWKgdfaI7RYAjKmP9Bltn+F7WB5yf+rkXD3faIxGqE+zpZvrSApp
gYr/zVQINo6KLVpHhcRKtix50QmWM5ANhm54UUlqhml6v4xN/EavsVrD+AuGWp0c
JgMNv0wJKPAYLg0bYjFzcVpsZu/pOZAsWz4JOrioS6C+1AlxHDokiVe2LjN5VLq3
+UtyOreVx0Se+8Q7WY69at2m37EzgROxehUXj000DXERGwlSiDuVvUVcUb5lDGu1
hMMybLY8lOCfE4fkX1Zijt4mvsjSjpHhKyQEpDPIQs+fsVxQwtjD9Ozp+WA6N/O1
/chEqn3/6TPjoMtIeGop4K4cZdVtGEM1xpROKnCoCTvdjTXCEadvALdNxSUrZO0u
E6aMLyK3f1tX9I+gCXVbCQHw/UWmpn5AXA/Maz2lxcoBwvLYEMWVnRIKe3yWf2Xs
4f/m5YKvUtDdAnJAfeYbaALb1pp5df1z01fYTZNyOclay73POh5E8qZPw3CF9fxV
XAfOq+9nMuNpvBKDu6r0Ei0TKEcSJ5fE6ypGuEx8cAL9YiR4rPEG4jC4X1HmE+hZ
QHw/zZrlvQcdvDn1XkVMwg3lyVvVsbOHpqzsx8XPnnFXT/AZemihL0Ynl5h7liz+
xKrt7AXjPPrqmegGBZJGBmBUFtXcF50XoD3RYdrT9wQoXmxctngfFR/LwT/zchle
vFdRD18iDq0UJr7+IYipxxJt1BnisZksfezCAcOn5Y0tKP5tcSgRIM0onUHI9DHp
8N+GAoDs981Vxbz1SvH09WXe3QizHMFXmLE1LJsb4tQQ+Uw7oaVS6UZbM+XJze5P
1aAY4p9bwgFITDXDjjmb4Sb0GPrQypi27jpsZUNDoyMDSHqthUgi1riiSh5ZTTAQ
7KiVprwpavJ+9eC1LeOtdrjd1bWJcFyG2cTPo289NLSZDOL9tVuoldYu/O3uaHGn
WtWCs4idOKDL5ZG+aEOYgX2dkYmf/WquMNgk1aF7wMTfIzmzEDi2jXjvC397OWRJ
MWFfY+ruLQlf80+Cu83rESxRP9urrVT61UlBgzieYfd1HWQNlP8lfPQbOXyGWqv/
0UmsTVz4S5rp9UprFA+XoxBu2lcZRPvHau6sHMz2fWToUbmATw8ogXiK6+tK30is
gXcpWtMat7yCFAqTm+VDWgRT2G41U+FKv1O7Lil7CdrD51RxQ/3hfGaf4PXAVkg0
oFxQCNNMWu9EpoG4/FmZW0nu5ZI3twhVAjobpN2t2I1nj8uAFgz955d6vbj55PE4
yoc0lxyloJsy2us28J0etiu6iyqBkq5/ssKfqabgfm74SXWn5M/OV4dd0bwnn7Gn
uzvWyMrxltih2hETddJlFBN5/uU4CrF66X1OMQ2LAcKsTeHdulN+wVqP8YdSfX11
LXYZIKC0Yk7qwtFaWqTTjXZCSyxHtfnEmc1FIHymBag+NibnoLE0f+UYZLcYOa9L
2ZWNqrzwmlmn0UQfKqQMWsvQ9Q1l8Iv9DA4aMYe9XszboCfGSU71HrMjUNWPxNOB
fzG1eH/IXVUSyQoRzUD4cwYlg10M2bvxystefRGRO5DiyU46qMYrg8fRsVqw5mHB
R1jOGJ3suza6GHIUkcXuo/sXCpOBxbzj7iHF8kf3MyR8yP0kxZ+eO3ACWw7PeD+6
DydKO5rFG3tn7atAlihpC5k/azpw3j33QedbNdyuJ1KmUu5HuFKg30hRML6Li1kK
umbkE2MKOEayUh4hoCaw8dYnQ0/ZYzJ86FUDqBmsMn+ckzp4kQlQ+PFCwlvazk0s
hhofIuejmSCf1Xn7Ivy/JcuUvtifs1hCFVS16slHf0GpDDhdCC8dCgBqgeQ90zkP
1JPf2BATbJYemnmPDv3K12SaEovotTY0AqhrDrclhaRH2ZUJTUerEq4lqgtqVfn/
wKVnyliLYBKFxWHkNvwSTx+BH81gWo8RpNybtuoQZvH3p0ByF96ZPKKMqC+n4wCv
H98drohQ1o9ddj2POPJYvLG2Ah7Pzxc8aG9fCMGFzzLyskyRAMoMtlm0Bj3md7Bv
46iuDiBPnHV1sHGlPjTZPNaRK1X9chHnGYuk5rlF9pO0RH7akVsTrY0e6mrTXO4A
04ZVvyIeBGeLsrtaI2NTinu6CP+ZXa254p5H0l04bxCVCRakF0gj3Ac8sSeAC+1S
dLbP9AZC5IH24jGLktjOgSwADDnbcD/qUhuYv6/ss1y0SH/YKCZPfxG+XcVqSU4H
4I3+VWhB6JedLHd//TRiF2XHmCtgua7vogYSXR4zGw7hW07nV0Eg5vsuOWTb0oKN
suan+SRUCxE4zwW1dvZ4YuHwNvNhZ5uyBoaYFnz4wBVpr8eb02f037GEBnT8Uig7
F9W5ZNyeYJkpjeyegnK9MtdMKmqqisOYnApdd6zU9LQMg0o6m4O9fLd72qNV0Em+
Jjd8fNS64Jsmid0QG+8zX0T6vwa8t8zhB0jy4W+eBz3W6cp0nKPFj4qlCTv2emvo
PtmANaZVFajt/x3EkLGs3/WCKctz0gQ2mVA2L+HjMK4QXzlxDpktGV3877hrlQ62
h2Ge4LI8XpPB7gLsX2ohnAUeA9wJcK1vBocUV9e6Gvk72jvuoSLcgfL3sVAu4nRA
IQ4G2rvHtTQ4HOh3KR2zAvcis6+h5OGM2ku/0aaQd/bpGNrNrJMgH/vjeYPABxtM
0Kt2VktZbuk1lghyx4+od5bhEcwpcAAxwdYzpdyjrxUSUCLRuwEZ1vJcmM0e0AtS
+Lg+zBT6ZoK+9Wi8HLMGi9d9XiBRMUDkIoMllF0Z+4EyQupbL7hRKr/RjYM1OhYx
Ab2x5AiU75BPPJGggXbv+4QimUpz0dZ/RO+vPHUfePIBQjB3Akiwg/lBhC3XSq3I
Z0ORjRAoNbWM7VgIqyeW1egh6EhSoSh0QIVVFNQRR1ZpLTqdeW2BPBk2oGJjNjFU
fvRs6FM/NkF+5cgi5mleeQ2UQFhvg462m9ajhJErAb+BGHlZeQaFyRwqnU2NQ+hJ
57FZR2rjXEpwI69XVRTNWBYWSmRBkIjvcmlQ+c52ZNnFy4/10DBZz0RitE7b2o7Y
xCEyA6DLgyuyg9KB7u9MsFhsEHLEAEfKmt5LDmEt6yuM+LLKJWBA9X1gxE/I650z
Zhk/TZ8xjrL9kbK8WgXJfa9wihioeP4FGw8yBCKmtIll+rhtbaommdsoL0n98GI0
xkz/KKOhvl0oeRgfGP+U1j4YkvPavubriIyOCMyH55g+uGS8E2mAm7TgC8dQI5fo
aW4UlNLKU4iji/xsFzaNawasJcu04susQb7HOQGE4GdIrRIbIpImp1EKM/bf2VmY
HBjIwG5xVW9w2C2EB+vk278eN9HZKEWtTIBUyPrZ2FiB6XBd5zyP6xj09HGpuXKm
dlb+5hFwY9ACldNrXq7jx51q0XMlYMYpQ6k3sleq+Wk0bB56zsb3H2rPwlWZk4Ww
NeF/CzCg46vf6agNQJJfScIM+wRdFHbvy9XzseOWnTfRUE9GhCdvX4eAGIpTM4sn
RjCpe2zLxvTHZ2qvF6AFwaebqsD87a5Oz6myTkrOfQKiB95EwA4A4guCV55fpbTr
AXCBhYBOwKa/HN1ypyyvoH96wbsDps9s0/+YuN0JJ7gc7+rKr+yyC6jzmO29rUy5
Su75MiN7L9tWX0xHpS0JBWY984qoy5Od2hOaDV5MOFakCmWd6BN59B1ADoGbIW7s
frz/iLLfq9Y0DVV9L2WkJPS8QzghImb77ZN0YNjOdLXZMuv3jLT3MrXBZvwFT7Km
7Y9kYBzmQ20WOa/9ZL35DEs65RYz9cKzRD4wrNoHIkZO+EBCOfUx6FByVBv6OR6J
GzYqH0CwsraJrDfxHiSvrIVFouc9ye/HxjbhwCOqLFEdyTZ0vkHy9QTt5TgdZHv/
F97k4caOEiVReIEfEN+HLxua1Ohd0p0ZWWJoZAKlp/VILZ7H874C5P0uEB+N4EkO
zXO7VQegNQNA1pqiixQPnhhDuBw2Fp1DExQ/sd6zWdRYPeXwE3wbs+s/TGlhxjAz
2sOo6MtJviFkiz8qZFiTWXoDtV0PG2CQQaPFbPQbhGyQCfOvHgMk3rrSz2FtWZhD
a6fPkY2nErf+ZrpIHJKPeG8AfwnZry+zJAPRuLqt8ThMQsxSQpylZWbO44kZBaaH
WR9f04f7DOFckM7F4vFoLYvZveXNkbIf2Aj2qPmHfTNsn+YcBMgXGZ8sJ1Duhmiy
44HUbTyxnesA1RSHlTRnOeXue0OXW0DBfCziwKd4OYVZKTCKEM7felFU60TpiEms
CuGsMTSqU5KUmL+05lKmu+65+kldxRn+BMPCvN95GuZSpZHtQpQ4QCWbQTfgRKA1
CXndpUfHK6rCr/w5ALM8QewBkoFfsQxu4OnQQxlor7ofS4n41L4ZCS3AhXGQpVxL
QXsY8SF75GykuJZip8dVMOKXuk6w28SUCLh1K86HDZPK356odxORg4RWkE362QoL
o18naT6kUtvOFF6a6Cay7lsBKW8RZ0jLaPAChPCpq6xkflGqsFNogvaFmjhMnV+c
SG3dzvsQ4bh94BpVMAF7AxSqr+LwCdAnWlQQ+rRmV4my8sMIbRn3/DBKI/m/fdXl
sgsZuWFN3BkHAJtYPc0M3G5t9gTK6UheuarFdUi2yK5LJgaiaTC2pUJEM7LaQNGJ
ADc45FbQaj4v2V/e6d8DTM2nQt2IBEqUaXILtBYzUWgaQ7H95/F3Ny0N3axijOAN
GDEY27O5M5VFTQoUWopFxawFwPbj3Jy04MabWIBYsyJgic5QF7+VAGvgf7nhAylP
+bRT1YyZGcA3iM0SS5iQ23Q/zoVz5zjptYZtLbkHzBYFgW+CIx37kkuV++sWogH9
5NoktyMfPGcO+PtAjnMZYKz1vPXDDu4eaRz7xaVUxC2w1vKmEo5Z6R3EyVCFvV9L
0NskGsAacJII1ETkX+IdsmSiLErneImUinRV4OBeop5K6gHFwwhkJNGGmUZFULus
2eT2EtynLP9Im185HfRk+yc4nCo48apP/QgQ+vvh8nidpxTF7iAkF1L6fVvk5yi+
Fgv8SBJBmK7GCCY79wWAmdg+JQmVyF6JuUGBRnQoh67dK+5D2PRaQbLiYYtJJQjy
HqhRcOxqBMFnBSpOTHwUv16LeP3zwXCUW1tgVkrMB+XKL+gy5lXd8gbxUT1STf2w
t3nvXYcd4FGs008SVx/eJUDda8KSEHWXiqu+JZ1eXVTAJbT+AMxyQvQnNQ1QWyht
xsOkzGYvuZCALCeAOHHsxO1pEdjc9o/RIxx9AYpj+WGtF3JsXHqlgkCuNnDH5ydi
tHXNLNHWvFehkhQ6AwKT4PYMRZy8gxa3jpyH0esLK1hd4BtwnhD7FAgI9O3uwlHV
hQRyAi7drhqRbIP8wGBsL8Laa7w1PQ8pCTISNOyWJgHGr9RvEn6lbHfEAmZ2MhLm
5YORbG6A9KKzKxqH8HSauthuQJZ6MDGIJ/3jNUQflTW5Px9RqNNj6clmk/Um15Uq
AL9PkCaFsjTUd0aDvcHSBiiQNyH9PEx4/LtJl9OBdW9gdiiVsgOxuAZ+l9dYwvMt
+n9XKkYQx8B1YBADHCeOEMX1ENGwCTDx2iJ3VuSOXPs9uRDTopmnra90tQEO5ORR
8NWSaWfoHDiRNzZ4VqYcC8y40LrmM3rpYIU4UMnkSknxvhDLi/4pofofgIlcf29Z
0Vu/WTehS8mFK4vAcezXs33dkagpcOPXKv2aupH609yyqKKc1rXShXFnwuWMDxL8
/jVdMSERR/uFY9mtdF0dOu+6LGbYI/4SC+fzbDvPe3q8+QqQ/2G3t9Po0N+v13RA
feJ3PS+6+KHEYpnK21kndCAchlObUc3xj2XBZNAo91nIZmo+PmhR6k+24h0j4d2D
VrSyCvWhREyS9y0vvwdNyz04JOzBdSxy541YH2ahc5c+XtDrNi2LIHqGWyicyiOL
Sy6Ol613R1FRKa1cMHnMkW5ftXW0SgVssG8rpakec5ouzZ4YoH/skBBsjXR/C1mB
3xvOCZPbd6t3QT/brtkqinvYh0lJij7blKzYMily1Gp8a9aHsJvnaELsLkD3/tjx
SgDicI0OklNRh3KZPwOptp48t+9DQczrzLdc1HKQ30Dh8uzkbGkWfDW40TjEQ9SF
W/MMo7qRYgRds8GKTdTM9ZsDN0hJX6txpEhE6e/rZrJl4EE95DgWjo7eJB95z6Hi
rfgd+6vZuJPa1G8qCUO+94v7704/Qcx1KFNxdgyJzv0OekzXJkK/n2exuMsL8aTb
LLNFy13rA4NAHFGKt4x30/8chQO/re0j6RWNkGehN82s9FDvn3b2beeQVnY+EUmx
SkdWzGNj1jtsMOkHW0EJFObrswXhz+Q5ju02zaJichuSaCZfMoAy6fe+SROn3ZI3
g/XeV5K+38TaV1/xEiFy4rVP/GhoWb93X98FX3paW+Kp2fiGkt5l74gnWzBk1Oxu
xD8lWSKFkJ+G7qLNCeP/5HdQZ4doVgNIGqyu5OOH4OcrzCDSxzoTo3eTM1OLUiIW
Y8MLcqrxjMvWF2ngwBGqvxqQ2vr9vI6nOS2WcIDBRrgxcddXjZupwcdgw7b8v52Z
3ww9LTGIHVsW9FggobLIbMoevzxfLLCnWFq8I/NRrscOgr1zlUv3nUeA4MQDdyv6
UPVTwRxJNu80AdfmiM4Ps4GyXaHYPEHqg7yrz2r+4NU2yoMEjUGep43sHqvbYI7D
iRh9k21pJCuqt+WlyrBtECZ0f6UejnWvFkP5rHguocm0D5X3Ocz3dRG11T4ln0Xj
vGhLjbNKx8ZeC8I3+RkUe0/YcpLT7s50ULIBF02/nBCV7/NNGOWU/vHRuCvmy5zt
ThwL/5cdawg4qo1Y6YhoAGwHuuU+1c81Mbt5PjTwiPbB0DhlUZrqobwHo0gB082+
T4HRlOrHnH49FGMQMX66id2uFWqIv6GMAxgz6gwKH8AAbeU9XHCWNJuZyRKufXUV
4DZhGQY29DUL+eS3RTNVK1sJfUA7Za41YvmDUmz8OZlW3GKT9XBXFIgh3UTH5dOJ
A1nFzq6NCrlFOIPJOfGHI0qxAxwZ/cAXorotxgSTELiRaa3hxBNnJpdKY5hLXDB6
+JvP5jyL2W+AIvaNl9P+ZImV5HJWrWnb5WhtqW9rU/TyWm/L0JsACGW81pqKcZaW
O7G0suIYPM8mZvCM7JNAb74xmTb6Xvq5AAKUhcCxSGvnelbA3I26Koo6dNbPW+mh
KECqymxViFBWHK0f5DDoRuJGeFDqu64jGfppeRgYtTiTZDYB/gRLKUI0eLQMA7+h
vZbPz6jTuAwShQPGk00Yvyx4aPt1IyJpZOEqaQS4ptvTlV5/sSaqkywUrSJhiNRB
dVAUt3CfZ/6cJf1TK2jEGLOze8F8FgKc8+QJ5xZXxErdFVdstK1s0gHS1H2k4mtG
R6Bi/3z0J748OuR9JwcK4jsX5CSDjggv0BHjlGSbWd5gCmfOJV3se4nJBRYI0jQj
EUznDjMUAAV91Z92dxFOq5Y06TC1NpB9TA+cpIic6Ch34ReXQ9MrUN7Iv9mBOwdd
v/BNmp1oN9YJVdLKzgFADjlUnfQgAphp9zIDZmCx+RoCMmtSbATLg2R9hjK/VHW2
iE2zm210PXTgDX/0yjvNKyHvxNsBmJiOB6bRqRO0OKfTnWyRU3Motx7/VWu2DEBO
qf9fdV7gCvsR3o2imtOtKztT+3asmMeESLkZQg/WlgKW969MyDEqlKlpZYqhvc+C
OvbIeiSsG0rFEBsChaC3Wy83g+h86TAKI90n5atqs93987pqM1epygX9y05Ao2rN
t9wOcLmYjKxunRbvTpnBHdXZ/W4R8FzMp4X95MxSlKiEy+tIrx7TdslhjuwLad1H
qs2HOE6OUB0IsAfe1BLYCo5MYuYHo+oi0eu87lR/MS8xynkmhdzajn7XO7YEuYzP
lV2/uYvhaYkD8lwTjNj4GiPDM+uQ9o52kq91gvTi8CPRWguDN5vhQRpAVEugY49K
WpynLi5RNT/MNk2HLaVWue23IxhpbTfgqmaxqS/k8NZtxAKz2cwrTPhDUuotWVvc
wyNdOsLNkCDWQOxVoQ2/EZSGnAp0LS8U7eyqedNLXvKknC0Vk7a3Np+Yh719lqKA
VA8uZReXVuG4bcnrAa2vr112Oi41NrFQCuqTnwm37orME9YDSv7ER4VAOcjsnPfQ
0YmCgfRZ2pnNR/NKG+JTfqifj9VNwxyITFeY/XB35t4RH7el+muJU/kaEeTIx8E3
kMeYQssLwAYEgg/bFmbHL0yS7luBtt6aLav2aSU9srDg0f5CmSiiBLhF4ovE0sW5
3m81d+WFN0MK42LWb5nT7CP1VfpDwhca2QFp21TyEN3E1FhJchP8wlurmz7ygMt4
mD5MxSR6COf7r3j8QcRh9M45VYBVIVMsdXE642RmL2y8i5VP1MYSCYiaA8x5kDLl
zxbYxQjv8kHm58eNj5geeSmeaVprWnfGP13tM2HHMkyFteu7uaUzg7qE6e2OANkp
Rrdz6lxTCweJHWI2gXFcW4EQrpTWExgcSIpQ5qbSnUS8Hb/8CJOY4r4xttf3Y6gu
Mw8t6tILt0U/fCOfRupaRAIC9vkTsBpsKX8njFcdbbI51grRXhElRchJ2dZs1pqQ
7OIrrP/pHn5S4Fl2qW5MW5rPwd/iGelnesG26ms8FYnE8tY7fK15JUfpLTp7RgDi
0T4Y/p0keJocXbaLE5TjK3gFA0DeEhWpmXcggOV/3LVMo8pgUna+eWIR37IuPkA2
rY9LdUIdfo/vArQV60Wdhr5sUvg3WNEsrpZmC4ZAovHKKrBWYhxpHp+egfJFWNle
TR1ZCaOdK36AP8zlKipqn0VffREO57ls8QjXqiK6A09QSoFLxFWD2ZQLU2hMc2af
R1pNzGyGzGByEcB+uUO7ywaUNC6b+WOuRB/Qt0bLC5BaRdM83s9I3Xw1fgTN/2Fo
sk3RY7ku21SOtYyV9TEiI+ixSkz8WB8+CqIdMY2ZjlbYA/dpMPOnLeB5ziTKXkjs
YEWYKgAgPCphdiw+wIuF67R1Jv2ANveF6EUo0oL38t37AkBiTH9W+D1FHqeTRTD/
EH+qEJXGlI0KiMxRYbwQcqGiqP3zOckbu2uOeV55STxAsERiE3roK+rD2aYEGJYJ
WF3acafg7NMwQJqaKr4Cgg/uVK3XHqRw1kmwf1Pny1yckChvRlxDcfNzwSH9QFpL
lq30GPdnYmZZok+/llDufsBiP7patDFob2rpFRO/3y+79HfyOYkWMb0I1ByUaqiX
uRHo6IY5TXdBNd78pNZQ8QaBqqNtfa5ALQPAXd+h4gNGSp6TqkKEZyxe0zm+L7Uf
bZ77D3MwcqHyk20mXGlzU3fV8KhkEYaMuwG7Bbf6yNZiqQoQI0T35pvIlbLOCutC
449SBeYzA+Y+J75ds5qq081xvglZIRJNvFkgyc38gobe84lXMTzDvq5tutzu+Opf
YprAyiCRvbaTrrnhIb0qimdQljYST5tcyZz7FB59u0Bc69+bDTXvcgePxEoCEqlG
0csWvfB8dAx+Ge8ynjrDlt8DliuKaLwFghrpuBYxMPGxVqKM09NoEBdvN0SKZf13
9KOEbtBdoXHPWoUlV5RxAMfoI6oj+hIr7TCyggMXFsw5htqMaFzJGdRQy7v+o3TN
KzD/Y8kXF10dzQ7Sil8Q5WjotgZmPc7pYrhM7DVEhLMDaaVpcBDYUAc4RBK3hvJC
ZdpupCuPRl6KEFH5nh32XqvZYTx/8JZC8tkvpSXt/KAKf+n9xJI3zuDtkDchenEl
c3n3Auj4or1vF9EANnawgAwEWQMaOgRGrv5ro+9cbVcYa65ph62REct0agh5qvjo
uDyjoSIz5+WnKM7XAwjb5h57znnTmXz6LxSpZfMODvcmeR45hRsxJ9If3tNXD28t
WzITTitEqek7ya+I4phHYDh2qaoS4tdvh+rSxcUX0lbks7k+M/B+3LAVYPXsWFb0
392S1PsiWgwgsQsbh4kGNPGMNCUGJi6Wt3fOZjz9IkGwp9MUc2AoOdCXc4NraXol
e1AyHLXFgzFofxSsKh+z6lEFXPhklC/mhgbhd9HGdMJs86VmD9XSZk0lLiiKU6YU
CD+kdZXHkT2Rid5gHiBMf+NuG0dLDXRH5dN6pxOgHA0AzVTD6SAPMZxNPLbVxknd
QZ5ZI7tKjbHQNESvAAo3t/G1wwB7gqBTn2IFahS7zCd58ot1mVS5V1H6Orww+ZBB
6leECWg1ECr6IZ+tkNlkwwAzO/cfGdc9TZzZpntLq58Ld1nc5+HrFbeoUf19xWsQ
czzS10RJ3qgXBiQpcsJCjjaEiAteMJ7Lmzobf+eNOl+eQimKyKQMpDi5/L/ahJ8h
gNEH/Y4nXOExLoCn0W1eGtOgUoYQot/c21PYn3tj6oznHGdhRBrMBHvy6W5e99DT
VVFTm9w6l9FCeEoh55CW5Zk6dM7trBhQf2Cc6wkUcpsZ0ZUqZ40XKHB5XYxpAiPw
Ph7Mz2E9Ntvm/04I5LxHRJZToxXe4DRcQDy3/D+b+9ykK9o9e5Xr4lKNnyxDC6wn
KhKwdb5WiJxzLqbvLdfBqDl3cCYyAWLvdz3oie4RdyWUolAq51J1xmdSsD9byQRI
R4ZtH9mEyWUZVVxMg8zW6t6QLPg3IlaCRnWqwVeQ7NmEYRnUvj1cxE9hPR9N3mBG
CqKuL4GkQb+fItq1zO14CjPPMPGgknrSTuKnUsInarRoxSrs+9Ra85pWcROybbF5
guF9rXKBcIW0CNFC8nwfqdnBTjUCK+/gBU9cOh/6X6cgEY47BTq9im0tCIeL/oec
BNlqR7xHPP9qDQIeEpGMx4jgGCSDBwJQdvR8t4yZkCJQtuPzCMI1se/2kspXVBye
2knXAgh342sjO9MJ7uy7PrzIA10hvqL0+9j/9NMDiGvFcw/6pBkup/YEz+eQCzpD
RTHlEwnJDUmbCPBbyeHDSc6lE6QVCzcGkBF/2hQp8czEtFSmdq/ICaywn1Ki0G07
bBDKIlKowlCqHdfib4p60CnrGQ8OUop6cimkmPD6fwWQV2SkTqpRZQlU23Q9YWlL
eP+Nm8IrfrlgYaT3LbLmzup3st0gLSeiIffocuMAYPlFC3O5nzTfSjz0IOITWAqy
iXvMjiwJgnMCvwy5fVojbtGwOUJCROLo/c0RZqtEpArGJiDmU4CKEJDoXewftjNH
mGG+nTFMOt+sBb4ads1AfjLneXN7TJ1fBoo0b/xDuXEw+p9DjUbMz2eMohC8sOXH
Luq/jlg/yASE44/Kj5Sp+g3DUpiCAmXc412pHOEJAHhwfEXFm9vllMde0F8AaZXt
QMvWc1xLWNB4ITwizf2Aw2KjtqKeI4hwTKXKNwXypD1ie9S8cwKregVib+nCe0xC
FFmGmd7EXJBt5HdutzDE6sGZQ5DL/NmQOZZYE+hJG0S/xrSDrkijC2pYe89iZtU7
8GvD5VqBfgmVTZhfcH348WulACzgKFtTxFaL3D3f2B6Mj3Z2DNiOqdlIFTsE9nsf
UCr+KNmtGYe6rk1i5ofHt894PGQVAHmI0cJF/IQGH3plAoGxDmfLrIzZ0Ue0X630
FGFXnGZ45wHTduh854Z8swneuMWxolAInu5QwnfCQC53QAlfgh9G+yHci81nsW7T
AVrq4Nv1uElzp0quv+y3BpK9SNx+N8kixEJK6bn7+46LSlOGyfaehbRa61rJ/ysz
YccULUUsRIC1IR4LnDwz8MT7N8US5E4Yna6e4jvBAisX6p6GA5suMercr8KNxBeh
v8ZquYubAqk0KmKQjEd4mxBOcOYXk3uKFksDt04uz2a502RSGTpZbZztiDyrJ9W7
LDE7JnjuOUGVW2yHiiIwPbC/RTO4kkQXJStQEdwrMoeEd4HTdErvacVN3D1KJuR/
sx2LMEkk61r/zYk6KBxeHA41r337TWhewQjvRv/MqxqLnlaQKB7o7g7pkgJ3E43/
RgDCvi5MN+Ks9mdZcI0cgyUNn4+asCSqNeCgNcIl2+zdks32yXOj94tDFtSzocTP
srJSe9SMomKHrYbo4VX/sGAT2LIrEF3Ws7+KLxZRlGH/OGf+uKNNKMUvwVKgsy09
O0bSlxhbolGRfg67hM+pDutBVMGXnXMQSc9JED3U2R1Fg2X5xXXLG68vg5J7LG82
gyEEauW9auqLBpF3f5QXWrLrbLWT9KTEw4MsJNEgv8pGPcpRCqHTlg2AERZnvtr+
Ox5Ia1ysaax8pCwBO5bme0ZsEL3FJCmk3aqCZxC24jhl8NRNm010UEXSK/cvvqOJ
tsYNobEsGp85WuanVsrmw73hkmv44nK+IH5HmHhluuga0HZoQur2Htj5gyhBdjFH
ZNco92Tp3IsvwOEm5DZr3uIKtvoRp1rqloXwl8Za+5+kz9kq0hqxecc9npRKseNK
PeMIEIFR4oHZNkoFQk90/ojFhHfyovUcNd8C4YNWrPl7j1FIJC8Brl/LIpHoQkP2
clFFGEHTHbmI0XRFIu6je5fhc+AlGGpd4evP9RRaDwMIfSZp6c2QpohdAsbiklmN
P2QYIL7RhCzAJku7vm3qhU4mRGgxIv8Yauw+LbXqxz4v3TxMNRsMB6GU+zY77e8j
oEyZ+V+NzOkzET7AN2+wv4V/Ek6GR/UwZhZbkRs97zY1JrT5YpIguIhkOJ5xwFFx
+a7FcHUxgnsMDhJPpeo96tRkFMGxeyT7tpYjuSvebl9t7Y0ZGrsaQrz7w72xOI4S
HAfZhaLjW+Cw6I3G14WFeKIx+ZWqbbbhA28MMxWt/ppsTBbbJz8xiOWkJOEvDsa3
2V/tISHrc1clEFAozct0ykYXN37ocQDf8bqnsSzZr2nWU/XVammLNApBkQIeEMIG
+bfwbl1LToJeJaRiHcVJGhwHHjRl/oEBJKRvRMBjO0MC60am2ERwfGsVjJwXxdVp
2by0Y5GcBLsRuV+/iUCqO2htwBadz3belEJLsHWsgvqpDpM01nNJB5tNBi8TkgOb
9g0Z2H/H7RZr0Ix3m6eMQ/IjTvAgLzyOQ3oyRah8FSPLkCmrlVnVmJO9bUCGZUBT
648kRT3OCQIpybMh33eSklhRJklJCf2HBH8uaoIg4waURqVmOP4mQUt3bgvc8/8y
Ov4225FkEYZU53GhePJt5lQjyVL/bqnJZy/DRLd8jfINOdbcnA5zv1HjLFAsSxWi
+Eh9r8ceIzJn6E7L522q2uclbfP4KeR6RqMsuhcGmQsyFrgkr8nBw6fpLqNNUmKK
pG/1D5s94aR4gviUD4ueaujjv7MmQp0TNu84S/W14MERil+nYBUSeKIYWoZ+3BNt
nLVupuMoeKokB7jYtkHRUrf8ZztcPaW77Wic4+O/cpx3k7wN26x886vokEGl5RbB
/bBWG4SsfPIo4tqkZJxLvY5tAy8xvtq9fx6EwKz4kCALm0DRkDx8+yR7wrqvVgwF
slEdHjyFQE6ErSCExweef6ODMTZ/TD7m93dT56PzdtdlQUzEM9GXtDdiDgrj3QQ1
D7aETyKxOOoiyFkYoDAqwsbvE+OR3E64B4Tu0rrvFgt5iIvxJBrGho0LykGexGsx
JD0OtDVzHRJnp8yi0eTBUoTk1DGhj5dQAZ6dKOj9PpWKbf0x+PCYvvQa+eASlQLQ
INzWy0coRy3rOZ/0fYhh/xyAJyLWE1Otu4VFwC96IJP4zezkpS1B3vI4E40oNdfe
09iDxETuKnCHor4b7QZG0rlwyQALVv/ho8PUAOjcyqEdePPHrvKfM0k6OC7SzDBv
6Shj/a67R4u0jc4ct0ZlQMOs7xEUPaTzfOevLnJcNOM217iFdV+aSkc1MjcYi1eB
r7EUUizv050PzVRk10HE6kGUVmzWgaqkePYL5QsRAg8F5/keZWG9w7YJT1OYWyaX
zTng4/wYTW4H43veg8US0XVvRNZ9/wdxOHxt6JtVa3Nx4icgeGocUjLYDeZ8nMI7
JoAV4TZAABogYRc2ieSd0BvuyWdlnuLOl3j+nJDg2OsAujqMhcZbGOchOWsfFFsW
E1KL+SF8Z+f6uJD5NhNL/jqLpCjosfEvSDO56n/mmhX+Psz2kBy8agJmmDMUkvKs
P6q1uZ8F5qMqtk5gXPKyFeTTr+TinJFlN3baJ7rVhoSW1oWXaRNpUSRIaL4cHIC4
JqsL2GH14XjcEOEEdksJJdv9gRKVJaUieKfCc/EaXJh5jEUL9TNmhkR5dS9KP8+D
xC5sUFm6UnKBtnlFKLJdndLMboADZkmHHAhGbAaf4q2vdsyFAcq83CmZsGy1bqgf
QJwBhG1yU4BgA7JK/uMZm5NnOHui6w5zP1fwPMgIgfqpBITbuzd3i3TBCm3DYkbX
mpQQXiVUASOGEZgV1l8/AMEOgME6U+RkifOobCEmhxTSLggC0BLA2Okh/pcws3jG
d2qr2lXLWJiyzc8mTUVE6Otmx1Kw7hetVRaUIadTErvNU+e9YDfS5Rkf3KuJjd0y
8XJ9umlZwqon319LBsRe8n7E9npQXhaQ/RNc8MvALIYadAFZGsyP7Qu/vopApwks
5x1XJD04Swxag/Jd2lO5fGw8uclVlFn0pyzzq42Gy9SWL99Pm7oMQJXHA2y+/IbT
vSOv3S73iDImnjZFoP1qJF/V3RhMDjckGT8rQf4Bk/OD6N+qzTwIDTi4OSyyuuqO
wPB/xkLf7YTd/lpWsAMKie8dbPVkl5vb9CYCsgXmsZXIRwYdOuTJmly3JfRrrMZU
JpAZGrdumzCOlrzqK+aRbLSVHLd1tueEQcBz0lFIEZ+yCdivisqL6VETZEka8xHQ
g9MyPNB4tSyCadxDZL/icN2oaebWbsg+jWmPqfMURLFVBK7l30vwVwAO///Eyc+4
2y/Kcse2+R7Zz26hm16ZEkjAA7sO6OdL4vMIaB9qFErddk2pJvdREmIhRPbC2Ztq
z8iBm9D1Om2Id6Fl7yNC7qEe7tw3Ok0EkCsZQstvar8UAYJCzHGAuZKW9PBc2kaS
JqUKcdg2ve0DFGB69/e2RWdZFrXfM/jdfP4sraull1M6NtdsY/P2LIqkMQ7C/bNx
p5kTcTTHUa5ipvLRo4PgM0LJsb1aQwveFUnTAqP/M/NsjMu7Le0f0kt+I2I6o2JF
aSIelAtGVLCCju3E1ylSE77VcO1aiUvLpTHwAtEGHL/YUVnaLkrkR8cnJXUGBnzG
27ORomoiFiPWicpWHIzTl5jZWvb6Ta2pGOb4Ow+Ej8V4W1SMeLKGiXB7vChyGYQx
j7GTRpPOzW4pgOoL4HgnjGRi1N2OE4Ys4pR1NqzgJse2w96/BXIsmmLMa2l2kZg5
Wv2g+SLHMe1ccffpH/LfS7yoYAG+X9j6Po+aWmqJPXS8ouBFn+b5jX1UNzJ2NCi+
QC+wDcHqqu5Thl9QLVL2NLIcOK4mOoyTV7K5MnaLtXdrUt6kFFwGSVht93o4Pji8
cOZHUIjMRQyGNyA9L/3p8E0ohLBy1IXudA8y1/RnVNVjldr3VolSwqP6TSBmPzGI
4IUxiNZiQAvewaK3ZoJJuWucdipCW0o1sAIYf/c+StbN1OWNEaKXTKyLAPUdyBc2
gKSDdALO3wiCP6rcKvg8x5pCS17YAl1U3LQr/fPeEsEILWbiX8BI1G8TXnFRjx9r
Jv3XsxfO9F9/BobSzJL8kiX0FqxS62t8nnaJEnEUP9miCG6gapCWxKzUegobjaBp
gLpUbxytae6FY28KwroC7Dnv++G61OOyhqBk05QKDQPtmmU4N8wBABqFH9nKmptE
X2HCGyfy2Ae5Y2Il71RiMoA5pJKkrfTOKNvMlMBmkPqy6hdxnzL8aLP6eXcHQVbQ
BQgZS67xoqQMYEO0iVgWFQ+8GRPDPhkEJelrJkqpVmYVnK2fcZHZ0sXip4jQjmex
jZWzarCUYPQirmmVLB4tr95mTOD7HSxDJSoUelhRinh0gs/uteQrxqMYJtyr69GS
CyPs5Vy1EES04FBrsd3POT07MrPimlcYoB1mwpLT9TkJcS5wiIGsi9Uc+nFkE7K4
hZzWHLIctuh8HxTLJy6JB3DD8bV2B7xpWYIaShScBr5sAl2fEEEoX4G4oij0DtlQ
DrJn/11oW5D25dHP4sd79dTyKZ+M1LL5kZ11AehU1rLBSbdS4bmeFMBajBg4EoqU
rSmLYy2qh7iDq0tThMiuLzeocP7BCol0Iz11lGqn6WZ1+t0nVNcJXa6HXSBNDk8O
JsBRFPr+2Ow7F3kSogeP7IaIsvaWnPf5qE19DQdz8zvBRdZQpMuBHIuiMWyOQOf7
Yqp9NIUNokn8tK+wPD5zl+G9whvr14eEkL77oABVCVMEj148GH2DLbhdGu1VysSY
/J3jFLJsyXFvk6y62eFH7O5q5RlIWA6mirciWvnCLi/U0C0TbAatGlEsupXcq2nr
wfJbSVhQE8VZ84i2V1fsR9q5/Qs34jYFSV6FfHrgBwG+j44vK5qjRsWK++4WXNmf
KYRTDOEBoSJg+pijFXjbkEbar2Az7MjTFuVlQX+eHMhp90eCiU+G3Cq5AHl0yIrA
shm6G8EghiCl88SauKWIHU17TR9fs0IT6xodtqWYozvd27/a2/rSNgYUGPP60ct9
jj4dmKNsODMwsmPomrBXCpkUN5ezqaOO0aJ9r3v0vq2zS1J0KO6nNBg+LqWwXMQr
rbgKBkbqRpSB8HP/ZQU5Ik2dwA2MbkcHTCS4ytRH0/qtp8KL6XG9sbX8xmWWsc7u
Fv4viITWvNAOk+dhnS/DXTtraV5dy0QFm+3rhse3Y5IAt8cDNyZVuvwh0RHp6a1i
Gqty2kUmsvIaMEXuYOTPdKsQgYeCNGeJpGB1k0UaySnr3K20TDeBkGxD7Fc56gSn
LKY47iyXcLdWG2no8DHk2p58FEJBpmdMwiHQ02m+qNYQiVuAFzq0+eelmN4Z9Tbu
Bs+eAwvof5/eSz8uhX8ZDtUfceqWM1c6eACo29QfswG8pjI1yvQPeJqe7NN/qq8H
WIXEUXCdJUoJGMiTNJK0GocwGfD1vGzXvfIWeMWRKDRHWyUxz3Mn83pQLW8ttjvi
PLYUq1HbqV/cdYpm8c4fAvFSv6Vl0twKBDxuvxz0xyTUETL/yVGPpgAAizQ0qN7B
ZQSTlb30zj0Lniu7c2LCYqcPyL48gbemGPNfFXWY9Nx5c7PoWDyY8C2QD2fXT8Ed
wdW3fZKVhJBGWrQXQwTKjLz/4xhl98BOPuvyTNWaX+s2TMy0fskXp7o6Wgm0gtA3
OIHnGcGHmHE7FpnOw1bUcGvV7kNVX2OaQwORJToi5QfJx1WZGPKC0e09/NIhh4l7
9IqtDTg6VQtyR7xKNvpuPDba1EOYy1Bt+kwDdPeHtfB0I2bCBvO9iQzCmti09GUK
1E3EIKyPxC9pIc9EvA2G0K9cXfx2MeE4AQBUFupMKZk1hj31YFzSq92vuRzxUtHR
RxSEPnnTFFdP3A5hgIs/4FtS4beVieCYBulF2wNK1T7gqwqBQW6cWa5kDfjIgpDB
Rn5kewjRM2S3SIWxVYV7KlHgJOtNkg3YkfWTmDdwM8BtnXjW40S7dhfXNZc6zIHS
iDvRbzHWwfqaOE7uDrKdAhRHoef1CyJeDvyRXVvzNyzIhYFwJoQubaEhdNHh+Gic
Rlg/HZZIJ8YeCq38hNYN5hyFh6Z0pbqroyfyMbyxtEdiqXGk96F99y2tjlX9LYFA
eejj7Htnwf2AekVsUJ4U7A0VQroQBuNN/AWZXsHrSDSWzCo2ayoJwkKsGY00hhxx
BLpEmnqrTk/Audr0BW5+V6/LoL+c1TUuruja3zbl/oGi5X29Y1izOpUav9HveD+1
PashICDL7dFPLU0UOVKEJ5MnV6btbIygBrm7cm0vwfA4/uS8LonHqOYkqbGZFhYn
OkHvyUPUh2bDHIO/SxL+oY7fCOzt17I+bLWQfssY6+FW1YvJhEc5eE1u6WTJN6Fq
0bJL++OB25jrDkWbZBAGT2643jrdmsD6CUJ5Gs7mad9Ut4An6U1YvkEFuQZOnVfZ
Udk2LpCOriATn/RfMc9fw47zCz3EKrsGCfzwSFB+traYts6LOf3YZBpIv9CUq6Tk
7H/apxZBD6e0ZOHcFnMleQ5mJDdkAiCyj4rJoX1Fmr6jaoRDa4rTTDSMHkOCekne
QW4kwbEi7QbsXiE4lptKkqwiiVsgJuTn9HL825FnTx9ohYoZ8p9tWqfv4O7gjVBJ
7FHRabF+Ivm8tgszjRHHpeJwngGtvza7rkjHjLLo7top/ik5pgUna+xjasrcuTaS
Ha7cSY68LRSobhWk0oG1T9K7DCvdWTHS4OqruBRUO1QapP8rPpEEqdjho3Ad6zuU
3F6fe8vUkwfLUwkZ9aqE2ZbBczZd7D+SalPKZI8BzZYr3S6litT/pc5h8sle9+xQ
WA3iFQDDbyXwPNDdeuAZQ5PqpfvnN4UaWVpUcbDsrJ3sTAR5NxklTqE55BNwIWb6
aFKLWVior+RtKlGA5NHFEYSs6fHaUrBK8sSDB6swaarIaNgBUvwZseyqJXilr+lQ
EB+Nk4emYLOQIPRbKTbV1TvsS/2mHLAQBLcSxukDYouEjVaj11xbMZ6xqsGTI7nQ
FwI4jzFuBYnmY1rMsOl0Pa1t6ZJVYRhzliUcCIh5NHAsyicr3CfLw2kt9zIumsvl
BMpWGD99KQmNV8WacmV4vKVdUYDigPpDUfdItBCInzRxHAe0DuwYMPzccI2R3W2p
u7WMElM0ckg6j1GKODYOrsBFU7A3RrWY6ivrRGaHD7mwlWkfT/Sk5AHhcCg77wQZ
ksuYPLqiBwyPV5N0VKr/ZfenaY5ber4vcUYSnUNSQSaThfGAmGjRsIyS+kvNnUqn
5eexAerXVlrLb2H09TzZ0CeJcOtf/Ko6ZzQSh6LgTqzgp5EJqGpV/cjaauclIIx2
DGCoOMa/IGr889Hgu/52sMfC5kn9rOZQFEUrmVL043P2QTano7hTEM5LoBC5FtkM
Twx6ZbPEX8IyuhxaTCnfs6jCuvCvdzXl/znBA4CuWdKz2MWV+VJjcgIFobwgCfgJ
PsK0nPVzMUeeQWf4kwh4e3F4sbp/hoEB2P65BiY2LHdl0ridqEYe+iYX0sr59Uqo
htfyE7Qv91QjprbUTgRcZRGTnV0/+selmjJkpyv5RgXMnFHhQZqBUSuyudZVBVMy
LjlJYqAJup17s242d2b2Sj1+o1K6lpDchBs2RKMCsWAgcXN00zvpYSXVtRTAazVI
RaIhV6ecUPTU6bZW74IPD8H5LHikr/OJR0eywAyTVolGOGWI0XX59tYPgYYSjhkx
H0UYZD2nr9TCH70bceznjODxB0WpulkBV7KwprGTZAF8idX8aVxloGjPkNfVMHMj
FeKOMV4m4Iky8gMI7kOeE7gokrsVu89pXfw1MFDgfi3/J89zWKtPeHHO/T2qwMMW
neG/rUIiXSd7V13MptR7o/NCxoEnhKYIxbmjJ6i9qtpQeM08aAbt1zwTDTIqwSCs
P4Y/1xHmY3D51mBezuEHZEeqrgsfMJnFp9SuoYopKGipSnSK8HM7/BnL6aXRMznR
dQeFO2mf7SJ4XLZZDjkGhJ3rAE0DmPeFbFdmDx2PSrxfwe5/QFxvnsvBZpgbvZFB
W9DjwBreXXa8lFbxywrfYYuUvQbWKbjSVCHZvyUpi/PXzwnTS4lzRbN5a13VeJcB
G+EzqmA8xsBOsoCAzLlHH/jQM+1M1y9O9vB1NruW/AjojfWKE8OrpbPNKhYAHY39
DxuFQ15fsEAa7EtXUJsRffd6Y7QpNNW/+XYEJs0F129+nK4QdfcF8hJ6Rrliy1+P
k/vtKrB+JZGsuJFlFaepA81PY4XY8/yaN14ufMrowPlB+D2+CWjhILv7cYK5Rq7J
CiT/YbLvlaNe8VLzX1ZlmOzyCEpNlPCse7GowY16bpxuHx/rURe37aJoCa/V9Nm+
Hooj7VdNh4u8NJ6eTehfwXAsvj42o4e7r49AdcrMrxBG2Te+0GXUJjAC024ahITc
O82+s1VVruzUBQ+DLPD/B9Xjtt7fxVFoyiKzcF0lOtc3tBh39b7ZvQig5/LBviw/
elFiyBwC0mb0qrLa23V6yQKvL/FcZTKEZCMF5Dxm5TzzS8H1kK8I36sxXKvd5zjM
a2J5xI+QjllAHAwsy0sH2kazba+UB51WOjjyDWx6rb+zgn+FVsOPlksiCtrVkcNK
qs8OnZZWKGId3fbOy7PMIQDm9lRyNrHdQlMf5VsdC19lqU8MHLB/JRv8+Wa+bNAj
hw6dsKzojy3za9HTM5OsyGXOwlN7ZLYj39SYmKb37fbYV4BfFWln6IvZolonx+dL
/Hti2+0QnCOfVxg30OPVcxKDvPbBnPgXCAkUfHuSQHR+EMQsNs4u3jXroXhoAP2R
mhNkvjMv1dvOrd3U9FV6SbhDn26Ix2o+H1Iayxd9U0Z/zQ4NEjoQZySjup8fJKmJ
xQ6j8TeOhBQiVQOptshdLPuO/MiryaVk62tILJF8gihbIk41CxsNJZ3w/RWr0mfP
uVOtm8JQwILuSNY7hpYjRwXrfSUod/DdANQKW92wSNr6RToqXeaFJAr8QixGevNk
uK2DYEGaQIQkt4TZj997Lkzhsm3UH8TIuutIWZmTgztEVQ7GHC8H51SseP8ut7HN
IB9pufnPA5DZ4KYyUpxWH12vS/hzoAXIN8WcT2TCgtcHFsV+7GcM85vX/TSRUBNT
dVyd1ITdOC1X1+So6QCh6d9EzWrQajt9DPGWtBeyKW9DEVP4wLGZgtH2drK+hbgs
5TiThezIOK+W1vTCMAgzWLyQIE0pTHsyp72QH1Q5UZ0LYiGVSTFYoZrUCeQ4FHlx
NKj7gG5am55znqCFU+T2XC5NYZycbR3dipRovZzIPtn3y8IOVKkivR4o0OYd7e4W
u1Y68sSWfgn5zQ+M42XkUFNJzzI5Cm/U+keg7ttvuwShDnqQb/vbUbKidImSzG4l
f4TvrB95RmIh1a8K3iuiEQajNLU3CjWpsXbSWnL3m18M35pBGdLVG1yd0wwwyfzC
o5PWxnYnnCu2SX8CoetJiL+58OHQLSpl/yvAKE1jmGU8UXvsNmjjZls/C4O+fiSk
Qouxp41MgKrqilJFww3Los40xoTdO19Z3rql+QD+mbCiE5kMidYw8D4ZfRZJkCNz
csutX6c76t49owm6RTlQn7V52lA0VwWC2pou7+UCczQ/nXiE9qI+7+uhFAThR6Ql
5yLm01M/HcOmhgEeQOYR2ECG18ZY+Ppy7H7JipvfXfmuRfbnQNcACYYDSK91Av7C
bPKbcQyO4xv7QlCKWNPHonc9zB96qsdnx6dAs6Eaxtxo9O0WISMWUqB79HnEDxpi
Wrg7aoFRAndBHuOUutkw4WVlTr/GmdE5LXBOw3u0Uxj4IXJtJNHobkGqPg0TwmGP
wfbc1WKRheiEvffWIO88LgkJ/N+Uwy7rGYSw9EVyRKprKajJVVSxCEMWwOOKqXdg
sIjhU1mN+mAyh1rzAXLhBDUSb4MfjDAkk12cFCWJyr0Itb8jIzGK+H1ZBsz6wkXS
6A13S/9C3zA3IHZ/K8M4BbiU472GFjTNJBjUBz5xBacjtkrYtaofK1naKaGk6gIW
OO1cFaGj/Y1W4SeqRoBE9Yuuwq2qryx0XsYWOqGpFytdbV4JpFKgy/3WDmPlTYO8
O4L88B2HaMeSI7Io+vrKf20d3r6OEwE3xk3M6MdX3YY6jwoplgH0rJ7NBqcoK9xH
f3id7OnmozIzKOG1bD5+dMjqrbUZ5GdujOpTR10PE+yB7hSO0OZ/8w5LkiEjuYl2
rJC2ZefZ7Bf9gtmuAgCiPBOb9l1EcVQLLGrjV4M2w6roDKHOYzFZSqyXap+VfMme
X96Rp0vW/ZbVqVsOTEtOYjvTE19cbAMdsuesBPy/ylZJ763JckDBkwKJuVHK+oYt
qU5xWLq9VNgLMl1zffmXfzd1Bi/gKvUGXvQJNS47aPUiERgpmhEvfpkwE6YH22fB
WUogh4DMD+MU232DyzgaVlFrjRKEY7XZ6RKSvW1uCPq+4EmilbR/sKh56smSZLZR
l/LaS2mAtz4Wk95/iisZ5j1YlPfAkCOu9bOmM4IjxH9MtRDRWABNF+fJFrkA+UVp
3+p6IljgsjjA54WZ8Hu32zVNOJvxiVMfILzO1jtsHfE23ou6Os5Uv/Qf4wfZxU5H
shaa5Pbb9O2DTKlSsOgu0w9C/mEp3HFiAzq6UzeD37SosKmcP/UTW2wNlkFxcrL+
cqulM3j6q2zDy/iSbzTIiOmV//EnkBDsSNhG2CIm3snhZJ4HBGk0PPlQyVGIGbcH
2V4tTHBDmGdsMGzuX/e3pg1pM19ZimakRkPIl0rqE6Ov6X7oXGGdYOJH/x34qNgJ
LhOVeOUd4geHUUt8thq0HJKvn2psaIMcOma4yyAfNlp/j9uaInVwCsJYopvD0VfP
bg828adcXt9Rg5pspa0Spgn3rTzTeRvR2mZ6qqBsu9XyH3sL8CppeDUDPa/pyIPT
Tnf0okYDm2NegN0WcU7SBaFm2mPvOilSl7kLgIVjafNt5HbWCia5v+zht9MWtr6B
QO5TWaXbWey1zsEW+gR3CC/h/VD45qVK8WCyejo+YmfeLhN9Wu7CA1TidO30HM3f
BPz413mSW0senHT6z8bTmId5U6udGsp+t7ULu6fsmK86hGXajAWiDcmBITp6adta
aAsznfciwddPjaY6f9fksnGRHyLriyoyw+e/KjlCnZdNi0mJx8R7RG+YY/mGBmlu
MA+IjYof/b30b2l11/tX1p9kwTgjSi69l9hWgvuAMb8WqpY6ACEuQT6kqAUdVfTF
2wPm5wc4aJqVUuqCCNetSpa9qHzdjyglxlafb4ji/IEmt7wQ7oYivp2MjrwshtG3
wuPGLMK7OdE2fXrx3Avcp5+5oa/BOTCgAuAOksrVjAT+bQ7ieDkzGoMJe556OE7U
Hk76gnl929n6HBLOgBh3P7X/wq3aymXWMfIUb5PbsJnnGoz1ztWGT7vhIPE2sGZ4
Q22SnrWQZBAMqoKWg9yB7FADy/Qr63ARKLFe7PW7GxkYHfHPI8hJrjlGEYAbgPgE
RppHFEI1CW9LwOU8rBOuZfhE4wiUQ/oP2+Ledk7a9bTPrZaJltfHo8yx7LbdtxFC
YWJUWPH4g7ZlBtd2fv0xHfR/X7PqxU/NR01Zm+Dvf/mm9b8obO+pKZ8BQljTRvWW
qifvaLKo5R1auADiLP74HYOVofAuznnrfhKTHd7JM3xpzcbewf/uFscxV0/HCihE
1lI8/Jjryoi9wxIy9OFQSmovu1QNGnNV2hIB2AA0YO+9WPV8m7wQ44ualrlwlFe6
oM5e37rm4LCkcfOSuLii3BjNqr7bxZaEQKFW/cdwXmCu/PBsfXh3mH/c1q4oIorf
/nwqttzh6QWt8xsz8XBSntjD9+GgR/RHz9qYJxRgaxZ4xbjvVH2zEWTLHsfcd6u5
aAjUC2jZKHPhnXHsxdI3hEstuHpgqkWmdMMaUvPjZ/7wKa1qoC/By89pCBW7Xhw4
7dkLE7dsPx8777aNXwDzx1/jczLefSwkMImwy8nChH6J353bDKfqdC8h5n1zTEnt
siG+XSXN+4D9kTt2DrHCpKutUMPVslE/d+Nvy9YS3yQS65IBft8k44ZNMFftG8nB
hthSYtpFbDXcj7jCjjpMf0IycuvcNywin+pUR6ftfJp+Dh+Ywl0fekv3zCmj1M3E
RwE78niwOC9k9B00BfCLPgndyp2UWp0PslImP0/Dc10xZaP0tjj191bCGDUfL2xT
Oz+JJkXtbtYxU4nsP33Ha38fZvy5bzdAsetSszcpoYh4UZUymAfz4rijtlAll28w
KXY/qylFeCHfVIY45wM8VdUoPuYVmBXsSmFvpVoczlta4LPT3nnrd6DBiB/B46sm
cdLOwTiX2djaHon11slha979mMO9wv7DGhhyt6SrFQPtIQnWDuQZ7jc3A6VhNDfb
B3l2AnufGk4RGIpQ5aLX3WL9YsJEoTyvTD1Jut+/XbjStyT+fMp7pcGjuM9B73ug
GKVY4IhPG9mXXyr0j/qz/zvjZZR14f4fWxIJVMT6sNDiPBWPkqVFoMwyZ/u/cI+j
Az7+UFoTKArnCNdzR7b2/DSDUxImXu/T2ldAP1J/3G0yEBy4PC6CplWE3P3MN8wK
vnJ9GcjgrBvJ/5clls8na6NfPEy0yr2V4JKbqRckNO70hS1Kff8Q8maU15WkB4QY
oVvBH87c+gj9/q/KYcvNsmrRzTNsgjWtVftHHF8zzaAeEMw70EGQ9mjzwhn7szcY
jq1t0vvkfYsMk86s10M+TbcUOs5/wN5xpFDq8xtmLsz5Hby3PfBvdKrpmCwSIbjK
8x0k82oRutPC3859ZwcPok++e8gdd4+wjJG+k96ZJxy2KJglZPyOcTFWbEJrZZHZ
xLb3tjrbpMPH096WXCXrx+itEQ9afIZWkoWJF0petVBgsRmXnQRPGlQtLgC8NXtU
IN52t4uGWCUwvuiEr5K97vWEu/lBMnqoDYx5IboBRF5yyTb/WWjUSkl5WUPkb/cD
SXtU3d2hM+5Qq4DVNXS86f6Enhr0DrAwHnx/izLXhgahOt6sXU/vTrxp+bIX+ihF
Amv5QtiuYFlbzqYSn1W+XlHyVuDSSWRQFMkYnGOj06fJ9R5R1aSoh7fhspj7yTdx
OLQ/exTdwrjl13tz41blLybUdNSlaGjWN7zvvFy3dDjkCJnSxLQIMEPLHt7BvG2T
tSJr6mg5HnzNCgiV1UaCozrEVvJIMabcqKGnyIEg0PfN5f72AFRmyEjayKF5bgCi
PHeYuvCkgDQ4fEf5vywfFY1hr9tlVxXaubcPoz8lMeQ+fQRpfxNYBaHRiCibUn7J
HJWjC9NRwbchcAi0zrwWJtZHB0tLj2QNCHIDGzq691bSlj3g4yRG6VxPxJSfik6r
aeACKbG77F3/Pf4crLKT4HQv2kFAThL4+kPHtoa6JrEvxro3FdxOUhd/A0mFWN55
dd9lBFGQNnl5mH0CG7PXiXE0Mm4mYHQ0QMFzbESeYndxAhv7NwniuoLfP5Ad83wN
Cbq16/e8LzELNSoq582g7L6doy3wZxNhkNRnWY5PplAHX4XYc1NDnaFBgScrbyQw
UJrqBobuHyMzwfEeJmWWNJ/cJdkV+jH4lXAQ23ykyQTSDWL6bUqfy9cLo7xyiqmv
EYV0aLFwcfxvwQBqnqMGGuqzeuq7F9ecfBcwAS+APLzOf6vxYPg+KVRdRqTnmC+F
EgyRng7GQkdJjv4oEzxGV67Ck5dhaHS0Iauye+g/KM8wX9n60TreslDMIaG8MCVq
NI1gDanAhOeEgLLnUv7ZsMkMfh3g4NqNprcDrMue2YzdjAMsYyyX1RcHTcJvJeMp
R8AmkAhc5logucJHtEHN1cLwhA9UAObOU9oEwa23jf2GlBKY3TXmyfmLBk7sojjm
vrNUBpDoDjcrlGjVOlfYpdTY6sbTgBo+CSSOJMVLNgTqjn8kafD1cvBzL0IptuGH
JWdqRLRdXqyAk3BNYH/m/ziM2uAyacmex4x+oluZKbhtAUI4YJnuYXgxcnJDfKck
CkLhlGM0xxTHt0Q/+a5zfCeHxGtQvyzgi6YyjFNWyxnSbNh0KQDsy4O797Ao7z39
E591tdmb6262JmtaUVxMx2p/8SJKZgymNFKjQ6Au1JvBPmt3SIQQxUps27D/VWfu
K4j+tl3ilyLPEPfoRVZpdp9JH3FYVmDREl1MsJPRZwyD+0ul8PTCSxjUqepxtzP6
C1Lh/w4Luc3qaJZjYco2Gs071gvm4SHmySnbNGxLxZiD7yH9NL98zA8PoHlu9xFw
GnkhnvYuYGOOh89YaaRMd5sftQJ4JB+ytg4uk9pyX14zM2FKf3aO5xoHx4uDpJ/4
KymTDcrKjQms6JAPnZGrrorg7Y4TVuYirnEe7BpgvClK5OReWyi7ZfVun+lBC5KU
JWFLVm+bx2UMZILIphIo2gUqgcNW3GPLzFyj6dj936UDuROGjBwZJnFcfYNhihRl
xuF87qRFp+3HB6+SRwjmn6/hrzo99FjxqE6k607vDufdUSdlV9kBxJyCyislmYXa
3SFRCt96eU2tij/bLTJ8m98FxPCpiQe/9VcF5VicTeZUz/aJoTMAzTwJMkR/Tn6N
UT0QWsle6JphXB3W3cqXkyEPORpj8D74KOP16Vv4EDrRzDI9ulRRgzMhABrlfUGj
wIwyaNSdcliLViIlBOShLcnm5KoRb1IysTH/GjZ66u3Gn76feEa6Nv+ncxtSMiTN
O7Tx4maLgRb4vAaLiMfmvl/yK3hA7rUyvfT9P5SYfRaJNG521zNK0Mxgy2dL+KcW
PN91oYfFHsd+rWa1GjWrxSn09qHE8vXr/FuqaqzDFmAGpnb865iXYdwVtOK2lmks
Piu9ANiVYu5UfeyHPuIh5DiZxTW02snJwgCZl9dYbYP4mwI0NWMggLeRDh2vEPsJ
0MJHauGu8t6K2sLs8lAl1gu0Cg/yajkVe8tPuo3VERxb/DRvXT5VRNpCSQP1wWVk
gTKb/RFm15tRzihnDfc9c6e5cTr85TpiGBOmOIiDkl/AVDSsO9hRDCZe5FIthPlh
mWcFJu8lAH4nhz4/3U8rTHYgdzOw8/vgtNF0MmopGBb5FHXgh4OeNvRcZxC3yko2
vfogszP7PnzDfTHEQaByzdMCI0dAxjP7RJtVqp4AvYvfZ+Oyo7VmCVCqNSbUVF2J
GnH0LAyCmY/iygvm+BvBh9rj+O8rmH8rIeq49YN9UDmIq3erByHftgUKyRvRX2Kw
qFreMtJlriyAapP1G/IZoyRCnzZxyUyurj7iFFKGR1CTZdfhL5EYjBCT+RlKELXL
wTOqbcBDKt5wtvtlFzmQ6sR8/Gqykn3LJvrpxpX/a6Btu3Mo5/fPd176qEgZe1AI
9rRKcq85udclvBgMtDpRiMYIllpMoaixEbSikS7rzIUYab+Z6gdFf8lm82H3R638
TFMsQaLik3nJqNmS94WGgbtE43FFrVp7MnfDxcIVVmvSwYwFL/djIZ4nKbp3/1oC
4/wHFT1nPj9zIlmsWLbVTSHR5OVR4Wd+UZ3mN8M4ZNuJP0yNkbLItXakjZhTa8EH
V7/Hwt6FDjulDsIAddoQQf1SbbjtJPxsN/6LvVNGf63pZdyHHNK8Z1NFQhzmAkDS
nhdI6P24BrZ7AJCuYuZiuveCanMUG62QfE2SYQqVoCLjDZcPF6XnXJ0ZsC+67kg9
+J4YWqpSAUsLmjo2OcKy7UbzfQyd5E2y+OkZt3/NRVmXnFkRC/aQk5J/utYOKUj8
vNQbItf1BDUMfVlr8Js58bVZfFqU6BUya0mDPSgf3VUM73Sy0Ah+QkaVuHQbPwnd
d/S3+ofzu44p5fckwS93f3RXLd1QNdwDl7xfMh/P8XpDajH8DkjsuTqc0BQRGs6b
MzmHU1txFMnmj9A22XrNBdLhc1IuLgx2rI//B3MU7l747sG5nvjAtB6xXtTbvGPT
Xbq2s33wW7wXa9te4aUZUWzicfM33vIVNVkRPEP33rUGPTgiZxLMxEV3yuIdp2rq
c44Yr5FrM8PuvlflMyivodDe8PTJNP+t/v6FvhTldU8OIpzu9cb5MO0YB8yOX8eT
4/3sOJBIVezNk+YKQa7p10+3ljhQFsd3rgGIG6icuvaUSV70dbiDRNnCs4A5iZ5Z
lfPIE8fKtXqzefddufrCBpjldGkeIXQlXjZKj9y7fmQBRc7+3rNrspQ7mqIjXQga
M1vSke9haLoFka0vCIIVyWP1oXFB/lh+iPjeUs2OFyatr6CQR/Vi3dmldJmRBgk/
G1s7UfFcq3Hxt8ZIt7xFAvpQX5w9S7AytDbw++B0LeA+ml0MDw3M1mxccTJQwJzI
6ixn9mIamnM/3tQ+fg0taD/xArWoTaWn9ELuY3fsYmjHSAx0f7j5TXT2MV2FbhuK
keb6t+rAKVo6RzHDOi2TIrrQSR0fmwWidM+7W1nqrP1B9c60zh8gliOwgP7OSEl7
A6AgNaD228ZN1zAFLlqbu6tsYHMy113yVPBxb7n56mSd+gTWKrIaDmuzkVAXQYVV
PMFtr/WwrC26qzwIkOBVmK9CQA54dvjr6yWthD6Nk0+jMNCMaKCRiLAykXHp2z1N
9hiNmw9GbtGLOmnCy1E/OEhY9bt6pxV/GbnzMvOc7PCoFjG/0YzkRLKcls+AyCu8
lPAGKwGGY5n5VQIQaZfXQPYPoDANspEltK7/tgIlX02BPYs3JpPe/TfJtrAUfoAP
Af6Q0E3mNvZTEOq1Dqu6ZhjBtdnTf1WFv1JuOmsCGpcJoi7n6aR0koN5BjFUIOUN
UFFW9Z5YwJAzTCFvJJpFHPEwZzLeiflQH4eQQAuDV5d7PNrtp3mtRtCGu1VV/kjT
0Ro6EmpbJWtbW2dCzYvwRU8l2K9T/vJIZuyU/ZUujG/+HN1PhZ1vUg0DDPlfxQBj
YyqyYOrOWEQU2Jm2BvK2O1t90UPsyRreAwXDx+gKpGPL15I8uV9VueRbBYqY95zc
MYtnmYSh/jfg8Zey9lARKc4O6i4X9Tm4QpX5MfLqJIJ7vplnakWe/SV5AkCicaUD
PxU7j1lUrpAZzjFdAm5GpHiHb5YlT9VQXux5cycvDoJwiC23hLgM3oI6ZJ1lNgoQ
ugTYJR9WJLvN7TP4HnLbzbdiKsPlMr+EQoQW9siBkZrC3h1xKFsQ8xsS/zcltIPi
OpsqsQyeF2Bpw0N96P/nhCAcZyHrDpXEfvarCMORnwBnHvDd559RL72MFuILBKRT
DlgoK9xORzYyzqjbmH8h0qvfA8qKI+pIT+eE9s/Nic1PEbyBuCk3POAlfbKu6yYK
VeQAnKNoStujC05+5Q152e4zxgvgplPX9jaUXL/sD1yzhOFlXbxLkshx9kk7V+Ei
fIN5+gL/9IJ6V9LTMitR/uCT8KHnuR2M4rHy4zSr+7osS1PCilj8VeWvxS05BP3j
14H8Bi50vPOWLBghVdleh9ih2iyUMkOGSSw1fyr8uh04ajE8/tn4974LktRj7aFb
OZS1ZdCKKPs+qfPQgQ8g4NojwgdKFMxxc+Jt9bd+R0POllB2OFgDeWsYaL4FYXke
iaoEKHk0LVRg9e1KACgtSMyjQe2CISeCy81sHBmOx9D4ZunIjtQu2EOSaStqKbTv
67Zm8NYRpGjfIB2nqRLEAetDSxpFi1bnQWmv2IldnM67BEDxe3CfgN3ziyChMjxU
wLmn3e3/j3Ij7S8Y6h6KLzQbXdObHnQ+grtcGjtI5UaneGb0oaOlbw00h/kjpP7J
rVknaAaotf9BTqRNjVJnPPOl1kuLcpKao3iCGGMTFg3dczgOd69W6i7NZ7QMcGNM
D3PAGhk/PA6mg/pwhqWBVWApDxLZcrTBul8rxzV98D9kskVZsbcOfp1pFwV3It3k
vg6j8X+G2vOT1AFCoUivPl1ZWZ4hMcb3hfDUH26/4ZuXZ5MKK6SM2R8ddNWxVzJp
o8uBfv1ruFZMu6xqCTCaxgF6VHszag8JVLkbKXn9MhIIWkhIBuJ5jOcCAe09xnh2
0ypSUe3bOs8eZ9IQa+WBAhMejCNLu7OsMFhNSYqTVyTnsGhkc0tXQJh9wvuy8Iyt
Db5nvx+ba52oskydu51tI/ybU+m4Lk9wznnZTXp8KB4X70qW67niOwvH8DJqbJRU
WejSkVC946pX4UzZiL4VvWlaWycWls5Tqh2BzcAjV87V1fpWI2a4isSNNgF3L7OV
MCGQE9zgGccFT8lykYphGN8CB+oVlwjeNJjp316T/X+MUoIwceKPN0OkR9L23Qlq
Ve3P1jPDK4DvQF9Hxk6EwGOrQrH7ozD/63rSQ1MtNxI60MG499OW3CKzjeSvu9fF
mff2uB788OIjarE6a3NeuRaUJ+QMBY7cN6QNTWtBzilNuevUDTQp6I3KMJuEMLph
jJfm+/4/IVI/miZVQMbMIJkmr6229v1U2VlBNw5zWb35p462PyUUp0pJVBvZ237d
InruWlVfUkrDXr+CqExOshW0KU5tTq1bbvjw2nviHxUGK/BLH9eKQaLIZ16r7s3P
F+uJyzB1MMlQvy+GrvR+4Wjm6ipz3xwtI0tkJpCeAhr9dNzh1Foz+AC/grmxC3D4
+6pjSiUIalwyWulXaaj4lcjFyPH7zPi7Tsn5BRna+zpu+PJYylv4pAh4RgACU8Qf
RCCRmUjw4dEB14bsIq22Kfs7feKIZBDvF964Www8YPIroI2eDkiRa9Mxx1maU9lB
tPRz5JSwaYxrA46zCeBiHeJkKJZ9qHOYg5bfEgjxNOr+szZl6W5A+mrveUpzNG4C
mnwDcCD/9P/jnr2o1mA6eRrWIhqSirmf7aGokzJveeT3fJjrnb/wHU5y0JvuNmYv
xBSmL81ObOlsR0T+rO7lzP+3UOqjAw+11fPFuGXIpe+t/5S6qu/EDMBuTcN4nexs
Bx7kACE303k+QFknKvUIGYfK5GQtly5PtOIoKc9VFyHKkbBYINIluIcaXSxTWqpB
m5Z1gJVQI/hp4US+orMcIW8IRxSUU1IFsEdFKFIZlvXeMcALkWMr0KGqS3ha6waN
WQcKY8+9T6Dv4SQtkM0unuNtMQFsrtE7pIxCtMv/eC63F43xijCVX2TZWt31dWPi
BuXjHgU986KlbmUvKw65TfcAIbD0JJLNHZ0vyOZAYtMsRnqNvIrE45fP9MQkZKgD
9fJbkvGm1Uof996/Pp45WAhTRwRXUmbeFXc8JvHJeF+7Yzd9SGay+O+8HPN/zuHt
9ZYZ+AYrc8hTIZYum149OyohM/GNyM3QnN86pFH3bnEPLC0wvGtYN7dBu+awYjah
+787ExxSc4unuk1ZVWftAGGm0NypF5xeTiPSczFBNXqneT3vGdN+v3ezOb6XhPP6
Q+Z2lOirIFCe28hhxDoXnKp4AoTvwI5CWQfveOXtB+wEwaGYFeYYN7WSgjOCQq5c
h4zSEfDampR1mnxaW1o9c8KepSybm4cODOK3sO8/DorQyaJBbTIkW+IZalGMD6QY
TbnAvOBUry7HsK7qK6lqGNJo7H+GLF24o3U9SEeonEiUbKMiwYEw9FRHUvFKStT/
1QyGflxgrgD8PhY3Nn0ObqqzXp6yKzLzY1+68IlZohOjTyF6QaffrTkdloyGPex2
rsdy5rw7mL4Bte7YPIFmFIQxUU1ayznZ++OogNmRHJIPv5Up6kglFxXgTcm3hCdS
5GU9mn1dmTNcNWFagMucGodKQYk8lyd6Y3hcqMt46QJx0zvUc9dWHIFOra+K+AG0
4+iuqnVYRD/+tUR2MpyL75JgBkFUwbUTMgcFVJK1B2vb9b5pyCaYkmp+R2Eec9Pv
XnlNaySQJxPCaVbF/sH5VQTqtXAU1sr4phoFEBPN/39DRm3Zb27TniUZBB0/Y5fc
JrxBUKhhw4De3hwUtRSHOe3t/BLir1XWkP/XwpSlK/O0Oo9HRLuzOWnVXOfDVbV6
NDDRcYah47BwOeyDjAWu0AwOmjJPnfhuNRZW2aS01NER2C1msVG0h/S4hB5RiFo0
847wxaJbbsIchcHQA9XXVcwgQhTgObcwvzB5wKN/Y6UW/U31p8LBD6uwsrLIlo/Y
ysfvd2+1wwbIV3zDLsBGQopv3HcnD2AAG8W+Rm9OEK6wqPyJtBP87EUfGVR+8rk5
Cyi3cbbcUEj1ltEaSUaNJmZvZHsHWKDRMm6cGF36eBAe5ugbW3o7O424bTSA+vfN
ktUlggkEVR7BeLKJctX79Z0uvVQerYrCnvJkuwZrYaYNW8gtoYo1SMqvuew9jB9I
m7nHvdv9MzdPrM7FZixRLSpv87mUCUAo7mmjZ2qBAL8E2m3K1Bfva4RMvCLbVPKJ
sjWpS9DvZRlQ6IaqGpvmGtpr92IUhY+ghJC0DKg0O0mBgiqYQbWLLJVQil7kCKVQ
gksnbZbBo0Z02qcv2E6fC+LFk29rNGx4B547P4zftTbFJGvEogVw/wOJ5vuvQmnp
BZV7CasfIigHV+iGuCH7bv7kWppA61WUNL37//6YoX507sh/66AvU6KLXKdJhuYw
9MuaAQXjkwy0XWqUz5TcoNvfauO07NvHad5bAYQlAiAZFhJpDt3jwbyDKaf5po2z
3fExTzBcoTODxefOF3gMw6PqxUL/wtRhgAP9b9e8NrKaxnwMrQS7bCwil8cN38WE
hWz8A7YHXgNXfzCkAEdUSZ4vKhmN5QI4VVxnQIxHfsa/a5lr9oN/hCH2xJaiS9DS
hrbkiFWVCcN4kWPGWIBZrJ9UaiaSYPNSIekxksGwsxcOYwH/UJEUwjwx0Uf12vM0
WPBbL2KFkducERiOE1lcgulpMBiwG0kRgGRj8fLA5opXC06iCjOlLx7esSTOtT+u
pqDDlP0Rtj22TTYKOTNZOZQLhNBLXvGD3sKzrsAD/x5lcuUZUrNeNCn4xr+bARJ6
B2ycYhg6Ew5TNpc1KyqCtODiCQg3hb3k1Cwv/eAKbkbhuqFg9Pc2yj1CYzgFsEwF
1ysd6gZ2DdJSZ1ztw5xPW5AQlNdou7KwMDN3XVtR9XjBxByY03nMVPgTuWReA72c
dhs++P6kX8lzOaRNb7+VM0Zc1dDjSzF7Q5OJu10GnFi1m3AW9KWmvpbSvHrE+jib
BnL45DYaAHbexXYnDSBenj1oRpbz6xMl2HA/XxeuKJYNBDdJLLhYWLSkgTNORnbf
Wr4LkMX1MI6xzrg472/WcqFhKLhADba02bOL4qlyCs+Shi7qi7hx7F8bo/6EKlCV
0RUQXAwEhcmWkIzUrgU02v1ay6GzP5zPuRpSbiVX5y+LvRGmNlwg6vz6S1QjMKpo
VwdzEsmCngZokTxr9k4PTnQSyJ3WikidzpWFv478a8RjaiQ/HMVjT1fp9J5FT9nx
k/2iOeM8U0z6CMNG0kcPWrxNLSYyvUFJy/ck2AFRYHrJpKdPu7AOCOyn+Iz42FPf
3Ruo/Bj/Uhb344xhV0eu4KbhGuyT0tLdZNfaF1gjvtF5IP6ygUq82QVo9uU9YrlZ
yK3JxcLJ3YldKwrcbB/Pct15mUO2l+DN/kNPIcZkVgg7FM/ZrwzPfSk6eAmP4Sle
zJmwiZDAU2603OcTtcOLOp6pEQ0LweTohu48cyT6wYPd4daO+e8EcP56ecpd6y6I
p0AxrSSoXbSB/vd6g/kGTqKiRxyJwbMTvcUYXZP5VR6YFeH6qcYVH22oyfFrcO4L
7IeAU5dnEyn+mHLNSoavzOalBtAuw/AlQLBtDSLLp9SwSJ292jCdmWeo0VQ59MLK
ivzbJw+h5Rlq9fM+UXldsvvKPtIKb6nVjC5Zt4TziBhL14QggXQWC9HNc/9m9tRQ
p2EduXHSQWgTmuwBxoTqWvZVI+OctYaP2h6NTNgO4UxRla11oPf66WagPFkcsGTh
YbN40+Gp///EUA8/E8Mj3JxWSVKyvzvhwM+kkp+edAEFyetPvVbHFt9Cig0P37eu
7FFBUMehI90m3OzsKXq/UhkmHbq56rBsqShex2ZqsbcLHpp02JvUDleETvDkKpIK
CaYIJUWhTMnrQ94eht/+PdI6mpFalDsUQwjdpz74qtooqVpcoVxqiYF+dmnBOEP9
xn3vSJYAAajed5iushft8X4E8bwU9m1tlNP8e3qt5Ks5LQZ6n/svCVyz6/uug7c/
rCS7JzMWiVJE5zeAH1l1TL5W4+7XveTJ10m7J8H0G1YqZ1fgtFwvw0AtmJvW8dqu
k+3A5V/v4udz6oGJ6ZPNGWG6z/3IPJk/CtEHsSly3rrtpHLXcgRXr6LxRbCDimvw
MkuJGxN8QEL+nSDzmXyiZ253uP4B3tl9seACKNvG6NxftYcb7kL9SVCUb/eN7uWZ
QV6/DTSXHeavuDHe2zkF0h9KC1Ir6INcgF1ON3/doVUhL80cy5FyzBizEVBCillA
nD2hVwWwKCQLXDO2qGbKDBT7pVZD+zxNS6EPeUwFwIyruL4dHQOQes4e5m/Li4R2
+N9Nhqj5mZmurCUhrd72jmMT6KdNK/lQnjG2TZdjVdzIGSEC3ocosoiPdIiHCGU/
TBe03XD1tsQ2r27yzcEDgfy85oc3PfYAMwPLkTOnTPe73tKh7hcPCp08ZNZxRjGQ
Gy1iOGOSl6Blz/IN/ZyUCh/2XBfXloz6Ac9lsGHALGokuaU0UNbRvK8cgQbG102D
2Z1Ep2W+TVv5HueK4/ntF+DQxVF4+C1MNoiXJaG81+SRAk1PEXdvPamWGzr2ww+N
mZjoyr/M3LkdbiJ70HgjjrMVRPqgSo3tsUz0fHYmukYbr4OfUffzzJQiIEMWEnn4
06Qv/tzyqrEa2B2wborFK4DSJMcShu/0Q/nmhKa17XIBlm1R8mI+ReWcxFWIy+SE
xfbPuMNLmmdMtx9NfQJ9DSRWo/IshLj2wld5V3RUntkK/kO5N5mneIwTSGOPkmeF
rBs3KcG++9YLfz4emkKcpF/rsidDfsqM5HVwBPMoe8FuqyLc6NmSi8eaWLEJxeG7
L//4BRRrddcmk8IC8psx0OMHrBbmbyoozS+8bXPf1TC0SFHAeDNHanYmSzQc+Ar4
qMZTqHkgNI3mExA1T+pxCYHMkOC1FxQF4HLaYnxSHusQWnTiWWIQz634tNeMbdZb
QAbNeh5xZCNIBv25aml89LP/xcuOgoiZwuhrfGva9Rccp3p7NcdcQbWy+8BmiP7X
zRfh672kt8ODBDlZFmfizj5fzSzWfB6xr1dqY4nUEDaKBVYay4TnQ4TU45uYYHXi
Pa+FkESu7ksDHnfUScuMyN5Kq7yTvg1limnuQtAl8f0gS1BCSmdPcp5/UfTwEIkZ
+Muss4bFX4zLsaLQCwaSKyxjwdCLfzrA86pqhiu7H6pICkZLwz8EAP1eHvu90P66
vlRNNbD5LDSg964DPSH1sLJswce5mmuGrBENQOyt4Vw1aT5SOlZ3+I1iNaSZ4grb
xNSw1HRHp5XzqwwkVdQnyHwbKXLGs2JFhkhJU/i4S5jwmNGmgNqWvc/uPIzy8YGP
8VtrKyrXrHAMwtNyCWZcP8WpoxyLARvmZVrELCzc5AlRxMri7tmo+WVVh5JsVAk9
w5Ls6oIbnxDbbbC0wIABnlR0gVLJ6QOYIVbHH3XheOwajazxbuYoPmI7HeZh4my3
M9OGIrokneUPIdZfICAM+jLgVDV/NroGq6bar7qrvLrdD3HtNJPXycw2YBt+pC2f
IKSMaRZetaR8zFWYjJVw/MWZbEOBIJD6EMOEHkz6Ql5Xp7sSMcYAT+w7Z2KFX658
eohOXw3fJmfAERfyYqfahJpEZaWnk+8BHqQ+VuzXjwIl9cNLiyXewAo+Qp9lSEoY
hW09NiIR0hd9XV40vw1Y9AtIoVJdtimGBj87FjCX/OX8y/7GnHPwFjNJ7nZ20pHI
IPPhRanjgc+CzDKwdX9GqTrGZW+pTJhNGJAruKsks5Qjza3mRFJk69gHRQxzFGcQ
skYj0R6FKlQpZ3z/JiwMNoyBu13IxNemkGPzH5uLVya1x7mL3NZD8yJNjJAq7UUi
f9jQNoj0jvTvunmr8Sf97GMkaXT2AxHB2tbx2mVs5Bm5j99O4+prtmXGWbWBPvY6
4mwdLxzkzMki0VU5Vd+SuWY2XPNWGLEc1kE5IMYELUyVvH/ar8G+kiij99GmMatO
vawvhjwWlXCGK7UF/FKUFXOS70n80EwqqFzkIoiH9ERspXhJAn0uZqGbA6364LlQ
LXnnf+HFfpTZ7n4VbR29rOL5y/QviQDglOpPm7rug8ppnhOiSYF39Ug+bvkzqCYE
SUJecN8dv1HrJIVziGKw6EQ2YGI+nyGposYtkm37RcL9zn3gF+4TYNFEZYMt5D4w
4njnDG5NRcSkckB33ZLmNGk63+ZJhW7+vY9gVHm316dpOlf5SXB9/NBby+mu/Aay
qGc7lbyCLyl4UmvQm1/qV0dGvUmyorGh4Oe/R/VHfzcz+tISfcBKi0P3URFebi47
Hig8SCBBOPFYj+JaYn8hZ3Fpt82gZmz8DBZneDpjfS8ji77PWP3v0NXICliFJ2pR
4EucSR6pmZWTDGL1x9JxJ4N54tH2uWkTILhRpiBsuu3d3M8IqJ3lEbGQJY0nZeIv
556VSJbPSqLZgywVJm3P2zxCeQ4pEWaA4xTF/1aA+a5mTdKY7i/XVL+fsx6pnd76
a1JHovRuCQBhNpXRcI44/d5IDNOQbQg02pN8HnTi8BKXy4I5oUa9r8s8lj+lGJic
iWNsC79UIrQxGN6CE3fk+BOrNOv0Cn0Nl+SIKj0IgPJTl3ODGhBZI9NG5FGMjXza
HKvfCXskUr9BOjIvESWrz8J/DZTqI1tbTAqhSdrJoyF7HYv31w7xo5sEtqayJCTA
OG05NPULZtEOoJuIqz+MW+4/0TahHuzkhbEXdCVSmc1mXldOrOMipnbkdtl3ArAx
GibMkAOqrn6ZW0NfAUrwibV2L8NiftNNRBbQIvK/A8Wd8Q5fGLie0TeuhLrnWHU5
WI+gX1wabuzfkNQIC9CmUdvTrnJIY6QSwaqt7fllMu2EJB+63+aUT0FJR8e9rtJj
zyk5iUo9qRCOvrz51dfXDfjEK7f/+RhwSYqKJXOJj+Ma4EeeNBK/jmR8QAEMbP3U
3L+xtB7sUaPqMSHDPB4rw1sUAF6zNZxrp5Pn6iJMZ+J+qRWJVPzwSTZ3XzJYfZum
ScFnpuBOo1oAU1A+KIubgnwrQy6DedjXRY/KHeShrEYBJNS47d6EdrGtTX3FTxpH
hYVEBs2MJmoyxO8d3eavY1bO1L9n5Cq3PXoKPSERkpUVZ+SMwIl+P3U7ahVDjjcK
Y8yOt7EwnkB6qgPMTiNmCSZCzvoGUyy8yKelJc0X0I1rDzKnwU1f8Xiu00eOkLOH
J8+lx8bu1HXbQvJERYybil30oFuyrDI/nR42qfdFoLrcAC64SyfV03oHQmIpLcWY
wSHJPw8khUeKMkFjP8LBEl5/pb1dTDsxYVheU+SE5icn5kcCh15GBLxwJI7u45bA
7a2KVP8V9YOg2VoJ32A5SNoQoZulQRj0yJCWdyvooQu0AfV5MjDJD0PgtqWE4e53
Lhm40Jyi7Vh9h/j4kEeuu8yRPtbFUpzqR3c5x/RCVb+pssgjenNprWoaioahL2XB
dr2TndqZ00uJx9vzZ28iGb++UtBHTnMfwUoZzky8BgfyjUwDymQD0TUup89lwsU5
zWEq8S2o3isHh81uG5BxZVZQqiweSvbFwYlWtpcgvLky8YEUdnZzVXXq6c5i/IJ2
g3c64trTfZ4wEG9kvtJ5UonJXpPAngtuUrqvXhtepM0mvdQRBuHywfHa81tqTjnY
7FS/7F9WnROsr7zCU4qhJSOsxkFiUVhJA37ZYCqHVtZiry0jdMnVQahbTD5HNfvP
1LIId1IeZWF8Zg2InUa24MkUZ1/UrpuK7Lev7q9JFgMIwlIalhbcJW6Ga5s5bBhZ
Txi64K0N/6rxoEaex7SjwvsD1JwbpUSJcfdm1vQYNtPZ32iiTfss5KiEg5M5vLpg
w/D69cneupJVi82oEa9dYUSAFD6t0Oe9Nrm0qCjseomYouKn0bBc40z4b2Gynjdp
JwAWlcLmCyy5d8G0RXOz+GSZfTU0EWpkcfEYjDoZebVBxYlkgWac+kzVKp8NYP0r
LbamVlUOAwBLrD6jyP4We+6rb+ooBoDyzMQKaPe0UCtv3CO7UYJpli2XvMDmiRbD
Xw1yAsS8mibsA46X34zZqjzWcWSMOGrQ6g54+DqbV7XYZVttznHh36N7r34ukcpq
SahoDa7RA47Q6TGsDcWchyNV0GSVLDRas+FpQyNKraplJgNjzj9h3xL9xFPTd1R2
F8v6zwgvEeuCbrIFDXkkgv7MoVh9xhCqaILKpj4PdDYBSpdD69GCDukmedujDsvd
Hjcv2npP+mgcaBJQX34D/SqphyUm5I8zEjmYdIcD43nn2OCa5GL37Dtu3WL3IEZG
ji4yOrudjfhBtR/NlxqlB+N+oPWGSBuy3/sELKrtzGlv2E+dteOtuUP1bZMGffsl
8ljZC6XeWhu7I807GR+Q4gZRu8DOT5j0sM+DcGBt1YENzdTcwkHSrREyVffGte50
9m9Ab/yGLY5ofNhLuxN5b08DJOvWaWccbdhIG85TRvhjvQRphARpGOyDD0L+sxxK
zpINITlhk6LJjUOjqq/7Bj7MHzK6teQlLmL8qraDc+wS8qpwnUzU+G10sfz2qXFO
xC+CFkHYYLNJ9QWCMR+KUx2ifm7uX5l6rN8ruH3ag5Cp8TrVwtAoeibLFz86iqVc
t8A8QYVf+3EKxw972BBAD6o4licn4yd0dDvb/n5jFJ4lOqILjFURFxyE1NJiXq50
RAnLGNuApgd55nfgrU4W0x1EPUozQ8V8BMuet+1fE5qOuJBLOQERslWurVAz/zsp
1Ubrq0MYbJYeL0B4Q0LnFvJzeQ3kMznZ8dSzglb9xlhP+5YlmSAc/38fOXLudVB2
KnFafef6rlNMuBOW0JalEoVuKWdinxMcgSPoWXUyPeLINvOqGRJagOy9tvawZa+J
mm02l9dgw9RSw7YdV5HVFhW0af0+lZW5KWMt+kzJvWufXt4k2t6wEnX8VchaZTe4
wBiKCdPAZBRSq+puAxFLhlPKilYPmStRIGp5Ox92B/aejXvQLG+MkJdX3MefuYXZ
duSl92Y2pJgySfkcy/Dd/QO1uYQH3xM3QxgEZwaj3eBgaZF3CkaAHLcVTMwTZBQK
Bh6hyujnguBvzixeav19z92GVevmB7nmqTGqdKOGmrivmrh/W6e8Nox5E8f1Tob7
s8G4h4JIShpKSOWXGwJ9v3kDV7zDQJJgeYKnnAW1Pd6re+54jByN4VU3w4TjYJlk
ohDwDpV1y81uNmi3BXDWP+IUV2geBs9hqeKWLsSOR3wowDK8zSVhmLd4Mddrbe4p
8oM1V8kXpC1mtu7DrMXubmm3GPfiVoG6NjbXdGmOautQteGEFoXFL/zXcOVxjr5j
DkyPe306yaWqUlvdXaChh+tzGLN/4/4LteUYGBSgKz5bgr21BNoaaIBAtu+vEbSt
rM6mTYcW0Wv5I6ApD7DUwnlG/B2lqU0HhqGOBIo+umw2PCNWlvL0CZB8TGqBrtMz
7jb6+tQ/SDyytsQqxPApWQTPg4esVibB1h9JUpFrW+EMlqybj6MxghvVn8Odr+0m
QYtJka2r0sLBEC5zCLeLkJ61uvX37yioGjazZfbxo1YU1jdMoqFf6z06VJkVwt9c
6lTywwH6xmk5B6nFpLg1CmzfiiQn6HINkFm7WH3oc0o1vjU+KZvhfv3JeGHy243l
arRHb2S3G7wEGpV/w7Bg957iEJe0DYjXolm9k1RnQT0vuEEOJixv3RaIfMPsdsUc
CAD/RcSZ837eWY9B4T3Y7Jt+ya5mq/3kX+keJ1doXRlcxwvaoLcuvtSnj8fccTdZ
ywS4+u0tmUt6QJ1hLJKR8qvS7e6wfaaIPk7DKz6mjcaptE/7rGjW2YNg1FJAzShk
ESOYAUf2cpyGscCZLuBMt5G/Dap4rNPzw4NHFmOFt44DMgaE39XkXL4EyUHKjpQl
MG7QADgNCfvfv4Le74uc36ohcRAxeVPXGm7HnUJIU9za836m6l68R5mtbSRFETaS
2iqQ56onfMc80p6m7M406Hvi6yMwyT1mexIBm1f7PMRSKQ/0jFBDe8A0xI9d83VK
nH0gbwu5zKOkaO0suxXCADIdzFUi0SK0DcT6cYCs8JBDC3AhSTgLcgqIwjr/TsZ2
ga6fDUsVSbLYSFQxiygIu8s4SMcJI9QcbSLLg4ZCcEYp+W0ikdmHSV/YfC8ml4HZ
gFqwtPz1PKgJFCkP+ArmH2A3Cta1DQ+fL4PJoNLwEvwEfVQi5OWvDBQZeluqHF+K
Ephlck8nXD30/l41FLPxfdisfczJp/rc/l9LoPVEiCKWIJyAlAlyUdo1iRZilN+N
P1enPqFxHag/QCfQnXoJf0KEX/IXADJTSkgHajVg1Pmsuu2av3124j8/3aKMUFD1
KxxH9aEU6X/iZchsHyPzrKTEiXVszTzUWlVyQ9I9J2/+oLfh5e9iPxhIL4k1dCfw
UflipmRmfOjHDuPcKmttyyPQKr0J7++rrxS7h0u7YwPMP1PHJTt6dUkh2VuG1LZ2
yMDF2UxSqENtEvEIeOWQ8LtJMF92qcS9OV7L/5+I0Dg9vd1go5JgrCktHRRtLeuy
meVxOX7B7e5cfyih4v56rCFG6i/WYCVno9FrDS1Se5/rk3HBPWccr6LF5oLFzemR
RTOdmbwRD6yrLr7fU+asUYXWx71GMTGgSRi9qZgE3U98lO8eta52NJDDzP4iI/VE
ydg3LNFU1qgR6TjB4NsN6XN/NNW3oSrJ4G3WXmTfxUClIgyggePwsfWw8i408yQE
7bLux/+k0LR3gdxWZ9KoRmiZAr8qnN3RZ2TvxU3KjXZB8UcUICERRBeU78MspUh4
WfBc5IczVkEeCiqPY4Xv1bUN0JCG7fnVVFirV0jSoW53vbQKtzre8t1ZvGmoswcU
7mXes1HCtAPBTe10sQi6TV16GSOnNFwUeqnEwoAwMw1P56HmGkqrvFIsdfhf84Wq
SQ+9RbcycGRPT0IvbTbscTtZcX2tOJw4v95A9na6Ua067lbslAI1UvlD8Knc9vf3
jZBv8RECE4o1fF0nSMTcrupmX75V2m2ji/2Y//b/6c+g/OIczRaGXSDzPo8VrjgV
3LkHftZ1kBRtzzazx2RJm+3IT1R8TX3OLwR6+DaXVFI2PSwsxzkgz99ktOID8yys
6UJYSmKzUv+A+6gHfPkKmXD6uBgEpCCYXr9rpF2W8As6AvScqAGDsemiLTigY0TK
eaWalpUf3QUnMQFa41w3bt9JJ9NdIALWb23DMCIhQxmgRydZUzN9ftCMApqIko6D
j4tDgzISr5w1GUc2QE81cSClrQUsUrqNFvZjxPmHWwHFQlOWk6HCNwsWyZdtRp2B
eSAyaV4U4Sps710ycO9WtKwpuJz+lG05mxZNfzaDWapHFCQ9eds18X5S5KFlJGsx
ntxAV/SC0CiJQyxICBR+afLeDia+VmVb/Xj+INWBK5VazY+W/xksYUz3qHUzK3wJ
An+fwIGez56zfk0sYS3PQbmnThc+a4Vfu6l73TvBwAtHOx5DuNrAnEOr+TA96ZWu
BS7HcfRUY5b3LEcm6/E7Ax6TaS/qWGrzvt0lb0yG/JuN31v7vwlQ3ggTYbXacTBw
Lm4yP0UoB1+XwdcUzMEeVLH/IghGJ7arMyzUDnt2m3E5wH/OtXWPFgeB4OR3M7yz
UieUDcCPKGtDI9jOvRhrpA5vPNF7eISkZb7R5uqYZtcObDTBBKYM8qNKomBqSC9A
iHZYhYtLrL4pZZbyEN89x6jJquQkGiO90+OfoG2gEm+QQkQW2iPfasLuHqisCe0z
xpRkiltWNudmP4Hg3+0MbxIEqBUzfZtAsdIGvGRuDS1HlO8+Qi5ky1WyoTxrCVhd
zV6u63sk7dSTkrGxtdAwXN1nmWmlFPr6CJ4Oag6SP9HQ9ls8CS/kZJhdgGnK1HJp
efv9IHeXWld1vGNjfw+TuRYpvjVV3OOm7f6kGC2qeqxv8vLb89bhXzv0NpQeNXDd
pm5rxPFoGUUllal7gfA1UTp5zwTehkkZZJsX2gh+iC1J2dufKBNXJo0coBFPfCMh
AgkRkbdUh1vYRmLus2iEBC7zo7qLCMn4oj79ddobp0VnutuKewtldkucYr6JthG/
cP5Fpv5TyGFa9xVgacW1lu0AEYZoWS490pIx5CLvnFwAtbdqrxnZ0i9WqD5SYjIR
qCQrLxPMnPRVQLlGkTbaJ4wYUYiKXRPkSuyTyBMlIZ7QK2S4tLZrTT7mAHNP4LWM
wF7QzZIxGKCfUihKUDGPevlYRNPQkNZutr1uqsTMNDsMeXsuh54obYJ7BSklw3W7
tdkC+AN+7no0LYsOrhevVKk31mxXztAt58WUAM06zzuE3VL8yhrt1hNG0R1E5T4h
erTkxjVJ1E59UlUx45FZBjzMpQV+Bu0tPcKd0b1LIP3xkPpbycYj395C7Knn2WAx
HRTf8QfTZOL66a9ClU3uQNHzgm2I7Rn8xaLb7R/7LW5B0m6e7Rn7zIsSkAKNqOgK
jE//UtXNtgwrVT92MG85Mu6EKXwbtBS+iisPPyjFAwP3O3m13F9okk65Qkodvdk1
QlLNpxk6kneaPZj80+JElHjtJ+CZ4q53jblMvx74cYkWSj3Q/k5p1jwq4NX9PZWb
6ek7rZfX7FR/iPp6PHiaozDEEf5PxXHeVzpJU9TbiHv+pvxMZRTQQuQ6lSJUjI9s
x+8VMWAuDe4kA0xhkj36OZT++4I7zU9iOOgHKAEOb1sG/TmsrNLCxaThFkpaj+Bl
+cU/eAfEsye2s8Jq+uQ2xsYUMl7M3qUr6HM3v4qbh4Vu10FkwHMbenpg3xFZPwR+
VPdKJPlpa1Wp23UcKtke0ZJJszSLt1ZRhH/+9MOi8srAEpHrNroQUFTMoxztYlxz
jkGvzQSHiLWz3WT+HsM+rmisusa7LKgGXQWW85M21AwzUbI0/a+OizY2BByWl/Zv
Gg66QFqQeXRV7kuEF+7cpPdEAlOIigX7nLVPC5v0TiRCUxBfjJiZZprwmlO0XxX8
mT/+zZfH4nPv98wAeQccQ2gGSm7C4d5lQsrszfLbcWSXwyfhMLcCMJb4dhoPVVtB
DTIUFI7JdkKS4ZG+7Uh4g16jd24IfPrOA0dw49VGopPzz2fGKaIzCTXW/isxk8k3
qHM3eZqjYTt0hXD8zo5SzUnOjDDLeKJK2ZSIwQDYZfxhM25SxojimadIVh2JgHX2
xRnCwwWvtdQ+kUg7sT+idLzH0xafVb/YNq+MwcvGf14c88kgcYXuNhcBbCeLU5LG
KZbDdZsnh5HAUCQh1KWBaM8dDGhGKamcTAuHAVWegL62aJnyWCsmBl4XuwCDuZwX
rTJ+LMaC8z+lEyAlNnXyk4XuOYErIf6SyLWoVVGxm6XnlSN45CaoQNgR4dOFu2ID
LqvRBcerIIahd9ORm8NBMH7vTJiE4b84uP7kc2JrNM3RkZvI5pJJySZhokCbFghO
dJ31D1pEdVmtFYlP8RiIsbBkRwmCdLzDUAXBu3zR3TVFr2pa/EWcrVnGZxbGypEc
GJ2x5q+f45l6U42dyx3uE5fC/SQiWcPdhagSgW4pYQn9BEfWf05FJWSAIYvTmRrK
UTkTjM6vSKgYhmAnOEzxqVrNz+L8PajfK8tmDTUCiRtn89aOFa3vKZT1zuxVKkuW
30Nl2T1a9zdHZkF537mK8pbTet3AfODzMH6Vnpea36J9/1eO/v98YqAoBP+ENoU+
9sju8N7dDecqs54uSI9C62DD2oyJEbg8qH+y870W8dnVq9NE402+V7roGWmBQlKB
4drE86N41I2c2jlb7jTiKsuAw+O7IXpLZH/oiPSVmbX6g9WnXgXuIwsREQZ5wUDE
QuoxCuZjYoKYf0fgOQFhaNsNsprjBkXfLu0LXY2n1de8qNVqC3pkseH75yrWzro0
2iQYuQ9l8tSfwBuu37cfVZHe2i8Bvoi8bMMF0aHDyW/at5gtahqahpDOiltUq8dV
AbADnaUd9bdIujNG6tHKA8EtbMiIVuahzHfZt8n18swpwGD8Tf7HmNwYlJfj3mMu
a+PqAnndsM3vLY1CQwqPfQ/JUn/DQMqgzCOMEEupvBNfQk9rhv68UJBI4quFJf25
Lntdkoyua+8upTwpZEb11Cf4Ee7mSU+gmZ101y8bl/SV6fvmMcvewP+2KOKgTl+L
Ado+7YiaR+214fM7QeX1x/IcZnOVclh7f4gn5RVZHHaLe4uQzmxnCVh+0Vxpvu26
lPG4QvqFpmnv8cjKIsoDCXyTJPQ6Kpgr/s4xg0pQQLNxnGJA5lridtIJyUix9lSL
Hg26knqaXOezJDfMQvMy0GXdmzv7UR3hx0SINPGLx5tX3KNybyGBmGG4bAyPegX2
uGyQUHMtdLLjOTBFZqHZV4Pe6SeIRz8htnguC8ypb82NbVoZnVqzpkNqn+qP4xvT
Jga+E34MnRmRWcvhEpyFD4ApLcWVvSFXkFwHehuIzt3e2IoKsvc4EcDWrHLgCuHq
2KJ6OiDLNgtM8XFGrPce4Wpvmx0kGJzfLUGgvOcWqF3O8u5oUUeDJNKXHf8+NuR4
JC/Lijv8vq8qSjbjqds2p5/yny6kVm+Vo2aXE3BVjtmS7SFvlHj6boWczAeHAsk0
9Bqk+59cRJM2m1Dw+l3VIQWH9ZKvtyE+T8TlMaXBhhK3l4S7//ekXJOTRit+YR71
IVGSa1ZnSi/sKTBZPXcGL2ZB4VjXTbpIbxVAlaBNWKIP+NbZzIYI/HYYl11G/blW
1QFSkheKAo3gqrwQITjvJmqikQivREhzwZFleW5My0Pfo7JjPXmeWmi+d/JyUy5p
H+kUbI2Id+I8JFNCJiAxwt2DDH1+3/9vrbsyfjzw3d35LNqd2GzO3K0a+DFanAv5
MvVwgUh56DulNTei6wQ2T7/8sQtayCPn7Lo2INoNQpkEfKrksJRNm4OTyC2HxuEt
TYgkkizHGj66gx18W9noYtZ2AKgIHpMDZeoudWINbvz/7M+TA/NDVn62heS+xoAu
zcvTsyU7aXNM3KwAT29kaVDfBCI1TUTA2/S6yjgaK5aZDeokR7UDcgf2zq2OwXaR
aw72CyguFyxjo7SpOufAr6Uxbkk1M07wwHMh31gy/TU8wykwQawqQ5dSw2vzUsHR
9bCV+EIhl/vVyiSvzrJ3PdwMVBdO97efIjfShAd28PXncCwTWpx9PkWXdfXxxOfj
9bpSgavkt1o8mZNwUrCA4kzsHxhAnsEbOIErnt1rQwFRZXiUS5fXG1ZRceZD+4xP
5Ab1rV0XHQdv2WoV6vm6l+z+UjOQ5t1C5S7QwpOTS+Pqn8Z64BCZ/Q9PEhdP1IZZ
xw1MBbo2op44uwVl7uEcJdmBCP7HBXm9fxVRqDPQ0OIo/PLxgyfjyARoogJRGs7y
v5YBlJygA5R+d4ys1KJynZoE9IDCgAI/rAk/cRO0bACb/Y2n+eVvAOsdwCunuKdi
Bz5OKG+XZRWUTBtg0LUK+67proAoJpopSPA09PXM8Lo+EVIlZ7vDZcyldGMH/R55
V0HxAzUxb4zscqPs7Ux91Rp3Nk7/i7jSc+DaZMRsH/JQyIPtklAg9M69hBhs+q8y
wg/yvCAklN+ic90tlzftsi5YMqhfTK3cr27TyPOZHFn8vqZN5VndhfAS1AArWkwv
TqDEAGQAub1ZJW7FTBNgi3dTFWKb1UH7/YXXLCtXXd5A7is6GJgqzYMBnrDXIgLj
aBrMlHNr3MR4IPh7QwLSm2CKsb/120Aj4dZ0HRQUM1gBTgOtAkaw42yTR4hyWD5y
MWNm1uuK1AaEsKHWLXQMWZPU0xTTw17FwU7NJAAuIv8Kk4+SDPXf2VoKVAbYu/0R
Abq8BbknM7bXeiKlF6zCKILdZkWFgxQh5250ZcxCUdoVWUzHUknQxIm7MRAkIayu
3yJv2888gAhuXjZK2Bdjj2B5ZLPg6F5FwRPA2/LAqlRYGoYpvh59FRvAYiLFIEbn
q6YbIj4L17gayZa+1iWkDpizKsao1A5BtQvQu21Qgjyclp3DBlr83P2uZ14+Zg88
Dtgy0VG3+cud/tMMcNTNwtk1CIIfXx61R+T8gJPSJSExuVpI8yzog6KB1teMQots
HrjTOeeC1IWprPo76VRGZwdLNtJnhPCURpcQ6Im0GccudkS/W3bW66XfJDqMnH7t
dh+Rxp/bTwCBM0gLo5tDlkV2TOR/aHjlNMZ8cDGp6yX5Dgyp9scS2SJ8Dtjsebl8
LZpIjFcnEkPH2iW5nyP3dsWY2nzQl8Qv6zvddZ4+QqTlj6CE7IJMpUd6zzENiXbe
tNRF6/Co3aQ+hdL/XKExZ9O/yB+JzxnrFVesFUDNQ7JKJhrV3er15HCVAg4kDaY2
kadBPJgepT5YeAUJnxnSaMvwKVzBRU+EBmtWc1Tobj5dGrKMtS+BF77OTZCc280+
oeOQEBODy9eHIc6iYyeeSXMYX9adgQ7v2kPunM/p+5w/JxNeETTFwBGZ8YLbO99L
wok4HwJwrEiiW4CYPkX+QTHhkUXOVORcMRYwni8LqumNz25DAP/+Ey4ZQMAALlht
8FiU641SSHBFfVtL64nhZp7k48jsq4/AvfPrEp3z79A2vUxJx08kBoWsXn7BdlN+
xLaxf9DP18rCqkCx/6GGGJJas7SFN71PMuZdk+7GNxpYGUdDoFYoh6BKCX08LTs8
FRZd8V+7FmJftiKPRS661Ik1pnvmVJ6IHSGXS6LYQCvENzgZgNP2KiGyG8YgdrVS
bLcEUHhNPf/n+MCdu5NTd2UI644jKjeZzlVRE2xP6kyvTFQlrXo7JCy8bRCtCi7h
TFTbghrwioscojYw+NbIHwSPhSs49wQ3Mg8crgjepzCOjLmq+gM94q22Fk/kkISp
IhynG7S7FWPkNeN+i8yDO8ujpPwTWzBujJGW6pshFhzUUDluiwYkU24x+QW1aJkv
mcykxFl8rr7ravB2Dewob4yrgqImDLpl+C5Sk1Y5VJtAwbx3CFTBM6DbO+aMtKR4
9rl1KfIrH0glbczZs4QdvAJ2FeUlwcC+NDz3+PTW7dYOOBImluu8Q+uUCkH6cfYu
X38GOusUU+dkYIdAnUIxJb5K9C5eGrXKGdXACBbzvBi0xmN+Tu0sFl8HxTQV7lbN
/S8EL5s6nOTJ5rTTXkEL4OOslIsZvpWuEw3Oa+Kt3RfjbLBq1YEunOe4L+SXTdNF
LGKW0qGbP5VWWphWIAMB56KiESfRSCddR3SNgmHZo5OoryTYAf0C6HPiobYf0twM
i2jG4IR0wy/Nvpy/iBISdfGsuPWyEdLFz7yadYHR3LrYB8zCXLjSsr03XyOF0Z3h
drE+57cBoAEDRKOL7FqaLxCvwA69yYyLLHk7iQMQNlWjy4aj0OharTnZ85Wk59OL
ovU4Mrj6r2HVkWXsJrIqUN7/ACdXCxDUtsNrIdWqdMsmQTqaJBjgVpwEtolTjUPM
WdFeFHc392Ja6CuVg6tfdHjt7rUhDfySZ2qRdvTvW0pZN/NiyJ74L+Qtwttt4R8v
Un5KhncrTGgPL+hzZ9Q5I4RbZ6OXmseCv/4IEiDnQg/WUKlNqgo9+J82Vyz4gBxW
/yKAJsNOx7I1vsMr7wt37/PZbVi8Klo+eIfhd8GQIZGXxPSUmqksyTvvRmjXxUnW
C/eHYeEv4+JkLmidPt3cwf1OndWPWRM+YUGi1jJp4ascnRrg0IVjwjcZwXq+Jb9k
olMk5LqilWGgjlME5sI339nYxpFtJmQ9LVqnoA1J0/Bzrn4QWsQEqPsrXpkDYGc5
u8DcRlM6ivaS0molYs+qw+CI9cUkxBewCJTP0bqaIRfxE+/+lH0Vz626UFbODf2K
5vvv2UpOmD2Jd3Ba2dj9uzjQ9nC7t84HkcHJxvy3zJlW18yxdmPAPoANjEY5XpWO
v5/E+0NW3JdKmwXC34X9aqQlpwHlvbkPRcO+c1mUgKNOfy+M9B276gqPPX3iZkvQ
YHOiH6DS6J8jatyH0cKQzk5rQ9mPS3MjGGDRbyxzlLEQtRLhcpc5SbZRe2P0oydI
38m8OQJTc62eGEd4ARWZhGX6xt7rSQVkix1hArkJJijzkF01N2RJeFe4rby2SF8l
wLF/kC3JraoPkVtJxPBGmdffVmNL0uWZip31zJQX/S6OYFI0nyFiV7McXuszoSgl
h//pdXLqe8w2fj6uzO6afy5q92DIB6oJQu/Zlc+fv8b+Kn8qRffwkMe2NLBWKt0G
L4plYpH80e39y/bxqa1iLMERQchkxaggUJ2HoZpxtCu/xY/VMkTntliJcVAPii+h
hYS721Rhz9AszBVAHjuwHVh54aoc8PRWkY3zR4Nv7f+XW9+Aj3dKs7LRtPkZswZi
E20fhR3Ia8G80V8UVJ62Z/r+Bt50azE3jpWdWzh0WwH6hT66rr2Rx7KpAaR//xU5
o2EbBhQhlp/n5EydQhYJDRBAyJx8KGxxyPoOv1Th7LPQU+0cbiTOtHiZWxwMuKJd
wP6c2kgwbh3HUdJol1div8oGBFCa7KB//jtp6psNmTSv8XAeC060gK+R72BmZs16
3uTvrygPt8G9PudpqXKsS4COgOZG5h3xEYEE8wVVBcqblbzGpaVrMi5UsoFU98vx
4223ZM4su4RyzMocH9mTcpLAaqDTEWe0RloJBqAsR+IHoeMYSt/PjwLy0IhJjDxO
t/g6kOyt3Pre4kftj72TTZ1HfcHS7bya9No5yx6j74bhEPpTEqFWbWBn7ky6/fWT
9X8ziNC4H8eo5CaKV5OvaMbFu4TD+/EzojV4EsbzPX3J6wCbpdv1DyGOjNXGTOMX
U8/s6nEK9uxXchfFX9wL/3C/WB2Hb2RT7YXwZ/rcOh28CZuFB8WHNRHh2hLdVAI7
9Py+mdTv1tteeTEOFUCgVtlh+BPnv+Cc+t/bAMeWSLbv0yESK22GoSMv01UkT2l7
kgtwhZtPTb7nbEqJMHhPYEmUfHNFk6EhyMxzJKf2ySvbgMo2HEQDebHE3umvOVEO
8bNX+GrBTq7eA3fWrc1w47e2mSQgXK9At8/UO5lgRQ1zvhLAHBYeD8B4lOJTNPDH
GawpF0FQQ86lFHpcOpJHiXhMA+9ooOawYOqOL1stWs3ITjiAw8GsoRtjtWwmyJar
wAg5tmDn0M/nTzR0DXUZa8GHtUy4RLPYDYqMgpsi2Q7JfDVpaSXur/l6vl6hmNyf
JGKUNpaYBLXRF8FGGe+/+YB4AN18sh7w3iGbQRlRDpJqeKqF6GRKlZ4F7CrHx1ls
tkRNP2SD642R1/i8C8AA+qPHLmifPIemEO48dZ7oWbGhZzuyXFFOPsmBKpMtcdva
erMNoprW5agYNPQksfhRjzBar/LIbnEaZyXUv2TyMxPB4BJF8t0x7KT/Jaza0W8R
ye7aonwgu/9U//eNKKA3AJhahyiU/vhTEh0N888QmkAIf3gyp4evKfw+jRjWQ5n+
9eeee8ALoaO2X4tJ/SzUg44s8TvWxkOBSvp5/Cifnr1No3lkcUk+WpjN1BCfjdhU
hle5Aeqi9f0HOJZXYGqKOG1T8yY9cJ22x74ul/ZXEAX8+QvPQoaKdtu5EwjBPt3j
LB843QzcWUrVDZCZ1m018QypzhqnG1Ug1c0rfryoWIQvffHTGgmzIp2HY9HAmjKq
3lS9QYmXDlZNFXTwlgIbbxUx32zVWDrfImmzFDGlHz62Ro8iCGglfkJjBFq4NpGm
xoMnDzeEQT46zQHPkjvvHbPBHm9LGVBxel5nT+nJxu4nQd7Lh3Niv3XYGcfWQ452
MZ+qqzefDUcuchHnwAMxVLqAyVDhC34o4OmncKShHsBoALL8EGDy5GatoB/QaNC7
eHKm1dTbw5dmoPVGpTtHeWVyoviMUBnghfBJYrs6Hmkoqsu1Cu+QfyM+/mw8bVy8
Z9wP+4dOHa/EBT1kenYprOuWdjld0543V66vN+iIhzI9H0zvP05BEVzX2mabzH2S
ejt+vM/N/bssjLaMUJ4YfI6ynjUw4eAoR1rmxKABAeaGgX5y5IUPaoQuvAn4ZGXs
Xk3WupYRFEXneWbEv2cksNeOcdktc99Lj5X8kb+iXrnZXEAg7GRrFWub1LEVwGbn
Vjo8RUpPnANp3kWg1a7G+vjXzpMjJmhpqNdD06qph5q+HCqwy9JuIm7Sxyx+v8ei
k9xvEQxSG4CepcdnyiRvLvD8c9L0xC4lSX2FgN6nDxaF5DT2oJDltcm4kBNYiCF6
wtRP0l/kzstNicYINEfMQ/XJHyCpZOgsWg4B3Mgdr1kC2fqNnXYPRmdxLrh3b3kV
uAzpagg2nLDcRX2jqPa+8heB31UtIWHoNV9keN6jOSugqrHrNTkzkTqDgJMC6sVZ
MYHFvyvmhI8Lp24IvTYZAQNBbDK+6eNvZX2PPScE+REE6to/z4dtejejcQ+cwYhD
bjcamQOrr4W9IhHhWQfG9gJBA77sXBICbVexJFEIiKoQVcKv1LhSkGLi4tkdQ4e/
etWuvE+i00lNeJvz0Ja4IG6JSlRuhfPXpue4ZMfyK2ZzPZnJPmyo/T9tl8tDD3Sv
lbGR2LC9WHV36L4pQPud6drSR1uuzTlwcFma4zrZuSHrbeZc1mKM7CRc8HiMEeHK
DSgcF5EVgQ0kKVA6jQBxG+YIrktdT7y9/p96Raz9pIzeQ63xX3VDbwXJFO4hfBfA
g/efPzKvCkPSW5Mk9h+G2jucIYA985XsWj24jKbfRg+lFz835M8WF+mEH1x0XXmL
bYzKk1ZD6+0KzG0bDqNXMommM8GkUcjL1z8TUUvyXLrh0dbfGgZL1nLmH9ayd4g4
bk4qImquomoeEJZEYn5vLSkcUP5oJp9+69fKfqHpsNgj7VHwuXfTKSGXZQ5MHYXY
Wwx0zzgHl0cT9KNHOXjBCXhW8gDYHOXSQUMtw6SMO2HFEgWWEIj4cnONNjtDlaQo
70JkDvyKqxREprrw8w89nGSe0waIQ9iQD574+VP3uH9W1fW1P9uSraG3pgdvQLUr
hOtN1TqFha/rJ3bEZ3eF1jGbUUlTg8vfCF17Fsx4gt7VXcy6Aui+GDLRcLwKDF6h
mphdQv2yjEIqD59nPC0aRJIJXCsS5jJaiFLmLmGtiVTOlcTJ/EIJjOh6VsudIpIR
kcNjRuPrRBvzCV1TSkfhlFP6DFZfRfi642gkx2DVaqpSFEUQjMJNyFN3LVHrOW6d
GJuuSLvmFsOXMDRKFBQiTlS7tQfnRIYo+IWNIkvcJAFkmOwDru8iayNCYRyUKsrX
J7HOE9w74qHbV1oF5k4xp9MOW1mpc4UePIDF0mktaxQSw+oky6jJoExyba9Kw6ez
xMAQHhNvXR+UiKcwTtRX/hVQPhIsAmCTqG2UOOTFKZm1gVPrbLmQoEVGUksmA7jZ
qqlOycqhV4PdZWMSX8aGV+vJbZKIKHqPvEzlZ4+FVrJPEfK32nQrQnzCT80q8tiH
beyvTJzQ6mz68tbjZ0zIyduOVSg3+vGVhx6qSIDTsi5I2/cGKumiQuB5pMKz5iII
x3TepVWwQ5mh5aHytSSehug5VEpzsXpp6EQAsFOu8W+B/N7ySbKW4ikuJH4dTK93
bvMAIhrWNL189rc/Ji1SxC6sltqMmkFL/GOe+MW30LJQL+0BQRPVZhzsDReR+GIn
yW7ljMj9GWEpN/SBkwvKUOFA5VgRzU15a1RpCXwR/JycDpAgK/kfiImzlWOtdmo2
HwTq4VAs6nz9J0eiEIXjx9RKGbN9fupQEwM6OrPHhO+QCq2NteDXpNim7/Kk5pBA
l1COU3kCc0/o1kBB+/bW8XkF8lVrqbATDQVrKOoBG6fSnGeqKUviS676HeyNRSVy
h5XWPWqPtC0nod8kltSVpjNa7nc5r7dcGLIpkITMKpl8E9fFozv0zv+j7H+cNtYu
Pz2Zy9X/6EWkHiadUuYOAgH7xfTJtNMqnUr9gNge1hZpyHHXGiPPAZcuX3PCrcCD
caaQbqUh58jPDWVjbGTgwby9NkN58t6tFX6sQCuYYfEGRKEJMUNhwBVEnA4NpzNM
zSngqJVMtXY6aMWSUg4S7kt6oJzlKRlFuD/OuhcnLZjpzRZ9iWBYyBdebcHZAXJX
ObA2WEwxrIWDq8BdtP7WMjA/2fHScQ7XMH0ZM1UVhcsHbswwt7PKXVCN2JpkTQFk
2G4FnFlsDvTzKQgGxzdpOeMS0XzjrHy1JQZErcvvw6lXOyw2Vlz6gzIc+BN9derd
BK/OCbtw7ZWKZITtWM/pLiuhSX2ZqUuB3jbIBD82Xkz1RTSE9RihuJuLSY5DtUuP
JoWLC6lPn7aIQXmO0MVDAUD7VIvtl3IfXDFGxy/YmsWjHIME3hbF1KDOC27mh96b
974gua/w8X1/kQ8Nr3GPRF7BmrLYV/CdvLNnR6KW0OY3Mtn8Wgx4IOkXBaWpUH6Z
jPVoUyKVniSlbn96bw1PgzPqMorjpR7IxW2I5vmRihhvaPD556OpuGCcUli+w6JO
gGJvIe+FY+7dzgcsEzAPJPDPU45ke6Z6bny2xGLJLd8Edq5W+diBHS9efpOfCdia
xwA4SIs/eAPsAW+aYVHnc7cqYkrbzVBjGH9i/A4WPWC9DlrKju8mDEqPIj+wkNHs
Ozx8Z5M0c60jiYmuSJmUSCLtUgM66dM0JdVrM80bxTWSxUpkfXJpaS4Scj+/CYwt
cMb3/w6e5yLe3RatfAYgx94WBWmZ6lhT1OBV28wXIuTZel2tA5lhIHFBoVHC0whv
FwOf7EPICW/cW9pztUjiQzDFZcWjneXTnmkhzUQCK+zQfdYWzDIOPBsUlInCuZqs
rbym2bQgYuAMFno60z2wXENaDuL/jOx7mlXY+P1Zo23mWE+ZUrTrP2yKioKwrdeA
R6JIkze4Efe4KoWtsrBR/4PCdOtCB4Js3NAjcJNP/KiVU/YgD20DW4IfI2zhIOnE
gLMrXSzJm708CSyrtjaCiBrQ/BBh23T8Duo2w/4aa7Tjqlqd9BlwdUh3sSYJ5WGv
g8qcTqVmWi5JWcWbzHFmMai/nT0Uam1knmHQRcPVOkEQ5vcRYgGWZSavXkaoBoDs
+WXZ7igj8B/QW8UTqIj6rVjyVyH/ZknECuEdAFbSLuB7d/HKUMXks8ifVO4tDHCG
5lV0JVutcoH3Nx4uIM95sQQjM0D+YLUVXlv0+6q+JvTtXPt//r4k+nuRjdAtL8lR
QncC7ZeHvl4DNGFp1sQX83JKkkLURTtPCvWzoUZYILcoCRVEJeDqGqkTEzIo9h0s
cqfZNoY6IMggMz5hYqKFgqAjpSEiluchxiz/dfGnM19Z/lT8l8faM8OK+z/aQM6I
w0EBxPycKaMDKa61H3KFgVMdQXXyF1IDFALJ+lXYatiWltAhCGhAR/0QTpHaJN/Y
0wkJ2zx1wiN7fWbUSvtJCojAvneiYazMyfWXeZtkW17nbZ1hcDtw4qrGqA06njpw
ZDf/x0dl9HNad+WruWRmqfoPSoCDQLkmfiqSD6Qu3frpyCARMbbEKVN9xNcC/QDK
4c1e/85rrRJlWNktx+52ct8++VjG2lkr3pNazLe+X6MJ7eXuJJdyrlVBIgaLqp7M
GPzGOli4UTYDI7Rr6kijvh1Al5Bq5WyBx++5Klp7TB4OJ8ZtsiJOQ/PziiB1WiOD
yf31OTdLgD7bKq05b9U8UbfdpwYTSzZ63BEDf2m6a1rooHqVNCdsEGnXdq52qh8o
lPJGkgLe0aewvyVcWTgwkjQxxTRD40rve0ljr8idzz8lNSiYF1VT3WlMxNZmuRwT
l3yqf0Pbw/6jj0gBpvVkeXbD+oD4aJ6eaBrjGW7z5JPny6S0BtWR1qVbJW6hMAAJ
AA0/HeS46ARgusT2PBo89qJrCLLRGt5I8T4TdJXK/K1T+kqI6fEheyH2O7SDeWnx
weGGpBdqFRunTsP85170omlRPLSAU9aYw0HOOh4/irZpX6h2eLg0Y9bisuF/HQ/U
xW597l9nPoyEwD4EPP/cL8sa1z0QmlKFJSDl7z3WrwZzymDJ1xo9Xj4YWPlw8Vd8
mhteqQs8UWD6tIeRH77boDzzGxKnrY1mNwZlgEJqodnoL7LkCNbMEiPwkBXW12WD
dyR+fgd0+S2bN7Ol5r9cMmo85gXibC2zmz9BVUbdUtKp0uBExXJbbxoZ/Fgeh9Zc
AoC6rK0ZQiQkVwfeDkvq+qTsHMCEYwdJgls0PhpGuoXhgtSYFfFg7hNrLtUroUYt
+LtRxC9T3Re2NB0GhzHc/cn2ZP97JWuql1W8SMMEEnzEPtOZfQcF52FoFcaUMW26
7UCIS34T8QcnQO+SawAE7Tynd6K8T734QQPnyyAR1zs/L+7mB7n/Ac/wXya9nOXs
DFbcfb1nDFlLGasYyse5UdZ3ig4TcIsmnxLscfm3M/c06LnjuEDEITqev9Kq4ATJ
qTprTAhN8YssIOnkNBO1/R932clp+kXDSsAOx3h69UIfe3UdfjLS+Xup1hzLg0he
DoL2MoFP0uEPQcsCjAuyhp/HvbXy5d/VphUexii47X1naq04wd49C373q3o/Q7kM
Bv+WzxDeusVNF+JVlXyi/QKzzU5XW/xDZN+fIpTt5QVn5n/UERAAgHK2JZEkDxGt
ThGyX2NzB+m8xel2HDpWYpNJ2U8x3rVOZJh/Zkj8r/hQr/51a9sTAL1/CN0RP3zu
X9JKQNa35N9Y8faXQupbgdEl50ZWOHfGqROmpH+0KR1kR1lSgxIgvcjTYZv6Cbvd
BMiiU3wKHthOvEHaeN/VzoTd/gzkKxHNsVc/Qqv4nuVannfwhAN5H0yvU9ZBHAXV
hCPBEYTzSGNwAFONbqwPj/d4g3DGQDbv5BnFF/tkWvskEt0UFLJ5Jc9T0T1Sa0Hu
66Tzkk6wgdxFJyvv85aytNzaP+BivY6fvph5v47MHFjZr3heq3/7VS4+wvn7MCd4
rjL1B4IBTml++pDQ0W4FagZd33I6MkBGLKPAC4iUCQn7W/58IZEPMhhfECKakMbK
KX0/C5+pWrJlREmFLgNZAdaf79unfP8Ofwvkx3Xb890P6Nq3LF0dksv608FCJ6F+
UcqGqC5VD4387HsXwjhGLYOMaeMBm+ddXeXqOdl34UHJo1BqB0aEjBSQXu+eFFz+
6X6VlAfdX8SMuvgUJ2/8a43mgbQRy/c4NflNk5CxH/kksUYd7gNMix+r5pPsbpu3
/gdTdE9XRtrqn3xqUxmwFMbBioQyoJEushYrIMVRsuD+GpIN2bO0BoQKRtCzxkdj
7uwRxo/nCdRmK9i7m8hWVtYYyKnjDOyUmoD4PxQCjRuwM3cWAiva6GNw2GXt5bkV
ZoKQ9jG+zBlke283sm1XB4s9VIdcr6Mzavogve7wTxJ1WtQeoP+mCzcZQLdSZ5Dp
F+7Q5ctYDkh/fBhsCHc09HNAYzdmdwX6uIHs9+9pcZqZ6GrMZtCNB33pWWg/sv6B
GDjjri1/AOOYJKxRMK+p2hnuG+FpCXj1m/XcrsDZuT18RGSVF+VBhyj7NzVvLIRq
bXuCU4DT96eYoPifY+9pcY0WT1qv25Og44IXXMyl52Fx9SiXOWd7fUAiKRASwkuB
vcaXHltzbFBMoOLCS7AUdjmye9qySZndBoQ3E8EQhEqTMTAShctTuIeHdCpsxMVU
gvlVbFOkXRyco4kHwg8pQU6lNNUjiQ54LzyrRzaCmZ93NAxNt1oWog7phoRDHSkS
OrxkilFpRe8qFjMOu7Fk2SGBqJKYfdPXjTHxj5RJReQJ/wisJL0OY/q+GFaGFiXd
cDUiN3bCC0I/WoMrq5wtnB07uZNRNd6vb5GYv4kwHREYVdsCeAM8Qa3oRrTWWHXz
qjCZtwyc3EoAqMa3wFa/89gluR1cktuvr5AIngx0OyAWBXqBtTt2+dz6PLfM24YK
+sIGBkt8wedHzO74hVeMmERMuZgrU0mEFnHqmP5DNnEB2LlSt2eefevaQFzA3Jp0
YEO8WgM44HkHwgemIFiW/YIssSUT093Rx8XBvYfkKCPGk2GXq7Pd8nKYMK6yz3Gf
Ib8Ti6Z6Zx+ug5h8FwgjDDUDULi/V5QL1OJfmUePeo/8tyBzoWLhavRDJhIVMxUh
hdMq3EeXkbzJvU3dnVxCVgiP/Hmj6Bxq7+TtNar4Ixli3BWSM4kDELAq6SpY31AW
r62XA/x+qrtrmhj8proJMYj5wI8obV2f1GxTryzE2rH1/NrF+LWBJ4WEDMZlKzRp
/uvyzjWwX4A2pPJBI4FIhfVzRbT9s036+ScAl7QR62ZhWKgOZyZ9BWsPz63igg0H
YmmLFj0vaTx1SoUP4XnGoTA9oDwAbBHbC9bKmfQpHF8m/E1/JtyiKFf3PMm7tgiM
ptDQrkKThg+O5bZKT5YV1OWqffVDernWynF5mUazREt1AHQeQ3r3psWAMrEX7Sa6
Iuy7xtTGkHbOYBrBVeFl/gPqnisrbbn6JOtEubgbveWbuENzMoDezuksbf5zonl9
pdS/IIJjTLgRmtPAp9jJySxdzRzcxEehWYFPwzi1HcWSplqzOpHCnkpP4QJpnM8V
bkk53SDW30QuebIqRYRjhxv6UGn54mdfodH+NPLzxgk4afPkbodL3DePMrcFTeKG
3YNQs9BFkBGLjeaQIln3/LdEu+lktNy+CfTscF8mFy/RWSLhJWx0z4swGYGBqsdl
x5otEWiET1PPfqRvqXjhxiPTNp5gm8o31of2PaETG46+6mAPclK6vpCJOTlUhXWJ
IuHZGmmT8JWTCRvUXZaS8unDPcmAErXNWetWaykqczEJsR0g6+6w5hwaf8iIBqiP
53m00JQ/hvh7YlBh0PISczkffDaqRV64vwH/GPeJdiPQdHx38ywUVhguaUwS13Ub
KUYImUw2rnI+74HPRk3M4Q2/yURp75eMlpjMTrBuUTFpHllks2NzMcKOblgwANlJ
qdvpXb8apmVb7ktIGHkhAkkf6RZRAsohJDyif4rHPrX78Et8B/nQsAvs4VVpp5As
Wl3uRvGw2FY6MBclyARyD0pAJDj7HF6pro1EG5gq8+2Sq9NUJGj9M+vVxPNR4r6B
npB86KzrRLjtNU6+XDb2BgwNgjX57ReFL62/O+LlB4g3pMa6Lpa0Y47RYh2C3EYT
DZ11AAyJtSgkZsP5sao5ljGQ/wUY4sM+3nlNviJedmLCcmQuGZzp9mEkvSQ8QEVa
Q6fztIHfTsVTiUFx8Iuhap1Cfj8LpQW0ARcE2PMcL0VXxYcDLkKsVICuraQJE9q1
ALF9JIoaC7QG1NQZGEmcxDc4YRD6x9faOqFV7oZNqMPbMb1fv6/3hpdvFnsuzxuD
eddwqhimnQHjUpCVAM3a5q8hGXqlElIegaOsE1dzOq+OP8VSNlu16dkJEsBzQ7OE
KypxCPZYvDahvXN2m8qx1CXtG/shUCQyQgE5yUGkW9fe043CxE+zdDe5Kbg4y7j5
NAKoV5IaXKtQbljMn4orRC2WV18txRUghMyPuBlxJQzaVrrrt8mSKFbaiXPiYyzv
z0bmLoubrJxZOzBjY+18gc46epiWVNJQiBv1AZQPQRjqrQI1q5zl2IwdRtATTdCF
8M4R9czoUAzJLk5Adr1QL/aBVPW5jsEepAEzebRwjwgOBGlAZGFo+1I0dBe0EowD
4wz+tU8IeY9bvTvNm0bIYOlWKU0S131DIVwp2UJ3ptqX+0u3zWOeqtFRzk9gV4nY
p+I2xK19KPlYinN7/bUZNHZbHDj+7lC2nU1hFBmSOf8/rH4J7jWTuNkF/JbTdIBH
GkkvDk8sS7M29O8wi9xHZlMhF/zQHd9BrGr+9ENWPx9WL+1vkqeQHZtd0OcApQWl
UvnYymgtZ5XLz/4han0qWAZ/33wJ0NOPpYwpuH3IBwmD2/ph1mLhxRQR/pFdDidC
NH885kprNBfxM1U0UeJz34xYKfujka2iAx4U2lSmQaCpS9cOyBPdU4JvCe+q7uNs
+C7Wgf6sX3xMhz7iBe2ddWC1sM6CMk2TCBMAWBbOeEBFi+X/B7oETblCu/HtIute
Rlu9xt86mrG2V9M2MBLubAmoPpQ0JQm2d1v/Z8tJDOqUDVuZ1CgyYCvB+FIR8Qe4
+uwCjJrJMVV6RE/KTC6OonzE9hLUKjALNXlAH2f9KA6yVGpQP4HQ6OSLv/KfX9aZ
22eHvajPo4CqtKJw8OpR2r8njvmlZ5vZf/g079SvHuyFUVAXHLFsKCHf9xxaYOE2
Tl+KfpsDU+JeF5uPGhtwfAGmKs8Q2D62+Vd1FSrHq0Md1amSdTdZNfF7XY/tmmPG
StqClJnufxbYsHP5YrE27qBA0BUSmG4csZ4gS12q9u4iXPufoF0opjjxkoDo5wKE
d3t0SLHFp/EKZ9Qk0r5EsO7zEgWspaU/3F/4DDT8rk0fvpwt9pQLT5SL43yQZjdE
Pnpk0sQaPuYn/JD+cH6FMaYEfrYHvJqO/EFRJv6Ban9Kkr1v7kTgyK6EC4abcvqj
gnJSoiuoEKIBHAjug38tBo2MadNhNn20JDm12AWXN46MN7Pz86Rqf3g9ewebwu0L
X56wtcG/vaCjERV6S9nxyy2ftJNLBijCejICDLe4+8GDpZwz9/8IMcBzm8bWn5k9
26Lgh0OyypCRoEgKWx7inl9iCyu8PGls2aGy2ijBYWuIQOM0CLsG0Ppf1eFDq6OA
KK3DiG3xmR8Hf0XKsQTUjI7tQi0jrtP6gyBdsWhDL7iFApJjam8B+42IbUqVDfV+
BovJh5sPnhPA1rg6wJW1LOH7Mz3U9vqmJZeEdO9U3l1FzXmStAe5zJZNF3kaCdDt
SQ/KBDqoj0/cOfCzoVxQzCeJKkYIY9KJA9AKKkyaoEal81pkj/p0LRSFQD6IOF+N
KAlj+uwE4KjwFGN+nUil0sMV8DTkKZ/fNLekCrUeU/EBP3bXjmBonw8KkaTu2PUz
ff1dmodcaysO8nL0xXcC/N2DVzCdu4mSQNCzCDU3/q1a/t3yRgRRezwILYzLvc0t
mrfH/Qx4vDLHh06LZ1aBBDBHKUWEaE+zDcLZ57W3ckB0S2anzahqVGj2688r+hNg
A3o++/bdAg1zJ0twiDf2fIXvv4MFAx9HdOuuKzdINjwi9uCdmJv3mgZFmDl/E/lZ
a85D04NWx466QdbHblUT51//EZbbBH6y5QdzSEOcgYYQ8Dgpc3L3df/bk1fEfEwI
EqSGbv5rsrZpi91RBb2inzKjrduwTNLRK3ezpveYBkUY6085JsuVNcI2J2PaL9Kl
C9ux5DIROIz5QU5ypH6F+TscHutDr0HdxEXxFAfdYe5aK6kkp1WuuWc7bOS1+jTE
0aeg+0wvbXnZtH0EBKkoc7GX0/CRb2oxXODW5URGFTarcOim/x8Ul5pwl68KPvex
PQR9jydoDrWBTkEpARec9jRHA261mDjQQ5aVoZSomXGZqDjNwnSY4m/BGg3gSQhR
NlSuZR/qret0f7m7ekUH/qTEkOFtufA89TXnXy3ccgwnMaX/So65CXshHCDHtRJx
mPzZRaRwg3exnYkdEy1DH4w3fD9WVKxWQKcQZbjjZR7Chvet0ocAq1fyOL/q+OrV
iWpu3LKmdlMpVSpfPIOM145OhmljAhzOp4n5/Bd5VdUMHYMgqF8Wea2novzy0dXL
gC5tYvYEy/vFFrFV7d11C35Tdt4jVRqzs83x7o1KylRiyqjGirRG8GHVzDK1wxKU
Twr+m9nY5H3EMS2kP8RDV06yfC5Lq02hZ0LmYAkbzzHca+3mdtYvBd1+Auw1gbPm
GQnDzF7iDLb35tUjuxgGuUCkbx0agsGQRkd9Xk8e1lkzEKy/ffKC4Tye7FXUb5ft
hICh8ULu9AoYUfj1VqzF6rlheRj2PMVRF5sWLQbP2GdyJQ74pZFs3c+vur5/xn9a
e0I7wdfdiuuHrt8LowWUr3jYF6Y5eLGeqOWwR+CwyTcM8WN3YxxNr9db8ZZhjjBn
dSq559K1KjeFvYPrZ/3g/dA3YDIs3toICe8/qW/3ijS74lFGKlCgGTe1dhafdvFB
2LxA/5nW2iWH7fv5/AFQ0RvwPszdLlxl7BVzB42WGH3YboV+z9rzGcY9AzS6CUNq
iw+V8yOYtUo4Sb0JSuX4CnBCJ6MDOzNiUH7IWp0diAJyYZLCZ+L+N/yZ8X0ArDw6
Kq4JSKgvaO2y0qhSp7fOgI/N+2qPdlTd+iT4E1C2vEFl5xfxxMGLN7jkD07tHdRV
y0zTvVcZBdLIyYLWdTCqDZXogJcQJ/atQELrdBGxXy5ZpUtF6gjoHiwPI9Z/NYr3
qjKToQsTC7KuRbeKt4svG634HVPbMXSGG+nxSWihS47bH7L/9yyzV6dBY33b8wP8
P9Fx/0hrG9rhuxv4v3mp0GcGNtrhfiIIA6R29JuxIQhBfuH8F8upWKsbiUxVcD5Q
+kXYuLKIlRBQM6smNCqPpebrg+bem8S3Fvop9X+YukJrPL6WovixEbgiO/INCFoP
i82hJyNodaxx4rI53nXiU+clKTP7p6EkLNosKHbkxUc2DeN4z3dGxoq7/Cna0GjK
5KT8T+lJfPnRUZEbpSVBZQNGIYL8oL/kKY0syU4Lm7BCEt6LV05URi2NTRBFfPEd
oxJqcc35yBj/sJy6S9e5T7T2ut2RrWp/Y7akDasvhaWaZukylg9ayrShNKms9QoT
iMhkzx2HO41PXOH6lQU0dV4BmX2XMXg8H4qGw+Ld3sbm+/dvl1VdJNxFXQ+7dstv
qK5WgpGL5uuyvVxNjigc0jLO42gy7v/1WdujeWz3UqLw+O/v5ZLq+ZP4lovYJbA3
w9ubnyS2JcTR7qFaR8K0idNbO5WzX++KXA3gdASp6dYjiRpwo9g0lak0BhaRtzJO
Pmz+3Qmbs+/h+sYOD3GvPrwGCzaQusyEQPMWVipSoC1iPtAJQF28z1jOn3sku3W1
c7zGPOdhv3zz3XFgvJw3tXE8roUStMzZuRRmRNg4eAuHXL2L8Uf8nM26p0zEnQz0
o0wKkQ+zl4Uu5ehwLy7Sudb6ZXLUxyOwe89Ef3h8IFp4yTZNtavdHJKKNgwMvpBT
hlB7JMjeNdlWXjw419UTCaBYY/nUjf1uadTn9Wkqj26v+Zh5Vy1A4dKfE4JMe4ty
xD17a70XVAiDCTNl1dHYz2nttNz1suMebABqdaIdLlyrx/0ut1DutycFxKzOemz2
jM5CN/DcrfGyKGWHcNlprvkVMR19ii7B+Ucjpg6HnVvC1vDZhp9C2D0eXh4gIY0+
pqG0QJovuk4KoH5COOiZ4Xw5H509+1AuHqzDeP0PhXCYoOELzO+GT1HjFHoGlmBF
ecPteEmeMxhy+/PWtxK9mast2hSGFFC04vKuMqE2tsCvItSsLEgTQQJ+OSEP/n/y
iDyQyluBjgHy9/n75tzglfH9V9DE+X7MkZQwBvmxWngBsIFo096E/UC+bZoKeBbX
kIWw2mIqow4ctyuc+FtAauFnuq98TN9FCoDFDSHXtY4IAf+cLJWnyfvS9lVhvLDC
IFSzwUOXTi6PFHmnwxAMM4jNb8MhScLM36ffNYOMsVdCVzPDuxJU7ynph3QJbg6P
zvvRFV9ntOjsXeOTSj/cM2yYPGh+Eck1gMQrW/pCFbe0Gvgke7PDBS+yUD3RAGPs
/dCu7yQQYPrPvYb6pURlhc87/s/8uzXBh7ShxtxSFsGZ7tDiIdgOCeiKM2U37qxd
CleY6OhY8AzE3ZoCqsMHQuiIL8hO6BtyzVaUoBPkH26jGrn+WEouvkXVoOiNkCcl
q1xB8bg5mSYhRfR4JcbGjV/6XIxogtCIjsLzKF/3AAvV8hMHflOh1M12WyDgjTkF
Gv8b0agStrD2d8adcisaeSbutjoBbqWBRBs4G41GyAj5fBiKxi24M8NIpErqC3U4
749TGpAstHksakjoeGvOxplupfziakxt+mDeFrHaqOgfocCHf3ul5oz0LLRLZYEQ
0J2CBYDVBHpCf30pb3ztZeuO5I63FtjmP/YNws9MxIuvnAJeRRKoT/DJcWCh9SNn
MkjHfzfwDpuyrLXb1S7qv8f7m+kz9kvqj9JHy+m0OpLskwbJq34eGWTl4cemph1O
IwJzhLDtA0vU/HWuagJCnAtu61eS+pEUaNKKEN3LV6qFCyTtfKVZsDtHc/lROdwy
UtLBawVI43PcD4NgG/G8LcXySZY1GB1K9wtkYPAcABSATdwKq3mu+MUk+9SmRL5o
tdwM+poH2ruKlB4Uro4Jv7neikUiX6ighBkoMIxJJ34bO/Cf9H+7tF5Diki992y3
WFTXONfiMWFgavh9jAEaIzt6HxJ3Fq3SI5UviiaChoQ132LV4wt1wCMbqjkTZx9D
Wd7YrH/shnr1FEy42BrEHmRlFcbDyNqq7rl7FMOZocpQ4oJydywbLe+KNtboF2Cy
zNOJBzhTs6gscR7GKfgJxVZrtQXcggNkPNWRj1geOmDcbT8cKuCDiLhU6XXj6fN1
wXallzNJSD0GtYE5VXq58zdn8pK2v5J3w66NY7m9N8e+x3imCULY2HsRSPUOH576
w+Hszt0k46wpMttHoTo1zWcKSlJ8iRG3Wp21IfhRypNup3VrlDtLBKaDMEsbG/ru
6xO6l7bHgm5SPMW8CZWAHFE5QMDoNZs0vx7/kbjXmwQ0Dm7boSHl8GKBEKP+PciB
2XSRScCT7IjuJyL3HsB/hxc5zL6tt9nKT5qIAP0pkFbdrqGEIpQiRSc2d4l8Lvco
40ZMWY+dsW4kIHSh5+SvqNAxBLeWSAWpP5a4iuV4/xR35Kjlfs0E9m3PFFTKU5IP
G52XR1qLNuIQtVj2p9VPAnOE8w56isXe4wsgwDINorW+BXIyHQ1MwuRO4Gt1Lj1j
p0/5OxPpaxSxQ7F90lFseNeH8/e8Urj4d3HMcHblk5NWP315f6B3yd3mwGDjEcpW
UqNM/DLbcwrdwAkYaFRWgOEvn5yGOcBmy/KCPw51fhLKUJqVK9oNI+rGofWa6eVb
+eINNUfJah73yccmd94z38eY7dyR1pZvF6DiO+ztMib8gpdyThvM1/fSgJ0BbPkh
Li/KnJRw8eD8rbw+le1k0MSNS3CksdfaceDmDUwyWmXn5TSCICvfpQE9TW/+WJZu
Vf+H+U6fBYv/H2hUperv1tLSyO0iDjBNBpXBp4weURMCplosS24RYHs7btVu9rdv
ZYl1HxY3PGFv0aRHHjXXEkepfnyxVGmpkYANBkmgBEW9kb9cPP/SH9W04lNh9cZE
lUOOotMkPhGe8rdtq+ei9RNgTHQthWCUJGQ4/sQ9+C3Tsq71fNBEyr3QN+PoG4MQ
yOTdXxMkIokK3GzRmgUW/Mt9gmTSE9kdfPKAxaQULukJJLsUEwrnwa7lW4k8jyhw
iPlqeremUAi7a5AQlTL0DjQM5k7Yt/Y2OfAS90MwGmlXP3XvD2/AwvCPETU2JtME
7OyXEaSoD2+upiVCoUxNysSSmtcVWWYbFdt+vGfZepbvgGnI9jCACTrz4c5pdpg5
j23Sg+x155iQI9i7KNq1slj97/SAuYkza4ZtHyO4vk7ZdJtvcB1sKtc12HJP5fO0
bu6KZycgmT2ii+3qF1BBZtewzLFKROl/vS2OCDX6NHP3SptuB9hHMcNN/ioPlyQI
DT3RWmspRMw2JGd+C7UU5c1XPNweEm2MFObA5K7v0E78fquS10zA4Vm0ugUEut3c
Oq4RZFAC27YudQ6u9xaDJ6wgahSADiU3uPcIdXt3A+NtNrg76itoxd+0gjaxPIMP
BSMw01ejIIsXarEWyD7kRliNrCtjPlkYOcPoigDV+VSLOBmaUQi7EhxQ8P+1KWUQ
NGSx5d9cstxa9uELKSfvDVNBneEMReR4p5xG/MZEy95jhkmtzxWsm/jjzAwCLVMq
ITTucrUF/ltE5KeeUDTPZmbN/PVcDX0rTyXieX4rNaKFwhceOAzwdHP3G4Wa38CL
PnLCEz6THbRMwCmrEE7oofUE10+w7OiAbDm0Gs5eAhLdnw64oli515laf++ttPdf
Q1+sdDXlSCnqJrQudUHXuCoux888QZgTh2+KXR+yx+qdqyk/REANCsxZOhvRYk/D
4jTdsV+1hdbruBYz6r725Chlv5B7/dCNxD/lTm/EtN47Zd6OHM/Sk1y9n6oEkdc6
5DV+YXEGgYIHEkL1k5cK8IKiS1zQxrIj3v2HarJKQzPtexcgfXMpjID4830jC0OB
Ky6yFzTV3wWhLVbUmJkHkRXr1A+uCEVlT1C944m6syYROhxEdY/b3j0OmauxbVBr
0re8WJMxUbE3rUU5JLCPOhTSIBhzzegQ6+hybU+qNIf3nDoXaoWXANDaQXQvS2SB
qPGGX19wVlR83FLZ66JN1xAD4rv7scy1VuTkE3vrC07HUDSK3tUwNGJI0Wh5Rit9
yE6Ov6eYF6880N1UW0x9NQLQk1fAbT5EX+1eEbaqCAC/Dbh15wsQ8t9b6D8na8HY
hrj0YrgpXTm43A3PnGlYYPIZj3YONLQrV5F7Jiwc6oT8to1VdZURoSN8BPhet+r0
Nmw/J+jCRF2SpI6XagDi4SeZJw5wKzq6/CVUHCYvRivWaogSX5+yAPZUQGrs9u/7
KkT79QJ5GNbJEPrb8PQVZBP94YC7bfVrsYjI3BLJagoZa4rr/S/PasEybExQLSd7
3vxA5gO/BMAcLG+nkIrHyZKctu774jx6lVAAyevzahP6SJpyyMwIZ6c87ddQxn2z
NI6PzOtilaqCnt8n69dD4unxpbkjyRmeCphhRVYwWSnmf4HLjbvLaVA2RZCYQrRN
j9dI0nqDcRlPWihV+UXMnoQ8mmJrSzhtBJsYZtXeLy1kRd6ZtUlP65L/VAGQg8ci
CVxjNZ4NJMx4ncuGduOLjdGTGvNk84CBT85wyssK+HWjYvjlhszV20sXuSCpzu69
HwKv/aOhQABbjuMYT6zBm4woZMETRC+pUHdyyr7WCFAXXnAVL/cTxHvAr7PGQ/iE
RJS12LE0o7NYeGV5b/qeyj6Lbzk+S6FQdLmcCgN9o+glVVtnLCVQzfqwPKH9EL+s
P9i9tRFARslcSJPLkMqGxUsoenH4wvPrbm3SKEwYeX2u+fWV2HIBHhFA07DeZ34A
6Qq9WjYPoGTaQQ/jThZ7TxVAfzavLf8v9Es1hQYhOtcxL6YPsq4ttIjsk/aqmHjB
rOjOchr4sjqto4UbQFI5Tjqg8dg+N8K0kVQLYC1k0j3XFgeFqNXEJiHlPstcb987
dPNknWqK6UA2LnnT1D4GzWqg66udxkZwD+gWM55R3z8VUTSdwhNypWY052fMtf7P
CreoipJhllAnu0hrYlpQp1nxIgkJofjiXshnX+5fljJd4Zq4T6vK77lXM3tmG1ES
O+o+feto+yGwfI+qURQj8MlcK/QHW+PJ+3ZwkOLnArqKQrmGE4d4hgjXcEtI4cxb
JMhviv3jrH/zbPDFRezJNjaIsFjEayT9HUqEUe7wGJ1MNRffufEGSMUGtwOuti4g
avNNkK23efNidJCS5J/m8ObzOszfMVlvWQ3TimzNSnNiGNk4TVbdMbPiBq+h0Zmy
4//waJuziHME9nQN49tMk3LvF8S/KTUVwbIyTcqrVYWpZwUwCSl77HFmk4a6R8Cp
mOlCp05Dz8JTvN+hllHtU2F8aj59q8HVwMTjuXK0m6bUbl83J/nb5nXh+qrZhyJg
DJVvMjO3Qdj1uUEOBM6J9hQ3f50lYI9HR7iXBrmZ/3FkNgho28o2X7almBhOm9G8
SWCxZmRqxksJI0bXiFK6M8ji4SOl+WB9aPDo5jA9kXwI5VUyySHTKVNQrltR/vAy
zVEqoFDaC4RLz7KBjB1svq8+TKswF/aO3H+ixPfwI5vTkbCjDUXuDn/8m8+9T+10
LBsmznyYWkzzKteMHAVMtyxbs3s2jmAxMVIxGvk6u6HcIzHhVPQXhgrnSxV1YYjn
mrJVnT+kivR59Z468Vq/RMgfGKYlOYUOS3L8+rc6wwTGuut7sJUBd6Oowchm/ITF
TKFACm+Yh4ZpS9qpLI5XZMJdTd4Ijj8S2Jtd5FazCeepL38/RqEv4YR8ekyW9CEu
Y1GONPXB+RS3Bavzeu71j4r1CTnnN9Fwhr+NlmUqquTdmCEB0D5gjRBgPamntVgW
kFrI2t/hTzalqKvgbLIz0hMNXzks861Vx16nQU+tny0TQU3Ks2q/ov6ctcHkqXH/
WLLHFROJSvTE9zw9ei9eQTZs9q0ujNg5FDxL9L0y9jDiTMTBVpB7gmel1w3RoQQC
BJpe1Be6gFQuGQtxOikB3mlvfBsOZoVdS3puP4BYDwVeXoUNhBg/41qPb1HJpVER
uoAsxpPcUv6RLgiftEmKD68ooPowoy1ETvr/rZ30LOzgp/19NS0w2xolRRmnsMYa
FlbSJc+A6tDVXBGfSKnELgf6lD6f5/yifvf0Q65q9FoR5kuFAkoMTYptIa4g4nRN
4cnfrLhfASf9PSKGbElHiFwdN6ueRfslUsnvmP1ZzgEHrnIDIrqKwZn16eK2JloG
3tNdCwsoDAkkoC6o2EVPWoe9z25Ll0c5ihAn74azVVJSCxAivrVLvR/GHVinQVCn
A3kxPZ0GKMKljPPSky28RZ2xQMaKIIoQwmFxSVyCz0rlea1abzUOFaIJHixf5kBn
F3RkbShYczqJ2SGfupi3kf9/HbjVLXe5IoJ7x9tcPnHx6s5w22bzhZQ4HCtKIZHO
fBrlA/zpA/GDLVAnyZl45lmE4KKdgLawoOhByBWsPqFZ93oocKXBiYyZrDsD7AV5
nsfh1VuXGspnfLPJbXrqhIOEBoT5HPVmzMQWPfHb4X5hjNrj0H2/EWFbmi9AayaM
Yw/Q155Z256i2tH3IuRqt+Cb5uzedXxu37Q9nyE2GH9Sh1DTtVTwLRvEBR8z9bCG
kmb3zCxgi5oXpNqv6vSSkowaJIncBIYGbfKVPLKd2/NehSdRo7TD6HGw4/+bUUZ1
1lWNaYjFrmDmbSIKW5RKQcrB+jTRim6MCumAVlYNqDOuo/3HdT3AVfxwxJwJVtIq
RVJpRp60/fPjS93zIX17D45PTb2yhcpcyvZZCsSnwUBBBbcxN1lSGIEo83VofKSY
tmpaa5hTLa43OcZX5nnrkJpN7jYU8M+unLiQLSH0gSUH3sviqtjkdb2at7ip38gd
D2MLJCeZk6BCcj/XIfSsyISqpEo3Xa47LX5O4rK0GvgHDDnYS8OORjeOlcEVC+Js
4JDPG8/UlhhFiA8Az5oaJM9Q51UFhALtILPMbU+5BsyecvqNuvTMXJLuhOT3fzoY
fEeT6PTzI2GwbTq6VDtv3knxC+DZK9oi0cNBF02DUs1eVP0uFqHI+RQ7laQEb71t
K2yhnaD5PCqetZzEabFrkKBlMyWkmVlg0cWInLQovdiA16SVftqzHJeiT/Jf9poH
rMMsgN4ggiUZOyehHO9jaccQ+KC6Zk/yq8uLpIiBN3PnsvFlKDpN9nAabEfb+Ryr
nlLGmwRcr9oGZ1YqcZPtrhYDPV/R9O71WCFMJJOYryo1Pa6YLGzSZzSSVe+ZQPTf
SB4Ke7KSQGG+wiN2AokdTyn+iFN7S5yfjBBFkTTbVJ3WMprpRWqtN8+PnsBD55E0
RtLRWACdQUSsphkxFtiPFLew/7PlzzihHAKCn2gM6uUc4YvA7EEdOc9exsSD81qy
VTJc7qUrWXRppra6V4sd+Zu36kjcFmzb8ZR2MBrS+1QvjyTuuLRP7EP8HD7lZD2J
Aau5+hoj/3Im5+YShnbL4XloVRC/z97Ls2B/GUaRjR9SRhFqs3jo1yaQ+PhOAIan
X1yfng21FYJr04Q04oIoIHsUwOeo1QLh7gThtHUax3CornwZfLpQ40I6wvg7N88w
ywfta0BYyn/NSS4Kbf98n3BS93QoiBINdCFgDsppxJ8/WwIjgIZSlQv9ZUkc6uPs
Lynn4Hxkx/eBQhOsOftS/YDCX+gx4tXgzHgHXJbIJj8Jk0s41oZjDP+JQy2kisFG
dob4l81p8BAtTZiYTeytav0jC8puI51xeoKdTZNI7R1Kj/CHUP2z2a6wi4mCUWE9
gq8sthDwNtcIyhp5dEe3g5yRQXF04RT3ATIwNcC9LKhV2x3HZA9cvI+iDIonFsOG
oGBIEMju6M6Qg4zOUofpfbp3buWKUeLP7tbz3AH3ub84dNrsCT6zvdyrc0QiWlXe
eTY5ArZV0E4TWFI5rAPprGZ342kltL+lWzW9uCwQybCN6MYCvDYcDF8Sr+uxVnwR
Qs6SDSamy/eY3+ZfbVqoFvq5ERvGnlWZ0hQ3OAWKeknmLROjPKNzrKMbzD8npLxt
7GNhH8/y1SNZfEe2dfPSh4PQ8vsP8ye5os2Q8cmOwASHEvypJHWpWe61wv2yE55R
HvIQViCcLBzNBQWXlloCOtZ53Y/RbsWYktl4nHnMVLPNTyFCUXhZQBLJpDVFOu0l
scCnt6sdAwgv8++GPitO7Hn7LqcioVYVNaAcyhGqJnFcT26nbT1dzeSwMkSu1Fg9
WfuBgyHA//GxL1QtaIAb80vYJqD82w87lEs0FLbLYW4Av0Hw2tbhIixPx1yXQttC
3tLdpweyC11u6klXatWt9dtTtxS6dym9Ng2h6882O6GyBHbHl9GK/NHkXi3EYpZR
jAPS8x557TJu2HfDvb7fLxzjUJYP8IIIPvniF03F0Zir8taV5IXckENFjs2hYn1Q
ID9kxLcUEm2nCWUXBS9eQoQD6xqCHGUwWDNZi17aEwQU2S8HMDVyP9CyLjzAdJjt
cpvn9pvXBrXyXf92csFV6Baus4ZKzkXa5abiqV0XHqK/Z/vI1i0LOBEuG+SKn1m3
ZwnQqTUDVqw3xt1zjEuYAMa0oIzIuP+sZD/9vOEMEg9zYM5c2xzo1/E/CpPtmiEk
ll/dTnSYwyQhiSfj6+Z1PLoEh7y33I4wO+OkTdlIivVwDxE5Xph0OfpUKgg8LW2N
TabufYwQtZBRKZw5tczPbd5cpouVFKE41z61dcKuw7aPOrhGnJ/6O1434TH8xP/F
n5GpekxiQ7+UjQa366AkvlMErKwS44iCvmc/aKi9ch/J/maeC04ceD5Lyb9c0kuk
NLlrDOGehPq2OoBA5/TOOsHP5SZfXM/6ww4VWsoWqQDkkZzRAWbIFtydijowEnev
baku6xRIH1ie8EaH2cXvN5yfJwfA5pahUIBk0XMwqppEDNrucNUr/GVDTCFx2LN4
2BvaOSEtpfHUuD1FGm8NTYs1Yh81sLxw1xOmfuDp/IPztdazOuI8QZJvPZzotqKN
X6xH+QIk4rNcmAXJOS6PhxEzzOCgT2hfNdXhrEU8rkyO0D2m7nwg+NbntY60j7yE
3Qul4WW7CAbY9X87IzPIkxdujBrUy1khwVobrWY/z3t5FWBbk0YF/z23DS9LEPVs
kjyIEngR+eAY4o81J1iDR+dYz2NiJYpMjmEVbkHoZbh+96BQa6dWO/nyWjvkBE7P
S6AFyoNjFjPAbiB4cvrHZOqb9+ofBg0ULmS57ml97hOhWWVj9wRQ0Wa697ZGpXw7
NB2Jx9sOLsAVLUzhke07ztskGK2t5eqODMXiIV4nHBZuXQPdQhZfejyogA8CUCYj
Tc2irMeSOiJInW8l5ljd8MHDOUZiZ4lvBQ2SpIhXRrJNVudRCyGKebuhXTqPURrG
ufKHo3CVazTXl1OIzYmXUGUHQ/rzttQd8QjPg25nL7p3Dby5JWHN9u6ly9fvHvV/
XX1iz66CUHLR++Cy9j6ZwMHHekatLJGEgWprwfPWeqBaRd/zPlYnbuowZ3ylrohw
yd/livwz1jeT7zEOtOV0hAVSO1nIAjrKLttdIgQTEwJAkrGvEskrHkU+Bk2bpNtx
71ZzU0yKCL6K2FBvQ2DepD2FHFrwBn9/9qx7VUAMbrQrkPYiEacIzT6oQprtHmbW
6oTKzrIsOys7nKzP5RE4IOpMY8Sr4f7gpeDu8wM4KWcFKBdJriFook7iT+qTxade
H/KLEvGl0IRujbNvIz67yOB/vrYExwafOOZTzplvid4COCKKBA+d4GTSIQQc8GOt
ilGZZ1SdoYTpxsgUVdriijGrhDzPnWE73BXaLYCHlFeF+WRG3sUFFBvNz16B17P6
u/Liwi5n1U0DnuqDJkXxjyq7SkUUq9gePXXyJ/+7dieac/v3GNWorwysFKC/K2L8
yt3j67cR2i4ldZyLMMfBxHptN4x93Dxq4l60aUoTZz+JUikogAgS9YE2Yhhz9/7+
utjEjRZiB8ZvOXOY15b4hAvtv0N+0/vY+aAVhlx2pAPdIO5/o09hfBzn+ZUUMfsW
w3Itbx5bBmatIPkM9N9E2H3oOGjDoxU0f4cedh0AEoLVXEj/TKWmKBogu3F4RTdW
fSVa93sxaIhY2j/WGwQM6PPEmjsZE9oQiwl6fWIKUBsfWBknZb0GkcT+PMwlGxiz
LYC6E4WtrZ17xm+d8Sn0XpM2HreAlA4A+/953X/iTO0KUNHyHgGG+UXkREAjXXnW
7oF0bnEMWYbKg4mVD8WtefFxStKFS93aZDSLxYXY5K4mtT+8bzrZeV9f6MK72GL+
0Po6ewYmNzoQ2oOmWjrzCiUkf9/82N8+Zh5epUzX6DStMIr7JBkaQgYI/CEDKdLj
MdhLo6GKguTCfe/LPCALYOzowqujmHbpbkxI/LDjzlG46WWUaPFmZoRrPkctROEq
YIouUpegot0Nx7VHQxn9Oj/zqgFBwf6z35iPtO2NcpLTAKqG8ZuwBet3trSoTzT7
I49hTPr+vi1HcHx7nNqedQsZXSQw7wgCSBPt7s/BWKWf7doPPxYsWC+BQ9DIIEwK
WpIHSKhaf3aGu+pY0KJWerVQrJGMrdkAGQrARUaSOHsS2jc+CrO3hwIelH7UZnRM
IJAakin1AplUukNYBwDWbzs8KgMG88a061vB3YuHqvE4uErSvekOuoS15bDOKrN2
KJbLZVSJY9qBZQN7I+cuOdeFLHUOHFzBcm7A2llQHZwwL/Z8yI9MsqcRuq7Dpvnf
yZC+5zYRkSnUYAazSnVFV2YNf0w9LuPF8sAFsctsY7GUKskxCB7GUkIbSUuikMbt
hvQU+IN/OkahraftgIqxenuR9afA+p9eTMkEXuPGNfdi7DpWYnEFXRVfLzz+HzId
X8hIf0V5JqSIjhTaF9kxBe3csgPfJukm1Bw1lawIAjG5/C1F+eIsqqLyK5+iF9d4
c+YzUZu9/KJK1NhA2PSyQmeeK5fFv8tUruEM4WSIvwMS7DO6VOEZRaZvztti1fBv
bjhWgdEcegx0yJ3uRgZGo8jb4/LgJvQHZ52DtktW8XKhr2i5QcWttSNEbGML0/jD
+WA/LherJ6VcD1+qGBEuem3N2HCHL+F193ybRAMdH95QltqnaQw6XMmrumcIvpcJ
cSS6hwCmn/xzTgD+4bNKuZvQSLJcbNC0K5ZqSzpcaIRrqouJK1xhekfxSJvj9oUX
iez9haoFLWXF6DaDAJk9bniBFklHaq2hq7Gof3Nx3guRXbfvT5yYRzGhBKTxzHFh
cdwr2Pky0uz0dEiMnB3MUr5xkoRmqFklX6bTNs8c+QccXc6b8eUalc2GhCkdge/t
+/lI/aKbaBPRj4Z6m1TNo8GHgt1sCAXwrls8ByKzG5+wBAaX8Dwh84GiKII38X0n
ZTnomBkwB3KKjPwXD5Y/RTBp74PX0alKc7IFHRmeOirV7Vf6FaL8Iyu+iTQWhlAO
/7bs+67RjhdGB8KJUEWoaz2zlKHg90ln9v5BeDeAPGSP+RThebB1RZZpV9sLXSUV
v7EB982E1Y95UUpS9ZhfXH6Fj31eZeunKxZbv+aMES209dvseU2IRZBk47tjuc3v
XiKvhxqbDsKtbS0rM7Lk83EAePYpUNlo6nKHt0NQFno6FLpdFT5lDw0+DgUtlSfi
QVRZHBoSoFfK/1Cds5KTOb7S6Z8WOQ6P3RuzlIDa778qdTRmMUHk6RUrjg7hXfAu
qqPISrSChOrUGybZUhTPKePfQ5nAZwZI9JvJ7NlAEHEAcH0lIqWN5tYUEG1xspmG
E6LW9Em6+az/RzEjY3dEQdUh07Vf59xG++RdqIYuvNH7RZsFyjgmIz1SCQH5zkLD
KdV00f1A/bQhQQjRtfUmx2jG7s3NhaRZLjz0i1mtOgZdLjII4YFoZeyMOgfBUMNd
jne3hnO6QyY054JKAYQQhRI9Y4CRfvLXjW8YoOmygIu1WPBJcSEfOuGm87SC164f
iCRaxS7G6ZYTl1Q9L0ursqmLXdFoKBnEIy2c21xPN/zuV4nJ+ATWETRPwUCx9Kkx
oa5QFV/UPQa/5JPEvrWUFpLdzx/2E8gxoZFS5/pmCMyf1QUO2MDcPfONMB8p5oaM
PVPwHZT9R53oZQVgXB6sQX17ViUbMK43wAzb79P33kCdh/4D6euQfXee0q6oWtqG
TmUEBDFN8Uix83uBArPSyJpD6vRf/QK/mLCz6R2EDd3c2/FdF9mw9dGGHgox2Asc
G242wOO9oLeFYdhbp8GPmGkgoWYl7z25VdN6gnzhGEDIyq8tugpJFv0TpK9Yw1eB
hSQWKmgmVEl/yvKq6lP/wxbPpK56BzYMxQL9GoGwARVddlGXhh1d+mGQzvuMD0k3
YqiBxssDuqW7tS0TAzqoKgFJ5G2J4aXnANyW9gU5p/VpPx4mJNvppu0AzmTV25fp
02L7Gdplh/SSgVyb06hCPyPbIBnuZaIZ1VmBMHYzobXMpc8xAu5Fj+HqBwyWEIQG
Z7hZJWSGARmevR/OadqmFOlZVH+21oOuvzQOD4lg0lyUIT4+0Z86Au+ZbwidwkZx
CGAqE2M5w1aHv0wdQ1O6zICX2dv1dY5rlf8WZzyqt4gC3xi1LihYRmHuq4gzelQm
8XYp/0q7mD5j1NOJEoCChHeS64q1s4DVDrc/dbl30k+7IO6z9gbUQHM/ab4Lafv3
J8IX17Y3tZOEGNc0NhwP2b8wsYQ1XgKVgjuxgmvQCa5NsqHOssqAn5iLCC9HYR0H
qAmkSnop4BhSlXG+IgPAPDaf+LSTs4TWM/fb/e1tFeQuyslomI5DV95iEVioHVc7
AwHJlfnVMHTv0zDGWtcJqE1xaWfioNqyXl5edg6FCrbZH+1wisr3wOd3CKrZjWeF
fB25++36+knGnOyaStbxwKzHqVLLjRrMKoM+f76NN7klYx2J70FvvyaPq4gmQUVz
IP+X3TdcBgLcafzPMogkxRhjWcv1LukhSVTqQFoDus6cv0VwvQpA/rZHzoUMqURw
o2lTnw9gR3Q0pwN1+/3eQbbWJJSAGbeANNL0/V4GRrNwyNrEncsTGdKuOGooyYm5
kBr6nh7ihFtybBta5SUEtcgNbn6AZkgtY7SQ2blOW3gtJjPmZrbmP9M2GAaIDE9k
1yLojgSyz/hwdZ5yj7bakL+z3ruDRzLZPug9/2P5LIMkBrl7CfesQPbQk6SLdNGH
CvHKfzL8yERfxYlj/38Aa1+6hYF3+K2EXm1tAgggiwLtoNCn+xXvCu3WyfBOn/UP
QouOl8t/KeHusIALYyAj1SBbfKZlaAF1TkBA4QyKAflis64JybTtvUxgrOPeFiIW
LxpEKTwQhOmL6yH/nqtUj+lVDBLzYs6WbSFGDmLTOGvpEx9ydapcNWnRbRApbn2R
Um53ypVN+C11ZuqvcoZv2JCtGdWxdlgs8kayn5Urp2pcj8fKxDGnTkZVATNCAqEp
dA/eBoB+Gw5G1L77jo3vXxPdWIhPCvEp0BEvPy1Vsa1FcS6X7ahUp6z0eMCBtJ+4
cFZHgQcHsqbCjW1Gs5fEbVUrr4JmEjGh5RlG3AXxpTWU2y9jb+6rrTnbkgs4MNVV
DV1AquiCAYyKptK9PK+WfUk9RjZ2nGm0ZbXv41m9qseFhnJW0xV/9z2fV5eTmm+r
BiSrsI+JK1Gw49nRn8h7gwSNqFYELNyTMmFZ6Q93LHpM08En7NlT6/7Ym1GWrJ5m
StKJWcIMsCbSYHaZPP6yumgugiG2P4MRQkjZOpDRhu0kSx/nv3mpz5kuJKIYnWPe
RDEpzpLvUzAmdqPCywAQPXUjNVByFk/LB/+/m5XdSPjzo4e1VaMYkANT3zQkoGag
nlQTq4P27QZjPfuPYNGQFWg5PGgO40nr0iJ7nn3qMwiVdhOwiJbjF0o8xTT2ygxx
bKdgyildXm+urRR/JixUaoB8TJ50UXg+8xxKYKI8C0zfMUwYrU3o1qCkWOcYbAS9
hTRhesZkZWjBElCjLSO6wEzSIP49z7+aDaSTcR3G2wVO/gI6JFQ/86GuKvPhPuT5
ZRbexXZbweTAPboLggaeu4VezWSYCi2Mb/BFct7i0WOMHUSjNiMgQpqV8bnzdAkb
tkuYgLxuosptj/Pfh1F0YWRgGIjybpriB+jUU45FP7UPDqxnpA+ighKVbpI2jajG
V+XymrPt92+fxSTC0dUF7QhcX1SFI/j7eyOjywMEdS97drxoxIC29F4R0h2QIjSu
xvuJf1D0ujzhSfbYEHGcmVm/DWINitSOrbfUEaPMkGCnPgs+egX3ytsYrhmOt5OR
i5GnkJOCbiKIiDiMRjFzHNuEBvg5/3aZq3FmUZJvqGQd+W1XvbLwO1csG1ve5uji
9CBlY1yXg3WabLS89FxXZzMtkUrf1VI5hmVDuB4ESUH7WQ8oV08naPykPAoM8aiC
65ggRdHNVdBPLg/GUbD5Jek2V/08fUik2RLebrL+dU/xJV9lS8gyT/Z51Fro2x5C
WV6+m2fHbKURSfAk2vJIezlaeBsnWHnw/DDUFZGkHSIhg/NHZhTxpaJlXqj+rshY
PV1HNTkjoUAdDR/4sx5LYc8UTprtpDirbA3v6jcxu0ftHVfdAUT3S7m+5q8nY7/S
Ug29QC0BCra/Wx4HAt/QTRkKFJ5NlcKsHIksW+TF5GVf0LuQy6ebZ6W+AOu56Nci
7hK1YhbXwasOADziO/+d6K5FemkxxWMXUJ95thlkuN2LWFG0yE8KLhBnYXeILNB+
DYdtN5IMG05ZeIxVeyO7EDe/4qhA2XWLbFQnbTqra8cD+5ekcmqmVvg4Gl0iGlg+
X4Op+JO4JeW/gn+6/d8FESDV3QVuklTO4zRWyz9Jl2vTcG57AH2sTU+NFv/VpLMg
TeYFFWHWEc2up7KfZ7tumx0juXpmB+L1ojopOAsS0lNiA0TnMx5qS25uSq2q7/Ir
UVlyAYTI4IhzCC8h8iKTy6EqIkYPQP9hCJt1+4bG+sSDj4puGA8TicBKh800r4Or
AGBENywjBISOzE99+3riDULBctM16k0+Au+3rZXBbBM7OGAwc2fO+/FdOXP0TqFo
IazXVzDujXYBXmGtgl8HV8mfLE+AC2G2tMir2lAPZapzIkh3whiIPRBlxB6rVF9/
PjJl0tFi8eWDF56IU/KZLTagi49pBavd5Cw27lWolT2MSGOBJx+VplauP9F03YXN
OZS5h36Fl5hOTHnp7BfMoMZA4K6IcXGsSTgbjv3V2fTWbHef+Iwh0ZeRyjHknFVf
mjExijVjsboh4vaYkLwL7I2wPdDP8M3dZDS27DQQa9JgUpdVLmLctYAgcv6oFVtn
kgg1z/UEZTA7axEysscD59zZgaXP5VJvpzjzoI4BKFNTCT4I5qfkZJsnlViP73h/
4KtAhbYe6S9mxQ1vfttaWpXWxF7h/rCIM3d37lT1kBVk0wWh5ZGDXl5kow1UaoYk
1nd3qc9LxuAIbpEjxQfd9FWCAuDUY4uSn4//QHqnCmoWMtr4ouI1Ye8VbwZr7LJE
weD/Enfzz1H91hp17J29i36CMJRQKLQAJ/Fy06FuQNIt/EuYX0STog9CtccySUXO
cELvIf5+S6tLV91yazwudFMa5sGW0o/0Xgr1GP6WSY3gba51nCYr2XxU90jPp1hC
rghjx9LtnLWPQOdJVaesHXMQopb8vxCoADeajEYBjm4wj/Ds4EPgVELUEHh1kHGL
HH8HPKCovlYPSgIOgcDQZXbQVUq6kPj/b5JERfDSWe8k28qjwy3gIeTzevObFW9v
tcz+gV7RWvYxRmNQjJJvtLTrzFUhXG1ArIxo3jApI4d750MU8XP7nYMvbfznDupX
XxGG2U1HqGbnWprHkt9FXl/UpYFqoXmUSMgeoWpDsna6V0CqDnM1C3thAlTDANeX
/uY4Tsi+l2FkXNjCjrgyQihxLBKukiISNfL1EUwjgwEeK8DIcUg4wXZu5H5brl+8
iKX2GWf7cMMvKUUFB+imituDB90PBuJVcwePxWPYzl/TTNsh2mMi08/wYehWJdJa
Ay9e/xizfa5j/gGpMDJsIn8TddmtqXATT5GgE56lRvVmkFCmg2tZ9UxKRm/352jS
TLictAaw7RjwpRNlD7dWA+Fvc7gQbVUmU+thIpl5qzwBOMzHSX5l6Aho4lcCe+ll
mimVzBdGXeY6rZsASseX26Lw8OJzQXKosC8TyKrq9XoBePh1KTiC2Pe3wTk7JAHk
ptbyD7TOeuGc+MOY1lvgu2514gdzrphypvnfGZGnYMoTe8D1Tz/fJaTb/1hYAv/Y
Eok2hRJgFNjxyrXsiZbBrxfWl86XO4P93ZPYqxTWMv+WgTGxDbH0Vso+G1eatRPj
6XWvHylcfDJpc/rx8OUvj43XuxneWVMcqu2mZVKERdwOXjePjj849UdcfemZeMjq
XO6yhSLlipKO8I07eRslqNsXWh2cJ95GtW4Iw2RB/tvKBrNKhj+9bTLER1ldFZKe
GgZeKMO0amhT0zCio0YndGyJSYfaslv6v3oNz8IIyeKlrdXmkBnxRii+OPjGTlji
Uf+LWObOnCmwjpTo7kPJ7RX1+NXgXfmgJWtz3Kz/zZEbOwhfIHSE07svxVmaVvtB
1jX9sELwXNpZ6Q3GCfDBxh6qMipnaHzr5coNyBjc0vjzoKIILj61sOx+gghTr4Tq
2izNdUbx1ISgGHbEBrfQuScVxLR7MAsr7BTsrd39glTCTgYFAOSRxhKXQDD5lRtx
Mnw+AMw64sLMy6AL222+jD41v2HFdzxuqsezOstkoeoa/oQbwU2s4d7AiEcg9cp0
+P/MfC5tm3AsgmkrcevUHhXGnAUi+1IpQTjRC4RDIpnMMJnbCBkcDQlisxER2d38
MLq+Yy9HnJgpEuY1btk1e9oQkK9CDKum/zRHruM1z8SUUxRThBsOPeMadVInHYiR
CPC5rn9niY9lgeit9Rfhiv7MTpM2hPTtl85/hb1kYCXagSYGPZKNQgbHJ632L5k5
vbQoPFnQ1AYbTbButRiNAXc097fypPTDVMUFhRNy+K75uJiPfOCmYM7AxDxn5mRO
466+Ox/atZ4p44iziXbLKTH12/RKmaJpN+PEri736HHSE1H2WWdld4BBA3oxe2FR
V0jmve0Uxzk93ewowGdO2PS5nVV9+bllS8vwqNT6y+Kq8Thc8z5w4/Q7AY2aU1+H
Y6eEQFHhACiX4WE/IqpNjD70NETVcq6MamjKrWOG+tX+8et+oGr23bo2yNoQZ/JO
WV/RI9OUwzzkdrKhs4fleyzj7KowBEeoKsvDgdR5j3yQYtjXx2uo5gimCIjXrW6g
4/+kcYiI99/EKTeGdBqNh2R91yiB/m7dud6Jjhl7rL9ONY2A4bZ7vnymJKzfHtFc
GN7TMnLyFW9rgGhklqNXqUk5rxX4ucG6I4JCjzzLnkBCj/o42pXf+n05x4U27j9W
07WYBtj4v7wccQ3fBKIj0hotdt2wjo+IJhRMeG0pP11pv7EGJNAWuaXYYX5siu53
U9x8J88kHUzAHIY7cf1qF8WCxEF7IIZZ1/IFUNq8A2hq9hvGf+BAF1g1MnSnNF+6
PHswOthFpOdtxDkkcX8lb915G5adMs0boClexzpJePXOeBXqLZ618xu7B5SOQmWX
O2DH98iAADnLBOmQ09AmfVrKMsTsDUoIHHi8vHdE7IuU9TobncboWApeo7UQ1vTE
kDejrUYC884LN5U1F/bFQOVpkgPdk8xBY3nbNsF2AHncVgiQHDoHseSD2q5XSHf7
k61r/b4GBemSC9XFcZT8iCBi6IU2tuXQ0uocupHr2Mz+BHmjNAdwie7IeLmSYHN/
PUtf0VREdSqnL24OdgtDPHT9bjQmUguTOZyea6bctpNvYKeZVvwWuFfNDAT/ufbx
GQIgoqJj/gs3FqIIeDmXncrHMerjCrTgE9K40dXGVt0fD9vfIvTRntQVTJPTQKxi
Wgpycfcu5X+qGO/CPWBdstXTznpikNz6aII7s0Es+BqwF+mJKDdyPbYELRrbEw14
x9+Vq04/RnxH/RKDolEf+hAeMZNBDUrUKDOqEvyBRX+2garAS6OCRKfUw4kk9CuB
OXePY3liBMuKOpMLXxqHeh/2HgmgTuH2ViBnyBLws4Ofx7yDg/XKUe7JcfLDtogI
y9RyprXaefX3cLUAjAt3A7K/qPcVn/L+JTxbxgJCx707kDs6+01lAr17R/yYmh+D
QW2CEj91TDUKQnl9QK2pZGviN2mo/lLwpa/34q7wFb3t5pl+4BxtbXY1JlANf06N
UwmmWKjaeJO5B7VFkquGZY+BRVxCgq1bD8hvurcJwA4JDmQgGn33AaPvNq3e32G5
1mynqCJJFAGuHTtg56R9OBQ1ybSW/2efFm+qQRIqInVP/idGYjFYY1V83KLxFmBO
GGll9kIuvfIgW/EFvrwr/cZphI4r3dyPYIW+meCjnAe/pUpSp142TXFoehFu+234
QGD969wXpU9r/lrTwaveptpJpSG4LwP1oG+NoQGitLXvmLFXAN+elNopMJpqoLhA
2UnfYjk5KhIgZ25XxYR/ygr82I4iZ8ZlAFhIfCkFwKDHIsL23WP5o5kKbLcIjKbH
eDb4bgzLbudFEMCKeggnEzw/Uz+jdGti1dHLYOlHDihEl/99ngUxQ7EBGaPRrERN
Yq4EuJO5LCmdKIytFOHIrjVfYMRvpwSatHgCMovt59vaZqlBWh+2PQcLUHpf2dtx
uJslgFkDSWRfI6LBKuKY5SGivwXwLE8dMRSWwNOahTdCXKoUjvUq3Ze+Xw/pHzK/
vZCWYTckfc2kNi0xRIbfa94KkESHi9vt96uR2tkTOudcRMtd25RcB8x58jpR6tT7
KD0uH0R8O5iL7x/ZWJ+MwR+2F4oJGiu94CUrgeucYvAoA8/64lvXNL99ud1d5Ilm
vc0nVn1p0RxkIfBFi+Gxj9rwN7BdkIl69qjbj9luBjIarpqfxFnVZecSvAaUDFvT
ibBKB2rp7IyVrGkzDcyIZE1PedmmKjyqQqZDxpUsnNTkmDLn2+/O24HAgr8Kb1Od
ak/zW1tiiVpIXipTxPVKHsiuEkvgrSohY4PJNDcxoujnMCOD+EFVPHDL4n6hvNnh
agyqeljhHZjMPNaZvjGNdEFcD9ryWMQb2pCd9lfpuYPn0ubkCwvfBpWy1EXQmRzR
bTqKAF3XyI20/cIa2NPFFcWPpRn4tDWD/1HBakATkUyqQvnsLaMqA38KvRqg3icq
9SVbe7QIq6j6Ih3pN4XACE1rTUw6lgwu/NkbOqP6GvFml+8ifEKHZBgubhc1KcEy
rzQTEo7IHu7+UpxWfS+nNxsXDRnJKt8tp++m9p1kWLb96ROuLhD+3ZAnfATI7eng
iPneXUn5+uyZBiAWwRtjr95sKLkvYM/KLhEzzGD3T3DKRAC2eab2P1X14eYrwNlG
C0hSFd0HHpp7KJ2xPoLFhv2v2Xhqjhpm1NdhezloFjxlzsKOtlrwtSgm2PVZiNe7
U2qx6SSOu/Sk+XiNy3EbGfG41KJADKkUobqmN+R+xrjhdwQ87QgzRh7ZPJmri23U
lgsmq4kbmj9UIwEs/GKpeqi6t0T9ou/S1ljg7WSUOLy2DRBV3nj2SO6WI46zHmlV
tdtvT3vK4G40Xqk+Pgh9C/Edp66bypETjtXzGeUeu7Z1r13MucbkH1HoKjWQnznH
EJs6N5F30b1UUHiJvGrdD10JLZw4AVe2xDAeCrObcdY5hr6NGh9Eoi7oIiUEuTjO
lQX7f5sksBEJw1Q0ajRlyvQowalWv/FVCr97AVE/6z4mWsAxzn42FJsJdqMHfM5q
Gkc8ZX5iRQqV1Ds4Q4zP9w5PaxtzZA8hVg4nUFUZSLoNDQOUUzuUGHiKbNgwF2HR
bBqX3v0Kd5gP/0+J9qXaYpU++RLPeQDkfiah3UiazULVVoBnA/VA21A5vbAX5qQs
SWU4EcDFXjkviAxCOhY68eerQLpXEBV6O3k7Q/+ZQZ/D34632DvsjJ9FuK3jpuGp
t4aQV0EfdmTJbmuDpfV7pcSn5iNWRJIHkfiArTlPeLTHzRxhAePfaxwUfnaHadxt
ks7GynXIaR6jYFDb8aJexPAxa0JRSbMuujWXcHGh02sfvE51yGM6IHttZ9yC1/hX
KbHBqTH3+2wI1fUFUKslv7CDmuNIMJQmJTLYsrjEdVJuZP4FjEMsQZkpxldbe0bC
IB5P9jLog+7ulIcq+DwbARRIeq4sSqKw+UfDXF7fygQtpQCg2jv9Jt0SR8J8Qb+H
OO34bY+cLU4LYiXN2zpbEpYOkHNkHV9LMONa1JVuHG7OGsMzgmwHi4ygv2MVmE2b
RQukD2/720j6/PzMj7Z6R9MZ/5hFXZ0fRDoguhA8STMQqvoKtymTDHVbLN/9zNsy
U50Tfh35YZiNy4r9boeTrr9/yWCqVEJi9Du0xhpUH1w3ookskJDf9uWaz+ks5k+W
3whJcMQQ6FPni23ystcAzdKhfCJQ8xWDmE9n6yfbDYvGEWowq4KUC2ESv9n1hlRZ
HStu8x5xRtyNDwPAXe8XYSs7JSoJW2/8vyS2D0s27raCJKmlD6uXOSO7bITTWuLB
EPFPB1KiTZ6MoKzRVND3/uKcMcacETjy2lmwyRnZiuc0W/TxvCUCTnb6nEMQ9Q7b
u/cYcdUwfVpNz0KThr0LJtLuiWKrq6U4Dfoivp6DaDaOUApvA2RxjLxUe03veS3B
1mbawCAKZpa/T4yfAgC5XDdnrVWPOMcKhSMsIut2EG8wAC0KhOu95OzghwgF3x0W
tGoIYoFyn48rNY9mbClifItbi78uD1HWlIOhOkEPW54bAlFpq4mpfMaUeLMLbF7i
U09L2xu5ABYjJpAlfE8hl79X2FPE/w+jkVHQRWdIpxgg2c6jczNKufyPYUHT0ctN
R8GM2/36ZSCLimjJct2lhovxHPT/eZAWq+fR0bxEt6BVve5NSFdy+F5tM0RAO+EV
Kpx16UUZeUx/XCktOuwbE7s7/43u6Yr7sefmGk7+WTEpNesdiR7qUI8bZ/f970gF
VklKhMmrGZLkL/OE4pL68ynd8EnM91GxTcjBnsEBAcpNUyjYwXzOOHlHLJt549mU
roC3MHIqY+63Fs3FDht7yGXHUnWjDmPmqPGXIehCaVm3ctiZNjsWY46EQLQIw5aR
qBvWyZcVfwY2IjLafBTxHm0DT1b5AmQXcmSOKul8AZl7Fho64abkLE4u4QepVjt1
kBZRS3DuC9jlw27NA4LEzrXaNLWTPJA5DmNVm8+5+WQOT0YMQjRizcnJVz2NwbSa
EDdIit5nHois7OA8gYoaBmvLjcNWtz/Jv3KITZoKm5lVUROq8nAN+ZMJmHreyvbw
sDwaujlP7AuKqRTPkaiCqq4j/DCZ5dybh24lPHu6l5FPV8fClyqSfanMIZjQK4R8
TDVe0i2UrGgS91cRZcexS/ZfYqxXHRaW4IKegu9qpn2oZpus6Wow5aHC3JBMlOaT
QZwtEKGpJFvdd6IgjSQ7jL+gOEum2B2APtKUs+0jYyzq9pvt34y61vApXrbDbHlC
j8CkX7ro9jSvMCtbugJiFQy82syoVGLnPrr51MQoXyQ+78rcZcxIrI8KPU0EYGb/
ifWHdV9rvSOi+hz1/f46YeuU3ma3Fed6cL7PYLu3HZSJjROuK8RkxcvKQ0OXC4At
x3ZQ+TRZQvfEgh6ZNsBKs4clfTSrRScJ8FK1AR5sFhMxtNynaamvUQHmryPx14WN
6LycJbWImDNU9fqUqbvzFMfPU5TI00zLgJIMT2f2Vc1eAGfjhU4I2PD+E1T4ZUdc
rdTt2KdULHYA5Vx8J1f0lmuW8Q1E0wdIZQgkhKKokSMpnaEyeyZaN8YRm5zFuewo
IVeHfF6iRsZymynUfbCoS4kmijzvKN3MP/7C3VajiQ5Rt6Nz6OmOzbolcgSScDP6
+gXAuSLYxrN8G5h2k4kXNUlHmy4mtHAz6d7zZtOXdsdVHKHkIjG8cwt4re8sxs6x
TQ8RXsysSDbAfuSJz8+RB9dwQPHLov3TTuoOARM/Cd2fRZBpsMT+RmauoE3O/IUb
rY1mWDnosZRSFoetxBKHkEEMpEtdwindVZ2DMMOi2RdHxh6qb3lQdBuz3/+8hOa8
mLNwES8rWpetbgkc0hE9qAlyUtrX6N7Gn9/ZY81PXMvh7LtKiRPdx6D64Y8MI224
my6EQOjutb7b6+T8sIerRiCQz3rozRtnh2wzIxQ35fbBsB0SZKrjrouwT7zpfnV0
D7N/bniBNkAvOTCwiVjtcWWixazNYzGBABXj2vYQxHMFaRb6Rs0Asskz+Yo2V4et
IAsHYj4GVY+D3E8w12SZNMG4QdA6SzAytONxka+orWlYcTq/RVV6tUabQR7Gt6Yo
YZPHk6TcQhHR60SthPlg0jgC7q3PtfXZPKKbOC57Wrh8CW+mnsH+lHDf5zLX0dHX
YALKGpcHqnJS76c/imhofSgY8Z3ZqYDKkIY9BZVhAxkWHQ5Rrp8LkL+fs3vzIYc1
fBhgGDahUJFAw7eGWi+YXQ2eD8YUalcvJ1h2kiYJFQEs80MXHC+12PKOtD/d1K6V
Itq0C9NNYXApksav3ntEm5M3V/Am4V0/mrmETrGWZiFagJbTvK1GWxwQlXzMDHnS
NzFQhYk1dEMgd8v/drnBW9tqLMPabKELRBSQB8SkUZQKAcmVwzGa5M+AeqjeoRGp
kAlvMSueM04B03bETt/+ddSZGGfddWup/ZGy+lxDl6CNNV/sXi891KOAEzLIlUMF
cT2tl9YsQBakJnRozIKxAH6KLnqB8C1Mr/ZGs1sVKKdgYFdjiizz77BmBavEGPLM
1qU4g7/hJzpKHihF49zXGsdob7Iarr0xGxi4RLtVq2ZRkpvLVmvKQxEShu2oayvf
xzwJeBZO8IuJPdD11XrTTeTshSz0gx3YRPn+g8oorsRAOywwkIi31TT/S9VExqiD
d5xwbNITrY9BGMbtU5hGVP/VoVEhj35iPb+hoYwDaON3rjdi7QAEMnIZjKEKWibI
JiC0qMdEEHidKL00LXhND9hwuuZO6WtxxnXYgxxDX5Dtt6AEE+1QQFb8IXPbMBKa
LnuoS+HWoDkXeFcyHrXEFhHXf7IR83p14nVDFpbtTs+4lpll3oegmNaAkpcjhLm8
eP2ictjnUvhJkWnLx1XPfXDIiO3xDc14k4cKwurWDFEQy46uP1ltvxI/nSC6q+n1
8CA6yQooSqWIB7WpkdVjhz7+ggww/NlaToQ2RCxobdEnrbe8t4bQ3ruZ5ixaSTRb
twt7o/EaZzNbWn+DM48V0PoGOPhRej6CDbqEPcy7r4q2yS9OekXD2+2HmHC3bWp7
KFa8IcwSMYoy1S6WQrVswrqhbTWq2MKMeo+yf3begiQgGMAgentrCsKKfigK+unG
mrZj1MFTxNy8U96qZn0opzPYEj+p5zuUU5J3rWTIy4Gk/O1a/4HGpiLLBY6cMiXZ
42cFHJuwF2o9niiYUS+Igdv0hB3sklYcnCm84cWf2EzxUYekPCtYiXH3X1TKpgYH
o+oh1K4mH/Gc+cMbT7aj/D1BjoaHbMmXrG2YmqZaZI5Qe7K+F4ajPEE5LK02c/7L
yfAO/gLE0mKnGLM6RX4izV+jP/0+UEKHV6yJFeblKqBLNLpZFRBsKkUNdeFU0AN6
Syc9Kwm8lEiN2u4YYD2ykD5NSM32GVzvyL++objzTaMKjrYxUWFCeSoCv5e1Jhb4
jSMyPQAEzJJDta+qkGNdxD8t8cDXKBkF6fPMKa7qb1UlJWGEP5unt+uwURVbbXjN
nMx+PeaIFNtGkCTdXYrCuWXHWh0ozT3g4QU9/aKabSmvTg7+ou25QFAPV8xqdoFm
c7R5iPiimmmtCPbBURgBcbdEv+xMo2tArGokoLO8mm8caimrN79SRtySGP1FvLB6
y3h+k2O/aN/3kW1JEOuLGQiEDfU0ZAtAiiotdH0BcH99dyuWAUEgetb5tyt1K0XF
7yL820uBd5HPU8K4b7vHQbaY4iwyIi3w9Zm/oiWvgB2PtSF1eZd9f6JQBZ9DP7Nm
nqCDLHgZ1F6QZigNgOCtb2iagtRC4I6dbXB27aJa8LGn+dOOrSQF/QyYvk/kYlNM
lJJcvvcTfkJwSndwMcXA0OMF60BAY8GzXkSYcYYhxwdl22SenRVSNbV2Unuce60c
7N4mYPPJtFZIRnRp3F6Uk9rvCQjBf6P3GTWGFBlAs45fmU59ZL93xWvGB/pSboAD
iZRQ0IV4H5n1Ipha6r1oin2ZXac0MZqsqwO3+3Hoyef2f4Qxhh8GBBAukSSrY2S4
m+zjpSc4CRCrfkSm3wbVkZFQvtbL3t7x63Op8y4zJmkQF/pwAbtEqTQ+5sgeBvIq
6ETCKUAgHXLfahMfN+tE+3jv1KNwKrOjIyh2Lme3YmdNrpTozPo4IzNhYuCLd+Bl
DWbewCM5FRruGs9n0jI2W7xLtTpcy7APP6suvx5XU/Bcwy3cvbiDnYxem7iuy5PM
uqcDEewskj25IGQhDuC8vUL6TcE9JVlK+zUrKgZ17W8UFxkcntn+00MeAWr69fco
D7U9R8UUQebJUPtjNO4Ae1dJv2EatP+lJn5vu40+jDnXBgEDggg+eZOJsvDEHRxA
BCFOPx55+cQa0GeFOBDuK0in18cpYBn+mrO08FSG9P4PEK8wYoBk8eo0vvHySXXE
E02okr1BWX+TYgkqF2qMX0mbLSTIx7GcJ9rUlfFBpF+Ls22haQtxxNwwNn3xwbvT
cjBuPZToo6YFZ/QrmupjUaW0fk4cFuPNDsk2E3GH/5ys+CG1PLyZnKL2T6/T0na3
XybMS7/BliNhx9AadO3xUg5MDeqIfgzua5bhUF0gm+x11SKFZsgEYwpygl3fja2M
wyGNEeaBOBLkcC5PpyOYIuJE6A97ClAZCj40Bt5Ie4MTNNSxpEpmGPEbUR5VBfgu
z4gGkDYCTDJXb1HLrnryoCR3b3DeoEInbs3MfgI7ZouXaF1rDJZMccKsBsvFDYCv
iimoVR80bxA/tUalgXiu8SCi8YAQ/wdPLFqz59B5dF1wzyTejM0bJr6KWwrv880d
PpTr9TM0j7h2FdGGK7j4wK8pytjK0kmO+S3VGHUbuX6wpfv5aI2nMEY+rp9dlOCd
RiXsKmf0xKuJek0Dm7K6wT8toXlf0KfZ7M3yqcuJWJ7xiz3yZzEj5i/xESKraA9J
eGtA2eq7ETLvtVoTlncwqlPnN0bzvphlyalAbjQWhCg7ShrvMfI0s9UzmvLKyPRN
yGBgrg7lkexSVJVXVumN3sUNqxppXNp5T1Ezzuw0k/FsJCWzt9mSqsuJtEDF89qT
NVkrhhLTjpj4EyV8U4DRBEX8nZDe6UG5H/+WS01V65PrjapvyVSQKKF7OCkjhTGS
v7f2tAumsStE3kuW/uPthYV+uBoLLLMhouMv/zwDmmoiFps9Oa0FczUE++tg4BkD
mhqao/YYZb+mJ33xE0XlPKtDN4BDHMwV9ih1nw+TLldi5ZyLWKVz2JZCj2Z/6x2T
9xcYSd5FsbipxlXVVA2CGeOyAnXc2Lw1GL+R21c6YHQH7AVMTslXYT9vwkc5FBr8
Du7gE0v0GeAZdzC5r/81L9ULPu+aLfxt8GirYqcUpJeuF5+ItORLEOm5BukGriaC
ZCscTMGeU7cPCmhd4RlmWWv04UGQakkK3d4qp495Mo0/f4tTycVViwsYuNV4qAFc
lCjIdoc+RZk7BDFh1IfJvNxwZOT7upQUabufMPrGl0PGskI8K4w52hwm1eUP2fkW
i4kAKlVHzue1a4s3VzRbqZ2+XeGb/JC4kOFyBxc7rcBSdnoyuPMrMVFH0A4ufOj/
sKUWbS90C0kpDSIu8LHVIx8DXBONOFRlp12PAzAGR72WpQESFt4PwvfvEYyJBBoE
IGkDCUmnN/TbhLZK1VVemeczR6HDC+QsPrMNZrll5SNHC9Nk+NXJK7UV4RUTDMcK
L8OSUw7fJUNt9aAwJ98b8DS80XSLhUl36bhokWVQnbpmonRPP2b0jKw/KqA9eH8/
Eg5/Qb7lGh4jfX1dxS8bbPNyi0AKWT3swIq38ylZ81jqufL7DegYoKJDuTTW2CSY
HZbAP0s99o8N2b2V8mmMhy3C73LYRajI1ipagxvme+AIA9CwFxLr4bNaxo0jf9Q8
2R/4tHhJX95eQ9lyGZTax5nsfCN7DRMH+cAfvyMLVJZeRO+9ErN02qYF0zCSe9D2
oB83QR8HPGPG9IFtoFp9sXhUPtOuPTgXEJ/HWTii0X/QQKh2amyTgGTea8oo0pux
CmjJNSZmyQIKuiIG0n1xtcYy/HYwOasTDUB6x7db02KdV63JMK/eK7Ml5fspOKJ1
7t2dHOsoSxetNkt2WsY1S35hwM+ub5l0r94pUW9+VNt6DRXLHLb9WzDBf7DIWtju
BGvlZ9xAiHbw8QRaCxYzlHyZrad3z7Kb/qlN3qDx+gqjcURSbeJkFzftxjlq6d9H
4ejTd1RW6BnZ+KSG+96xVN27Xutb/3fRbPV46BpBwWwBRRRFpZ+IzUA34Ts1A6nL
84ph8wbmJKlG37dvm418zt6Gwee1nhy89rSvrfD6i98U+RqAYZFfzytfjRotup1C
b/wDkvMzyQvOkCMa7+6rsak+oztzCLo2fIrjNvUy7aTFMYjboTsUS/huYTs42ASE
UHGwkaKjDyBdT7UAhS2NzTeEvAvgP1/9lR2U2zMwlU20Q7O330g6LB/T71ZM9Hqk
Ruzhf/dF9XTmXUZQUuI+pYLGP+FGJHIbEKnmlhK2wmvZtQG47lElrVb06rZ5kWcN
7wKxXDp6bq1TQE1mDax0Z+T2T7up0ted1YyYQwZwFlmtWHD9BV3fXofhKMtCyuD6
z5RlInwF4wMuF9T7mdLn3oAkQ+yYdh3EIMYZJbIk6EkB8DZs9Il0X87wk+zm/w9+
B2TIIvXNqP2bZQQkyYcgjNiNfAQLhF/zfwPoBzkGaqNDcE8l5KLCjA1nd9ktuenn
gEdx56Vqc3ORYNaScuyDzWRX0G7QBWJO43j/6AcSMlUUJ1DUtDHvn/Oy0xum4SBf
h2Da6LtjNwqGbzMAspPp+kFzSyBfGoO95GPuMYHZ2tvV81xd/UrbuKRvZtsQxSlH
LL9TvVUyoBz5ti+aHJ71vnPRreCukg6BA7VO3o0aeg4UcpmM3Gl/09wFoT+m34Jm
oDo18MBfEXsFekGtPNCmBvaHLDVzQSr5GpTjV/K18wQpy95LJcXrysQguCfg7g8c
2NoQNFEgW2XY0AyWHv//ZCEpPf1kt4mIkWMbK9OqUFkiL2K1gKxv0l3lbZy8yQcQ
CzHwU3JNZdQr0aefv42oM0B2j0GmjlXebM91y0m6GBGmGPXm3W2fw4bOl39/olFt
3LjoqrGEAHrjteTdY+4dYph7gFNikXMjr2JLJLS2VkyeaI2ezrTmfYtkv7Ln8djx
TZDDQiQF2jqje+s5IXqYKGyKUZwNuHE5BUpL8cupakgOtYxs37+3eapZYXL4Mxq5
5/G3DCt6Vtk1Bx6KXGA0guLBnfTyqcqpjqYt54jSTvrvhxmFkG+MgW0cRxsb9J6g
H1zKqYM8b1xTCDvblBL7kGgxjMfaHzOwugrryw/f6K+nR23ac/5iUpTYUZi/H850
8d7XG9MiOnTe8/X1Kik3D0bf/oL3z3v3UZGDzB5PluGcaPj3qLTtLIK2aspvOIMw
0+BhIyffbapvBtR+F99AzJ2tbjRUFFbSf6VxCRKq7Gp5Pqr7vUpSYPDJr/aZX4tn
4Ilt7y0KZ2d1Osff5122eOCZyGaawjLT2Eiow38zdrIO0veN+DiRPeeslGPKns/1
40Uy1feGNZoC6UEhxXqw15hEu8K350HlmmoOIVQ1nW0EaWaDUZRydueh9LU2xXBW
8Ur60nv5rFG/tHiDyvpFICa9lwjYMpwjLYgl5yNWB/bc4eJogzbMGcAhsp8utPWu
HD93oWewtdKo2gTfj1DJ4QpnGEbYOyZbLwEeRC6mzkiU+Lka5uEXLNpJfNgDMPdv
IN4x1mJ+Pm4p5eN0VmVhgpGtdq37k9oregRHwDcV3Dq1PhVHLU4c+I7E4YBZMZ2m
OpuucJbS99eFflIaKm64dXRa5dUcJWY3B5C08+UeBorEf9vtwCQN3r+Iq0TxXh/Q
YEr2hsZlLz5ZChSiufXX7EW0dqi8SbU01GQ7d22A5UKDFeJB0SO2fxSxZYSDVdJ7
wltyVRSGFA0MSyk1VlLh9mMgjY/2K2KK1Zgl3bSWVWBdnvk7HrhtPGwDnHzuAAZM
aTGrdJO9D7FCtQ6u/V8/2T1o0JtxTxUwy7zzY03NOWqlv81eXLZcl2lAfvj4Tn3j
cEH9HDj7PFDtbS3YYbKU5MzHrc0aYMdz64ZXffod3+Lib35nVTx0igL/ruuHB4ZQ
2RQh73Qk84tMCkwwTLqJ1Knup/g8pTvRdWbLFfZTgAWeWdUJmekSHLTroWZGusUh
Gs6tg4INu49w/TRowTn2V0tJ0f/QlzZ0hZJRiUlzR2iolELKlGFu4ynXFTY7sN3r
YqRSXKV2ppCYC1lcf0UsklkNUOKbSNKBCsYpn3b92zjao0FTnqMu+r1eeEOvdids
5014xNBsuSzcxlvsnXcyi2p2o0qaE7E7n7F2+iDAvVg/LbLPNlQk0qqwgqmbMQ5h
qfFZIiu4arFr6vOaxKvU0pNL5dyAg+BEkd47mT7BjtagnrVu+zLDJo3iWDvqeSTb
G30WlFC8FJXYDdgKsPDK+XDQ3RbJNKB9Qcqv8OZ/P/AsBtl6Z9hTYnd5HK+lcxWF
Vyc/osPsUO756QeOSKtsEcn3zXVk8Zk/n6YjWSWNbAjOsuerP72xDOofNGuOUIf0
SbA1s8f+YkI1wKglFDT6tYAKeuKTAlLWd6bqkcX9Dqn9zcFmX8hA6FDfVbEdsGhw
f2Wzj/6z/zev35JH4oYPx0DDmadBi9i2ZPGWV7CVwG7sW/avadlAdhk+/N8XQhv5
ebydaRMRr/TU+x6CVQCOxmAU+GXKZyR7bTN4zm+UYAhnlcqmH1JwCotaUGFvOYz9
kFNQUjwCQFGwK2j0js848q6ELtdQx+BC3mZpQGohmx6RuFRdiIMjilTKWAuSO48S
unC/WpAO4Z3T3Do64pJTgLtLCOsKDrV+yQ0Lvcjy4gZAHocM5DGq7Eqzt9h+DUc4
Gk3nF5mWpVRe4UD/+E1NS7LtBy9DYsuFDUl0MBaLMFU4gsc0wB2jlF9nNY4H9X2N
j2QF9xw0BhiMVsFYA5PqMuJlo4t5DDGlMgeDbjg13Q2OzRsSS+inbPHpgl49yjmo
t+LteUqi6PN+oJlp3OpoZV5K72LRBekfXssT4SMxqDPffz2nopXLN8y/ocGtbt6n
O0wHjWKDbuHK+ZzJTW9mr0oVqqZnnWS3brLWg71i4y9bDMz0mSJ0Eyk0VnshAQqD
S3XcZv517XVk4ITz8uxrm6Svc0t0gTEfFvzPJP/RFGPre0I6rscs38gvfSATE87j
kV6LmeUm8mf9BdjQRuZG3r4re+yTk5vvLNFHHtf2BupZFSrhOF8tPJ8YXUEen5UV
TRtzDQJ5e4rlhnHqypYGYhlHUAmQTkJxYO6n37EurMcGjUMFdvduoJuFwTqhQlbU
B5iJtaJkXvO4RTYykIvudDDfqF8xzzh7S38WDFf900N4LYaeIvCkJrG20X9lngAt
IILN84aTP81O6TWGDHxjeqriKBI16SOfbcz/sOtBpGFkDx9XMkMuk1fO0CmEkONK
bfWud5xnRudo6vdHxED4xD/0QUoMsUD4rvBrUyCWBRcrSxXCkTjUN3HeL2R2qF0k
OAgF1CZGgeCOuY/UUhX7MkLRRNwYkQMvihc1QFZ2FqSxNNDk7A2D7EuoqGBaALo1
ADplrGLu1vsf+TFzPZOTga+JEc95TGzjPbGhCmeTcov6/CankT9Iu3LeAPM6l7Sx
yQYp6cIkbhswe7p3NtezPQoCgcBRgeYn5HEz08oBRy9QwdtiHSEHQSlBBFnTSWzJ
pnaGwjIdJuTBIiYEhdS7f9IoNniPgKpKGLjMwiQWX4rdIm2r9xCT1aJ5SbdjRmpa
mQdY8xeWiWsYHyuT9ZhWjN7ybchJzkbGjI5sJ/dr68E6lc/xT7Zlieo8Dt8Geue0
padGBNBMWfgc8mXu1yaBBP7C2Byp3rWQ7sV09i3blSWU8Gz/uaPGpz/lRoxWhU67
YzYOzSdgC2B+GNzcjs4vJCB0VX3aSw7EmIxK3v1SEGWXwq87dYCGYt1Vl8N3aLG/
LSsr325tJzp+/4qSKnZb5bFxHQFlLcSpNFQn5/q7ADqS5VFLNJFnugjDjB7S4umq
beu6ZQK/2L2+pQPV97DezWDgbhi3wbHe7l8bmB7ICloq8fSz8RaxIP47VFMuu6zz
UTo5en2S6pF+bF1WVMXlTPGdrzs9GeHaSzJxglpgqVnCP61UXydhdbktadD33WRK
rjFPaEuGLqwx3EsX4QU2ivl6DeV/b/OvY9gq09m4Vtb3PnrBZFvm2sVytvHnX32B
1bRVLTfwA51fCmbTGNwEmn4/N0EWQIVLOYwymQAv2EzPViJAYAiRgipsHSoIw5qH
kqlUNYkwci7e/HUZeY+ndJk2JMqn8UsbrdlrbBb2K2OK+gSD+ik6CAh2hcLYkD/c
gycxOjsrtbUtrqqJwp/mROUhw/fN1CVAvDeGKjAKOuoSNpO3mqT1bGrNh0oANgCu
TO6/feDTrMGXkKq2zjSkMUiPFsdeqnGBCPjW3WsF3pevxs2mXUiandeKzQFZc8xp
99GAqjyia09q0zC0e7a+JCAe8YqgVTGEJqtSsO+qT8YQ0STH9e+67iWjL++gVx0q
SwKgJRg1Wt2myXEk3Uabhx4Sw8V12Swb49RXqD8lxYqir85DsWkiSs1lqyX/sMky
Garja4F3+0U8jJNlzJYfwr4N62CxWYCrS5VwEy/bCRqzbqn5haMe47EwZmSqbmOu
lYArZogRtmyPqDKgQQRkBiPLhzXsjXWcVJt0XqyTMOrDZBS6bq7QR1y62lfhGtKO
vKPxzqOUnJQ+RB6mVAZj1d2K72T7d8/oUcWfOKc463eVcCNYSBekYfL9rpJroNoC
lYOoHhCwX60BhV8YgTzpTWMXQNJaL2zt2/2q9pF3ZazzrzL6S8pfI+OCFTyktHj+
LXyjheWWI8zWubDrrkChSkBrl88DokygyaAgVg1znD8T7YEc+iAhkYsIc+JRaOZH
n55efzRRZX52qTEwJhUom/8mh4BsEUoSDEktcdoL4UrrlgruG+VNNsMalG/oYAdc
dpfPdAnwcbKLPijGU922m7/DEZ64B+JJ3AQiuvVf+26+QohlAI5/kh4ATFj/UH2g
XR4fVhrNily2XuE9XhPdRfN7OKnvuvel6SV0ncaVl4bJvcCnqhwrWvKiK0ksZHnt
oxIfzVSas1rIRYOyVLgzx0lTIrb2MjMvrmSNN/czAFjo+2SaNFhqMGrJ576k0nNq
IP4zAuH3ek6f9WvFVr5GqZPgd0rPCh9ZO+RAdI6irzy9T5ZAXYngachnzqN9Jfuu
SuxZGpsbQC5oQK0VLVnoCGPO1Sl02H2w3N0Bd5juSchTbBR/CxzRt6iLzRZaUKUu
sN5xSKnKu2GL2NdsVTHlh11TAG0WmdnbjvDqCtT54/JXMJFQ9t4m87dvh3TIZE9/
feQlMRo9Am25UBJ8gK5qTdXyf2NBbUdS6YSjv/15i9KxcKDQ3jD0pSSO9I3zL088
Qu3D6ALzR3As5fFk4JSnGkbye39VzIqcqUIKIRin4/ISW9xL66osrknp+Sjm6cnD
cA0Ogsk1R3gOp03sUrh7AJo6jkTbZPNiQVsvU4ZX667jb2AokLu3e+Tdobmpnpme
h7XEJnkSe+V/VcVMs91f/XfQg/X/RilP06x/uWHybdj/72U168nTY3jRGQYLxw2K
BMc0CMIe51eUnUHI4S5krqDbrKrAyyO2kw9q3L419vF/JvEd+cfWUcgW6/T2tfg/
bVK0CU6dWM7bUZsw3/LkBIyn1Vr//mfapFiK36R0xrihAPExm2MxDHFOI8Cdf5WY
LexJMXTlQbC8OLTgB0StcrdaOCytxjOreEUN1IiMzNATJNI2+eWUnsRW8HJhaLVZ
rvViS2ZFYBaKA04c5TlXtGNvQxqZ1jCg9PWMx6DKPgjlE1MZcWRTJkCKVVsiSbUO
sKQU+8ADl5vOxacy7coOr0ccwBlciC/uqM0WT+auxFS72FLAxCOoXuP0UJa15I17
eSOUhIRw3ARKQlKJVT/W0zRR0wmJ0ZxkGTFVGrPCKzyniacfcfUoPKb+/s8o/eus
Ln/c+Zl6jfW4myDQuDnAfXUr/oZgI0cOjoun3EVYp6LcvgHKKkRZLL/k40wBgAO9
e78J1oBwvMMOgCb93NEUl8XUlDdfuM5JzbhxCMgkL3cm8JHLv4dwlTKBGWb7ig5v
Dj9AL3sGmCi+tCFO56sKAkO9Yib7GyzZV8oKy3VWVuiDXS3lKW6n0gI9Kw5mNTHn
vLXLUm+vHb7opttdls7oPL7rHy7zkTFrHFMVJNtYTPESA+pQvodk/CqH+JbmXdp0
8qnbs70qxT0kfeGDEdFWYE/8ROqjq2lnFw1A6TvlRBf2+BxXqswpvtEo0Q1r8Ky/
LU8nAQvUld9ywq3ctzxiaPpyOOA9Rw+ESse6QWcH6T1E7Y7GKIOdMXXeuYp9r7tv
XtO+3IWchQoNsGV5605AjCQ7tlgTq4zqI+BpVbxsTPBCOUlRfuRBTjrGpa5MW3C2
Dbdn7BxJdTZyDlwYbfrqDi02btHVn6l1wthF4nw6xofJ84hnSe6QFdJr3RYX2YVA
lj4ymE/z+H68xkowcMXeq03pROpmPvIFVYHAJ+NJbDpuB1cz+dmcKJTEeea3qd3w
1Wk3oH6kfuHCUVZg8Fq8n7jqOcdFlOQQem0ToL+U2zykLd39LMlHxGaMh4XiedSD
CYYm+FU3OpmxpmgtWhjqjg1NbzcIcXz5FUrvLwou2jf3t4Dy5igO39TXCEjCNBM3
7SicTYAgIZRLCcLJLrfMAb5hX8BhwmulLvbEWRds5Uw2uOUNNkt4g6Korw4d8jUx
LoKREx4QiVpXdytp1H+ng9rncQkdv409a1fo68k3cBlfc4AfZGy3ybcWb+n9GhWa
o/MuUekGDHSaGqPtjSiQkrq8EFtKXSLLBnEGm9uVg1NF7Dp2oADU2HEYZatz/mM6
OWsGe3JGYCvZ9EVJVi5+s7x4UNBrUT0ZiKwewJK1x5tCo3CmmNMZzmDtSdBCB+MT
oNjjVbXJjHP+vPYkYt3wBtNAl8GFJIT+7CV207Us9StWKbUKX8TPmZBHSc52tO5u
HLIYj6grrxFCWupEp8CeF+CxGhXjPV3uPXihBtnPID8LGcrD+L//ILwYGW3oO6Su
e+mnFZOhcrevPbBJkw2p2Qh9E8bN2ZiTE5BFRSY7uIEofbyrBhSte56AIpi1Ztjr
AuhEIsw7yNHSFmXJbsJ8pAQPoEAuvGA5Byu4kLZarNcQESWEq+eJClRz59ktLGyp
DYC3SHAoUYhaXxm3V+OwPTPkzkJ7OYFhSyIyys+vnNGgjmBKnRfqRerpZ5vHSNk2
YGLUzuL78xQEtKL9YQowt8jNSFIf2ReQhrGulU1GeHWHWA0bh1dRhlX5oc4jzowM
2bNbIdv3puskWK35ZifLBa7ek4PtNwfaUlYjSyAK1mTe6Wf03djBn5QnGFwrjDUw
qIZojtoNDD439Xi7pHJbE8czE9VI8OH0HZtKn18SQSdEYVnpNRlVBo/taPUvE0b5
3fw+UKikkVrZygzmkBRmcQ1iRWpHToYGbushg3G/bGVv3tYMxTe0jZcojeQTaA+v
foqZOB3QOQM/zKdj0r/btiO4EkfQZiBMoQvTfb4cvDUo28u8Tj9ztknx1Ku/Z2Gz
J54Z6qKMyKdA35HRcO9Qv57in+Cq7g0QedvZxDs75DOSi8hM33lOqbkEmkXQaiXZ
N9M1ceWeqfsnNY0I2QC2BZYMhI6WQijeEIT/k7x/K00ORWyjDMZB6XIqiJP596EL
lhNXz1/yvHJ+5qGO4fdJ8cZd0dDmqBvkalmp66xCEkDKaVgIwE29W69ySXA0TihE
yNFBbBT353PmSDCYmZjLmvgkPi/Do6fTxs9fOtlc1wlBJLy41lAjwL+qavc56SRG
ZIBwIgpEWz7VxgqqKLMevu5jgb/Xx5W4P1w0dHmF96/u+G3CGShaGrTJHUWAV/iU
bXJPphM6u29FNyyj1N7KIFNsunPZCipfZugaprmGryoH3E2/cpFd1Jzca8DySr5G
arObVq2+NC3TPuaz0mkU59B83EspIRd8wseJqCZs4ATlHc+zLjlSzjKUcl3AtZIh
p3zIK0m376ebOo4l3eW+l9SrTYD2SQDNirfq8/02SYGS/VtN9juGUQRddmla3XHk
0t576okaPV1gvi+avmcUCyXwpEavELzn1Wg/e1hLbjpFy0dxLFTr6QkUrI9hkVwX
GPhZaZoSpig+Z7/B8dzEvB/FiHHZZGOyBGW2aTobFgSwkA4LUDWhNRYkMA1g0v53
3dsyoD+gQbN0XaUfOQR8H65PzjgD+LznjxMgEq3KPpHbtVeToJ7gNj/3Vxkow6+X
PMQzCwV6Zv6srEoJpdA9yg8+qiiUimVLCK0ZxbwHIE45+MHcvoin49+s07iGyjLk
hOkYYF3CB88bVo1QhHWsOIk25/wCdGFih7Bzq7ck5IlArZt2vZ2ChfFXz3ZzxlaC
7tZZfrpA2SaF6h0gostVFMztOiY44uzlX/XVtO8xAww1/tHT4LqW/Mvp2MjuGCYN
aYLGXwIXl+crWKM3Z/+qnI65m3zjAJkpoPYNg5A62OOa8SI7tg2hejY4K0LF0zT3
QsWOgH4y09AnDoqP71r4NEFjOTfrSaED7655zOgvWuj7vW6yO67CzNHcnv5/MTFI
HJa+VcYVhcafaKDqdwkPq6KWDsLDDNwF7DgN7/8MuVo7wovmGzAe8SGv1RWpBYhs
eBkbxw6OF3CRcxVOHqsL8xXm+QBaXrLmcteiCF+R9cA62bD1aHZ1AlG6nnIReI8s
0M7z7YmlrxgR3GKxGtw7dwjIf07Xw9hISoFQN16/jVrclrgevfWPNuI4c4PSgibO
qF4PLQrJZRFXJGaIBsm9pXkMTJPwEM/C0LpDaljZui7G/UUD0e+TWXT6/GwHHpDO
oqo6exeyfofrfM/s41eAITCYhrmpOvLTtT5ezHQrilvV5G9WI2gYSsV9f+GoqpYz
feIRYZnMjgAwXlwm9UOaHF+1s11if3McBAdCNWYho0P5cmPl5h6RgSLXIkFNOEDB
GngIa6e9dLi0FI6ugtr45+l6Iyalw9JS/AGTRmjMfeZYywWKW0ip+dFYM1l4sEh5
ShfO6oYNxS7T4IjQNdQcEjkQyhypQ+pRQYscniDL292ow7Ox8CayO1bWJSCAfLNp
I3S/v+E7Cexa3LZIYwbbyxdP44QbQ72XiLI87mlpUhq8jj/3Kf/sHI/4iBzo12W/
GDQbNbsdaqRl3HZicMVZfqiKgv8SwHiwSxY1KVtQ1TvAFDL9+vD5fWSmuOk390y6
QyPY3M88e2ZW/UlhD/fJlybPxJkEscccMaRLsZNc1a068VptjFOV1x2UeFRJNcf9
WiviYGYtokm/ZhtVYzgwTAeiaKRAEuBkbMI/oGFmRjjjJcO5+o9zlaYMMaPJiUKc
WHDabpCSaB+4RUEl3MsZAkeELTkYvYTT74pYUvDpzqOgcJZnDeYW1TBGbJ6I3mlT
Arp3XlvflEW3SMcZldphBL6EDkYJlT1XL6oXfn2zTrjCbjUuM8rfdaTqW5JoM1yk
nRrSZQvxc5Omvci3VyfouP1QZOItIU9pTbAtdSytDFo8/y4mBDXZF3y5xV3o34t2
ZsGxj7tlp5VE6IeXIN/s422XAa9PwHRnRU+HW7yDly25ij2hT5qVwwDEGjT1Dh4p
4uYxjVAPPVoFbZNaA5YrU/ztxje5QF1wcFmDNNSHDcTk5P8ubXLt2eWMDNlL5FLC
Ezq1ZNimFuUJNqRCD8xTceo2JTHLI+7tDwAEoSw38n0hfm2Bscm1kWrvHOQ0RI7j
e1yF9+8zkXYgFgInE8QVc89v62o6EOvsg+L+PS2KrCemuMmnl2jyeVYPWjNHl4R+
uAPrybPy1dMP7txDeEYvhHcFWiphXxzG89HFpdmOMXlrudOFSYkrIyRlOs1dPaQ8
5zq737ajM3Tu56gcUekDmxARSAf/LnA/D+oopiBs4zxDGqw4HBBrbH1my1VJ/0UC
fyAX/en2+xmWq6tDA3Berjy7gZHJYskk70m8obW210u0qt7lShTmbrBzdxT8FMjA
mTP8wa5FyqWhdP9JCJpRxLyn7nc3IFLc0lOaetyuiGfsiKIeXIqi2nycMse07Tk7
B5vK+bE5OssssFefcoaxDQia0EJPZemMsnCbH7avim9bYpLRvwgB0vh+RoF40Mta
/OY4cvAPS/sr16JtFNECTZso8hM8dtTdDi5XZK/srD/7x+AAGBZBxJcf3m73KrVq
Bywz+S3me8En3uTvrXQpL2ch5uJJkvfE6zXUK8/YrnfbqjzThPpJAR6NiSC9S7Vn
6nXPttaYFMuadkw6j5SjFya3+AEixyyVObZ0imGSAd4jIs0FHCrj6q2VRxRfwhjV
yI1/67gYWjJ5hW6IC+uQKQ8bH4MNCjNF6X8s9fDqNuiTi/L1Bf5GL1s/JNvNhKJ4
TfPXQIrFghPQj1/grsJJrVKJIm3OuwOVtTnd3geBF/gXVE/VTH59wWfgBSmyTsEt
G9881J0L6DeIyQ22JM+MlFldmsRvIKleYXmMfYTnkw2M3YgjuQG1Q4uQffRU+7uS
alfcZeeP1L3pewK5QR2MSc2Dx4IxOJT30jNffIfIzFLVElnjYLq2hRrzKn4N7aQ5
dApuz3QguLGFX7Ea9xD1q4yWzUQPx1f6ZsptFdvR3Y21CeEnCtZ+XuSQw/51i1EK
Rpy/lbX1A93TmvbGoxBoINSyo7FV1DTRYYTJhKYRt7ICwZ7nfei42C9n6HOo3Km7
B1Z9okqUFi/3qK+k/iDDZ+3ltPP8TUOFVcyWGKJiQIjEbCweIMDInS8liaSWIbms
wPsfwSqhM1eX58Q/Tu19GX0Y547Q9wUVeQIEsXz+iXdh+jnW+Bc+GMGYElrJqCuj
ulkZ5gMwvTtOh4CBOvBHO866mzvqmhu3Xu9o5Vsawz1+Q0krOMzNnsuduWeWBRJY
UVVxrgBWJ0DyeV2S4UUFGq25bpRFwrWaeBZYk1WZWJnYs9/1ezJy5rimbVEtKleH
6IhAZbZ41aYoQrrzHDeOmt1l9xpGlBL79gyJd6bgbafOUz5hCdAXP2LqvB6xwzLa
ks4Uh9EeE461Nv0sEk8P8UPrbBI0mZBACk7mO7GzFroJimKZcc3HKh/gj8IZPdWs
odJmJ1D9uPVpnZ/CyNcVkjuRJ+IL9G+HyINsA2wZxQ3cvJt46IOBrlmDqF8gJwIr
aCQ7pB5/S+WPKuJ8chr37+Cvbs2R4VflV+k5yb52nFrXDmrtKxlGbnvTjrycMhqm
64MXQ8uELMMlU60ZKKRMub3CePLupIUHAEPp0yKJcBXTMEOIWJZU5OIIVYWiiJKW
pq1li5YqbJL8Gf8UQnxV7xnG1hJiiPIuxgGxGO03YxQEw72ES1l2FDmBOuTR2R+i
8pDdGZqAppPlml8DkZCEIvLnUvWseXBTqiSsWmeKMnNOWaoPnOMJMgqW0TqX9psh
xXcY7YHWf/0KAqhXKEebZd8uw+dYVK81W77APAGhhPdl8RX6z75zSiyYWrn6eAKG
RLqdMYOs+MnkJxhqvFh7vGq1ogAuW7Pxem/13mqvdstXOAsWxsltxxrsyjWhwe85
t8Xq99C0yPAi//MTNsnYIj48KtCHkNkbWZHjKcpU0ymAgioWNWPpf8DRSm0n4GOn
btDN2BGUJxhXHFVQpC81zxwG72caAxbY9u1uPCe/LPowHx6YxqBlrR8hUWsQnvaL
QM3cmiVJNlfr1Dp9wiyRENMUetGc+97e9+PWrZC7duTYqN46cBlB2+VdNPVCmBwD
GyX4l4CWu9DViuYq6pFuLRM12gBPYNv3bhETFLKysyCAalozL2ArfovKs4eYo2NG
zWTTU9ABMwbuS8m/Oro+6ByeU12Jx0oXafBBYlYtYWVGrUgx8IwFr4bjB8w1UtPo
I7t3MRctMhxiOGFDuR9VYETUY15XAu3njv8fCOlKwsNduDqOtZ9XhuaZf6xGzZF3
7vvX18OVOV3YuHWwD2Jr1L514FtSF10/V/Oqo4nKTMXRN417jwFWVu3rVRQqSiWQ
B7Kc0E+KxUo3yb16iaS0gYWliwsxQ06JKxQvAH/wP6yVZeFeR+J5SYN1ZrO+Wyfh
t0jOljSaZ/xc04cfZCVIhYmVsN8qEGuKwog+pZ2ALiaLGIV/+j6oJW7oCDn81jz9
6vvH2cL4QO3lEIdc4qpga2ArRWXXlXGXRSqG3ZrjS/HRhpRzUHwEnZXlgGxIIPrA
+Kd3ijwBLPCYnXgQ0BX2+cQ9disMPjVCqZoZGIVCj4Gr43/8KpgJkOl+2+l8d50g
wxphGNv6/VJvGBcgd8CRSEcjOHuD7BUMJC6pKTO8ZNXkkjUjAvVN+xjfEO5Ww+h+
CULQK0kQKqXhw05GHHNl/Qegyxr3hZJMSOAN7xJdKlK4rtaOAcKwNjJt0l+f3ljv
JfKiUH1oPUrIpVgubYtuLnUwT61M/IBpxIkeMj0VA7j0ws/6dRMkTmQD4ng2EF0c
+SS/uL1fEo1Wdpcfl1fEGXpjI4uqluEihhljwdqcudDX4XGd8v9gKOT11wqFhgHs
sj01y7HE6K7nGG+poUlmxhAKcRuGKxzjDxbSIrOEjNwd8/KwmTqP/qUZv2TG3lyZ
uH4g4DQYtfBR2xtsh6pJuVmVOy0p4Qy4vWdREMYZqNY5e774+aT+dKmuExSEI1ld
pqft8rI/FSj+JgquT7YqgGi94dMXhtVRFEMM+wsFcFJy7DeuLmCJP+agtUzlqvHT
R3P7pDYtQ7QgCNyFvPneO/t0xhBfattdmcmGi372BMkJ7rBUlUlSX3dXA4qYzRQM
yAKfSIDCwPEx49SJwZHK/DaeHmFTndiRY5SUybrAouUuBQXauIYt/5EhlLgwYsgs
LHgf4UOBk7i6IAK7blZi1m+iLrdb+HBD8AidQFe2hlFN8G95owEdmDDHF2k6ij/1
jEo9XG4uoTTsauJGujsuB9IdeOjZLLDFYy6GsmJOLiFy3A2Ee2UKzn6Yz9sGJTVs
7Okb7Oi60iV1e/FO/1AzOGtXX0zSWIJydvQfkLTtoH++mx1Mh4ttopIY11hhsNi8
xwOlpDtOAkGPsM+MFXFIR36Bfo07Ild44wYBkIZjFCr9UnBsuIMajuD6moWM2DmB
4YLJlFUvIEgeHLpzadvTTOKajnfTRfxi8bpA8wPIjT3yFuqV/KQxVeVwK/22jYEF
ZRGgYcdrxZao0lgd/iC3WNn2Pzdq8P1MSzCf+d+yoL63QCBySfNWFQU8COZgTyoe
UOr24dGEk7OhwDWzqHyK2Fo7FUA5Tqmj6caaIdWQ2+FRrGgK4SUIdkMfpv4eEPaW
Tu1hU4q41OQbbX5PGfZfCDaJrXdLBbrUHMsMbd/rr5vlT24osrokRuH9xSBh+p1E
DNbCBmtqIG6fze0NyY5eeH1YLz9R5/la7sATogsmEAUrqX5Guv+dNnq43zZ/6aH5
zPkKxbIVe7Db3jvDwV2aAtoyQHbTgqRbY2PvXfV46ISbqi1MX0y7OboYbm80npYJ
UlVo3atEq9Hs4DEWTBehHbFncAHUiNC6747I7wat993njWqcg7YNKmUN+7fX7iyo
InEDq+cRV1ohoSdJqpPkDGwva64hXJ5qZGd/j1AKHO0bkS7cfZk5OHSEEfDBLC9q
rlKiLljkcmSPaeobVhi149ulKGWCv9VQIJfpT8wmXvNui903RIGnJA2QlTQ+ilAN
9WjoHyyTZg+FHpGoSzkGzHIvyTyBCfzqm0ea0+Bi/fX/92QDdoUG9NRT0pxF4OXC
sC51To1FWYphH2b5StY0rS0jJZIrA6o/mjsFsuzes51chDQWQt8EKNvLARXHFd1c
YoUgN9MJA0j4PjW6Y/goJGjbc9NjIFf9BpSmd3S5ZDk5VSMnoE+b+pTUJkKoKxh8
Cjts0Mfj4dAjJCUSxUpZ+d51TMo/brODRPWeeRfvz/NfP+7kl4Hq8QurWBRkZtXB
ughGCM30kQ7yivTiuVQKgzIvH1uEb4V9kp/H4Ostd3BYgnWFyz7OdNx7JS6qBmY9
rymuBPRBXuOwz1tgjSYcWhF915qwy0gGnrVU36KfQrwymNn+B2XNe8V2NxHJjFk+
l9fvXj9LsFkoh8l6pe0Tk4fLr8fnhzV/qrLEwH7GdrISkm7ieCyH3fziJ/F1j782
aO4O6jIuEc1lmt07ya7Qn4uAXgIUZcUIN5UFmoHO5731773ojFOCd/SK3YIpHhvE
ufuQ0tJHFPHDFx9/PQ/UmdqcPNPLy9rx1IE7UB4zaYiFUAoX4Sc4+gF3ZJ5utOgz
xIOgYkgiZB9SsjlUgPWCKGGMebueJwzTFt/Ijts5hzJkDLp+rzFBBM3D7vDtirR3
zfKRZCgY0Felgu15/Rtmq9aBEfDlG+TJ8xHsexx0QW6wnJ5n95DWZENJxi1JpF5W
c6BKtTmS7d8X/h71sjL1vu30zPYMQ8h12emRoktCmFgxxMHZ7KXaC6wT4qfy8MaY
gmbSDgZLkCm7peMhc7ZUx4qzijQwgms6+bJEtZdrgcs7r9nppha6OmzEPkfH4AbX
q5QrlDPS22+tnRhA7KvgDKhr1HZuOVKmV1oi1IYECkUxwqZBBovHuuvGQfJ3g0eO
xbkEsQDr6ELEq2S8DsaY+62LHF4osW7vZT8LEca/zFU+t9cyqrzNfCGP5leKcpyc
tujBEOCKVkRkNR2UFEbDZsJbi8dz0fZQpOmTFifUidHg5CxC/0cUFbXNQAOHNH1t
MUs7ReiSjqmTVBscqfUpGtd/5ruqkNNdi/ivDc7EfRNJUJJhQkq4C3BtzbVnm4bX
DpqkdcZfPNuB8eirDmqO39O1UnCZ0LSXZG7SBaKtzuf7lSe6JzX0phbwRCBswWTD
YZi6icJvwrsFyYkTp9c3uiohTp96yVsuNWp/3ziiHGYfTlj8aZx/gxDNDZSpPGIk
VFzc+WU7BWsn6OHT+YU4hn2W73oY2HVomydF7/VDVujUNvuxZzPN+m+xbDb3/UOK
SM3D/QO0zwNX1n7f0HmuhXVMVmW935jfptRijj14UQ3RAGIAhOk2TrYFq1JOdTCG
cdqW3H4us7L8n+IBb37gl/7FfW9G+B3zTg/o3po0f4kbO4RbUiG0M7WmbehOXt+H
0Gvbl++UQSfFGe4/glSnFsjQijuSqbGQwrevkDx2KLxQm1SNjNjSegbFi1vl/sr+
k1bTR7nB6Woy+z+CFMLBgIYXDUWhKIOKdT0b/4t6nzG1+bBhbHm7u2IxdDvvDPYq
Ms7XGdO6tPJgqZG2OmOrhIz5nm82qSRt81L8oWwt+HQGq0J+W4etid2hgfUF7fKX
1uhuNo0HTsTt8hctnzjn0kXXNBEYOZHRhbIez4FK1mWYasfrvCWuUnMLnmpx8KgP
SJvD0L18jwmug4Z/9EF2klt1mrJlik3i4Ikp7y7lKYoTcMQ+Vak++nFPG51ce+QP
nCDRTpyWGR1ULeFIiF4lkUmVFTG3QbMREjWH9/6hIMaphoBjoctsWO2DdzNeweIp
Za99igK+HttjEdGRhzN0JvtIYXaorarwIJvGlu0A/0RPUTmCc31tyH83w84iEsrJ
Z9RM+I+9Bvo74QDBz0qgAcNQPhYOswB8IY6IE7RSN7R6hO8hXe6eNLcNSNlnRyBj
58EYAtsdXZVKstGX9VBHnvmu4mc3NLPBC56opsfYRRXtKB+RBaRqc18XtaK/ZUbs
Vnqab71S88q8MGHWOa53wUgMxhBBwIy33STvwA1jfDNylQgZfHPloiJUOJtSYdXW
KxBWR+JTMJCQsAUteu9NDZFZcsId5ruQxZettvW7o3ib3dqf1Nqb+A3KoKvRnHG/
Gkk/kXjVZomRm4sdLJUhHPn/i3/DdNqMyxnKzzEfYcz3rPSHFm6gVYTKfGjK06vW
YQnlptOoRfDgsaIPyqLdaFtNxyxtwVj73trRrEquTt+nEaEFuAW2XSvaWVq6jJ7S
gcCJpSBrA7QD6qE0t9X0PfYypSeiPqYHoFz8SQkdNn9cJlDSi7yUmUa275Erd+kw
7hqvd6sKd/KMpdbzsBmKpSo8KJZz+7cUUPq6w5DPDu2yhS5SKGwGQx+ODZv6JDVm
TOFUXPMv51iJxJnUX0JiW9QLXL3akTe6dj+aCSgM9hu4htOIlILLn3esDJUQ95fp
u7xC+TkvjgjA8G/aAlvPy1qEHjbWJ8u5Pg+LBVco58RcGUndoXqt/sIMf905wMsR
lDUo86oIiBVnMVbfheQy2roiseQt4xrzNaWsdfJvwrW5ol4QSkvno9IJVuM+3rVa
JmKhT1k4Y4UxF1QG7imdEEakGepbEozZzJSn6fN1hqpub/YDnhkeM99jWtyWFFrt
QdiTyCysbqLaLvGD1LYKbcdI37uT+/QFGZS6NL0gcCaRAnwfi9Ul2SSOg4n6uWMB
OyU1HXzod4ICvKz8pNWtbCwW/2tX1ckAeyTL/SjuHjJGrHZzBYyryLtqmy2Mv7+0
PRa/svUU1wzrlEkDHJiecF3t330TZCMMQ88RLMfQxyJM7WYLyk8PSqNiBTIC6T41
Jj7S3pR23Y3OmTQgdOp5PKoD9vuYve1qtkDetNrXaJ4pZUZU+xw5kz0l6fOKUpox
wmZo9Rc8h3FnRtsoAL6KonmUsZF8TIu+DJchbcR8QCLyqM7kmhrAOBeMmvl4dHvk
Ga1vqiTpJt/rHTM8jQF+3NmvObbxk0/YpoQWSkhBl/ByOMVMLw2vl7/XUho00fFi
OWbodNOatV9D6MqmjzaVcHq9d9QyoUd6u6F4YyyoabTh02oeiuQYw+IQwcKAtv9/
trXBHLXT4BIazk4ZhYReJXoawuO5Jt7B9SDS10kyH7PBRjrSp9WDhhHLv3jjCmAM
ZHub4591YsUQ/VONXWr6GIdAaEbB9+P+sND6b71XD/JjD/D4bvfmSN7PXEwvzgXx
/uHmzQMtZGvu5G0Bg4DWW3aPa3LIOXBfxOZCd9Zb+/lSF1rFXIbbq80+vLY6OJXV
JFUvXXU2w2yYSqITPkKGp03qyGZR9jUe+ti1HHEz8QaVwC9g6mQ+29AI4NVgiQBG
5R/AwDZ8x+P9PR96+39bHnwGwLNLP2RcWACDTCWDOl4gxt5Z0x7I2ass8Q7e0dmV
sFFp+ydgM2Hpw0hQ2Cn+JBk++UqzkFCd330pxvoVVkljYSWKSxUrpfdz6f+wVhDo
4rRs49QKGc/wcuc0eEZp0AYOfOOEY1t1I8DHijx3iebd6oHp59X4A1SCRmxxKGY7
w7uMyupC3WOk6Yqx9eHOEW/iqyI418SoS/0tYMjgzg6phk1zpw0sxm916bhnRdKI
B+svnlOVjzVM/ehJ+jsNcL+yG5FuOSqNbqGTTkNbyL+BLSv4g3afnl+4FsUANVus
H9yMU0yQWDTjUnxjPhmz3y7hNXv2Lng/49y4BQ1P42UR5/5AassRgOugxUrlMwr7
o+TUQSmvCX3k+xBfGoZhMygWCOQdOfxE5MnBL6PTq8qbT4Y98QS3DHW0uM5Zv1LA
ulUy0R1r9HiVVXjJY1vqFtAC9RQoTy67ZBHqooQ3/9mRrNb/26vk1Yji3pQFuTa+
pn1gs/q6e4+YwRnPa5PCZd1PEe4pw7BvRGCTa3vN4LGXYbvVrLUlNZrWdJeuQk3o
LvQ0hvN08+R5o1zPFsERqUWJrfNsSbsoa1nOEcTBhGr9NdK3Gglh0u/jRubMbuv/
HDXLm+2IAqqNLZU+LcO5JC++nKMjUJYdZTQm1BMAk6nLa362ra/B9IQKsfdnAQd+
jFdsc68sUgTns2ltGGPatO7OxiMZ2Qf3PanNreCmH9lgM+6yymgdLuewnoeMWgeA
PUpm2mAcQcYRQnLFdkOdZi7mkympbxe+tw56q+xRkpfYAIJAcB76JQ3l05yaI7LX
ECaoCEBNali3+avNtz1Fot62Rwf03mf5xjQRAYXzI1Q7GBqSdGAiE7emkR1djWBr
SNbp9N5emT6SymmH/TVwLN3R6/IuPT7eE0zw2D5YT1Swr+q1GZDiPbRKSyxAajfK
GT8yMRl6knXdZamdaMEKVem9f/Vk7c5S3+HiZGZdPBYtmdW4fo4cNDqn2GVCUz+X
q+q7i+P4sgbrN/nDNu44HXIChFNpY6UNpdRArROrEmrippwRm2V1W7PV6fVaya8m
GlamvEMJ/bMm6FKLPDcAYm3TyKlvzImnD7xRMxXviaiXdez0zC6BX3UJrbcSi6Md
ViV0q5JhbJdeyOWtYl3zpYRgfaxin6dl5S0wqw7gncT/E4hIdcL+wwJY/+x08ONr
8KQ8DWOd+hFA8V2wq5QRnHupFVg6ZggpXHuvDrPA13Lo6ObSlTfv2qW1wD5+vZK0
cJdmxRIvKzpXuAxWYjYOBs6A4jq4HJ9+blgFqZj214NbAv+W+uyeSQlf2WLkmOlw
PprtB6yJaMMmUi6HQokFiCHwfrTnMMk7toATMblhhZa6fRFQJ1yiD4+uIip6tYCe
eHonMUUCwK2ujq1OfElTYPuFM6/3D63StcOGHEyyLke0cQRCb54pBgczpVvmT8rq
+JVpZrYtEp8L1ldrqIteSt4WoNpfrEdyk37nzfBBurZilzQItEKnbPQUYMNKvsX3
JUF/lSMMnwTMMquZJZLaeAO2D6cDZzUwQzYahDIGLbRe5h2+eQkOY6z2EaOUspF0
kIJWCMwLHZ2OWJ2jruElLoU7gQPTCZN/6nZ42t6Hd9vKyPVeFmctrEIxztjYQYTe
g4hGruRiS3R6bBnwWmu40ZTJ0PYvnPVJuiw9Ldz+tmvwTt1jfVmM4UdCrtWVHK3B
et0vcHAJM9Zvt+eJIF3Wpc84QtOe4BE0f91Lu69n8OFR9Q3aj1L4JIN9B0+Y9l7D
ev/feAZR0wNHxCf1IltVwfyzd8yMRuRUCfVtGXy9W4TdagEX+6FWkrfpDqhPjVtp
JoGJUl7xwdwTQcXOvRlekLjTc+pC/PHt8mt0hnqZv3Du31fgnBF2w/I6+edcpOme
9sqvMeYCFoXlLTuo52yv38QkTygtmPj+iO8Q0hwLAeT9PxPj+1XV62FK0Mg+D8A5
+yiRNTJ3ic55Vd+J3ifERfrUXj/TE6GfqpR/b2Ip8e4Gv2VIv6gNE9Wu7po7OFvn
Cf0aWHv56EQzPfWWZVRXQsMgu6HBb5Vc43IQSnCEg34qrojlnnNUgpoOI9mRAXt3
mED3T8w6xdOFtwFnaTx1mw9gX0PoYI2l9udTAQat6msWFiWuloQsB1HL8uuqK0iV
c+4UVzin62uVNREKxoT1FVjBpSTY5sOoa32912FxcUikDfVvKdWnxtMVQeM48Z7T
VTGTnAxYcZ2iCFMbUsXw2VvEskkiR7vKtU7U1jpH52N4W8i4qH9hWbRDUFfifIFR
AZBCx3/4l/oQaNA9uPPGi3WnEDcRnsY3GG7wU+YKtc7bSoYssjsduIzEXtqQw7We
+qwQR9W6wDeNb0bcx0lKeOY7uN/xYwPENpBrncaUL3h7qweDnCJXjYy2KLiZ2USg
pd4/pp8683/kAfA49Qe202p4FmVgr/LBdsxEdEubPCL5aY+MVk/tLNMpUpQZ8kHs
ee2IF9ovxIrJvLYhY0dSWY7UF8jkH17F33MLX++fHRZ3aP7N4atWeFzFBdwjYdp0
cCNl4QhWdgAZbQXtQiCJUDcbiIBKsYiQnBScmjdmKGcchLEQeSKaHkWuNInFxD66
fdZY6+XnBXCyHLR2TeEWX2ilc0hsmuqyNQImpCMVt4lcVdwlIbp/A7dgQNsvA3SG
4QTeEGUVIfYqGw8zTZmNkWFRWW/l1pHAI/jD1KVZAsre+7kWEzctgSFajA93xCyL
rGWeuxsX7FyoMcju1VgKVmoTPnoE2g05jbiNUjyNA28TGgviIqK8lvvImRJjq00X
OI4S4SIRrRkXNOQKbMffIu2YlIctIhJVykdR8t5oF1yGAFtEo1hpjURWHqeBm/0u
50uF2Y6MaeNne1KGcbhIPxhWEL6s15RJAVbDz/IfsHqziHoZ+aqlcBREwhP3Y+oZ
7g4c3XMpp2O68Ei6ax37g7/vRhxXQ+JB+wfuk0LtrDJO1V1HELpxFYNVdOluaMma
yjvV9klgQXMldCYtvaIBJM4HCkeP/hhayA/X76b/PvYp6/04Tay4QSpJ0um+erkl
16XYlc0j5lDHyypT4hgmKrV7AI0n2LT+M2bxX/NGNj/XY/z9Ktv1HlCVrrMoxus4
rXTWrfgw3Rmg6j8dek9Y7aDJZzJNZ2X2R1nuyK0VqEh9LgolGfuk73PbhQybuKFP
wb/Q1CuwpbkUVTmJJ7Dck++m6i/ZJQIZCJDjx7SfHa8QBBuUoMHC0Oe8HrHTk8JY
/tSvWWZdJtmuHnj3axmBeklUDcsq/28mttVGspFJcWyCxNsRHPMATwCQI8e/DWEd
XipXb0oZrTcIihwAvxnHRPDR7IkmDglrO+8ly24Cv1MygOo0Jg6kxmubhVlDSE7Q
wr74diyniHujHEc1uWc2zRx1EZ+aEK1f6aPeH0ys3trnTMAh+KL5WHrmw4Eh/reC
owFEVocsQa0zf+JfTyKuyCZ596OBbRGL3+3oADPTqs2eKgLGEKqIcJrl9zYzPEOl
CqWBv3KxjsxEKmKIv/SpDG+CCp0eSgidpHtqqplW8ekZJFqSE/z4Me+i2A0aJHd2
HuddIPreB3Wo0jEaBZkIDgVszqSpr3cU8scrCRuVqzuki7lZ09Nt60njOyYxZgFK
VMPC2cMDGzKQLUv01u+QtWC6nsDlZsUJYhCQVPr8fonEY5XKnIR9vN+sqO4f6sdH
znm2q2V8HJ3RS6LhpFV6eFoeZB+vGTrHEz9rngK/Js4iMm1rmDeZYcHAjRiRgkUq
TfWcKKVxBAJdtGLjfGF2yFZIIXt5qH8OLCObM9ZYaB0KP1nxpGZyzuIYN7hx+qv9
w0d59Hvoek282eWdbhPpMSW3udO++M0p8EvcubMtmQSjxb1l6EGB8Q8YwJKcF9s2
I7zVfwF26hdWh0iZsjIUI3oLe/JA1zQF962zWaDFUEd4GkPLq4ockFbNrutal9SS
OoC2hUe30oTV4hgBuZl/37Izmvn+MOxDyCEPVHourTLRm3+PAFNcQ8w+ctZbQc7p
xrzvN/oVBGu4jUOnK3zexrx+8ax+KwZ3Ok7Yru8Gv/yD8c/wQlj88dhw/j1o5xv4
Yp3UOrNG7fiHTjeIg2OoUOOJGGoRh3ek3p1lF5fxFDyOm5+Kp+N5ZdE//Jo1Zuhy
tz7P+yyl+OYe3sOGUHyTkhN4BUnoaHepcPBp6qRFLMRh96CNhy9falDuFQIAklN9
He6uNhhH/xV2CXgoak17Y3CUXDZ1zypFUHtFN/GfhMZrAg6VAJcGxLg5uNLfYIei
Vi4YsKqG4bac5XVIjh714CT5djb6keJhY9/yoPEmwRzOsEsWxoczlmZPK6A5+fdK
Vs4hGh10URIrjfLA9LvJYggdsx3SrTSMffQF1xlxvmgqKl07ugFPW9HERHMu7VZ5
C+98qn3Wg8sns22BlEAJLMqF9Yt90JOh2N/LH+mSLKUtiIebe/NxA7ja+/k7hTTw
dmoCriMY0vLEaPhD+4RtTIEnVUHFZ60Nh2FrKh+GNm5PCrX3n5w7i+u0bmfUumwH
Rm5Ug69mR0Q+7SeY7lGbcO3ESRnqV0paiUMWnu/9G1FXnYF3538pkfZR93v4ay7N
V60SFUDHkSyIjjqALDwOnZAVjFtmKrAJbQDOZTfdF7R+QUmcrLAc1kyUwY3KXbGl
Wa2Ntn5VX+WF2Zo5ubZxA3v+s6rRAB+zDyoAJ0O2v1RokSF/OxdKhNb5oXYKMOkc
g5GoLOOPXG/bFc6Bt1BzTKAKJNmGJ3JiNcHKSzKk1kf9a94zphM0xLl4HyiLFurq
DEu6MJTs3e3mmGIymzgBhh14fuM11vTUxZF3mnvNybfgDUSiidWP8sfVdsz2jFl2
vcQ/LeDLY6YAMDj6PQfe51dFZAB++iMIgZav0JmvTk6ClssNxNE18dnwul3Qo1y/
TM6BUYziQRcXhn1bAq9rksCYO4SPUeDPZwfNG/uIK4agvUxcM/a5AKOg2j0DTUO/
CihU2qzNY/Nh3Tj6A++U4GSEU2w5ASXVJVt9i1t71U/EFHz3rsZxW+7i/33FEE2I
UNh1r60XTxz6J0MdxcPYcdzg/dnG1APXTnae/rsHmjELljQTieQHjhGtvQ70lqAi
tBCiGZj4Rc0UFx4A27+pA96ha5FatbsILmTp8FT+GgUcfd/shsFa0zZx2qJnDzSi
squ+fUl8oryTQQJv85G45Yl2402tCpWKKMcr0LoP/cjd+GtbElibjL1PVtQiSiAc
A5SZ17FzjvohCqWi1qp6kVJ6YTpY/Rfg4wPiNpv86ZJkT6TsgogV8j3sjLfw+HeH
LeKoN5G76OwZOz4vaVJA4vW9AxHulKonFgpKRRXxx6D/Gu75IZVG3LRB/TA+2zQP
L5Hrtb3pwBnYijpo/mRZNKKcmR/Y6+QbixC7YIy+VzBJMgGy0jadDJ7Zb/dfg5Dc
u9czVrVfxMPwxfL3wuA5JzR0BtJrGr8a7ZIrxIbUefHCDG5o1hle0fQ/EDe/ZoDa
j/O25t7ES7++he0/KZITkguYaBFVFzAgQ+DF1QmZ0hnoxeaeWu2xAnhtMdGzGo1N
AITLpTot5b5bB/3mYEaZOIPEj4rNPIAK9AVwPoxx4+EZF18st2bxhTrDOrgyHYne
qxABV55OaT8T5j82OZlsSsMguuwfENHdy8kjrUD5q47FxFikfDlsbGD0pQ+ZK2WE
f6sR6PRQtRYvQaRBVr9by18uuui/X3UoODDWMOjghp+/8ilCJMsD3Bx7AWmTrBA9
3Xne4g8PF4wl79vB+OXun40nN3TETuScKtVqfKTnso+6C1cj4PSM6c0k3lZ6TrAM
4X53bR9CNVkcEv/xe/aMX1AItw9j3US1u31VcOnrVtr9f0krKRlNOsYNZOiyljTw
BLUBwB6gvTcKAN8SmgW1A2OOJSOjl772pqr4WQUm+kwksFfbJlfJJsVLtmxvUtRg
DTTTwmGGZUm9menoHDyGe5C1VxhnG3GyX+rV749qzaRiJV1JIypp/T1VjlAtwakh
Q7pgXgbgUuUI9a10ZaA3mtwhfwH/Xz2MD4EQz0RiiP3jIXcUKlBSAf4H37MZkL3r
kygLCv9vKfMtJWKhUG+kIi3FLwX6kpcRb1qQxZo/i2oQlAGgD9cnun2bL1iF7hh7
VwdeChpIS9dJhqL0dKVVHhFdR/VMe/ipMUmitsJWadOB3QCC/3qkkz3jjaWQU48c
weSGVDo/dy2b7rdRQiceXBB8kTKyGwAmjnWLrDuw1FBcsBHYO65rZS755svqTsFk
eEhKC95jO0SLZFn9jeU4BSav/3Iv4PwRG7fLVVjHWptf+hjfsF23rSOOgHvMjWSa
9Jvt6kPMjjyZDr3BDOELRKP2HuPPV91S2pH0ayASh3CfyNvOSI3iSJhddsPKT8Ez
6Q3UPvz0jkhaZnR3uT3pZx6t7inC/LaiSr3FsdPbB3NtXzy8zmtLcuYRuT5oMW+C
z3KHCYXa0sBHWlNnkYUXfTtIbEepfuaXCD+KwL1nt/Eohe0O9vpj9ok2H6+mV3VS
fk0CPXNcNXt1GmEhmmVxdfh2LN0SnNDX3c62KQpRA02Xcl7dmVAm0CohJvjhYEkU
qbmrdXHtOR6IYOlMufS1JBBfZGg0TKFIkk0wKKI8BiZl9mplDFs26T47wnSZHvxd
VJIaziCZTdgOBQuEkcM9NocxuqbUjn4iU/0lNi0DRxOIvKrDxXUx31Xvz/JL0Qv1
oUnAG2BrgrkzI+uPIMlWlPRU423Ajoy0QgGr0aoRHY6CYYZMdEqZFlo3WNY9Ylnp
T1wmE9P24AkiiiL4GW/v1qXhuUubNQ6m1vqKP/s5Llsy9mV/bjH3Q//qWn3pVery
kKWEUPwrmJy0UA1q4JL4jkNTsx/C/PeND3M4P31a3nV5LrtBCW2w7qQjbqSnXOCt
eRVb2uLW0X7SkZ7ILdG0w59zLd4agHHL9zZEx340PBYI87NXN++BPJ9Va46gi7Ig
XRikclTjLWY9bUr9NcaqA/sXhJNJEiS22Maux/1fePgoO7aS/xDYbxj39B2MQnzQ
2Yuck2HMbmGTyNI6sczyO8IGr+Ig94a9sy2lq4ds/+z3mcZhOlmTH+ymiL2s1bz4
oYTDIgf4R3Xu013einI7boWxHBcwOTZA78+YGmJWBiWSl68tLGZahnKUcip8MVm3
+627xCxTh73MCCYLlxbMP3RRCpsrAKibezLDIwthyNWrWEDSpAWUThvL2NXDSon2
zzfzr3h4VlJPTU+H0s+4rRtH1jOSanQJ0RVOZXAuewBvJQtG+EsPBMGI7lVE6Ayl
+zyETCReCTmo5wGVjs+iErNQJU6YYc+D7zfETD42CaTyi7yE5xFJycAZ11awrc7q
a90WSnlbOD+RvnsFzawR3cnki1d9AISHjmtTnXw3/JTbK5W3lE9RWR11N0pIbFeG
ZHlGXaiUTO+3MX9I6BkbG8PhnEASzDygAABa4N920J2Fh6OgLyLHKLyCZcxRjWwa
QGdZkoICKTBXD5Zm67EPzNCkFxqg6OfhLxcYkTkZfpr9vbifmWrgcoyaXJROmVrn
g2Dx67zMhj6Apftzvx/z5ijb1pAAL36M+XvE6rd0n299KuKHsvhTO4mYXe8ep8py
V2XjxfgRmVsstJVCpjGzl04h7+UGMOEWAMN+/mrA9N/1tEQ6XRPpnONy08BRzsBC
i+14tvBNMgz9VWLRVSkWcCdU/ogcB26qvoWlaiTKBMMuHBao0co3Xo8bTf7sBf03
U/Y2aqxkWJ2yxWeNGOnbO1sz6ZExhQdUysu4NBQaLvTOIcN9zb6lPfF9hsRtgTtV
rpIE5RnpHT6Mno8A6hTkIR253VEnUjHlFyUVpLgmkRq+EbTQ2u3oKl8sXVmPxoTS
GbXqWSwdL+AkTT+0zeRvQQ7C5YWr3oCHCPglCIU1DbyD90TCawRFZdisvmdWtnI8
x808oHMYGs7YgBPtnAnX4atxajKZsSM3Wjv2YlORe616IFEVipGj7sQfV96ZnkhJ
5ZS9a41WouJDv8bt03Zc7PixatWFbyo4MrKHLSg+AmiJBnhUCBXAzZl8zbsIr4Eb
so8JaXD4rtg5ow6v+UDBHZP6go0SsLVZ795hqgVfnNI7AlcNzY8EycDidfP0YnwZ
/djHJcwj1pUSjyxspNXi8mKtC2X0IX5tFNyrLWe1yYG+r2v19UpUG8fNlfeAVoxe
oXo/RTDcQZAvz9zwkutxiItFz0fo5xNyiRDoCHUVKm1z5i5w1eD/j6yxhj2xAlYq
G4Ri/u6Tp3Foxm/r/Lv6ISFEn/oDbmy3YFcv19f/7mpZh+D6dweaZ2pHFaNXfKoB
a0vFTbvPA4aue3eT3yza9qQlZlHbPjg/dxShlC2IfJgUcAFUhVUOxBKySDyqmKeC
rJcuUU5MPXWB3AENYAm+MPbT80/shpO3ORqjzFBQMlKnBIIsRThn2QM+NfwKC6AA
qn8lOQnLC2Oqo0p9JGDL+BMiQMg5C1WAjVnqOxjGsZJug5Y2BNZMv+pTUZ/PJXCs
SXSYfBlja8Z5MPiOolzQJ1WI+nVRI0REOaMLvYLZRT/FS1JNz0DGMkYyjiA1DX3N
XLzdHGoSar2+ch4fn357XE01bxK7u4TonluJt7heZXMGFNHJaUFMwPluW8E9EU+Q
nqoEmFMZzaOd624PQShg59Q9c4Q5TLx6HETml5NESUDX1ymmrDMJmxx4edlFYQtM
ilNyuoLC3m7ikKLVg025klOMSOkvO2Ym+AU1hF5npnD4yfTwn0Er781asreoilLK
cWpl671GiAvBK5SiyYxOA0+xU2FuMv3BL3hHppLwzZWdWpYEQagb+1oSgf+2Vr5H
Um7CMU3dsYUT30FyvY8lBEkZHHh+DQEUBvNwetCE2VLixx0GGoSx0s4tTuYHibHp
GocEQMAvQl8KPhMTRyavU5J2p8k4gqKFycvS56Svq/hvN4a4KLVlI3G2YDV4F3/Z
ireoMfg8sOaeQkbQLRvH0UHRTab5aafhp4N7LmRznvwx2fmPpdqub/tQa9CRc3oY
bYz7hBFQ5ZV+a2ZIgRTZducCrzuDf+Gr62t6A7Vwz2Ul2fIrkG423upEZHAwMre/
rGHP8i7kdB1AwDXZJ3YSDOTJHY7zus8HoKTD/+yecP1i7pdD/9TeTxWGoFvGZDa7
0SqwEc4jYWaR/LMSSV8ptumlwg9TfDdK4mH6xluC88HRnSavq1YCTYnJUfbgwV/6
FTzpJ2K7i0e+MoPgNuxXYqlIEpRucJ/gdMNuaPzxTXeTAd7IWyC41ytRdwz0zHgP
j6jrfAaiEUPPPR5IU7oy5uepxZrni7CIbMV/zwS20mNKyomEkF0c1c7WC/wbGmdg
OZGhemiJIo8E3n1mXrf/kU8EPyy+2zchT13XPls/hRU8GIjSw7aBrFZMz7g4aZt9
PtEO0y6kg3n4s6RPwZnunl+LY2Qw1Pa/JynMmlpAMBl+tl149K54vmMzlZ6wahwM
jg4mBQlmIAS9fGxumJTSFmb+X1HxgYsi2qSiY8yf2FF/6vwf5cYKpgNWh3MdLeI3
EagRDj4/xUw/0I71PKJsqpI+clMZat5rOmKTZvBtDgL++RwauMY0efVISr5vfC0w
r1xZPkhgwsh46O6ezoBsx/xd1aCqh9BPCKJxd/AvhKgwGWQi8vdh3HikQc57DcoS
bpefmbyOzxekAE+hp8Sfu6IcDtndy6meOXq5fZZu+CYa63PmoimWlDY7KYA+0YVe
9oX/bfZVzocOD6WUkeD2awB9f7qKri/LPl0ahg89rhPLlYxhoSyIRPwxH1qXSMm6
RonMjXSiACrqmWL4k8L6c99B3Sy3HopTULI4apUa+rqjL2R0RmhgaVabCJMECa68
cuPHFNxNSrA3zfa5Thc/bM5SCXDUjHEwvClvWKh9NL8IFArsd7Mkf+0dvsC1cQzQ
dF4DTWgTk07gEjNT6ACH9+fig1Tk3Jw3gsKDdhF7HBISCSIBOhYD8yJ2AW3Py/kn
gZcsfmlwaSSaKrQD4Iz21jhsIHEBAemsfFYdj2AUbG1ykX2gJpbvzlH4F72D7mG5
6y9r22lnKTq38cz4285is8xQPtqobe1NMFv1e1O34uc3iECIyWvoOxvUUmAH++Lv
QA+jrFLxKOtacAqMZC9wxTVzYeNk0Vm8BxL7vYV0wv2HvBzvvHqSlvJ8W2cEF98X
JkxKPiCbBYdcnSqSRi/5HK8SfQ7dYS8ysWgMz78qn9fFDGDSpzREBf+WXVfOxZ52
o86iYMkotFbyWph15GhwsASfXua1Y9hNe+SWVw05N4+UkjjZFiHQrxE+nOK5gp66
WzoFj0V90EQVFs0i4jzsMNPSalq9Lo1hmXHCNfB6rcqeRQsI3KbT4M9M2ZjTPqhU
NRYKES/QDahjHiO8mas+qj2jy0m8kwpX/IsTm2UJKPNEbsaiq+wzF56BEa6PfF9f
phT2SkxD94xDOLqIrgtMXepfCQIMSoCSUj7BSQiH/B91HVwcxFwi3GcjMRi0xX6E
jnCfDFEq1PflOUnCZ4/82pVj0l0lyZyhVb6gqsjC1vHvjAyzQcu/VUwfbmvw9eru
aEBA2r5IMlZbJiqrTqMoVgnAq9nR2jq7MJWmHqFgv22UUb2hAeopM/xrtuEW7DF3
HadIeAdAv3bZyWifeh7F89FSky1UEZ6nmcCNKn1aCAeY7YZVvy4EGIhTrsvAK54p
mCbNB1X2BJeudfT6z/SOcsclPwjDS7e0SRywiI1Cj+dgNzwkZEVvO8xOAkM/2G2p
IP4aV+tVcq48ltOf6x+EH/efhXwV3lxu2v4O3GxBOiT6YN6g1x0jdnBZ5tGs7nW2
eglmMjVoQAqK3ts/pPxgxwyg42TLRvVJ7Bm4EF3Q9IakDFUPmf4MPLK0ahoQKLp4
2pgGVqwyRUsCYQ7gRwCUZmhejtuivD49aHJszodb0PjMUxxQkIUMoZZdUQkbSxw6
c3j8AkVapRG0r+et2jQpGADNYpZcovTdjPIyjjKLjoeJ5FJbnIQTOsQLFH1z7+hC
NBb6rOMV1Qxhs+7DS3Hj5WXYEVadePAbYw7Qp3yqVFjnnJ+2Cv4pm90bDVdeuAZF
uGvkAmc11e0v137d817t+FAKonffv6lU2eS/amc3+4s/SwTlRqvDnC91NMFHy9C0
1mHuwO4f7DSnrO4efOyyOmRATQC/02RUCdw4wbpxumJBcsjccVg2gtOqSM20vnA2
GJsbyxKCxnGyPlxFg4iR0atRBa2YR9BPkBohQ1AKr4lXPOoPFONG6Q3im112Penv
heRthAlPI3HG8E69rZF6QTC/NkAr41kZceC2ixjUR921XdRvBKfI8Hvj8AkKW0/m
YQa9qU3Xjq3zuluMjI+NMcSoeXbezYEWIBppVgJKwv7azR3XVDnJm74JNQ0FrwRu
x0DW2fC06Y/Gaq/VdB/iy/lWtFBy/j3kWJnvLbsV2i+Q01R1IkbWdOwKv1bhs0Ym
1z/m/RATsqTPf6eKcHe1MtQdWy17XGK6MPtLVWpyTKSFrqslQpmzrKZWrnOzDU+1
reRlDjPlEwrJIELvLpYGTbZ3xfBUQ+BWYcmba5D9TLdh5H7n4C7U4/Q0P+WnUv+H
mkgkakED4OhTGTQFU3TyiRuVJV2mvtjdToF/xTKn9OahxElKEOJAWCh9CapTS8xB
Q0XR6Nt3W2IG4dLW5+aX2ik5Y7XCRFI5BR1TvvNl7wI8CW5OqsPA2LO4P+bxTQMq
hefdsDv/m8aO8c51UsV5CuDR8F9LCjliY1k+iNu1EEgaAGrwyZy3EX0hWMOM3P5U
85JZI8Tt/RSpfX6Od/fL6O8yITbl9vgO2MKH9+YhAYPIcbEM9C4J+NJ5t8upWEkM
jys65+0PQG7dVYCY1x5yrRrYGmdyr38nmtdvTfY08Kmaqde87DBjJWqjace3jCZQ
crGZ33T0GUUxYaIXWr18thYfLy9boesBnuByQXKSaAa7kP7dWfrHyKNRXasUHHSG
Rp3a5/XIPFS7lpAal9qfNC5np72FmVqPmKNJKutycFzJywJJL6xt3ZEmcqET7k/H
+M1ZKToa5y69mAkOL/6mJ0Cfc+AQ/WqpNn3HSc+c02SfAnJ6TKDZVJAsdnQc5rK4
LP7LuPkIw4ZFXKbHV+cYERq1wsUwO06OgbzkylOcnYrGWDMoGn3l6K0ZkFHXsA8d
Ib7DRvWqRgNr2g/Hy+h+OdtHnUpHVtO7R5Ewy/EPwUfQ7UGTU0pxQ77UMuD7UZyx
2LqZGVWok/WJQYPF8IuxgdOGpVhIqyu0tHRnbQ3QMwHbUkFcAeCnTJfd4ad4Ay1P
VMwal/9uXMC3xlPS0mfN4hnjrT8g6WPucI3kuMtDIlSfJf//TzTZPqT/6+lniTIk
dIle/alrhIvhAOZnYDQtvI7jq5uZWYLn14sjtgOm5FUvw/Njwiz5BRlmqNdDugn6
PD3sDJGeSNlwKdUxvKQxHGdRC60srcyqiGmNGCjO6SMCtoi0xfEPAh5Q3SiLF/hs
fqIANr+lIYqHSy6Qt9H0FCrRwIIYO4sWuheZIgIjBo8rPuYUP279ep5jEo39IDib
5pF38v4IOULzBekRE9UQyQb5OzP7Oc8Ua3wI95tILnMKr0z49ZWFtZBGgEfD+sah
guAGC7xNFL9Lw92Qk5OMGzEPF6o4OAsYefGutcKEpBKa789DNBGtaG8rDQ5MMi0M
JaaCsiO0fGXYZE3iMUF58p6eekZcSV2OKDEOXF0V3ATO909jfyScn0H5aNfo6M5x
Ve/Dmt7JXH1HnOFMslrSrdp0AfXKzUX3qhTaOX2Z9EvDk/qe649KSfSFiZFeFBUE
fyB560Xe43PJ6R96xrgXnhxmjCCVgITlKzuB12Xvo1g09ii1LdLGmXrneTK187sf
3G61M+2GyZ2DfKn2SEQsVYOqbadHPu3J6aDAzrZjHeiP9R68w1cAgij0q6wgv92/
HRtQQ35squfeFPP201okDUWFJzYOBtxps+d1K+B3rcN+uUV2z2kJTuBSCEd5dxHO
uxPEliqOMbLG3h5idiPLehX2GrA+89uBNS/AzFJQLMqSqwJJs/duqYSKp5XuUVb0
pmS0CGOiPGK3Bz7O/uQjOmwLFJvdZKlJCf8DCZxJUH041aJQXGvLmn2siQsBhkBc
pV6vZRZcKCIxClfSF2NbBo78uY0bA42NBG3A5++x4Pay+yno5qqJTFDnAJuVtq/I
ifNpVIJV3izG8YwbNCZXrA8kZZT20XPYdU0uyQzsP81K/CDdIyCMvFh9tqak/bxA
ozuVNe99D9AduwOTSL/Ijuf3ByewtnqaZ+mz5H7tcWCYepMIyZ8EYaU7RDdGk0wJ
azXp3uP8wxBQdgrURizca9dZEd3KlRbUtwibLtoMea+F0KrNPLYFzEMKP+U1opJ8
Sl5ehG6hY4KsCy4BzVfxx0VPYmK4m7shapokW4TC4Et9rcb5zp48vshLr6E1ACEJ
jLhDnKJrO7yrhuPVH6v0YV8VW0u9WCoe1C8pMLYeq6TsE7IdK2y9jzqgOgOucXQq
pEDvI/wOt9PqTV+/y++w+3h6x3DulGrVoFUHYPUOQFmsw8hqxCzoBgGmnq4/PHsd
JzynXuAi7mofitx8pYz3D0TEhBArdeaNug63SoISK9TbkS3nlS7XJCf44Z93Lw83
ikpTdu4EDTzmiWhXcVnkag29qNi1U+d1LZIAYkWMlOmRW81ty0UD6fWZCRTprzU9
ziewGQQGZ8ai0hoWZFPv7fcBqqXnvjVjXMD3UdBGUpKQ0XvgakxFgRQ2jLPUwK5X
2FIVle72MmD0R/vhrJQkMQyG80/dlgSqAAUKjhb21vkqpcLWt6uYSds5X4VhXsME
S2BBHlfVoBUd1oJckDfxErL7vbuRHHr9/UgTlNd2HM5e4tH6tKqrnyHUK5pCnhEc
F+YEyOxojHnUMHrDBhQcGYzELgq3OTy1qi29thmjY+mkZ6WwNjp8S35/HSHwDmb7
MkHtneStMaNvy+jiNMynw5clwMt2fTHGx/9/E2gL1MdtIDT+oyAQXxQX6MJUUpTM
eNNIaC1croyGruAwu53PohKMoMPSr8oci9jWCSyJ5fwJ2j1EXk0YvGYVd4Ijrwtk
WjzRJLY9mH+Wakru9F4OE9bIlrL1dbaJzPIbWuRQFbHxVTl3B3qmBvmpV0ES9OKR
IJ/mUoRwJeJkwYclsmQ2SquxEhlsteUJdQxGAH4k5nNCT98nMx0cf9a/CDIkKlHJ
pJ9QMpHKIEImoAYHIUrEC7b1zrqx/2Zud3Eod+6WTBqcqMUBqpJ7oOScpRtIWMHZ
1ghEBZT1oaG0frTBjT07ZNRF6M2GjPC3HwmkPdKKSFWuRkU7LpO0FCWZlPuxfVoE
c38P59ZBLtKLESC/vTsrDOAPCJ46HbL0WphCnPgeiyPjuEwYYQEc3zJ+NgzZAWRu
RGlWxg6BYpCBDxzFpcys9KKKN+lGoGaOoZ0mzo2xd/HsAdOn4h7FFkykhgRQ8xxn
TX79phwqIBSeymlK2X3RA9wvvZcpHUNtF52kkS2wbd0HEtxUuHg5BTEnjLYQShVM
v8uRJe5Cy7K+w8LWDz7AeJb7vdFXEARdXbQ3xGUK0qv4DKSp2Tb/VE4vgs2PJo2P
AAsO3IVC1NyMSYkRQHyyFyg8izJBXzskC3AvZOQT2oe7LdfoJhA6844Pu676Cmw+
Q/tm098XhX+7KAUWNryyDy0aAoqhtMnXTO7DIjY2qp5yo7gsIQBxwlZdZx6AQi5E
1GRt0lkCqHtQVEUiwK4QJsln9bs/8dGnV6IFU+7U2ASTwLWGxlVnwMe2Tcld8G93
+amN/B4kuiBNV8tmSHXIGsszpycxWc29s8E3BEEkNnXFMkwS//uCUqHFP2B7aTwt
QxTn1B0qDfpN6bif9eWBgfGZ+e5MY6JFov3CUgOQ4Mxp3RXwj05IoIHJtQZ3fTZ+
m7rSPd11kUamQZt6BfmdWytQtBFtDUAZWXFtYjVzlGqNbtCpC58fXynRMxQJx9PL
jIVJoDc1Sqk1jmoy7tCUNMrpIrfYwXbOj8ORygfv45RuohKITaM9drGc4Z8OcLhW
YiArXddxVizv1dvLh+5NJc3UyCoTRSsPrZZkBXUHdC5CSxLiXJh2wiKN/hFw+wLP
Qg3WkzY/0GA3G5tw/WVA1cUAzVTVh2B0VrQbJRuVa44Ndd8mGYBFkXortaiP85Pi
WWq53YXSJkIn6C0bJY+IVkZS2KwmkrRTBnZHvhTn/PFm8BUV6Ts5U/6d0+ctAiTX
Gfvq0DeS5AwiQMvSRJOtU06cDaHrFcI2m/gHEZj/odyf6xDzBiKngA8UB+4I+dFV
YHtOe1NolvFFileEiFiAbEX+buO1xtLI9Io16MurEqbjzR8OrSioZDN4O4Zj7jrn
gpWuvsHi4CY3WGYgqIh2jdobmOPZ2MZVNHC2x5OIR6SFrjZCRl2TBJ4IZ8KUvTpy
+tubFDjGp8D70nTRj7hgjcxvF666Bc/tNpwn4HlTwBTOzGrZSH655YcwRvxEst3K
xwv3HKWflOdLWOaei7JQjZlxNi8oBjuM+XbwvXGP/HHDIkCn3Ec90zhxLaU0SS5F
Sxxx/Oq4qACfjK6vjbgskazkLbn1r8X12o3QVhpQ8/lWqAsbppNNllNRuPMnVKn3
gw82BJRyoawGMks9ZSRYlk4Go4TDMhjITY4ljWZLdXltaVai7WIDDpyVmy6L+hrJ
hACP5QvuKitlDbOL5mDdaLsDzC4Y7CNGCLAamQB57AQUmCu6ITg+lX/v1EIMOD+n
KRFvrcxGMgxmjwFGevjY/EasaG/EnjfZ3vKkiC58dHyGizsO41nWDItGxHbqidon
92SQkNgzPsIBK6702N98/U8AOG9k9IORoiLTb8Lg6Jq5bI/F5B98TM/FZY4KBbKq
FtW9ECEwMPqIvovnWH8Ss6pFfIX4d9dJ8P5/NOYoTMrCoHigbSTvrtX3lijAKRQ3
GkrNjXfKd1dx8O4pO2f0Pvfm+FipdsXxSGeqghUd7+VG/taD5wExrXhoBxBzang+
pk7cHA7bE4Hy7ccRG14C2ehSLIedMCwe0fQMujOgADHJPrx0ZsfzIDLaThBSjyjH
FSS3qfra/D4isAW9BImIw1CFowrgTv5gXlvAk9GSbUbfNv0Ry8Up7L7eyfE4NXoF
ze7QCzDASDBzgM8RfEiWRSM07Zwd0C2qLjOw2/9GSYO2Lnwf/3iWEWBlaEiQANlJ
+c4dfQeau8z4CmfoA8JSxiZ9ICaTOwQGf2BnVUE5orhUvBjsqFQkKvpwBGpW3HIj
9NEZdzzNS7iQMBw5sOv02qj2ROpwKdqYXz7NKl7qkMk3R/HxV4YKenC0ynjofCgQ
3t/Ye8yXTHmwNyVqv9tHKjOtXyX41c+juBPiJz3YjN6aZQyhgXXuCxnbbjZiAWO/
HKX5Kn8rOEwipEnzsQvdlnAHh/YqcMAQAPNkq4V5lP0MNCN3u2JbOcWaJw5gkuKQ
4j7CQTvk5Ruaa2Y45HVy/mLUcH71xCXLBIrMD5OBtUyfjt/gJ0aNYtQG5ZOxB81h
PW5VWC+ELCu2zXHSvDpzB6LEflyQcxtqC/LBydeu7sqjj1unhi7qH33Q1Z1P9f45
k4+jPnKXEJdrFNNxOnUiJbdAG8zyGSCnJACnSLcqFcod4tClZsCBiaNUxDkaut4S
FfT9ny/q6lGZTf6YIZfiVruIzdmDeQshoe5FUcWuQ99/r3+7EXJrszSvbMdmdKcV
5pqDk1LqcUjRenc5Twtt80P5TKKha5azMuXQTeHB1DoO5zLbd1siDxi+wE4mi7iN
fMH2V2keqb2crw4DUpafFuhnXxERa6C4aJ8g7DTvmHERz2li6AyUO+OjNgbmKhK7
W+dk3vT8trS3rzScYke8io2y1MvU75//UeMAb+E8XGY4oUFoHQ4iuMoEYO8ySJn8
rqy+JaJg++I+k+C+X7lwY9uC2UmOiDqGdZ3IaK/gDWQE7snCwH+Uz3v5KMoMR47l
RhTxhWPp+BsCl+KeNswmQcS1xoa79GAw//uyHETkbfSXfEuaNAU/5BC+YLf7cIN9
cNW+4AD66tuXrIaQSsP7n8kC65qzBmtnXFIZxlxzphlHrbAQdgb1DWZEvYLsUY2W
aknX6oED5OOxTun8g5aaSeU69+5eQptSPEmiSUTzz0Lx97Gf/APtCmTbzwKw64KX
5yTy7pdQvifJ+In5zo+me+e6PS4MBf1xqTguNHT6Dp0F8y91Q9IH+mohiavVXZW2
IxkfaDvKMAl8Bg5MrAQLiYwPHflaNRi1OkV8QLAFm4HaspZRGaDByovwcpGFKKqA
Y7lszTDfOEQnUmVNJMQaYolJDMJxj6scseZrIlg/pmRXWTuHNHiDwyw/X9lAgM9S
PGg2626KgC3Y+Dv8MFQdm3VYRchyRtUGCMIwdazGZAns9PhfGEz/PMi5xUe4BwYg
i3/tfePkHvTxW6oumNPv++uSr6ujlnLVoqjGuXUaQWqCXP5aPnK2TyW8ZLAYgHmU
m/EPD+t+VBYBRzpSfElKuEcRTaeSEva5L76HXW2ZoIbz9NBoTnPstVwPQpPDT5wG
NSt43MK9/uiJ35ngkDvSesHio8OMgNdgLSauWKwfJe4iyJr1Bc9c1HGvkxTlHwcv
LegG4sYGf44p0Rodd2WUxbbi09FWOSiUY6CTYm2O4hXmVGu5nRmmLvyuPfnK+IDS
59YJBJJDVLAAhQtyCDihBguhxJHs6XscFc4tSUW0mF1w+Elg+VmfnF1JmTcyCuFG
GDkdsV28vcE62Sz1V1493erND0kzG4YkkBo+uvHHNkcN1d9tGmmg5rEoK9aKEBim
03zstMh8ZPGGIM03BJcneSSnTfnutBldXALbKX8qPkmx6mASiSQTPsA5TgpK9O8G
WPPwU9ykIO3muKiijd94JvJ2vsCNZLRGHCaK2d0tOknoXs3Do/CjOtHer5rh5Rip
KhWvjLrRcZYgRg5Fp2N4jVUc6f16SYFl+xlJeHF9mmfq1y4iyGmkOCwLPkvTNYsn
vDAqz30jtL4NoxkKGk9EF8Ex9RYr8w8l6bqvU+c928JBzSvHG0mSR008zfcx6eWR
9ftMwNTGoNbG3B/FyyKfCjDMSwaVIjtq9KzJ+zJ0KEb6X1f84ww1lcZIyqrdYKZx
tfJuTjtd742OFKWQAa2RDoNdtlZ4WCC4inXT7AQXe7q671poqPWp4doG4Ao/KIE+
CcSoB9jpzUCyEjCGswJKTJQlUJg3EeRjkX4I7DFI//2HRRNSxuG7KLTPy+t60xzM
pIRL4e6gxbRzQvUoEDbCjTeEf2l5iItDOnckojTDP4wGs7Gb4xkOUruk+m0mYe9H
YNAk0cPNGudTY3rCEUy96c9vxr8VMDEIXLqWJ5cSorFWsaEbhqm3PGBAV881SCEb
rOT4Mp/wxNyjCKcP8DeR7pnzRum/uKWIUjlRotRsXmFvHdHOSojiPUxu8qiqXbw6
7Pma7ezUNPdlV7vFu54I87WQVKj9vZbb4vqHUbEkIF39pcTyaCojvnkl9NF19ysU
DRopHxnWiVuJfL7SKYLh+zDXc2dVXrUDjcbZYmYUWgN5JOB51BJ/xcJhTQBdv80C
F8pCE99iekWdM7mO7kikmubrNGs1yCZrmCsps7VkDMQXg3oWsBzbEJbEaa+fBpa8
cwD+iN0uVyqEiIBfSBtbnOXw9ulUanvW1zjRVfwngQMO90bpCPJpIbrh8UTMFwPp
Lu07C/Txn2ftfk7Ar3PfZ/BQWnV3fHgE8c829rPZd5NG6tjXJmeb+okOriIvXkA3
TNMJQynJMARuGnWmgRZUkxvLlJPqTYtDdOr/tqhZ7onoLse03cloPce8AIqBAe5W
2Bj7PyRRwupa9jP4dvQknOufTW5bOecHQOeyUyg6can4MynzhQfURdlgRcxnDuGY
QMRUGl5q/iuW0NaE2MWORnEeJqqH4Sxzcxgy8QHE9yzO6DXTGIZF0SGzHbT1C4iw
DjSv/t5DIbeGF6JDuGN9jdFBEXekOasr6sTmJPzieqEYUAOpwsg5nOwzieIc8HDz
Mbuu6YCq6yGaxvAALWbrwciJtGmokejvr+YQKOJaUs/RA7zJg6GjIsGEWwhV/9Lv
qz1aLLHBf2zk+HHZtl14ksww5GfZ69eso21gkPUW5nPI5FJDDDY/4pye83hJTdKM
Aqo3AbY7bSAKMPGb7hkYSUj4jq9xKVG6gvQjEzxcpEL76tMr6mbQfSTe+3nlRJfn
4O+2A4VkprFTqKxPYKhIoXUdw4XAUimnB7xRnbOukr3ihib2UbBCfjVhWRYBQyhb
GKiE9xZrw5AwZafTtlfDCJ00kpq8lJ4lxj6nYydieXrrArtvJwgPQnxR9EsgKkaq
bvP3e5R8l8S7u8wpk6chxl2hmy/mGEwvN/V15pArg3VyppYYdrWyOBiWYSnDl/6X
NLA/LGsmuPy2vfCOur/2Zd+9/uf/nfeSdTkg9YcFW5BzzNBUZN+qTmxVUm+O5r2U
kASau9qg7gatAV4mjdgNvG2DMaOLYpyYM01lppFPQS6Kvr1m8FA8EMW0yT3eZpJk
/tVpVaqP8q5/+2iQX7SponBWX+XJwzBfOdzmGKGeiajLuZ+97Kuv49TZjxgoXGbg
A1MmYSChTS+NjBqXihg6H3JUSLjgRWK1dki7w2nS7+/AYPbnEUOihW3gKXT23Lec
E5bQ4buQcyNR1seAMZfS0qJEPrX4v/+XeMd/2HN2pJvXIK4+ioA6GGEwEJ6BdWrV
1HC1764CFC+Sx7p+59lZuZpHT/7bcUDryFDTNsdJd9YnAR4pHdzwxG7ZBSuQ3x3k
mNA2j0Ko3Ok5I3h7WTP0gzjfgG1VoZvm/PxfRHiVMXtRji9mboZLRyOR9UyQxkgT
ILgCQY/CfdUdTvGotbQkoXnJMyB751wyWcqzsWHk7BysXYuqKTHXkZ3IffE7nWtd
FifUaMNxXKlOT284Z5vG1w1MaGvIqf/KzjICyy2seUu5rvzTBcAWFZHSFcQbsfyO
WUi0nX1/sau98qkhPnxwaPD2GEIdLzev4cOit7+1zTtfoiSbyVkMaFupK+h8Z5eA
sKIMX/2R8MkNi9R7g/PQKTzaClCKud1sllgLYyKlRHabLuzTLkhqp/9u+h2VfJpg
7OYtiZG/KxBYPAO54D5FYuerw8noDwnGN1DWDdUKdfs9CXM2gwH2N0trt7b7mNWy
Ac7m6iQmrZLFdnsS7LxiFQrWC29ADDuupI+VS+nCZ8QzsvK15E5f3npPAMnpvZJx
P2DF1t88Kz5A9EADGG3DKdSuFGvTNatn/C2budzu5wkUJiYM4IafFU/PvhKB6u4Q
u3mNkucIzTgUdrZvrne/vxPwkTS1qq2dysTHYuKqqQvK7MNZI7mZeIGf8rVhaFoa
t3Y7EZgTT5YwNfrATXQo403t6gQ7t8rYqrHhfahlgN5Jt7ahOatM9xHaQfoIWXMi
/EHhuv9PgzQV5GfcXLrwMuT81Jcjc9Ivk+j45nFBTO0cs7JqK4gob/jasTZuRbHR
fkKcOU89rDT7bgPR15imolVdAecGFQ8bbhCNYN9oCeCKtOO/ruB+DTN22zJZSVZC
4kqjgXVp1+y3KrFyI5B5MPdYCKb3zbrAx/ulHT0HPDm/DP14dVXypD75DrzXzArX
htv+a3eFZ0IJsndtbaGpa+LLyUTieIR1eL/NciecB5Hv4Bv+rhiIzIwT0nB/7jXC
EE+CxUGtoLhc2oS/CLjeiW6HMNZ03DssC69J+g7PqujU/YYUXE8n8XNnC96iLOlg
6wOUqcJMJ1lyLsAgcYEYl6ZAD4k/YC05ZNoyNFH9G2gBBWCR901FWKgyTMGGZfTk
Ly9oQx6YeJx1vdAODJTpD5rEenHx/C/uM/GDsObxlBAU02afHKgoOMrTAwJqJFBJ
30ob3Oyib2bnIv0J7r4c/2IgjWFWhYfGgC89tr4o2rJ14wTb2P8AUejkaG7waka8
J+rKo5kn11rhBr/OqVbDlplCWyGmC24ULYb+DcZeN4tSdfz+C3OjaISK4GBqIAp8
uy1f+Q3QUnOt1lfTVXgSnqS1orVVMoPdlHjeH57j4BwIH2wyQfkJsMQEwCv8cgFY
4DbvX0jtFfGkF1Gfx9Nx2d3uk2xb90T4FNIOovTQzQDRzhj6GH//gHOs/xDQSf8Q
U7aSAJfovr7YEKcBuVc4iUeRiceP7yO7tv/OEsCvjoBsbndPyYSEL55jSCjXLBcZ
Sy+r/Q3ljQJd5J1czNQ2nHCqQWBymAQ2UebCDXUddjgzidMGewky3R/gxt0NB5Dw
y0mk4hnMPL+AyHbEY86SRHndUSi9dAYfeIjhe1aAqJQUF0vmyEZdGsLs1E0JAJRy
Ph6XyCNMIvRWFGZOXFURZWSMsVccpJJz7aMRtbE6wV9sZNWE09ZLDDZMSPoGff32
pRud1zOLJqWfR/go2ukUJWgwL4XbK3vZDRZXwfkDUWByFUK/uY35kOfPVi3P5SGD
BjgwygMbTvPtyEAxwNvTVv374iXwQ6uid8HBAlbfT+mzHQ+bbsTjP1Kgim458Ioa
NNpl4Y58+m1As7MH94izGFpdHVqVOHFOQJWSwxYRTwst1SXqgsYsF3JGbB+da5wU
IW+neVMKjWbrEs8ZqFX3os6eFq41ASK9lyEWeB9zkvZmr7a+coV63wKV5ZA1Pl+d
5n+iXToDQ25exRpGmDXescrKbnVmWPMJAn6tSB1I1MieFYWwtsP9rDgUlXFgp1qW
owOWITd53DyEGUNCsqel92OgNJsjMeNAMGqgZAVblqYI5halx5GCpXXRhlR7vBrf
d26Amr1w9TYdMPRTpkvTF95Lzzv4VsnMM/6WWQ3aGZr0HOgBq8VeeaQJtHP3tWkV
0Snp/Rgjh1v0zPkiC82xq4eZfS2md+uG3U+LP7XrKusCQypyA8W+ut2mnYEmCtQQ
CTRMY4Nfx3nV/dgajP4REi/NxIsY+zBooofZ4mduuNtzCUh8z5IHbtbsdTR5e9sP
XBk4uIiUfzK0biSx7jvJBajpZ0IsfgqGWybyJwlOzc2s+W6TMcBQbFcnrwiIw8Ft
S1JIiP331dKHXPdVoCCplQoFLmCTGBnG/FZU6sMX4h8YTOhQO3EscjTviZ8JUAmy
vPYt/4IL3Fyj1NtGtjPIp+/bbUo3kia1G4/rvv3QM/r6+XRgQK+glwan7//jycIi
ic86TyTA5CydHAzbUw8pkJoN9ggEU9q8SuIi0mWhHXo8OdkkNpfl7UgjdksEJ28c
zHGs7fGItI8WOsVCDamawNKAoS1MjUXujzak1xDeURHGJ/i5avOK3DcRiJvSe/3U
a+9pbmRDfJMtnrVZEPnKd6f38AEuodo3N08DwfDvvocLRjhEB8ZKtJxsieN8P6V6
aZVosjDbtboZgFgvnXIatKkG+fsZDtcZS4CZ8nNuFNoEIeXehElVxtF6Ss4PQ0ly
WSxsa1RexQbFkAyH+bGld1ZtSIGvCxxsxhpTNG2pdJy9kjf+NpkzVkJcd5jRFs14
I0SwYEXmvVrWYXnsF66q11ahgQutQElpbeYOTcWNEsUUN+ReS9Cl/3QSmlSIHnLj
kmbuE2zTOtu+E4makN0VEimP5quOJ+KCwsqmTyGBFyTH8mO+fPNvHRFXS4iwcnAY
MiD6k/I3rZiFXaPAeY69EJgd9FNjUf16kzAJkuwTOp9vsgVGsqZwqD9QXStys8qy
p930fXyDhP3nmVF4aDOHej5GgubzUIObr9rha+rimNpO6NcTFiu9IUIa1qTpXvbW
wnPUR4SPExthjFZ3sgXyt5KU6wBJ3Abo3eLYvRRAY1aPaT2HJ0s1oo2DaWXcvmKp
EqkQWl5n+MpHU+nRG4gUze1b9RPDy4XM9yZSUm70UJq61qbieV5s7MY/QF5308cc
tDCuZc7JCjHF7Ms3LPOxlY+fLYTC9DBya6TXwwqKg3Vt8EqYV1FNw8qt2RFjbVyo
xJqsT8fkjT9T1cIMum0K/yy2VbM1AXmOaj5gVRNFJy6Mdltzw7uOrm14ZSMCqZfy
7y/Px3ZVV1TodX4eWu0/glMWui4frQNJHY2TO86XRp4lbPkwznNxsvHQ0yTevsDA
eCL32mDykwfeStrCHjA093NzArCggzvaL3MDwzpPQHyYqQ/yXFkNUoFib4KJg+As
uVX2yEgIbRGjEszACXn4+ET8y1uGPsQIt66zXEBD6IBOeQBzSZ+D7O+eiP3rWhws
4PZ2zMLsWiJekncr/a+Bqt3CZT9T8vX4spWPE86FqRAN6FrYaKf5u14KnzRbF9mI
tTcq/RS1i0+5QuAAC+qxeWT1MQ5qoSA+hY6YrL+oXRZIZhKtXY3t+LIxQB8B17hZ
QEg2sMTVmKJKe03tLRJs6Ffx1KTodVjMFzpCB23DfEC9iFm2xXb9InBc8piV6/UA
BDsWj/k5DSRPX04o/b4XbZLt+dkqGfdjbmue8nnhp0CpDvVDWg01Ay9xY+KYqsvi
pIcAc89ggLIXPoteWDsYg4cLzztANMtQuHR8eX/EWzOtDRkkpH1PjGs6eS6VBEkp
yUcgFsGjKHTBSp00RSjjt5Ch5to3e5KGYeLrY92OBfo+rpBam31FmIODMqWddBse
/M3P/R+IzDTEbkKpSYvZ2fC5732FAzJBkZv60dHOoDOsHgNEEPtpfSBw/S/MO1jH
/bJ3lP4qwMD8vYrbdHvb1MhZ8wHpx+GI/tpk9k9WjCy57YgZKpItg3YDnTQt4RNb
qI1JO6aaVfr1XhwtXovcoZsBZHk9L71179GPmnRay1UUba9U7b8eudV3so8tqTgo
0wdxxDLdFSdqe3ZDXCN8HXVGC9tUyM7HprU7VvQXha/nsgzkzPjFQhxoZTJENXGA
imtiW3urot+xO168mCyl69K8qFRPuq2Wbc5UYQdc+byiS7PhL1VDgndhsgNZQUW3
+Zey01gaFHjoW+/d14WwHJ9CzBb6apaY3PkM8HmFaYr9Byur6SMlmS3mDmMlaQzv
sXxE9HdgOIlU0RRyfSEL06L1cJQjxO4zSL8S9TT1A/Le9moEya8aiv2+RqBwWGIO
FoUgcm9o7bOtFiiEa1wLWUoKtum31WArwO6e6JLZlcU18QVoVH5mual0wuPrWOXL
ZjW2RL6Cfb7OcCK9VTKAMMa/uRN2DgcaA9KKjCLl0esudAgwomtx9qzoGWtKNuaQ
DOaE/bURSpOgOAVz+3Hr35P4ToDks4bPNuKoOlRrrrF6yr1kzMBmc7ldq/4j+YF2
x3YnU6Tt7yPAEOTR+qFTIEnjsdz66D59Ahv6VqWxOShgRHx9VEdzO7p0GF5S4f3G
LweaWQjXCJYEc/EjnFB0f7DY6eKPC8k77NhRabG3R5r5Tcbjd3Njln15kQ/B/MfM
B8kv/VeItZiz5oLj3srbrojRBPByS/vkNgR6ppFpbAChhVhBQ/2tJYU0VqwCN6mw
hReY6D6p5MXS+deJOgY3NJ4FF/fd/PHWz+uIO/bvha/+H6weQny+bVIikDynzWN+
9zD04JFaoxP6/yrnO6e95d8iLNgjyOwwGkPL+1RbutHwC/N0P9QCvnYaYQukZaA+
ED6F4gkQPDpsshJE5hEe6puaORodnuV1yzMq7pzAau850UHfQQ4oZwTZmVAbMU40
kvRmXp4IVm8LKTuoyoKVEDnE8yvJhJVzX0wTFZfO60iuv+fujE3Pae6teno51S7I
P1p7M29klVrLd/XuNIZH9KI6gPAhqaDpv4TG981FXKF2GPk+oqrsSUiT1KlZd94F
/6nHGMXOckEvNTCKaDhdvy+UMYEtNbJmXWrA2DLevPR2KoX3gBLJzq0xfAfGuFhl
VSYLe8QGWtH41W46Drnco9vCjfsluXdBMiFP/Va92kgvftY8JEevT4k7G5TVSDIj
1muJEaV3YPoiRI6IFqkKYdZPXtH0Hq/74aC59BY4AZVIX43BWRi6H+gZ0hxt+LdH
an0STd/DOsBlugawFYPtPfPxbuAeBkPHDLM+dQWVB4xJEZ5gI26N7xZCxs4PrVkh
Vfjp0L9jUC/+gtcnrXqh/P4FVtWIUo2b63aTKXTRxCioiBp51R/ndx+X+spEvROi
BKFCB63gdokB53CruVMZaHeA4hA938647FpIxUZaRHYOXQB1vDsw1ANABUNc5fQp
Zj7tyO5h5/P6FeQPZCtr6PA5CCoskG3E4ALi4Rjevl0fwhtSw4PDJpSuOCRh9wOo
5EY/wS8wLAS8IZuLLibgN2EgQy9QRRN5uMTVz5gxOGnf3crfcV/KUWflm0sZgJbM
D2KNYzmarEWbd9kPwVkkII7A5jbu8QT5HC9L0cFfD8s0BD53h+lj+J85H1ltsolU
3zdsGjIbdmNF5Pg2Ae8GGtbsUFy/4PWUVZMHSXv8aU7QyYefqvFipoBzORfhWajg
Yiu1OTu+wv9HSEKTVKnM7DPXZueNbqh4JgSRHESDBMVGI73u4IAgkhXe8R3rdo0P
gFWCqzOE78o6mdE2MaEen1wVOuicDU37sLjLeEV6fuSjmJv+WVpAhh7kRIQ1frMv
SXuNV9fE/l1QRy7WkFbaksWoWBUJAMQODN88fqmE3Y4eP6StzlBVfA0d8um4lDKe
JM6ueWE+4HlKjpdUfT70EeC61AUnViO2dih8kS+j2a5BioPz9r7DCtemxhyk2I/b
nx0HaGRYrw5zZR9rDuLJi/5+S8Tor21sj4FG+7eLwme4MiCH+myLS0BLFizYY0wG
CYBomfRlMD3gOrUcUApSk8JDOm1r0T0kkuBuWnLbKM8MtfLObX4y02/PtaZIAlVg
PkVUKPo2Pg/xmTT/WXveLTTZaLlOO1W0OTweCWk+Ov1OiM/u/pT8R3IsyRREiIRc
IOTMWsNIkE5LnybY2xee7V0l00fIZru2OWtIt68Ew7ARrTTQo/WkQcQzEiRpG3xd
Mp11KdHINimM0w1Hht8QHl1QOVWQOc6sfI0V31hv8n8mK2P24uIpHS7JBaR5KMgY
KGhSpUH9y5ZB64TL9N6xooylga+IFS3NfVxhwFAOclHZDDD1XuAyU4mHEMaOUrTh
VMoyYwqXL6N2uguJZl8R5HOb5HFg7mR/H/7KA9NWcW9yHNl6hU4nJJTplT2C2+zq
o0ezus5o+MoxdQw76e4Pms2iHh6RjE1y80SbPbWHh27GMNy01EqnSnP5/G8ZRka9
CwH8f20u+/qQlJMFPt9LFh9hopd8dp+AmRswriuWtZUOV5g/yvikyPQQsWLRlULy
GDxYzkGVZ2k2XoD9HXktmGhUiFEka6TrO/LGfJ7u4/92isyQotX0skY+pEZtWsXq
dIxEfurEuZWrj80uQbmMy98tCDDbmL4cvRzqwT2VHK7d1wnl/XXNfxzg51vg5C5X
2/96iSi/aImV4C2cT6bvqfMWQBYxQdS9GXGvg7dubUcGE49cvCofCC9BZvPwYw32
TBipTkcRKTUaKIFiT8z78ZF+FqxnQdepWqPxLsLYULP117l7SwwQtur2506BX2EP
zue1Io6My3N9IVXEbtaQvJ+p8rqh9JbK1puWP9M04XmxYoHIQ2yipDViJ3f6RJYx
yB983kmhQTU2fqMcZYRXZoPgYEjNTc2Cr4+IV0p21FbMoUGmHbm8dxtZPyw9UBGA
2KsGJmAzMar1itkJAzH+0aDFDQqY6QrO66e2RuXdWut3Dzu/tzMlqKyZ5LM6JJuR
UT2Wns0bMvAW9cQf8MSG1FtC1GTxnAbfo5JjJh/lsY3mrbL8aRcfuF3Vwc1MG5r1
KGbuvxK5nsacbQqaoquJiJiTKLSUdL6rsGLV/Cg6mMmHHXy56J+PIUXDz1ObQ1BX
0BbLUhX+c+QAWRBFLeQ+wD2SAO9MaQ/ntVpmWihgA7O6rFl0wzFs80v/HhURO4GV
OUkqEMv5/9XSrYJaSTqkVyneiVpef8awx9HXbzV7hX1CX+3YmkxpNK995yV8mScy
bk0O9LMMxXb/6dpRtNh88svZsbI+KWffzH+YviTgSr9zGXRLbnVMsnwp0FjkNYC7
ChYvlaoEGQt7X+5bAP2l7HE42VcaCPa5ywarUCI619QHKZmmtO8IotQ7qE2w9uHp
aELzhHP9Z9p79mgic3n5VhBZWhPhwSUZ2TL11Kr7N0a2BJ86bty2iRzvxV6s8G2I
Tp5R0Z3HYG1QsORCxr1TQ/Yvpl0py0WNQx2WjpZEUmlOksryujdqxQGApPT9TfRR
2gMdrf77q21Nf1BIrRwc851ZwEsF4gcv7QMZ/71+C8tR8UgmA9gI5blbrcY9w1sU
Mp0wg+/VyDFqxpH9WguCzSb//z7S+529o4vd8WRed2yLtlWZlJRAQJIlquFImDA+
UwfVB9ZAjGd2xY4ZlCMU0LPUY9mLYRvJ79ftIImkYlhcOFqKG5DKHJmM1NmrmJ2Y
ENUcis7i8X2VE0moIt8VLalDG5hIyu4l3fHsdJ4UGIKaNhXNlxdMy4dRJ4TLA5OD
IZFz/zDR4vmcLeSuKbgLs1sPPaodAlc7HgiVb6hB+hXRZHQUHQFrLLLVPIOZdPxS
/7hPnLp9rNvpGeu+KbrhfsJF4P3GCqdI65vTjaEaF7Ql5E57wAuyT5q9Qbkvh1uv
8GkN1cb6ITEdMbWYnlM0jUjMkzKQKQ6HdXK6mY4uMqjLATPXPlu1ck3qDj+l8JKS
EeMibDuSszgMorOHpWv5mJVkv+3m83CWieNnqoAmbQUVXhvCjqi4h7T+EgsjP9wh
LovHcRMmBMNMLNzfFrFs0Anjx1UmVQtYOasMvUp3rigNBgla5Unu3xQCcDasnyak
vD3MEKSpJWJv6ERTEWYkaUpgh/AcvmMkfOM0gwzC6mMazwteGhTPHVK2QsUTkgu+
LTlQtCvUm7kAdjzSuAUa7q680JeH5/WlNZEfidle600GOb5vZ8eW43Fy3oQDNR3/
0oln7MleMeVmRtLl7J35V5IbNAaYVjg63bRizvBMZi/KdacnMGMRdMgq5pLV/JLP
u67JSTVr7eSiIV26DUkuUGtye9tyzB3Ihk8khz490MyJwPnPfyEZqe1IBUdbUd/D
1epuk0ItdPZlA/soXEBONsCDUib0DNnX9bCvkGk+FmV6L/fw2mAh6z5F/JKjz46L
7qqWTQlldi1lhhYSmZl1pQClqoxI98DRknV3jDDuiAoUSotljDvOsJroVlQPuvvO
kCWk9a6K4C82eAXC7yhhg7InRUMbrMJ1JPMvgKY6v79qbk8zstAqRdLVyIBBmUQe
4TrzaZR8O1mtubL+Ke3sTrlo3U8QjXHRcHUcOMVeHAR2klVPav+VxYZjfztHYnaI
6iOS93ux8Dkv1TJh22DkKQ/FKLGq+JxPzcw6cNXAQvkRPyifgGoFOnyf438JHsLk
YQqnLXoGIOxnjvxmg0jD307WElMeTcFLx7UbQFIRNDQc0Rruwsz7icwYn5kEcbHm
CCqs6eFttLrS2JbBefP8ZdSGfxKtsdPfXa+uaoBwI4UcZ/+MUUF1pJnCJ6FataZW
rHqo6TZ6hVvYwygdwbu+U2Y1iJoztksGsNLBYVT5Yfh3S11MbcImwZ/U8ull1fqE
YUXp5COoXIFudUcLC0EJcF1GB3e5oeyh7l83u4tDtYAhIOmY3Ibypq5NKMJPGYEp
sX4qbmTrF2VMgeXXi9Ljxxae0jA8+4xuHmatDB8+SfG2YFvEByfcp8ggExBn5Ur/
IhTnSHJMl1SUMzKyANtcJ4mUDvmKPIGoOQQIMGJ8wgASBrXx0zHoKWe+isbL2ry2
V4wSJLIqJZeidUF7RpOEq9teoLnt6w6Hf/zPnPHkY8dJF0yprag8MSkKdupjN+f6
kYHy87dH5nTCrTrb99+nn22Qmo00AlzIDKcH98JASeZhT7S2fTwisauJqC8p9JUo
sX/87LXNg3QU4Ieja9cnwhySVh4E/SycfRvo4tlUgFhVyizDTbTNWtueXuiDLsnM
KoTdKCDSvfUEhJ/ABnXNO1sZD7yqfwbQwAAk2RAbHey1QZ7SJX+XlgmBrkQXtUf+
fRQ0vw0niiKa9dF6SJdrE1zDMT2k99+/ZBTRXwhPdj2cbem9athQtkpzwgVjWozr
XBrfHFxTD5h2kJBU+chHDMNy47GaAA2Hqzq/34NSTH34X9M3vypC9AengSUpR5Fx
3zFAyvC2V5+MBd8DuoEOguZbZad6GDBteUWViwBhoBwGGrzqNof4nj3NxN7z2igC
eqE4e7ot6oV9yMX4yCieh0j85nlE1UPyKYzWwn+2uRD0ltUr7qLWOa+ysJtkr5RP
UmcrsNXnDGfVWt2Lf/KUUAEYQd24Y5qXuzaNziNsKJ8xZhgp8zCqL+5J3i/sanso
HOOCIV02uv/WRZXl2Reg/1IHCAqeHN2WqATbkks+byQM8LCI3nRzkDdRBPV+2A1T
v/oQXEjVVK8fZDlmX6wN7Xz7SftO3PoFQ0Fvm+22oIGaZOCJo1jGz2yrqsgcrr+c
Ugas9kbBTNSTMwTCYbfmPFJJ99BCYNoRc3lEotN881//RKXwbHn4gfZwu30DxO/G
lwFDTk3VVwq1Mlv+D6zJG5DgNq5si1qVYRIlg6C9sIaiyfEW2z2lJVx5h48TUekH
ckUdUqBrXPKrtxAE8KPTDUU2cqGFdc/Lr+4vvWvnK4d/YQRCM9ttAIvpv3QrQGka
yPGvnziBgkjEdYTBdeNN92OBPV0oxy9xlRPEkiB4bbNDKtoGpXPjZaCzfWVYcULX
bCv/SAhZziseUaYVoDfk6RUqIbRkf/rmSXsLdCUXiPQtahKyLkQ62Tyt3eB/rZQh
kDKITXOjNW044JIH2yiZD24CQodaOAPisaHAPHS8l3Ahm8m+IkmyciwG6m51zi74
b2mblGwyvoHNb6HhDzyjNlO69ACNNHGMbNuiV6BY1wRpflgr8PZyHUbx3r1nIUY/
2dDGjSqaNEfhbmphHr8LojbLPoGvoOv5bRNYO48FPdY2WfgM/2Otixr+cGEoPUv4
zMzcIKO7xSu5SWryHLKHZr7CvI6J5auVlnK0xy820emS72r5Tsct+G/mtjXhRsNX
+Bbn/EHBB/fb9iI/obfgjnXeG1DsHxixBxnAdAG+hXXMXSi1QsC44J1vNgLEblNn
aMtmUrp5OlRHsGqO0JKK4y1rPmoMmQO4WpAXJw3DIMuC3TCTK56LKWZQvqctucAU
5Yk58UusQW4RQo6OXUI4sNIlK8adTx0QWdPnmez2QjmzuHwgDRVDG4VVpuxOg+XM
8Bm7MEg7uPCOwijRxrE1NKtjgTVJC6NOyBYZ22G2Q/uXYlQQ/0sj+tueG1AtG6dI
o3cREfz/fOBJMHzOYaXhTqtCvwV/Ee/7tY9agDbP8s85LtEdpvIEkoaG8+vTB5UL
bbMj3BmaehsZ2V8e8kQb1DgvXv+iTRjWlO1WHHvSj7/f9dt9WQbXlwxn5B7eWoPn
sf643mCkpIO59smjjXwC7jL1fsoybiaLhYPpqlNniXPsznJQ9YVCbRJJBZVhkn1k
hNn+yHM2TLojpsekgnu1hZlsOyIAFttIqjGMRzNIJgk5KdACUsauJHpPyXzR6eQN
hZBaDa/HEg58H4C2PXDyc9YBCW4K8DzRGSCsESWKlGXC3q8eeK/EZkCYmb/kVSiT
zPIhM2/vzDzD/9rAROpHVWOwG0j2TzESCr0qqJIQI9dCpfuUZnGUwj63ITGneXBf
3MEGkQ+mXpxRNTyfc/f9nIXNOq8H/z+fzcXd8wUL6byQCwhNmqZgcRHQlooWjl3t
SY3ksVtZE6jUM3t9I6EVz5TNc2bSvuFqruQ1MJID0NgKixYeAQnFbHMmd2MK7TmO
m3REshD0BhvymkucwigEp4VwgpSomiipl9aEZ7qZ7yQjA3CyrVooxy71q4zSIceJ
8PyNR0CU1YwxIu9wihWB9TRVgVKNAYkgFnvNd3J9DeaG1+hkvfsw84/zXW4Nf7+M
ClzScfiU6Y01hag4J3dQHiGZoIZwKHXq2m0KCbKuakqHAIEHPE9rFfkb/FK5I2/H
GoTxlCrlGnwD8VwvMsBSw3RDN87ViVwkTOqj18FkirsBr4UAKQyXktIYFUBM8HyV
/3ixNYQioiOJU4jdnuYc3sQmCAdtqGjpfFnnDfkLsIOz+gV0pz+460TTTvmHEf47
zZfXxGDaYWUN3fTOUa2Dy8EIoohXc0srf8C/uH/q7aJgsyW1UAHwB2E9s3CiePpQ
QQiLw72lzw04jJgnC6VS3OXpz/A5P4j38VzmlWO/KtuL0bWevye57kINiw03ty+O
TtRYFDPu5jBxUMzS0OIH3AqpIFMbT1uWLM2cOVRUoC5S0fbsHhtymhevOvQqU/5y
r4hbwUBQ1389ONQzRxxW1DwM0dHJOsJW4Y+neRPhtLCHjCt+tVv4vyWGoY/+DNHu
2q3UCswKoGxNkBeVxQDtce2UmXfulJppzeQ+AYc0zg7xpciOClv1Zf4g2oDMQ1mH
TbrpRkmPwqTHxD1mvw/uVyf+5ub7GJIaUWWmETE5E9uYQ1cwOo03TGiQtePNIfuO
JFWtZDRasfZAlsf0e129VcrmaGXrCe7kd+RFoRboZh/5JzgX5WxPFyMf1IFog5mb
X+uH5qmLDJJbxxdfniFO3DvYrBNejhitMPAS1YUVfxVe+1GJOfT/MSLb2DhYR4Fn
Vsvfz4eo23IRjqlD/+/0J0jbTfi8Sd9AIY06/W04CH5NfsHUMBvNV1Y68zaMU3O0
L1Fg5UW/xagwfJBtM2xE3n4Lqz8SK2zoNTIXRlTkUylgLDVsNI6RaAa+tAalIWYq
DAmJz94C0dj7h2Is0GN4tgsli/G7LHdDNVlYw6/C8ShRieKP/ZEQWV97Hmozbn66
hctLnc8A6Ho2DLC2UyqOSgIxII+iL808bFVwV358kGihcu/nrDbGCeLSSL/svuff
U58f/rI0/RFWG4jnsrRBMk67TZWp5oqopp6FiXV2AuK+pPGd8SubndklycigbI7s
lr/6OG2Lk5aKP3KnMS3M5m+088HxgFBeMUi1WYQHlXMkZdGYKtrcW3zF0T2CGQsd
QprESzLRPuLxzmNDK73f9WeEfCcIYSrbg9GunX3XxsjjD++KHwVjJ/d14YRuUnsZ
SQ7LmXM8zif3hMXPqFhZ/TSBUBBRnm2yZ1PvGeGuoy6SpkvQ3j9YiPd/JOJ0MhMp
Na+8TSAF1KWm/l3+1sKEbGW3tUA6wpUNH5K6tc6meEa03yGofZ7arCrX55jxWAYW
CN6bS5l1eOfRDGY+5n36+ehExftonwtWKdA8Fj0cXqyIPDzTUDA3eaIp86pWEVRQ
oyeNg37ViqhY8SkHt1efvwYukHdrsnfz/LlEiURtSWchS2hdOEaZZ5nuYnJCjbCY
fN4/BRQ3MQW0Yb7Nz5A2nCyu7+PDiak+m1oSpuyQQIgA7a5Aj9jF79Y/igsVklim
lypvCP5ql+p15/1fKWv/5G4Uys07x7Wj6oKnxGcao3HMKzRFkAzKELAsPFcVPJd+
cC0uEfICHpSVzeGJePYAY5CtyAuw3phEUvBFHoqb0TpL+9WovMPWmULQ8r6BlZhv
FrjybUNo6DUBAdYjsSL4lr7ftLOQ5wc6yO/cFsW0cRcymVStHZ1p0YbW/UQo+sBM
I5AS+KyUEsDQZK8SR3SxnpPqb1UZybyE7/mMDgRhKNDPbzAm1JreF4J/Juc8e0jz
kbr9BQH0/VIyXkPeUepI4gPEkQmuid5OmGEHLeemul1gy49+heoQI2HeD0ZMtk4f
OgF6JtCMvUuP1z97b1fmqKAuwS1U9MWNYP5eRkqjEpJLbzT41Rwtw5OtCoWzG3ov
+O1gdiMWaQQASmB8KQfxXdejIVpVmbthJQ5q+aoPt68zyacwhaCVPoBMDmlld0kO
H3NiIMb59HqkdqlCaODdYU68XhWt2DWM80mF4POyW7Rhre6I8ixWeVgMCaiIK2Z8
1jULjwpIeSn9FH2p9IvLoz3MBpZ3mBgn1/zhJbWqShcjtC3OvjQSqmrXLqTdDK9z
8yOt+AoMMPnHjJoYui9J8EvMbwnPFeORpk7SO4w3/F+jUmOb0knzAa7eOtcOcVvz
jLZOsTxVKNwAWdqjsC14S7c2aWz+dxxey/SkfXzWr31nEqfSQcPWRb3DYnR/VxRo
YG/vjZrqTRBgS0xHIkDmkveAldxIfphtZKaJPE3izxWBb4CPOsbwh4s87K3uh/xm
8J1AgzTuCLubi4L9jn1iJKcijf/edYVaqFZuz1Bjq5w66wGty126RjyQOTqfco8c
+KwZZE8ak0NE95xAIuHG1uqiYutjjXEK1NV33iKwY7sKQAMxV3Ne7zRSzt/2CRTx
bVGhxO4PBCK/yqM4pXzuuDfWdS9hMesytdN3dP8NaHe9SIwm9YlHIgXAmXTTYL16
hJ7hHh0Fd15/xQaZaCqSA/J0DXa8INx4f/Qu4N9fwNMGKW4Gev0ycanry4/rc7eD
hYkPbug2LPnXcn9POlCZHNf4egUoUVyEs45TUTEoVsm4GP1wsr7mVPwk4Qd+Mmp5
SwErYBhQFb/CEFkG/1bnI0wZ4uHLzdyRT4GG4M4YCNMq+3y2ndbWWmiU0SmESNfP
0WWEiRBCrCy1scHbAzC66V5IPc+WtsF6JDkocpnNVuGLwOAbfBTv1sRCsXYuotas
QxA4XUPlP64rbcF2OiFf+HH+SABMKnFjcXkfQMmfMs7WObjFS6C6AQqZ+eXlXF8Z
QfTkLnbiBdrBHn01cYFb/ZRsxTiJAtlzYN53DLi/aCzCDkq4XX8jKDE/LuaUx52J
tb+js3kDXT61idpGAetMDlE0Wg6bLdECVKn13klzRXVJn67BmVaaghAvTJz9DFYk
2Axvs5UIGRg+wcLORrUEqHI01+dBzNM635DKhL4YBRfIwg5/PFgK3MGxG0jL8cWy
KN2Zz/H7jwpI1lm8VPdgmrGkL8LG1HM0MiY9p4Hp7mBxq7tI+dPR/NnFJXRPZu6f
/Mc18gIlftW3xiYTBf8l20M7kYtdGk3pGeQ20IorDsc7Y8BaSr30ApOJ8umiU95T
ensoUsQHm4Upq4XIGyCvN0wF3XDhmS5nTjtWh/rqW7re+q3XVq6/MfFFzqz3ho4m
0ZsdK/iykdp7NMPvNrgeyIOgemtMx+ZFtEhc6B+z1HNQXRzjndOgEmDqJLgNsNF1
EdPAAQw8BaHi1CErPqKVDcfaJSZLRQC5AIXLZr6Tln0ygyMk6sJi1A2BJA31QQjm
0A5ZJ/YuPzhDKEnQnmUDohS6o6o4inoOQX5c8O1Tb3RSVkMxPwCi25O4s+5+T0Nb
Rp9ZqkjjDgr/TQCg8u1dk3KX9XgM2XQaoP0AhZK0wSzFAXg3oHpLMZrRLqBwbsT+
24JOCDKRxQ0jvmvq17bq5YcoKQHS0ljZu+bqGpsOq6mc80N9UcQwMF3b9bfH7k4b
mdE81+CjI3CUa2FpwHRxTKmhGPtm5UlDHv2ublJ0gtySX6hAKSw/+SGVMYI0E9nB
Rm1MmtWNksjjqtmEbY3Va6iROTwz5QTyJz6UDo0v+8bN66xLzPtSfXgaCVL2oZOB
1D1xbOaJZ1/PKryPvI+pCkK1onrg0GFvOKgEsffyzf4cDpG6fHDDLpz1ifUUnamh
YNuX7Jv9vg8BBykXPq3djKiQb0jmZwJT5JWJ62t+S4ADPgBweuIVVqzpyQYpd0qh
fCHqqYFZix16unpowrLmJiLnwaMGBf4zjSDWsGCCGxqeK7/vGbqYmIY2f/XyToEs
fHcjV7P/M6T0+vVtJ0u6pOnrIOJIlIBHQgadaIzsnY38SWLA3cfvOuCFn3Qkw8q8
WJiBxy+ak1ZGE1qJTenzpWIeeLHq42dgMFmqo/XTXtyc4d8njyRRxTzgbqasIDCq
oym4kzSappITY2yVc3oSfp+zsYkv9z+X3qiqnUq8W4pCtxet0kXlqA4r87Y8fakN
YKea7V59ZqX39D84ZGmwfGVki9w135G10ZAJqs7vnExnruI/HRBxi3n7Ap7KGoNO
a5y86esibfYgHWmqejHPcCX0V8x/GdbF4y8uLdrd0rYaOInCtEMIGSwiLAtM4v40
UWCcfq1fjKU+4prtbYaCNixzNzdWLoX7bF0fbWI4wfXkwsDqQJgdvK0YK3Ygp/3p
nhuQqjnw9zb6yUgKotexKykrECVpOVAJeDD83bS0WRY3yVdBwyVGXi/xP01IPwZJ
9y3ezEsSZ7AqptSvf+ver33yw/D8y/ghCShj0q9Ote9fVD8pVj5qfhdAsJrWKEmn
Iec20AxjkX3bhgN3O6KcD0HhfVhMkKh1J27zFGub53PIUzQx13TTI6FaHe6g8lNd
xNuqOrhKoqoG+Nf4kWMiF3ROoMQoB6x3K4wQDS0jKpQ1zGGi1mhO9KQw3CsQ6xEr
PClRMhV9uqLB/zwpEFaWl/LPin6IhbTnERGqYfv21Vmk6q0q1rAX6fb/ANl9ZCWS
JOX09DS11Hg6v0YPE6covA+VL08+eKkzMD0Hzw4BxocuRYU/ExwlOob8S/dJ+YHl
I6JbJYHqg+Ki7SjgCni8sposz5WxlpxOPL863gvjUz9UdfdLsnF+HN65ef0t6SdE
TXTLP9wAlAL7OrWq4/32oNPpcctDeYFygfnGeXof3ZUdgzl/Hj2XZZ87V8aqmmSe
ikBhtusksCQA/9BR3vORfMMPcsLz51Shh1eDOKecb3LnFu95og/F+Cvuj/CdYoNL
MUNloC1P9QGxlsFg0oJpkLX6SVY44j8lqKgOqzDmwCBWItLqUYk+Ed+qjx8Ns0/f
lBb+ltnVCs8ZmZNiVfwYF9xiCIiVn7W7x7WISOeCKLuWWC1TsKhsCDioGU5Umttq
5mpTKiEL3ra/WqhomciRI5veLpBwZwa9tig4ey6s1W2KEWRth4U6G24ODnvgHEbD
/qURN99i2ZccQY++dGpVRHDlAVh45EF3fGIuDePiM3oYYENz0ucAyo45D4FRDq/r
/NPn5Ts8ZBEvDzz+Ihw3ttolQ1PE7y5aLxAf0pb6CBaUtHMP6eWB+ZJ2N5o7qAdR
+4d+QVAFLc0Wdke35hmR7A+xRztouBDJ4AIYQM2A0PbqlM/ejrmgeFi76dLMzi5d
QntT7MLTOPzXjRRPvXATbTwPR4zAl7RLdmTOjD95u7RGl2Xf16gWbB1OiLOkvZOA
ML64RnvI+3bArb2Dq5FK2t2HhGgsgixDdMViH8YgCydtnBXs7ayHeAsYekrLm16S
BKy4FdXhrghhiH/vCldtVr0QRQRQTGQz7mUQFwxSc1/shVTOabZt43sBk/00Xa7+
5+30vrXozbZyVQXPMZT6GAzFFcE7IdqTFu4+3Td+mk4XHpUuWoVA0vt9LxJ0ngnD
8NvtQWtJjGfCRvDBXSyd01ucXEdPx1nlieF8+yYRN3/iw/gCj63EIsVvwWIc4K2g
D0fXwdCt9gRd8bXBrrL4aw0jWfwPSvDhxJM1IblByIkcJKQxpHHO2qld0kplDcfX
D13esR+QiqLsXdzxnqOrc2TF9OdZLXWjOfKmLqgIjkxtesEHqYuEzTb7FyMVUa6P
fzThYuNecEpEC1uZ5kURPaWHondbedPAX+vgP81bDNf04Iz6itARIfPH1Wsp+plm
a1773IhOL+HwUnKNyl00uglONGcDjkuqZvkn1En5wqNHGHm5Qmx+hreDsMAhUKFT
GRGlOWyyMD83KYIQeRPGcybMnHL+GebTklJqf/+sumiHBGhjF3oty8QYzi6oWFrX
Cptc9kfO/OmXJlr3pYucfi3MowtrcdHvaIpQWYbpBaW/E7bY/rBgL4BBDklAzVjb
dieIAVpjE8jbR5ObnLBtPU97hc2ToP5jq3eKqo2u85FG4j6m02HZuUBQdznIEWoa
Axr1KW6WzRkdVeO6fjTWQJW3e2QHW8GrHA5F3Kyrud1L1NomzUjA5GhVf0IRSR9u
3ItJLqMjrH51kDcyIlxk4E/YAc9KxGrhvJwiuS2gzu2o5aTrcyI0jIqXsUoM30lv
xMccCF3HfsMatZkSvYmnq/5FErHQ03dExwT139uUBSfBN89t1AJ+ZZM41UZEGacJ
GqOhbVu8tshAcYk07A3fzt7PDc2P6lZ1qv+HNODnTo4Cui3d9IQ4nLZsQB4YS2wb
eFulS2mOV8qXjCE8i/RdB0Hb5R0hD7lwri8NhrTgrvr4Lh0zDG9bTwEJhcOskyw5
ihP6J5qPhEiWkf3GY2Nupb3e1Uez0aL3B1+Bu2DGeemRbNN4Ixz3X1pRdYiKySe2
5R5X2nfiKbWZOhfrSf71sdsuICjqho9/lE3Fd026jEjmI1fdaz6IgHhFGEIguPlp
QZEirEMlrhHbO2HbIFG+XsntrTu8xHnsJHqCv0vBtsFsS+S/4H/2Cm6bQ6/Q1evq
xHbeTNZKamL5DCQObhy3MNmNvtOOMa5hWbH6CsOZwdWv1yZ3tsoOOQJywYEyt67r
uvYMNGpumQtNd8wrCLiyg/U7I7ZIz79Nk76cUXBwrJXlYLnTFJQfyH3gdQpjjHqY
ACod+p2eW83JTHaOu3s0DhWhjixxJIgUVZqz0/pb8EQDDFlJ/TRCcigHApZZYcgb
LkrHN6uoVMfXo6Fa0q7e38fNskRZWEnu2mK9xLf1JYk8kqCi+DpX+Y2LnTov5aI1
1HJdxb7nQ9XlLIw55Yrq/vKgEH3G3J5uzQVQgtbMOs5xk/E1PcpLpDwaRSoNDo3q
ypKLl3LBdwqo7Fv9YoUx9DWN4LEHV4SahBPtv7xRTYCD8RcjK/mq6blRiMaGn/n8
fp9mJK/g0dHzLwDkhiR7mEaRd3ZiF7MAPDzvhp15YRA/F1Lc8c5llOj2AwdgM1mf
Wy3QenugsZBjysqm0zpuDFDZrXhE7E6N4YRATiExxuFpdeyh+mmEaborQ7okS5Kg
YaQQx+0SoWnBML4GgkKjblidQeETgKNyv3TGluvFTtS4hTGijARMtPmmJua6axXq
mrC2xiJI/+4DTapS+wlstumx5mRAa23zaq76v9beSD8zY5eBAruZEMYNSiLjHQdw
HKimw+hTA4yLKYmBWyffWhlF9zrdEARm73sDkxaSpojFW85XyniuCtci5AGPKxRH
Ci6agV5gOqLXDHdqc2Oz0tkZiDzGf7HR1Nd9yjM0ntglnJ4gIxtoQUMsMtg7LtOF
2Akdot3ZGqRfucEBFbhn1QxzDDB9+iP19cQHWOQpe8D/yvc7vz5wfVjsfBlT8R+1
yPfIaXWSY7x3PZcsP4P/Dthj8noi8LdR48fAfEmgJZUOfaDDmqOtcYLndqPYBddH
GeiRWmgMQHVR0b4XpJQVHgQMg6uUkYOBKzdwIsqeuXnD3mVy7NeBMh/OwjX+x4hc
a3kCIkT6K30vuuV0y4wzVgMLqaRaEdhWrS4/LnJU5JmdU+c7kV3e+fXMg36UYeek
CAXfh0IJvf/+XRccGiR3uPQMEukLmTqy39BqEnM0BewQYYy1jeEavCFZ/PHp060O
nUBNBEHeZR5CEyQJCuNJvn7t5tUcCJhxQZ2KBelLTxv/9Jvwe0Wb7s/bFIOmBAsp
nbWjHFV3O1MTcJ9g1as1CVV2scgGeBtfUuNpdQgK+9TKPma/bJnvGyUVFcf5unXC
apCtdevo7eQdylxgGK7mE0OLvz/rBwEAzhmD8QV5tCPtp4xUtx4gtQa8R+j+cIi9
rq7J+r4ohVSZ/s+U1wGUiug4tnkRtMA+57wHUTXpr/6hmaKSZJ7cM6YemzK4eopf
wpmWhqeGqUuvcarwcg+ywb9f41EMp8fW6BrxdX4XQQt87VtqB0JzNNeGhCVaA2Vj
OPVvKv9EV1+giFSrpsBuh+2UELD+fGdIyM3JPl1yPS3HE8Ei+dJHOtrzX9bsHyXB
ytRQc+UMtyhXyPUTa/oiXI6jEAmAfejOJJSIRbLTHTz94BQCi5orJ5HdI6sSkXnS
CeHxoFu0r/+d7ujmyerjEggmt0EexpZsTc23HBhjlRrMIsEm2BRgNv5LYVTgUWN1
P2IAODbsAW0m+msptYQ55NNjqO7ugx60+DK5XVNojB/3y5/OuAySdwKnzb+rvVYm
nDfk7qa6VrZkn/xhj63TOEIrjtSSASqCrhj7SLZPtQcuyxwIK4D59cQJh9NQrENz
LujaaPjK5iT8Qw6wSmr7B7jWyljo8Wx5fENcvh/vXA2UOEGgF0ZQmyET8HQRefL7
HHzdpH7IPxU8IYg+4rspmq1TVTt0FquzM8Kfw8zMGCB9eTiGkIOpSc1nysrnuwdH
1jnrZCBYW1MqfDnKZ6/+pxPnsoFubqC0H05xGSQFy0fXGOdeo+VlS62l8vBedXps
8OvC+zMf55NyuF2S92bOjakYCInRh1GuZnXIGuDeQwnp9U8VIUy8NdXDy8irOzEV
0WGU7SI10oR3yYBzR/CsM54Eli0GSAfNgULEslfk0YKBoK+sg1bnXybd6siiooir
XF5b307P3EjETlwK8G/lbIN5KTlkwQyHZlMaCybrBOc2mBhzUUYFroAG5Dm5uaqf
NfN9cs7YNcoVnlYCN640zBabzShhpx7gmCTn9rTjmN+3C2TR46w2t0ztL9yiDdsX
FDTBYl1ZDe7L9ltxZK4BI0tQ3+z8lJDm3jjd4WstfD5RnSrBpUGLOnVTO3ZqZoEB
uVk6QOesufh6vHkndeDFUKd/mdSDuA3C42elNAVL70kmNKI60VrGVG2zCQEphIzC
zL2Q/HHwdNoT+skGraZ1u1E9qK0zuPMXDoSXWlArIrzZS8iDFPsx9CZmybdOV48G
BmTns7lu8sBsQszUMCAIg8DFyYVRMm4c/0kT8FfgdkRl/CEiE9q4bVeQJ8flUHT4
uC3XcudyiHdWl/+j1KxPIN3G4gveZrFNhzD86ze1vYpz4cpTd69tzz4mrsCKljjA
F9dz84RY//DC+cnDbRu8xyKIXNqrKiZJ3asXqtX9Wz6PDlV2ih8epnCCwsc4Q5h3
5u8nMQ0qDTMXIe89yUw5WFMqHJeHgNjWtKGZOzyeLBxMqWH342SCaRCAOZWXZDTm
4YEtj0BR00F4/NyFEhXxh2OwzkWacI7unOFLr45kfgKHvp5nD7SWR5oK2IfJLX97
oJfhP+1ZMav8H6s5j8Io2ZnutaJq1wQ372+AnHhQ9JYYucZuPSTMg+kuZhhjTjxE
FxIpfZPYJMEo5Rt1Idq7CpfMSXXvdv2WlzabEf4m+n6ecnqagzjf+PelZejZiJ0r
YZBuEcb+lBso5VerXXpgULkqzktN9aFMu3LIP2MZoZn9+V3k8acUy9c5Y+SxJw01
7064jb2hh0gRo9RJWAlEgV3NLXKlgi+1Udk229cEa/vQgDLBtjAYTzHxeOFm6nvy
CmZrkxhOA5Usc3TGEctBtflXlb3LTcLHMGhqEKk7r+JnsW/PtfhoMcJmCncLZoAB
u40O09eYFNVdm7+ti5PIs2zvjcfWG2PGQ+8e7oroHpd85xOOQcfQANADDFisAm9j
H0bMAcNcgMlwSmCCxi5hA06+NZ8BrCOUatHrIFHZWMeP/27Tg7adYh9ImvHCtEec
YBWb0Ag7fPIdu9f0qEqcar8sfmWGJFA2TdBy6t3x6q2PhKeaPC1iyDvTxACJeXwh
w3r3Rw/19beDXNUObhL1G8kxn22bhDIPQyokd4atceGeCl84qL0ddhG6jQyCr/sN
4Iy+9uvz+VtPYdnWa1Dssu74Ty9fM3KeDAd4HRJkZAXQTUCZUA1kjYSlKxTCA76G
sMLqyP8TPrH1q5GHa9nzBuNp2/xwMukCU/qnEHI/MQ1RDGLlZwqQI1h5slQ4qggq
wK9GdkWO1m5plPVieqqXaMFtuZ19i4l4hLsI7Z3ZravJaXLvAWHFReujkab0/TVz
zynHwi5LRj0DQnMVxIJLAz+kM+coW5NAPOyOt4J3kEy0yMVo0TCcNNIeNsj6fHVs
u2h1to0Lw7tS9UvR5OYcypQDnWXDvU43D1tza4OqpLIEC7LLHxZh8XlzoKoKdDc0
xdfqLP9QipDviyJb9zx/szEA/yPUm2S6WG2XOq/gfwMsKwmDfOjzzZfs/Rb21AES
zQqV6005aqK7IC9p+C1HKrPPduK60nWILeDw3i8lMeFqg4fg9RbfM1LNN2cCux2j
jxJZbtrv1Chxc4uCZA7LnxgX298D9qd8H0gRafdyh1eZVMJ23c4FnmJk/G7DwLT2
qWFPARUuPKmMFI3ptwYGXwdLW2av9fXAsZezZ+hvjNu1wuNdq9LxdFN/t6dX7FG5
/eTWux+izG2rMJn8c3Ig2SsSZIrbkXzTyaUM2Nc6Y6AAN6WwogEFkeKdW48b65Bt
1E4Xj5nmvPXqNeKr2jbyoJWcxyIlDgtOvEwzVx/MAhwQRfsAjbKYSlbK7JfLgI7D
oE9IwFglkLFKad9KInLQDMi2nnoLCc0ubItDyNXiYmilxdWkhyaMHfiB05CxCxxv
vHHT7pww6JIG04qkuo2M8m0HoEiwrQ4Js9iJ3HNeNuRClI4HQAeSYbVrHQaqYQRv
JvQNKcILuj/GSb9TsXsnw1zRrN2AHyc6Q5LAl+k2Lpi4bdyidS62sFQQ1mOWhw5V
lZgUvp0FCBMoY5sFjeamsZmanhb6Yg0D7sDY7sa/fIRKe7AirQeqnfrlkmlhfSHv
sZvoZ/tA4G+W6F65XQwylpEPvHkAW1XnIGHFyYwu5oxNYP6dTDShLJTaBbj2f3B2
81AaAb3zF3beiic4Tp5w9DJnngtNOg1FrPdlB/8Gz5ZWyBfa9LN+mVPQdinYwJ9I
6ohxVsH5VdIpXS2Mw8zxE0m8FjOQvkYUrPgHbIJ2874e3qCYK9Mo4/IMvmlLOhs+
mBUYm2bKlfdztF5wZdFQNS7HTc3OVq2E5TXYgEEDZ8AkGZ5e2bsDODxL1SzAuUrL
Xlmhq113Kn4KH4C3sxkcrxjfD+klIQkQwpwo9TsFRGC3AKi1wR6aaMgbIg1KUT7x
zJ78HbJvULe4qxspaswz7Nxpy+JNmRGYjGtoIRugrbvzKPbHbL6+cqFGk7TO6fJQ
foNNiKxEcrHVpvvCiB2GlUtFyoRDaGPPFu9QdVfCIQ+a0RtXL9i7g6r0sYW8cv9t
z/20QQ+r3p8QWo+OU53HorMoNDfAzt1Uhuhj5tNI44Wc+J8gp+FnErdNVcmH1sM8
j8pd7HXtHufl4mSX3Z2OV3bbgcTkUNwEyiCAJ9gOaPq5DxwDevkTybEej/2QBlFH
u9GjwqIpTJFV9dtES1p+Y/5xdjmtyYc2bDcta6j6Bso9k3R4oAsfjcMyJqEdIC0p
rrmrr2On14lK57eYkRaoxzYw/XQ5gEBCZiWaDYbx+z9MzAdlNJ1ySdrIiFmKCpaH
HKtXvcN+h+TkWCsabavV9bjdgxg6x4dSuy4VpM9rTzxlWfS7lD94ueYTnsYbFuYk
1dyIqCsVOkc6fnWyEsRbvPWfvNhtko93BImKk0mwW4pDB3C9BnVoDUhjfRUYsb8J
0yzLbnoPUMHsJbT5wIvCBXKjdPMCBhHG25+jykHDQ4puzzBNmW/Lall7vfWZlJFa
/EzPDgZTBVAsqkSIKu/fll4iiOTUzpDj02Q2Bs6zJwwDDFbVihQck5K658LG2ZJm
MLdwWut/UWhcYUVSbu97oo9XIsTLaGjmPsftb34ebwdIXbt4ykdSnhtbLQ5F+Ze1
jbWp2zLYFvXdRN09Q16A7qtRQnm2CmXWZWcC3N+PBNiVzhyySAEpFYGYvJHqLl44
wz/HYSFLlxRn7aWiI+olsOLOA2rk5Bu2w47GB/QMENedvyJhyzvTw+i/3rO5vncd
6a99QJCIy59Ii4MoJeYRmUHwQF0m7gcg15py/smUADFhvVcr6eHO4Q14qRNS0n/q
f6i38gbzsfocdcs3yks+1L+TuvVputMsqASua843UOVCMmqvbUj7rUOEnPYQxnp4
7CpvG9P/HRKb7R/fDoM9AuRs3jOsnfpgUpiGxXnM+gj0WTW8ZfiOwL9VyX/DCyav
RLBbBXr8s0Zt5HY5btN7yj3p6iJ9ue7pnia0EEUimDNTYXOX3FE9pmO3AzAi7dp8
0n9KUGKIwcAqGBhdC45KpgEyDtzYSWgA9E7p22fPHQfEUHQrsBKnqKLuL5IxYPU6
BczQ+allTCZNrPF/8k9bF9MN4AM1romTXL8cIftIK1h4GogFpEwTlLKNf34wISWS
so2atDoJFaRR4204EmLiNqkdRqAN+OrWHMayg7kUTTPf7klz8GdDaPtAPafbZj2I
9HbchxBeca//XwZm6Ygmk1mPYXckSmVljkjjkJZQqY6OwQtyuCT823lgyE9PTQT+
src0X04h78bhiR8xCL1pdpYnIAdiYxdLYQ8ZY36spZTJDhpkBlPnKzaUyl8g5SFY
fpXppDhlCNGTUjJKY6GHefBvjEbw72dXCDn5UvLobqpCdBlL8xgiyk/HQpakbNcv
KLDMK6n+AgEHmy3sjnd5omcKjI/IoJg5xXKnVPm3oOaalJHMui3MgS5+2CFD9b5y
Yg63ii+Ea4LL27CeKUqpop8jYjPyMPZ9xXfnm0165YiWnDfeHgVA81zYoGLaMg0I
SdVdsajBRxAxoFhfZe/XDdB4n/2ONGa5qfylRT9LzlGRdA05Afr2Qn8aTBFHcLVa
nUXUOjqZvEgKtq7ipqcSISfXdRWRLTzKKW96cqMZBAadBvDRCkBAYzShcutSCUZf
y7R9zryIgR5mjIqFutzqoBTwrMeYHJPq4WHgrKc1rxCAbwYTjH+DP4M7fJP8kngQ
uvLIN/ByaknbH480XFvhrDUluqEuqMGKS7LOF9+VVdEnyC04uOf5wIdGCI6988Py
sFCktVJjQ2eFjmnfnuzbk3iUiH6EGa4PRzKxwx5P5eAk6S8a3Dpl/q2OceVLTxPa
2y7PieAb82ilf2XGwppd68GaPhJK17GAbJeO6lVsEfITZkuPuZIGY/Cd6hVyqrCS
cgaDsVw77ewIZrAvdKxzE5PpOH8RsuqIRIzVXDKbuw/96hhzS6J1x9AvTW/7ZIHw
EcpeoCS633Y6EInUyb5xz4sFRmxPCiwBtGu/YAfmhmA0AsDDe2yt3aHevRqzZ/2q
L6U3e5ptU3zCTJe/qANYKvQcV4AiLIhNXQlHsYL5sZ6uVkBr7SYMu6C3zcX1Ew9a
vrW7oPnuAydt79TObVlzwUO7jY4Z0H/nzN7kVrw8SgZyLqS1Cn+6gggGvTRbtk19
4QEAwZ7t/9VHgiyfDs8ukr7m5H7lG7m08rH/MyySwUvwjS6BsAPiZ03KVAoBSWbq
FhjRknm1C4F6qaqLSs7R0NEAT7aQlZ+pV966dtqCD0BdJlFWKxcFMbw/ksXtkIxW
1xtoVRV1TNNNwtyn2Lw0XJ8vyUSB2vv7mMKLDMJMpxHIcjEMbFF+SjyunVcMYBqf
+4vsJizYf7GdvknlMzBdsSPa0zXrOYwa361c/SmfZWXS/clUmPxUABXQoueFfOTJ
TQpinEDOlso0761IqBp5Mz0FNAAWlMYlskBk6/WnSubsHaRVfr7W0Wwzzjf2eOPw
8GTq9mVCLsDNwC4w82URz7R7+CPEjOLxt4jb+SxRtLvRGoGEk1OaKSwIZQFftUWk
NeQ0yBXqwCAX9pzZmpJgYnF6NCiGQJFizRVJiXAVCPDM+4GupFbnZXR7vZQcVAJP
QuW+xMJaFTZrG6ggiPY/bBzHgxeigofV+Q0RIoQaTfctf55osrmUn+RBNiT3xFf+
OvkU3VoaGSNDwtwLF6nHoqYFQ/igK6fHGn6fO98xFelX88tVAgQfEGf0AycO/mGL
1bMMscHy/lK9bU1z1JaIHGPwHCenl5adRpMo2GDmVYSwl4p1M7jG/6VJQ/pc/K05
z3fmOCArCZJlezPBXabbe7lzujshidYQNYX36E7xy8QnIvPLyAImpJf3D7d4OuDy
c8HisSHsvHezLXop6IyYR5XsQc8MtktaYimoFxXapkJXaqABfz6WZM40bTwOTUDk
zsfUcysx0mbJ7QGtm5LOYRG4Sd2s7aCt5BGGyrBDXWjxKrE1LHzHQyIWD1O2xv+S
aU9oOe4HG+9PCdT4bIaN/PtX6YaMaHYNGdy5VU8U1LAEle3tR7iIDehKy8Y35HCA
O1i2cguQYEP7xr4nG6h4Rf66IlEXF4A6MdqCCSk8LLCG+FO/mweezM30aXxGcgFY
uUv9DZKPBpMNdttokl/AZHIXGXKtG415DDo86oxNoKUuUKnaPKzi75B/g5PyJ4me
574Dy1pHCz2UlZ3styc+UdS/rhtshbJQVI8hGLXKWD0/yajdznQ7l8Zapi8Z+pGH
5iC97fFKMkY9kYJadkYMScCCck5Umh1L9jdfIu+s8JmNhgq9+6swE9zLRE0fTqtK
J3SfGNK+bvxHuhGTID4hoGge0QYfUJkOXr+yMhJI+Tk6mrUiDYKc/oY0w/ilayEZ
MyHQx3u3SHz/+/lN2E1cG8i3E3N3JPxyJ+G70rtPoUloB/YUcGg//fGDUSHHe9yt
qMqKFeeqzsGZIHDJJWFSw3DB7lEY7FXRZH+cTr5jQ9GEk2UbV+SasoBbpaEvjKLp
TNVK2y1L2N10NWyRN+CAqGIdiahLhVolfpuNDXv3+jkfbsMD6i+Cvn6iXD8yVkSk
XUL7NNTn0dt5tXcrtc0o8xbdNVyYuTkq0W45BOp6FLZGblV9bsK245+CHkNH7Y0R
XEGob9NFjHtWvahbid00POH7UOkskyh21t/p2GwOvHvKmgUN0yfFhEQfULfcKDiU
6kn+DlzmCN96GFOkFkRksG6dC/IWFZVDUrYmyK+YyKER7yd5L55WnSh3KJHfo3wt
gCqUKWJgAUV+5XyFJJGtbP4jgma4mrQdrR96ZF1sXqRkkNvyM7c4EYxedR9cxuKg
Rg45GlUp0J4G2ouIgJoHxuIrQKXF9Jl4VIQBtRNHzpjSB7MWaU93sGLLdgLcvnP5
lpmrgrNQPJphVfS+c1xSj2zmAc5INWMAOBSdMQjadQLR59Z86sAPHDk7WZDfHLXO
dI65w0CYJbxxAeoKI4vtjWueHiXfnDnX91YxmJt2AeFigG3H4a2v1jR8on/vSMPh
TDMvo1bXwfv2OvJU/L0LcF0Lxete3Np9JvaAy4qFiuXWGh7QKOpr3bpFV3aMs2KQ
/DXBgD+7ZcHKeWj+ZiOhwg9sADxzCVwI9/TDNloHLxQZbBqEmBvRrX7p29lu82Vs
ssW/VeIZuhEgcrEV69CcMq5O3DwjbyJWo5vrvGxOQvBAf0M+dgNkTTOGfhachLjM
13yeFpj8CQ48SEvGOyNvhvQOcAsrbE4WPvXcCyu/BAjTdktjiuMd+o7Z9b/ygo0J
6Wqh/fMHi4OqJnI71cbYFhYUoWpWbDLAhh4Ghb6aWRtTymG68zuHqYApS+Gk6cIs
aQ52n9DL73Gf5eEEjLuRLqhMDE18effEnwBRWWUqmH6IHG5PZ74e7SS9ZGulo3Sf
jw2tPWebt5xVLG7UAOMoIGCy8GpHTxhzzTVDzAo17LJ39zQ5SZ8n/MbnivkRCaRe
RG16xfVgHh1mdNozoC8zi7wNA3pm0NllVtcUbE/Sgqtke4b21ZBBlMn8BmdAfbYW
h7qmwkXtgwABnPAd+yXQjXs7+rOLhvEkUQlBvqRt9OHgVn8P9ZzTkhQ9Oy7Zv3Rv
8VuGfJdrQ9z+GTPa0XriTMdaDXfD883ToQnOm2v1IB1NNy+POWi3Ry5rUoMj2Eo1
QBq47bKjaFugok/JgTGcFJ2bxKwxmbXSL/tppCSlkcYUVYxnI6oKX/WCSAq6S1fJ
fbuRU0eDExCiLdkXgGYFWUkIAhkvPy9+G0pY9UiMwvB2rtAvc+ZpjoTY60oekQUT
Ms3nbvRjja7VCyWA+Sd0pjIRf+KmkVENxU6rLaqiEEOGg29IzNG+/zLx9t4wtDyl
2JBpxIY8NIMsKVnG6ri6tvjc3PC+iHTBdb08HOHm4TqlQ2ZrM9tMbeZTqy5yrjt2
B2CUBfmLZCoDSpT6qC3pzajHFNvpJN/Ovd9wRft4pY7/zDz1SNCWrx4iM/NkVIyD
1m+utoqCRtAbrCRYRqrx2Lhzd9uEAK+PEPK+BLJQAVZpmFdHybG48rK/Acguy+Il
aEJe0FZuYMrCuDuglyQ7iLke6uVDgMEPRAGLeaa5LAwvEZEKrtMO7zHXzlbrwg59
6P0DUwL1q0JXW4lK4iqrQEhGl3RURXyfu1dL2s6l84Zdt+znK5XJqo1GDGXe4n52
4+AJCeHSLxir1rY6IjSSnyFu6U2MMzCYyRPKQNBkt/Lzl82FK5S7xD01szWqyEO7
2rqu7YqlNgcm8AhOeCptSVIsOrB9egsatzIh6Q/REEmFdeVgbapeI1/8xZOkVK9w
Z/UzRj4ueA1GWFJzmHM6IJiJD3eo0bTglsWJEc9mGHk2ssLm9t867gOv5vf/5PYO
BvHskx6VBvwR+B2AkqypvL6dFJaHrNJVryZHaQj3hE0dPyoyJ4zgtpi53krp6dTU
14tBfMEOFJH0tLW1sPEQ/Vou1Ds1VqhCQzNZ2YttqScRnl1RBu/HOGHX982W5lWf
mlIIZpn+4KAiZJOiKiQPl3J33rv3ONutHeqqtsgtsOsQO6t51u8wADXKG0qtu74E
t75bNOzHQ2UQsYBCspqbykc0r1Z2kv1+WCqCxDDWSC2W8VNHieECjzCfYAKOKmkM
ONeubsv+uwQlGsAoyFL+Si/gGxCTwPIjxJa4pCXlmLiVdkikY8ZOumcciAXc2boV
hQCTXKMIMaD6wYWtX2kXVxCWELP8KOyMK6sQCtiN6u5tye3l0GhbxGPkYF54iAcY
vvIRlzaLxjigiiiHc5OSrMHNGCd0q06vblM7dyURTfc/0GMhqzn+HcBKDoVwYQOe
Ll0DvDFOSenwXbHnmFZHwgICYxuy8MSYr/z3hPP7zZtQGjKKukGtTJVFDJQwUgCA
4XATP2FRlSJ1HwYntE3u9v1Hm0cmhuglykBj36iNis6iMvLqcNS/FqeU3GdmuEAE
cC8Mq8Mf7hS5MUmBNkoncEeUcXkQkG9rX3j7d/YNyZwtXvc9uH2Y+7Iqyuj9ASOV
gClRARJsV6T7JL8SB/dM+UA/qYw8E4IOI+yBZVxTNzf+KBpHZhB1F4S8ljEYqu8J
n0qml6fvTR0DkhT5UDMDkHPEpjP94BwHh4aIh4GgQMQylwfl2B1BniM9iF9IJzuI
PJAR4/vdgg4NODXsJGEvls3iJ9VPYfT2e4kFeOfgpp2E932VasAjHxC7S+NIatab
2q4BUmLrUFeke6Nlhi9nCQqiEXGKVzAbcTzT1slB4hH7ZORLPdvFZFQwGcRvPCca
XBYnr9xtyxPC9PaLf6M3uXLrRqLL4NOmasNYrlsfGA+X2PGMh2dUx41LHQgsa4+x
zs65HhJcydAzWLV2n1jAuqeT1nAn00vk2AcZLJmWUb/CSitIv8NHkhPdoP/QIhdL
7FaNWfx9xbCizJH9lvnwE6Vok+4/W04hFgbzc+BAFPBv7MvTkNsOOyRD1PdaOBE9
eVtbPGgukaBXlNA87iass3wtMt1DPaVyZKAuuVn289q1+UYFy6nzQnfY1vO4c6KO
3vlLCfkXiYm1Vv4tApQKRRaqfK3rXWCIowQxOFk1WD/LLacjJQpRfUPAvDWtXdPh
wBKc2uMOzqmRtaPDr9ESIa/hrU7czspB1jCDmMts71Zmuevhnf/TUeaNanSxt5Ht
/ftV7QiiBl6bdNRrNqzsEQR52JiYDmxMUvCiDjF6Hi/O9u9fSp2AIazmr38zWrgZ
CNaBsjRrSb7fxF7YodFVzp/LAx6qe/g9yiX2LLMMD0MtZh7f4HMsNaiETleMJxTL
UeHTF0w/4Mgwscsylcg7gZBIwDU4baVx4rIm2FTI3/IvnhFGPnN2WkJV9v0Ihuch
kboQtW6zP1J5ZUk0l2BH8fn3dqzU6L5vfcQzj4UD3b0n1PfYifyO2H+FCqLvK5RW
q2BwA3EVV1Emd1IV4SpohryRvqwuWNVla3nvdu/kxrSCdPZ9lzttaCklpWrYCGgi
Bin2lsr01jPUEAxFCvV+ztgO6dP0CqN4JjjO16qQq2SARIPp6Bks/B0ssssRslyh
aEwk7JmlRWLzJ4wRk9hcBz8GUPdPX1baeeuuJFGSzv2FjX6xdyzubt6HP/wBo0cE
FEQyJU1PRzy92uZwR9/NMNhu4sDsm/YrYrjpax0751CZU6g4AplfL6L0oWsUXz/a
xZAv2hlH2TycWkUaRHAAbVrGySNcJoYyQkJspktw45Wvpqd7uk9EiWLDcD1aqn23
zrQfHS7Z57Kpmj06RNtDvVdzejJ0gRzZNpPb7SffdMNbsRzsYUTYJEagnU87KkRu
qaSrvBfYGGsE//WOvHb8x3PBME5ko2I/+VDlpBcpIWuG4HVFGffIEnUiru49gLe6
bdFdBKJ5DBTUEr8yL6K9F1E0Pamhs/dWHkR9WG68N0eQx/YbsCZXMlZj0IxGRHW/
9fHxB9NLF03xa/idVI2OuxmFMmj9xYXck6ie2IqXcLuouOaJwiznFNkxGQOOPpvX
5Sv4kfcoJ2K/g2SODd0c7aYFFW4rDCnkkwDcz/+wEgq078FrH2j2XO5x2MCNzymg
lK4HobglF3f89BmA13i/H8wez2e1/9V1Ru1SNwvLV/Lbivaidye31BdP6FivjJiv
C9jJbh7VKZHp2xIV6AGUh8cCm8U9CBho3I1j1vs/P/Nm3nxoV0pTcLBm9FT8xp/3
mWb8x78FnEoz6zMH5WMwrOFmB6iTA0+RhnuD4LdIpu0anLqOK8UtC3Mkf7T8Utpl
kqnruotzy8AoS+itLBFnz+VwVOHKkfSMLfBzdEIVDZMRuVs9Oty5O+IoDPxCrE3l
bVbFbD8RpZefs7XxX7FglWuYufdK1W+9WexrHBYN3yNhMxD2hXHsLVZbzkA0amlc
r7W3JrpNlVyz6+DTgocpis5duoeKYWx0chAKXhygwy/pnnGiIIcnHqiIVCYEUxOj
BNHwn3277iCp3uML8zguqgNxs3pOoUsk6Wx984QVhxkJjVIzZ+uAHg/7+7v14pKT
4RcAjJNZfFM4iM7+aUgDH4d6i6/7vZ9LvcUP3mIFSD6GW9awUpKwpzpgHF/rRaKp
c1sChGAbzqUbpI51dbl7tw/9guclnELH5SidwoZiHq7v9UGtE4MT//TrMpCoPEvj
kwt+tpmVrKr84MA51kO+EHLV1lm1YhkUEVb0JLRXkVCZ14uY0GqwuHhoBDSMsJEE
28Cc8hndhqDRPI50X1s6rsty+hSIgbuwmAqi9W84nnuVffWgDts4KsGKfept54Zx
ivX/gxHYk2XaNlcLYPg7muGz3cGn9EEslupiiYIkXIh8TGV0FlenSz+1bTpp8vnH
IG1FV6I49x0w7buDfLREuiH8qr8nl2TRw/biqfQEbKl7T5h2/+cUIbkMdtjoqa79
dkXKge8AuV+olejRSfEBfVPOsGp0MZzm4L8DGi3xkrjq2JR3/JRUz5UCus41zFpr
oA6goUabgS+2aBEDEDnehbGPf4hkKCBidbUZQMhplrNlNY947ygehCc5K1OUoorz
OtrCYOwz3R5Fo7hoTydSnlbNAThoTVslAyJrULVls+jtb3WbBbUJtwPfK5zyw0DD
7u6ALB4eCRN+ezXWYD71SqOUUFrEB59eEgqBFtV+0hkIl/zxEAQzUKGdUaDabfyT
5rBBJrSeamnR5uiD0/pDv7w2PWHF1iOiAtFUbfrGd/dTUoSRC8eg2UrDEKGmO9hy
fNn4jJAQ3RJ2RzAoKM8Btq/M+XWxeJAdFcZKQyOhdG0Hn/5sSZRzdfo1PzVtsS5w
hLhJxxZYXD+Fwz6oDeR4kcAzv2Ob76JdF6zneFUANZnIE37/M1bNXx74B81jX5Az
87wC0meEKFYAoOGaTAaGf4zzz507D0IzK3GHQbp6Itlcoa2EO1MqwlwnfNWo+rN1
CeTner9rHmoG/WploNbUrTmsgsJXdJXkU95P4PmL1npORI55CTLrQ8xwRtXvPMxw
ZHNb22fA4ByhuvnEbr6gFIJoLSW+/ZRBCikpGCLzfE1Is9fkw1SlNR5f9xzh1JSy
64nsFi7pd0gJ4I4sUuoialtJYlgh613pTiU0inbXHlru9k6IP9q0bzqnMXuiPUWf
7cFOggVK8nll5RZjzPYryW369HBU6OfcKz+Njow2XwVMalYRDmDqHM3WRZ8xvLg2
N/8Qjuk1qUAUntcsFCskFrnIPHG9aosu8Ol31E5jwoIJ3pdXkFPKqlAbMPAMeKKb
zOzMK8lUzEHs/v4MEHNC5vwx24ocRZTZfggmqR/5TB3QdoF/tHe24Dj7sznO3qlz
7LDtAVhRLiUGTGF3NqdZsh6+4zYQxZFdaWf+oX+A+/4YOhqz+jVStcKbDg+pfkO2
VN47Znidpx8wXNZ/7N7Ois0bOPCpWA//6udPe8rLXUamlUxsWODf+Eq+si9tAX9z
Xab7z9FKsiK5krM7wYnht5zNY+1zctixFyn6SazKpKgA3PVhq/bXfhYQl17FHnNq
R6GmSqmqw/gT8PQ173Tp6ST/LVfuiN1FwHpH/oWeAteKFN2zIpHev/r2phvtAxKs
Dl2i28dbNSwXBP3nNMVlW3lGfTeA/UL579Z2IxsocnP0kxLFUU5+RXDVFBU5UOng
izB3lXBcSojesYD1W9wp2BEJc1kGcg1k2CBV8KGCcGB0WXuBdF1VgJquhwMW0t75
viv3wy2rHTTDplI6cZgPPlJg79kGf8keUjkxMCCcsr1oSAZczNKY5VUx2o6idTEN
SWQYFX45ooy6modknix4nMr2Nsg3a20uRNZjXwB7PTmUdV1ydrqtHus55DSC/gcq
yWO5dbyDAh8RS2x3iXxHSxLx895EmVNgy0QWjzNobA/qp2xocrsCKfcCMgs9a55o
DhW5sPrFsMh11o5bAZYBtZpszJZWIVuyIS9bsiJkX0yvhlUpKebnR9kSuEXe2F6c
WBiuvrPf5gARd0O6ezOI5d6qGjdHiKN8RlMK+LXDWtHp3B6nLuG8zhKWxLDLztd0
jAoQ82AANUrPgWRkWT5cBh1VvQo01ZPke3gVIJtG+XXNai7JM49e3xF4UtJMk4hT
evKHLD052SK5HGLy2mN2Op/DhAid1k5UTXAozMrINQVLxbiK/jx6XkupOEv2dJik
yJKftNq05jyVGAa6WgY9MVeoinN8WAkw8ZEa+ZYcoSzWDV15aBdZ//V9bm4HWjdV
CUrrBX4L0UMgiyZUDlOBDz5mLXPeuXnI8JkMk+pZfextwleUrouwB3MLzNLI32a0
rDoHiJUmmEjM5wiJ+QFGYcTGZAGwBm6HCh1fXuIzGmfwgpQa4zsc7kbkC/gmod9G
NbX0q321gbxqj+cXySwkcvazX1izvBWjm6XZ20Y/SF5H9j+zzHkltD///KeqGKeS
7uSGgMK26zvU63CJsSxN5X2ws87BxA9fdJL8Cnkx+mKtQhIAFcLuFDSuwxnsMr1v
wvT6GlLFWsoptzawlAwiQc9GLM6433lZcaN/qwj62GJoW0AGcamlOd4uQdFIEaO0
r0Npc8M084Wge9G/9zaYQfw+n5lbbYObEJ7ETIoBoipi5JEau29NcO1fkysvHEBd
0OHBPgd3PWyC6/dyYgj/8NLk68j8aSN71iLn3PkEPMynbtWO1eQ2eCCJEY6pFWkU
yEAB5+s3Csny0RPaKB85tHtVfoKLy50L20j7HLL6annNw2hhakDmU1sm5a1QtNxd
safd8VoG24PexYV5+v6KzmMen2+GOWQWV4dS/VeFaVIulrGzJAn3UhVcmYS8wGif
RPM4r16oqT+iYcASLOoe0ycef72IqtUP36uvdpms4A3OShIPXf00sMMONNvr0iV1
9aP7hi9aTmhFPR1h378oHkpxMYFTNnEOJLJBZz0+/izaUYa8prNIEXEn1XJ7PCCh
Ih+CNWfsIrYH9ud/3yf1mLiGdBPdNA7oM8LtApVN+Uv1AE9ojj9JlCAsFUGq6UHJ
oNNVmyNlaIggIB3a46RG7ZFFPahgc6QK9UgrzOv6Du2RZzPai0ZAxycsSadpgwhS
x0fmkVsejaGW0AezSU4XdfkBNaSHo0RkEgZ3cOZ3PSiI3xcLdL+c3lzQsTQFr6i3
G5phowkusXJudqiPU9wMTD6ZNAFwcDZmwKwmthR5/wRJJbP1R3pTOM2g3PhI+H2U
cPkdB5jWy+XwKwWb3xAv+QIYYNvaEJn/2ORhjeRiiKxy/gh9sDpkB6J4K9YZRQeu
3Itdx3Op9wyCD3SRIq9wt8WcvF+YpTWvjo+4rlxIqmiwMEK7j40NfRDfNK5Ly6DL
UY+YaP0Zz0/doS0DJG61o8OIROBMejvk9PCMUSaGwWgVYM2q9jTVNw1TF6klma18
GpQI94ddH1WqYggtEyP3KvxzLnZDver7wrp2hsryFyF6aziQ58vJdiyUy5qcz+M2
rnPmL3pzxyL05P/63s79qTfC2Zi+CCgYdiXeKd1ojlbOWhbHczTQ5xGEdOC54ifC
ltCO20GtIcxHv7RlUTRwj/gtFjjGU5Aw3+au/RyQNYrTD6e+OQssM/FjjNls8F1V
/CjVj0rJelP9edtTNXwAKMzyyCPPQirZbWSzY98Ty3rx4pjgYGaSfEoLkaOD7WzW
BHOvrojsumfCdSRjQ+Gb9SdoezieRIIrC2B/jHp2A7iH8LvwnCTigE2EzSw6JaSr
y9lgFlwMWU2rqYWF0RLHBU5+jlFWT723yfJ6Duz+UzSJH1MLO396yh2hsL+LpPz6
S/v99rC+t0qnAF+5xMLZ8MH7jfTurhJm0Fc6ZjENfmiBxC6Tm6XBjFNDdspHn3rj
TDjWlr1MaxepFE5rDEpzbipb56NU3Jd6GwHgHp8HosTeIrmiS7kLU24VFRK0yuSx
5UC6njEr26xdJYITquG1IiTOL/N4blnsool+cMLlVU7yLx2lKAppSbpXrwa1eunJ
fhkm9gbKWO8WP7jerMbThUr0ar1DybHAu1oqfk75pyg0xKquP/haAA5TpNZRomAW
AXnZkBCoqnO3H1s4LSujrDssfieOn4nrU7U/QdLCXttch/olu/+mExuCwn/4r/AW
SmpfxrGAN4bS0Ngiqeq1a1F7rYnjBGthP0fOieTTXhrZmB3Xq28bbi9hSPQfgCyE
IeGgssMDY7sGuec6376OhiMtJCSUc89MpH9I+qzGKSGenAfhysGCo7OoDE4oDsh6
WOhFfvCc+YvnMdVDx+6xgDoXQTPoIuPnkTr6RiYgFFiv/02uNjQLRZmI1B/szqVr
5CWETShldtLrziLS7V7N32Eos6v+JorfUIMvY+8uBQCG1Oiti+/GpnJEHltGrv0A
MBFbaUEF9HanRb0UwMm1FZgKqo0ICnKsSLEv4gCHGL3HwE25EXOPdWm7zvBztbuc
StGGL3hgzPsHn3KhsQCITlCshPXmQaLqTMWfaBngBqBMiJKjMUgDzn53W7LuBRXK
TwsCaxsJyxN4xm0o18crn5FcG9f+6gNN+fj1hYDxFWA+3fd7ZuBxgU9PN8eLTduE
/qTqcS3xv9txk8zod8C24wogxOsj2dXN+jGnwZisgWyoLbJoq3J5mD6QtP2w6I4w
4WJFjYz6oa323XmJxHiPfCzStiSGp1hBY5Z5lQDQ+CMfJ5zoVscXMF54ezn87c42
JJyJFLKuYmS1ozlyujlTSiyZVEwygo8HACfu9Qfi1zuszg43bth79ZLHlGVBFJ/W
ICE5BXYvW+RL1qfyzqgbW7VeetNt7J2O6wbjckZ9GL7KU/gWcwwyn+HWuHxXsH7e
S1SW/E0Zb1Xa6Zj3vfzrJ1K36Sj/Xtzq0rKhqvdtHG67bSbqKfuo4PWh5OGLKwBI
S0k19joSAVneeOfV/MMLguhtqiwbcxih1/vJddL9Lj6FdTa1aRcjoJDjaXUqxDlb
chE0B0jvM0uVuXA1AbBy5zujXpk8eQ0/pFI6u0+oZKvY4CwoVqYHIqnRMhiZWzeQ
HDY8JDM4NX5IRWbIL95ABaO3xnVUNant3yQO9FkWGjWitpQkrW3N47Orfga2uTPU
0ZjV2krsVV6wKGSaGZ4I/N9cEgHcCxQdyKEb0puJuUSeg5sgIybNBA4Ktj4S1+fV
iQv6PL4T3rDWqewNuzujYhP50InkjWqpl2SHXMH9KJZDI+jTnFMKoGbwPScix5H9
r6cjEK8Dj8F1SR9VRDXMqex92c5fA8XPcCmAFkA/d5CtcmMZiotLSOXupU2cxJqI
m4l7MDyCySopWxRGrrgQrHwjKCRbHgdayv8VYm0oBRq0vc6dwDiaNO7RWrYJWK4C
DkKXLZzqyLkP/XcaDg69o978ZUzVHwV5cN4uoW0dTugEByBxfENEhUdo82/4avfc
FJ7XdIzcQtPW61gZoAnLIRAg+nlsub9gIlseKITT4tcNPddtj1Sin+PXOG+2JmA0
kMQ2hK4GlecZCqk4/o7LJmCXEkRN8x8ITKy8LWUhHyA4ppcp8oWPzpucr3HgSkWJ
o13oZQUDh/sFcDnf8n1V8nmG54jDX0hySPAwP3F6fkHd7R62TfhLvFegeJm1bmLm
QorLh7VJlNArSiQL13HL8ZmTn9tjVU05bNdDFuO5nhn7a+DkrqzwDJi9Hg+qLzrn
6gOrG/C7BEhPUZgw5cg1y02q7CSKEtwC4gClbRlqM7iOd5TUi0ISel/tByaAE8fI
9oizwWDxeKhR8SEytB0QDrpyyJr7yfbh9ELb01S1Ala7fBEbzzaSB+JOFvmJFImq
YAyNiJabf+cIC1tdDqEH6Do6mYrHlL7mA/Svh350EdN8aCDLJBENPirvR6cKMv+d
/qaqlAiaAhGxwXyaz/k178NO3SX81vCt2iNUfQlg38uUkdi1D8W8vnxAghVpOHM/
0HcaYV+cOsoxVdjYyPVyUHDEcdEOSqOn/1M7lj0+0XYHSgbg0Bk/lgKB6gEr5lWC
3P2GTtsEQP2uKmSUx5Hid3QeJ9BzbG+ciQu/8oz2U5qgoY+47XofHKFiWmsQPtRJ
AJeicTKkNwF3Lw+IQ0GJ/Q9DvAFWvSuwT+heJGGs4CuQ7GauQwF3xZG/EVHcFcPm
ptuOp7U89/gnMbqeuEjxmu8eF/H8JYfHPkt2STepcDW8JhnOCJnkgpVp4d0KYN4Y
S4n+W5VDu/HBAOOiMEp0+dT3lvOlRggw50tF68wYvT7S85uJifbzt1U/0HYN1jDE
4hHKhKLdwfqb6o27i8h9NWjJ8OvPmVp6KEyfmKsO+j+3buk61SP6qH8Ct9ts8YIv
ENmEyEA5La5K7PXvoXvUFF0jNfnuy3+mPEsLwLv4K5WjxW5wCwqrFxN8ekQOse8N
hgbZgDtHpTW7Hdirg+tq0+7xWTZw40KMHgGMk18HB0P/kdwW1E3dPDxuvCOzVyhD
rx+bRGR//v/o4BZu37G03iO0WsSzkDr1zRG2+EvKBnkU41VqxCweoAHcPQljGNTP
KVDExhr/oxDdRGvPLG5j6tUWXHODfKV8NoTYVN98rwOEiOB7JQYCrXVfCqdPLTu2
2chc2D+sBbdd5iIK4IwYkPucrvUm89GHb+dt0NcvCIox7Rrb5bxr3iT06JUHQaaW
LCX6Mnu23vSohhQDY2SfZ3lcg8eh2JZ83uwVhws0tAaaAmbQYy2Sn7lbCVERjXoM
oHHZ2rX2gq0gK4LkihfcdaFBSgrztpEDVVbOGOltz3ABpHdmVoxZ1YjlgWS1P0YW
spi5sMeWy0BZcTz57cKTaCJN54jibHC3v3HmbsRCC6a2wreagbNORb/BrVnadtvS
CB6c9Iy49sgPp1zbTJN+YF85rsdT6a9JelWgrdhwUCov4Bk+WVY6OHJBYCfFahdj
I/kaPCZG4NuY4iAr1Uhoy/3Ql2R+uqfIIODzqzZ2XXlV8j4LyxgOLCX2aV3hWdVx
mRtFAjt2R3CF84+rM5hYTPEWPeMZgaQpW6pBh+gaWLqqYQDXEkYj4dy/iZNOMGbC
ZKSrq88fBb+JtyGl7rrVBipTyiDiNgid9HyQIbqSHoqJEsxZ527YrjWMWe3r7DOt
Ue2Tb6o9PUqIMdvrwae/TBWjXgykknmGa6XSifrXSWsrvTI0rXsAqBmvGKhjWXIV
JLEU1XVYZSitRgpK+9OWfF5sSa00a8woI7NJGtNb1NGftuAjSj+s7qHVJ6G8gbCn
u5qYu7QErLiPTpyM8tRckvzaeSg1bLU5AKfPIjFWrwfspZHLyffVyTc6EcwFYrqn
TpILvF5sUXuJuStIjAPub2MYaIj2FmXpN7FNiD1TlVk9JsyfOAnFuvu9cKlkpKPp
emFBiltw0muK4OGkmlLfsLmBcyZO02ykPr+Xr7SiaFxiNStNzWWt4apSlGmGgius
ebFGwalerVMdKAjHaQQaPwtXAYvrrnvBRj5ARVGuILzdsCnDRgW94boADDSQmgqh
UwbrGrWfYWA3c+nxwzrrLXUzlP1Zw+kKg6tPtu+y9lncXz+2UScCKrOWgA9I/lgA
zXytY9wKgeTfgsN0EMxTDrUadMSNs1wPitgEbxfanfsqIEfXYGIIulFEJGodyvYs
MYxB94g9kMOQTi2QWLf0JEQ52E1Ro7aZs5wxN9UK8Ub/jPSHrOhxrR4+Aun/6YAw
uWz2kdvp1TEiIOvqT65KX4f9TFQ2eaU9qoe1NqXXgN7Tr8aBzgqQNr/ZnXRkadOT
4CTPnakVoDYui2fIFY5O/QZmwaSOK+KHwaswb1+Xc1D2Rp30as0zZewHC8SIQOO0
0PDHyU5Ub5vd0khOPyQjlTR1HEM51m2E/7pIvPQsHXmUXHWx7TbiPc8L3awvaE6s
PBCLfKCaLbXkmJ2xCTyGFGllv1hW2EUzJlljqjtj7dzx2EYFg9K+TT9h0VV9Lw0v
+YdgGBg6hyJKQUdxCADPMF6KYqXf+pU5u27t8mTYpQ8dUufVW3AVAsBT68sBACJp
XRS2M975waGWm/Bx/p9p7fnBM2fvoaosiqLS7bC13LaruHXJyIEq5Yv5sVyZfU5r
xI6jaWCDfY3hu/5SQJWGICmUY8AWGVOT9sHmfbeyr4Pb0QgbEG1NdqrecEMBxcHx
u5iulOyMMSQyI68Y5kRhhDSCYDLOLUyQJOFQEpxRlGqrT2kuH8W8Qwp3oh17G2OE
+4TuilQEAz8m0noYM08fgamntKbC/PsbzaqI/IrJgE9RU/3iE1h1KlOhWzULsRVy
hAs3RbR0fbMYquEDVZL6y1G0rWgNoDNlm0EfzzazNs8hmWRychmQGWugTAf7Dslj
V+xrpS+aRI1MxibToT/8eZCIhMLBmyJKN7YK13SCGdAHthi9SbhUp7PMy7GO/490
ph3UCLMa5DCEesuhA0QJ5aztaNmMZ3xpGVJg9CkvlNQEWD+eKZSPb41SOTxx0EJJ
2gQ7kac1jpbhUvOJbUy8l5kZZnUK+2ZNETb9GIIU5+awdtUUKt4SNFWdH1f7mf9P
4bs33cJhaDXtFIb5LikBZFShT5KaOYdWakryDF7FPiarLfE0+f0IvlempyCJKM+c
vsLmg3w5FZIs08INUfQ4zWZIIY/ApbqV4Pp10hQdLGqpQaUtCcGY0HlWltSRuebe
Z/gML1/NCnz75Dh4l1Urrux3GrSO6S3DxDionSstxwDGpIGZo5SVaHumJAppRxRp
KUTV0HRkXlqeqkOqTSyWm5nn9CUjZLWMOQw64HCQ87S1D9Yu8q7w7Rvc/2NArHgV
No6mp9DRFmM0kJNubKMaKGy3Lz+ChKSbNceGBC7GuC6ra6iZOkVG/VoKP26fQe7B
6u1ucnNQpcRf+uo1NrVU2QQsQTmRJl1p1Cl3OtWlRj1O/wdCAZVoINvbbl1Ay/AO
VoFL1/cIWPw6O1hISnyvexpohsD9jFXl1/Vn+dCzrUPf4UwCAdN4JAHL+2jTye0I
hl2FMASczZ7QpX0DzxGYcqeuCBKsHPcPQPg4+vwY73M6YN0pJFFaTu9iUX6BlPgP
qhlNQoeF32EV3IrlCdF3N54Sxm3kHiuR4Au9vtGHbJavBRR1up8WrZcVWKc4J+wa
m9sojuormg9fXHen7oLcjUyURCp/CU4bdTyx7PDhT8wIsMHxYsbG7MgDpr8s2E4u
rf+6/CTMM0CKo6u9wxSTcEj2KTKfAI2XHHwH2CqeR1xIROS4muRlCa8atWtXcDTi
PTvklAZWgpT9UtD5ujpuGm+TlEO5djhSAb7KQWk29g3Rza0iysJOFuGmLJDs6d23
GX8P09aHTSjSy0JFJ/38pN6kgUDX1exJcRMGpnsz6nJhPX7IO1m1JmdW0DEQ8vLw
AsX6UqWIpCQzAntOcGgA8gU/xQq82MRIwF+eovGdRqhaBzQZ2ApOBrrXG6Jknwlm
8uJ2Vd3EItkOXcdcIjEbDZ7KsvRR0Mn1jsLk0EWi5Lxa2EAcLkFeZ0vk6dPWAbhm
juzgz6hJv6KwJbOEn7nUOsdQGldGVre5aSQpBdzyc48eEaOA0QyxAX2ckhuY7ed/
d/NYkfJ6oZZfbMVXItbvT4sGME7X+pyZpuBIdyplYX/zjfYQykVKvk/Xl0ejHRgr
qZYHfBVTTiYU841d8NLCKS7ZHFF8Bgi4MCvwyQ9cQ8Sv4eVQiSsAVQrMZLbQN6r4
8IOl7gApG0nnvlPQ24d8cVIstAdOAteAUbpcgoMLMpng+wWXE9roFNJzhhm9Z7fz
6eHGRIv6ygBWTk8fbLCjDQxNvLwrldtemfYkQCtADQ+Pbrluk/N9wixhkTmQ3U8H
GNACgjUSklcyx7JmaB2ANIXOaAFAg+SA8XNllJeRymoBlSkHSdyY2o0VS3IhDMR0
LAYZbPz9/oyTNUgMZvU0ZbjJSAOg1kOcEhkI6hMVSYm826YdUYF2Nchj4E/FkDKl
U5iaZikf5x/uSn62N0QYttHbwAvd8PnM0VWAV9BHfMV3F0SFWAVaeKtz2K4WVas+
PYsetSupIqvaSzTMKo/bDzpIMfsNOh7G2vgiKeWu9Z29+ysmPhThaSvHqGhoCY5Y
N8IvW4DQHMZSzT5EaFbTN1ho2By1LOvcJOMCyuEy8XsrRPIJvpdSCqYKF44HEZkE
wPOAxU4HbcwBS6fpEw/FiohxpegWAQP5Q5jsvs4RnPmFSxU+g4lfWEeIUxCxU5VV
WP+ixHqGz5v27sMKO0vmjepvGPXM97d/JsTVfGc/zsgaaGuC1Is4Wq/ZAnKoD1pa
Bc89ymYCRXKXiRjSWn+2Lf1Jn8dLqol9ODwGFC5QLHaYbtPfhk/zxOWd/fqAz5Tm
6aCzZpvT8UoXwxtMqUjHbSqAK+rywdrJchNYKSs5W+Xjxx9AQdD5Jm96R0E4HKKK
5y71ZaRdfadKod0K3C8n8FJ20EIimV3Id4GXvvaDCT9yhqWhe0pUbG8kZVCcEz9C
0jAM2jeD4IC1JknepGJ6R5B51SwWrMRd0JpCyqkkGy4QE86JgR9gUYGfZMWTEW2c
4W/ePw+NWPcw3+Z3SDqXGzCAyb/veg8iDAIMg5PJJmT3yshuzOdjpvLucupe0W+k
x1un52nJSEhjDuNsKvf1T121vOn3vGebs7fWidEFr0qzmsTBNzgVSKFFs7l54mf8
64qECZ+qpGj9yU/FqOFUg1gdzQhlmM9sP7qvGmnHeoTLbqPlVWnYNI+1U0vf8lbY
5MlnEH0HZRKFKvnrF8bt+2SQ7okvlkhlf1Nd57gbCdN3MOeZFRolv02zwGEdhvaW
JT/dFLmmYpNme91FkS7ZOWj2Yaa5+LAHj4hXMHAMQm6o3txXKGkhmXsoE3I2iHP+
OD7xv9hzbW0ELos2RtkumjMZlgiJR37QiaXXHxFd4duTXb1M7f3CyMhA+sucOlVd
BdUCdTKEReBzbLTBb+wOL+RN1RLWdjLjndequWhoIyxqL6vhvfvaUp0XXFA811af
R/mmoJGOqEmgcHWS1atBmd8S4YSnYsMQd0vmVg/XmUztp8WJ8O1b8mtFeOkRPXE0
6u0brKPSuoUtLvhidvD4dXFrzs+M+z/EX1fFQbqJLoUbUN0Kw1GRWcB+dXngKS6L
DCCb+C2RGnClHcklG6d/1xtOasZlCcumUaeNtdMYglf+Jl6d/4e/CLBoV4y0hicS
2n6hZ7/TIxiC4g8efkIoDiBh6DpoN3q3L4UNmK7DR6tHLdFd8GSqY2s53TwbwwMU
CGxuoRRykDEtgQPsIxYd04dIJs1gK/W5bVeBcaaX40eYXzLX26h6AXTdAdZYGgpZ
tgE6J06hQ6guerczBFQL4AVAxKXq7VjAyBnI9QJBtJVB/EMTPJnDJm87VIwaluzb
rNH7szZDKXx2FjMcS56AnCHs5T9jBAyCfu3IePpW5IEWHXx44KXYfIre3yi4cJY4
rdn5m9RPnwwJdGlq6006HbCg7qK/KPgdDTaXTEEiEYWrcgGVuGkkDJDA/OlFnCJ6
Y8cBIzukp5J/MiLIlMtM2UAaGUmH//40qyecI9zvf/Gq1HXsLBNT/m8vP39n/Wn2
KMXBHSp8KLHy9ZybpGSOcFhEdrK3nPTcQrGtyEGAcjg9IUZk2G9nhRY9JAuJaWbO
wElFt+gyds7oD4u3SRUeIDk3DsqzcpeS5hLwzqYPIbLZgBRbSvRDqnDtujivWF0K
/l/Vx4JvPSSkP2MXMiJxfTife6YuYiacvj/tiNsOsdY0NaJWbjgGXOfdiZeZQCa4
JWcqKMFTU2Jh8pa5A6bssQ17l/1WNRdv1eRpiDtFBZKrbgZ/mRISqtkJ5PMgUhef
rIR8AhXGHvGf30xH9cAu0LzmcL4v2r8G+9krOi1OmEK5Xs7QAcQcqF3s6SwA9LNi
2oDjOYFE8dLhc5XKQbZaL4AKV2GeNvvcM3tbgQ62LZGBuB93bLgqnFrIdV1OKB8x
QtMRDnoZx3o1JYjtYZGLau041kbC0gPTsHU3E1gN5LJJ1W/2vimfh7uOmUjOw3pE
+nNpMcjdtzCzkeaC3WUafelWYf7ndsfiiLp0qGldsVgTHUSWr167WKwGqARylZE6
35/bAjjVo740RTmDwcXZbeeaIPAbGWC6Vh+tfbjPNFO0ybsZLTg2EG75HBDHonCL
YhRKNEm5Puc4XBNGgx5l3lxsgP6742K85fDhPzSFiiDfhyYJUPlNxqJJGW4d6I+x
7ln2EK0V5t2HjGRYzcZXClsSol+y29tr5NzgBPSIXM5Dt8yjbo+j+fgo3dBnk0MI
fsKy38sb/jINx7+Y49LRPpnnhod29MrMK0VgickbK812m0YZoW2T5UNHlC89DbDi
FwE0ypr+FAOrFmxn9eQG2hdkkjQRsT4K4/kn/cYnz81qJiLzjLMu5l00t18JQUf5
sFX78/gFD1KgBQZPAQap3s2+I4Gjif9E0MQFZPrPlqKj/Zk2PHo9WYCTuOKVX/aY
SRD6Ov8vscqXbdW8wvuLQJuZsgzX3luyYuiCR49O1WYhSez1LZQHrootpE6k5O9D
Sr56zDJ8m61oLqQ48F9T1pZ6b72i4LR8KcOuirquZh6OfVZ3a0bDtOvwKmWpYhx5
9/pz48NRLdosLL2KudWCaYDJt0wvWhXvn5i73aRfIFxPtNv7d39aNYEcl/DGomE3
+HG2VoH/cIC+SbTBNY8BF7OZjvcJzFWmjJ8gWSGr5fTBzBoGNtIWl+2dLOqK1LQ5
v/a2MgIypGPaulv/nnARIb7QKjGtRQgYuD9Mdw429ob80hr/KA7HfJvsPFlbXfaL
hpjiN3P9ZWYmbg+vWqFe4rRhxZ33H1In2DOGZ+4qVhzSkOfahXT2cEqlZWHyGg38
cQpFEO+mupeeMXduRchKVndTEdLUrTnmTcBfuqN/Oz10PLzLiNzCcw7TF7pe+pfL
fm/iAJC55gIxAu6KhwsP3/jkYK3uK1ZkUUTLzJy+hQHOv6ZNYDab5DcTsaOp81Uf
f3ify4JGvJdpVWVl0+UEX+lhUyqHTbPXDpLUZTu4Rlo9CNg8bYFCmbI7TNW5xl8/
6cIAxHO3neHqcDy4jq1qCf3C+FZ4fhEIAitCOgfyvD7dxySpXyO53N1fJJ1Stuaf
EW7RuFEFSIUjZKaPsgIMqMzzc2PBbb1TGvNhNaFXlNwrNm7NcGR+xOvSLhIuKkKf
EzTRxgWBx3Oc3T6rtvw4Q1Nr4lxr3aL6U+ULTj1qq6Ia0OfqBCuTqjQq2vb0VqrB
lwhJGjavyK3ZYX49YA+PyiFmDMK9OMVjbWqEOUq3gcSxDMHw5pNxjQU5LL1X4nA5
KCgIFyyZ3PD5ty+1CYB+1WS2OqoqCaMn+MDBidOzPmGY/PN1ASLcwS+5zzmKm0lf
NwL1wjB6yyyqiLlqQaJ+z3ZM2d4mKQ5i8Hy9KW1R+LBYVC89kYgSur2L/1vZegFh
4q/gVBIpiw+dOft0g1K42wGNgtnKWRKM9YsrGzf9w4zoebmnfx/jj+UD8a7iE5IP
uFavGobU/Zh/MhGtbzPDRvhmGmKH1jxmuFgvo/W1HAD6TbjvdmrwzzxCO+T4BiW+
Mt5Z7PLGbR/nDLiHvxKVmVfb9eUVNV7dU9ZJ7EOEqvdYUXW4IeB4rO1qEWc/scza
zWbAPvAYbIFmctKh4YPJNbSw5tk1z+DZLV3uLwGU4qd3CSuu/IWcUwHLkcSGxRkT
OE0JYpvl/WF/4fIydy0Vq9MD4F2keF/lmcvBHa2H9YuNHwpmDDPPdWIhdQbvTSs0
Y8iVhenuWK2qAjFA3Pj9IQ3u/h1Hm4MaTxiAg6Tl8mVZ5ot6hCJ4ZmbWa89Gx1B/
0JtETglPWMd7RvywdMTYg3wlxTk16GeBLTQTLK0T03E/AgkNr+gVOkEweHADEeaA
FgUC4KEeaCsgfxzHA7wUUgoLKtwaffy2wtOb1rs2LSGKre0Z1l4SIZq7d8gzLlsh
lMaiR7TFr8RJfzVAbBTPOeiqp+YgOwmUc6GFgba+nqmL79ydl/rUUHWmZakTY0Dt
WOJHT+zAVIH8EQq2MkZ7xvQVaokBWTJ+mRRmYJU/FRpCDNBO9MYbWtYZhl2Vg8+U
2rwUvRQA8Mg0ubAw9lnSQ4XgtPwhwF0/ahCJegus/IAPuE2uRMjVdoT0D14ByF8l
2dNJp3gHTNjf2gporQr2Fc2hC5tZzySm9QQBkHGvJke7bFqeuC6WQBMEcunRkEvs
8myIZYdrxqwCisbr1c4/mmJYj5Ov3j5wvQn5zuAu84pJW/jG4uWWYjYBuee4l18T
5LK6KjAYU2Q7nr0BFcUKBt2/uq4mAW38LyxletPCZcgCxsk9YI9TafaUG3KMQWPO
R4VeWImocK9FsYg2FMW79B0vS+AqcKvhRkSPmcF5trkGegzsp/rFFqhOdKrtAhFJ
Bi4P7BT8avPeo9hajGWCQFiOFd5JWgurgdWVa6TR4sSmRIK2Diy56+6/PGNXdz6a
YFCxE5PpFmC9zldTmflDHZo+9M64Ed4thOI2RdIctJKJ89YeE7zYMt+7pUd0CCzt
XdurJNp/hpblZ0GLZXeCdiApjSzjHZHBlKM1iNnCUyl5zu5vidI5888jhS9/sdR8
EQZKem1SaeUr4NcN0vPTYrATuCL0/BDdnrW3pEH1IcGXylpuVutdf5B2WT/P8t1S
BBB/WIzKFdR3+9ruM75siPbq12nXCZfCxbC3Nwc2rXwBqIgrtAbBsr8Vbuv4b0aY
fUHRCNP9zzC1t3BnHgrDhqpk7hWLIbQMeYpgFQWerxzfGVSK+KvJYRgLKaPYHiOR
5QRQ/I8XnA4r8OFDgGFg7IwwvVdLj/FylpkSHUKhuyObPKFuwhYmi0YsGMN9YLvV
ADQq2PBjcsHVwjs3R6U0lU24mM6KKVVrkQhZ0tdNsUP5H+mevaRAeZHf75eHUGY/
Y8Hn+U/XPkwBqCUVaLYR9ez+TsFDaIXjfJzsBjJ94J/l0aXBJiSWjXoJbDSTbEu0
UCzE+r+rKkGcDQYMzegnWaBlrhiK4uJ1IdVRJhdmZ6WJ4fobulRbD2J5VQtnt5pq
rmkA/ofjs/yCkfQj3MUB+THXN+9n7QQIqlh61s7ibtOAv3zo2HfCqCHKQNAEkfs/
7QT18vqlDxAOonnD1wpoRvkUi+0CwZN/i6cNPlAeoGAllJh/KcJrQYb5KIVB1DQG
aTOz8yuyzlvj3VAA3H30u+G8m8rF/t1AnsvpQWoGgj9CBpyRJaYBIPq2aOt5ys+D
cuuwbTC7DKCTeQ/FDlD5z2Qy6wWI4UUhL8mCrcZ6ls68HJvOVmfDeA7WFRvKsdSb
h0rPEUN+ObqM5xgZrESgOqM3+SW22UEAYQ0GpAlJM6F4qkgD5lHV+08RLGHXdkoq
unF8tT3cZIPKnRJIwHQgy39415q6cZFdpBgC2NqZ5V8gwIElzdO+QwrI3tEG/NfV
dyEh/Mj4cUmfgM5/K+BNTjYHHHj4DAo6SfkcjCPaJDKU9s5/XK/NDqZ0o5Zp2+8A
V2S53qA1NoQO8d9hJ+ucZKF1GKY+e+ZySoTkUD8G3zRDfJtaakH0MJBr5Z/LTnEx
Pr2SJ0Z0VfddaFJ3vjVNaH4nmbQNKSuq9Efgw0xPCr3DrwKeSzVd1JJZt7vIFvsW
+HUcbsshrIrvUEzriWnQvZkg9eupQfK6AgA8Ike1Wn6J7qtWqdSFe+i5wQLYUHYo
vNhp7QWPiG4JfYG0WPi4pmwaGyYcWgsQK9uqQiL3Us2Av6a28perTNR1oRy7aUqR
7LxyWeY6+7z31UP6cSlmXPDegU02Y34QVZBewAkKn7ZGo3YCt/LD/59SuRfVhEu6
S1TG5KTDg8aiitIYejAiP/AfwzenqQp7areM50w3w3BW18iwhIETwTfYrir9l1op
59Byy/M7Jhmg6k3PQ7nJEd7kHpbtEtTf1aNg/B1haAqcAvx8UNuOxKzfHUo2EWJV
ud2HEJ2ARWw5thdBKNOak5/f+wdyu66K2AG4YpPF2Kw0lITS0z2AFJ8E7R8kb8Aj
8jWYClCmXD1gbQD8Ouc2R7CpNqv+3ma1rLUqYVJ6B8BkorGuPXHoZeVLKQ52xtmE
OJDfvjtv1oM6OL7hVeVKXn9g2G8B5RKIpO38DmhY8WvB67nqQmP6PsT192ClCQz9
ttZF9a6ojMEcR4O2ZQnwG2dddWaLg8xnQQV9K6kGeG5704ejXkOsDW446RIMy390
+f/2eOVXQHUATCc3A5LBj2u91cqU5su2tUuLfoTsFrBcQcLyM208LCl1GWSRUvoc
+DP0JNC2FBDi2EFIEcmssHPmq9fXbjpeAke6FhLVqVI/XTufTetG3dk1g8euJuq5
cg+/o/I4/YEBqaApDUIpJdX2UdPSdmY6yjk6p1m9xZ3AxI9vcZByAzFalqaZdsNY
GukrTZUbsf/Ht8p2DxjZ9c6Y/WYNQLf+EJLPkplgVDZQQmgsjqxNBlPPZi1HI97a
vAZlPftuqDWuK6DYU4ADYy23zxLOyyCXrH3WOp5GAlafN2rQKJ+glOA8TBz8ZL56
4lQfOBN7t67K/nUHGM4ggT/Ut/KwG5x1ggVVmfDAeXcCz0VqNC2sopcie69964IH
eSJoKCClCucR4L+rcUJ9jyN+dwRiLWd1gsmWCWiXzIxs4+FNVquBu5PfFjObGM1a
tcak1vor/55z9iKdBxADre49Y6KvMKTLj9we2AabyH5xPYarbri1QdLWjHvZeyPP
FSnRIhr4vDswYv0Bt4QJ7Fg818noRoltYMv6ck5x5waFUHSbY+MTtqsBXWMVLtVj
dysyezLKMihlZUU6TCJJRvVaQ6JIpPwHR9eAPLBfNwtpFGVqSA1Upnm+IHlhy7Oq
Ers+L8IVxxLoCF+bANiIZLF4rQBKVA3l9xFd4wZvDJ2uoYiKnuxXNM9L9aawIbcQ
M3Y0GsUXu2hooiL//3nvfYWhfEM3MQGjFCQR91dchHSfRDYp/jPwPZju27utiDtD
aKqdYi6cdTqwSUYSE4zUPyJjtm6uCor9ju9d6seOLGV6kudTFB/T5vbRA08/JMQh
GPxsHrbs8iEPG2XwJBu54SZ6oFQIOggKFgIQaMqi8Vk4uTes4m0Xe9tWWOAuIk45
PdTXdBStRQ/wVFTcu9ByFtGQxgNunpkSi4Xbv3SdIWwMvtArmUvLlTAkkQ8ZBOcR
g76Z+3s9l67WgLXE4aI/T2ob2pLUmp31IG4p2uq9eNNobCZnm+fRwzp92yFlSG1d
TaTPA/zOlHF2n/Kq300nHojb/jvdiaWCvG3ptsGV2Dqw6BXyfdNXbGT9OplEW97A
lL3RSVEEZooNjLK6yxFfOmE7pUhCZ4zIKsnxQ7eM6HV4wwoH7KhQpJcValWtZMU3
hk7+IwWnlgPiEE8XhRhECAmFjJn86i90sXGXDc8PLExW2v9anIOmNmekZcSBNAfH
J1YtU/zaA26S5myhrVpRbEoQU9M55ueRxG4LR4l2xPotwvwnYCpkKFaze08ObLiq
/sszwZU1yc7rxp4+s3m72xqkwxYQk03oygpcX5t87ZNIFY/CXSbLtTA5SabGnuTg
QsqAjplWwejNoAnrHBvQZ/MAL1o/uZK43j/DKm9JrhT45NBysfwiYQSjWJvbIIQO
3OXNNguBDvQs3sjXM5PUB9BC8V6b8HIc/W/QddQzElMRYv3y6TfAwhnUvzEMk4Gp
A3yg5Uu0MqUnKC/p5LvawSMh3b2iLkZaJo88vbf8Aq5Bp4NEQ/4L3iSZEEXZcFLA
Psd+SKzjbYadcM1nOFKWHrgnoWsaHtlaVC6ZTt0Bzg5GotlX0Bmuwick5l0e+v9+
iRI1276MJ6ijujD9kNN6bNXMwqRLdUzoCFafJN7hhWUrU7EO5o9VtbmYhIjlgsH1
g2aBX4l9z2krPPuZldmu+Hr3CiX6owbrAJT2pRH/8Qc9ujssNB6awfsjP9ph4KO0
DW9PhQwNZOvkS4ZD8XvjHVI2euOtbbmMKwx5N5EAy77AU920+QyCUzrwz9dkeDa/
kKSnrfx45wR8EHrcRUD54WxIPu6SiRMo4/Qmk/2VvTBSnFIhS/I7cQUmrbUgLxGR
lesTPhZ99lbtWW9bR0EPPntFLE5UEV6FFJM5AWaqqhz0/cmT8pPAnJU8/LTN5E0H
RGqB+eWM0+PzWU9i816MSjC+DIFJTYMSN3WhXCebnvkhREoAGkyeusoIhTeRiQQO
gzX67b8BZKZyFAxriA+lgwGPi3AYsFhTvJ4RC5cqg3SraVu1vynB4dAK2LUlQ/uz
s2/DgYZoaF5zbzFNDbIyiYfTcIsE8NOv9w5y8RHsiTSa3zAzGtnNNnY11hW690YS
yboAy/eqr/xqap2oouP/sOeWKtghHd1WcQhhwvHNo+O7WxS7Yc6QIx344RjHLZtB
HhqGKdMxL/qzf28DwH6hYzPtfpQhP2wjCHHaf6y+5/RUjfRPRr/Iph+ykDACtxgc
c5Cncsg3GU/Mcj1JSLZ6JaJO2WNogEx77j3FFnE/PBHX3cm53x+/hsxeSrd6teJQ
KiysztRq4E/nnTMPT04je3xpF1iw8LDU7vOFdkdNas+ev3PkZWpmpd59ljVgMG04
9gvm3RhhnPwebsSGZ15QMSu6dGNz0BlF8xpdYZs1zfIycLRoejOWxq44w1N18Nzz
E2qhlVG+nqAUKVVal4/8vMn9Su2sC70H6+hGnrO21+R6Y01HMDGcaoB+PuvWlQo+
x1ADcbBtBQc4UmKmhGlP9BgasYX6y6HeAQgiXg/WYEWiwy66aIyrsG4I4MYv/9S4
xu2ZwrkJwqrqfhLrc8VHHpGgEZqXJrq8u9a38UgPdfjxC3gYcn6NXse5kHdmMnJn
uMWmM2Y5UkQ6xFA42b/MJ92QB/VbTMsyaHVw+urDKQrYh8RY3lQiHblkc+vM1gpd
IsneZn5gxu/XHP5tjRWOWAhNTWG0tKEymbIuy0bLRBKk/aseTJhQWdMfzhAAY6dJ
Fm2ZV+lbXAQda1dLM4VTchfu4xcrZu39MlraJxuHB4snhTBbFLgn+kMCFnBInppG
YbGiya8JW+FsBM6/2/3nv73hjtUB1w/HuY+XgT1XUvXb+Zrlwhaimio5o6JAeH/f
dMEooKyUqpQUXbAwL+FaOI4vVW0WePm16mjwmQZUGumw29ZB1WJMGpc89U53I9uC
0PxJhhBnWJDiV2+LTqpUvJL+jxqq4rcXfhzOPK/NnF7Tw6gJIoX20Gxem90qe3X8
SKE0tXQn23hRbb2ESRtD59kG/3ZHjmKoCVM42+ARCNL/l/hv08CC8p29CWfj0iTz
as4c+fST+RPILdYNhzuTRjXxIcqQeAQ4d59pE6RCmVRBq1azCdhht1VSjLCESSdX
42si14IhrqTFU7hnXM8PrvczDcYhRPo0/SMC+3jp+auKWxSeQ3aXY/0kXO/yOzre
7dwFsAklFbvL+9cGUH+Y7KyMVb35MtNJtyHIgXYeTEUPWdDzX8qyGsat8ZW4aH0p
+d4xXWrPHOgIgquvhUGmgndR2bphZsL1z04BOWMMYWis87rJkITXwMSfE3dZH1re
pRsI2ne/JqR6wBl9lwZ51yJsq96CKsAT87ZR4od/C81TV/4GlDPGwkA9H9H7EKhN
Q/gjf9IPKCPZcMhvmlMPlvsfJjfrPEZd/aZXUgD8eIISWYRzsLuc3aPX0liRCe7M
AzewJ+vR04knHHRaMl/nc+ffiFcQJB31/583GuwRznSn0cOGP/A1uoY2X+kV0F4j
5lzjhHGUnG7DwKLi9ySKSaS7Q0E9tIgR8/9L6eLFW18sYNfIgwiL9EI7NLM4Miko
HWH4NVq37kdD5ihxmEHczzB20PnPvffEE3+FJgfTuQg4VGWifXupSVBnmTOmN8Ef
ecpBFQ2nuz8UNoJB3lsWocSHeeOrBwfNugSAHtlNYvWm+EeYec2flynZRgST+og3
NORlldvJYXcelf/0K5XKrcY6Zz19cWcQcexk52qxALhOpzfvt5z1o8WJMz4e5TzC
v+lnL48Xrp7/in7ACFS9sz+86fKbjm62xULFY+UnH/5v13FGz0cuNcskhgzKkc9M
nPQDIkuJew0T//D9Wx+BGcsw9TcQ0kxLCiaRsPdp6XXbqMnQp8RH5m1sh452wN4/
yv5knaSh4Ei1qHinFEOEBbVwxMhi9VnEuYWbtZnvVaL/3LmQoxRjeVaXmGITO9Uu
fl+c08IFiZYgS7GiqrOs6X/p7aDIaGzq0pBTOQq1Tm223hUpiHALx9hSJ5qyxO0k
Zkw8FyXDo0/g7g5let7XnbIyQqbEKCacbGmipYFcTIvwG5GUcgWmmxr2PPrL0j+T
ynoadSYgfDYewt5tJjNS3Heqe31pBvV2UL4UnaI+Rl7bfsxfUE1h7jBqLLT1Qvgr
3cPXgTSsCt+JriVRdfAaJPFjTDvqflvlA9uKIYc/iynEC2KmQ6eNaHRunTfTsPdK
KITZC8nYFp3mvSu4xLMmXM/n0WbpGW4zIHWiV9R+4AVuNgP9/Mm6YAu/RYLdKdwl
xLMoL2n/cXemEePKnJL05criLyYCjd7B7WuEE5ksK+pRNQu5Otsq+5LjCIzs7GGZ
25GjYi64tCwAPeXSdRyltSCbfOvIcSMKhRAOdpuS7DAiqD+UH3b0DEVA0ZrDb+39
0ROtG4O3l4wWromlTwr8dwHmwiC21zEYotpEJyotUkNGFMCGXxDBgx0RaUTH45ir
Z7baNZ5eg3Kpt3A726ScDOfofeLMRQtqF29aSfEwilbs3VHiwqqwOjR8hA+Nrtn4
pr8EUdDA+py7iK1doaGxXpo5I/EdQFxygMNAk8c2PHnUcYmicSceaBO4a0WEgOsJ
b3isNMKt+CEuoymYXJRb+DXTME2+cOOuuuBI8D2S/KyAB1iW7GL6NEbe3GvSP73v
uyl3Sm92ze8Gt7bPnYxvJ3l0QtjCS7aI1wcjKIKZsMxO8OU7n+Uz7kjiEueYyvhZ
xMs7lKiXC3taI4bo8rnBHKZLJScwVtqjMPfNdvZuAQgYHElL9rT6HXGItT12RcRv
hwxEupMRF8JjwcKFmZojlodWBAPkRG+D61x5yF/fXxQJbaxBurHak7LiIAePFbcG
XTzY0+7wXvw/oKbJbWgOlTAiK2eBj7sFPioGDod7KeOTExoBPM+gxHC1ZLx+9Wc1
DA/7fRw+Eel1ot0PiM0IUudLWdmx/v2QMdYSe2mFrZUVexSjk5iyJKTvf3+13Fcx
nbCKR93ioBopxuYPR2wOrHrrFBFWfBr1cj3O7U8JsqnLo1+mZG0Z+s0pUMDbVIQ6
rKNCk6UaJHNqK8OhWx3okmyw4rHDs4LXeHvN/CSDBesiPkvu3SdOH09MCRrhwPDL
TILZTPLQBLen7qxxLcLJDT394mzZws/Pm4YO1UH78SAOPU/ahNohE6amAE+dsQy7
4ZtnOu/EIc/TkndU56q4sS5Dlpo52KEAv7BwLSDsRgoqaerJxYdbOVxXshh83lq2
6EjfeS1HfG+S7TWbT9sffuGII6d3a9sJKaTXCToP1weKO/MwjRmVkt2aIdwYUQV6
DGAetEHhVRSsiIfWspSeniK3bwGd0NLtNLWLZBwJnvoXm5JZHUugIfR4wWwsFfgv
36L+vo+HIc82HpigGf4akjqP18N3m7XbbImEQwApH/uj/E3PlOcwfrFhcGPbUn4b
T+YSp7ZxdFJcwoekiN6vRJrP49aSsO/r/Y8O2nS2lRQWXllvnfgJazcyBGMN9EeK
wh+OBDSTlPjrZioLmpybNe+x2NH1URUAunD4lbF2kkxOXIY6kEUNsUFG6l0A7F+B
aQUVn3jlz3CnmhTBvKYwMZPN0MHQUkmVMvdBEoiHwmIZgeDQEP4jGZcrt4TVNHD+
vqVj+qw9RgeOZJH6f6O8jL4Z64Fhjnrx1IRx4n1Cnw3bP9lItKcN7YpQRPjvwKDh
1x6XD9eFuKAHc8Upapj3gX3xO4oj+F/1fM4iVWlMZikhth2c6/1EqMtqTMBoAwpC
hn2IRa7+wuix1QQbK/EyJu4lUCayakPFZ39TtetB1VWlcXu0KNMdWBhAtGAYRXHj
MaFJRor04aNrbmmFoZpOGMjuRpdfwGF3Jz7afbaOQAAMt20WK7eAh1E3+AzXNmyy
nBUPdnvVjU+3Sr+AW0kFJy5uEwUeIdB/nuZPKESmj60WpLsFsMj7QPxE3Shuwr+l
We6XySMFhbLzwrcl6GUNeeBnaSVMoUlP5SxWKic/bi90FuQWszwCWZSwpE74GwOb
HXhscxIOS7wTziV98+piO4RNLywHi5Hg14fHRaDVryw4eR7ZDNAPri3HuhS1SzG9
c4vV5sUYqMtVzD9+J/RsNonbp+f9RfpxpW4GCqaPkXffdHSOqUdvA17xJey5U7hR
VweqC7Ov9XXxm3eisGgRKmRQEJyJ+YiRxX8eObuswNuZGznMdax72JdRzWQ0QvDS
itXnf5ynGGwUsW//OFhQiz4/ekgX7dOTCC18ChfCs+oTldbWOLI1y7twSd5lVkh4
uBitWL2ncT9Rqv+ckhCyGP5wPIXtLZg/D2eyuSq6PSmp6+xrH5/B/KW1r/qx2Cxh
QkLjXLJVvDW7hPRoCaXKgN0pKT71JsH4uwvJVZSpdiKvISclmW/Zxaxs0IIUCxDd
mlnHMOQxD1R0PNaV2XIGZsHO8EH5mgjfbs8sEV5ifqi4l3rWBkA8Tc+IQAN12sni
6sDbI27mAje2kGULgN+PXP9PjEbrB027DHRg9/DOQG24RpylkeSxZpJABSYm3ISJ
l6uzJ++Er3TwYo5ZwJLGQ5PLbmLR6mWG0AUlsKAefWZRo1zyjNTpoBImW4Dl/98H
Mls4aw1AhbbZF7QN8zKLu9pWiH5aX7SJbdY+d9MALzaTGSysBMkBkeevH6nprz9I
6GY5+tV70TfDvQFYpwq4MWv1JSijgWqVxI7y9hjteuGq/avEPWJ3Wna765q9mxDj
0z5ndC3+ogz3xPhHHQG/CoCjBVMABt7KFyWMXWEghaSCIgCeCQHP6Ap1kGWafVZg
B/Tfryrm5i4EMtuBPbYkjyVhKRVOMRRtG4VtxbPfhffevBZEii6mip/ijyezy4hB
qw4XBJYkofsp6F+m+ryXEjuPDKo5jZOuNeZ+vNhTmLIh1xV3ME4TJHw56LdV9rTv
X7G7f9EqFToP20/597T3JgEqi2L4TQeq8/3P1K14T+uJfNT17TUQdaUqriPsp0ey
y443FUxJ1/PHJlcRFTtuT9LZdRVyWc6Je4dht+3IgsyK9t1GpoGrmjxTYkU1XI4d
0CU8GTtRso1dUHCabJl3cBlxadRLMX9NytGlI7mM7Rw95h0pXSk7EMSgm26ldStQ
FA3afXdD6BHX5gF4vSBL2osBK17J1KQ+rWthjcF/xGyYttL16b/oqIEEu2FeN6U0
M21hkW0Wgeiasp2oA53UayAXjy/5l0QFyhgdR5r3qwRvUMblCdY3u3votCiQZGM3
9tNc1YuunsiD+6kAqAxDlrl4DXgIbEmEzz6SDvsuDg7U9ZpMSf4LqhN0DwYRw11C
4bw2sGUws5VU/ogtIIExf/J8O7ukZgU5V3WV5AD/tL36a+P+/TOUO99TE8axCYrU
sjaBiJ0xOCMcbwDONb7EIgpiWwaNDDi/xBRK2lqT+jysVonnqd0BFrBlHiYPCeDC
NMrTBw569zS+KQJ9v4heWFK7Wnwl/XfedSE+/2fINTtuaqfgudheTFuVxrNzOwd9
oiLpI2znEtGd0YSp61S86IQauJFvCunns/CiCVYc+4tv0d1t78VxD9Fn/OnwBX9v
ObvsOxKxRpalZKMsYerOOnFHykOgRIPFLJAEyH2aHpUuXy4qZfS6n5P7iFxMGW2M
nyT1pr5f8pILEuAhVpQ2e6cU2w4U/PHn6ZLjOD4P51RuHjZLuf/hgeGfdS8gnU2W
+j7Djz8UT2R8Ah8jG++c4wMza2u5X6hB//kKNjdQ7acBATISwc5o8Tli/mVbY6k7
cx5/eQ0lSRdRzAVgyBx/AKZ8KcZ0O5h3b7hV5KU8gH9YVjum1N2sKmW7rGt+0hit
OXBYTPgmt0Glx48HZ8Q/99Yb/2pq4FmtV6ahKqQpKPXB7nNjjSNV/GsVl+KZoHmm
X5QAJKGrvRAqtq1E4rnftc0FU4OJATRc3LZb3WHv2X56ZurBcjRUL/RADmpcqsQU
+5XruO8zLDe2nXuGbneAmX+/jwkJQ84oUskUodol2tYZkFqW86XL0lJs/BYkOJ+n
+0+dCCzjN/MvOAorE8ZZGB0t5CbdPz8F2B1BrHWDiMD0ys8tdyt6cvUsiMVl4JPi
6BPDWO7iOhBRA2DSaZeTqdDhakgxnepZ4BsQR91OLoN7Wukrb7gjuNFYqbYH/0J4
ukxoKGQv+5rrZBh9j9c1Vovgd2nyZDX2kPu/Kz2YKWDMBte/uF2fPEULl3SuX0ZZ
QN7BFAoKZnXE6+gt8HbAZ1enVoRVb8HC1BaCr+Xua+aIMGDQChAI9O1EHW3RXwqu
8NUtQZlnyuTE7igDIuc6KaN+GjA23WbQsPt3c//hAPV1q7BucnRirm/kHgkIPZWf
2NT6ztc36FwBaWYNhHFlC9KRWtI5HEjGGOa3ZVxCTus7AspFA6N6YvMuIxL5f9VW
5VZAxGbSD+/Diop0z9Q5jGnoYPbN7mBAQBQS7XEXxwUKiEj6dw4vii8k8Smnx69N
7utGf5WnCbFPDdOQQwc8yO2Spz/MyH5jtOKB+Gxmk2D7j72yfM84/zFJf/ETg6vo
8tUDTlyOt/ymFf7W2uHBAZYJ1/Ib2mVLNo0rhCdXP3zBfFFuNJ+8xWNO7Vtfxz/r
J+miaD71hK4OTXt24sG6HldOZMEDS7uvwb43A9D1Y4JCBp7xDwv5jKxFmSpBFwmm
+4elmjeWksMXF8hhUe3V8fBBj5QExXgLnW7jcIe8hBFX/A0XwBFp7UnqUYHsqwCY
OOHiAKCqXLYUWVCYzVly8FXTNYkNXx4AsLllIbccQiKwCt7APLh/5a/+ZQyQVB0R
WEkKSXfZFkyD+PN2xP+JoTTu/0Kgm/trHw4uu0oJkG1cY3wsc0D2/IYRgs5BxOjq
tJ3uUbgdT+eyhb7wp3DAXkZrhzWsydLVVj0hCjoL6SAhPPH3EEhF9s0Rf1mRbBNK
iITMaMDylZuoXpkePSrmkqiQFiP1cHE5alDfhnJ6lDRsNxYoE4gsYbvau5SwaJsS
v668KXmJZ5JBiHW387+H/PMUePZd2VX3qrxuQbNlz35jxTbCycz/ZJexUNoJzI13
qvtI9hBJpstntdLSbnA4LEtuv9WSUfUFPnkMScRpCaixXaXalgpPwGnL314FI1na
/99bPvVz7nKRdBMylVLQ6zm2EJ74F6ytDU7b1vy3iu5bKaUtRcjj2F8K2gJL6kE4
+CyTxuCJ0asQhblZNsF31CX3r1ZqAJ66mAOptJgBzb1mxOeNnx9CM/rmBI0MZ2pQ
lAzV2kzBMJ5UMeD2UxPW2mlJt8wa8r1S+0sqs3m7HC7lORCbUXrwRNgmChRjUhpg
io78s5AC65RRWLzcFqf4tIP4enI+vq1Ss3iyqia0ftWSTDL1GoBAXCu5DLLaqjrj
qY1rZhwOyTZb3GYyjk06DT8w9cqDgJXaYMMGloRCNq9EWSVyx0IKN6SU7G/IvuWY
Ti4IHv+h4pe59D6XTSGPaGlLDMU9CIlply6lf8oiO8V2zqyrI0RfoM/ulq0TL8OA
myprx4Wuu/EVOV+aTqS7dr/YQwZMd3SixMc4wA1sRV837paI9WeoQ64+sXfmJ0fF
p4HPcNzrlWXijtJkcYrnMEL8Zm8FAmBqKuvd9r7tlppxCs4R+C1mcYmlidzdk8xy
B86jE7KKaH5P34b56M1lp1IXZGSOhNU2Xd6wdW7kft3Aj1hzMEnXHbtvKytvVrPR
064+kbjUwk57FQg+MKNmP1yJrdmbaRfcy+FglYiaer1LTp0Lmu3uPzwKwOlaKjbD
bme0KzNABqL4B0/8BDPIXi0e2eZOMPIXZ2ZpxdIY4lAZstPXnc9lfakr3qlwzSW0
bWOnkDbsHY+0wDI+ocH8WECTLmmlS0yLJqkYVX6iG9OQ1PYe5903smYVJ38rFUF5
RaF59z5dxT+qVTVEAMcKB/PFbrEBhn0dtj2sT3Fph6SXnaEUI8/DEwnT1XnbYdCU
BqWemMqSVgAOGX1gYMZXW1WMsm32wxqbVRGQDmePTbF0NJc5oLDcQiqnEAWdng6v
Q9LUTYkJqLioCkLfKzxUTj2I+129SFNHYfxGjsdFSbA9hSVgxC7OzOLfjMGuvSA3
uCO+egOHNmef2nA/wNLkeXnhcMsbTKOM2PUghNfrr0nmEij0fwiob6zhb9sIGLhZ
Q7kAVViw6WE1wNegfReRUkBlkEnkgsbK1dgqA0ovuF8GuQgg6Ia7Zdi8yda2CHtQ
niWGsDP+oYZQsOfMPm/JruU57pTx9+OD7evBACUcR0uLY2b9OmnGlNJVgdf62MIX
HFYp0AGiKjHd98oMzC8vPfPzaiOzMql1iZG47u/xSac0/QKIdYiI1iTt9zYS08XT
iU0CjELot1x3jcMTOWZBtg8wZuOa85uSt7QobXkyvpv5zfNEvpNg3auKd00zbpT4
LbXKAta+LpPJ8Y0pspbsaLE3yaQ/iA0eY5CG1vRXOc+6duzvpBQ8cDEfLvrQPqdh
jWPeuLcQeZe7lXShE507drjtsCayMq+1Esz5z7wdNI+UZgOTnT+9AtKius1QghQd
7zqG+K5nLO8uVX4nh2DGJ2bV5njBTYLi023tFrjpJ8VkJH5iLswnFaLGCOJM6LBB
cnz4/Hwbrnf75UqRoW/uWyKQ4apC+uAr7zNx6O6tx39J2qOmc6xGhN+IvADOhdoH
+n2GuwuYM/6IclUVVFjlFCXosxOCDJPVioWrWzPf9ATTnzbLzhs5oN6518Wwp5dZ
Sir1crPu6ABFnngg2iNdUK4BQ4yN16jfLzK71AnCCOIySjF9eqVPJXmYJ1G1zDoN
ONo/L/0+8CLAuLbLToF5/w4R2eGAPgq/BMs+txMtwnXJWig8mESwL8kYA3gVNky9
JgtbM9msyMED3WougqJpCM1IZmPGF9u6PX+fJ0Zh+b+3N0Z6Pv9vLIbGFEeWb6Dy
m49pvy9MW9tR+pUjj3whHZNNxs46CoL+uF6lSA6jCU8Xh2pLEADLpbX0DXneyJ2Z
ruVAs3cXIk8fy2gOH48CFoDO51Pt4Zfn2Vu8tSFMgZ9sFwu/udgTy2pglm5ZtNQ5
rD70Q/QXR9BMFDw64eDgAm1btCdyiZKEUFhXHD2eA3wEdcII8qMhri8DDVb5vaUn
Gkl+WCfHEI3gQnbRO/mxIcWIY/S4BN6kadIzjVcspDHaqkmJQXbSG51MGfYSSdLT
qtnfEjRf7ell+cQ4GhjqiXXNRYUfyDmv+b14PhrYf6bG5jW2Y4UfduoiMdcU+J7E
njvuTDu5X9d73kge6rkLtKrLIjg02j3fKWiAsdH/XzDEZC2W5OiIWci+4P/aNyVF
ODrapJpvq1eZ+FTN6FAhyD6eTEhN5xHThzOBLo7eeF90BVKFhNkYqFV98mYNqbl6
NMZMK/K06KEL+PBEpgGrcsqFIvSGFK8OtrZ24VuTkp0zsm7ox4bDWraPr6HnE2En
MrzGQjb1/RsWs353SPkfJArKTXKm34/4ajoQ9kgM1N5PqI0m+UjdrKIuqJZCSZxT
2JJdbUcfpXUWTXnX1SLpDZPD6aSzYfpUww+O2gJWAEA2hk+0IMfw/W1i/n4r28ny
cC5W3/E6aCRoWUAjOUy9uLsSDqLNH4Nx2cQvHaRoa9or90DT5W/6V/IhcZQNBzql
KT10dVqPl9DyrWIPd/nT1d612xPfwfNiJpAh9vFSTuqKDuS/vDhpM8x/qbWPWm1G
6itbVBwh/SZ/xX083GwNtlP+0rG36dCNGB/9oo6VPbyJK6goTbZo+ElaN6rzV9n0
uXR4v3EW5fpMA1U2oCZRM+GnO3vl0f9vXDOHiIi0PYgbUTqspjiSJa3LTyl68AZW
vLApJYnl8cJw4VGIpnz4XShgZMssdLpXad6iWDPukj6hgvCnda/eDvr7AAsby6oC
GKZvNnpPN5tqHVlKmXZnf6pJfYDWU1fL0KH7GF/Ux/aw2wZPDosAHWnqTigpGNjJ
KmQO4R1KttKyc1c5CWjgJxJbGSKN1J5nMXroKKyyjf/l/FgyphdclA32U6vVME3S
ApK71qOWEJwNXy7qEfbea8/EhnqVW6GEn7u3xMJkmjFb/82AgLni242hGuiuUOTj
DBfE3Fi3H7OOxhsE+w/begQcRT8Rfgze/+NJKS5RzhwfsQ0prgTJbPQaV7TRuIJV
8iHyqMLI4Qg4WhxA5H7D9hJTnTVxdQ/oEHCY3kUjOa7nn6+EtqhsTrDMxt9ft06C
z5P9kCE19Ug8Bj8LZE3JHslLdnfepyeAn/HZ1g8/hWqoa4KIBGGgqJObm99Oh4gU
lXXRLy6GHayHXqu3BwyLEny6fj1bzZ/1T2l2ZAS7FLwkb33PBNsPA3BvUOIxYavE
nh/A3mhHwBzHGNsiSzFQBMNwbAbiCIuSFk95E9YlgK83kfa+uc6rNBMgzeh7KZt+
xZD86kjYJEslxQiLKZdv2VOzSxWFg+nvsAJaW0BVqaVbMoNpYsDzmzEJt/Y6+EnA
IMzalZG1If65qii4EAmHeLPHwOKMEcocs0GVfm1CRBCwtIdMOkzw7pkFNiZr55et
wNqsXaf2IDAhGhWjGdWVdqyjYrc75pCFHvPd7Ja5CgRHlKWKo6iNswobuM/btGmO
AC5xF/WYzcgm0oACYHjYh115tijERzWBy0cWCVXG6OSNJE1WtLKHkTiCoRzyQtxZ
ZxN27bQ0QWUKSWHp9j4OA/tdZqKROMkHvVZf/vqBtN9C8GrecGv+7Sm4m83Bn+Lo
QipSzM8awWjv7mn6g+wh4CKVDFPCOoG5VGZ4qvsIw/gw0jb005y+PR08EF3mGfF7
xLxSRzVriA3HdeuR4tV3wWPOCHA5UYxwr/G1+yugSS1bv3c4HOHSW0kchYQBMN7F
VQel/9Z7ZDS7J7TiXcpyIHzwCheDf8iB+zM2Tk5XrUZarFT6/zO63DRSfhAUP7Zd
67UH+6xRLJ+4dusKe4IZHdz+H7yXFN8SWsVRfl2/nIYxMAhAzzvmV08fmtmgg1mZ
NTU67IJ8PQdcXe1h4VKnlhAsfQhTyzGItsw7fRGO+0JPO1li4xx7gafdmQg381Qu
k5xY7fZuyGGMPCuOwEli+xJY7iS3Ovglxcekgko7gk+ZbCVHmPMdOnLRtqi8Kgwf
cK7EJz9dXtyHGOitwNGxkibwhV/XAx7aPWVV/RXFk8CfvSeGBngy9yXNnQ5R9Zgh
yOCkgoaua4hubl+C+rFZFBVpCHNZ+OQANFj6MlHA/y6awlAytWlraxpENKENsbXw
eKMqe0ncAV/5W19ONih2s/Kvy2khN3J0OTKoCcHgwV1jUXIWkTHniRg7xJHtXVoX
zdG3L1dcZWI46H7tj8SMeQQcMJ3VrhO7npfjI8sEQ7pTG/xscsJjQfK2vwXQqgea
3meC04WQHDH8BOasvfte1BzMX6HRI1PftJCz3hvSSMaGtK6oC9KlbR0pYx4Fb8qu
K7AGqqTkJJ47qKaXli1oJhlAIY2DfMV8aJ/9sk/Z3hXKapYNkuE1UiVjps5ZuSXD
6z6X32Bgk7Hei98W/qPFCkiYnrIVRjPKUSpESTn5jVRLrGF132d3ADKIs4rb/TOW
4uyzymr97hl7xJSztglLSKT2OMQUNgXXgUk/T51ZD56R3VmwRRpHPtv1mvcLyYeq
30Bo8p/Ajt+tPvFfLNDiM7LmNs6WT6VslTaEdE4giypJpHc2y/DjNKWj/z1V9yfU
sKADPxD5efOT+OKgzUbwTQSfMiarGcXO5ODmZWn2JWfAZNmnEwRhFUvQqAOcZOsW
zqMqJ/7WtrI4f55YF9gaHJtks0BMB36bXOQE8dEH7naHLVEGOKzP0GdB9A4qqv/V
X8j5QyPhVQYqp7HM8BBTf4nWSmFKIpvmiX3rGQFDJH6mdgN8N9FNGkA+VUZPTbAU
jPrYaxFptG2P0b8z4vVrKv4/BfNitGhL9tgWPedbwtUVpVF7QIvsZteyBGNHUvKo
zNLpotcnwRKfA48OrMO3ON3tLLm5Ief5jDipCq0o/mqf2npgbblSz0vIimTXDhJy
Ew1hVMomL35Z7D2Qp8bHFZzKv2ghhR6vrxfWrD5cRE1x6zXbcqppqWSe1xj/Z2NC
LUjF+SNAatePuIrjmvp9/3OS8DDqYXiNTYJTpQpHsefCQ0vzGkNApzkRfxS+yB3z
erPqE4/uOJCl2HySSTvFxVNeR9V/E3D8uFlt4eF3o0dD3O9EJOKR0vrW3DpQBWHe
E/g/2vqsjD4STuKQl3kj7oupCuMdob3W+66PizdH6Y+3jfEBljwjhDIwjbYYIS4a
TALuYWwyvmaVMTjHIC65VHc+A1P9VIix7sAyJIkwbdmO/TlE+926+ZnKGJY0JwX8
m7t61p8zT8p5yICwWuqwqAC31BAanA1y0uhaXpH/bG96PFw36SjiHLpqBBQ4MwMe
9rHDcoMYsBNI1OCBo8CBL946xhurvtqq25N7LOOek57u5zU8JtsIC6DS4sJKIkVO
SGgDQQQTKwQ0BKQ4/zEd4oQaC8h9p2B1Lcnj6cPnjVVkKpAzIxhOkAtOBHNFpCSA
qTRawI9XAAHvzz+tNdwFShu2Qeakg7diB498ANtaJc2EQ1+J+TJA6s4QutFWE5F9
8PZjgSHZdc7N32KG5enNj9hYl7ZZxqK2uRdMChrzdTNLnr8SSAr3cgd2UYUgJFNj
G1I+KO9n3rsEnbTNHx57Fdalm5FntGwqX/mK2PrvQ0PsOvFXhUSdeGZ3XWD7sHcN
wWB+esmS80gxJYXPEsCfy8DM6qwtmVidt2lKtyuFIGwm0mXTmQBD91vMldn0B7c/
LvcgAPFFRuSDfNAxKlwWjN/77qv1eHZ6digc8vzrYIB0nE7Xb2BIlunNAuxk3U79
WGBHSBtZ0R8hIUDZODyiC+TMiLIw7BbPixUBCV+g4UiLX5xtqSOcmR8DI8ww0Lsd
yD3ZYazftWd94AGgv10rhTy795lYvP98Ll8qz4ta96Vb0h3pLoSeMfSZd1tx1bJu
NBEfvjXeip6sJ7mUUYbK58ivNG1RnmYDmPRllh+APL/GJtUabC1QvxYfe8Nin/ej
1lKgHvCbO7pZg/GDagFqPs1yJtToRWLFYkSjbn/J3UuAUFw9ejQnFmtKUFpvoDZC
P3vgWebX+GqAn+Byebu23xtRrjE78FPcxTFawhJX4YV0j0f0W3yKY8mLnMaPxvI6
PWfh2OtxA8s2F17pXocw2ktRjPrN4pQSkzHEa9Jr1otbkXxuuNAJFo49lQEOJYSo
oab37/6PzwQsYHQbmNwQ3I/cWjHa5s7Sp2h4qpc6DfFunrTspUdmE+8E+pid1rEJ
69mbk1LCbbekJj/ODRcrqbJYnDxM0aiR/AJIPLVySwDH/aZP6eooeR/F0e6MOo1f
nt1/Icy9XxRFaTraAIVH3OxXEcooXTXs+go0/bq6u38lCkwiZBAxRLSTQ2wU/RKM
zVcpvU9Tvacidl1+H97paY6I9Tnp2t1zyL9jqFuNX9kH7sRW5xOrXu73digKQqWC
55AnpAiflrobeDvk06YNLzT6A6CwhzBy7cRDCavfx3qFuKTdbWF/xf3Mdej425Kp
eN/+jOFuNt5wRRfR6EMT26qnR9pBgf0UcIobWlyXQeHN79J9cq4pL7mAzxQTgnfm
tRqhs7DW9mNDdpHIPDO6BQjG4wB7yEyl4I7ZBFvlGUfiANZxN0ljuCyjKxmj0NR0
9pPIYilJD7jEPOZlCv7fiLsPGu9eIGiBOfAP5Hw8Sn61vaw/NoziZLQ0BI89vIE4
T9ctY57SDcF+CjPDGJfGmcTeUyJsK0StqE3aS006ImfA7mhFUP3Uso5x+MkB30ly
aacj08E0CuRbDRdO4gkj+UMVkEpHJToigGIt7MgubkHBlCgaTF3NVHUDywFFahwy
zl1fncCOYzDV4quvVAgIY5lGOhR0owFCtD03UolQPlYyL8LA7scWVsC554xzcRjU
r/FQ+Hx5AEoqBRTFlSCclsoy8OLlVdg//MG6rx+aipwdng5Ay59XTS8kHC07808L
HtqnSBlwuZZlvqQbsttHaSwp5FjPSpPoWPdWmu7eZZOX66tIZB5bKOaMK3O+g1C8
h5TatvLQ0xzzqNmwvcQBlKGrROvaGi9RNfqNkNJUqANHoN82ZaCZkigg4e5B3sTg
M0KTImCxRIdcHcbOnJXLJKzOHygbubjriUvxqDCq+6y6Vuntbd7ESQGkPJJbXXLS
C4jA3mcTTAT3aZyXT+0jg654p9SIKrYT51Ktm+DFNG5FwRra0dFJ4fGSm34ez+/C
n4mRaCHbn55C2YVBsIUttIEI0LhoZPDF/Ey6ZGawQ69ne6TtyU32l2FFRHL660sW
oEmPZ5zsgJXGG3gij6Y21HEs+QxCgZSMIEMIqH6IAouQZrgKWw4BrOuQKbZqV6QU
z1HH9bIkoPxL6QahWaoJJmFDH4no7aZM52PvJuAJ0QFnwl2h67VWx2g8OHUEk2eZ
rNjqv93DWEyd9ZyvVqsK/4oCMqzav89+zahYzpMJczRVRjGRNeG8TFiOYMmxksGw
q/hhMM/vgNLdnlaIRTUr/0ZrzA68KsZEGS/5Hx7aupHFltgPI/oKWJ4sbfh4ecsd
4U1txaEvJX6lABh+R/gNBRNM9WkqSGTTV1rR6PzfzBWiwn4josB5XSLmgzJ9hwwJ
J7+gacOWmdmZ3iDniNGN0Wy1NELiPP0371IY4bK9LTlpzCOqdD8OTT3qg9yP9r+r
tQM1lWFsoKwRyIAAqnH8RGDqQq74sp0IQZ3b1WFDMEPkB9lryMQahlYGSqnkqRCC
ewNPJ1ATqxBLE2suCVXN6JP/dGxa1x3xWTGFN8hCOrTj33U5u17ztGTOnl20Nx7w
kAAZJjkKl9LYGNbpJ/7B83+OgTNeyQDWJWTPNFlP+wTXPT04KGTMlWY4HdIOmbdL
Du/h7oR83qH7cVVRFN/H/tICNL55jJdClnBjJx8XJEli4KwC5sYqYCuXQcWGuHt7
SbCDhZ5fgRF1PopE21L13l3Dk+GCGm5w5EFAiBqsF0x/U96rg34gLAZhuPu/xzdf
KoS0tQ5oGf/s5+Szitqi1IJ5DBhyq+G+A1T7tXFq602aT/gRrLes5Le7x5cdSoVK
Cxa2gXgCZ1mrRf7F1/NOZw2AiDAVnMMcbu6jPdCu8/F+4Pl/e6pxcl1aANlV7MbN
8TeRWoK+KwUBPgOZqUWjfJ5wCHwXCc5liz1z6H+4Cj8cg28DWAd2kues73EnS5TT
wlpq1cSWYgLmImSk3O7A2qSuW70O9pP3qM2V56nti4o48h507lL6uaDLP1z0Bd8j
U9SuB5ujlJZgRE4TyspVZVxKrL1bgVkXa4pwIwovQ+zZKlNJmLvAsInzEtMoXz6j
sqS8Cn7p8OYg23RlDnFjNNAmUGsB/i45IbuKVXJE3ttnrZpkR77xZ2PVN/GSVX7g
4KuqWYO3ny8Jjckf5x+r+KVzxmOSrESnoGUC+lOK13fHpmzd5UbazAgkaREsjHvN
A/4OdFe79w+9YTOZg+piC8cotcD9gL6Di2We0W2CnxsYb6s5998PYNOAmuRwULTe
0cnacb9aKMPoTfDxVWF+clp+I1m9YpaGc/7tP2OE14x9qR9wwtw4eWn2UVDKNIQn
Jz4XMkz1t5G/ErlFDfaC4e11nPE5A6+7X10wnGxgZl6r0U/94C374pSJkAz8lDeM
pIHhYMIQB7LLnm6aV/NpqDNyBfNQmgzqwXkgURQVKvg2ranDhOWk/gSHJW7uvNUo
Uv9vGy46laH9SpcQWVq7Ztf9rEXtRGdlWmWt7GW5c15ZvycfMZzePBmqQQLuIjmT
GqlrJ6I8Bj1ZN37SeeT7q5MuQAsLBIGzgtqB9rwoTSDQv0dbdxfkMZTz/Z6viapp
VC9EG7tYduzECI8WBo6sMh8ubPvroA6nBLDCkPg86k25V1fP0uHK0BhspQgPY/do
Z5RFFerKcZ96Hs2/E75qICc4viLE4k77fyXep4CPbPwY2LfqO853aL5KnrRklNBm
fGjpY30M+hy2z0enBIbRxZo2Yr/Ls4whCD6Kzi2EhKHFnpsienZ8P3kUTralptva
OMf+ygZf6KmAHOHs7q/xIYsngb8gtuNjcL0MqVM8Vdnf2clgU3BU05EQqgoXyF99
HolHU9YRWJDeAzXa4uH/yEI9cGkZmbNx6U9deQ0xK88yxmrXHehMSWgJ/nZJ5ycH
++8o7K3GobP1OcSGjNi6R4wgEjngJCm6Gu1Dhdm5oazy4ImSJI81MWVyeBvKWyCJ
F4sGWHMYLcTdWCRmLiwbjDPxC6GzAGo2tJTHNTBOXtvMmiwT6oIiuDCmIjeDTd9W
NdLJhE1TZBu5ZTeAPhyrYKK0lUFnk5CmDEZ7DFcEr2XveXU5FAX2yuUuDnHmgxJJ
52UfXfVWd7UqtZyqMYSWfu2S+5agtEQsXR1uKjfOb3PpqO4iU63AlC8ehasGHBuu
SGhRQGpJz2R8pWPPzh5EMAZURJqW5xN6EQLZ54+E/si3Opsd5BysxW6doBA25T0K
CUBvX2QYpA3mRb3qvGhYPl37sq9gOzrDKZXRbb1Dcr82pIceVmHhBP41fFtpiIqF
ojjfHyNf9gY+B1ysKJMfSk9N0hESaX8cIBi9cjb1Uy52YkIW/1WN/evvcbMdZufZ
VwgonEk93LWpZlqk6EMvzE41j62g4Mh+vW4O0FBw0MsRgpqAZiOPsMPVQ7JsfbLW
Sj0Fx979UgMQN21frMKeKdxMtCDoVXrrXooouqqf1Sun4nG9CD+kGpMlBQuaoAL7
aTFX0liahsu41mvAvPCKB0xc6GAjdMOcPbcd7x/wp7o3XHWiilPcGBdn39b+XZcP
lf3LhKXyOmIimd359M/4C4is1KdCpuFgA8Qpe6bFWtPohaUBqlyH+ASY7Cd8E3eL
a8i8uK6cE0We28YhefNc4Pda8I6iekXaT4dPRhxNiudJkQGcbrhx1MInrIn4LBl7
xcrOlDKlgkYK5N8bld/PMnKk96YCq1O0KV08FZYEfWW0L9Dc15N1+/bzF7fojofC
bQaM0RcL/6zy0AaH/daBDxl0ML1mu5oNOlYgUcuYxbnqc1q4BCqvXtZPWgE+EvSP
Fw1YfZ1ucZBTJoSVZyf2HjaYJZiDLzVKQ1PihmR8jDIWCopaFskGg0hvlSZ6vaJu
bccqDQiMy9jqnsadBz5xMG5UnW178BgoSvIxnHTEpkqnpvoYSvuw2jD6I1Bez47U
7rhhXecQybi5PX9sttn5jL3F5aDaS6FxUKcmANVLeV99RiLu8d8CDdifu6oESMMK
5Znyvt+67HJYJkRoA1Yqu8/GVkTB6r7GRzKmTB83AS4f65exE8RCH28TlATyuEMV
Vgl+SPA1jks1y6EeaberEWzCUowD4RMU4XFnoOuxJkvppl7acoOHZu4sqRmIzLWg
y0e/AvUAiVeEU6SQ42aY7BG1F41+vKQ/w0kOkrX256Q62kaAfGF3xtK26dTUxDV1
KC3rapkB3uxIW/sHDfOn2Axzl5vc08Dvq6RIeRKu/vY1fwXmVPEZu4G8QNsodGKw
OS5HcIPbs0vdEvleOcshJ7gyDddsiBcmcP17778k7VcFscpPmRmlFNMsUA+D3fi4
byT6fjV6nvU2cs38nXDd5S+o5QLc9j3j+oGsRg8fNcTWp6hcSLe3fHWe9cYo47gz
B0DzcxBoYbAZpaA33IpSEfEozYVh8V/AH9xtiv82O3p1k0ta1vSJHlLAbL1NVGW0
AFBJCjn0HYuycV+fUn+r5f5t24PIdMjeErzVScVB1jYnYvPB03Y23iWEPXf85Cg0
HaeisbVBUL8LGt7kPHRxcIJK6hXhzlUpTiq3k2Y4HOMeBi7Unbr9xdOvUjcUFnb2
hQSQ032Y5KX8fXuN8MsEVobedLY4e88uYEoB7bqzlSYlM9C6BfJ4x4mgpEpR0W0a
WVwm+EOWj9tPGXOUraDOO0jZdAEohdR3ArylejYgfr25Aisx2A+0woPwPKMs7KPD
5z9fwQaH95Y2X9H3tToRC0IT0akxUnJ1IOoyUlWuJZW+tM7nuWzlCvqkiR6V2lmm
hGyaXmdRDuyD3VLoV6PT/NPceRKCspieOWaYmNTz98+b35D8eyP+8KC4wihAp4MS
GJ7JAbkqeRifX3682gF8eNfxYe3XcfemgZIBcIRY4WVP1fgh/h1UuFhetKl91IGT
IUlJtFVfLi6Om1Wnx59dkV6tZsTW7xfcA0yejvhKOZQxQ7uQ0Jt8QvZARuIb2ZAS
eCG8r0/t0PFOwF/vFfHaajzZAqnaeMla1Xkw/ER0mrVXDsJlio6mrgQMLMxMYyOi
F874NXM5u4FwYeLZIaqJ6boxiyi1nZJ++DtON09qHuFissF6T02JUtoF4RoEi1er
j405z54J6K7pehcq+3Rd/G6qQgDXEidXJ0606ULBsJsw86Sted7VlGP+MTQF69WE
BtqA5FvJvqrPAhSrBHhJ0EuCJVipmKENlG6nZJBj7D+Dt8YeInF4YxfIi8xvIil2
cHylol74l0n0ccwqrOOaB36OEch55NH8SaUFdaOduHlIaSnkh/ZTLXRme69OU1mK
jGaTq5DvvGpZfXjoS0OKUd8tqw/DaVwiurEUWq7P/Fcpbj2n0EPdIYPWEvx40ZNW
g8YWVuv8H0oHsmmf5OHVcXK3XOHjHWfiOo/VP8hHuM+qqDPV12ipeiNUaXeh0XLS
ghIp3tdrOWctxgxzyku/75+bbKit3gbgFbWse175p04mvaV66dnuuXEi5ONMl1A8
PNb310UmQ6pVsVJ1CWhM7+gBH6HOWdPtbXDrnbXNmhOUMIoMMjNY+vPGPo7LUsHX
iJzYxQcbuPvQ8CTXx+j6CTBI2+IVBozjNMrBIEl6UshqXmgZGfwOrH6q4JQtcK/b
LeLFYLmeO33SdcX5YjvM//8XZvxYfgCyYn3OBLlvII60PZbrO3qhspC1Pb8EiSD1
PFr3s8kPXkKqrdRwkhKOSW4+WNNREkIwTvej8CN4N2/yqYfSC+Kj4lbXVlgYf6ks
hH7IZwfki407aIiz76Gqx3lL2fqjdA+/gvnvNge23fTJJC5CRWRfC/KqCP4YHMGf
3sGyzgKHELuYDOaRh7Ax8V94gQUoZY1PLOc/Exc+bkEe1juicP8SWfJdGAUzpPOw
PaHZJN1E2vVFy4EsnXKfAsl64+2LBN2OyYDle7bSLKzwt4//a1MXNj8RGFzr/PIf
uZBnQafOgs5mqHM7/tz1dy1GDDsvJ9w2tGkZWzwptwjPqMsNC3qnRX05EAqjBoFC
sLAVlY1q5MpfR9l2XnYw8KZ89tAZ3nTAyq+pT0nipHk0b7mYv6lge95UAi1q9GHr
IPTCR+CN9agXlIozqXXd0TN0eKPV71DNJAFqR9VlwCztBMmA2ibFTLnDJ1ck+ML+
jmONZlAqfZ5vnc9MID3b2wtmV5scQkr7zIlYK5FsICjKFcxBfj0lmxs4nIY8mlUI
/hKibqOYQj2l9g6lWU4ZIP3Wd7Xaz7kuebOXzH912Y+RFk/i3w90TsPDVHlKompR
a9ONiY4JY3OxxQLiyahDVKP+2HppRLPK/Uq2s5yqXGPexL8jAAA+oXM7bMCFgXln
vIvWl3acFMYB6eenf+iuUO2PfoWaog7pw68Ql+DGZosq3laJGJNALIT/OUagveCV
PB9jubJFGNhySw6niC0c52qC5U1yV0S/TM3gFumgWTR4x19pbFmMWUz/o/bNudwW
9OYcub0go2BIuCP3aMdEXusmtWivtmyrS6j9jO906UElKjRhP1GamZtA42If3lgH
llKBDDUAEam3ejIuXmrUT+WStG0+FkbrCGv4CQbvT0XQdPBITxEtPF1OmZlQUC0U
b/ARMv4kY48UGjvRwj4qfS6d6xSLYLgt7g8bC6g5oOSNdpSOggQuXRwKoNpX2GeJ
eBDopMSseabAyVeUOTyTTsuytst69ZakbaOJLLhMl2ktJBNon97HadjoMz1DjZiK
Uqx1TGcG2lu3m/RzRvmve7mwF4F0I2m4UHMpnqPizdlUQQYokB01dygvY0eXmy2s
SvI0ooo60JIdst64Ywk6Gkn3ITZV3i0oOOFT16SjxjXeDj9df8VY4QhySTEy/1Ss
qfQq9QRTBJ7vBjXdWqgdAoGxW7GDd/aLbTstT27pF6W24y7MVk37NAb5BS2MuoPR
v/cx0w/Yv+zWcwr3RSCHrkD1cQPmijQvE8dAm4gN919oRsXGdKQ3xlr0uHdtcOj8
V5h1o1V7e2ocXC9oWy0wLvBqODpN/jWwT3nO+IzjCEoHXzzPQ9ilQdV2PIv7hmz3
NMTqkXJbPXDTttbv78aV04nnJ4QCjcf0VUieloyMHe0TWJATO9FYjqqPWK0r6uFe
n0KdcNUFuklxHauyGTm8QL1keFVziUjcBbpwq7Z0uY3EWZWKXHnke/BGf/ZhSf+i
yjbidnfchSMF7Y0rXOmXAUSdqwMUPsJ+NlwJiOj3nX0EB7KdfnOHGjAFbNkLsBlD
JZjVOxQkGnXO00SISWXLlVqA5ZXq1fHAtLrKFwDITPk2Ll3YTDFUAfSFSBdmU+E4
P3H3DglX/9uC9BL7jv4J8Mxs+eMbepHTp9JJb/QNiDyRZgg8UpumpOKrcjH8uAu8
MxYWqhM7n8uK0rKMhxrxOQ1i0rDZw41IH0e0YHSMnJvmSvr+UnPtvcBZ4msFMSKP
fdR/ouXFX3FrrZF4d9dp1VzQDPPHK6pEfEiEtsw3HO8aJlEi/h1nrV/UcG3FvSU2
BuJ5dA6OTN92IW5eLGFJkHh8e7VodN+3gKQsZMbN9r1KHAcALlqX0O84Jxz11ozv
K69Z8g63tuMmq60NBZeDWJd1rlAjpXnzwUDllxbpK+g5yugl7w1Lc/+Y3OYG2bAn
EtBd1EMaM6FVz314G4Oj557ZOcZD/10ERnKfu4KchAV/ylrU4HYmpZqcFGYJi6fc
29qibIzBSIgZTO+KJw0o1oVr/VWtbH+Cba2cQqRL1F0hP+HbW/eynYvqS82cZ1Sx
RBDKv2XEMgPUSdwKc5z27UixooNrKOm9Se2cd4XBF/pH6HxUZ6MYXcdJYum+LLGO
F2SrSVs46a1LjFRFbWG3oPchkeh1l4ApDgzO2KUK0NE5NoP7cUt6nf0RAk74YiS4
AwEf4MLUgYa7e2Td05+yo3k34Wtq83vlgT/pTo8tICfr6N/wY0L5StCTUB+m2BXQ
waU9c82+IXigW9DAlEe2Xsj4a+KRmbkXDYB02GoGh0dZDuFvAcH/dJSuzL62Q6v2
9a5riK9UeSg8R5Wg1yWivyTKJu9kUZZZWoKi5OKYV5vdG5+VyD5DbXsO2ZYRWdIT
W12dHUwEhD4LvSAgX51P0zm3ROaEw7neWiRsK9ZQhIWfFr7OrLQ7Xa6s9ip+rsyj
gpOfN5odeWE+pPeR2ZkwzVd0FDsNK7HBGK1qExzfMAi0hFkMVVt1NStkNFGUQ53h
UDSD0rubOb8AeJd3pDWAD1xVkHyUD/AiXo7hT/jFADZqInJcoJoM2MrpigctbODI
Y6m7unMykrCz2znFUXNsadTY/6L2bxPp7MC+aoGD66GiNLmayMrUrRO4w2IQ1SzJ
TycVoQgyCsskYwp1UUW6WQliHnME1VxRzGHlLQB7rznfM8PyYEb1G0DCdI9m5EE7
GIAo129WOmng6JoS+CjNICfEamCYgqYOV7B/uUYPghZhHbi8n+3wKzzVsqWeMy0q
nrT4RM5JFNJz5EZ48N0GP5WCe9S/2Ukptv7H7vFunMMV+MfqzgUUHt5VgUhw4LHi
F5C+LSJ2NefVSXEd3hIyUU1Ro6FXTlY4oFfhzE+4dQqr3gR+R22NIaAlIVHQEVom
zvbx1QO3/0GTDB3BDX67yRPOmWOksXf3t0LP2uQyookN5WNftrD49pN6j561e3DJ
Vlk6nbp3blimFLgnHntdqBa09HqsvfIPv7JmsAb83GD15JLeAETHqzWxt9+3A8c5
5DFNABbauCfM7nykSlcHEmbSmlgC7A2A93Kejmc+Zz4ZuMe0nrn8Cm5ID0Wo7oN9
EemZDP2r59rxoSCO6VC+/i9k0mrtgK0eLUHtgTzOz/Ea/n7G19k1Lm9hW6i/Pa9P
9qoS79yZi1oIEcwzysELggSS/pa5zNYoAS2ZbpX4wDkpVQtFOKgHfiYPc/7S+IOD
b/WL3Msg5ok1LbWhTKXkL/YKYmkv8Xsij5PfIsLjOJkJVHHNxu13T7ys9jEDHWqN
wkUrH17fl2AtWDHCbMaxkg3OZWssXAlQZcvGUtMhDRVi7xPb++7iZXp2VPU1Z4/w
Wqwa7u5w7+NTpESOEmO/AdZCfM4iGYPBpzm2TACxGZo3z11WXioS3RCxYwCe6vrs
TzKEqtRP1kEluTcPyko0kKM6VD86Gh2k5R6h1r9bA86c/CkRyNxvwlO/JrVH/tPV
2mt/oDASC8zul1qiagr73YGIEhHNglCsGAAS4a9Gh2BsN40bowG9ihKeanCnTO0o
kayO3V/ScfvB7dYnca4AWx5+NcFV7fjDeXx2F++PULuTz1Upj7ImkJ9Iq5q41JxB
s5Ileo1MJMiJIznhlASZm6+n105nPLyYzB2eS1DFmw9oWmqNLf2EoGcJtd2Ta1Eq
2z8affDfUMlmVv3JiFxSlpn/JJtf2sNNs/26lVVwcGrRMSdqlK5SwPK+5HUCGtee
q7glM6Vmu+LJn0abJ/1Z/vovcgNZX0TCtvBtDRRt39eHZ1RYfv38tTRvFncmO+MW
peWhIbvYRFZNhOtJCfHEqQVMYhLvR6WPvw+M3zXUx11hgxUOn0YwD5bm90XxSzoe
Ik8z21guxs9aIJmZiyUeYN/3i1rdo1GLYUrVzFW7u/ph/0p1NqI6F8WAq44pbyJa
PpnqRmG9jqkJjUxY5WIkYnF9jRoaeiSxZZnN5BXEps9aFTt1sNRG3m7T2/toEOoG
YKRoktMcYVGxXzJ6OBicStm19kpEcNOtGgiWf3n1m2NQ85o1w4TNJFBOSq5EegoC
2jcpkp7aC3DLUOPhTpIVDPNRPZWYU9sLJDtwWLrQ0KraHyPpDRJw8aPxmj8X+xUv
i6qyBcXgJtkJx0rhVxfd/gw46HcFuvePgnIohWvDOqpW8G9dsdKuG3LvlbzCXVrB
VEHfJS2scASE/IDNm1uZJOrogACq6ihn3fuHyNBceA4DYhaPFYdccxJ20WD10U9q
pjAJhTv5DVGRB00GLOOdny0VIjBAiAQRMdo2IMp8PFCrXGlF5FbUeIuxxT+H/kkf
XM1YK65+Ur+u9NRsPpMvPp7pj/lR4h2oSDkX411XmHYX/TS6+3d0K1X+ZCw4jWd6
XWXR1DAYwZqYtNzpS5oXBYw2jkckm1vMB1qLgLqK6ZlrLB20pezRd4RxhzlGPaqo
6siL9/k0x60TtpWYn9e660Zce/8mjmyWNjVRPr4anSDeKW87ihllCBOMBFxBFUsM
IYyUo2T6nEiy0yWMu89pbu9w/5q88lwaLhClZPg4l2atof1plU8l8GtxiCwNB85x
SBH5KDsOTnWreYy/K8V8AxgWC/ORHY2RH5VthgPGB5JgTW5mOlQOXxKHnZ6mcefo
ltXWi7O4nGwK4gmd6Z/ngHV09gCIfy6Fde4oI2F6lj25cGpTyi5XHa0mbR5FBApA
hBAIvfy/UM+DKBnYC8Pp7jwufb2EUDHpo55EzUK/lsgzgKsfR3P0R/ty6n3MMLwC
QQ/uOU9BwmolQhLBd/cz23DRpQWLxXTinac1K1f8daGRtBHMxLMIFdcumXWfMAyZ
f8zDOtWFs+pjPQDHm/VtI0EbScpvdb0aogram/oiL4zYkzRa8CW7J87NH8l3qvQ2
4uQXK/oC3QB7YW1PA9rB/eFBVtIilE8H2n3RkIykacgLyXwRbXevg/JlmokQZrao
zrDZnIhU3pY0B31T18TjeFzElg+sSgh+/Kxxmgg0X9CzIY4XgnHUTI5Bzh6EId+X
wnXDeIoFSeXSb+oTS9LkXCg2kifX1t9QQQ975UTsoPeWO4UAlmlhSAygAYjSPhqZ
xA2MAsuM+Y0+V68laMHqmNcpcx106MUYfGmbUXU3fSgObAlkqLZs6en0sB3HRzaC
8QsTI+1DoxIZc54+eYiP6lwhR+x4xY2rNYs3IdwQVpsItI1rDJwVREptclblDl1t
tWkZgFMRapz0YO9k972b9M9RG6gr7nIBFhB7hFajWFZGT5/85PPGZ+3hHjiQ2QFZ
LAQSEhIXVtHqxu9y8ufRnj6gvpeDg7xzavUg0oAebAOik97Puj0/Y7mLcTdAVrjm
XWdVm4AmXbu7VvcDcLVmETdio6Evklv0OyV0scyg/eVNfdPJvQzM2wBRydAoOHiu
TjpFBTeq0HxRss7RwweS90ihEIkwgZS1BSM9hU9+GEoT2UMV1qQSc6opCR/b3SxE
XfZ0niQPu7P4rj3d8vVDS+lAUU6hQ7qN7CqOX+lCI2aruKDJJfksRBeHNWCEJyeL
Q8gjWKsGx/ohWy6VQTosioeFtYVknjQDA+u4ATs9Obau/Rsx6MihVDOVXqqhVspZ
ZljYTJXGmCVJqqLNdMvvUFGIlRFssVUN8QeALM2u8gY4ejhYyIQY93x6ZfftIdjo
3MhgpF+3/xTExMJZWZzqre0ezwi/iDeP2otQ8nt/CAklnaEH9fpJHEN5Rb9vp9Ik
6GapEE9I4qnjkUg2xuOhCkh2DZVnfQLaqfamOM4vCM7NWMzlKSy3W3KNx+nztfeR
vH9QI7oKSLfyEWCNg041ABS3J5I5WWA1LE3wdDBbG7paJGaqWKLnv1kc/xYPwTMa
XQFOiZO/O2YuUjcQN1cu9s4fhbxRHu6i4V0uZxhxpG2CbEXphRYTHpCTslzeR1Vi
NaLeymTMhaDIiLtW9qHAsXH8RMtDSB1HgdcHAT8d1gFRPgax+q9GkJf1XSrn4ilR
iM15OxYcI/kVjtnLv/o7LxCSy6WKn1zkuzBWXCynG790HSWdGoRMZSUIOMJ+BaoT
dE2+ZFZNSr8+L5sJgZl6MqREFsRoQgdlYm4uk0eUsH94syGyXoIhIW7JBt717/wX
VLMh0V4+fWRlxVQOvQCYVyo6i6QmA6LUXZYr4ifUVLk3XZrXX4ZMPAi7/pp3OFBz
EiVU20V9i/pIwc3E+g9uhzFN2aaQ+DdeEgOAS/jYqOJJkz7lJtWeDnE0SsdDKz5B
8VVJYE/6fv5J3ai6AZl7T9j0SAa5YMO4VIdwDB8YcJBquKYeauLPYU2zzOQn7GWy
XB1eSusTGXLrRq9aNFcpJJYf0uXFPPGv5gsQC0Gg3hIWIDBmAiiXq44un4UYYNlE
3OmxprIn6zdnTX9V/g7qHeMk+G30lWf9O3Pt5TlPmWLBjrKSK2dOonSDMvHbaItP
P5SHBUQ7eQ2u9gb72YS3O+nq0jvJ7NCBkRkaKzosZFPuv38BHocGR6mcOoc5/vxf
hFzhbbKrOBmrvmkKkgSsBpjSLB0sWogP/8cRD2OmHYMJ5EffVMI2qqOxNxNrKtFo
zi+842ImX0ynYmMd8gPvWqekCTFnETJTOB2CtDAyBV9j+Zy8p2W9qhBt7xbWf+NW
qdXw38aTlbV/p/c3eAC5oOV2y0jOlDexoSfpUzApwFFLdXgRp2Wr6UuAhfuyhzkS
zpVRqvi89dWrDO1ReMYEhsp8qbHLa4BNiAsSP3q+grI1YxICfl1rPvR9OEUDsv+8
aha8fBnJUveDU9QzXOkim3p4AQLdkGGzCc6GgEl/nIrTBzvGdxtxvQrp9cXLtLy/
i4trAddYStpjgJ1PyHhFTDt2oCPXL7u6ZQwjan3z/LEZf9QouBZ0QfU7Brw0tQnw
URPRtcG+hXX0MBxco55AlmFP/P2T8YzClVik/sMpiTDGUQGm28sGd3Iz2WJkCXXh
9pJIZUgr4dynC80XoqZRetPkhzgerkEtBe3p/XkjEPkNwHeS4mF/7SfSS5hVjxZi
TvBrE4e7hYWL+w8pZ1iWMngwDvPhp5ErOn9wkjvwJvrpuTIcpKUB0056gdfisUP7
Xw8puA2NllVqF0UQnSrcFrkzaajpx+X8KOw7q1fACcVcmTAZidgbSpjmH5ViZ+Bl
Tozv8nDG6epwZcM4YYomi2y/hEkcwpRSIM5p/OG09rqTzazihMWJ9gdzwfJ3ClL5
fqHrK6HJUFQT1KOCB8TX0c0imoK68SjQzy5vVMO60XjTI6ZH1okG0zlWssJdySpJ
azs+7QwW/boECOXmuPIdfSL1UFn83xCx66guOnl2gNAhjPu7NXoUZ7w+BfFglLHX
D6n7OSddQlyyXZoMwntFKQ0Wp6qhQrV9GUF5mpAyoWvyeqW1NJrV5b2g3Slv9fhF
9T6V/+2bC42ZXCa3JaBswnw8x/vucVx45eS5ixOZA7XtJxpRIarU+SLyMLHw+tEl
RzotSD1hHiAyWGnd2DjLlup1qu2CTKfE0vr9gNsA0nWFOs8ytMdjxxX59UGJxkEQ
9/gWuBnnVIpvO7wUQm4CJyeb3WJsp92M7vUkOwJLXqtHvZsr5Bv3rahMHIUzPR03
AqJ/8E+wL5A4APKdk8lu8yHu93VYN07R29ILn+Uk/szcW5dgs2cyDGIfmF9Tavsg
NMCyy4LQM0otohfuaRT3erV6A06gh7qSdJG/sdUishrZ514i2agxvfZlSnIdA1SZ
wWflbYDxyR0TkjIn/jEqU1U96HLKcDWqUVUk41tA3tQlfrdyN57HWoC93NFUSnje
LTAVjS56poUkZkFZUXtwhOtf+YD7KjsypSC1AQvHsteOO89UAkycCiKCuMdnNXTm
c+wkBwEN4+eM90qJ7ySnsGtUNOJmH7sG4BdPBCDJx2JxYSlgjl8pstEy8LQ1Qw8E
rSpOVKi1hS8VO9iCAgj/6miy6oH+9Iaq/xlebIUhwEeNUeQUYifIPFZuuVcU2ItZ
NnhRKwFSgyJxdA712VVWvaPdy3zglKr5S2o709b8XI9ZpJgpZMP4UckyaSQNZq4L
rldF9EqZ/5Ev23xmSNhju3leZEN7ZKyvo9WT2f/AXLMuuxVd4qqhmvkS2UlWI6K/
kFPFYnEi0dYxfae5YmYgK16sovtt9sWrK331LfaE+MqmwTg1bCDaMIXh0kdTGrLl
TPgk8E5YZs7ikK3H9sLJGzTPXRhzMYH7BdOkfX7zIUz+l7ntUCKdxxGDIVvVxfPP
Slj7n+XVhYLRu20iuFc02nJim5yg9JyoRrjS2nOF9pcnBy8j9TbUxTTyAf315JVT
hkpM1UKG7Z8P9DTvahWMA7VEs1ad1ZzcCNhcs0qXejbYfU1K/AgL/RkhcRfbzzub
yYOVXhc6W05NtPNMIXh1eV28uMXJDeR9T7uvFti9sO32EXjKNztxiMAO184qG5us
CoZufb7EGhYTSY94uy0vGpfrmYZuVaqSZO0zkMA4WaiAMaZcLvUKjUczV04wkVuj
7SVk2PPgT/ElTTJiL84455WYY0la3LgFzsfa/7K9btXyoCsFpS2+kueydscb+zhU
afwkqNRPeQUQMfDEnsg3CxRQFjoc9ga621/uLodfMDH6VVpgx5XuJMGCNcRlcHsv
SADV1Vcj9Nn42QxBeGqdCd2ZYrPM0Tj4lijquY0xD7iXA9NCCF+UUjyt6Ehw8oIn
bPU7Cbb0wD2Gm4DTPZ+7Ru6oqnR0pXD04/YPjRzDSXrd/4a8bcdsX8bqQVkSht4D
CJT9j2BaSaTd0y88vfCYkc2K/Od1Bn6jxQGWXjxjUwItSSMWlZbSVxuJbH03CD/q
8yG8f8bml8gy80zuCkAW/MKanIHPxjOZi9ESRlJvXqBCpASiYD2b7ytFK3NO0+j7
mxvYNtktz8/GunxDKNhBn+Zlw8g02UDYGOuDTBYhd0x6RSY4skYEwFVnrl62he0e
M+TCvPP6VKLbJBWQO/8fayzqHAXMVBPCRtRVA9gd6Ta3atY8hXBUxIRBVwPHCzBn
3gBgS0ULPrjroIfOY+l+xzZ1hfMYloSy0POBJdx/xT0Ce+sboNXigW6ptnEF1QoE
34Cq9DEyoUF4hIrwITcVGiMf3WmIRepENy1pGycAyxFFp69Tu6AzjAn3QUD4oK05
uQbij+pWxYxI9ue36a4yMO0nkDvXNL8a+fXEOSzb1C4+wegdritGzWwPWzH+/ttZ
YIfaUdwMKAvKr4OjJlNSBBYpEdMRuRe6SaEuEsBg+rxKsRyVeQIU7z0qnUgcNl79
Q9r8G25DWfzwysN9H6jY5mz+tMYNhEBYfQq3PpFkEvs3LNFFKXblZRSDW0rMomGq
rDdsGDdfEXnP8w8uESxE6wVpV7WhzFwx9XJP/7LqZMsj5Tjny+UKy5OXKnhJoEql
M022Fvl3HL1oqQpov8ypccQ3vAisfFS6YBsN7IyOYQo39jGtccAX1StI7l12q+Uc
FuUWYDyfo/KTDnNzifSmXf+wg27gBxuBn7XMdMYZuZe9O3i4iBPipacIWSHUiAeE
HNPLmFEsUiAQUMhgofVLauFAS96c0jehJg6UsmEYfYjKFBYHzCEViWDhBaw+im4M
xFc5OJ+hraHZhD5d4kyTF1UTm/F+Wx4GrHbPC3Md1gxCh1kIgnU5zoJfWIhKupzv
IPMLWQv4xVDztfXQ56KWrtXNb3gTTELGgEIJudNtJXY6BPIa0KjSww5k4lquxfJ+
SETDm0uR0WW2YUvfnf2i7VzE5PBSaovGbVS02+n3+wXkg3DBFQh0PEYIFJwwheLq
D2OFC6h0/AQUDpXxptPGLKL//E1jBaWY76XqhPprZq0+1zStMUjzKIHvOWPNhIV5
oRDsFAn/EIkL0+ZXGLU13AMy7LHi2FMrQkVt4KxDrWpOy0jrMkmJwWsfx3IZdXxe
cVaVFEaxNU3ZWBN9Ppml8E5D0RfqlMzbrYXuKCeh/yolxh+Nle0y7dCQJGdKgYFm
pdSJzYSUlHXpVxbiN4/J1KfV2nNl+t5Nyz4VlYwWXn9M9pBhTZPI84j68m4Pwec2
4YGxeRvMk4yvqCe3pW9sq3fR3rbl/S1KEtgETCYRJwV4RUoiciwY8Bcjp+2IIabL
aUYt0fJfq5SPJr1pCmsU6jY8ZBTe36slCH3DVyWNmAoHqnuWs6NclnIiLi/ajk0a
JAIYXk7e5DJ5eKE4uLMjxtM54ktK50UoRyEdJaNT0L0tVcRsy7+xUCI3gFqOrmVe
e/CziOLXFg3nbmKK+IS4qCVI3CJivk4yZhMWqn/FnUuhHz/EmNWpQ5JvS+JoUruy
Rl+lSfaJl4b9f3BgNpDxxlEiLtZxNECUuzYSAKN/QUle/ZjHGFmB6+VF1CjNkW+e
sAyAwN5jgIf5W/t6bfhDTv/y7/bZqXIAGI7zgcbzFOt12ByykYNN77zvKkNTisdK
xIZ4JHQTSq1biheJpJykIwtKBA9R1fgTG1OtWLPEa03WlsnW5WpVKlwTJelzxzNq
01rQtcNpvzDAupXHW0jrwwvrKktdt11iu4hp7HXOpbkjV+u20VVLn7Gd1S2BJdNc
lNRu2y+Yce+Oqsq12mi2J7WmNccWljIPpky/efUdFm1yC/d+VG6ZMr1O5nGZLGfv
S1yX1VDhQiWfghjbpyxZqXTt0yEoRwzkeARwhYpRaobm0G3UoscPsbdG2Gc4kFnM
EUOqp5yLfLHkk5afB/nN11Oc1z98sfTyKgFF+HoodEBoaw1Bj//M9ZyeaBSSQ4Ss
mrOOexTkh5ppCxT6SrKSQN+pCTFQFDVkr3XUFCmqFeb1e0gOTnds0OSXfHkzhdvD
fyELmWoVIEDJ+ZuoqwAePke6H8z+UPjwUJOeLU77v4/jdcJYGdJlN09dB4iiUFHR
rSAl4x/sP6ZcRsgaJIQYuWKWf/9mKNQaQ0hvj+Pc0yNOOlBz5KeMjpqi33l4o5Lx
2yiF7VvO154XnBPgsZfHSG+RjG3po+9rNmQIIUu59H0RhitFTnpPk73woOBOAx72
mwIkYmfmPerCwwvOFY+CNXV4VZOtANlRCNZfqw7XHP+heHb7iWJU40+KLZHwjWD/
R73yOWlobGdkIN8XFIFfl3x0aFkkDjFBh3SE1lLF9OFksDccKm1Ug0yQSu36gWlq
FHFvpnQrG+zBY/sXRiLsMsz9b1BqTD27dRazGo5Aasbj+OjNisghb8Pharn4lFNR
Bpy5T/PD9xHrbC4b4M38SqRrUQCGpNX+12XY9+XGUmxSH8RekbV3B8NC8/wqG+l/
ybk8VhRy32uBqgDL0iEWgdFFMUdO2fhQxG0BXnKT6SrnaessDQb4PvNA6cADn6wf
OkbZbKIw9wS0C4jl/2MDBxeSbcIrOM5ulxJhBvPawNZ/c15J5IBL1Rc8TM1veoiE
lt9ODPmJAjStr/pnlEG87Jlaei6wtoVUfT7fcohgs8lyHWnWQ6erEMZA+1B5aDw0
jpzCeJJeG35G8uhCckbFTovWJsk4oKfcg1r9v7hnI7nZssXTuNE6/spgVL/PK/Zb
8OBoBr6rRJ9rv37XbkTVeQhRCIA4A4c3nwj4AUqKh67t7rOzKlgKmk3t7XRoy6Ll
C+j3KYp9x+F8IOpy4w+IkmtGFBBIu1O7MCGR3SbE38Lefp4q9Q7RGMqhYiCN4xx4
6lCZ8YiIF/xdRfBsYspE6lZMvflTAO2Sx31UqP+zMB8vTRhGRUwbSZ50PfMDpJas
Yx5py5LphnbA67JMzASOFHxsBJILzfQwBnqPliR2iA+k2J60pdOBEvULziopPJg3
G4LBfsp1EzKPI5N/aX/8DeBrHhibR0vl+jEDIOCcqopCdAtZeCeZCs+Ec9DyuOGx
f+pbCTLj9W6y7+9xfaNZXmTFidp3HrFTL3k+rkWAo+J511BG5e3KjvrAZgHmFNWI
A963Q5NUbZ4XW9GmCxDCiDkdg/jfqGHpUl2Q/Wo02W+RVcQZ/epow2rQ8aCHIM7Y
sCdPuuzHr4+1c+d1Ccx6hAfZFuSgYigPUOM+irmcNCNwIARcRbNpANxR9329APOE
11uO7THzG+K21GqVXydpkcmj8UYbBvhLy3pSAHt8h1Qf6xFMnCr4AFHmAKFcWuUC
tDpTNZiYn9uKpaEaNa+xvPVVK4uZBVFTowb5Oj19RCy12fmIwXiJyJxm4FTYzCim
zzmRAGMfS6ST7RDl9dGDSsQmksURcF9tB0JHyanb8WQ7vI3oe72rkHq/ozYBBrQ6
2ZRrQcoTWkC0a8K3tv0coiwQ54duLQJw1ta/Dkr4i6wQ61dVN4KBRC+uomWA8Fng
uNMAp2O9srEt5BRlv0j6hzczOgFx1NQvMw/R3x23bchhppgycxma4Ycw5kcD0xXc
oyB+BKigdkIhJJHYcXweiO/baXP0QzgIsw4X+2lW6MJtZEiaro+CcluSk3P/kNdM
TKHcxy/w/RLsm5r3GCgZhSnAPh5WARRIf2RK2IU0A312vKihjTNlGu73FJGH7vUL
MfGw6gv8OWYyJyMdQco9clyFSpPYKYlcMoC14DaGmGqCbgUXnzjt2N0V38VbfPv1
paTRCrvuUvvzQiO3S828mep/NjBCJC1iDyKy47YCDVRmwaiq3unCkxRw0m6hZmLb
k08Vw61vaPRfKBoe8qR06l2G13EZZEAxPKITg625ujJZo842WarvuPEFmijC/ZAn
q/3TOxus/raMHs0NMrnbcEc8x4qWbahBcx1Ocx+5qbdsT8Cz1a1F+FM8nAvG3dIL
STV+miwMNQMVcHh4D8MWKlAnvY26vXYnXU0PhT904tMqlSu12J8FnxIjy+A3XCkR
RJqpZqyw08/fTTX+L6xx13HaC6LvxeVER5Ev9gM1wtRC+e/hTH9NcOlzyjOV9jdJ
emNbzkRjjLdD0z9ZJ96AXSfehjaW8w9z1Un0treuQo/G2ayrs5BhEp6K4wXBBr3w
zNTa8BOVM8AZ8laqaRfRt5C7kXlW68xVcjABMRKd1xlusqaE8zC1Nwn5prF2NN6Y
k3LQaPWU/enxjUaj+aD4UTx7+QZTtdxEKk+G8NFSnXCv4SoVm7AOWGcM4CgogaxM
qNa0aDot4cE+xet6znAdzAeP2hrijnNrpifQb8M6HWwXL9iXeD2sMrakiHa7m4JB
tFNcrcuoQZsRk7/s68TO5jU8gTz+/y7yscBI7S8uAIfnEcxAWSpurN+LrYUyRUgu
AJYWJCmnBopnjQ7xAQldkTI71cOgneeJg1ivtoaSg84yqeZFhMnI8l1y5JCpr4Am
9jRsXou0EuVRdh6d4i2LD+8d5JjIUlQGPERngtyW9ptvbiIaAmHFTrJTvcCVG00D
MVgtIbmljn6t+M59lrUtcTGHG4SWysRWh28uxyxy9it578uHWcY5BSJReyF1X5jn
ErI1huNdxCjr6RFy0riga8Um7fga9lO4zITq2xrafov2Rc5onC6X6OFCtRhxC4pI
CRvR1dvY3IrHBOtFXXWB3RHzE2WnO6pmYq4loW5ai0BNSvQe+xrs3lmZr92ihnAw
Hg2dxIrxVn74eYpHR11AwsAnU8VMMs2gDLEtfBkBRSLPqmicr21tBLqDLS9c6VhT
i4bB4tz9MCEHIKjz2ZiUvAsNB1t51/NZ8JNG1qorTA/d0Hb1xC9ds6QawxwgX1U5
hvCbOqX2fr8iMc3+1TVX7j45QQtz50KZtyJ6xosKWBh/NQvBFeVWy3Tsb4v3d7Wn
mr6icFuwoQ6tZaltWkHMIITamA0aw/dXM5ZIrcEvE1AGxwPBxG1BI4gVogMNEdxK
iRgbWLb0DIvp3cydEqGVcm7ac0+NTa2qvwWPy64iypMPYsgy//NPhBKLKczH+o4P
SE5gfdrizbWoffqxgZg3Fv9ZYHB7elBEL9/dYgU5YQ3sH9dYzLh8LWx+Ap0Xb7Nh
5JyQ040gIz8GugcH9+ATCa0QEjFLRH/n86gKs8tfnsxIVFpcymXh/NiaoeO/mM0J
itbo+78iaxqAI6I3qcyJAY6p885sdV/aCYS2Hcq0dhRx12FaK5XcakKPuMA6ELJM
H8KINMhbJW+37SsfGW1gfiuxzr25OR7xg/yR1Z/hD8S52uIwmaaDDHhtUHiBx2OT
TCjaeEWM7flIqEPpnFJA0TdTrRpnhKSDlGRzxRW3MH5cZ5wXU63++2FWAFUqgxJt
3UCoh8dalOdszEQxmuyJ51dZU7WTAMwAegJ9XVhhwDVsOg+m+BMFvsa0TqiansZn
SzXR+ZHwTg0J7KcrWo0ll6pv2hOJWwdVnpYyee0fW40ZUvbdBLUY/ApxP8LbkC8i
2LzvMVpxA6BkSgTI/TWem75ykz67XNTXpi2ZBfO0GPtLIltTLQ4+mE2grOyuu9Uf
dgihaXKm3Ij5vrIDhkDD7qX5rLGkMw7OGvr4FJ534c+ZysmYnwq9RYaLSmli+Awn
Mzd9U8JuDKc8Ybh5W73h9g+7hCO5YJuBE7qU537aMc7fjbQPFjkE8KIv+LOjq7nZ
c7Fp1ne1bQ+Rih/FrT/S5nm7f8VMX/KYGOkvwkjNu6z5uRcpM3R/Tg7eSxlaTG1N
0mSTttc4+Mmko/ZaAhouSc28jpE7GGj6UW7hoO6VGha35NmkRho3r2hQLsMMIKeV
QbjeXNqMOLfNvvNfGOuP/lbE1HMjwJ3+bn2p33dd1TuQ22BWKXntDZ6r7/mf9Z3M
2I7i3riZdhzcXCZ3FoF0E7CxwraOhXRqcqXCAqCGzYJJ/cLRY5Kz9xV0NZiZGDJ6
e+N8wAs87t6yKRX/HBd2/fYzMUc8N02uRI7McOdACtWG8inV5P09mExsOzuy1eRm
z3fq7wduzGPwUp8xxviGsCnCeOIyrHBKPWNB6OT8e9dHL5iCdf8ZXrrNQjQEjRCb
SHrQ63A6Dq6gj+eZeqIM2c98r2rYt2YKhy15Vln3KWYoAs3M+mdahNRZg/Je7l65
y3qGdV///QPWYNldvCuj7r9Nu76EU5FmDlbjojrVWbJ3tArs3Oy1WAmOx1wNJAS6
lejhqm1PF8Sgjen2w+lVkwdnodKQU0DJ9LHt46Pb6IaPaItliWQu8AzoQcUj3urg
MMApkeJ8ChAYIEot//+NPPh1bBjnltnti5HuLgqu5YuxjvPTfPx+QW2mgUFSt3n8
cFXrT8B4wqNEA169JoElSS/mNyhykEEoHxOlA7/AM36nSy3S94253jbAXXNxyTYi
P9+V+jo7iW/wcPTrO4g2puhk9ma7/eIIn1Pd6FrkcSMRAMIfVunyaGdI3isetHS2
bvftkbhkCkpCA0N6IrTot4TuiuZQmcH+uL/mVrCJEkLrvqpij5x7K6WKpmoJaoLX
LS6DmtIrX4TZ4NuIoF57eIErkzFWBlFRNsRDaT6HdrKRSljhTLm556wGJjMz195f
1tnZQfjUytAp8gDXauFlH46lnGE6j88HgiMoVvSYHmN3TpM6xN+UdPM/7Vj00/N3
zWWSFhB9IHu2Y+O3LbP+nMEmbkTxGq7TwsHbmd3Rbr1MQrGHjFZ3EgKuM8wxeW4M
SOu6Y/uwosrnC1xoCcgvPDc7Py6e/MwKfP4oeEBn5TRWwInMq8q9IkPYVTP+rgKr
VNWa071gjHTQoaFbaWP5GNvxxoP6Qa8aFI8uGZ42QVFRq3JekIWKhrvFg1TuvP6e
IDMCJHvKxsgLtkl5KGEQZWbRIE6XgMxnPb5kmSvMDICPsqRVKy0UKf4nC0OqFq1v
DQNGN23QHXhN/90pGYl/L23erj3uB5KZjA6jf6g0cvgKf+o3tElYnCJe5lDg2eHC
8r+P6aJgr02/+cdLmR0diZwHDaio1Shz1MFoPqvs20oplf/EC7olYXHHY5ii2ByB
L8tfijWb0oWWbGrf+l9SbfIE9GFYmD6pzLqzLZDE6W/tZ4eekYaBvdfn4Jqazjkf
mvdhFHryyvHHphqfoGyWoEiqiKLpxD3623Lf3Rw2C3G22u3vMWve1NFwDudGwvLN
YOsSMhEpOuKPipiAGrx4/NC8xoNG/R0Wo2wIAVMv2ymN2pRZoBhdD63L/EQjbEUz
dAPbDEozdcFduOEDKf1hvDwgZuoSKZd/inRBkz400Zyq/xbnlJdDSkU8NOHshTVY
jxLMJ98QzNVA2HszXiUlxkSV1rfCSRb2toIRxrpm/wmG5ljgNahn1se9ip9D2HsJ
3NyhUoVXBzLpkm4L16TY5dGBGc3EONnuq8iZ0q+wY+Sa9jHEPTTPFBlz0H5+C0qy
o4kj+cbNTPbMaE5424huXeeoi5yfnBHtCv7UQM7BoOHB4BYpLieQAsq/9Bk5spcb
niVxoDY/dTlQYWYp00ryKrCTbOVy43cg2e/nWTRTSiBEFo4lXlFRGjbv8LiBLUH7
M0q37+t3iJP9BN3TIGIdBMt5rRQlUfqpZf3l/lHAQ6v3/RF5c2xHWlY8uP0JUXlL
g7tNnwDd5E6KKLLV0udfHIKQKNpQ1EaNXruTPsamEtOz0h8tybqB8HJDtJp01qyA
Q/brMsl2iHiUtM6q/fu3llnjYaqqJKiFJDH2eywuj5YaddlQ2D4isgIDTALR9x/s
6Y0Qc8HiJGCgy9wJ09ydqkQi9ID8nVkenhxTzUWZB0qw+t0acy7BX3QsXVfqJpq9
RnZW+Jbs3kwyGuMVwXkjUJdbwTbeFtal5fSJ3onz4jvopLiEmpZ3n7agBL6g9FNl
DTpQ0NocQkFyFVnV3lokLDVGqeh1bzq57mPHq63ks253Spm1r1TmgE3y74kkK57V
uil7RER15XdgnP7KMmer9bPNF2IpjNaUGzxQU78HFepX2zOmeVm1c7aNhrTaFEfl
Y8o8LtDpBMj10WKtuIUnDDM+H++9/v9X4sLg6uperVD0FnY5JlWgPNxIka/X+Y5L
fF4SrilNEubLRmwA7kpvALY04GzgxU6iVo/Ya/eSTJf6L042FCvl4AafVRi6zbjr
JFva++wqjtxtvDNfR4Q09FGLGSEiYw+uJAQxGeiVPBSEsyeERpoxvlt+BGM/w7Pc
u6NJ6d1IwAV4bzngb1Gb85XXj0GnX14OcalmlHDMSBb4DlkpwVasn9P48XBm9S6c
W8M1I+Zejv9D4XyBZxf+UYJXhGdn3m8nUgvk4u2doRvyTvfkZpQ7kah3DRXbCHJ9
moeaZR+9CpkT1dJAlGFF8AEyNd9rNRvawclLEJMX4a1GgTgQ8uhmU9eLs6knEWQP
dM/O5PhjDBENcz7Q+C6ZtL79iIgiFY48DHjakU64/Bm6UUOueVNMY2VlcqvFpvrt
kBWy2R/GheKTbaVRJUccVzRXtiaYvmOhqq6DUBqLCZMj6SQPILUk71kmq2ICzc0s
t+3xIDl6GI6x8Om+FRgbmDkz11UU3njpXj/XIuxKHw0N75zSwv4+WDqFaOFb2j7q
aS2Ps/JOsicBJlVDXwj4yY5oExLBU+IITuGq9ZGjN/KtGKCeU+uiJCqC8/c/6twA
NaDfOWC09SigJfzhlu0XzV1S6Yj/YIdt3EOf3R4LvOG0XLJQyUdwr70Fzq0l5wIN
y8vyIQIYUCkfZhUqr5+abmD2Kotu5tTXzKLxR/dGzx2c1DUoIT5qh7DUmR8ZW2BI
mxWPIRBhpTdHDhYUoeUmWuFlpNBe2sjQA8j4k3JIOKaR7E0uJR1PnROyDhgUcw9A
TG7CMVq2GpjS7S3424FV8uk6WGI3n+JFrX7tW/Hu0mhyYzcBA0QeqOPHzi/hPhcx
jxR7g77kFiN0wjjwk4WVGZ/lMqCQCVW2Jv5bnH15V/q6BbHm1MfBhOCxyhVJN2oo
Iehz9mHbFX/81+Ft9uJvLP+M+UtBdjqyoaEgmBYVC3Ujvi4ZFq6euZuwoWOKo4jC
99HqkUgYgVfskGL3uSL9b3Wm2cw6WHSVdWvI7/+sdRBn8MkRnad5spzJb/dFH4Gy
o4FZkMpOOSuvxR/pKsS1Eu58+Seb0DUIfQqlyleQI3NKy+1cNbwttSMEeaTjOokF
yjMMiC1zyvsQaf5w2k7AwSAwpSvro/EBNSLtJlKPkOPyKD0lI8DD59WyCsMmlXqs
UUDZoHbM01ap7XhkE58KVDvEQtIFiW+MJadR/fMfBA2sALIHoWuDyYKuQ6k1HebU
qAUt/fSNCCSzgGguvoKLdLpPpAnY0bmFSqjeTsWgo9iNrhaeVq2WN9bW/r1omlzb
UWT+HNymwOVQxXu1THDEOLzspjF2FcKCrsT3xuqEHiVolz8d8PPK+S9mjzLfranq
+sVTOIG9DM6LctmMceoz+nFeXLmFjtpiDF3GUhaydnj3ya2F2ipfS4cKVQwU+E68
VDqPXtDWFof8YvnwqL7jR6aVUlGIGCtCFU30SbPoIKvaoYIiGu5GOXTw9XIAzNb+
ek/SCNfz5f0aNyg7YHWywtdSI0JfVLmUzvJ3+T5eA38yVMKxaIz/lLGo9/7FojNO
dGAmpB4jvgKzVFKoUJ6IL3NoDpLB4p/1703vzRbo899mLWHvZpUkXRCqOS78lEeE
JUZXuSYpQkOo8kcZcjUyDrR/+CaIbShmBkxg3PRDHu0Ho6xYFK7VcRjy3B5iMoYJ
1ugVwvhH3EWkXbf+5YQXhrDX/GUxh8eeIgmWS6I5pN09i9h/suhGbKyaHR8b2uCK
AqNaQ8s0IaBknPX3F+mp/6JrwtvpmrwXfRQpfdwvekSnZGEug6dcr3S1655Ui7y/
rLB3Gqnfno3gGSbAHUZy4ba7WKmUVL+OjX7nSVCo38BHP+jc1hjs0jiV3X6xGXoA
dP7ikFkSENvma5H9wfEE8tpZjq5o5OsJ4A38jAd57UB7I7M/hw6UhsuC1oncxPhF
uvWHhbyy4/d4KYJN8BVI+6ovExseWjqLUkOVsQeqwz7siS34TGfaFQVIRuDxeIac
bkOxUCn1ctdsuc15cGlpEJ84p1Us7ruh2HXQJliy6BcmWzwpkg1o1tG6Qh/Lgq4d
VCRnPUC2uWRkkEGVyeolVBeX7ka5bS0I1WajEiQ2t2kGT50eP7F9uUcQjDZ22GrV
r2TYoCb+Y0xNcOfPI69jfWZiQe5CKCrjT+92gN/2MCJay5mjBXXfB1HSeSkZGNoR
rTronPWraB+MdgzDmdbrp8AsG+QJriqVcRxgyQF4W0W1ezmdvhqwwYnTsQRww3H4
nx3JIZnI/B3wtLEAb9WmX/4kXZ+4sM66JnQUzUk03aTgSAjBi130AlDQBufOjN09
1WfxjLSk3AlyD5L9wFvemEhIxOFGcKJnWMjOqkex65gSiIhP+FnwFJ0MadigXN5O
upThsM9p2+5W+trxMs98sKAVEtcsFLavlZAT8D2lKHXRA8/u0gqa2isRXpG6P15+
TcEVg9TdRzDB+DJLJ8mLqTZLuPSb52wKbwVgm6BmcB+1+eU7OHF07a4RAxMaO+Vx
n7MU3lKLzbT1WjB1wyaxiEFZ09ghv1uDb6x4ik6+OjdAr5JUz4udLqnVlcOXmedZ
kBejom9PWq5gQcQtVIHg0FXNqW3HonylTOZya/ju7Qam25+GyDKB+KuRpld/buTV
lGZbcjwbFEsIWavtlw9fPSd3OPKAmvqt1zR57w0+0zTRStjocpIcaZW9xudXfqZj
Oaapti7cvoNSIARZdJ9WY0xTBa9M4y4DGdig+Gt4asQwdUiApDL4D+OLVEhDv96t
MBbH/dsj77mOjcBJxTM3pe1w3Ii4WL+Q5nzaMGPlL3ltCm7/s3xIRnqJQQYbqfZ5
3TnFdpealbcPxvMunfzKpaL488eXoYN2CxgMkO0gIYFKdOVnY8qUxscJ8nLsy1/G
c5OcD5J12jg7LXDHQo6CLFfUbcV23VHVmbcUfvYd81opU/biiRZwTZrlY0bI3RuU
N7WxEXExXaTtjUoYUNDtN5GbVmSIvLm3IqRqjgABOQxTl/rBFYkFfWHyU6C1NDWO
R5hHQlCwFVMLv2kyHC1yoU7ATD27nLMztaWtNuu1z9str847g2pI7uMMdcOG9FPs
LUqBnzB8CZKJnvs35lZfbOjwoxGTfWWJ2qUdKpKPRr/x14GdNiJxRmmFPqFreEcx
3fZBNqWmkPcjyRqey11aFCl4Pj14WJvV+txT5q/F3bE8Thxc716AeVi1ZWQj1nvM
/4jKKNn12fWdo1W9OliR/f+HPqAFJy7k9r4JNXtg0Ih3uENeS1RlnMSMCiuFCzOf
Mv7uZ+tIdaHVwjnXEGr46+EwuoNqtwfna8lbeSdIF0Al24ewKVLLBfu21IVkLn5+
rdYMEN+6hUaTW6mEJt78axDphFTDpnHIouUAoYaclrb4eIzjtXxH1NWWDaNk2Y8w
6NzAFKt7+bMQ6fqmgG/sVTg1TFvLKBkuJ9wixaY3hjvBJJDT0jrpw7AkDPvATy8P
m5wU02lYrsLEMCxmatFyCK5eKdi9B5AKvdaQVgAm3vMHrtwH4dD7FSnXLL7GNYF5
GAlOwDpxkA/BHER7IpKZ4MjsBz72UQjHcOnUSGW1FzZZpryTYfUWPxAZoVTvKLMd
908OOkvmhv5C675Ib2+nIo8WEOuGKQ46YPZzcMycx4W5Y4vmbW12k6JS2IK0lAe/
Ne4l+5JHQfUHeor+1+DjXO1rRKIEktlfKUIExdytMno4I9yPjBa2Ugw04xnhY++I
mFa11hRpbjlFHVBODoOnAPci03hnYGNToRokaYjrNm0Qlehw7+kzyRnen2p1w9tx
9dN10qpWDEBHFBoCivicqDO68wlLTCsJfg0EjNPaewXkvqpxAyQLPjoZvzOEHpgg
TxUvETPYUtn5SWS5P8JTP6BW5gNlHrqZBlzkLeAh4Dg2RFsBBTnuMQKtNzuF8HjC
lxtEkxamrpK5lhuyF4C2JbvAkJ2EJrjII4eH/DhrYPMDF0p4fOc/5NnWOy4pxSOe
ytQ5qTAc2Elk3atNJ+z80shQrZEVbCQVxtOk1Gh1fM68mWGS+SNfr4Fdt53vp0bj
Qa3w1KNOgertRwTEvzHBn2vtLv+YG1g1pzwIcaMYBA7FN9AIyfMfYF25WFA+efpZ
xT2rtbZgC5Cw59WnZsifA/qec5hhffmXYyzVFhZrXNDqf0Iwxm3+kh8lVKsKFsa9
OB9/SMip5ErDGxOuAFnU4c/I6Q5Rx0MOZYZLWiSmlAwuxOUMfQUgnW2aoM0rJb0g
oS+hb1BieVmfIVUygRWLXiLOBrwz8aJJuz/Z3VV2HLsBAdZ5Iz/YpR/aV5zK1fLY
i5wJt3Qd20C/uI6ffy68fFsgCn3+QH+RoLiRWmgXtTw0CNZLiaaaUDJrzELVNBYY
WCaQgZg2fXrWPoGTb82nFABdfZ2DOVAWTGM3x3axASVZeTT7Oc1VNC2tLQGCrq29
Xny3I/f9guvopSQ7GdnRQdZEo5WUqlrsHShT0YmP+T+50TtJoC1MkDWHP+ajtSN5
//Gw6K31OJ8XIqIKa4ALMtArC5IcaMj8ZWID9BlZiUEKW1mmF5lQ8DWYwiNrTEWX
tjhmkrtzKibYGHHovJsr2rAOEJnW+QYtzk+6Rh/fhfhcfdxE2tNHzV+J56lBcERq
J2Hz98VFkpZXzkum4uziH7RDjJ/BjbbZ4HBUBQgb0QZsg5VqT8zDJtjFhwZxxRT+
MLf8aMp5ZnsnZQuS5LNBvSHCFZR//p0jn1bFpBJUrlWDlNb3r8kFQWFcMNbqwz4D
jlF6AIVi3MXLFecsziVswLhI2ezWqtcq9SzUiUFXN3HvaZcRh6frAKoMkxouT/5T
rvDO6Q7n8M67GuOch0X5wx6C0Xl84dBN2KrcN0Fl7oQy5DYYSFCyEY2Ox7YAsS46
ZGlsi2mUBczrN2Vz3DNROxzFhOfELX4tZ/09kfKItJypGWy4IPUUujl0xbJSRKOP
9ofnBtD00TTWMuqooylgWmkKpAXllDFJXLOqtf3Q4fsI0Y4DVny3IcLZLnP2XucP
8SK48nxS4gVuOI33dj+ehybQub5pfzwonCupUkSqX1X8wk4lYZHEdkXmFigIMUuo
hwDltKRvLGU5yo4GAZsOzMVh0CAvDbwL4JTvetGImCxlc8HrqfG7xAwDHlkQGgRW
vutnRzDj+m/vde0ezyIvhelv4/NrjJos0rbg4+6Avw1L31S5vsX4dgI5PX0Ov1yi
O3dnCpakbgQohgsG2Pf1SjXzH4kaW4NXXWczh4jM65YVJHGNrU1Vkr8y4nV7MPYE
UVm3XZeVIOru9TUq2MJ552FfN0xN5Fx6N3W91w+Yae6N5or6KozUgOr6ZaENN4aI
2gQfHzv6KvJ1xHtNw4IQ3hBVPfD9Kcuux3nwIR0H9Nl8/T7456GlieOCWonR5Q6/
+UTZt9P9VBwjtqygUox9xE1r6nXmTUNcTa+Mo5Bt+0LATWfHIEG59BoHh7yhWvzo
5bT9F9yEKnd6b9UR3tVBnOaOXQ+cCb6gYfX6LUWYTJ5g87oYFMKEBNVu48r0tdMm
ObkI5SE5VX3kYrJ3U15Ummmto0Q6Aw9q5PbgNWBsq2F0qRpbhzlNpsBH3sr/2rIe
8Lk2brN1yNNFU4vUOdM4pAIDJGbqcErGPkej2jnUU20BhKnePRyrTVxXjgO/Fjop
JLHDXwmJ7oab7i2IkgYSbh9nmCZLrwlzGzgEG9bA9QRmvaS9Xv7N1dNRRPdJWo3V
/jC2/FR3d1AOvPX4H18Sd9rIRSq3or1EAKT5mEmJtnGemAHPWhC1fC1Fg66JW2F0
fropbPawGmWx7+PeoGUf0mWknmmNz6ttuvZAkf8Bg+9+zUq+xP9QHCR17LzpnOxK
kpAPPrtt5K3EdO1nq4dUVC5QcLA/qgeji23Vw/pURnqUs7+1zArNM1wkm4l+pnI6
JFlcobNn15UiH89ybNcVWVGQ5n5aZcf+3zTj5o6Iw3xBBPkwwoQwAoaH22vNG5u7
VLuDbp4qlpua2ZFwx7jp63AD5z+9lJaXD6InUngK/LBOCCJb+hR1zgT9Sf/xhcE/
M1XoJnIf3s6DfrVMa7hMVtOOcVaQzCOrwRYFxLQKtX4NEFyv9g0jAqvESKG7H13s
ZwScHo/GgR7ceDCRnzasFBwHtLOaOq+g8YQcJracCqc/4eDkLLZuB5mmOzWesg+V
NyuDDJQNNthhfMJ8Ll2VJEQU4lYU3FIOV66oSBuVRB6VKIHCKMqsRJVM3vgGtlRT
DK2bGjrRrcpufdcyrwsIXb4J3GecY/c7sOYfFADgPDqXlpMPligaKXacsZ9E9UoB
E5q5n37T2Aq10eFBYSS1/xxSpdII57+towVdUjXguRivdh6krUkou9Xi+vlp6NJn
C1zY9p8PoYdz+vHrVy7+0pjpaW2JmxgRWH07xblRkCPulcUH9NSXoSUwxO4RtTFu
bxAI4XC//0kNSxMEJhWj7olkA3FY9ZO8pXc7PUeDzugGAZrt4kyKQzcEsX752fr0
rOJ6C6xzWkWCWPPuwnhGEW8vDJ7G9SGRUMkKIj0xt9uyh3dVXYAvfbXcKHKWfKce
2WjA+2e6EOeV79M177BxE1GD7dFhZe0KG3NsX3sc9inmdE+3m0Y7KPbGsgufXXkv
IvkkGq6i4TdxQxSREOCdOf9K0gonEeWyA6X564ftmG5lGRbe9DjU7s+F783dHtJc
TA58Bx/1oExV8pkBeC2gCiOz2oG6X5T7tqGjvwCOekqWNAEqp9Ae1kPxQz66c17k
o5a7h4ry8y28niumrff+YnErlBpvmseJVXh4rXrIS/G6nGt+V4eBKKnGJuXUTtYZ
6duWhGbRsfGA4lef21h1i/kpitNVijFH2fXxMhhps38j08mKtSF05qBoIm9csztg
Rhd/gRklD9Xmr0KyRNi+1TEwOu256Tkjc4g2sTkiNCiP+IklXZx2GOxCVSOSUgSc
kepk6O/sLYKkniWpWjhk6j7S65EC/SA4mRKvqqb3BvNgTvwfgFa6TXZq6svfJr6y
ceokPGEQB02VHWKp7v0TSPO1BlInwC6VI8d7vxVN6wbP4SmjGb/HYRWoqEdvOy+A
ESCzHItFBZyZ6IfFft3i6y7CaJr9m0sUaWwfTQWErAbt/7nW9l1YcegAp98938pc
CVAkbhS1jExLhr8vbPSqUd5WRkz5vbJYCbpMBjIr3YH/0YIU0X7MdRdTzeMBugtA
zkTyMsr5CtfErvWLeMYnasx+lmayjSakUTtHdQHruPx9yo+/MhCyrp7nYh2oyDNx
o1ANz+hU1UrIZDIpeNGAmUXf7MGAN43gNEE6F2QwROHpHlY/SR9sx8Nu9DRwR8uq
BKi5DUtscsVWalRwtS0vc0lHt1hcs7KmB/4HRb/QBLJIF7gydcZWx01kh13P3RSo
UVClAdaAqOkAPib1kUZdKPXXVOPY+fZppF2PGJMRGXbIyQ9oCytGRpNDGEgkZrLk
daJocrgsxjx6iW7KykFkdKD3RiaCcfkW77RzkJiyXp6uluax8ofT1EkEWXjvIAfP
uoPJiB0TNBiffoI3RPcEByGgchrNf8s6MfYAqXhLiML4e9ISaoUCM+u8DgrYa5MU
ulwZ/97nF+dPE/zUu3iRIG4Ni+LZUYa4PbRnWC8Grp8iIVYTrNGS5f9e5WmFPsWx
SoPQxjvXhHpe89Luqm2D1j8C/PEirMyW3hnY2d/RIF6sAoNXk5YS5VJbYyN6OzO9
lHWoWnkxPqOzLp5W9PUBG7cor+Y77gw4Wb5kKCR9r69YFI9ON01TEz5CSFtAyBSl
khuIdlL1W5ZyAIvKDHgubB1ydFuTRokPVShQF5TNgmTpdTWiPZcWzeHtvRsunpow
EdUzqKj1UUJj4UZ5XI0hSEC9p22JIkS1rfgShLwDdzzZgC8JDIQOCnQZsmc3YA8j
Apj+5bMiEZZDzXbNTXPPA7YA2R/TFQcacy+DTPLRdtczGIXR8wtO4JbckXjx235X
99LtzOk/moDdUlWt5+7X+YPRcyJzxLG48kSiqeUOuUMnqWpeHnQqD8Nq2fjA8cfa
J65G3BZSdFE2Pf7yYRMSWJ4pCXi8b7xMGPC48s+Ki8nZdrdd/ksl8d4cEuKzfofL
3TDju1WITJ9rhu3wyr4Xeo0NVjMFZetbpAX+VFYPLCJTixRfV76BcDSOv9IMHxmF
Cg0Uilaa92lLP6X8tIhhFRCbcvcX9oMqilmBQOD4eJW0Ddi5RRr15OgSd3b0BDFA
aMlU22WbsfQQQDuSg0/qLDiIFRm1yapmtjKQgppOFFAJfP3JYfDwVnyDgurZgy8f
Bq1liK/wQ0sUNKDXmCMBWCVDlcay42duf3HjTz/91mTRXYpCS9khO/9WJclzZYhe
Sd2px3MTUJ5/jyyxfbGKJYrsMldsc9kwPI971boaBkVHtLyqA0bXPcIvUTxKyBvo
PQI5AdB3mzArN2KopKh8CjKcfdIZjWu2JWEEqbLe0rzd0+oexEjPQYbzDI8c5bNM
KZxt0RcYklQVeahVOsz5LTl37G5j/rSROwzu8iWj9DB8yjcLdhUEC6Z1NGI+unvB
5+pSbJGNxD9oj8GXdwmw6PW44jR96fjaCEQi0xG8b417kBUhnH+V0wofrSRAHh9V
EuItpOdyo6fmYZWX/sHDUjMbWjpp3sbFnJLHVcLXiYxbhbjAHFGwzGkBbbvTP+iU
GA8agjIZAk6Y2b0D1NttgsOf9uAw+7rOlNkqBBitS5gJnW5LBzaCAuVs++3JVQ4L
VLT8n9kuvf5xUAGjMXT+oZvPGwrpDPEgBfBgCjKP7nf9gm6x0TEYYYntQDvvefWo
kUUa6bgeFFlLA+Ltl0klPn6ck3zFBZgSZMVwi1+Zlg7AEO4aq92aC7Bkd6qHpM05
VnP8DTi69jQ1QCE27Hawl8QupFjZQTWaLnrxjTlsgSmyU3rw8mV6G8tjs7oOZdUW
eb0zk56yrSB+63vEQO2ku+HCaAXqCZ4c6fwdz88YnGY5wPwW8MsxU9eaj+bYo/oR
XovW2xA14RGGwwU6ZQfM4EMBy8wq24D8CvL6TDDjyoAM/2YXUAlg4MMDDaKW4qgc
SoAwjZoZ+vTeU+7U7gyFsscBqpGXGsEwVAG9ZA2fgdZMeSmaM8PREaTlf/O6Kj3W
Y1CN/5trElXQIfpMEjaIltGR6vx6txjxMtOLUTC8TDcQp0Lk+q+4ZSjn2U5osPtJ
+JyW8DErFspXIW3pxiTi1zoxa/j3rvyEIH+Fc0hv7Hy22WvH23zzbcqBFEB3WKRO
dw95EYTa/6uIuNwyiROWRia89rmH9zpJ4RJbVlUVkO3HQZpvZ5+4JdtctXDf2xka
XFg3xVpZkhYQE1x3bO5SZNzwWei2IqI+xFxN71/in3l8rfsnkSjEQSG7pY04YlJf
aQTQETvhmHioEpPCY71+arhiYxgaP0aOlQobKfuFqvqw5Ipk4DkgPwqBicr7d9T7
aayKaYztMKEkmpV4PxoDApi8EO2tHw50hPFuPZieqReoQ4Y/Q8hPVvw59VRr4P/5
+5PMjKLKe3RpR3i/N+vv6qAzkSKYG8bycvSjl2/67IjThXEMiE+9xu9C6TM3XMfT
pqZ9jUw0jBlMsUWyVN9t5EZHv9q4aD81un2L5nhhNUHF2R6dCgaByerBmzs4crKS
WAWP7rvevXNf0goPCl+HDUD7Y5aEaPwBq7l34nOucRX9NMbQ2viYfy+qG8U/FesF
XyoYTF7PWVWapfS5TIEqym0IKf0TntIuhvmPf7UTZiSGizdi0lW8zUJtz4yaIyEW
g+LxH8ukRqbofd9g0sYfFdp5OgIC1Iru5ge1dAaU9tMnySvTHA/OtYrPNCeX/4V3
V5eB0sSWFLQe7/ptVGZtxZ3aBXY+1/XbD0tT2NDJ65ckePP241Mi7JHtYEzL4wLT
VvQyoAgjUgX4ECX0yXthf4NpCrjHJrBDHgm3jpTGSHz/xj3IGwm9Y7s4km6MTB/h
Bnh/8yhJykKYKJbDyRGpR+IJLeO9an8hE7CtuyUuXW4wkOcJ/8EPL3w/Tmjc66T4
sdTsPlfQqSvsORo1S+QUyOqipU+glmcU5U5qHMGtPYaEhVyuWVEdbgChJIG+mNXz
DHqouD2pkVcYLtNqArWyEhAfgobnEs3OONZaUP538YTRHtVB4Px/xwIeSba2xTP7
4XbnnZZ2ll7HWwNPeaM5RjLpdVUPoKM20zu8abzgmacvNKfjHoWDtfAyLnG723zP
Y2ARUsmMo1tTREcMpssv519gaueim+u82GCOW17nw8SOe783MTcBnecVr9Tro11O
TP8LhfHJggmmbrwtSD5HPtJd1s1PBAypRFPrNcuYriIQfooaHpPSm3Sc3tP6opXw
bATBCGU0m9qc59Kx6ZiefnbStcaXGItwpxvMQF8p+ODg1OzwdcTFjlCw5GLpPyrT
QXJksKqKjbHM3+oakQTAdFBmBLz/d0EXqSax1ufRzSX4S59J/PaI7K0o0zVmIEe6
MaeJsCVojpRp8fK43jJXYUYBzyFKpjjA5GcmxcSunu4AD0d1K/9kJKFaUQfVMclv
htlwJqv8KxPyvN3gquxgndu0RQvMAK6+D/PnlbGPLHt564sHjZ/PTHzMiNHzZsid
lbD1pTUxZrd0M15a5U2c8bMr03ygDw3ggfNVTltbyO26YRpUnqj5VGSRWlE5qCT4
dy8NANanebQdWFia/BfNCaGg01RpwuHUINq3T1FzjK7mMjt3nWXD5sK1VAcxbBrE
UrQuoidXs4ht4dWUyca/5NIangYO/X/cNZCPlJCpNRaXuUP5Vn6zlWECn5Opaw4l
J9Kk3JXzlQkRinPYdlaVH37CZRxu3vrg4EwcFNUoCNKLmdEW390xA1P0zj+7V9F6
FzqfDSeyB3Wb55LosKNcsukhDA3+eCAJvZ21gkdOh6uOMi4PaRO2GqtymTBPJEdD
PQfq3YMCUXND4zPWtT7pucoh/Mmo2eVkqksNJa6XqPt8Ld3F9bNXMtqgS8MiB6ww
LNZG1lpAVqxfV4yva+TTmpod5GZCKmYUafRXk4xhxHJYYn9kHHRzEGmooipcWw3H
8eiR6DkIYKW3UtVsXjb8I3A5R59b8tT2po1r7EFW4US0FBoQlK5W9crywrbPDmoH
XjOpQsD1p15kcOfwcYyobfsBwRqUnSdWXv4oXypRoTwO/IHyF1SDyo/8ukfagtJr
9hrl8yD0UHyeGpw4drKj9NqWJ0jWxcNuW8JoioDBpz1RU8+qWu2wpCykBICjhKup
ZTpk+xQ0sZdr69KQ4wgjRBbl+u8orba15GNe4MyuPxn04F2IRIi6WClYnVIorUt4
Mx0WIA6YR05IdIVE4Pfgu4vWthIast5R38JTCsV+0SyXYf6d8ZztOmDqLjukOeLi
oLx2XhbHNlzs8ePaJzTeCE/1vVd+uicCYyni1JbmJNQktDj9yFZKr9LxCRyozSmm
7IWjCduqToCVwHq6+TmJyZYdaIn2ODWyyzuSxXC6tPp+CM6RRjlLWdl2HOY+O+bo
94MTYVP0YSvWzAz0tSL2QiGfihkNz/WbbjRI9Cbp0W/2CRPymZ0QW69KcTFKEBSf
2oQF38viZJdQvbw9GZAMCIMJMs/XOM3fil3nntSjYV0SHEazBevOI5m2r9/jVPnv
LwQcVLYbXZ83uO5tXYFnUCUyG17nzaaAsSkvTAII7Z/cQTppvmbjJ9jC8RgLWH2f
kwgotG2CsKPwraBSCyMm9M68bGqfCSzaueqcBnOipEQNBRUkRzUsFGh9qjvekfNc
VosK6Up/VeG1ve5dXhGcNClrWVBen7hT7A2fU6b3kBbwNh/3P+diAa/yqWezRceL
nruMmsRky/ureCci480nwVwxNN2QKrlvWBme3IOupQl2AuzS0B1V8YQ/Sw6lTgrX
gZEx3ABRWljGrQmIKFuuXVACj/b/S52wXcNcCUUyiSyXfAiR+aXCcQ/DwzY/wMeC
+gLEFYpQOyU5f03XADVSQvq/5KTBiQMj6MTaQshnHZDxNO326rzNZIOe8ME6bU/I
rLHf6gBp4dk7FbXvnmIMhO2Wm2faekXbPpuNHtZ0qjWSHStEzb3z36WT5LyerGHN
XznbRxZoiP/AcQtdnCEOGR9flD4r+TaUOEf6jC/QL1Enohbhc/Sw4jxS9tX2ApZF
G7K+kp13lPYVSMWLv7r5Iz+GbDGO/O0HwGiPQj/6qxPOM5/Vjn2Zkdt2zxscssLh
JSUQfF16Uj5PcbHkZChTLecS6iSJK0ItJq5su5etncQuefpa26ZNKOc/NpORtPZY
KCOLIjqcJ1K9S3YfsEV/Yof0aJeSbAqPDVQ6TRoShPqDaJduuouz1r3w5WMXWooT
9vchWgtnNN1+I1gZl2G9Ce+IF5BeIVnb9xKo6cC/QIrlfTYQQ9ncbKbUO7gLhnjF
54htpABHAKQRGDdKrR4yhqiiB9Dy1iHnXGMCGmaj3ft0J9rueDi0d86hsY9W0rsA
+ViqTJ5qZvsq3nBIhwh2Xf10pwOWeRJPR/jdzkeAg/G7m3AB5znsqS9TQNYrRm0g
9L9Lm3xuWj+dw+s2dyO/OhxmAdw0mZZ5hu/3x0YMcZLscasWZRtwilceDB7nKxEi
lSIkD5nEkdA1v9+gHpzRTYAyCR8wkC5TpWbsNH2LHKxrYkZzbSNX1Q65SDtAFl17
PeHFPRU5QiKirD73BKFIP4JE8oeO+6nu4LuJCdKFB/lPrq+0fLUc982TjoRCpBSu
eFrJ+CDjNXmjsudTLMo2S6yvaLe+1oEQTrsUEiik9iiueulLmbCPrG5hKrSHrpHg
F7LtgwN2/J/4SW7Srn9biPz0HRgcYitKkedwr9r2wxAh60zaAStrnzw3fSg2eQRn
6FEfqVaxSEhhkPZvxLwHwVAdJLzknli72pICSmGqyXNqlwpJqBc/hOmsamRpc1of
u2wguT6QZ3LGIYdR8b1rO79Znu4JEGPELnv3No+PcnxojBcep1dZVGP2NKIKs1dH
+qH2QGtDzPqoC6kK8+J4NfYS16Wksnd9RS9AlTjEUgftpS6JmfKfF+SBbZ6/PdzP
EsS+w0wEnwwyJGeYDmy0XEb7tEHXw595YzKwKnL1DelyRPM1YnhEmwmnL7/L6V+V
u0PQGdK2bKYAEk2+I2rqEfJBEE/XBrY7cs2RA66QrEUXT8HQFz1fMnYi1cQbbdQP
XU9Nt2dfqW+y/nhqVkIi3TgkxaWCPR6qeZvAyUlTjGifEN8HZeyrS3R2dxW+Bal5
U/+zmApVg+4EOlaYPSkI5t/uPM+oEHat1TUwXCsuw6LjX5CTFqaExlwc0gdZ4ppZ
Wza4XQKOaypqYCxJg1UPq1ppZJ8Y4X3hEcYqUxF0QzIdCUMETeyalRHj4k1V5eTI
eLkD2fHmsTTkQUfSMnRjPEmt9m5DsUtjs1oIkA39p/McbXiydqH5nJBnnwnXayQ8
fNU/cRZijd5uUrmbqrcNra2dlnZct/b44+u5GCBJWtpyM34nR31jPhkm39LEHdSe
9W782orhLPNPVuTpsdHW1U3AUGUD9S0wRiaDoQ/D8inqT9lyGovhZYIE5sS33q5W
WKaRZwb/FhInW1qyRFr78btOLG3YWL4BeGx7IfdGS/u25HvD0HSa6fQhdNgvNaaO
h2b6LyUBv2SL2Zf3fDF/vDfLGalsz9vtLhB93rdysG2/f2ywaCZG/XgyAcdOXXLG
o9quoFyOSKTxvkZU2p5ZqF3GP/sf9y+KmEEpvC+V6uXAkY7RimUoyxd4iQovlGwQ
YG9mjxp1nNd0x7PHyMRneRCOJ6v6MtmpbB1wPtRVMzpLE2lkzCCh7H5AlONuv1es
XUx0bJvrV/4oJh1WYrbIVHHXHiqzGYKCdBj0vv/F7VbxkwdphQl2crmRwBtTXK5Y
ChmLzb0i0pngKVFsWax87+iYAQeyw2txdHyitNV1FEktZxOuKJkVZWLujknw6HHi
nzKX5wygP8m6wVB02+Xe+mgY9BjlVx84a+/IZPClex1RO2pjmvWo3YVwFOY9Wfvk
wZcWZda5AAwr6SdCGftjqX51buQLBUY2Z9YOh/VoWCNrcZy4/c5U3Lv0jekPzgt7
87eNxcBB69bJy8wADkdT/QHSk7m1+ykJgAp2tKsNBWKI18DWHWQSpedaYclzUj2M
7uEYOZyO2Y+bp9qKB9858QWKRmPeXX7/Xaq18wSEcVe3OGmqzSttmXSzS/RSv04+
R4723foAdppDKtT67A+UT7qn5vXip2xpYyetWz4g0omn21XP2YkcmBf5RAP9SqOR
jAAvXJe7tiguu86DFHj0JW5qEo4GFGLuAIUko2Atz5ueST4AQyieeA0onjqvA2WC
zY1ejlx5bVs+ivXsId+4rX4gEH3SKyrM7BHrzkHcOoxZ96zRUo+AwKWElMuSXsNF
/Y77kWlcOISQTsW2IOd4ryAtuyUjRCGy6FqnoDPdGEj64gip6+9WoLf/VXgHHZGW
6AbexZ3kmtcKOsUk9sr/TcieHbuHc+uke8qTH4etI6OlTVasW2JS0VKOL/rujJsU
bOMvfpKStLSTl1YWNuf2kp+CXicnHtfUPyNcnkGmm9Q1zLQHATrXaBKcs1XWMRWv
e2HouIjUuQq0UMeIVd9yjGXIql7cf9Q+yIkKLh2pM9TrMfwiqf62LGpS6m43HaIR
vuZR5CzGyPXlCuehnpFwDG+lHeF8lnPrklM5QoXreObvmZ6pHMUhYA2lXOm2Vb3x
lRpRLGcil5TLfJ85+HlogeqDcMEw+cI5iQr1KsiaGmKBMP+JC8Fc8CiQRyz6WKQ9
FYeYB3Qzho/cG3wEScwSd+ns9+FSZ6VXOMgzTMNOHw1i+wGNzIc61/82kxue3Pow
4tZDC4+XoB4UBHCPMGgTUjcdeadPKoZqsOEGBKMiXSuf4R2uOHnLpFTLMrA5Y8Vx
cOLj7yZAwi0T9vTn5iKdnyphhyysDgd02g1YXv/uxy96K6kWM3pGgW5zFppfIT/p
ulQbH8rN08ycvRcknecjCzPWoq2M39R1RElC6tHdLXyes5Y0vEZbUDtzVNsnvGBM
I94Srd4cmkg+mASZE7C9/z/wxJbmN1+XkJeBlNK6PuMu6aqUCwvuzWHNDahqLpjs
iDYGzMz30/Of6uPlXewp0rs+8EvNND6wT9Knt6UxdXvGbuOcINAU5XFmlJmr+903
an4//gbPUo7IPTBSCOUxkvdNSwr8JMrFferOtLOPy/NB9UDLrgqYL3ITibxlVQkU
4JxuLPhqn5Qh2AIUnw33Ye1yrtnbAgiN5vMGqPIic/XXvEsPKnM/pTMZKoS4GtsV
+wOL8fFyR7wT6SK1l/Khg/83H3W4avD1xF14y7qpfMvXIk6kNTDAQFOpP0I9Pc3k
dF8D4/36nbgB0dX+zVf2iBX41VRxH130S5L0J9P3NzSRJMk1HKVeOXdUa3XhqZsY
PwIV6fwRqVuWxugj7VjlflFTaR175jFFzUP/nUNe4WHAJ7fFWJhHVesLKX4ezfKN
oI5TCYUvl6JF0WvVv4QshMBVA2h6h3lVa3JsdXK6WQMeOzmJQNGJs+zTA0GF3Lgb
OWWsXP+rvU+5In7V9GnbovUpIYzs6mDNXlo+76/hhuSod6jGxI6WivMF+1jJ5o/K
T83XOFPtBkURLdwhBoCkkoQE4RjXTSlSCns6ZsyNdFltzxingq3TpKn3FPgII+SB
jfDcy4bEaRQpHhieXd1q67r8nXuNppTdpTtto8X9lo1CbKUU/z71+1xZc4QcSsiT
jQ2OJqE3oYfDIgS1gszlSabNiimqGL7RDipJNuX01JF2BRe0vSdX00ej9VCLp5Bw
gkgeHjvC5v6QWDEGNnvWpJjg0qiEdmNvASGHh5+NFmrJfl6RxyJirmm3I8XZY+iQ
lW1eTibABK7JrDfrx0WV3yzJdZp3fG+GKXJqBQjbuOxEXbo+EisX9e26ohvU/6ij
2TeI/5hlm7eAcXtGc4VDh1B7LtnYSIguyiFqFldbVjQp3byQX6FIDIwZylsTAuib
nuIqA4zHACxwfMeEAmCZ5DjdniIGdgkM1brAqPP/+zUOnvLu/FVUKtPSwbECps3F
6FgCYYV7sCorJrB0D7agbmoQOZmMl5Oa/u4Ob9g+Z+k9P/65nIJ26qraJuWbmJcK
8e0wNGcENnHj1MXmJ1cacpMJ/xDPaXx7jtPS+Da2iVBoxwytxj9CXouCr5xBDpym
b9VWRGU/KM/oyv9vEhdhZ1LYc3Km89OKnh9pOnsKmDs8YSMmn1GMABStP0f9cbWu
6uTeJzMmjpLikTDf4tYhszzRu4gAvWsQRx3NslaitLZrIqxirfaqVTd3z8LMYoVs
vA0PWm8MMcPtlI0HZOLAUCOgeeDT8jzOtUwAOjFyLeOi4RpSIBL/dHQXL59mbWDA
DRlhXcCrC9PfPZWW5CzsSJ/MTWGNhT+suZ9nbe1t2e0NpRYMelGwwU7CykrcuAib
faB2zad4VM+Xja/Z6PQ3TGLdo50l10JzwyJjLxasp1eYhG9dgjT+akYaNuH9j4AO
SKPuaH+avbavcJYpzTCu8CKLuJ6iZIygzU6li1eUGHwVcy4QH50PDCg81Eh/f4Q1
6XmSZteA5+QDO5V8yChX5k2LYfVxD3p8zeq4F7GsjetkgO2WPKqaytsza9lrPm1x
g/+2YXL+I1PDsZylKMBhO8+/4nazoIfqBgWqy9HKPZrHUmMdB7L0gTUbF7tKTMc1
ZfDLZbVNDM+H70Gdnrk2L7xR8m9pm7JiNlc/221Dg1B9sVfBw+TodlCkmx0giw1T
s9W1eo7UzeId20pAvGYT69DoJf3SZER1VkqM6BC6bDfqx7pQwIQr2aX9HgKTuVIx
NFQ9c6vpTNMwYhuCtQympCMUCarjijcIZViLQ6ZNc61+uU6VZK96FHJmktG9yqYh
vyI9ewnEUnh7EFokbf9v99KaVj3OdhZQpKVGUNv8eYL7Xd1xyj4mRZf15u51R5hT
jteK5pDVQr+dk0zZsN8lBTaAKc26uRQ/FUTMj/A/iPBu6F/1VorYbvsYbFXXIswk
Fk+WkSkfv4YZaERfuy2FOjmZrpF8miANaWpI4PIx9qPtAutNBhmRAaekTBZrzxhb
O75vqOSf/I2vyABxRY9bDNlarm8UL42l3gpgIrDKZgvEnTlkHGCi+Er0vpKfnvo7
UezIwoCdnZHsRmoQcpDTMrCZL9LrA8t/PCsQdiWqBSVm9UuxocZ8ykHckPLkaBSe
354UroNucKPcQtRNDtrOyUiddLjLB3Ouytl4qLwIFcUoLZUsM2lID+7FgHDugvbR
uniN/cMeK4drykUkPa1DmfiQT5loG3EzR3friYGpqXnIdISu7ZjSXL4cOntEhE8k
f86dKceMg9TSrKXDXBYznfdWggYijk+nAueQzzuozh0yfj2Bywii3JismKcTcKfU
JJK4PSHR+YZSxtaJxyFtUNxxM/1bv/uMHQCl+G3LmNnib6R1qi/lL+zpOYJ+1WQN
c87uDCKWp+R96Ka+AgzmOpTrYcu7aivcmDru+JV+PXAYUQ3UQHY3T+8SuD0MZ+ol
W2K61+1rfVmrHFJP4QCTXVrEAv+zHw2MdwqmcA7pGSO9duoTdQwmKIRVIy55k6hx
ID7vUbDuwbep4Qb/IGAIRqpP/6b1prjZRJ8Fi+6RbZxkp5Sfa9kSj6Umu3bfdUuV
+eY7fS/n6n8LCwqy0BxeFyF9GbhUyp0LGzb4EWoKlQEuMnCx28GPbyGuAHHDPEWA
GmieybNgB9fBFiXmpi+UQcLOYfH3e6Tm97BYQhgdnP0fFG6S0cJZXfYI2NdQL6YZ
sNF+BneZ9We/P/jfyeGJn/qSteedngK3FhYbLGRgeVy8qS3Vl663j5uMmfHgGV5F
h3hzX4lTtjVmTgSSzmwGshhy8cAGj+e3UnL9KFEmPZ8Tg8X6UMWbeJPpS3nVNWIM
EaWGCgm2wWDo9YSPF3yVEspDPlWhvzrjV/kujmxkkzC7xptGRqvrdwm25FRkyZq/
VEkl91jLdzQJDvSvsZxYso4Af8OXtaLvWKCbjI2/Rdz3UPz56gJxnr6m5q/CcmDa
N71WaZNPGeq8Q+jLdGYTVA5v5Z2w/WNA8YnM8pvL+eEO4xqmeZFg7WS0RWtJfJDJ
3JAOY82Dj382QsZifVFMVHB+RHlAHIFH0KQap5ai9jD6iZ6QVBwUmT8MGxcR1pV/
RtY88klQzmHPObdrBvNUxWuRwHLQwc+cVaYosaxHZDsK94myiDVhJ2LhSpGwAY5R
fc48wLC7aOjMQH2oc8y49KpmheLTHuaM29kdNf4lp/2ANbJmUflr0GPACON/7wdB
m2MRSWdUhV15kjfF84rWBjhXBj9VvWP+yLx2BGZN+hDeTbuu0LPolsJCQTD7ZCoC
qhcMQfEPOJvM+D6JtEjp7n2puKOwDtMI8FPZ3iGIGIjr9iz0sT0zAjEQk+0IcbqC
jiJN97xBk+cSuzkF5q+dpe5Uwo6/VyaJ+RPcsyT/zyb77aTfLnxdwnGeucUGFUf+
dDb4JSnD0OKBkP6l7tM/aOcf2294KgwRnOhrMgXZisVH7IXFA4yiDSu5VHh38gGY
vwZkPIEzzeRQqgHYA5NSm20ZYKh5nkp79df52RVsqk2fFcm4pMQdu7yq8pyf+V9b
pleS5GzYKNCAoKSMHsYPDOSVxlwqORtsIEyUVkCYX0kNjTwqXqWxwfJ+FvHgboNk
CJ/QS0RC4pvreqHj+gZK0ylXE2aXX8A1EoEN3KvdQeC4lhT6ZanF1uOPpJmOYeF9
Xn6zPqiye5nUxkdoJUflrZb5GCtcpw2HaINeILY+ZEslrzLnr5WvFiL9ynC9+VSj
P3KAh/6KDSkCDZr7VulVvM3sAwTHov9idz0uAVlI5XlWtLMNLWvIpuYhqmx54lFj
otmfV7u03VExLf+FqeFmWt29MB8LQhm9yQ9jL5XUzqu+llLsYnj4iIRTcKecOWnl
cxDHr19eZFplWFnRcppnai46TC2G3beXMTuSi/7Mgb/kmCBHWhmHfvddTwtZW0Ox
YvVpCouWFlztVXjdfux51casYv2gK8Xp3Fn+C8dMM5ubui5MS2jc8phpEm+k/VGg
06RL6vTJYbpexcas19I8w+6UH0HDU1ikcQM8Y4GVLoaZQTAe5FWUV+dCFQOnygLu
o/Cuq74HEDwfgoxfXBF5KO5J1ST1aoIR4nmysB+TbqYRcuLvNdhCCyjuM5HRjAwx
d0JmnjL3/lZbQNVANd8tGFJhKPMjs7T9HBCLiuK/ONf1P3/iItapL3OFztNuQV7o
JF5KX+FYg7xj1BDaxr4uWx5ypR0DL89Pi2tj6PofUWaCGPso456Rw9CWDbAopFH2
zLwgEGVT4LkaEgdxEvkQfuVzDBeBvMiZ2AJB0he+E7PF+rxOFREGuuFJuMtItQZ8
0Iq3Kj4pq0kDxQ/aI3fuV/3CLiVms77opia4hQWahpSXrdY/xsEPyXOfXAMFLv87
lGh1L/XVtHH04ST9ltnaBkdZqf+8JxM1sJsJaxSH7fn38EGVReP+VQNUApLU+l8L
Kw33fIspDc4EA3NR2/nBnLACn31TRcN2OLs2DfmPPWtQApuQIbsjVwozspAXHJ8x
e3Irn8EVM2xzTm6aGWgKt5R+X3lMFQg2AsOOB3q9s6B9+28F/X7dNeR2cjJ/eIS9
8LamYlrkDW24egyaOwR1Q1j4+AOrLF5yKbHUF7UIHyX2wcPEMZsbb+m2WY9OzR2l
UIsyHvb2zOcyzhszvBF2+JI90pO5lRYY1uz5x5HaEWqAa1mWuxSCpdPGR04gDvCJ
OXLlqvMa4FCh2a0sSRw1EcxWEhRs9AMFP9xl2f6iiWja+AsHtc1JRQZXAMzDrW5D
x1mEZfiEg9RW+UMLdGu61jcYrX2R3SnpkC+7Id+L1D8YEBd2tkz+1kA+WSlnOLIO
70AGS3RJR3DKYo/YijwbxDdl/ahDzWhgmiDjAdV7HUVPt184ugeYRumJVas1jHGm
9dgjwt8j+6OIseZMUfCaLBQzJM/j+lbzZiFsm9zNv4QAKZ3j8e5DDVEBPuCpmzS1
vn9sme3MTi8qk1VBkt5uKcA1apFj5OP7DLf7q7gk8bXoICLew5Jjllz0eCijW6qB
TOUT7ZqwTk0jeqbiauotwW+Qi94X3rSo7l2J2oyoA53hNTQkGUWFA+lnKujK+1T9
zv2TVKwK1SNJmeomkdZdnMbc1w7RQ3axGUfCHQCfcjO7w82IssT2UvDq05TVU0+R
V1ZW3F4d/uIJnjx5CdzKaRiR1epTO2Uo8kJ2U0vhfxQxcDujtYmbQ+e8xzC67yUw
ZW3Y1ne30ytQ/48/hUccq8Z/mkG9s3IEgG9fujRBZZugdiGiuDmvRvrL7PlzbBT/
tU07aiTEC+o6mE+MHWSAVf6+g5aIlcCO5vHOdHY/4KolTBas5fjtU8mznBWHwxX1
wJNlD6gYeb5s/kvPBn08vmLZ8cRe1/xxSpao6OhxCTxc2PUnPhpt5RNPIo3CgyMw
iddZ46ihx+UsZm5gCQNouCiwD9OWRBRPzzN+n8naBr1jHAudT4lAaW+E+wQCRGHa
wD4PcLLk5h20cASazZlD+R000KAy0fTswF+IkgSbJaoZK13VASYrKdJio+2NSMXv
v0jyiGKuaSSgVSE/xQPG+zalVk+L4udGYgW9og5XcaV31Szw7tfj/UO0xOhhXkUs
NLPS4jcxlsVBH106msf9RMZ+9rMhvY2tfcxuRpfmYbbVR+kWAAaANS/BWHyQiAp7
T3SntsI0SisfAPy7UD11Ie7kKKe7LrMplEtBUy7F+7JLXLOBCZ8UUAcHcFGfldgT
1gnjgz+sAi6HikLsntvdmeqrizS7OWJX10m+RrP9INt/IGsGPUjsX/P/9ZpSqd7u
7DSkeq+p4+yAgp+ryrltLecOpiP5q11AfqMtVpXZNpNS/T/Zygi5KZYNIhh/LKCI
xxP+gaidgnCit9xrWKO2cwcooc/NF4rJWo7wx4DXYi/+zG1HDcOBnXirVvdOVIMz
Kr5VIOOWfGTUUVKfQV1qHghNcRe6NhSsEO4mHgyCX/JiZ/PwgiBaaei3oBtQ7VRQ
rYJYuPm6cyxyLMCqBxLZInGzJBW2HHUdsyLUBHcR858v9+JFl32ZWLje/9s8t4pL
engCTQ1gqyX1EP3ckwXZSwbguj874pZFf4+1OISLDz+SkHtUTggEklFb4YMtrkWm
VRGElBa8B5UJFuP3BTiuxBhfnKdDDPsFdphT0xJs/B1RmRtucWA6ejLR8mXYzEAh
aUbYNa81TQ5c2H9vd60iF+yUXAkIba1zuCwg+462xk8tIu6P8c3HFq8zjRQ2W9sy
R0C+RkK4JsTG7IcMQC06JxgNeS6QQfI6o21lIW8JxsaqyDNb3SAW+/7mxd8nRpwX
01N2FUAw2JedIZfWcqZ13WSMj0cWdLgHaI/0wPLKwp0MrUWdk/b/V9zFzTZGZbZB
Xn9rBMfXtrlMapOs5j3apYq0TH/WoIem7IW0TXodjWXFZarqEWvZhdK6vNCoe2I7
kR2NS8kZSkhzOL1FJX0dqewC7vFPkPJit3ia48eLTV8mWvpakCFUgDQaLbwMsYn3
hru/1wj/IxXyI1FF52qqQhQBsik3HKL2TnWHNZKR2UcQ3o7z3dW6rtIKauBZGpnw
0hJEWouDSPeMcYDiOnSnTcDMpNx6+2rpiq1kmOPeC7Y2lHeThhuUikaD7JzAZiZu
otpudEJxao3/4lofswBtU85WLzPsTFTphGCgY+8Z4tZxf+em75MPm6SHZ4YfejEj
1KcrfybDQa0dCoX+6JDn1CebOORnfYvgIeeWCYknDQECVWmiyL2jIAVM5nrHP8R1
YPk0pl5qyzRHv1FnfkkAQthgKcRQy7HWcB5xaMRlgk1jCmd6eg7AxH2r6P0KSvui
URIFo9/PMYJDROIIL9lguqXMxQMvFukULtFsGkjTn/LI3uFxG+OM9T3zjBXNuWQv
pbSJjZkpJSbSFEExl2+n9SDtC+qLpgo7Szd8oymTsMeuUIOCGIVVsN59/2uPiz3E
WoTfYOTO82nAjfitcmeRKVwOI2CHF26Lbv8tFd7Mf5n30Ne00Pu7qwnd7dWQZVYx
X7iO8vYvfEoONDw6Em9SlTT/iEFb8B5EK5oD7iQPbb9Wah0bVqXZMz2rCxtEzBC8
z70+ofjZ7mAkARvWblPyhzA2/NmISlzqEzPgVVc7cUZCer1i8ewSlnWz3wsWPSY4
9/G8cMYRCMgLtBjl2xQsHbilEcwTsLF/E6dRhY+qoUpppNEVG5dcxysL4Nini21B
KsfE8WolUoeitmcmOY9b30tux2SD1kiUDi5IT7WuRe8i8Q/OtIL1MGdbuk9r0Kbh
kHbgVCziofjialdpftVJpFVVnTEscYEJEcEwUB2pv2YZY/++sDuDFK3Ch0LK5vuZ
B6YB/krzR/GcQT9R7ix2OeFWbRseK9inRoUehCcIP/KUjdaMO9F1JKXo/zg8j16B
6w8BaETJSr4UEdUnkytAjYZCk5MbXKuTKTC037l2dc+P09kyfHBUlkx8j4q7tQZu
AV30F2DWNxDorsBAdyv48vyjGddXNmasLRpkuce7VZWaXIgBvjlXIuKV915f6+fn
EYNYX25EUomRCQgZCSctaXtGqBX5wnoM8X0vSu56cw9oMCmw5tedpwf4adSrZBAz
MVU+Assh4UkTBC/xEzCEpJQ5pLxgVOhHWQVRL/1muyKAHx3J+a8BGhrVCGEaU2vH
KLpmn6dcQJy0e03ZBtsBwILK7NXjmWuI/10zNUORnpoGNKdp+bIQiu35El5nhqIV
2JS8UCQ3iuBC5zr92e0L0ndJGVMhn7fOG8JDZLL41EgbsMGgG9gIKHUv02DAMk5F
5xV63U6StUrtosrNsfo8Fo0dwJbltLGg5L7iRQstOawT/BOi+MAoLzhGllPnVXjV
ekrPGq0PBaHpW6z3yPhABWIOYu8FN+7K/uUhd7qsnUJoo2MzbVk8uZOEG7RdnzEF
WMYuNsfG/i8Yzn7XYeEBRV7vY2wmFYeTP05EA6juTUrDdqLWf/DO5H3HIC4y20C7
Gl0yuDJy+AzXToRpooN68mIf73c/BQ3N/VkutEgJnKPXimPGDrMuXb8MebFnO+20
SSosDC2fKP957sdmd2q0K7JfkCFC4bAoekQENMDPmJ2d/nurFhHtp75abgpJXH2O
nal9ZEKEkypGM5Hl6QMI5z39lJ2RnpEX3xnnXrfJd2MPDqv49GbqOo23fKmQvB+H
bmZ2bAd/uwcgVEN1lw/5rprJ8Gz9uvyUX74VdUePZ4anVyJbyFODw3lUU/yLIm5V
/cH1RmstMb74hEFGCQ15Sh9GZoOHzJssYEFjqXEkim/QgxgutaatW+ICr3XgTOBU
dqvGCjomd5eVe2P/rkTDmN2fs4G5XJ4o4Omztwhf8BDTNUum41WRwm2SmS8B1p8U
OzF1MekbldFmh6AXhpnFUtA9WJT8EQlj7vIKE3DOsCDqK1/BHFQM4HFrUzlzWeqo
e0x5kRpyKGiy2xS3+hS4JBsexGMxJjEvoHvT/kyp3XuaoBFSe3+SCtwY6XgcTRmp
w8taOGRavyxgyPYsPZjvba1S0yBKPq8nALDivgzMYg6nw74pT8Wdw07m/CzslJg3
00Y8tl33W3+U9gnk1+YYSl91niYRL0CymR8bj/jY0yQiKOpj0aVZ1iQQQ7CBc9zS
tv/CHcB689OuA3pZVYKCOG3yOyTfvPjgKYsFTXjArpVC4bpTsLqQaeZVMzr48MJY
Fk+dHgTTY4AZGryxr+cqvdOEDyGIkdX27qNI+nn5+HAIL/YaErZSpk7IfdDCD6Y1
2ZfdtUc0dk1ElmtJcTjcPd7taPRrYpQDHS7qhAVhwBwjHtNPmW+64tOVtDlwvtCB
UVBOtlKkttlrKdjX8fhy9ec6qkYvKBG1aZ9lH6lBU+Pk2iuQ6t9YXPUoJ0VvtvKM
PhR8W0ok/6PjFfeDgRKxAmFePp1KFCuilcdRbIjDeexuIwBMyNSUm9r8egMdsyiR
sYmejSApVlm9+4uVwwDUzY9pmTb91cQ4jyB0YWF6EI6HuzHi12PiIZSvdmoFIFCf
zrkzxm5KhLWQ7izJZni5zQ31rlo3mPKW9Psm4tfR33Bj8ylVNedGsLUtJe11ByxS
NJhFPhnJdNbnnlo7MSoP41Fj9Ys73llDJYCtC3gGn4CPozF3ED4B5AdJLE/+1Oe7
Mv9bS+sE5AiM7QTyTbLi+ZPNPmhlTFdU+3r+ZImlOiDp01a1Zr5r6HRO7bD+252B
snQirorZSMZtEOP70yMZBqfblyN97KMg2Wio+2z7O9Nqq1Xb0ecWo7ZevfS2sAkk
5gAZnNyTdO2nhDBxK6LFQvs99KowoeP/qe21yILLUMw52nTWTVDYIMXwmHXkcAzv
1Nd87DKqmwnhJSzfy/knfK3hoV2pFPyW+AxIslW1stlxVysK8YOjOkksnGens/G5
9Uj5YL3XQd94sH/Okgk55ufgtgOkr4V5ImLZ0bN0g7LnqEdWamFzkHKqWX/sZKqU
c0Cf3vQbh+rHvzkmdCmn5CV8aVi7w8A955fpYu6S/PzCDkL8RCTVxZQkNTkpMVnB
crgMKhD9HHs6suZAofDZ6928sKleLrEhYPMCm2e5v88qwfXhIOF/P+cgsWnLMESH
FmQJ01wR69FBYup3TK9Klwc+pFZQue6w/mQTgn6sKWr14rewoPnyBm7roikvu2x9
r6C4UlLHtO3yDIspCYQzBwX4ava5fc+6n3aX1AnTXqXWB/kZcgUIjwOnCjuMitRA
M+NE8MGuQb8ozha6OxR20SHBFpoFxoyNjWfscXDJKk3cM5IC7ep3+p+3IhdlIpdF
3Vm0kKs2LGTzLVpi3QDmGf/RimQbOkd9IDSWQcnuERSPDAAXdafyPjsSRdlmrmBP
sx5/yEjlruZoUSl7dlWiC1Ykx/pxxZmOFJN7ZhSxWBcqfewZE2bCVF2ffWAqyODa
Mz85VpGRo6W7ZyTw2gIhPhErsvQ5qJWUn47TWze09tzV8eJFMaBOYYwW4ofdw6cd
yhVx5PQuD2mzXl381V9ugtQTdz2g4GjwyJTA1/aYd/5P+4ot7ExLCyCzqI1aV+f9
L/oduL4M96PpD+reNa5yEgiwTVR7q+ZLIw2EzMTbj7cVXRH03Nbsj7ILeDr1gKrH
sUPGWbVM63QC3Sfc9XpZPsLe96FKbDukAYFY4YcEWd5AgeM/0CyQk96nsMmZXxBS
mIurJQUeW9tM29s/wl1e9ZSZiUOdh0z0wefzW0dM6A5fCmpwXDdnxP3JC1dah1by
FRwlJiK5l5v3uF/gvp4I2tSv2LENXAvx1FPtlZdaGFpWRqifS3BofC9DWqJk5yJt
8+NInd2ws/4/ZVSYvCHw5Qlfclte3Bv/L7UDxD3AJeOo5Ky/tdS2FOH1jjV2nAzs
KFaRH6/mKaJETDBwtJek1LvFjhyMOjjThakXSeZVbbQbbK7MmZr9JQIzZ8GPr9IQ
B5rVc18koPOn8rCF4EtT/xIQ5tzIrL4L9rDhGwamhaTG+OKBElJPnMcUeSMjOjsQ
IXWbLMrgxXNN8x5iDPW1jDc6eA23HS48B6wg5oKLf8b9uDH6PGbYwp5GnCq9K3DS
IM4urOHDDKE/vec5FGOzBVQlMO8CHfJTinQZN2wIP5U8v/P+iaBqJLbB4ooKr7pf
wwCVojZQ7LKtAw0cQzjPDPdm2I3iShQOADhDWyeHN2IgCpT8tLQHXNs2ZhOtSwk0
7SpyplzqCLNkLgBPjQwPcZHInNUBL55ikAT5pf60LBJqJBMnSKFOJCxBNHfs/Vv9
Lr6eodX45dHwAHYYvnF1jebOVgOGAqiBT08IFTMCMdVO/HP4Ifv4ij7YIUhYXdsz
Kxw39KKdjKgWbQZR7RFuBHsaIZ4mKlj0V625j1xRAgIajtwN9ve38StgS6RW9PKY
S16utjYLNddD+Zh7kW2jEtWaiTCFp76UovFmkoCqUBFXGw2ATjJ8GqZYD10RtxGz
hqsV/QW2GAaqF9m1YLgZR1GbGX48HVqQHeL9aqyQgKisKpiLCACVLqOWahxiHOAh
7X47+XonjId0GdCD4wEdD4H4isNF7U0m+PBnTyG232FWp2VpSRAEiXNn6+vmn7lI
7HjcmDivTcebuVGNA+MAHGVvB9gQD+/MxJx91Q+o79bCsf28r9PULGROCWlWil0W
/fdzypLVdLGSM3GLL4v6B2Te83UnOg+UJyjfHyv8Tz1IsznmtwoZeR63Kl9U4S1T
Wy8wjKMyzeHKfw4M8SlBq6tiu2GHqNVdMzQYV53PAgmKv2EMh9t7+LHTwjkEIgR6
T3b2CvMqTG42xBxZbkFEsLPgO46mPTIyS/NBXLyHYJTBuiHVE4n+k0Q5wqKAkkGu
UkX71SBSElvNhFjHkynt82DnUtpqcJQ+cyK+AIjXmQYkJMJba6r236Qfu8wYlkPE
0X0d76n+ZJPd3b0pfLxHrJAM7C1Wdx+NjQbofT2d+3gqra8itnSFXMfXCIKiDv8F
IKqMW1IxTzkIgJMDiphsBURfDRruJo7bgtKSZBivz5T4kczMjPb7brUCuuxO32k4
xsGlxRXHQX+VErupkGHie2+wFHxoteZQudHuNHdNP8O23Yfph5ivwu1ksDOt6xSs
io+jazPm7gcMehzq+lh2frVHmTZY0MbJIKqpo7A19fNjrEzBG+OD0jf4wDUX+ELo
hnoAKUNVmcp0S+TllufIQjt4ajLmKCxzT+f49Fi9rVMEPoFCtl02MexLxIt+3+ZT
yJ1jaYzjNYarPSpcXWodJ/lpuZL5/EWvBXVw2vyvEYmFhWCNQosXZ7Miod/F4M0D
tgbxsVhOAvam1I/SZe3L7sHISmnldAwAh87JLXjE7hzYZnFV4sHc0xAiP7U1Gm9O
/D/RIdgt6BnKGXkNJR1Nws3gPfoZOg9qMKB72pBZEuaVjtOA/j5pfofzGotYnVj6
J6sHDyCvzETfqR6JKo9Fy7HCFm0VNJ/jw7Rdy8g3f5rc23k9/y3LoCvQCV1vVO01
F73nauWDgv3Nv5MDZWS8AdinnPjgN/KUuP1y7nYTn729WvtvESGhOZ6GLh/mKQ2S
IIHtgJ3e9DGsLI2T+kyEYyHtGIbRJiRSbFp/HPp+aurBBhbt6y8UEpXXOqFNZuXG
jKS7d1XAXxKSnm8Kgnp5OfBMeNYVHv8m6aOSkfm7ZMUn6uQrNL543Rops8WHY2Wg
buyaqEcGJMP0MTXvZ/swgQM2Us2uqniNahm3HEQg95DLymg9AiCZjzyiHb5+kDzD
7qXAcm2bGCQ9G3iYstaz7sim4m0PIXX3Dv5GxgX7FI8jVL2XCx4THY8bXw7igot1
kWLwrriyagc3Ii1bEsYdwehWsO/usVB9KUbRWsdQQUozQtMgWsuTWUZXkW5gAKRc
PoCWWHSXfuWd8NEcaE/AfAhOikx6YLfUS+ZJiF8JSUKc8FYEsnP4623nifVC3Kg0
PHXcOyPA7lJErP+0j7Mf+j1xmzGP4mCxX7E72rC3biFQCQ9gGvjxa0lUka110mM/
g8iLyZdFR0HjlS1On6Z53Wnr7HkKycyBeC7GiC5sR2O9kf15ymV8usmP/KuHuEAR
5PS0OCYjNol1o278pfgCna+HVVvz3m+WhyFYgW2wN51uTbIBwiImYnzo4w/rtRzr
qHlGo6/b8xjIzgJ0ggqWOqcih1ulJPiO6I1A3/Brmd86SCkELxHxL2wVDiTs4PDJ
3hf1bRXbRZF7oP848CbqeiarRqCXHU6XD702hR0wlEAoXDpvpnVRsH7aL4Nf5sN+
C/S0QYKzlo0p4eJAxw6G3VPPtQSiqDp1kq2Zx+qqcXrdNLib/9JiFUKypQj6P6Wf
SVoN3r7eI/WoxKXKZ9XzYppZtTp2KypidP467jZ0YeBvGBBkeT+niUAyQr0IZ52R
3Bf8yij+x7R95cN+48t8/SZAyfF/p8fqDrvb4GBUhjfm7S4MJEi9951LR0l1kR4x
62i6p0YZmhEzG6oFoBXL904ijqucShg0sIo2rWHtCW8cgp9r1ihpPJg1WpV2siF/
woo7LlvK2Ie/f4NGoNbfotujo9nN8wUFUezvydA4HUOf/1XB5/5ConGeYKC78D7U
0+JzOz/kMo2+vXH9QRQ0UsozX7ixZOXUvibA5mZmvd6pi7bx09nidaAfqpPsTF1l
W+k4SPclnm/61XdyWz9qqQ3ludsd+xKLg+PTMBOu62N0TJakuZQ0jYDs2C6dA2dq
H4vGw3hRyy+FRBlONM+s1nig+5W9v4bB/qUKZmdAkKF88G4AlB+WsstecquZwtsG
5uaHY+/WkwGthFITUwsBBGJt+aVdFQqMldujVmiehuvrLXBKXt1XVD/akM2dlQk/
uIKwSGcqE1Kks1UxSOgCfOeeI9WKYS9h1ZeDLrpUGrEiREVfr5JrPFZcubwVM/t2
HcGR/SiWBsCK8DeLn/tmL69r+DGigrK8ag+7Z9BQ/Vio67ihOFUreO8UmScLd6ds
fupnsn7UoomO76N7TVE//KwkELWYkUpuBSEJrnjW8yNn7ExYLl7qOt6tx/llZo2g
bOZpBlktP4iX9Oa1rwrqL6u3hCl8dm0Oi8zLFZsNHQhh1yiZIr0pBp1fFRn2O1Ht
b2muEouS96OcbNSCVMO/kSxIMOdSDT3a2KjWMVTKdG5/8BMmzemnSRGyFPg6/lew
2CeuoIiaMzA7UkWzSUBr/HHF1AhstiNfTGYbWYZ33Mm9rdHDh3zCOGpG2jnX+nRf
uwDJm64xxtVB2lWHp3rm4zGlyxX0Cd/nD5w8XfAwMTTAFmgfpIzQlcbItg0zlL89
eWgk/Nt2XYnmK/fu7U8Chl+vVC/qGFSLt/49rliMnm/BASfT9t5dBiYq4diKHu5L
5jVgKXRZqWwHzbHn5HBSOkFSvkMlqCKOZ38nRNAKnPBPB4sXBTspylJ6QmwdnKjz
OXRr1efBb0sVIbkmM6VxEq7rbTX4pDBs53mSDqr3jPV/vhXwnwaVgLv6gi/SDqkS
mEad/L6WApbCvQTmgufWSzRRt7+n0ij6KWvvBAHMJm5wy9rzTmG42a8sSt/SGNfH
w1dx8OYbMBCPz2ISQDr1PkKfRikveo8cUTn7Srr3bT7SwbT6+5kfw0ho05W8Bd6j
2SB7OA/euJZ/KYmRDRrwqNY2dq9G2qFqEDryut8TuC6/jozHc+wwvjxddNemu5rf
geHwJTQx/kqbLP2xxzz8T22mndOUb3ACpZm6+CRubHP6jwaBAg+SschyveS+ltUY
rc4+mC99U/jLzNH4Goh/BFRK6ZYuHfwrA0p8APQJMFikPvjQxY8Q0e8VsR3RjD7A
fujfJ3WUpz/CetEY/GaYmobg4pQJCpmSHopZW7+JGnGMvsKHZMBTBvn9RCLFDQgM
G5kstlne0ALSxJUOJXr2CFTcZLBNe9MkZSIaVjrJF/Mdttepks3yAybGef3zv84V
DcbO6gzzUw5tIC3gtxxstKU936kizXbC1wuIF9/lakhL7xE8jVXNRjRvjF62h+Ly
Ox7J14frEzNCtBcgVp3dn6XgB7X/pqkwo1o/9/phbjR0GXdOtUpaoulk7j2PzEIp
jpdE3enbDH/neVdEDbRb3/FWqRyUxX6kjKi6nKaHByUJ21OH+ozt9nXUrZDK5Qu5
WxgPWJJSS1Fg9IVOy6zoK1X1varaesAuV9vzwD5LUNuY8QAV9G9qnRdV9DP+82js
1vwUaYJJeGy5FxJllfSbn5wVbrQMdWuVzueIKpqNTsUz685SaShPUZYzxibQvKDa
jYidocXqeu1E6TTCThJ4ZdrsZ289kx1G8Mi6rPoPxa8K8fSFvYG3DucPmRo4gMDP
qjbbqgpoLiJyY9BtYs+/jIZ2yUlULBgsZZpzHFM1RAxQg0qOSp84DpLfOzt4Q7/8
pomu2fsEdd12hm0XhJ2gAco05i1WR7kPknCfJZVC9too7hrxGLlkSyGLcc5xwHKe
AhIiRG23KQDqQlyJloEH3oU8E8qZKfwaXxxvxQb0DjHTMfmdd1qmDVn61rM7C0LO
R7iuv0qr1G3OJlT4CaQMYPvDnjqKFtmp8uc3BBmngBOgVZzWQ7+z5/7SAJjWSjU8
FcYUbTxTt5ukAOwniGISDOT6GXkvXu7jaxJfTOnFrF6ufrAIYokSe62UIVmPMhxH
9ZmcKaZkQzRqeMPbhzRaaam8DXW0zD02/YUim64t0G1F5NcU4ygCnBLuOgRIFqF3
auzjSCLjosWDlojmrwPMiZQXb4dAu8BeHqRCrliNX1awf3EKnND+ncIcUVu9lPpc
eiQmW5aaQ6rMwJiQ3QMjwLOpuGuHuR2XFnqEsijUqdbWQ3XSKJ0BKfEuPBui0HQe
ZIL8KIKz8bpxif4D6fSgmt1ZhsweoO+aLejkab7YRNg5o7Ng8dW8Yj/wpU6eDYNZ
8wI3XxjKvVNiZJO9nfQZrlrRy16V7FdNe0RE4tFlDRAFoHDXzRl3mh0P50GmmKfU
fypBL2OOOg/FSyg/j8pE5sZQWgD6t8MMRZ9ywIoBU9wm19Po2ildoB+9kdVQdd0m
2arfvB5P1YlNWl2QJCwTacEIMRRomEtuimv9KztLizeiCRBFSzaZJ4E8ukQnYVtG
dlygp1qo91eQVuleJoTo+/a0f9gPh5CuBeaPFJClDpTeV+dEWTTrls7jsx5ICxFT
X2zprtBAf7fjhezDPLAPgBNt0QSkoK3s51S1Xrz1uoCPOim2O2JeU1jN3YAXsbjS
oYTW+kSAf58OT7P3aIA37m8S1y6tzsLP5s8TDyWKrYFRdJ/flX/QVBJ2f9CKa692
jvAtNLoe7COPWLDtj5T+P3ZtDN7mwlUp/rsHsvIvY4qwc+BBL0EdlYx68vF14mfi
SCrN+9pXPDJ8KT/BNIz1y0tc1aV2HbhjsEbcVJQJA1PVb1KWi/jXmV0IvM7DisJj
WJLwAkwgUfJcapRRgt30qG3U7Pcjblg8misqjJlrLfKOn2IHqCy79ywmhQ8mFobK
NvE+FgOz4lloGzML8ZAbpInlvmIp7QnI4taBhVaVx4KL4I4jlvv008AlZ9LFQiP0
vgPsCd+cVzYceTtlvvdJlftc+JufPe5NHSx53fwwgIrdh3t586x42f2FvGiuc9Nk
Kl3xHiTzYQmCZWnhHZnEZVCL5dzkLsEPafekhkXf8jVwVbyd7pFi4IsmK0hTs6tR
rPYC+6hlAE5TfAdfcUlHwzcvo90ZzhH/D3Z/YB4CNCDbp0mMZwgF0QhYdNFKrImm
6laEBtnpxtLC+2BP3nvImbjxQX/CXgzuiHKx5PKV8vcfoHFbEMv2Pn5gZ3pVdNLS
p79NfySJJxHRRNeVqQcRjmVnipiAHVDqWMvgzT5L987SzsmKSFuP0ILlVobo1vr5
0SCiDoC+iXT+EH+7ddWET0RylV/5qs4VGIJvrs9kTx5lNlGxGDOUcCuOnnCinHjS
8aEoIIXN8zjvcojaTogB1uVoJ68HY+OFpn6GsW9QSR6qmXDa9hoa+QyAU1RWQbcA
GYGzrhLm0ZHYR89Bw0uALjJ/KxW7qREtdWmmE3inUhSOMRGgBmYLmDQfaSjV0+V+
y34VaW9y3sYcFgYDnevFZlCwzc4zDG019o7XpbUmlcIG84k4u/fEBQQ3Sqvi11X8
3fGclsVm7ooBC1Q5pEERgdEJA/j1yDTai12P2TKvGHHmT04bGgje9DpNn1AFCRC4
7ic12O+RuTnZXZgK63KJTGn5ortU/kl64us6NCzdjF2nKUI4KVMrtcRnoUTtUsqb
LRDZb9fIRUCtbHkSp5TDWCa67Arr1GVpZDFsaB36zxyS+CYdTki8uZu6aljA4+jw
5cQ+KqgT7+JIIBSCcQAPRyv9PbiiTjseW4Wueh75/JKmeq05CWvI9PCbLzLiHSYK
+a3ePaJG5Porf5W8h6j33gFQkqem3Lwc/uX5K2A9NBC8Je+wafwVUGqC0teV3yGM
N+g9oYcNAknc5G7KZ6m0vgbEZ7E0kAdEfeBUM5Xv3mfj00hTIT5vBtOwXF+y6ZHq
e5RD0IUrL6n9JPVWRy4qZfQoSLhfGPuuf5yEkbDSboYv512lJT7rtXEKTQmYLQjI
B0HSsBntbJsgvczTyHIAxeZ2XRXywoxgB/HDJ16He0W0Rk0QFvx2GCd2COmOqq60
f7pSHvhTVTgrotmFHbartchx1ESHBj0lR5MNj/O/OcrwUvqmlYXS+8gEQDq9Z1bP
bi9ODKZ18Gj9ErGOwnTIZ+b2eAuoli670GBp1CYZVgphH44c9rwAVxbm9xaJJDFM
whIoKejrxGZuSJZhCy/nlqgRGwgZuaw6vIjElPpumt4EUY0GW8jEVmOgNkB0kYgr
3JbPfcvyK5VUiEJWe7W6W209C0+RflKDALtb1bFicLj5s5oMhjtEe6j9eMR2/Rmn
1ehwQM12WSF3AR7DSAOgNcvpuoUV4bstq05bcxy53ZwLDAJ43A5XMTn0PtqKYUkF
Dklt+t+z5QtQLN3qoefN95nlI32pL4tZvxVTkHvpwV8y1pExe/Ij3nCIHDTnXhOt
pdcl+uwkDUxrvPL8J0XYOYJdhECMc9Zp9x3IqNDG9NEW4BPuEX0cu/4FwQ+7WX8u
oMVsw3Cg52lGymDhUIYs5CXn1CBL7UfLQ+F9saBEtQgdEWqb9qg7o9HvwuK0heQt
kaFAPW0P09ddXFb9/C2JnEuJSzkJPp/jSS2gXSPDv7s/HjdjtsFcLbvkVKugwFgO
lXU3uCeX7hzb69B1H985ADzUC/yH+BhuYjHbhne9x7UzMFUsB858SOmhkDEato+4
bHHGkiCotmDshk2+X5QDElPbiQGk+91/T4YlvyOHG8+jnh/yLLohp1udZpgKOiHL
oJJl4clJfXbeV0+aigjOycW1hUTavhquWZh0p0hB/6+9GITXJ9qSTXUdu8m1D1h8
YFCiyg2MxusaUT6mYCG18QC8Lm6/DwyUKyO4OG0EUfQ1csUMdKzzwXlP4eyKMxBJ
aE4k0dpzJxyMT7wH0ycTEwLWszd7zPlSICEop71ubh7nb7nM2rjofKqoPCTRxs0f
QA+9QIM9V0BimIU5BJ3j3Ha6w+xgUqgJSTlhTl4C305OyvXjK2ijLmMTzCFW1fzK
UTValydIWQu3uxRfJC1xZNw6qgz8rOFDb2r+EHnIm7pJfHNSEv5JpJRmN3K9Q1+4
bKTFy9qH0Hqhx6jce4+OzovDr/uugRd4Rz13s1pFhGx+fcL2tUnCr4nhdDrtw47/
rIfYxscG6950OscCwmW6f2gJczlaZCpm4YiAv7GK+hcuF+tokkfDE1WXUAmIacGe
W4GWYbqpzx6sfJKaJ26UebbteerPaUIOQpkglnDshQw0IZUsCbyH8e8A8WOA9P4P
9twhPR9G+DLdj5Svm9vRnlYQwABFURO29SwMpOUZSeZwXS9iJH/08eoXMM2XLgqm
ARwAqdKr5bI3t5hZSLe3K/vKF3EKC4+k0MhmfZaxqQ66vurlwq73RQksNeTT3G8u
HALXX6TAZFXotAQFQDqyWTxpvqZJZLbJLoLq+0f2B7/wpayj6VnoVNoFnMXIWBbP
WYMvemE3p7qU/whtUW8KC4qG8IDWbBZwF8hSDx+YEjVJ09hQ8xND5QqE+E7iDWYx
Afcq0XNJv0OQwe6GvFOHPvyGdSndU4eZ5VzQSzKixtJw7dCeavCf5hvUegIq8RRa
2WbBaHAlObKk9z2Rwa1JN4qZTgBM0pSih+BJQNooz0eUcM7gdtQsW230cRZCPlE+
VX5r+81c9H4yXr6l1POfxBedHp89Cx8mwjhAGuTMJ8U6XTstasJrUv3Y+qeXAVE8
QjqIdke3aSKDuSRS4a5DLzmkfNAW9Gke4+7D4nirb3vU0hqM0AseJE/N4m5L4RBg
1qD9L965RKSQWy/GDL47ubV3XFrpL7O+SOMPBgflC23Ty/XRHcxpi7hE4j0basEb
GKWphrW/wO2pi1Po6Z0akYKyYwizf9wqsnSsTyBPqb6P+dAKPdik2iyyt0f+SO6w
9DwfE/pU2z/rZ8Zy4NPRIXTx1dvMy/vHOeZIBJMGLIHUB6Db1fCIAZCiNzrJFX7z
OmiaGMhT/iJJRPh4hE5diE5vh2sym3app7svBAlYaYtIv6A5cIfmUPneWrbm3vSN
ArOqRX/jtdwFIVGt2sfekEs7eRpU3S115v8K4D6pKABhDy/kDyqFMGNkf4dUza/U
TlCKePSmyRrYgJXBIsdsenPHqNzHu8ukxJ3QOAzrsAkgGHlIcxqu2DnIxwbMtYMI
TB7rXoaxpmqRMjabVJVq+8aFpM7WDHIGnPQlpre4Sdy0edqoBdBeFKXQmmJFmX14
f43tkZVnQ0YMdcLCv9WNR17JzYykZgOi3UEk9/m95xr1t2cPdEkS8eAZoQj0v+o+
Duy4bc5AXr8OweiifTAMr4bzhx5RtQUYM7UL/XYEsK07XnZPiybRw6Mk8kxrt/li
dgv0CfXTcn2JSjqTwag+6ofekbAFdVggaX8ne8CkzD/JOibODSJVyq6Ky/ZXftYw
22yUfUVzzo+gmIpL//3H7weIbkE+mTk0krYkCugjDMmBBfXMoZQPHRraN9/1g6IT
OXVY4596TpLEzwKo1kxS5KzHaCWKvmdihbvtYvitCbv2P35CZTi+8+8Q4xqgzR3r
wkIOnCjaqXvUy9mUkhKaQy24GDsd+Vuo645JKrWPPwWUvEJVG7NxU69rrDH5nrzO
0NYXiSIiza4xurGVDFBo2BEF0aF1AWzwxSNA+6Ai6YUQ52Bnzksnr3NJKn2IymN7
hlf/ZNH4BaPuMQvuDue90L6azvXarpKhiagtuUm4KxuLcQrtXMNgRkaP6V3PSQ/d
qIM2PdOSdCKO4EED0jxj1qBfQKZU/TCc6HwaIwHjW2a/Jxc9ksjzgw2+MpKeIkJR
/6AbmvG84gtIM7d3N8GWkFVnTDRwUa2h3eDDTOAYuY3G02Ojglq54XYgR0Nzdimw
78mx/eWIYX/TGteA7Eirvlc4/gFPvrQnfqI7w9MWQFaU40gGVZ/lsyZSP9qKXLr1
smn1Twgq1AjwMhPTotpay6OA0MXh5LeYgZ+GBY3UXfmrzUxnV6dbbrSZnShy+wGU
4DBH4eHTkBO1hpTaNzewV41PPoZsJi6YNVZegRfcOKgT7SaapA8AItrVuWMstZHI
/6/uTJ3VCI3x6HoDc+NETUyDQ98OQzLUDYIHjxKcJXTjOMIaWdCK8QAlPxcfl8WE
pzM+Yfid4gLvHbNftJDVRxc+phhJInxjfn/4oXCmXtrKU5hPu+gCLUa814OPzb0N
J5LsAqGycK4WT0zPoBPH2dMKEHZgVs1i+yVu0VpXgw1N3wqhTJWWbuD2acqcm+HG
kLolQvC8SvCxU52SqOE4vGfwbIj2OelSEcB+xcOOOgMBZOnZY1h9ayYMNqKC3gwU
Ysw8v4jOmEF1tol4K+bz30qlLCs+YYBDr6+smM5bpzbcD47VzXt4ufDg13l0WEr/
C5x6B/7CD3ssh3XhF6ytIi3SjK9m+16Ys1YF1woC6J0ajCxleMfFITQTCVtBoCvr
IyBPCldwPRiVAz3+411UjOESJnUf6Tg0L/tv5ADkJTuc4vDIcBC7p2tW756tlIEZ
ATVq1zZU1EC0S19cDM+kOmg5ZQV4cCVhKECOOpvYP+jXHHX7RKIJKHDDn3Qw83iu
8eGdGJMybw8i57AQ38RaWo8k+rH5ZJaI0R+pP4QbmB/VGdtXOIliibclB/DRsszc
JD3iBUkejRdruKhUkuwVSXQa9BQTLAGnVWiaugOiWCHBLN7Tc7l1xnJ3LXZBNs+H
LOMm/R+T1DRb3SK5VuVxDwSbd83d2FFc9XDKGyLTf9WQ9YHsaep1kBBUy6d0SAF3
QbwwmEDEJu26Ch5kvWQMifq6vau36CoGMft42bt4MV6GkBJkpP0tar64FTJ6Ufuq
7lGutoBs2myeF1uFjwY7xVyM8MCZUStDQpl/2ogzC9rjyjn2XQWs1yJfFYOAdOXq
PpzyO7PycbguMkQ4VeOZPuA2zApHMLZp/GRFMq+/3f6Cf+2JjivG1U9XnEiZIAmn
hgE8hjg+AembJ8CcSyF1/cFW7QNDodYSwF+fWmO5bZ1exXM1i2MIr2Td/fBRVxUO
umhw/waQ4Tqt8T0G9BwBHsxXkE+YJgtNbgz159v/1j69XLqg7LwwOrFlLzGgLECp
ZcDaXZXJmzXRjlzPF2uS/Wha5VUOUZaBvAjhFwMYngUiA2Q5wsugTR+Q+lAQs0Ri
/X3VEa2m0sSorQaWJUiGbAbiw5CQeBW/creKcy2LnSMfAt/QLeTF33zcDgMd5o5k
tISAQTBwZiajDlUvvpJHyLObj+yz1WyhO9uhSjCbDOulBdvuSDMGAAT1S7sthUVQ
SUxELy13afgrjPXrzYM7Hu9QAyS0dPVCPbQiNxnSMhTg4UGPpyjcJxXA2w8vKRhE
aCRKIas4J9BeysetKTUWJXovXVkXe/V+K+053x/QcqH3v9yPCrn2ilLKo0oedrsJ
II3CB6YYaK16lNiCpo+oKQAfuIgQqbyiTCK7eR0UOP17ktBx/geEU6kVxjuaIPPm
tuQJGpwnW0Tlwb5Ds/FGaGOw2QzqDAhXmZCsV295RnnWotGK4Ag4sMcFByDujBd5
ImsO6Moms9p54q+gshZsH2AzRwqeUrMCFnCWKIc/WFuADnzrzYRRI9KfpSTHlr8r
x7H6y0TJFhQtZYljIEHK/eilSWaMUJo9MBtEb52vgZMEhhMymuoAmG1d7oHMr+Xu
HRSV4IPlJl17k72agrVEYkD9CI5Tgw4eoTkhkheuChHWBeRMX1rCcxlNmyQKWOvT
SaVdpRE5d8xpegKq5jI3lniPsCBHUs9j7jZ8Bo9Yy0YkmdG+NtpeKxB1ebjZ9Zb1
S/NxmRvm/OxAxwb/IPf17KyhS2j8giV9TSfjWzrId4xwnlq0LlbwyU6mcFolSD5h
iGgL8wimBj6FZwzz3Pz5/O4AmrG45GraBFmPPgBBY62ypjEplZkDAxE9Gc2jjN5q
pBHqD4jtM44RdqZjGj9SyL/lymE5wbDusUIU1hHhLObBDpQ+U4eau8l+cs0utPgR
gjI9qCfxkLBEhELOT7ufq/mmBIqbQ4SxAN62UjfPn2k8oABxtNq59oGwOYesOWyZ
gw5kTwhosC/r7B93NKFQ30D01zkb3dDLNifDl/XW55uL8knYuBATl58BppasdaKI
w676sW+FmUInQEQezRv+wS3NheGXaVYowRyWEoSkR6Y26GlF7s/pN614Y92xsbzP
8PNHn8l2roTDZOOJcVIlCNzvPeZBfU8qeuoM9FKcfz2RrMWDJotLEyE5a8JXKK6p
rwXU0ERvWdXJgsawau0rcvMPTHPu6dMzNDoYpytv3cN9Y7vh1Tu5At5JlciGOtVy
ujFXVPg3HrOrGgoE258+ry3JDanGgk9H012fjKF2CqeFvKc6HcGnmY6fGt55gEv4
+blgXDRYwcaAavsfMQnwb7otQlFN32VdPKxiRAFwWuG/H0L6RqXBExv1V345nJff
SIATXQfjIdVcu2hnHfEM+16QsLW6FusWEHTWcJgl0BnUQO5foCrzic/zfaIU79aA
FuL5FSh8xNPe6AIX09srUgkf+5dOKMlqHmYnBApGHmwLmK1AUX2l/aDrzH///LjS
22MpUHfR2KUeaZVK5SmKWC3qDLiZRqhXvbbZcHMMH5C5+tmJtjnUjvsR46BpIp0p
awJHlrxiaNYkqEtAZZBksv/Le3I7C4DZrzIh58dK9sYoqeobqsu6Hr1KX9m4N7h6
EXfRMc7LRyDTqy6XsjqHZRDIa8yE9KCCOkl+GoCrGVBSoyBtih22kcaByhz3ImIK
se7/ZT5wda9qFas35rTvGQGudtMVAPcbna+SDdEEkRPf9yaeKj45cKvAr7GuTUUo
o9bNjfy51RnsGWFhpD5Cww4XBDxtYk2AmmxvBeVESrfGgWawdxkMkRsX8n+aD2cI
tfRhp1E18UudNsjOvM32Ti8gX51tH7Q41jPSBWz9HJ45koOa7on0Cpy62RpoCGlE
T1ZSyzTTrYOXzJYfZJGTpjl8LLcK2h0gFQkCMBIH2h6c56ptayz5StZjrsjh2PSp
6/n4TwqkPiMVcmXlet2mD9BuGwvqjSEYKcPjgrevqaqjFNbI87JjOyN0lI40o3aj
2YVyQJfuwZzcS/A+yQsqyP77hXHGMzN1qXa1RUXohnT8zrluzbjpPaYrXivLxH+g
Z/H47x4za9UuKk5CrPZSbHa869Rs5MfAspYkU+3BpvVrwPd62r7ZEBfPj/VYUaSY
nvTJ6V29aC334PtyBosMZtEBNG3uATYoNtzseyoM6Cl2qzZ3A+bSeXe27cwAGQPC
onFTi3HL3n9JdvSN2D2rz9hWIxXLJUGk3uUXk/W5ru35rxSwryaBu8kvRPakvuxA
fFe+XIuWHxAAOTSrXlW6B549EwAA3LgOBL2R1A/X01/lRBf74R23CovAmfCAqIhD
ceKujsxRU0GwPEohScQrDmKWEZnqfZfM/1QLejpdFVdpl0VeVMdpqBpEwEfz77Rp
UIMiV+c93gc1gDoFmryXYl8u7k00lShBh1l3Mbs7kjr4bYeDjzoKcNBmtEwput2N
XqMWhTk1MUiwKxBuqbRW/2Q+IccwwC/0VeMcVHRLPIXU/SgE5ofm6LOOySdT5GPk
Ie1PyvifnVAB0uZA5K95CZuVFlaWWHMbvxM3j7WXm7akIkknBh8QhDwMwfbaRiR1
wIbOwlvXyErpXIDV+He92KV2qsZFp5X0g/HhCZoOH9YPP9Xf/zW2GuEPJB/YQbot
X5otVXkYcGJaR9jgdI2ttqfyalZnj82bQktMliIhPD53wLwD/Zh6jAGlYkTrel+n
yaWoSZWDb2BRizV+hX9SsvrM6JWWhmlybC1nGBIzT2cGyPr94YVSXsJCiJsDlXWC
OerFAFCoGXbQHD6J9+yey5e2/mjawlN9iP5oLQCZijnJLOjh+EkeJkWqW46QwCQI
omNXEWhmNT3Ey1juToUIgAnbmTRsVzXBp6sUKEmGWGGq6wXnL65e3U0bqpdzZ3Po
M7UuZlC+oSVk/q2J7DcCt/Gf6+w10yDv3lFRHLH9I/FYAj430zFqTWyaGjfcg81k
XFHVjabS6n3Mc5P45yyNUqtuCBgP2QHBI6c5o4aNMNC3DlyBT34GOrFcGV75m4B9
5VCcewvjPQipM5qibVMAmAT6b3gD1eqWgdKc4eaybfGT1KqYqQtRkIwn1kH1jMHi
5msTyr4BYQveDk/8l9t7oChR58tpGPynHk7+yXrvCPG7K4H0L+F9ymX7YnsfcSmT
LxKMG9mG/azRPxKS1UGV2my21jaYcHTgpwEmXUc0iQipT37S80DAVP/jEIZ4kx5q
BKrgcrYwsCciybadD1bGjJQqtVqoIJvia7XASi9WFUiHlNAui24V4iXWg2/TgF4b
g3zGAePvS1VXouY6qVovdIXChIDBP5ki6m4ppCMakOcwtdaOVj3klrVZDQLAbSIz
yI7V4vPrv1O0VyiE6GPi8M4d0dYSkxOpomOm6iWJlyJ49F6yfW2upc1u4LQXT4+D
3wlABt2Af31zIqax8LO4TZ3AxonNeFjWOUJ0awnU8d9I8WdNL3SpWMtyqorPLakm
aTl91OP47oYa48rOsopuphM71yjPCn0yU/+2py7Wgt4IFIienyEhs+PdDnYLa6K2
EyXNy2pKov5YGxhjDoPFHNIMJ9SpZZcsqqZh9AW0bOG1uICf2fq+eENWi91LdDho
Ps9ZEpEZOiLAz4FAFN9BP6RtU6kwQwR3n35MSr16LPWn7bPssU/MoQoerKiAStzy
wR7z7zKtxYgfMaOjvHTKxAP6nkYphfW1K0ueEm7yiBQjdKmtIvf2cwnhlMZZNIFI
EANWuHBWSVSyxI3iRO2ifHq2ydnk7EGEwOzZmpNaaCgP3dBYONlfmXfqbQUQLCvh
uhJtt9emVcG60Bl9xPMJZIRLT7bO9WM70PbQF271gQH/wgAXWlaCszu/cnB418Dj
s9UC8a2QXYgzOosu3gCCgNiJP/IoGbQXVUX9s06xB3oSOQUZjYiZ83oPICiRIGGK
ga6D8s/jbL6G1cbDStH15Q08IRKWoyYcJjeSkRGgNZzb7RyKK7Z1fiS9vFYzSjvm
xUOkPvN+yOK9Iny01VwpO1Xtk+k3lVubXoR3x9njND8WvBO/B5wfG60myEEfjqvG
NnRVinQD3jMONKqIUTuV7z5P5iYMTaJ5wa3KeAm0U/C6S2gwfURTP/2m+KQ9uUug
HhTx1KvNK0c569XKPyN6FKgkWDgXiztbHShJFIT9QO8jPv19hDIhnHPeTerjuSgM
OStp2uOUwLT0UBbhprmwr1cGGDc3Q634L87QZo/01u5EmDG8s/qNeu7Gzqz9Q5CS
J4h4gOEpJAbnMhtiyxBzqmHtz2eSxhu8a1Fjoilj7tyf4yHUkuGse+HTpbkHJtgd
jE+3aMqVy9LMIDSOdJDbWVyLn6d5EGFV/cWcIRJNGkjnnSmJt2UmqJotd6TsaLSu
Y/8LSJrCtL0E7fYU1bfBsPjZNOITAmVkIYKhkK16Mizq7CNnMmvftt9QoiGjk9os
SQyFVIG+MYXIOrFcmBqp9s8BqHoZfNmq1vs98vfZ0KOUyWwNmXDOYgoyg9hq7lV2
Vl7FpHfuEXlkDPt2NtlDsHwGbO/fzejAsr86S+R9bGJrBiQap4A7psYR4Xznjsi7
eYdYajlxL25l7RjRkduRfHw+v2mTjVRHUUn+f4u9XPZPHNHKkbTpV+fRtNYKz/EM
Y+fOa5chnmnJV9j+RYv/WG/iac8M0HNzkIzDRf7dRYhaYezoMjBeWsYTxttjYHWm
YJaozmXRMjUgPI0El1/E1yk2sGQtJJv3dNgMU+WZGZ+SYXdpiVNVHpWZ5vrGBUQF
s61Brih6bVGd2nCvvcm+anBWIvFKcXKetStB66KqzG5hD+aOOhy560ZTSF08iPs4
KATdMKgEq9OVI6ta7JqheybFY0hLXdqjTrt5CPp32dP+Omg3jodD3iStMYxr9xHJ
SZI5kgEw6mtcrEqzo8IZZPpEUIGdqw3TY7ZtQ70nOgOCYddeRtY169k5Az/d9KuE
Au6vz86DmURMfwygoXj1Uz1LDKxMw4AJleUh99tkL2C9KSzLDIvTcpWouN/eT941
5IhROzCa7jkS98IYk6bz2GrkIldpaLo3BpE08ymelO6snMEqYcraZp94qGrE8PgL
hagNcIeYscxK2dMF8W2wWwrE9Dw5fgo8+e/FdPv5ZoifNJ9+x8huK+6ebNaxUQCF
0HwvQ5DflbuHOk7r9QGuRr43/EDHyFJMS/hrfIM42k79holHav54pV7jE2FuTDx8
JH2z70V2R/c7CWfgj5eeEfTbsaQzg68/cUTRHXYZY2vLHgxlitECP3XohlbXdTKq
nm8gr0z+Jd1fkFDp/nZ3Eamaa0BuzpwvAxoyLEFE/Szp9uvRhLuAmMQM9ZCn3a6A
nfTE6RdJvm0H/uoZd4zJBWNsJ9gehtAZnDwSaIBeTj9MTlEVlIQse+Npza0btPPf
DHNw2g/iSJwoOblrs/kFybaFJGCzNWEF8HiJXopto5uqm8OIP9Vzl58FISV9xUwD
m5OxGhBvf4PZXWh8RqIjAN7ZSjGXBqtfynaBfFEggEerGird4FQIkxsMhSpTCnXb
h31WuegitlAkobu9bkiydW3OPyeAHhEP49NqYKVAG/qeQrU8XkyIt0ZJTpJWSCo9
Xzl4EQmeEYSTWJEfcP5Naug4BNMI4W3Mc0Uaz1JcIKMKOqHWXTdnWTvWOMUj58zf
ZKld8b/WKAfJfeiC5RyAYk2ig8REwug14PSFAOFQE22LCvQBJ9+EGrG586mRckv/
41y026wKS7bZ8d2oOU4A5vzZ8sTtRkf0IBwRlbqazBJV3/gKkY7NwhMeAyeuCBVk
DLVa7UdAwNL3msHLmsjySGRpc9qenhkARwOB0xq5TAb+2H6mfy70xkYriROw/GjD
nQNH3AL0duX4CvTrPrRaJScHOwyESHGxBtLqlfkgDxamvOanarGF/tm4JAsL2Auv
g/hWhtTGzUdV9tCoEpq2qaXR/6KS5XTDnZtnD8zUFdTnyTNiW/M7b07HEav4hVod
BrX5Umj9GorCzXBGB211HhwGRy/RBcK3+/8iVIeW9HZLuxLkDf5TpiVFVCH17wQ2
+tDWGLN+bigOt1HEUCyDTeiWA+FAKSJ9VU0K6TPxGIw+bZznQaP1zlCIz0ijs3nj
SAThN4qC9GpJhRkXSr6CoDbtcBvXnerw++I99pouAtUEdOyUp5cWSipviC7Z/wsV
e4CeH9hA7c6Jp8tayc57/QlyYDoei8OoYAscWeOq+hlwQ0swtSfR1+fyXHExe7yJ
RQn31HNE6WpnvVdeDIp8DDHfjRwRX/xvyUK/Zex8BMI6bJTPCV4DraUtwaXoZW4S
bjef+cv20kabRuX1ap6JG8FPUUWqfFML8jRi1nppfmMTtjYgdopL922a6E1Cy+Xu
c69sE2hQBTI/3f98WPfcSY3ska2irar86absDDVnXEexPS+UUJeumyyXCBXbJcHH
zujhVpyTek85xJi83tPj99K+07cnTYM44fNqVH5xeaeXMUTGnMADciESs3Z+aYTF
5g3/Wq09R4jD8kAZeCOUwCE8Ea+GjDcVa+7Lq454M36f5lIGVFNq0r+EmLEiqw1r
MTpJzVmHbm4gfUWOr/P5goMnyGFp+hX/AtS8rbDUV34iMpI8Hf+96SE9HqywBE5p
kCngrVsTWPuCMz83Tfi+Q3PceAtB8YKuiHjPTDScVxHizGKVuq2vDSYl9uOcTLYj
fP0pRybjwGqm7Wc1ItnFzXbAmF0sUqTXwqrNPAICtPo9tYZZQpj/xN3AJe3/cy9B
CiV8bh+UtfabABo64N02qAkaw3TGLWc2S0Lo7KJbUzaSbz2STxGrKDsQeDs+2P+g
LFxQ4cmpzViPCUO/HKjrgzq6t1TddduEviyZG41RhkcE211scxYB826HAPp9Ay3E
5SELw6XqYS+WlHHsoDJFw+8dq74Oa8BlrLxFjSCEiLQnVZmP16tY1iTsdvRhyZhm
QEBJk0lbqMi4u7i5M5V55ZoqaKmRKBa92IRx1DHLTW7GlfoamSc4ZIyCWTPHvIPK
QOEjypgwWbIOFTJ9L+yf+a7wWmLiD6G5Nj2Hk/RXk7Z9tjx34R7SsJc4e9YVUlJU
D5tMbuPfmTKpo9Hc7unvvQH2N4SxXmsKzSBsOxLaeny/StYfcaGS66Ox5Bo2/8F8
lwWYb597qZtAWFJBBABwE3pGcoqQlcMfyuymiFpo5liKwwl/Ay5aNanWI5+3j9xI
zEt7Lk9VNquEXzxbuwuIeLFw5/CsvCTCZDG1oRftpPgNjWp/fIxHkRuULmppFXMQ
u/9hkzdTRheNdTvlr0h5Omc4abbKIpXSZbDbD8gyrADDl1eUOMHbD0fUZv+zVb4n
Ln3/3pAse/zICWk8gkp05viqFPqnBwoc+4yHHwRozg5406OtX9H7W78XPqTaGbXL
nWrKw1i5opEpEt9zFn4WWSVteiRStlzRTtWM9/Dr2ekW80hNlwlfRQh2DjKhbGQN
82JlvOnFqkH5rTONA7Tub7+Yj0lIlfAwlJb6RsECA1dxeaVFQdrOJhhvEYpNl8PE
jM0NqIjh0vpBMfGFsW3unTi4N3ZZIU4ZEx2VTUozAmoZ3ic243zPiudx6ucJ7xaD
ywIcAqMISsmq8qxN0nqpPHA2Cr07v6xE51Hb1xcnoFx4+Ip8KNYHcKG5d2fmkSsX
jdNDzHKae1PbQkRDc0znxE0QB1iW2q8Ovcz24UfwHuHQr6M6czKBzcBm8d5jsQ4Q
ytM6d7E5o3UXpGfeajsfEveTBF6fJ4L4QA7C/AHCL1gs7UhZvZBR37BJNbbny2kA
ZEVnSO2YEYmm4q6UlygkAocYjuboLP8vFYBAHIsMglcrFujmTyzx5uh1th0z4OEJ
8LTv0ITgaeviRmAbMaZGUYd3jF79FbGZed8vXP1zUYf1nGGGaHvQjFBVtmv53k9i
jgWjvDS4fULoAMmPdEuy8WpRndoTJsHiW3YKs+GWXsbkPhq8f/migp2UlymIUBgT
HY2kY0smNzcsA13/k6c6yq+oj5YdLX0W8KE+0bOHpScbX+2OeEnKMP28IT1/a1IH
9pFnY5cPc8G0nBcDhx3vn7Z6FJ657MYIOg+/8EoqWsKk61tnhlr8d58tQitJ7YSz
plAi4NyH+P9H8DyBn40Xy7aIJKTReuIeFV230ujkAkRB0wdMcPhy8B67sZh1taHC
/nDVkg4evW6skEsEN4/iBYy/L8sIR1Ax3VqoJv4iFB4Eovk2gUUk1TYYUTRO8Sen
W8QObiU5VNvChGrTpAfjvOb69U40P2RUsPXktZWrWqloq/MoYQEfhNOCAH47ChlJ
TxbWTR12ZiCGZFmqG5gN3LgWBCyvmyrF2lww0TxUuM9oTgnPHADG62bEQmm+XcE+
VC1GQEtB3e/pvwgifRqWKWUbnuMLQpZ58C6zrvPzBSLpWy5d0608YdYzQDINh7+b
LIkDOZ49dXw87ArONVp/onE2GPdtpcBhkFnDIg4MWCvIwTVcMPHvU13zwkS5Uz9B
YuPjPybtL6LxT9N+CKTNcHW5MaXwQUaA7j7w5fmHgcdeMKXJoT1MxQqDRn3yhI+J
8gyranpXvcBErtonsclzAbYQfexh05u1V1AC9u6i5I2FbhvnZ8hABxdODr8q9lw1
36AaRu1FKR4/jJBTct8lPsNhaJ1/xro44GvqZIe6KDurDlvYUXVxCpKcipq768Hr
8XPgG7xrwGRuvtHewDqptBz9uj0PTQj/4leT9SNIYyD3CXge1091lSP5AnDNHzRJ
lHeejYc2icAaNnTnXydjMlSShK1M9jGv2dtlgvbXBuMogxKQuoaEDRb20g+GvP+N
iAk0LxSukhLTj1gPf2UiA3aCS7zpAlfIFRLz8Ly6XK2SCf+XuFAvcJiEQTSQQ6A4
BlFOn4nPR2L+eKh3kVwQTBOWEUBrHkP/Vp4I1lSzZShxHr987owCb+rat5Rup7P5
vnVfcw2IZmf3QGkxTVNgxHjtEcUzVdKzY3rxl0cn0EjL1zXYQgwFMzwC9seITOaW
t0sDE+DKozOVc3ZvVzPgebQMKlNHZW1LKBZJV9Jh/W+/ObJwcIDuutLALxjQG4GN
WNaczq046IKI0LrxyEkKztdKUAYNbkedrTEMBFGpfbWXaG0iDE55IpUr7Ww7xnH1
yCGzDfKwqKNQfQBYQ/9qIjoRh0e3+uOACydPIJt8sGdd1FRna/T/A7WRjRN+seJC
9kIQxya1E65/4SeM9zNvoXtgkMuu+fsNe9VT7R9InXhemLIc2l67dgnDqEP1g3km
Nvn/9ZBDvRDaIk3Pzjz6SB7fyMGNuaAXnE3iXnAJOXk3gF5UmX2UxbyOZ8Yoq7d6
lkTxT0NFMnRHKlEOq0ExjXWvpl2jRfV31kOTNsr+K1YqkPR0VHtoPb7z0EHtgk7G
gf6ffifci4+zVGTq935SAAhdyDj1aSJHCm7ewKmNHBDG9XwZKAXqf237NFWF5OBz
4cpKppQiEDK+GAfDtBrYL7/oK96EwXv7hh9+IlE8PRKARFuROUIS9kpMsV0X3GBT
vQ3M2r+UiyLOJ9YRb9IlisTVjcBYGNtn/0dPT8PFbborM2bnwjbfThuFvmh1DKhY
9Ah2MIc56iPhH2oTvJGCiEJZRusN0vddWfYhINRRpe9WGa+UHlRiqmz7J4yYzUAg
wz3mSOzw35G+67fSv7Eb0zd9NiJed464qtIReGgQXRk07lQe4WUpb15mJCzchiUu
cHWCeXrbB9wcO6HrrllJyk571ODewSkLVdWKGYQKerFaGmN5p/FfAENGR2/yzSGS
zEGoLAHH5+hICQ3mOzczsPQ9pBhncLTiSqPbZJ6CDIvXo1mUggDPBO8fDkfpJg8C
UhR82FR1lvK07Y5cmPjOu+JUZ9+N/zo69wzc2OTKnQad0yeeeEMwivTynNdmXnl/
YLIxoZvD/HpCINHSJ8JShaFAfMkiFnAQZAFPitqP1fvm48qxgVJJhd53Fmxs7ZBU
n0dqe0R/C+zq1r46D2ZIOhhQ/Qc7y8bP4tY0VR/TIPr9vBdNK9OpddznoHI85+GE
oO2I5REZDuISD9BS5mg53aKTbdoP/6wtANs/5fL1sOddTvBu8LKv60u+n5a3/mOF
2o2qlwUS5lLk8lrfUutDOQyOh7chZWXnfh0HhAow9NTRhvUAY8nBqS8ye+S9QY/J
EjpscDlm68R69UDJsKf4wBiK0FVHXOOz+I9FJpRjgDW4VnvUCffuxKQ1MRwZe5FK
U+UlRgdtgWQu6jm7J8UIRbvXvgtsDBLufJb+pHNvwGzglbFaC60fZGcUbRxJfb95
kBOgICtOFYsJ0/fkZX/JCQSyrqdcQsSnPGKv684kDsWIf58ufb99WnWIIAo0y065
PGWTPK++oBRK4I1Gvo8AdTItJJfwhi9OODakpaDtnvyhH4I/IDNeTpvT0RmS88Ys
aPlqWwkN3TJ0FyrB/LO2mc6k5BiZ1aGvoB1fQiABpGZklzBhsMVTS6dNnBiSU/ps
LWAFJM6mCY9bYAbTs0h7yN2arXb8wVhFusHRCVTnHbKuMEy+XROuH4FHonj/ffhW
LgoXp0BYdXc5TfBQikWrWse3T9EHEmj1Ey3wk31kB7eKbHlegZkJ9TP+3aPTKjXj
6MjqGaWFwfitCN/UfK6r8mT2KV4LETQOp7se4bfnkLbMeiG9cSFv4iZYHh4PqHQ3
GNuN7ByyTe+/jGghkl6L6tuD22MP+g4rCf001gnIMq43nVgfTjeLRAZ8QCdRaPPf
qNXrqLBTUsqvjI59N/wn+9P7Nu4sEKC5dE8a9P+Q+uyZoY5a3m4RxyBNem7Aoeg0
PRWIp1Rf3aiZ9Gv4NHhSI6mJvZML0eOjSMOPaLFlsUIGnmyzuVKHK9POLAuUEcIq
PpgSh7SVUcwXu4by46TaprvFQJ3KFWNRM1Te+tHCYfzvzTNYQWc37Z+5wi5LJWNX
+n/G1M/JqkrfwzaCAVQXM2/z7sUa9hTeqj6gasrJXGbmMUrzXp9/T9x1BcHLzpmz
Ev/UKqjdwKMuZMGsxGkSvA4L1JdEUUN/3vSL6ipfKXBHAz3wmFL4GvrDD4S+9lvM
e8FnQif9cenvNpXj52FmQypXEhyvzM2RexPmBqxAyjKohy6/D7n8JSHHE4grO5Bw
DupzMyT3fPIC5nhZvKw5n6fpB8gaKaEhGptW9Ojj+ZzMCel+5VofFI4CNLgbBzo4
FBVxg8hD0diqdQYOspfua1UY9GPmS1dHzIUL0k8csibn+JKZQv3UP8QJu31ZeLw3
2tLAthUgAAobEm3zKxLbwB0e8nI9jVQVD3AorqSo6/p++5bPqTbMPXYY7/5OzpYq
wK75AUn+6G8217dVgKwgv/0BNZIgZIxrKU7RgcoKQe48T5cG1aYp11C3NAHXbHVK
jXpaOEcTvI6F0akOZVs9U2W7Bl5dDrWZmXWj2ZeDLFjEqHBhkuAUeSYaB+KaNtlD
mUYs2JeI092xfTQQMoTAjETAcpw1jSHcE9G9mg3L7mRnweUdthWZIOE8qd/ojfhJ
Y4OHE1XnvKPE7U4VI4TiNhaXH1WWHS9gAxIqsHQm9hApAmaFMA7L56WHMgWLc6V2
OoHSCiQKwEeWR2KenN8RMakfF5qjJ/ghTqS03rR5Vq2iZwArZojOiZVKA1LLa8eG
6kHy7KoAETRooL8lJy20jrGRqiyfDWDbLtn3kfpm7YOX3LvIJmy2zpBKf+A8iwHb
Gg/gAniFkcKmlIvCPkC+0YIy/krJ+67MEr6jA+TYLvHQjESaTihCSB7lUTNIKFYA
suXOSEw1OUwn3mc8fZ+Z8IolabzxOTsR8/zKEfP1wKw4SpLZBxQLlvi2dUxhpaYv
SiwoE5XEPMl+1NYQZlbTF3jWkPIWu4AB5dgpQXgfEj9XVTFY06dlwOKhgIHpKlS9
GT30r18lV49oqPdWRwaVBE5g5RdLFqH4lXUKuKSOfRaeTdE7YEqhVdJYpa5/SXwD
R2QlT5Upx/u0utgy5F3IG5aDosteuvXp913Qoy2z3FWtsPzUEKqm9MUP2IWnyLo7
2bgL+xcrWUTW790JKBQIhs4yZNB2OkEpKtN9QryPW3XYft1Bdm133MgvYLmA+FF8
weOrdapCrT2MmjPg5BrZAPyL6kEnydZ6W/FLdMMmB/5kv3WFVce8tDZD6C2xGN9S
w3g5awBtCm7PpxJKclITvlTowIOiTgHWBgt1fXLKs5vDgisepqXhy1rlPIs3+QXY
m1A+9w9ZhCMmGzr35/FOzJqNAZ7AYPx7SU2wPanLHTQ8ALyiHBXB+iYeUzIvKFay
DYF1+iaLxI/EFmqdG+g2/5/3vbgm8/EjjF4G7yMNpn9ypyE3oL/JWxq5gGAKI0EZ
99nlltMZRcmPP5+DSvGYMgXQRirY0aCWGXxaXY9/OP4NCUGWBrCJvbr9vQ+X1ivd
A19B4JwBVw9DkFJsRLZxyUA3Z6ismzLSi3viK/AiYpBRoKu0N7Bov0mAMjOwziRt
z9mMb1Wzp04hi20rrdimGdJiyMssCpUZhsAYXC3r3Dey+1kOuDDfUdSOnzJ0tsaP
7BDVs6SEaZ4m3CcIU4EJtn3w8kN+NJkAcmRowRi97iOwZie62wM4AAkr0KvXYbic
y1pjFK44/JFYVvQ+L1tnqy2ZFOQJ6hxdk/XdCfRJt8fxmYx1g75H4Z9hywvVSqRy
PzAIyq7PS6wv065bWcpCdhhOF/pMo0G3VSdQms1CpqQIZ5ScYIQ/pSubqyRMVItz
Qh5WgbYZVTycgvBC2IAVw8r+aujuK2wMfvdpfm3URCioitkxSwwJgJS0c8eGGiJo
O1fx4Qt6nSj3cZvXjaYXeYQP5hqSZz2nAYYTvBmLFVd/dNqHub8MCfB6nb9OANeP
Kwp0GEXtv1Poq6BgZy8O9+2u8wwXEuAl5jJtotiRiPLRU6mXpTHhBfy85h8RjN/B
Zi5rKSb8dR0iwvXOp79s6UM/FwjhvVJsJcwAdr/F96xeYtwgOh6emweE0a+oao8N
ZRf5e0c15/FSq7apcyos0OHZLNhUC/k1pt68CijAdRxluIVphBsQ8ewRzx+tZTLO
+3eQcwDTQt6MnrpLF1a2f1P3KvFb8S7NnH0J/bn0gWJ0L1vRvcvYcK6/Eoia/k9u
Afx+u7QcB6fgYyTM23f+JpPCEU9DxBM1Wo1lVpavdmUy66uxMligtMh2DTE7vUzl
gQfuqRTczCH/srcHP/jfoEiKkwy2igTyNUZEg/lXFwM/O/U5ivl4yU8p4jch++6O
UQZq2fV034PTj8NaMuWTminyq/5VEVkXV5PRNQOEHBFdI4ANAmIJ9GgaQZiQMtTO
JEYV9dd7B9t5FZFHostaDqT85UgcNdNC9fNhe8UaOaG18llU1BArWACSKVTocyh7
m9Bn7dOrQEzWMRq5fRYft02NMKhuhNNcbw7nn1wIZQHoF+g+Z88s88aSh8fOq7wh
/gzWcnRXExxFomHpz3iQai8jgufPDlNq/PwOYdhKdUE8QFE64KJvJ7cK8DP/DC8d
CvOQYDFKiDTN2h5BC+4NJpmg9FS8oghReCELo2Y7TcSIa8I3Zx8DRu3gRHZqokzP
dGg6OBioInrRBNB09Kws9Fb7/NcoGmExMSjwo5JN0C3l1Q2g1y31pAjVfr1cmdhF
xAUbsKhTI0z7X0mgdQtkq0H4gpqeFeJqNPSonqrdtFYndzxdCRYNOVGFU/ZkoAqg
NYPgX/9ypkebvfgb+QpSK9bjHonVPMXgAME3M1kmgIQ+vwDuXYkO4d5fxQaAi2AQ
IMpG445pkK+39E5zoErem/4NI9k9sXNHXfIJBJP8eSsMYKeoNgjp/jhZnfheNuoH
ld+n2Q1K+oNtMUAAB4N/kjt2Ve9tIkGH8MefiAGcWvXpEGrilQCUDEWRh9GRCH0P
CJWiWsUlmUSBnEsQjcXhqpRRsHaycHPMwRRpNcH0GwAPRDJfV2zoFgp7tt5r+N+E
MsPCDAibMQhu9OPPa3YNixAEb2PWKebjgJTTAJHWMviJeCfLfolRu34rt8Kq9E3v
bjGt2aaKtBvt5G2z962CVoq0voj3ywsu5f2Ix7TGxvISbkvCHmdb6WaJrSVI5NpA
3mZ6WbP6Nn9gny7UpRtEHb3WmIMqnq18+2nKdOAdT9Ur++0+rsQAPqs3rVV70qdH
3sblwW1Zn0s/wPLHvDqsKFJ+kmPn1tmEuqmv17VMZF4kV1Ws/VjWpLIdzzmXu3bT
3bqO5JXl9okBY+a3Nfzi+W/mqeiZDMrmALmXcLCM+zkUF98RM4QLGmCMTkuM+CfB
RFDTMOQgmU79skuwrBQb0JQvhAgBdJRHGr1LNy338DissrHvReWY4eHeJDf+H8ur
UGcMOZpMDLuFnypD3EVMl+bJdiWgrYo9EdtgTaPUraSeiQQjtDBq/I8NMYjACxMk
sjEeZvESvMrHtP12nQskUZrwFWPmQKt2lvJRNOWtWBJTf8Ubh/AbTmkcy7FazCAn
sPT09QToMVRYlYfcZ4lYdGR0RN3kmhfZlPA4W5XGQEgK3aeXZgQgTecoJvgMcJtN
CCc/W2zwk5oBwEXV1hJUoCgDg5n7+KMB1Ve1oh5QWW6UPXrFpF8opK7ms/yuDH+Q
vfC6iXDI6mCUD5kNSVsQl/q6QGvLRfafOnYIDN897Q84ZeoWrsMCi1BuHCT3wBG2
xUSRt8EZjok/SBcnq2x/2a2pry65FMf7ASLr3vSl7ogahBz3SDPHFSoQQLj3/7Bp
d5Msw+pzs1cTJG63L+ofBqRs2xR8HUZPD5W8o7mE2Q9K+kZKlDd1zxSIs1Gv+DMI
vQ+BBo1AD2M0kRHKEnO9KIUmQMsfBH52eD32K0TOBkiQaSsAly1imXK8oDcgz6U6
gJzMBVILW06nNi5UG6RHSIGBKtaxxQhKiQUG8TZNE7rdkvQCdmQA+anI4jgNcB7a
R2R/+kGoSPRbYsCy82bUkpyVsBv30yv9XbG7SrtukLylw00VOhKQMbj2xLQ7w0Ae
T5B1cIyMnDAMcjMBJUs7xv81w8jBRPWsPNaoTox+pek9er7XfCYA4/8vJoiTuP5T
BPDn6U6wjMekdHbXrjam8p/pTtKtRw4no7vCeiZUGNPTAM5oUuGf8o0AtEVmWVTB
ccTqRxW15uYE0GSUdkHrt/qnudoXJRl1tQll012GpXJxj0lPZ3h7ddm53xEBRgFh
q33evlu52QStp6dDnal1l6M69vdMKJQ4TdqbAXdJQ0/MnfmzZLSGqk16lTUxA6ec
NU/EIeP9CohzYnzMz42U7edfjpJW3FLRXr/94086Mqf5BIPermB8P3T+H4cF8p3N
ePk6hGY8fbu6XgENjThCQSeqpWj8fQoOtV4+gj6hV2sg9dsPcf06XjG4Cy7q68+J
VwhoutKR8iHh9qTgyS+hkHukloRochNBLGUWqUDrmAY2vdt0s8G1BNSEsiO+nUX6
5381dLfqU5h4wK9+xqV/JY1qgv/db7Ii+WePRFKxBSRI8d52m78fNMx81cubQia/
B+eAkXDfmKKYpw1kAPdwqPnjj9fZxaGO8bkTx2q+efPUiGHE3XGJwdUwNzepDkSg
0n7GKRMDH+k7UXnVR1mfXqzHN/IE8aNn6sx03Uz1VZTSCJ4LTMDqcwPK7CaHZSnC
3X3k+Xhoru9bM/baFp0t1+6iwf9QVqKMTJpz9VCSKjKapAe8LLK5rumCbmWCZ9Sf
jCq617KXWDVr1t1kwmX1ryujVy57Co1o2YXV7GB0Dcu8V/9iA0BgGfavYkayZm7F
aZZBXBWkAOP/kD2SDn/wW4WxYvpoQewase/kJnVZOYAPAMBT+qjCo/cARmHN7Ev5
uhRYNsDtoZ20HSLawLnmLaLnOEuFIbc8F8KlGpfuMIzWg3T6ckNyo2LVy6XdZueY
6zcla9Y6Pt4I9tpZIq3WlgAqv3KftCnkVdkBAlBWexdeHYstOhrJrtJCDGyCnZZ5
7CPKRNt5eMctlHcS/p5XKq5FtKDGPKvNKjMyt+kcPvc7TLMN5ZxysjMp1sMpWbr1
fqMdsM2+BmJKJ0ximkIcadDQ2ypjG5ACphxo6n9YOoFDFiFUvIuE2ncS05+ioyaM
VZlE/6s+JXq3/qWDdx3Zkxe14s1AVaHsSvG4MpmZ+zBSKR13o8qv1jBIrBV2sBsV
Bw3ijpAbaXfBI8A8GhQm/1Jh/uM4D3e4Oaw8qPHuei0CMKO7VOLsZq1yYUXsuhot
r6HTHmrbEMlihv3Rd03VAG4BwGjtPhlqa/S5QBRexHUpqrkDOVtK5jEUSpMzOm44
mSXBUFKVERtROiw33VIH+WElQfIF6xQgTzw1pSRomkar3OZcIZBg7ZgVnhTsCTUf
na3gb3u4dJ9XULb/Barvf+yJE54RKSh/YB2LvBlPhtN4Ai2jVxok4ngjLeqCdNlu
nbF2psFpFtBViaKBJgInDeri/KyxxyTs9cyo00Y00aTfirdQHRIpdrlgraH24EUP
xLDhA0j8IuwfQz898fOi0sg+FV4IjMRALHAibbf3M+hxeGKhMwVjZK4xgLmTsNyf
ZrkNgKlfz8x9Nvf2lfaDwaT1xOnFX9uUU8GFRXvwGKQy/n0PIEIN7lANfawxJNus
wineFoMrXLE5VXekR6Xmlusq1TYlF0/VnkxijFi9P1HLsQIPFzygTWOUlmIabwRr
hvkQpm5VkgAQtcP2ZhEBCPqjB8kXEMWHDbHr7U4IfcsTELsgV8dATcx4BadBYrvl
XmFrtW6hRTGt8d031MEf1U/ZRpVCClnHQ/HpMixlopbrapD9pRRw28/hg2jqmTLK
yc4UYybhmtiRpPmjIoEGenv5ZWC7i5voHnYw0EsJVQaf40T4g6HXpWSNucaBm2Zb
9ciA2HjLJx0iAiqRAtQs283EBfKZJfHGT4uHiURfe68x4gXtkeBl98zSPS82fmUA
wNZIkCIf+jHyIU5KPvPJ+hVRynSp8XURERSrEvoz+AGJRROhfpa+BTsh0kmsasMH
uRQiHDRoVPvNCJA0RqbNFit1p9F8u7HVSYby2LPdnXDIzyI+fxRBw0XUkelCvnnW
IP0ALXBByEGDWKXETnnWEPGEMOv95GCneCxyk7oecN2X7s/boxmG6KvEZ7qhBLjV
/G/hXIiSkk31yoQIN78DIKX9l8Mw+lJ82dld9RbOmef1S0eNGQXkG/Vx4cLR/yso
kKBkIAYoU2oOON8uVqlvDCNft9eHghhHEwdzbe47rYJ/8/SCDoUORM57kaPWjIlf
HSxz7QmLajJUqyg4iECmmqDx+FbfR3HrmPdIuCWb377vTa7OWExmAcSW8hhIRB65
dvaAQ1WeixNQEcoN7A1uA+ehIQ/mDZe9vyHpEiRvzRWaStZvynh9L5u0rQm3FPnq
2OaJxUDls2btexoxsZYErXIJiF5Zb7Xh+Ydk5gahSNng6UkB5sO/fdiSnel+It1E
PHuzTNJQh/SlYvEb0I2oBXMjp6oTZeUO0skoRkJ9gUsF8cOxtDayyWM2rMjiHU2g
UdQpA2YiyEK0wSH2tQ9XV+mqdvfzdFm5qSC//7dEnQbB21roFf8Wvb6xI93E8asQ
StN+1Q5WDJenU3WgtoE2K6gYbHvP3pXibQeqdAdi8q7cMRFFhY0dBEBnYyNokS24
pTW5cyRkbnyD5lxLRhn0SSkQfDxO5AdKfRBRif+9qjj0CUOG07xMgsbtlFhBJKyM
X88l4uahirXYdbHejsXEVagyA3UrTI1qhS9PHukTt2HQP/Q4PTKcJu06RPzHAvxk
sJy8JTwIr3n0MGtvx7I2V6bsnqeeFmcqFZ5f2zfwQMFTUCed1qSEwUWjfnLI+YnO
yIxF0Ev5LM2IBqu3H1SFWki5p0mTmBRxEUIhVJa0haAMeqZ6qGjc+gYCyyHrFyp5
oLv4gaQh5INQNSBp2XZIBWy3STThiHyw+T46li+44/5m7QJ4JwDOMWi79z0oyzMl
In1MXBHWvKgtRN9cX29+X/lbQAAYHJNWs8TraiML/+onmucFVgHUexIzGJ3T9jCk
mx1ec1Jg+mNkYuhfDTCt20lF/DxHpSHs7nD5tcNoUhGyPRExgZoUNm9fEI+7g2tJ
9DAVEE5D7PuToJYRr2BF7GLJWJYd22OcKoomMK4l/ivVbNwmMLhAjSC7beGQ1EbE
KeNO3Khp6H0OvTFBgvhvU9O+v08d7B6Jmi/qJxebLWepdXjQkoaeJ4pZ78U6xnkG
3BaqLfnGQBc4Siu5uSzR+uPQZImHOoypKtmCbri4G1Skaxlwi81tcNJW6ZeNXHBx
oTniwlaKn8LP3bSJkbJ9YNfZqJ3YkOb/DCIqN0RAjQWsoEzqRdCLrshTGfl8x/oy
qE1e15QwtUTFQpYusOzntDiyPSaXFtZ1uhNzONtCV0LImH7PgLbuYJf0t3e1oGaE
mTwF3evfL/ZAx+pAbVSjcXAnoXsmAfRCd6j5a44RglRLCz3TAPOtyUb5hlPMrTO9
RDeo0jlTTIrRwpKvqJgMjMN9DQVBIXRPwn4bhBIEcLnpOQeKCslaYdUVFqdyD79O
6CRStIJHByFHHbmKTZ5lv+CrKipD5aKtyCAxTnjQcaIpgQcv/yt1JcUOUAiZLSYv
SujLr3RWUiGULHIwBHTm4z0TKU6/K87jo8Qp7+hexDvjxwAD35mN/L7YjQYtSH9t
5aH3Mq94dc8+lxLPmenDz4aSaxy+7tU4ZaPL7HhkqGj0gNqSxmHazWPqHGHpq578
El00D7yK36k/jCYenMABDJ29oVJ8I/mzOxH5fPTd0iUEsYcOiErjHb6wtofk+Nx2
Tp4Y4eoGkzTJK8UePYjmdUDkGI3mTCMnLjXaCrKMdi7lkll4UuPCxyDyaGiRsHQu
E/DuoPTe2ocaI8uLcfSd2ZEvmdPJgcJKQaiH0IZ1ivk3RYVmWEOzax8vF6T4Wfl+
m038uMew6EM2UgGjK/cGcnjJ4Hh23sRkTHqJPejghl8vTFWxcKRanx++DGgZVZDH
DhRFGeGqhF6QWGpWhYk9TvXEqcpYlR/7NH3RNye6ZBeeCgEGYwguiQjSWPijbBYZ
lLTBGvo3SAPT/GyP6b0KzntMF5xYG/Nl/0KqVtxexTm9lEuktOXhIUPBtwiLl8TY
bYCkPdTNpLWUtucddCFPw2bsinOTgW+zMUkLOpdc4Ddzgfzntex5qje7g//LaiJo
20NZ6ESN6but9OcViwwjDV3syQj0XIFmisoIQFUw0QcfTIb8iXTxKGUbMQeIWq6/
DK/Agt1uEWcD7iKK8x1XlV8UnHNV95iGksoQKIXPfIj5l1ISC1bJzIBAmUGch9/W
BeBCSOdnRw27YDG+boq+PTZOeNMIeZy6bCzIlarqp1byEkmL0DMSPiRxW2x3Or1Y
9rVUOs/5+sLTnOGlL4UVl+W21G7+yhbHviHfXbdd6AB7o9iWtJWZdgmrvEEZO402
mJehLMCAzg2lqIgnpQqCz0y/sLtQXFR9KBTxeEwcV227PTyEwLTnTu/vqKMWRNHq
3CkaJzGgQCejEv4UgOewERj879gZ3Pw0tPtDRlKyoljgsf7peYA1lANc84YoG/ap
ey8uorCOdcrkreWLN0+ZcdXroNB0CITxOcvRIf9P/eLK7lv5+aQRr44Cf7vWFE19
j+c8DlSnNwV8v2Ua5VMZdOo5YQU3vpjlwM+xQxKL4NhtejKqAa1F/uPBEjiY4quZ
20SoPHh8OuBWAf/6oWHsJfwEa45UctVAugfj/AKrfj8FbjrCxdjmBeHgoG+p7EI9
PQ1wbdFBD7Olac5DY0BA2bvSpX8kSHXqvdFo2jf+7M/aE02w4MnTnjNYscm3iHeL
WUbdTo24lFYsdN6L5oHlmCYcB1YJIyDsCc7Ku+5eXjmOkSd4dHEHGkfzlIdX6YYx
fyVVPn/H9L7yvAB7a5/eNkJSaLxGyG+v8qeUjYfz+THNS7tSYNCl/3cdH1Zc0tSG
BS++KWB1dhHkvgpIUaiK+g3dpGRHb+vCZTg1g9Es5iBqKaD8HEhRJU4ZWjQhDYr1
kkTQEKKJK7OBMjAWirn96rLor8J387MgWV0DKelYgpbzkj2FTbdMUqW6VTn431VI
pBnL1p5c7H5qONSlIxqmUUd2CRSsHf7Tr1tGn77uwKnnmzmTXx7SB3WOByOz33Nb
SAXIouvtrqtwIIgT+HoNe5JW7vSXHDRau62Xo2x288atQB/W2z5KG76kc9CYExx+
2uwQkPYlyPE1ajseTYDyEGLzgJk9Mye3GzGvPzTbEoJY5LYPG1AsCUlihl7w3JrA
et82WOp00xBJr6tkHowHycXqei0ACQu7HBLZ3fCVzGKxY/q0Qmno/l13VYG+eNNb
0LOTTEgP+OycneEKxt4djaDK74D8xi4z7y1YRMax8wl8yyAI08fz9mKQffbdYm2G
VHcvZJFO+BWOs4X5cCRJ2fsBvOrq/xvh5iFhMZw4heTgNnXclddzeCKtn27o4q2m
+WP0fT0oX/2a4l/IjdKLrtrQt8X9IN0eM6C9NxTJtqxH7lb58N6hA1VpL/iouAZ7
qUXcqbP/uWAW1Rya2z8mnEO494VjM1qBR/l+rZ1iYRKuXn/7GhS6ptWBEMe5GvCc
6Zo46XBsA5rlbjsY7w4Gp0kyJV+4t2kSlX7KnU7dNvn4p6Au9qzhl6W3LwmmrCWN
TxpERaj5Z6RejnHJp2zZwrBYOMeLUEpGuN2v0+pfX+SisYJVWLotGbfiYHXj5Of8
Z2btx7QP6E1chrYRgUBVKXc6ceHLRYfzoexXe63CGpaVp8v5v2mnkUGFD8ZLyt1f
2rLEe3zF9ED9rENsycOKZtyNVJDzHgKC3PrlCMyKDsOy8TKsN7doIN1s2fAeMJAT
4GRTYHHqsGMhmwB/0gNPB97SrDJjNWthkTAdvoMp1+HwsYEZ32iyY9xlmX703pWM
F45D7ohIFksHW/mSOCy2wqmOZV4nJ5BqOXiVMN3t9H/jG/cnEOvnzFqZlxwNRfhP
Me7JI3HqBo8ceNtzQFqFTvxpBoaelKoPRA3bp85xNJ/SI0CX3UYizgwMexEJ6uwK
Ga+vPphLxbSV6SR+3kt947VD4GwnsRy3ShkeLf2aQ8cRmFv2dvJZy8hWTzgBtgx0
zznfLZs/hFZt09PdNVhEyS3sD5WzExbnWA08lwUuvQXxZ1HeHNRVlvD/LNiHmFBh
JldWJQsyRcgVbpMdTogMakHYzWI9Q1D5WC3aMCuYOcNSOYlIStoTP0SXt3bw8SR+
DVBlq+Fko5C7RNUuCMEvgKSKAPYv7cZuBJcjqtgO/SUcMiP9NFL/QUHzyLyiccWe
Ix8Va5UOtdY3b30xb5hOSK06kQIZVSi3a5msvdo0aaSmLfWOAJTtSzm7FvrMA3oc
fuvaf5A/z0yVYXxBL2QZoVBLPUPoUu2wJG9mh/68N1CDvyhn1OWQqmPcMtRVcJAX
ODG+zTdIbbdjZ8oxN+TTKyE9u+yZHIgjNbfZcfew34byGz1J52QguPkSGJpUbtJJ
rf+RT1zhxDJB1kDyuxlmDc1uIbqpV3XKw7Rwi6Rgh35ZaiTVhciN6VImOo7nNYyt
WjH8sRbmCO1PhX5QDsJBFNRVyrAOSSnhD+wHMF7LCDgKvCB9yvg7lWKd2mFQvldq
iZhqhytRznSSh+6EdoPZq4VORQoT4y0C097ouHImp4BXRDlwQ3wfV8U3qQjXsXpd
ifQui9bLdSe7D+UqQ1gMxrf/rKvuOAK61vTLXyDRTWoB77ARJePHR264MTfdEyM8
pYV2aUtNCtnz5Y/7oESWwCTsZItaGmr4LIa+OSlibdQYQdM6lLFSYa8a8AeQ3RyL
UtDyOeEKkzC6XWhDVMOmj6xaa7v4tS+cHvA/TySOTquQpi2Cmwl1Ccsvpo71jyGi
M4OLLenp+bHeI7oNFn6RJ/oDblyo/R1qns57Ho9Gi6+truiC0njrbbQML3pmbcCJ
wzQgpq9XqJ9WfzQ3uaZfSVPdtzpRPOb9SjPekJsZ6m/mcWS2Ip7Cc/SSSPfp2Hla
wlRIpg3maCJkdlLITtvDseqFzi2K0i54YPUJFYA3T//sGKYWoFcgdCI2Xph5Kj9o
qc2EtvAUSwaKWs3JWauDTr0zq+wIyUKAdpImz06bTeNN83yEGm38ohcmyy/vTrWz
uFSloVW3SgtjUd64Qq0fC+b/eSQsGggO+n4/44vRUyx5Rm5aTsaCISxexoSyCBq+
DXVQk0m/e4lKxhD6dMQE5OnEqksUYcOecqSm5K+690ZARTaRfLxGe46drFuQx3bD
uwc6kKUztMehFxHlBvaVLhKKUH6AMLifNUj6Ea2T4BFdIZI5g39X66w2WE4qCpQY
ixq8AhSX4sUDtWIOkhThtZg2t6wMO60tKa6R711hY4GJ5u7HCdX14G17QN7+kVG5
NJ7grQlnk3M4bPaKtKcE16QZFnGGf73mg0hGbuGOPvimt2qU5oxPdn3hnHfgqFAi
aId72Lhw2jjFnVQ231bjiwMyPHe+EiaB2CBqO8CK3Gskma2cm5AtY4cXgL7Dr/ta
DxU1T6ro/Jn3wanro2VS5DHuKKLQQu/Yo+QZ4zUScuW67pGofe0ICtCMPTNHOvI3
Qt/OdnL/9O5YS3cuaqZ4fn+XSfRNBJPkH+PY//1GyxkGL12fgkJ/WrBDSz/2vklM
hzUFvzPNz4SqOKQSfWl/FSkDIh+2LlWQakzbU4olY4OaTv+yt0yHNTJw1bMyv53Q
oK4Sev0NMrwiEDPZ2fsQmlyroFal9F7CG40qQsUslL8D6amCBvadnrflFFAMx59U
P6hPA4LOUqwM6mlDj8UauBHhU1cjqjWV5rvOdsLyqYGExW+oU0bb0R9X1jgthOL7
BS4J6SNaSXKMbwFIWTX7xilY7WbzBlfEzop7HBNx9YGFDoIx3Pvgu2MupEip1/nh
XXVFGwV8n61E4gxanfHE+vFI9yasv/74MA3Ey8leVs+bd7Tf36uNvY9ScIcH0V2C
wFkkGCS2ddCH9chPPc/xtA78lWnZw+gmQ8aC/hoqbTxGzRg1K7nk4aZfC2CCT6D1
nnSnEOESpERxgOFQ4duQbKqJh2cIb56Z7tq4uNmXCYNK4PeuWUQMyw0cV//Pw78b
ltgqTBNWm9zpoZbWlE68IUxlxuRouhbw6eApvusoUKkiFSB2Wjlj7ev2wAa6Gj3T
6JrWVyA+2lWtOdXxoMOr/hXGgIGDhaM+5/DoxKH1EJv63dj7ydNjO5/B++meGVd5
CSaOWXY9bCN8a/qq+dMnuZCnU7eGWaUSRLCwBjaMmWHboxAWj1Xt+WXebu8R/q2h
XYLfkIBRuZ/fO1A0h8pwjlP9Sgq8vdEu2irancHIAdcilawZ4HE/GuYCOQd8+02x
QcILty11NYutvtjWoGMMnJU2HrdKIXs4APpwf5SdgHbwXweZ8jJyxbaKTBmfXIje
E1tzWQ2GwaJfz2UWo5FKKodA86CLH+2fR9XYj8hiWDFdN/8dOwrfGRGTx27hqVUV
4M3WUEdr7LG2327oBOzIWF4+iieVgSrH4CIBG1+H22yEuxH5Xmz3a2yuOFGJcKQA
fNrihOXHgAiS2t90Qmz3vPDuWVvMxuigqD/s26yZ0ym8VvcJdOj4fpPGVil3T7pd
OgjDKvPhSoV5sIOHAsMfKXVMwkXNpP+ZoT/STnNIrSXr1bGAivk1d96C9aYNKdvD
EnsIfgwGGykXh01T0tqnPwowwzz/SbeVoRS8nFPDSTfjgGJ42Fh/2fOfQwOUXGUV
R6nBzAk5m7q0uwxP6F+KztAY6+s3PrTT8HK4hLQJiHU05UAiPXQpUHSLH2agGBfV
m7V0EF+4f9Xovjf1uS76V8eLbbUG2oih+huCcUZ4vGMyetnL+uG3SZcew4N+s0ZD
SWCTbaY3OmjM1hG2osy61hYXq8am4qPvkMOBtAOkKtgUGE4yYmFcbIzxZDDzjNEv
ywj5mda6wHgxRJ6Yi1zt134GohPs9JjEMw2W44s4rylgxhVKF4HvW+/pggCf061n
KFkCbcrmlSg65AUbMv9kWo988IsapXlAuvuN/qEB7ZFv0WW+3apsqx7hMg4bZuzi
xrS7Px7yCoKap2LV5B5cprCfahmHCUXn9zbBAKrG1nDdABxFWApeOJwFgIFOQgXt
HqnY/wqadBcYLYZnuXArTWsheWJMhohwU5P6vtJgic6va5/LX3MdkUBGCAYm+h3v
U0WyK8gQ9H+JX3O50tbrK1wEmVPELuwfedRM7PBEt1/GlfmD6EGfVyebuCj3hFh8
JkD5Fa5GIX9b0hmwttIUXdsAibdLtS99l7QJZObN3rr90wvdXUxc6opj3fWwVmuS
SmuVrLl+DCT5keapQVxaoBMLpF3zQ9rUZfRQ/hUcJvxyn8cOflZL78s6NB3TU+rV
3YdGWIgghN6jCPnSOCMOb+62mQpK++vGceXz8noACznWDIhse3V/KsogeIWQsizF
I/oyu838SUmmTCcPrFLWy9eNEcQOeelGt2DKQL8g7En5wJQLr8M49FDyHY0z3PZq
BHxrhDqlY9/uCC/p0H7zRf5pqsvam8ft8W96SybLjtC5uqw51/JeUMRWazCgMlTw
IAOkVY1YvsHbyPKTINOCSN3wAcL3Ijp/hi6QXZp0kxUwNToVtzO5c42tDEd3Jpo0
CpkXc0WnNauMgBI4b/Rlk7w2NIstMOJ5PiT8ROsBK30Q6rhnYiQdPBeFBL5WOnGU
n3iI0U3FdG0z3IwmKPnVJ94dqYRXmJ3fce7GOB6d81GO4v39pVRqw43fHV48QVI5
7OlCaELYSOZ3cFSIKdw/MsoWd7334fyxp6z178AqHgr8fAG5K9ef8EfOdDYCudA0
JcCeHtatcO1j4Fu7tJikgoIcspa7lAL+3IbMRpv0EdXjbCei156JBPG+FnUM02Xv
uA/l7lKX+EM4s79/Fp/ktmYrfpgarLG0OlIuYJeosBkDVGKCspNYADs+qnTDtb/o
mnQqqMzSctxva/1zq3CcH3MIUk1anmiYNDWyKC2CzBI4nytm4oUZNDSCko2RCb+9
/Qu+qnBxR5Go6kkIfJWCxuVdY19SjjaybUl9LU+HJlJBgu/UBb1nwO+15MQ1DN/o
37obNLRQ74yWQjwE8SHoGYbJZGTV8wIQdZWf4VIcaWtFK7gSEtL12rJHNyETmlM4
xG7kKxM5aISQoqwpc39/O9iSARCTXYrb6oNPUHFoM1vj/5MnVM+FLBF8c5WVENoZ
H2XoGDCQpTPDa3jDvmpabN0zmSYmnifd2Oa5DKS8aa6Uyy2KfGR34XhB/oDCBj7/
VkN+Ni6IFZfqutV9SpLmfyB870yk1oMVg+f+HbA08F7FsaamCKzdeHPiuU8Btq2B
e397btMVt1686pY1zPOEbINASZNmebqKPCjVLL7QyD6/OHts7jrbjpPhA7VGa7Z9
7bpY3j5y1wXfIv2jGIXTsbM8aPKHBv8PINP+3mK/bvPsqSj5aAZve5i+PKdvTu/d
AEwNVgsjDbDf7D4va86OFoiLkb6gPu/sKR/EZ8lNi5aXCeEsOF64VTN1kO9MMG0k
iUmaFRp2tiz1ZbcHJTdXxqiVqr4yid5V3HtzwikpZ3I68cxo6JiNX9ljqzYK3YQN
Nz8ThPGYSghgHAmPagR3O7HoexXCZjgDMz7nf5uHKssWq+gurBn4AWwrbnvRD7UG
0m6idpqGFNBYpk7kh9Jzi/WZoLebA9HTJy4crid0eQd5Ui5MWaBpmpwQMQdtIzoj
GjAdGmRQCIVIIb+F9TCdA7MSv/BmzuCJgNJUWl6Df9Eco4uJsZ58hpZAqkTmvvHB
scJ9zguD7XtbXgUEF1snybkPFA7dJ7Pq4kAaEh3TtDltirDUwDOBbEO4kQbGierP
TXYAzPyA+4f4irmPYMJx2sSxU6Ig62gYfBvHXo0GscEpRbswtgDoBbvKhLDZKt7m
00SxCEEFKA2+EFh81XLuyqjO42xHqY7JgoIcY/F17yABtM//ql1SSIe6oxvrHhi2
U+htc3bAlUUP9lF3laV5eHY4VLr1xyseW0Z6JBfZXmGaDbhvJCGiG+6Ks0ERxagA
Cvn70mv9RdFVt7w8WzqoJ+XWDCiGb8Vrfx71PlfDr+uvvwsqM8HFMpauv+gL9nmR
B8KJ/3MV8bjPgdkb6M1MpUxbQwvXW/2p1aZzbOVI3JVhVlMLr7DLuHSSFUmW1eZX
btiM9t2GYLWtlUcHffod8xOBcpbSHrrL2HA5zEIy2Xy8JoO6XEYOywQ9F4jhMq5J
AN2KGBho8kR8bdkfri7VRwS+In/33QrALAiNBKgTYrqRDBsokEqwrgM2mqsr3HFh
VGhT4aRXP5iTAprZ2wIAQ4CFLIQSJdMphu/XI+EoP8TgJLSSQBp/q8sbl7y54+Eg
kOUgo76EBn62eNq2Jc+7JH5oYExVK2iq7jWgTS7Bn/6vvYr4wUyPsLyDVVE4S4sL
eO7wvXaiC544fMMJV2Sgswf29z9ZASOLhNOC6LgdWaCDEWcblbfoOtJ0mXnVsYCu
8zhi7BBw7KQAhxLG+gxfEvYYNwoczyg0j+sGI5aXcNmexviZSfs/WXJO1ram6q/g
xvKNZ1OVRNkeR6CeygZMY6qN/SYlEBGE7IGrVQdLqs5iGWM7g9h3iQLgTj/1c3l9
p5n3zsmdMprGbnPPsuAj7j2cpRZGILKjpC+9mZTQ81oS190/UDgcHgO6J/nYUV1t
IA+6+5wPQJNI982FaQocWDbcfza/3a1Fr5Nt4b4eeI4IaNXSFn9rufKaEjmHkIgj
D3or+pWd6qyZ4bfLbgdV7Q3V46nV6AqghxftvzeKMLNwjbee4wcLC/qVId6RNlHG
94j+NDbE0Mvt3248VPeNX5CAGsawr2yk7t3mxtvAwA/iz/7IL54320SszcdXhssS
OQeIIJkTPIN3b/KA2TA1OmbEm+kcp/EDWNYy+JK326qEzEqvirjMypeOd36aUmeD
FRU7AUPCIdicN/StT/OJzDuxJ03I9IZ+rTV8tiknwBhs2U970DqRIJrcCpULAoUB
isOgTFkmIujvRpVuyiKe/vtpwj+S6x9bVFx7H5l9zh0FBsqkOq7yPnRbWSezTI48
Lqkow7y3dcLWjch0yafWb1aQRFu5vHEA8WD5YaBP75uzhI4HsfV7oO5jATzSStO/
ZU1pzNJKeZPrgI4Quzl7/DJWSbXXBv66r4N0ncOvNOVn/eFzTX3GjGTVsvbywuNe
dRSiLNJVtEyUCHlCEHUHTXzI1s1ZsSdgkFYKvjTRGwb3dbI+MxzWFNK1rr/vgHJh
g9wROaSOdfVt5K1YuYlyglsYYqyOY2cdowX2ZOmWt7FJIWVMsNvOsKdVFdtk1+ou
331Gtxtg5ZG9Jt0Rv9N3PvPI/BNVDngnVvdvs+gzgkDwmI6lGWNmMYJavS/Q5SZL
0SjCdcjRgc8Roy2vcTneWF/S83sP5Ats8dGyxZufyvuq0A3jq+z4gxZeDDcd9jXT
LQmZ8baAVXB4wURGjwE9KZkq/vNfL1VfjZ3VyR0E9VhGE/iPjrtnjl16H5Z7NDVF
MGyA6Xvip5H2FOtz6OqH7I6vSF9RiYKlNTMRI/9KVMh5UoweECb8mLW9lGfUVK+9
Ya5mYDSWHGDN8J2w0moyWhBszpJWVtmvpJcsv+R7rvG9Pn+WQGoe+QUEWN3kUNcR
mcJna3Xrc8uyh1M543JMYlA9ezaXOcnuOlxOnkIm78iZhuwQuBZorLSYsL/18NNg
JIPoudClBR3ZD+ckCG2OVDNwKwTMwVfsdSQ/olmg2th59S7RsTs9mOFGrxTb2Z5T
D1MufFYlcTKYo+giw6J0NmtpzzOTmfn1cXxwRFaQTSukyvA4UAttKJ6ewFqJHHKl
CLGn8z/ewC+4+jCiK1NqvvZ9wDOxyrcZVlwLU80FxUzyfa1L/f/MOkl24Hg5FcZM
Iqo/1SPv4rdgJl1LXp3M3eAE5e95YAGSRGnyC6cGpmvwRBQvfxWrFGf7dOfoJ5yQ
915jhBgt+crBPuQHz6BFJJdBPwtZWazT9t7u7PmbnPDfKMB3LzsbBppGbFWlPN+F
x+jzQVsodM9FPq+n3sBqMrdrhLND2wmuqO3jnPvy9m+1Ei2Or/4lNJbGlURBH+Pk
zhpUMENm1feMp47MPNB49+vrKHiueC45DYnxzcFuEkkeGeLBMLX3dtqW4gqSbP01
9gxl34KOEDsunshm10W7+/vYmSxu0I+YGRA93rMnrWhIocMCjyd/z4NuG4pXnVOp
00FSRurG35yg/RSB41SIogDB8NyTaM+qPSJci+Um56y3B9wMXW0YvAxJ8cJlHkfC
YovvKmBOsko2oQLM0J/Ymf3HcSiNzIE5i0ej2zawGsOxGgaHETcNVvpDtOqsWCLT
d72TFGbPbdDYCRUWUXPWTj5y1MsQI3fISjEvEpB1zuGEpKP08KurRrdEp8Fp4q/m
mPudRUXESEzkUMOrk2RQZY7LPOG1MOk4+A3RZzRA2EK3CcnqafTO2a/YM4pvfBPy
SPLv2BPhvVH0ZswMlsJ6tfRVj/z8UFdQ1bv3YFcv+7EdUSW5QxqGtOSnPwCMN4Wi
cEvFnzeVt3gyI+hvVhGaQ85IrY5F5Bw9rEfLLtCZYvOTIt/YZQBV9H5vOEbV03ns
HLb4Ijl/mJSKE7CdcedmiYsJ3byPwKGob6Qx6x/XvW9NpNeeCRcAL/A62Li5dDKt
DfxQ7QY66yB5ADqMg8oz5x0lT+gDQHY49OX3L8B384Rb95LY7bpj1k+QC61JW8mY
J/tYqh8cjjMPdIQcVGKXRcN8v86C+hsZgJcd5FChiuZ3Rkd/VWCxN9fZQPw8jVIn
2s70/ICBgaBcHF327iCVtB9vQnqmwvGywEse6IVR6ICSfzUH85MVdT61I0lUHe4x
ZS2O5zFBfHJnMFIJCBwFDxO2+owWDdEQ08uakHJHk6IysXDjRq04vbkRudeB6FGI
bm9ANVkyG1rYLnyAJtwMGt4Jvph61vYUCIdoRSO+k4exqHPUxb5pix49BRtM3JaX
XALfh5GpgHnU6VfUAipxKLi686+kx0LB6HfRG5rB1/L/L/mYpkt1WliKqhxXu9lH
tS4tbsDnRA1ma+uJa5i1qA+9MgeHkdu+9xmWcpI/fGQu4ORQcD6ZjHfsll968vf/
jvL6HDbFGn7WrL1rXLqyUtt3e0oL4JDY62heUZiAjMnepbNCzU68+VCBaUthvxMy
Q/fDtxyGV6voXzAMmpwS6apDA9yP0KrpmwACLO7EvYKd8O2nJHFVDurunkUz0NF/
aL/ACFN9McYyylSXgs0smJRgwp3ukVgLUklcFHtHVwwUuNAlprKZa5Y5xQM3hVOE
6zpAPczmtkXC0jBkcBoS3vU1siyD6w3Ux2PaCDEJV4SeS9+CXp/uvPX/xpTZC51H
woz7NKoYaqrmNfjC13vm0QmvUZz3Cf25BlepaqED0/hgnaStvUnI60RwRR/Q+FAQ
e4IINjirm2l9s718tpTW0RpSsvzhizj2L9oY8i9cnEa30tavf0UK+8hfwiwwh2lx
+9EJMJANg17MXdd8+xWcyQqBsl3gvcXaBpO72K7JJtexZVPw6zCIzZrWP3/MN+ER
TbxuzqHVnwCYn7wnvfr5yVPi8rTIltybWxbdHXlnxJbhmnQhhKTCll+u8SofExuJ
ubJ+mNNMLZavEHAh+KgLvVlLPh2UqofaFqM8lQ5AuQauxY2E5C5zHRrGKrxxW9Sq
IuldMmv6l4jHcAxid6kwJ6f+g4j+kLjF2yW6ipBBFPk5HJc/d9JKVwi1kuLMTv0M
PRG7m82g7nJCt6Mz1mXK9vlASdII5TrxWcuLtID29CQ7/ZNNa0km68N+iFaHCzK7
eZyTTg7HQK9TvD8w9v406gtXJcgqX2tcgzhPccj2/xs/zzaEg9UzQKVa0fcZz6Tj
rjcvydLrz76poGQeVwEacXeqfVP3zgyKPxvhpoNVGe4l0hyfNDgpMUOkdxjs0esy
NGlCdhWF3BtuIu3/izbrl+DIP4dyt0eq3dxQTWY8srNKDXuzS0iiHFoKAz5Hcova
WhVbjwk7WX3KGaEDFd1oyqyyv8EOl0SV21N7BCrW0lF6koFiZVsRrdUxLq5ZHJwq
sAwGWa/SnT1dnTnWAErgDyjSXekE3NadhQOOxUhJE7x/cuzgIVkaCvd3Iu5PhP1f
2LN7OQALaB165Ny84SFXG8D3nrZX0nkLbIYRcX3RRP09GAKVlaRg+3iNHE86rQB0
QwrLa7Wfm5rdT6PjKajOa+4oCduxrhqZVo5bcQ6moXDdSvqqy+NtwUmyJRn3F/sm
Ydifm0vFDptaCtb4n0T/jkSaKwFQQRlqjABpC9ng5Z4azcgOD40tCoDiANTSwHac
Vd+cbzPECG86OV+NouRQvPipY8FmMZzirpXhQbJDW3cSkUfWaI/rIUAnZ8k7AJwI
PZoKmN/6mk+5llQ1+EWt222AMEiMvLhavkda1VcK9xxRaQYcIhNvoWVkEOy7SbRL
yDEZKQYvblbP/UV7TWdH5Hx5rRK+kzSh007XFwM65FnRsdrtRwv2fwnKIa6ONZ3M
4gNeouy5XZ/YNyIgpOtAnjHoymJaRuXR0/pwh4FYdNlFXo9KCuf42b3vpQusJbOf
komZLQnfLfEnUYojUxyS2rV0F0TcA/3OYAZmfATgpShvnfsRAItTmwJniQZwYsaF
RfeOhLNkV3da7a0F6rpL57lEgKnTIR69ctw7l+nCfqcUp1sV7lcIz8aSHgJ9ybIv
rrcWLwX1SeUOYBmfxiqp9OQgXPgls97heA20xBJwqfDb8Ewib7GSL5PuTyTIjR4l
j1vqyKbRV40Qf1f2yLJel475nZJyv5WWVdQD2SHgyTUoL1FJbW+gho1rpJNe30qD
Yv9wj5m871sLD/faePvon7t6NV1tJfbYPSBtMnLAHtluM8bQ/vmmIWIY+4orZShc
6gxY9ADQLhg5G6I1FBLiQxrs/R67ohgpQZgAt3hDKePj1t/tP8+Ant+Kzk2ZIwBP
NFfQN+8RedvjfYQddThcNJr0bs7eRrfwCJRmsQZ4sFcIqFvFLmSH/JuB5GRPHQt0
il/iXJPph6IaexQR35Hp1n+1t/bgXQ5LA3BI/XXsB8TwSnzXOxJoSsvEWBiUJ1Kb
3vXBvEHRnQx5Y+L8TTvHsQtsiXZ4pd8uPT4ZA9vmzURFx8ZUThJE6wmwZH9JGLke
CHQiMUYt2w+Eh5ckKAE3fSMTY2ud05x9Au2gym39qcPdR2r6JwYEm6N1q0gWxeeq
Uk8OI9LTlX8kxG9yo28aI+8PAgH5fKDeNouoBawlCM801AvD5dWg6Ays23b/sQmf
5jWuSUFd4RPYPAVol7mMilSuNKCHJvZC4uS49qdgo0GMNJTSKt4wEN69quej41KL
RTJBa5SzNxeDTffOoa+PjHE/URVPSWIWj/yALtYQ+TFW37Sau9bTLpuVylBuqSqF
yvh7MgMPA8fiNEVKoAauGcE9QAc8N3x0d9ifqKD9Rk+ud180rKxBaXE8jYihi6EZ
irjeQ4p3LC8fHhgThUzpypq2aGQSwC5i12VEUWs6nw7WZ30ZKw7Ha/U0pqGWlZMP
EwVoUE9rwe6e7dvGCWasfJccwifHw75/jElEOl2tLq4LHOFvN2Y7HNa9Ht+xWEGX
LKR9TeFZRUQoo7yrvh57cSRqv346aIniAB9cjXrdE3UEFlg4x4TcwN1ol59Cnou8
uXONLEbYJoxmkpw2tu0/YslDmuOg2RCbzBdoRnAJtLt9oejFQhmg2ov98n6PnAir
OwcYpD9ITnNlGg1dhUmOAIPn2wGiUtAA56XlhXIHA59z4byS8m2DnKHBQeb+d2v8
+yf1i+GxI80oRRtIhNo/2Xlra/0zFUblefqk4qXrPzCNchQGEHfrobj0HsfxmQNx
ddw+mdTS7AUQCY5vVT9ejtqiG7EIudeJI63eImFfRzj9HQJqvksYM2Hnub80MYQR
ATu/uCSL2PAbK3FlgEKb96O74hbaYU9KjAKX3NzIdBZiMvhSHvzaWSyNFbg5tWqJ
BelYnzZFOTRnyPj68eO/N0/XaAXvAZVHN/Fg7Cycw7215zyaFgxYEDwZ/9orwwBH
3fxQxHtD8DyXA/beuwt7BpddLsAdTPt4130hX7+Ac4QWU4EZyxS4CfEAVc8kDs8H
RfRLEF3pc97E3DXFnGbFK7RcxNh+VkiL8lgqdGL0EohGxvNOtReWuKwIRIHYsC4U
tegArBfbU3m00Qtz70dJEKQO8/tn7aV12UZ5Z8e1UWRmTUT+fOWwSF0m2aRpATZk
0qIiQQ6zixI4EbU9yblvfkEfbdliibzEyF3Nnq9GegAl44fHvuu93j9vZb7Im155
tEN6IO0nIrPLNnStoqsko9MCvWHqCp/PuhDzjv200+vQ6OLYciZAXzZjlWMOkCHk
wSXVIGlkhznak7SW6ts7e2sU6hfX09oaWiXCSki4IsGSExq1J82vbm0bmbhQK8nR
nJOvfjOtuS3HlvPdjqkkCCr57lShQ3zq0X9BdVR2DRA7F4Onog3/LSrD6OTLQsk/
hhaJcp3SsKyoNf1ZSmUGSkF/EOayAunTlVIZ01d5nnhqe0MAXsKJLyMObzuR5Uk/
oAm0Qj1vtOwa+WItyWcxDgTY7JhEJjLc5Fhyb3w93uAMaGOG2TL2PBeohSbrcUlj
3gbxoH0Tpb4YruDDl5yJEZ7bUJnFqOBnt2mya4ImL/k86fvC6Kxvg9EGDfSCZ0Kp
dzwyV9Q/dEWDolJdAER0eSs5XGalw2Qe1ytYuS2aPf9ZAlTOYnS5IYtzIusa60Fy
9lcSPPtN8Fq/cwIJm4rOFZM5rjkG8lxlWuctlYkvs5QU6W5vMy1jhDfFLIv6+CrL
mFyTmCOFubmBSzLzfZJ9pkovHlV+Tr/s2bhTAbx1WWOS4N5YPgoUsxtiyj+E7GaO
q5LBnDRAlbvWBFtqUN6XwuOojVFyF9KyEPyj08RqhtjucNv79IGvtrRWmtCBwI+F
0CBRgsoRmYsP898uoWD3lB67cVyfWvea9F9t2ZuGXT0m19ER7XQFX/xEYGwpZs4v
uV/9uYI8NvoDc6gLLmcePqgia2S7BV3Mo1/zoCcMNXutXU8x+5pke/SEPA0NVWdg
p+OERRhfARxRfn5XOdppnOm/QD70fLXyZ1+TNPXveIKY8owBDvYO+h8gUjEv/6j8
Bb0MWytwWUagWdRX8jDkv8O9JmBGxZmf+5lRD2tvI7suCa2UZ7JJ+HeNcHtJ/HTm
oyjbW4pY/UzMKP0QAT6//zycgySOoErlF9C3HBq+XXViPkfPMwhI5IY0M1LTQwof
8TNiyL6Bo933ujYfJ1IKQ9L7MFfkSQN96ljHmuYMi2E9ApHwYYPAJN2RgyKZWvok
+Xsk6/Mm1kxMucdxTRxEhGTnJZiWHw75RpU24k/0JB327rzmXT92DUf3F58it+UY
t6TYkyvArlK78CJdhu0c8tE8cHiLHPRFQP/lavMOon8TlAqFvWXDDRTdlKh0NVrz
Eabht9etYhwMXK6ZZBwrEh9bBdaWt8NYoSvpOYpTK5TVtcENdEkBw03JbONUCLa2
O7tEz5sG63bp+8a4pvhSGvF2eL7nCcqafFgL1QdCP6iE+F1wCWdk3p7iaD2fPQQy
7tSHH+PqISF6BYhdqgTkTwfZC7L+UQA+/T+xn6KjFIc5uscgNeDjFjbNFjeWdhWB
2Q7RW+9HMtzuGcwfkWD8TRjycFhpFbxU60B+EvHrRfXsZk1v3hi11ky9hVYy3r3c
ptNJBP0dmIXZ3harCRDrphaQdeeWMpRYVfDVwgtR9n7S7H8V5wO5NhbyhbSRsF9C
PLOgmzsTb3iUBOvCPIpI3u4s+X7Xzh5BISKc8wFHicNFr2olQkNDZUZ0yMhbpXoH
TnEGn3Iv72Khztx2qtsguuyy+z1PldPfyVaVHtiqCqPRCIC6+kH40vwcaBiK8A09
uL+llmpWWCRt1uzxaSOZX+8Fwk/zMss1t82FuRRLGmfErO1eveIJ70Wls/Q09XTt
/kvRLJL8XnfdMmdoB7Cvxg6smAEuvJUC31zq5ZPBpkaefPfrBqjt4Q/o6O7yXf57
0i5Fs5gVaq3nVa1K4zJNWgQE3VjG3m20bO0dCQ+H+zKEvNMU0n77Hfx0UBg9Wybn
CH7uCT60df82ySdp21waGhIw0bB+ILZmP2yqoSnRzff1RtWVPV/0slu5G8rCfLXF
HgNnbYPKJ5NRvyzotvFa4RKBWrteaGhLoOcSmR/nWP16RYbBMWEi35WI8eXcqBp8
VDN2brwcdxMfINXx7fqogA75ue0AeMZ0BfAyc4gcTu70lx9p+yB6wAGxW7Hoe4ze
ldas0PtUW5lwr1Aw/NrAUXDwkZc1rcGXlc8VLdgdCr5f3K150pO5WTy3vviM2E97
jQkzfmA+b/Z2Nrk4b6qoJvwIfDfaXsIcG3wc245RuqKcYYBI3LLlSmtFF4kJcZWY
bhzt5atT7cUq+z727S6bXgVLS/aO8vOxrDj62kDAMwfpmmxAPVwAKEcJBi/zQXDy
Vb7DgWhaihMSVjfqqZYuPnjPx2Fhsrzo1pPmnEZQMG8RrUqFzghLSd/Jt5jLClz8
zNH4tZ/xc0//78XLA0P8jghYqJeKYCkpxO951xkw2uU4yE2CUZYuI+GMNFZKF8qW
jnlOT+BhxCGnzk9smszrSDgoqdRuCHSe9xk3iGRIF5AN2cG258yvFi5Mw/dYIbbr
LNdW7rUTxqsBvxsq9NE3bvxblztSJ9G6qvrFUVpB+8pV/aOa89D4J9F7EIKWlB4c
U3yrZiLeUXI4uUDeKHYpIGgm3RV4CJIYaHrEBXbvyGKAZHYgYkbuoC+6bwXWW+l5
N0oo56bONyQZxYGi5GpJwezwGmAE33MgIBlgot6HyUh3VY3aUHvIxp3BXMgX6bwV
LjDoAKDGQyhnhXZVJtkGlbLNCTWt80oLEeTdiqO2NNZOQsOH8zWWa45RJsHyOjB/
DIEWFdFOapJR20GxB6y01BiT86qkly85r9M/CJT5wVwKC7Uf2o+ZDfy8FRVZSX+n
SPrdZehw4LiFE28RLpIh24OGDRiuYs+0m37OrMojKgM0qWewjlsJS5HNXJ29YbFh
CK7dXdmKqQ+B7pw/9rUY8sTtD/xr3lphKAdKGlAKhdddVcIk4Tr28S5DnAu4K6C+
sZgzpHed4Xdg3VW/EjgiMdgeRe5ySDLg6tErCh+UQyGWSONG2tGjTxOF8qbORen7
KVj4Tg7bUIwmnCXodImHQk8Fzr5NWwwRjnFHeDx3Pml641d+fXiTUNF1io2Jsigh
uyZHsdw24RYu/XrPqcSQcOUh5BaZOQ+/t5UILIiR2XqCfIeBCv62dIVfXhysVexX
xUtfOAqsDsAt+GjwVjaCr+x0o9Qxv2CTw7yOhXMrcur0RvY3B5PPK2jWMisEJeef
AyOHQWfJpwP76d7fv7IHcDwZSQCG7/nHPabERtMPQIzepQZcSzH1z8jd4QyZ+eb3
d9tmaZSO7TkmkbnUFVIJ35gQd2LD62SLq/ngCE3GQb1BZVvfkDE4WWO6BE0yEZTr
VENzUAFMihQxW+JSq3Rsbg01J8lRoD2m3r7i/nhrArsoh8Fug8BwZzHv5U3ts9Sq
Ou8fIxKsffVqerXQQwPGKo/HeQUIdzVRk9ym9g+uRZ7KmRN+YcriaTB1fwjHLnz/
g3wsP6TRfRz3vnhTzGszatY32RVvPwTaUlH76tzNhEJOLv58cvcwXd9MDuECq653
rm2hH8qMUD7m+8GzcdrkpskrOmHr2+xXt49loc3UeedjRzHCc4TbegkccpIg+Bhf
rpkvhh/XCp0eLzhhlNPkGPDaMeK9YigK5xLhvcI1PVmUB69+JOSb7OZva6/RijLJ
kgrDz1FpAZlqljllh9iVr2HP/DPIh0x7+BK/ZCctSsaDwHjxyVVsUtbXoOp9YQSV
FqWeHx9tv1wc8ykHq+iPVAqf9CETMldCPzrEIxr8/o1M1SUuC1WZMr8VtPhkao+b
QnlzJwsiBT2ntVsHMzULTEbdXjbUMponDtECSVolr44c13mrMDm7MyM337sbXba8
+HRHsmeoD1UpcdPDKSeEjpE7DMesR2BabAm7U6mKi+koqD/sFQCz7uGFWRQ1rxz6
sDLbO8DNph4lA2Upj8Z6jB98fXRCwUGTqldQ1QpRDQmtVS63uKeKsFQS824Aa28Q
FJm1AUEQ8jofJJie1zRHJdlVk/3fE6aHMEbZMTusadYQlxywZLzwNr3UGRnI1Ahy
kJMndpRYNaxGah4NEPWZREkwXfKwI2sPJF70vmnSahhZv4Lcy0Nik6u4JPLCMZ+j
AGqN//y0dQEmy56vi5dE9OE/zlQ2Y758TqSIrRmqXeV4cFXOqnghPibmohI1G29C
ZiwWsiC3k8r7SULPaqniHsuAqmuKW6XjpCzTNXf3/mPAkSwxI2/i0nqS2zkLSsGA
sfTl3B2Ew4m827Ke4mft7uOlihQI6UmWEHgJqPAM0lE5+ty+ClDcS3Z6xLbjVi6x
lRWzfmgSqIaVsgs+2BfaifU1sxFsz8xDwk9AG79dc8ZWgIogx9KdLaewDR4xhB+Y
9Zj43PZuOCLpkFB8ltb+NA+smAZbPV0d9wDzY+BakZBJzPUyTg+jh0/ycs9peCFO
g2ACgegCF7A9db51rRlASTp0dAsnDrbmZtuSSqdfl/ykB5MSubUR9ySlW4Cx5pt/
lwCJ27GVGQ8bRTosNDcEENsdZo2rG6B5cXJg7SnRsmUU6TpR/AhTt+75cDN7Rwqb
GcSOuIYOGGvHcOyTFyx3ubo5RfSp/JhO5TLMbGiTO1AR5uyTCp6PAXbAbxSRQAd4
sD9Vs+04Nt9dpu0XbrQLCVD9OyLDEa+EE50mt7a7EbhZhy5CdAEZTq9FMXYN6NY1
kPHTE/NoOXpZTHAqaoRENG/vrXWTdXtoTeP4AgzakLCv2sKTE9E6WdNwCN8SPH0k
kF4hDozcG2DeTB94Zfo9d1BIJXz0wO/EaBaD5CiuGB81wJCqgp87QIw0lO82lfiV
NOihph3OOoDcjFN9EZjUAKALG26GM8O5KVddwA8m1JDxwSbBahIJplFoYn6157gf
j4AuRGJCgZqsKK05yN7uoTCvtb+PBRNMv9I3yu0pPvViodfZDtgEDZloIgkobRC/
QLj7B2PQriMmJ6L0pOxSclT3aHq+yz2SH8sj/DIQgl2ggfFhtSX5x5ZutRMJmoos
kcRCHCeuC9Thwia5MglUrMiwYDCcfeQAGLFgvVbPk1IK0IjJujz+s8T8qKjPkwMz
oXAPC16gD3jcxTCHKa0lOmDmVjk0wsXQC2a+T8HXLzPAnMDDBsxZW+64oSoTQkiy
l4q8gZkrfp9CObwEC6Cp30Oe5iJeHNADAUOR0WUzoeLGPc+x78E0JE8b5s1mqY1B
vseAUl56zQMPT4WnILk0/382zf7sbDPPuia5u8auZdwzYOPJRQ+JjLDvTZm/+aeb
xtAhpwFLXClgYfeiQSfCjL4FT+02P2q7TL71OLe6XI8cZJ9PgfSv40iLmT6OA5c6
ftVGSmKUYlzF/2wbIDltf0LT9sI2kXFZ1qp/jzVFe3HJTFLhu4czxAa1Wyw/NKa6
OqultuuhhVdMFvdz8m54/k9codDLywmz3xBpiF0jXzXzv5+J2hfKsPJTS/484VPT
EhaZx6jwCsTEXZ8pxctKXG4BB7kQYD97NhuTRKj+6RDX5h7x3y2AOd0BpRGAEtsk
NPpL5KE6Jk+v5BGUZssCe89yxpknFxiL1kMUA9w9QDjsaDZF/ZT8fjr360x21QKJ
n0ZE8M4TTz22zJh79GaElGkyB18BbrXTqRjo5ZVfcGT6mDP2BfaCzl0ni0RRMUF4
5fK6i9AV4efhNcuo/mHCH5BtPVQzZZc9EHt9E4o/C5RESek24oP1rcOix3djkRvq
cvk5bLcrBEF/okN7yKhqbzb217lPtUjiopdg/SsChAwrFIlx+XjkI89TPTxpZavd
eKTsCyncEMaZYfWHAJO8TOV/XN0EFTfnZHvqBXbm5fUGNudgOnCKgm5XHAtALsfj
zj0ST07+yq2E4Bd5fMyj4DceH0deD90UQqYkXykUbwgv0/cXfaQPahrg2K0Nw/zv
yrSZK7gK0qCzyErTyCrVXMFOcA71gfQvTUHMatBJSu4lpHC6zEdeQ1dMeBqUOz+i
9tLHkCMOJ+G5u9XQopwGiQK5qhOqB1vpMSqWgL2gvcMtlRQk605cHTOkZ+f3m3/X
rIm5iiCy416CLmG+HW5934G5YgtPImRr2ouGGf24QLukpnYPrqVXWbsUS+RYj8WP
3ORAZX8U3mb++0dTAYfle33uU275Srse4fMRJHCZ166YHb+wclUQAEzflm0LF1iS
ccT4Rz6cRyfwZcv2VJkryM2e47oatOiwfMuIPIX+04HzGlX2q3Pa1dSrqemKG/BI
nYqljcfBrJ91T+kY2V1Tot8SH1+Yu6ltcbaWVyM/GcwlqX8eGZKEkqiDfcK5d/qZ
UZzWLid7PauWZT2f06vBiiBe54NRbYoDu/1DajBJXWfhdgvJCqRrXe14/SsJGZ6l
rVgkTNiiDUtsp0nNcVS8LfR08IcMAqSfAvIc72jJojsn3PRiGZ3yqqQ5VTZgEEFS
9OhalhK5tMbxsvDY50KwhYDjrNYr2C9dzIUnMpPi3yB4pQ1ef2MehZe6zlk16Kp6
GP5GUdKnagP+wD8EmujJPwdvP1dUw440/P+qFROiJYziCfbZPAySmZ5OpWLh+WGD
SgiEEjnTFmRAKoZgnpJCpw+CzOIz41wCcms51YHzUc4FUv1e/nB9llm/8biLcAKp
GbhKqzqx7clGZ3LRHCPHjtAdTPYk8JDxFX1HXyJSZXCSp5FryHEiDRkHBLPqzhdj
1RUUHTnK7cot6bpsuLbIMeIOhlF3CFNjbgStUkFpq4u+UdPE392UCoyq8TH8k62V
qAHatyt+3FLUqlAm/QAchs9mcp/HHJBA0Kt+WRsiV4SKybneRjw6f+c0qYccdxrf
dO/4Bw9U6LPNWDyDGuBo/VGDNfX/fCx6Fw6J6EJaSuK9Ya7jSeTZ/vPRhQ6OXBDY
dfZl2gBSRLPp/ssJz/6EGOsSF4KCJfaTKeRmf5PQWe4OSqPVJNfUgm8vKYSXjkMn
q1tzYuWMRz0PxrIqh8uusKoMS8fmy3yFr0CQk/fvL5Twjq7lUG1GHlHEsPwTxf0X
35ikmiuPaX9PT2VjkMASd22NGOLg9A976ncd82nUif8F7x+cZQySlooPV8XgQ1Ya
sHwEwMuYQuZElOBjzv8PJNW/0aHd7iJ4w99iGy5VC+oJuInWyYPevOoveqPUloJL
/S0B1iR2DzjU+07FikmDiVTq3TVNUxJAcDbouK7y4CVGJpJwODVv8QZrUaprQFRL
FppwbBWG1mTQXFilq7U1YBAEJdiE4dlsf4Wze0/Bafv8gw9SuN9AidUdvzpHO81/
FV9LNlIV6rohwq47AEvwmmdwAmgLb8WSuU9sXzkcq2e1yM45+zcpMr8ZXtevHlHq
z2pk0Cwh2UBxq6pr1pG40H8ZupB7CbTpM4EhO9Q8RTSZ2+S2F7O2BqE5z8zjfpae
lrn84R2dSyjat9E9xcUqQA2Fx6+70Wq0IZKt+5VaetJO9cUwmpJ0ki5nsDNQvmYn
Q6JsBEtTdjg1OCE2fJvkkHndrulvUHd+4oqhnRX2Onw1VFKqkLqVh7LEojYhlert
FTzpJlzXKXlyeNv+DHbPNpzl4F01tTK1smpIVy9YBM7OvRhrrN+22ZAiFOAaDrQn
qpMEyPW6Ky4mN6ziPGXHl20f2Lnmas5cj8gt8UZ61IGlfm0lH24dXaSJ/w0RnDzx
TC1J+XpqDkoWepM4Nd7NLspV+MC6GSfOnMC50FkpTKWJU029ZERCgbNvvL3NFMIW
KuZRGktVSRLJdkkpixnJcZGq8wfyHG063pZvEFPLSRydX/Y4KRKtTamzk8N5DfaB
/7NzvzX6jhNUow4rsA/uao4kWraFRGKwQoajqTVr+m+8SDraL5vK8MgOQFnLxTdp
3wB3Q1NcshyjArpvtNkTo5/4a3oGFypEPpCwjkgH9l2oiMjuVGYRJwtnvTlw1qjk
xfwEpuFByn4Gjx0W4NyPBaKcNE3V5JKHRKVredNO0YZJVrQ7OtHxbbYjry+8dfv0
tTxwXXRWtR4Z6Bcm694bSrJjzM5eXz8KgenppWvaDFbr900yQ/U4s3kLHJC+Zo8g
oXoGpsstfVJRA0Kas8wxB7EMzMW/bo3IZXP4nWVYJi0wyZHe5A/RCUins65b2cV8
xbrqNXOyZIux9XBrQvMd5w75+l2wovG0QbxxIG9tPAoUkNxYPColLYOfHukzqiWo
XRjeYLAG2gOWQbHYfRxlxoqhXKrBgdgX+fuxx37730SRrQqxxSXZGNpDG6DuCB3h
rZQtaXE1xAf1ioA1ypJk5CgSvlIxwtJAdcrkNvVzhsI9zgkZT4e5IbE7RMiY8d/k
In/dLNFqICv0yqBzWXcHEObg0gvKbLalIBrRWT8vIlSzNhyNR60aekJvMM/+/KQP
RojnGr5iTcNPMwft2eiPVsX+jDIFhhp0R9AZTYFCqC3xtwxy/Y3WqPcHxJAA0TOP
6eHukB4xNHuBdZWJw9N1pmBeKhMTQL6QV9acpGrhJVEk/oPJcmm5IYQ/356R3Hx0
Tib6rRx/yPPQPt5S2XD2KRUxPvNETteGjOYfsF7eyb47osqRBkQA2cWaC4Nzeowo
J2f+EcYADsIQZbHgB7o+S2PtWxtLc//3UfNBJmDv9mjYlWBjBnC93mdfLo1ixdSL
Fs6i/hc0L+hzVr1E+mqgscfC4F/yofE5zFV/dG+agDtvsc43HsjUdxU4d5+Z1/xt
BLuGqkYRfecNI9E5xG0FXVydQARAu+/tiCpvQhqI+bndDgncppZGC0PkQpZ1LYy5
TPWUNYkEnUgoyFGSF8GDDRVjSirbuxTlEPcpz+ax4eZul7E0g/YlJCcB9QgZevHm
+4xWRCbSbTyA4TmNy+v2NwAU4F/oJqgPawDo/WNLCUZ25dpZmhVb7nOWGVxIEoNW
yQpxP3FqoCSU7OljvwoMZq8LtR3J6gFOTLIWrcqC4fuZGZrDxgW8+VbcLItxTgXH
MZT4WvdfVhM8rw3YM9oUGMPWE9t768IDCwKZyIGQT777sJNh+fGN1/SJCJqfZ5h5
WNPEVMDiTxYWkBGksvtYgSdOsaaSv9Slu0Q5+w4GxjlMX1opXyGdEnfet1YZrUTg
ma5X0mUY36mBKeJUA1uVcKVrnba8tDZXRMaYK+0F4FqFfRA/rvij4XycHa+LBkWy
tNvVU7yrKY2aeMFlsEPjyO/qF1h6H0MoZRkorukUgEzcCz3mP+jglhLwNEHHx556
rMpVrWTyOjKTU2Rq6IOPMcAvfA3VDHP8Z1wSfLNAcOoptZ6H0o2sshlitW0bmoC/
R4ZpySz6s/7xQsmdIhecsPeZsmsdZwhmQKD62oSbL3ltphTkzNZWshYV72xO25q5
C+Jj3i1wqRJ9u7cY4yl3IpLp3iTWnfsriBdiOhiWokby/7MkpCnYtxG0OdH0dRjC
ZE4kGJL0imsmCDJAbcvZdzUXy6W+Rm/Rfytk2d9lrjpbZWOJZoe2lmawA4rDG8PW
JOYo7DP11rNBX5Z2eNyNWJMKyPSrZoiTmeXT23MsShMhozB2sM1K5WRyAAt6BhKr
ei474bx31QataQ5GYtjHSJOxizxHWzTkTfHqAVBXZ0FIq0Pdldlz43PW4ZDAQ6PN
qBfm0Ighnr1Z7BU0TpbWmdhPEkWLCulCGvS3zuOABoI9/OZQrvMNdxDrKr32GA1x
gfWY1ggXNUZI2hpSSvtQ5KhjONQgKFvr1XDo0wmLVjiftmEIMnB1PT/H49Y/CO0t
JAuDiSA4tA2pEJaiPJ8qwXGwR+qE/QjbZq9VRWkdYQvnTx2fQ4yKm8UO09703rbC
bdRbG299UyXW0Mc8IoG/7Sm3eEusHa9ZLikdRONourltWEzmsrjAzdTZ64EFKZf7
pwW8kveXylPZ9Ri5BLhP7bi3RuBbl6UiC7Gi9uT4PxCaPmzpVSHwiYqa598iPRHp
cuPNjzSZxdOSl6+d4ER2yonQ3mv/YhBPhKTTqydJ3L8Rm7w1+KsHG4XiKExdaBdb
keedvtf5nYuBkuQXpGB0hgOdruhoE72uaXvvvQWDK5w9eYojCFi96SwK5duBPyUX
LDHZ9+ul+sFVJvx0ZlBR9exxVlFexIzkn/qpxLL+IXIs4LQ0qHGI0OwEHcI4kFU8
ZXbi/hSHQbqw5mhCu04vPrvDMFBQtm2EcCo2dBbzCsv9y1r/Q8NMWhxIOeoTeuFY
Sx4sICVXqUtLifv2+E9ikA72fG5l0igARNpzdaIgCzBbHBRK/C9uLEwqwo0fWuF/
auY4P+5XtkN4UeqnMEw/G86wEtB1zQ6BaeVm30S7YVtlVh8UiYbLGI659fjwZOSd
AvlZ9vC+qtXIt4vS5JBsIp5S0NRD6VRiwZtkMN5pFj+oT4INUhNh24Uhfp87mbjb
XT106ofGoKGQ0wtj2vvjVA6Bhe9yTWHHRaOL454bguSyzAxQs/T+ajrA0nZy3a1E
P+PFuuEhknGDfnwCbf+Ojjt2WBXw6KnGLFZY6m95QIP9NziLt9/RQJK/A6FXqeyh
6LLiwEy/p5HFfc5kumrUi/HM9QFlKIZFPLEMiAkTUuiJazAy4x6jhYrIHewFEBlp
uQQ5QyCsTNNDQjjkoo99AnD66TCp6JuvMa/r2SUmt5J6Un8jUO8PEXwnP4uStub3
/iB9k9BrBlUcv8Mm5C4aJsnC3pW/SHdvkLQeSu/OUiLiY17yS/+BNdLO9JIKiRJC
LV999h7BCS1YWGult0Bnh0ECaBmyUXySN9S0+HZwiMJUvT3bqv2XKbEZjZ6zaKpe
rDH8o15ChRmp4SnBStoz8NnBBhY/K7iZVyrIembFfAwQHQBVGDpo60OrdZiGMYLB
g8dviBxijNCMXHyD+dtNq5kU2Fi/HdaDeWIQKwN1EPLzLf1qGH22wv2wQGXdAeWA
NqnmxWci7LtTPmE+Tpaz50OmhTus0etcWtYImVIozUoaQ4KBbwyc2NnFr81/ZeTN
0G3cpOkpjOxIceJ5aCUWF+kjTuwLmb+rElJeFc3ehnOQtoS8gw0jprK7Zuq2GMdx
6Qn0CnmCZ9Pss5KTKVHqEfVifGDpPeK0LQDjx+2J9WiCrehcrOYZelxmohfqEIyp
LmhoJ5lp//m+PMIrfZX6K6916UMLBEjrCKglIXolvLKUQcvMEmL9tbrcNRlkdgZ8
QwDqaVRw6WfrcAISzjPFYfXMJcPzsnzF5lyGDnDxLxIbqc2WAEX8ZRoly5VNxsmC
nDShZRcu6zAk+7WlbUyPKZC9pDHZCZx+eHUvgX7w4Xl/a7CdEeFBsafzfd/x3oHW
gQF7KqnWQ0+8WLpn+8hKlWXp1YuESPvXomkIB5hs/Ichl/1Ebfwyw+IAY6aoxlZ0
S+Z4hXQGJCIqutpr7WSDgTWjKHr3DmCvjaqcHcgt3aUwyPKEozHPh5Tmj3cksYRu
NuXf7CeDPEy5vwatZHBIotuxMG6TlLjAJV4P9iZ6QpTgfZQdNCQwoRkjkS7CIyXQ
zZMDPvmLFkNIJ2892yhGwZzU5Ij1TIcwhTc7lD6vWeL2qgnKSXry3h5bm5yaRCb3
7y2wCw4+hDeUPz7sRsxDlx2ABSy+cRAL2ZiVTdeif/xbg+4ruv2E6k/khuV6Cg/a
n3rqFNxWj497TchEl3vTb5YM4bEUOHS25m5Qlbd1CSWHtkwbFptemjXK0EcCKmez
+ffft87AT0+mI73tAd7s/8xgOcR2cb9t5SW48++UvwgEvsuevnf/KtNjZgJEK1vB
whJWzOW+QjjO0JjD5blCuJwKpb8lZjIM8hfQcJi7HCnxcXxbDvpuf8EtCbXq+6na
S9cAKarN6E59TGVzridmdFtE/oreHJC/BDudb8I2RdII4KtBUf9DOV/a4NbBB8nY
RNO+Bv/r8z+e1EL7k0Yt7aeh3j3azfiSty6ZX6lzflqv9WsuVcwwHnnv/Tzp8hi0
cAxCMODCbn8gSJqC8fZpjTBYk4IocbMutQ9xi5SOIhkyK4Dtr6fBGhpSNe6GORuS
nezc/fEmCj0xaJ2ekrB1xD1b174fVmRx6km29lKqIPNGy9LU+ysdSzahGqeS9ghu
kmaXij8/xUXnkG8jzVMZK4joUrh6VSL9/RaGhu5Z82pEaqQoNKkp6ESYgHNIp33p
6r2a01/SdMXmSI2DC+UBUyigLhuhsdbt0hPy9uSLT8vOof0TrBZKF+75gfeCrHat
GrfG0e/gM1elv76RXVE93PxSxtvX0n5zmw10P5tlDRdBu5lzgqwMzwxbdcThPvhI
34HTWGR3pMH0H1dwD7EDMW32Foe5UeRb5rc6ujVnl1T6ovVy5caFJXL4+SeQ0fpu
OFDJqwlNvpczrs58nVgNLUk4G0Nh+ayGWrPIUW32EiVG6f8J9D7EAg4QJIG2jTb2
F0K8EeanaOzJivpLJg1aX2nKvRuzZG9/byGPXNpOO3Cybo1kwyiKerosNmN4YRS1
7TpuOykjWcmTclS4hCCW9Rzr8eztIPK55P5N68uTOcGnZoazJY5uiBqvptGdFz7N
nnsI21GmCz8T2IFZFRq+s0FBWpITfTtMniyBR33vtRIlB6Xgykhs6GCsEVkwxEt1
P1fGzWIsU/Dx5SXZ9/rBZPAIL0Si+4yGiXl4WU6LIL+HT1Bciiu2WD6A9XQFq/V2
pXwNPDNaUx4MEMkGkuEKC0x8fTbhS93ThNkxPThRn0vy4fTraU1RTl+jAaSremVq
LdOvc4oiP8NKt7Qp5jX+7eNZFquZyT2KSrzFRq3Gtf0D6iOVq70zlZzFP+eJdbDS
VLGpLpngKa3dAZrg+ATzI4G6THumxLBjO82CGraTemxxtLV1lh6D2KPBBhy+oV7S
BMCftCXFwx8Y5rP1ueRGPdb2pg0Gh6/UiElL+ybnTfzr2KpuwBUigwrtoUZcX3Mu
y920GRuyGtnYcnd96AVTtadFng7DyoUS4wf0G9zqjzcv+qVC+i1lY08nLSyyuEf6
gRVMgtpcUJ9x4xuU4JC7t+lR5yIKt/vNIYL0g6c8cQC0wcBr8QBYfhpsTpa16LCt
S6RAVIcSxZi0yxSNcx1xCUetsWhb1IKpvg52as9oMx0Dy+H6FT4idP7k6oaqAoL9
P/kHp2eYFcmkkG68XB9OEbmbgCyANe5n06Xo7o0ik6I9/vDt0kzJe6PfNpLlLN6m
FE8g+VEjPSV7Ynez0gfM0XZkR8+1Ahx2ifaE1SdGk4k/TUF2TrgAzd5sPvcagHSM
wDCxglZNJMs9uJ+K+HQuHHn0MtD3H4hFQdt5s+GV4DWjBy8VG8N8TD4SrWGZXRuB
4ly3qKZmC83K1BcO49eB7AqFd3FwHleKQCk+jg+frCT0JB5SUC/uvkTC8isE8OwE
UD8fHnhQd3v/GRf8NbN/tvNtf2szlKRcwAj1UAHExzgvIMgJZIGrkyYP79mjyM6s
HePJRDwNwtxEsjsu3/s0W3I4d/3vB6QXelDDyiVcy8KSkOu+JZwadXdUKCrWmOqa
so9Vs39GXXYN+LMgMxfyE/xT7Wj6Ip6/A36ZMJwujsEix8sdcmrHN+Qt9tlUOoVj
VflkGgsHT2IoKgoImcwUIXxJ155eViPkhY6x6UbrbvI5V2aK3AUKyhlHp3xTSsTd
HsbJx5x4E49USFCRkzLhRjUQh/tsgIDde6vdnykOSuVB5TkTNgzkeGphCpf4KQty
8O3vEckUtQxE8xv+Fw73q81w6pNL8kWsvu1Mk/jwYcdev05cR9vviHZUNqqcQHTM
dbJyufBq3axBmb1SkL/INAbw+Tr1F0OB/Yc8u0FJvB4HEwiaA06eJo1jjyrgXZly
4zqYsBDibE2J731GMQhAo4zyMbuoZzsMJdo9ZI43eI0uZrX7eL12AI+fEn3JoZ6d
7Y5pMXEpX8dGMToZv0V2jnOY5fNXPFGUZTF6JvlT0zL86km0YDpkkxdx6zs9Da6M
yjNDOJ+ZNR+MO8gjNJ29VOcJ5CyBR6hChIU/FuxBgyfqZLzw+Ksi2KF57ey5oyf9
HAipp2ZbuPksRfV3JoAM02Prn9eDeCmwrOXtWrvUcSxDPcr2gE7RYMwEcMm1Cl/0
Me12DX111GHen4YdFDGNJUHa+parVz50WT7UbR+eEyPMd1vQkj5QxuKOBv600PMa
msbloQDPXS5mxhbGoHc58EI4jHj1GN5TZxhZqIZpwMyqS27sjJ7Co0SyYEa+gBG3
ya8Ia8PS+URs6I9w22scv4WeUcakmV/Tpi4q+ZCmSpa8w1lcMmZ0rdVxMAczDO3k
dKi8thtjoxl9JN/Z46QVTUeSSS72i8a0Qjix2rSyBb/+ihaOLYB3gwLggwxT8UC3
JhREdWJ0xmogNr2bMcH+Ii5HuJr3PyBViHXNfbSupnoJWo+A1LJSP4IfUcwC6/s1
vQCEZige9Va/w8ue5y5ZuWaiNKRCmyRHiEOxLBA4173Mr3NOXDek5yatb5aTJZkB
Cok6S1pMeW+rXuBnh+Pt8sOglONqxSRMIi+syNKW+6USBbFac0kjqzhkjvJNjEl3
lVFjDGiBWToeEQmX9IU5/9eyyP91iEqdwX6yHImIFh9pP/wts4DwMQSwN6Gu5ZvN
wEPYTDDcu4H8P33AdeW/7rBXTeggDfiPhW8aYMqGtmKlP9H+DIwdnQQtWNhHgvXf
4bjlMACqZrBDxiXOEXXSaVkq6W3gGRQu5EZyBxZKqnx7WgSm4E8qAdwWZ8Uzusic
gKpsAIy/PEaaHizTzcfeJNjGLtbiiDzTsfONVEYVDIlLfPtv8IakG+jEM13b5UfP
kUeKGIjT4ZloGNno0LeUiGhvtmMymydW6C4dTCT5OI0wA77s1Ou0l93l97kkikbV
BgDyqegG6dOHMH1ogXxBMah1binfWqHtII1G0Rhcob/AQP9H+cfd+aVGyPNXibtR
KT6VgZ/qkoIiSLHzlrrwm8msY/WfOPNmRkdB1zeapM1JcJrP/5HAFYsSKapMec3M
OsKHU2py3CeJMNkoAY2j1vJn/J/v7ND5TzQSylBdhyZ0DWlwKCGI06ofdmyLrtQr
6FXxQqlmZ8F4J7MIxN9sB2mhJWuGBYowGKyGP9AuPafUZFEc7sH8o9CgeM3Zn9z7
7FxbipnT+qiP9xE3lMIbKxjtdzWv0y9kL+DiO7F2WIgMaN7cY+rcfmha0CSjWqPm
o9eCE+GCRnyx3VMXCMCQ2Dcp2kz3p++LWbBUALlWjvgvEfoGNMn5Q04J/A5/BCef
p1PM74aXavprJos8CZGjfVPGggpK0mapOH++SWTZc411dLgyRPar3q4jBvcdxacv
IF92jpk95a99pLQr9pBXv5BzZpy+DrI9rTwOw9pwGeZWPlr3xH+E03kB5DllHuQc
mddJsBRpaaT2K9IIX3EgV0RDaNiyTuGkMkhwWlbYbHPcGqppXpPHQZbzhJqyJyDb
Z/qLXHKpkzkbmleBc3nR0Lg9iXS9OK2CvesOF2vpiVcQhAZhLRoFlS5BJ1dkFxqd
d41JC6inil4/RCEt7sD00Np0ZJXpRo7x8Ahd8+qUCub/bVNd1vJUWrSg4ScBH8Uc
/DtdXC6SlPrxHDOhGjFqY/dDz8SFtJ7U0YTUJd9rrUOMe0sWL6TEkcctLrijgVu/
TolElE/0bw/DSCNIlHZrW74P2XFzSK74sR+6lcGZXZyfWF9JqzSg/lp3iP7xR3LS
mp6iOL1jIrkfGUymf5vEmNqXYzNtFPB4vvBKHDJPUdd+9dN/B1k4GEcZbutRjuU4
FR5KJkHSLBucDf8JAQqtdEeJyILaoV43NjUdx7wr64FtIFee5VnDF0e/XT453+HK
3+nShG/+llnMru8gHc+zPzpz1VvvrGH9LSHHLMoYwWsL8IZ85Ya7ChEu37Zo5t9C
H9RnZ60eEV8IwhqJ6CPYEnJu3/MJt/Qx5ha13YEcADmk7XtJdWaLZdbzGqiMmVYW
JuYBFhaq4LE+ahnH/YaYamSAJquPhfWSy+oTXKm5e0XMkHlQHjeWHP9x3e59TSL6
jZPM55UZr0TeLwKXkbW00SncaLLBkD/sZdbEkAI5y2qLeNq/fyse3t2fQuIU7PBp
sKWt1+hyY6OCV6brliN18Yyvhnm+hLc0nl0ckh2Xbk3fJXFl5Adq7L5flvV2vvE8
v9XDKW+RDh0bqY+CgsTI4yEFGsUBUXShU7BtFQlgXxJeZLd5RBBFUzPCjBEgvy5l
RCdotbfI2zAY22cjxWmnihXFSmkxGucpF18qvG39o94fhy0zGD8aIXIrkYX+YTMB
VylhpZeW1kyb/dD3fLhcL+wwbwBFyOoPz0OeuxuNNHx6NQ+6fPXN0yiXZPLft7K6
T6ZksQ+BaF+cQp1/qMwNmJbNmpOfKnB9NupnsM5FeNs5FisF44RO8cAxyI3aZC5U
PsNpFugzbzTLSQj++bK6rwbXgS9TawSbwCPYPl35YAn/UhjZyFA4tCeG40XdnPI/
uKwpQEoFFxFUeVI3Ou4Lma3eJDALBIqxtKeOlcUFxw9OiFozLbm6YYOY6lHAFLES
ER9JSyZRsMZjKLfDV3BSCcRRCYCvumZ57AjER+GPJuzmyzLBYWUXjmES7iJTDIUB
wilpETrTSdFaudKaISjIHqCFvgwFCQznRbteKG/aOVfLwhLtknj9bh/xtSEwJ2WU
nBn1mEwmq8PSQybyvpD7Hwx4/pRCWkL1qM4XFjDHP+1DXFwbcJawAshuasWyxnEG
mQAUtAx1SuQ7webggbtO23kHqfFaT74XVLlL1/pWT647bEC4Quw04xszOQzCTDzc
JLjkHCpdZAQEgTBR+ifqXf/euTLc7kbbm1owLu33lkJvCaF5L1K5Z+pnTc9b55/D
yDge7WTt4L5V+p+D80e2ro9R79luoBYFxgAaM0E6O60oPCmalsrfXY25e23QBxTO
XCuOzXxoMTcp6o7NqEDygtiJzot6yB/X+6oJ+Kp7l7BOmy35q8CTQxwVVs1+HP6u
JkVLcZefcUNh/VZA6h3vREt4UO9vp4+1+cS6i7mpGBj/4c2MRCfum7AavvEVajJO
vx430AHR1fzNqhAS8zKpxfmdubF25Nvq9dzR+fkHoa0fbRG1lpbjNU3Z4OwKttxT
xE2qRTmmpJpc9L63BRzsdR758TNC5AdNJh5v3UYB/vtSKMPupyvBj/KjWcmeypph
4pRFcRgeCRMaEj172hgGHXwo7ntvi2EJ0mZMniYHNnCKJRsFGE3+Wad7qoZXqkWe
TjG0qtliEJ31b+rJmW9WG94M76VmiT0nBPeMbHl7Fo6WVNURMOotZ/4l9GsIZSan
1VdxmcoLms0kPkS4eIKGtUPXh4Zbcb3au0ucY6jyJv77GWam4A/DLy3oe9VsmqwV
qwPeEJwm0m+AG0IYvzIlamC+sQL2r2Qkl/TYG1eKXFEjGkoqOZ7yw3C5aRBHO9zl
8iMsf/T+Bo/Djxf1NdZHh6zWvRR38o7xmpKvcL3bex397c5BcKxUwL1lCADDzkfT
NDpMVxO5tVesE1rRV29p+6+LEZlwblmuyQUiCkqhmKO9ZVHex2ph/oMJWjmza1bN
mpusLgrCK1jmfCosgH3JU2QS3f3mFD+20u8up2FKQOmFBHKSisJ8T8PrHrEUff8H
te91hWa1I63VfGgTaUaUo/GY0cYWO3stj6Y8TAMQr2RbkrTMcMcLCN+ZvsMazSMl
exQMCepZV6O4/5/n0XWkOikANbfshJVARAoq0e0YWgQVsM+ESCSHzVLjfN3TmM6I
h5YGELC1tGucYYCIY9dAO0XJmDgypkVwiz+5y8Zo3+SV4lHPFQAGhgDzF4+jqqAA
iYZwCuxRX6EzQU2gFlFigCW563wjQwrUo6NI6ILFSCgsEv0KpTFN7Kq+AW6z8xVf
guIQSLmE4vT+7DMYdhijnn+VUsyEYch5MMaL4OQFnu8Df76xy3dOea8FN6/u4upP
GLdD5OxkoDN3NOJtNZ/JvxwpQXT6Z88MYtt7/4gnhiSPeY2aVgzKY4E8Jphe7HpE
nyPjkCRzvpwB7Zz0UMt7dtMU81kqIHyueo2u3uYnO8Wfwa/vQwfaHN8+ZXGCxLRy
9g1afyZXbN5x56z/vHdcJ3xBnIfxHBfjmVIZoK7OcMOEqYJzxnn2oGchhdZ2CCNl
/0REg5TtqqpSY0dDEf479NykbpyogH7+MJc2fRNy3gkGMbRz/PBLn/ixidrj1g/4
M92nR+zyQwFJfsJtxoxnqQc92s6PmJ01OFG+X0kz6D4erGi693qpHL+Zhh9qTG8Y
S8HPqRu+A/rTNNhOGod6rNs4B6MYaDr2tznApn7vWUCHRLnH+d1da5bJQA0AREFT
mHpmiFOUqBqYQT/aZ2dwH2TI4L6nxlRajeKTFR2GBxHVVb/Ic/z2QR0/ViugOTUy
tZbEtZx5T6hNjdc3VOVv4iqHY92CxnLCnCI46a4jWvf2FgY9e4wqpx7yAsraBvWR
du/9CKwoy/vUp2SaC8buDXlWHIvKa+IeCi6ci2AChFP+bbyUxOiPuhCie/HHdCKJ
NJLpepkeNu8rHkaBewgmVzKHyjiHQNDBawmCuliONMH2ayUHAfI1thH6o1pGJs2p
QChInIwwYaL8T2yzmWtHExqxAA8IQ66us+W8IVE418IXjY7r6PPdMQfzJt67Wk6m
7Z+0SBcU5QYOt0E8L/eSjvrTLbiGQ2PHzUFf03hGnnFyDYkWfdpXp4t5JvXnRcmh
lHSUl7kQf7iTyPVAq2Z104JEEGAZ4/0KmwvmD+BzjrHVQjrdiPnXmWml949K1xAb
3tnyZ6DOgA73UW/lKiwSj/h37IeUzh4km6LUhbTBf6BLFUEX/DgiHhzSUSez6f8Q
6FnVDde46N5QD6iaH1EsrVnoB6dAn8ZynpPDDNxgLWCKbqqFn0PFmHH0beAoW284
SJPquH900Ntp5jGR+9fapPWMfIVuhqd09sE2UT69VMWE9myK1/TtRKrL4EOaW/V6
ZcyBUbqAJDltTatL9c/Bcu282A7iZIe+to8E/N69L1VPlRDZPVjMaODP55VyRyBN
dV6tLFIKC07uVh4551WcgewZuN4XLkcTKMAhEy477nSi6qELjsUgxlRDnD1BTDyg
fw8UddMrjuBy67bMbJypGZHnvDUfaC2l7L2M/kEHoW8e9HcomhysOtDDvbuiGXyd
Op3oBqkMqnUfj9SIxp1lrjqjnJzgrx50qhhKfL9HWWD7cakprB6eCDk5kUD7bTtd
fBJPVX7jAtpwCs5i15BXhGklnPrW2YgS85Hyuh6CzfUSaxIxD+UgWsLKHRUBy6xV
zzj9MIBWRNCbiqrxf02OFIFTqyVagxWPXDTHqTNTcULz06JxnOBAqs7vIBHNgRKd
razqbtRIgut35E7HRszlCBL/GQS0AT1F5V8XMkpW5SC5uE8USWO8alLKVq68LIrV
fJHbJDJopuqn09cyoqe3VEu1MnuhLRx27IK3p7jwA62CTqwDWjlA78YtERN2ceo/
5JIREt1LJd+XBues0oNWIG7057Omhxt7GYeszuFJAA4+RCrnD8ILQktaGtv37rV4
Yqa0v8KQimKgho0oVID5iwPqAdUlYGZE3F1xz3J3fxVpvVEe7pO1SrkYyhZS7hqJ
XHmUMjKDUsvBxpwVHA0KggNRjaEGu+kjMhptELQ7SlRwZNwxF96hjAr411F8Gfgw
2GvCbX77k5FiIYudVY28rHUEg/B45BO3sxTH26uCvWpQmjG845hBfBL9/CUoDE+x
P6CBtET8F6VR/FS24SUbAvshirfPfVaAX/O3/oJB4fCHxIYZQjL1dIhg2f9nrCgr
RaOaZFiOO3L9foGLyr4TEDGAammuPe67kWUlFtZn5SrTk90d6L7CoBwWMWh3rdMN
P29gV034bDtycQg3wLBTsAHj/QqnIKLJEYXDhhu3CeqdfSPoQKMgvkKjZ8PTUveN
dbzOW17p888eJSzr7b0O9cdL1NFfgiLM0MD8KulgjhlIdSDipiIas7Uqm9a9l3/l
FPLfzw/0vE0OF8V/6Yz53YLTmam8erIT2PuYmleMLLwqA+4AHrKrLNBczhBP/hYB
p3NmgeFl2JuEyPEwLtIHAaMaivMsdqHWFJdHEHbWVMz9jF9UYuzGdTCy5hWfq1gk
zz5FTgdkVd/7kEa0E5sltuJqSD/s76KGCdc3WuTVryx07aBCTJGZm7LSKY59x0N9
LgLFA1OLdY9CD2bGbw21l2ESq6pyvCP1xwxa6TRLHOyQag+uNQ0qrdGLupTfBEYe
wcQVyGzLR7JhFqwheVLAtLDwBGGmKtoMrzkVW6+4IQDYv89gae455EEBYpXcHvP+
aAv0HkDxAVRknJo4f/D18W8UK+xXh+88U/aDJaNQNOZqbDW/tgZ36Frg1c3YhKxR
ZQzVNPG49kqF1XdT/VtcnPhndSKnc+P8N8chcKrXxWWI/mOcssr09XKVhgcessIv
e8Pqb16C/c0+Ybh/RVVrkbhdj9uE86CrC15JsV1BdJypruOgG7ZHgRzKXoz9QeAu
kzDl+yq5X2+KQVxM5rn/DY/2++1M1EtHSrfD4wjWcMyVwmFBfbEqiJm7K4+pREKo
iARm54Au6Bbp1bythpUjYyGjExUx+Mu0q49Qqi2Udq45GmDyZR7mLRVMaFmN77BW
aeRWlkEjjLAnhvLaU0X+3v9R4YunKWTFGEC8+v1HtXMtnBqKfOf9c1wq39ljvP4U
VNIR0imweshymG2o4bXQdVostwzBaaJtwn6RQ1UC0ZfXbY7RJD9rVkO0m4SVRv0T
6GNjECOpFksx0xzNaTUR5durcir+Yqq7aJ+7m61+Svlk4lYsDV9S2RoR1NBM10H0
m4u7x83WAtbQJ2KWLca+AhnOivqFBBGxLepeyrIWQatvkmXwKloCrARpMPO/C5hU
FR8E5UDFxlgnCHygi3jMzueYSByQ9OEuZW67XdfMr18Z/Nzbu9k3+BmrE4ZZ2Qlg
7mm61RyH9N82eDS/O+HlSVbQyII+iCKAZJtfr+PQe538id/8dUWVJG9nwh42GKWq
0PQMrSg+52rJ7GABDNzmt2dm3zq1xPGyEv9kGfUCuc6oixE5m9DaAuWCt0+AyZit
BufytqbhGp23MILpAean7Il4iZ2zPiFI6J/h6RGdw/A3rC9MFJCchs6pXZ1s109z
m5/EYGRW1+OGv+1hEeGBl8J8ZLdJqlUwBMyTEI5N1KovmSAkXZ12dEjQZWFFKOpi
AjjTciTdIWejRTe8dmFjlmjBvtY6vqYS3ZweRgxn82IYhTI0ZjEovLvZhQc47n5H
6JNz2qISZzuqHu+2wnScoDFEhRlpRQI7VtrqC5xc7eCV7wmlmOA0Emoy67/zVdzs
QEHO1RlR2p/pa1Hv9WCZwaWBLeHWf8q0jAOiQoRh8DcNPyBhzkWu041wD1v84AD0
DfgVeDoCmm+9xHUMWrisQQfEA2V89Wu2Yz2ZOI8pWHXW2qxR+LeYqnrYKrLN6yXr
NFe+vmCHzuZc3X9c/dEYNOj2r4G9NSoDQ0PRh3l/QNfNXexLgAvGosXnIChz8jB8
SWlsG0foB6wwWCYS01yurdBq5soAt2JB1NWYLi8gQ+mSclxcuG3R1xi7/2sv3Dkb
osvsYO4vQoLvPJoVwVvgoptRtAgpIHQXDTDfT4qX5YHH0MrLbTLvb4cAvUj3cmmw
4jR4kMQYfxjHrynuXh00Unnz9PQ1cam6r9T3QprHjOG8EzKBLIYnpaZrSTpXvJfi
g31vbctoWi8RfHmkNs6y2jq0eKGRe6HsW7kKGBv+vHDqUOLfcAgTyqU45fRcBbzG
wQEJnq1WTKuNG6e4mBXUglBL2KyYmDMGY3O//Yp19ggPzWeh5iFmdHcWwOouIckT
OIvjYlfbwp6r/pmnYoOH+wvgUNffz7VebWQYoqJTMoH03R7YvnSmzoXQtKKxZxRH
e6riTv4z1VlwN3SRdybDTynTbYVt6LvKIy+psszg7J/pM0xTSJqv6yxVYRJvMddy
bPaKu6YVGVq2exQZ10gSutFVHH68Sz3kIaWY+XNAIkA3qC0DOfEMtgWGG5BRzNf2
tmzAmRdI+o0F5iF3PoaMyZKhSx42ulu/EoO3+MSO4IlcPd1+HL1oZFIQ/5Uum9u0
koVtyEAcxCU9F6b/Orv8itQBoS6tH/5KgNj7CDyMU/awZg4gpRiYP0T6hdvnb+wK
igXYBcEG/rqmeVDmnnxvigN5cRlSDGDh8VbvWBgvUqb3US5vVRDIkvSPMGmIDfCT
1U1bbDY+1EFj9hPzTi+805IieauLminPgWBscitbdM75SFwVSdP74m1pGbCj4iWi
HIpB9s8yFhXSf4FRLoy51Wf2rBMvRc6qNu7JADksInE10oey8ErDLAnh3Hcalih7
JaY2wHHn57ds38qbDegNm/BAZm1NdNfgc7TJAsRKDV47s09UPKQTyfdz2XW/lnjE
6g3V7utc81pQmFs5/+3JsCf9td7F+2680QiAshzLhn3dVEtM7aL06k4BM33N4yLv
s0GCrvmbKVcxucbZEe/RP5kfWCqUm0fzECS0dJnVy9gRX/tUv7WhM7Q3+wt7YXwN
yRcjAx9pUnNR6scNybLBkOdEXzfHL+jyX1jJ0AWgD/E/RT8nPmu2rI31Sy92zUL7
Kuc6x8WmV9OcvdVKKJLB8XItt2ChTokqdFkTNYE5aSVji0WWqeM7w43ibntpjX9s
beLkkk58s3kcZDbiyKJ34nVCR0vZb92zA2oOOX4JfCzZMKT7FsKYjatFlOKZh++M
n3BYiUGZg0OHTChQ2oSgJv376xcC2sMxSn1IwEkgaea9s108Yn1UTXmYJOlw9nE4
Dkco57u3X5+Cp8+cqlvg3l8kVLdWNBIwgHya77X8hmrTc821hJP1SSJsfH6Z37xW
pmpuCiWa5IPbSP4s2nvUWgH0+0aS9yX/aZIU5yjDTWnIIfePJebgjt5q/RBRVtA0
5egr/G7lhFtSq4a7tPXRQAT4ln5v5ynGwcqYdmiAO/5qTABIx9v8NwcG4kFhu9hu
D4jjYn/Gn+XKuzZx4iQsq6Yks49t7K2gIZeSscHMRDJGEvEp7mLjtUiZYmq7smS9
L83g/C55OEhxrQCNW/kOtpUVx4uzUw29qaRGjo4T9auH4a/eBwbN8fOXaKjAhAcV
aScOH6gWCY4eTUvyqZTY89xoJiHfqtcZIDk2gjsqrfdNCBa33W4y8rjX0bjxbgzA
06w9USSP77svQKi/eInWJhXFtXOc5gb67JFH/XGZpGvrkFuIFxGsnMJ8ORwapHXW
i40ovHr40Tq8XTxrOSYkH5w8ex7axPl73mD5C5Aq8dSAmqVIyIR8WCMQVmBXXNQS
C+cgV8Z4U+7pNfZhMj6uqU8eWrEosiO6Pp0QN0ZhY8hmQvml+slCtA/pj10Oh44A
VWc7KTEjyimBnJBmqe6LfUM5X5AFkmOJvxykFdwZSkX7fyL+4fIMPTf/pofVm7ov
fHLXShzMX4GjFbVLIp1SskM1ik2FGo3F8WdNpwDecE/jFwzjDjEe29fqH0/bn8Y8
ueo040pke2De2BLUAWEVrPGOv8UA/4oJbxlx9lI0llupmXjUe4L+fPRM59IO18Hz
YjrBHFMQMCQpKqNniwhT4eFT5PP3uYlLWvRK1gKdcTThbfJxAx96KOeYisvw2Qsg
SCjbpm1sE+1K2sr19AYKQNf+hsV4LbaIoLqxRyiQABPxrf4eJpT3MUeULjIWuT4v
Ut9R46h1CstQ6LgYbmpqwUN+Frcx/cXdnJ1vtNFspEU8WSWaTh/MOLvgWp+Gndr7
wov0wbTlEuyzvr0cZHyGpuJOXKdL1dH+BO+5ghxDeInhcEdFqVZQEQEm6rG5Z+yv
c2n+DppZORIMIvBd8S6L8V3t4m8NTeTbKYuylqSc1pfDcUBvLJ9E5c0Laj4eq0gV
f+eR75eeA7h+qEU4/mFYuPQB2kYKeotriMjlLF2sIiy5yZbGEjkXLjuzkc/rAzwS
aSZRoZc7LB4kVSwGphb+qQFkB2ZEVbYYG0eg7i2GLd2VJbvyxD+uYUxjP9cQyvtW
CHv6Vmm/RHnzv8DTCSpQ8GVZZzinMT2QD4VxlEINEHqrhqyeTXLbL0Gg90mi9M7U
u2HWVOBOnpHGtlGFnpRpHhNkaI0PsC2yAphRT81MWS95u3zxOUOoNetIzGLOuyQL
rgWL8WplmqqzknhluCcK1dkqZy/GRY+Xhi5+jnf0b+fiPSBqVNhoasLthnzNT3Q4
4FOv4jADQrksYDV8SUzqtog/lcSBs8Hvc69jIUjXSOq+C6LOiZevup7ecgyQ/w8k
mzAEuZq7lSzhCYrf57GYNYtV5GxIqui/5WIGpgcqMXBqE1RdM5Gr1mN7OBSbCcif
pjs6WW29wDjRPZa0acvtrwvoPiMJnCjBqkTt95/DpPGvEDet4QMm8MXEcdTtzhM7
YCOtQy8kBRP0BRZQTA7lJraI129ySCTdgyOSpOOVxUhv9+ynrJtyGK1N8F/6ctu3
YLSFvO3b0t4V2o/tYJRtimGR8kdLniV63vnaLwkl4bIedXtQ6/EJ/XbXLwdlAMqf
uKZhgWIpfEvJdYWO6L7wX5irD/nH4aPEHry0sirm0gwXMwxVCpk3uGPXk184JJV/
XS6t4KECaD5iSmOf9U2gqB1EYFKKClrmBTE/qITvAKkM72QiD+YgGuoAfyJvNMzv
TZ7rYQ4bkwQn3J85y1MbdqCwIN0LCa469q0ADsC3vZBTrBZ7yIQrkXU5dUkNf5ag
91dtO3tvNBK6HaTiFywZAqMcbvjnAkBmBui67/ReyAbJQkmGJ+dfHu2Y3DyHd415
Jvl4aCMVhGI6KACIQ8JXSoKKFOGvCZKTnlccL74S71VWAl+GYjOry0bjPVFAuhcv
FvXNabV2mxc3utgXeVkG64OnYb0kk8QLPH6Waw/ZC0FjuAvanDs/AaZ0u4CsBV+U
8wQfo9p1mzVSfSiDWXcW4tEdeLbR1R4xdytn2+xoDnlAJzkDYCbJdr7Hy0IO6s3E
OyzUyZz1ux7rOnVTtI3P6eXxHSTL2cbbHsh9G4ZbRWEZqyN45E7wMrNf2kKN3Kj+
WFQwBlOwR5618xVxoKyQSWZpMZYhHwntiBo21lijG29tcM+Y0axVd0dPSftR4oZr
Q5NjWLICfxKMetaXrNMRN3dnZFxy0Wsn8GUENkXxh1LZlEO20MhMgq5bdZjEkdSq
zpJbgfokhvPH8NKUFZYYOHJNQeQeDuRMNwSu6yxTfm0Wz1X3QLRCYGeuMSr6ylSv
CUQG3gmC0K67KHyL27k0nw/GuKcah9c3yqTp5gHHo4H+B32R84rNL2OekrPqHd9o
28NEzlbjuoHWasuYYRxUE56hpkyO8b43UKAZHcOyadTSYPtpL0YxqeG5GxMSyqUV
7erUxLuP0wOj1pZMYNs4sPDfMRjRQ/OT5ug768ta7XJtoMoimHAFce22wh9jJpnv
6GdH+SU4vcVjPvwQD/ZNdLtaQ0M9s81XaDOBZPaurlX8iWmznOK758RNErUOeqmt
BnDjYmppduza83tNIKcPC2IWW76gMaiXyvBOTTMKbyWTk3/MhQ5Vik2wqjjV7OW5
3p4pZ4nLGEep7lR3PRJe3bqTZylevDTXGfjicrZArzSZpPbUOvBCWsnmGvTEsOSX
5rKIw/TXKWXCveMhEHvZagmKQekx/USFDP6+wpUDzgKuEJbBxjsilXUUwpqfQMnn
wlM/gFFj/393qZFoALJDO0KXZ5cDVmbRMfz+GRvy1Z/0qa0a0d1oV679EZp7kWCv
ji394dQmr1PAL9PA3BeqglcNgy6KT2Wk3DmJCmbNlm78oq3jRDuVtCdCW6jiB2zD
xsk/YbcBHf7aXIpKmjUym4aDSbgpHYi90znFz45Nirg6nF7z7Ms2GnNzvX9cToA+
8LiKpRX3b+ZwoVRXiW5MPTQVRuLz+MBefr4NLMkDwmUkzBt+VEdGCECCLWkLe7y0
osxHeLezgsvL0DA+QsxIUo9jUBWbLpZQ9ERzK+dql5rehiOE8OKi8jmQs+myxPsj
xQnR+quMmzCYewVsluNN8bcz43gHmxE1BfUj20+IFGHY9RbIq3b2nYgExvdMtPao
K+0Go8nHZlNH3ENywlbN/XRlE/FYfIdBuyVxoe1hXdxk+L2kvWYeeQuJb050j1i1
GlDyujZ5ftiUJZG0UhPNmpnshfHArahS6HPsBR3PwEk/F+PRQCS0D2zVSpL52+gk
FQNsSRWlajz37WbYdZ8xal5XCCLFfwbaNuhev8QtjZGlaXRlx+wGE8wv5PxYk8Ae
srkXzxWH5KdBY9CoL0gUeArZVs+wJCifuoNVotPtpuYLT7MXhUFpWP/M2lIMFwmg
b74KooEbSw1V6rvdHHWQVPVJtxSvIJSNFDMyqBH9mu+pGnzIlf7IjoM+j1fJ/E56
fYcvtxTsBxUv80tmh6EiHJ7Mk4tPTiVJshVJjjWuryorEbHNozasaWYl8NIjnNTW
XceoepCIcV6pdb727ms00PF4mQf+N0LkCQDLq5yNzIsQXUAxA8natErUuMHQoBtT
cfp6+P8R+fDlmGf1fNiMRiJMW6S/wm4DdMP06/Sotobdgu8Hib4AbQ6649Usdlph
AtCXS7PKGMeiXgGgr8Z/jC7Ca1Pr4HVkRWKby+W+2PA8fceTv1OaJOn6G0y5FCiZ
bjV43oHWOM40Fn7BrwdDiXsSHvXdSFDUg9v/G6xD36w03OT498H/oO0WM5uJT+1v
2PPB1Cahni+JI3UdKkPDOOcH6xL+xeE9SOrTU4bXuIrAzn9+n//RCrC3l66G3XNo
6L4Gw9C0RgI+ofIb4R2UMfTU/Liw0EMpXf8G5fiKccVbn1Lm9PzvTDHQ5piYFP9L
BiOqeQVvvTXuwmiHz3TDGyXwdFuMHSq1ZKscx6CiVdI76PtoU8EJWPbDAHklKSmt
q5hAPw11j1tQqqLsEj4G0IL4vSNXEt2Eb2sASnYUasPg8sWEZfyvo24i2emftRNo
Uga0pOaBYtt9Pc73Im1nxsLz08VV531PVDvtaXZ8wLXEywyJU+0Zoh9AfavL/qCU
G6ZesJLqmuhE0kZ3IUBLcqgDvk6hFMbVU2gdFy2wysp9qlSs9sxsZQI/PfaFVgs7
pVWNgTBozeVvpigJga1mVvyxESUWxLCCpeLAtpQsS9oIMlDH5y3sBGBMH6MQEZ1u
kFzubXyhR+TawSZX5aCrPHkciNG8uSGFr8WkN8jGYGy1Ub4iIX9RTYjuuhH9hIzc
HWRvqe1NM9xDL7dKcpO/aKkCoK8qfKjcExy+jSHj6iExDI+vo/d+M18UDiD3g01T
a6+OCfLzaL2B0XXpkXF57rLlzzdg+FCSSUzEUL7nAnlq0rJ2YrzuBeA4vPxPzn39
osURAWTEB3HRTJJlsrL205Ewlbv6ETkW0/xFoIZZ4YraaW8fM0nPIlOSpBRgBbKl
d51m2rwFdl0EtxuNCEWbIv/PgZB0YdsDxtDNzKj7+GNWfmWzP4Pd/lGvQuH1krWM
YLiIVvDteUygdFreHB5dlg7I8EfvallXISNu1mImZ9pHVGp8j02WKg/9/WHdKoOH
8Wv3fkziE2amtnVFwrJ3cM2ByIvqjY3DjbWFQI/nw3kDgx7XwGvPzANlj9aJJten
awzc54Tf8W0GWYzfJPB9kdFHS3Fzv8mA6ZzvNJuCuYh6chNk7OJCrHqz67Jt17A7
VRs6qrFQc9tGA8zrx1gaDHQNcr/OQZv2y/STfPf1c+cVEo8Ses6+YlhDBBblTZ3l
UpLXEKJsX4vXlFaG+Kbu0EmWfRevHcRdT14Hk7nAruKoyEUYvIV8gphk0sDk8TQB
kvJzgrmMkGug3Uim4McciCLrt1qTFSInWx0wjSaqSVs0O2INoAGRnuyYqu33/nlu
c3EpWoOsY0pGF8/MF6vWs1jSjZ10DM2n7Flam61GAq0KsvQ7ikHk81/hE+BawMrL
mrWrdNyM9dC+ahu+Z0waznplRDWithB3LqLmydZig6LxOi1s5Mbblhv3ZWnPB7av
uEYFz/Ii1OnhH57GnYa8PDtecVdTTIJ/Nh4bQvG5mUN1WKs3vu0DXnNHPE4buE2k
PMPJKMouGj4SpvWoUp6sNp8RYBbsp2VqFrhgw90M3GfeHfZWDmoHrsF/ZT7vmtkZ
VJzQSGILLGCLeWfhqLP8EUlPrgqZoztPr1Qzt+9dT8261/H3+A4DCza23eanyN24
3NSv7CpilikHqACJWSfQUau1yvW6r0plUXMmUFcCgSY/Zh7jDGCj4B/w5cinrKvW
DuexLNUFApmvyr9v2r3gR/M7zv21r/KWcBSA3564QrQd5qe1yjnULbpfq3e0EOql
Yim5SzMtZGWNcn1SPg4RojquQ24NDH1lTgRu8UOeyKIRhOEOUuZookLfa91DZhey
JdiUO2dNlTYcTPnIPzgNAhJKJTczpmJRE1kDxkeRjj3c4DjY5/X68FO20AcMWjWw
ONyV8MKOy9Rd7cM/6VZvrI+NYGaGCk8xUqbPwQnaO2wupLG3+STb87bVfgyyf3VX
DOhaNRIwXjzTzzkqzLLV/FIViqTL1PYEEd6lnhX0m9/4QAVhEQjTEDEivoazxFeg
vyPmCe9fijiUIO7i2YrxaMf/N73dkBWOkju8fWxQYKGLEjzZnHYnAFuV0WyFLTDn
TFxEtwanVm1OH4UICs/2RHdkiy3A+ZCa2GhpAvFsCRQ0oA5DfNP8QatvO5HETpl0
bikuwGaObd3LsjwqIdE2C7aZLFtwHTHCRmqoPcO4vplPXWoW5hGoVtivQmEPWh0I
nnygBIOH2In9HAqQbou4G4XicRjGVEWxHGZJosUeeYsTsfI3FhojjdqMrBkorOTZ
67sHCdFQ/1oYs9qlHWgule8Pb+s70fM/zE9C/JSqwUv/pizmemA30b9AEilU+sDl
g2oLsvmBXTkxtFR6j4/5YSXY2hsWmXdWtNjB3SKVNQx33nkHUxngZU3kpKi3bS8g
HTOt1+uGpcQP+1qoJFIhGeBo55i8+P9SaRPom3hLEwwjx/2wIJAVBRozRJ0bwdw6
yBIkX8DPkq+bAG0U/D1SmEG0wK5GvogDuIcIVeONUdDKuNFjjZh3XUbQUq5Dr9Zs
2GRnDneAJf54tEOxYHnQQ9r66bTzkeyf5neI+fut9/GbLUwGvZjWd9klYwo2pZYm
9IiKB+atwH4onpnHnTG7SHC2V/VG3314e4SkvYEY3cEj019PTYMHBsMfCr4/bnMR
MZOFbYtqqCMJPgf7Dsa9Mi6s6LylqK6eC+xrCjuVrnzJtv3I0/xwT1f8dQGGzAM7
r/bwiKjSX4nbTkdlANNJJHBsfb6ejJvzpJEZIGzI4m077JX5OaFwJyZIJlRCwYQA
sJxcOWuBEWAiTodkylJnpY79MPL9CDRZlfY9wOYjsJQKJl6PmKFgO6539UXvzhs/
z9l3geZPFBynBsNLFcOH85txmCNL8OrcCgCHAP53IBBOBSDxUjtcVFISRGStygpw
oIba1uJF7DcBhdSKc+AYruTqaEfpQm3HoEysrtvbS4v5PGYBeV98ltycAwxAYjyg
CXllL2aStiCGy8kx1MBTKm2YBH/e1Kh1lKcR4iB/K6SqkHJmCslP1Jy9lVEBoqpQ
ccNsw2tARWgfpXTTndVGSVQTilBuvDwSKXcLWWn/hVA18BEYjIKJv98Od0gjm2SR
Nh4pkTjHoVNzG0NxebU/Ei9ib1LlIs8t4Jb5SbIQxJM8/Lbo0Q2QPhV9ipLoxcHm
GoCwyp72NKSDiHLY4MgPBQSAbMTuR2cPLe424b7ueEGFLwT4VOeB01zI63zmPOr9
nuOHelojAgiaSUGke/thzvNyYYFHegCpumsgK1psW9PIEc/DQIkXEAabUu10NNCo
BZmqt0WgEKY33SqTwVbf/2kJz7z/UYHCFug/u9c47G/i0iqx2QGPRQ4R0kZDWsJE
6/eaUs7LG3WhNaldU55/3Kd7xgXCw0oxVQlCbADGCWi3VNe9wJI0j0yiTc/drMGw
LqnaLn0gSZHzTngGxa7Q/Na6FZDyjVJHXC4Ohd+eGixUsM4EcN4lm8HfEcZfb8vJ
kZrBqgM+iA+gZSl0MbphhV5QXTckA3MCIHwgq0gWSM6ljJLtHeCajhbYMYUszrzK
MVNdGdcJxg/15KpYlJLhMU+zjtxB4VfLsxd3jiEc4df76olhxELPlY9hUx9iKC0H
g1otTL86AHlPLI6raaehqOlYJVZs6QDhc26PhHIqoSN5POabWlUgVpU6wDN3b+V2
vbqzAP72FbASjcTrIgGnTL00yWhXQobMTlNqdjScX+UbtwSNU7sO037hNf9Ppbmo
ycc2uwKr2U3lXhQ2kL0BSf/QzBPCd0r/uiBCsRPxzfi71lZCbN+JSY1vJkxHt6co
FyymkPu29EdegrpwHltk8/uYCsuscK0cB1C0QyT7BJM0XufeajsjzthCLc7G0+Sc
gDCMS0bG3YjA+nFFCLYhxvaCKwOfNAagTkYn2hUV/jGAe3ukUWMBJWyYjqgsXwn4
eC/IKqAUxKpva/Tn3GNoaVm60SnCh7h7RoK9eqMii/yrWI7nmmpsDw3SX8hJF1qq
MJFri22QtmGtEUvaHM2g+2fgSNV66b5sB7IxZqAmMeH3cBmTGeZSURr7w1gmN5Qm
LyYIlQhr+FGpF/FOAwrDkkhdYb0R08xZP1kSF1YRUO6jk8hX5d4JaDqoijEk2JWy
5z2++D97P2rbUt3+lqkoeC5mZTUB03iL+PUB+9+ASlN/Unu0aqr9Sp3C0x+zt5iS
SgQPBtheym75aG4Hne3+bzRR0vF7bkvEYRHqLCCV2cvZ7gzeASFNSiajPs16Zhyl
tTeXjSoxFbMSD5sYHJ4b3fmgXHN2q8cITKedfroh1g3Sx0mnobj29BAN4iQ13uIw
z9roVrfqS6+euF/wxZZ8QsxEPmfL3KpeiQVDEf6qkdQpCJmV8Aa3R9ljjjICK4kw
X5hWDIC0OpjIX0wNgEBm9orHI93+LuWxPwZWHXEW9MkiMg1/K/eqRYBY/uNH0L9c
0VW9dLwb79iCvycbjeSowpQXWgTEuqzU2NsBG//NP1sPSgUmqayZ9MknBwn9hn56
uJ/ouZ3zTboAQt5tkLw/UPo3ftNzkix5X8x0X5N3TWYux+vYaJScVZA5pWfNmn3B
Cs+jVgZ5ET3U3B1mauC3dviRoYx3Oskfvrs66uZD2hUsLyOMG+VqhlbvK8ZHc87T
50dvZWuppHNXJZ+nJ3kt/VFhimR93k55nCj4bWtz+PKdJK6FEuT5iDhXj/lz9ZTh
uoTkwYUnZTFdKn6mpIIZlZ+Jg/Q93JiOtnH6CJCo0aDd25gpiuTLx7Ov+v3mubtE
dZNwzdDpwjtn8VrxbqO1XRPDQWKCsdn78mDtAE0TC6vlj/PwAczIh2cGlRSSNYN5
i+gPiSZ1JNmyDYcr6Um9JAON37rL1Z2YNRXFjGWbCO/co5Jny58yjW3IiZ3oRbC9
nygLkJcDC5zCinxIWJUJ0KYxV2q8UE47BYZBUVyzIknwbp5LzmKWtFgnLn4oNubU
HNbrYd7iYulBe/6ZVxJLv4Hd7dNHI80/qs+xUIIbIT1NUpZ9eO2PhbYibUg1Cqtp
rhht/MQBjFVocmzhqvaA0QdbVhKtfgpJA5EJBgRbRiucswyoI2WaXhq8VH0hQKcL
3poZ5OfQaaS28trCPf8BxwJBj8EbgFxhnILYVLOty/9OlBM58jmbW2UUxKQ/PO/i
DlBXNsgUfxH4Z3EwZPqbWLf1sUj3THaTTveA7rlhHN4Q6TI+Isf1ZzY3wTmhxRAw
Z0mW8LDyw1ha+5+rdFD1MMgzjImtKz9XFsS2k7iqr4tS0LE0ay2kLKp4DX1dzfZ4
z8z7xZWKrcutI9fWF4u0vBpMfiWK3Dp1Q9RxH3qtAgdLlOdTVFGgtBAntngtG5ed
pcMlYLrn9WGfqpDSO6SiePpj1STzDPWs+KoyYdgJKcw85yO3QohEPPL1TJBAmCHG
OHebvuFj5AvyKX6v10370eTlnnWiaBD49GMI26AxbqRyF3oEZALS3S69bsLQ5uYg
6K1oivi6M1nAuZbu/uETbeFdvgHvMstCeG3TeEVHuMH6jKDObFIXmtVyFxkmY2vR
LXBA/g1ScvJ8xhNXzpp2pl3Eyv+QWZcWok12KoqNu2DlGK2QTRtmDtr3Kp7wVjV8
7zT771liaT1rdge2dntVngdnL/ubuc2HAv/eSFUM5gPvdiUk9HuIyj3AntKMS/dw
Bl1CVN+U/P1EOT5cWo1gQ/Nunm4BcjPy7Et5DEiRKA/6vozMDHbcnkGGImK8BkH1
z7OJGvSOQCKpmT7HQMg1I6SCvuYADPBItCsNaOvZIs6dgtB2vyfuUgUNoLCFyJQp
WB/gTg7J0tbHvaC2nBr9wcWwz59r3evaMjRqH6XQU2I+R7WunPmuk5Pt/R3bAVU9
cWWvjyQqx3+C0pX3RBwd4h3Jgwo2nFwLw61o/fQ9uXF/TeH1T1LV9lPXuvaAZSsm
7oZBANYS8YHGQdII9GB9BiaKIgeCi7xkCQMEIquLv/PhzuvUF0+G1TNnDmFLnmkl
F2dnesESkYXczY7ZciiQ7reeNE9Z6GKg5fsKyOPEnh4CGri1lNHJjyfsUFo8DaGU
nkRSKnKF1Uv7daQbktPm2ecgWGHSmTC9X8qK0CwqArtXBLA0yAv9qIvyLyjYuDI8
GzZ/v0AZNt7SnSl0nnDWOQUbmD/N/Y6rQhzcSS2PerhYzWNFwJLWc7qz+GxcZCEm
LX6Hpf0bG7NSCxLTHJ9tgq8NbyXpT73eqW4a/2KU04MFrXDrvgRhP3EkBeddP0GC
+9PmwtK5PNce9ibxCb3RwbL3f3DAiqOL3yHWY3QOrNRaakcamLkusW3Nk/GT7Nsa
1QwKoRZuH06Fhw2KaVuvTeXLMZqt+15G2XnFRvtgpe7wB76l01gRujobUbS/Wmq0
YTcleJaj8zvmYojpBHNSRGwPdrqeskSXXPRON6YZJEJautzSKu8VfztFdvGvCEnI
h6Ur563vWfpED72uAjCyWeYspQADHyNvPh7qTLSPScmO+tJXVrVV/992zBCwzjTw
qhwBi3Gzw/sQAd2NcHP8jxbSmHiXuuA0zPmEOrdjWfOCTI8/fJYQNED/oo4Anh/+
TGR66EYpBo5+NexkjcspUXSXiUJL2wLo8KnZwA4ezqHOY8n+nKDoc45EA3WW4K9z
6Z3JebYVX7dI7IG3js3AfFSRXyMyap7i6WoB7kiOYA3uNYk+CmFJ71e9NB4jXJx9
H0LO/gGJRQKQRNQRN5G9YR1ggkITlrYSQW/ZN/ytHlvi7jcvR8oHtOqPXSOM+u+v
GvSpYwS944cnS3DYx42hBHX8gQd/z0V1r2tMq7sSKfvhdbAJ5qzaEND1MQg62chW
LbB0etV15rbGEI6h0gsGx6sKhYIWY2sJv4VyLxcwR1dqFQH3e0Z7JRd8+eMG6p4V
dfm7pTLxrEiFLebW8TTa3iYci7WC71dmD5UUt8ljH5EB7jwkO6VvsDgMXqANcMUw
evsOSDRz7PjPjhPfU87/YpNl5auSzH8preT9CODnBzNfmbYaID1v3jVnFw2UVgAS
0GVUyOSUSxrGhGA/HXoDgppj1LQd6PCC9tc1tdJ0SweRCdwHsREZXzRXzBNZxH5u
CzhH1VovmXEVzkOBpNVgthkJZU4DS60J0KQXsFjhq8V7y1BwGBCiJ2+qmEBJwoDf
EPELNL0QoBn0//9EMle6ShOz7T+46Y76bHawhwFNQgQSBiV5Q64gZIV8HynrFa6h
PJbb6ucl/DwoAN2aBocyonuimSIvFJDuC3Sg6FmIIRc36MA3Wxg4nbWV5SkrmKG+
r0ZXctORySzsxN8gTq7MWNXBwH0HSLrWqyzFyPt6BGZVxltPBJXOLh0OG2+hNRyB
0T1r7Nj0THf9vdg9iGc+llCnij1iFp9+w+2YidQjOhSLTfoc7I94PCdhVB0gNZr+
SB8xRb29whcOEMKklt7oOhdqKcL0Pyze1TfiX267mceHnC1Bb7Osogt3YW33FSbx
fcQuo2alvw/o+w4qru39e7RELlUyyIbp5pri7O6BL19T89T8NxivIjSTSpxuEoIt
jPvFzoGcyXQJfcPbA4/GGWsgOeTykJ232qrtX2cduyseEkpdybHfFmOffEt7k+h0
+eYXtpIBJgxuTmy9kRnPgFsv9oVhKDrTfRjW3l1BhRGeIR0XCkdNfZGSxz6P90pl
S+/oPl7XJC2h6d/9bGAcj+9Newg3Bn8d996nAK9UujR/6Wk5TK3pfbrOyyQ/wL4P
n2oZOJCB++M3uXDglqCW6TdFS2W/3CRuWDzy3yW5FN9U/y26J7TsyxQGfpOK1lkf
ZnJOGIK/GaJcTHryui9kZaA5WgbbLT3be0gVU5w4JpaP4qP639kJCHI7qfwp5avW
JzCdvVedKyls+o92Uaj1EJ+kbFGigYbiYNZwpGjdR0/b1rZvEal/6dFL6cxtum+7
XOT3EUakYPc0rG6MKiBZXstkdLHgzK5ah2r1/q71kaVV8Oxco+IpuqB7mkP7HIy4
YwiK2pMRzM7XM6oUrjn7/vI6IIaBVK0mbSRTBs1VKg5mxb5UWmZnA2HggagqnzIh
zsNv1q6FjRejDdXTjwYyO4Eu4EnPs17+M/nbdld17JePpGtefumAXdPhk4L4C40s
TLQ0R/eRXxorXrSAP3eFJTQtfcH2bolxKmBPiklKL6Mb0l/+uuzGkeTR6aoQazZX
sl0s+TOd91WOSJ1TeX6Ua25vDyX2TTprRTexbRvWu1kAbltUzHyRCTnqNet0dha+
c3XJvJD5DWWU9mPtwddjxcPaXWuSDXBHmoqEGy0F7HUSu+RC/p+1Q+hBkbwPU04F
cCJghYeDY4wXwfMRaXj1j/OGHA65LUz7EuIfA8A5wS7N2w2uE+vJYkNFbdMLDahz
M5pEPkFmBcSyt1I3iQBrKrtAJo4zRFotMk5Hs3HO4T2rQC7vY7hV1PpUgVDbV5q6
pX2pzq6sMxB9QY9gMhph1+piKm2VGf9drehcEToK+gF8RwYthXJhhT7wsqBSlbGf
ld9/I6Dwvo9irW085vZlJJxJqdTSyF9Fde+z3DXuRfl6YNfLgNLAYX57cxuHRblm
PfCkJw/ZGLsFYsjWau+q9ow3rP1pFxE1lOe4LsuHdh1zFMHGYXWc32lWmgwpWFbn
E2SxBZ/S/SJQt+dGjGwS7fzoF+M+DRB2fJlI38xamSH+17ooRgVCK2278pPDS4Po
gZsn4S3Hg8QqkNCn1IkQCrad+C3BO+AellBnGQ3wdH5fhwlFzKitGiH6plNJ5uLw
5S7sut6onOXG330POpF+7phoxjWDhORxHtj9Ly3Irxg9O25HxsQTuFfRKkIPWyFN
a5vmZWWfaUUbhTHC/dbw0y8F/yWYRE12lkMdPThy2qqEs6Ov7NuEoHXkN3KXR4pA
XflQXs6ZX2lxu6JHGl84+72OIShmqBBlbOzgsCb/sH7R2XNcptE/T1DQ1cCXDnd5
VoDLB7sHvkQPlk83ZVjpxWpVA6wsBNRN2gypQVQvJEyIufIP8aLEI//vdruWVbFg
DsgDHnkcOR0fb1U79iuR1eFKnZ9amM+TqLOlu13jpTuzPxWKIcMQNL0ZOQif70W7
2OiyVHRkrg78qpSEchaVAWp/IL00KwsZ/KgLvi/5xrddk+Qo7m9STMTWHfkmGHdw
dvDTIDCqlHytFO46m8OljL6+YUlOHBf6X/aswoSo1w0hSHuJgy5ey6cNzrkvSmK1
Gc3kbd+d77N/HfwS9ZM2bej0ILQirbDXgX9v/v9Fq7+ze52BbUhC4/+zOEU/zmxJ
d3/vhPICzC6166bEygHhSaM1tN9cePsTX1381cXNlTbUbxXuDeHthyOrSA2sU3UX
sZIeSnx269I70KeQe5HZrGlQsZn1U88OrrI4Rb15FGDzLs1OBb1mXByQ6CkxNUTI
KFKZoGbLwmvcHEi/YZ+6bUnimucnfpBq1k9sTdY3RiccrJpA+F2iusprI+H9Fw9d
MXrMy4Ap5ws5Epjd5Uia53/+TcQ5yWSFmF076/nYd/jTX3xOW6UxNnAbmKlYSs6P
6wh3ZUAyj5MAgxMeeH/OuZYSM0/LzV5ugDX7iBUv5dwft8fHWmDwScyVDPHlDpiU
nob30sPAfh+AzDROlIV8iHjFI5oc+4o3Bz303/fX/2ZJCbzYYfpg7AfWmNqdQvAT
pnCrfe3w6TZe7k84PAsLC4G6f22qLnGFduvmCvvBldfTMrNNu/T9QpTuuq8/pkOR
5uCiZE1Z+2UQ+vsUCU4bUsr1LF1em/EhLJhGunC6omF5xhkJdbgLHw4nXyqagpRI
Ir1kqEVig6sjXdmboLGD+7dg66Gzl9JkgOCtugUuPVSusOM1d2Ag0gJy32Ydjq8t
ACGFZWXHztYF2xgHCRUGxefuANiUvpsthiHBMxIsZEYI0tx1Mrd66Z04x2y8ghSW
RhaYuQcqREJzJb3XxTwE8DCqh85kpVdjX/TKbzA3mlyaEmkW2CzIaL2mSmYp7hAG
uxSd2aAOhgoNpwAIK/WLwAAjZPU+b4ZNCOHcVOIAnVp8Yalv47CVygTofiI+kxwF
EpZLLzzFwmpwa2pfwx2VydZXASC42f3Hh21jOxcv6Jhc6+1JUCJfvSCC+T//vWcM
4SQVMR8P+JO3Gky94y9Ty02x2moU81y13a8yeTq8pPSD//jE7DsBgcu5jgZxFeC/
a06+lUbK1EvSVHqycyIPzDco2GTY9W1yOIu9UvM9+dyu46ZpYHe7sDxn2ruzgTca
yxlxXfRyPAFz44iBuGJO1Zxw0NH3bNVOxhYtVZSXkBFxVIDfIn4sJLal0Ofm7zuR
BcHsqD+/Yl/MKlkE+1YYWKj+LEwMuIfeAqk5A+bKvkrDp078tNh4izIytfYBN6lt
+ZPXTdQ4e8f3kRub8ARpeXxbEvv5gE+a4T+ymSoAN7hlDgUTUy6ec32iR5eF1PaA
M4xP3Va+ruiQfpDFqI6EdM+FcLHxq0qkgB73TUlcYqlkTR8v54yZXTSbhVEAKRRd
obKrNmlqYiPOUX7am2OMHGkBZb1+Z10TBQ+jMKHdJur80Ts2K1++5YATaca6rrea
7cs7/dtGyBMVMsIcwY/u/6pKTUo9YL17pFUBeqKFAX6jFhDFIRXpAB60D77+LL3P
HJF5eqDuiiIbowPO3qphEk8uEZCzvdpuFDy+Lo8/HW5iKuhL5Zvp5loXEQ/dF2n7
ke9txGyChbXgJh+IwL1Ae/YCEcjYKUGrcaqHTT+p8dqTSklNMOEnS08oBjEelGCW
UNXbtXtDyjg3BBLHtiD6LY6ruCGRLpBhpkCGeN5bGij5AHIgYGHZ34iv6JYOO9lx
wbUTCBV+US52S+60WtGk668CnLeTeu6JGrv1cJCS0u6tdu49AagvXrQ8VBkttWTZ
gm2BTVM7nX14Rx20vRQtPt6VpCpMcXz8UTbjX2o/8iYCipz+tQl3F7xWnzerWCaj
394aYfyFjuAd/JzsWJx+xMd/CNSxV+scA+kfA/1sgxOR1ajwaWhDju4HfoaYjFVY
9C7LV1yzUkRaDdY8Lwjqkkxjfsap4n5nq8Siaf1fpiOK5Vbf1DMxNZpq4P5C6+lZ
PlJRRD7m054AW93yxRXVhD0DC6EuVhQkz/5f9XSLK6Hscnv4R17pQKXwY7lhC4JK
d0Aw9sVY3PyadfUsq2Ju9MBsl6/ihfd6QrTuZLHfeLCFkd1XeQVzKN7CNlzU+pPW
fNoHWZBh7uO+EuYxjAPPrzOOfZvZNZZUTQw5PvBjfN4qwnI+9Z9814vr4p9gQdSs
COzsNnBQRsz9aos+6YjP80+I0s2+Nzl2hHwiEFYDpfF82h48Ym2dZlLyXMWUvUxS
1udzKD7l1Vlx1TIHFIxa6VGFeU6Bd8wjN9CfemEqc9+ZLLArl6ven9CmvEEEpY1P
YiEsiN1YCFm42rE4SWQwR1fp1nhSqCkjepFJt96mY0r56TqpRUZsSqhUlMZzQcJ7
iiWrCRDNHXjaa8SoSXHA5u0CQrspl+nU59B+Dm/J4/yxv9g6W37TQ+HV/eVR+8S6
LLMgEd7m0eyB+ztfLNoF0SzzY3cahUOewf1RQ3A/ROuzP/SJmJlXYpnqC3idWkrr
BfbxDkduGBkA6HU5+sDQj4sC/l1l9dwGGO1acxkzHLgck5oI+gdNEJ0KQ/aSpXzw
nXQuNqZkyVWTWKJegu0c/EBdUQ1eIKSUExyuYhPIuaixv7aSk7aE/A8wjdFr9OcR
iohhaixobD7pb1emP2C8P4i4nu01L0uraIWGPfCybmXd+itFi6KEXj7ILgxYpN2o
yBwK6vZBEYEp3pokdLXvFwytQjxCgtXHF0akb+KtS9oiEBmQDJGWEUyL/nVQ9iuD
at8tI4Mi08ZfIFI3Ogjhtn5J2rjJD40aZYiYCjAD2VBL/uvKbox+VDV0TfpksXbq
liSVINQw4zr6BNYFGIrH/OKEY7s6mBdVkYuBUrGcoHKAWgVYd/VPpOYrUJ+ULdp1
kW5Qiqe+dTVZFcWF/GQvEywxUk/ogym5Y7MiuJuzRYwH+Fe9aCSYJ7C4GTVrKNHZ
pmyEHV9ZZH2lY49VyeGbDWWufXFKvwmECjkQYItmYcwJOLhyVAkEgt09GjnNi5nR
p7b7vTPMPJMgMq1W+2nq3Jx1w/OvE9M8w43i0ExEJ6CUY3CT95F+12LyG+OHTlHe
V/DhVSL7oKE+QI8FzxFl0+B1axI2XyHR8YU5CfbU8cf9LpircMVoHpG2Kyabqn3x
xspsIdf/4fI3Po4lrxlP7B5ylJK2pl+B9lu0t3arw+1JfRyDTB1jbmWusd3ll/8W
HWh/Yb54outIGH+9Gr9Rra+2xYH4+J0YJSr9Ced2BgszIFvglKQW3AE5cYqNH/m8
+sUVIFnUe6fXl2qgMYfNU4NWoqrengPOXpbGRRJvoW+aKEBVJLxDsywJ8sYmEsmI
xDv1mE7vkpbye1dPELNS92r9jykXg7KQ0mIEjvSNiOAkDwjGNGOTzwAx8g0VVLsQ
ou6YoqMW7lWTeRgBUpRCPF/9XulOu7QrcHTGmT6LpDy49EIxYC3FcqolhN5zkyly
VkU7eIJXJqP1dNdCgEUfxqkn7d78q/OLyjYlK+y/So2EpBWrnHPtdJTOtUo3GEhE
cpz8nqmWixmw/z1r5Q2D1LSLVaTMlznBIg7OwjrDiyI+KPihIcg7XyD1oI1Ukd4z
FAeSOX2kk0yaSd0/82sFuTa43xf0ipTMEEUqLuUjtE+bFTqCzrlxz8fEHyubVSq1
DVeDVet8gf7xEvkihdIIs+NgJdNI6ntpDm7hlbJ8nJqIIqRSPLiXwzJ2AbpxmkAp
ZQALQSNFm6RCpzn9AjlmvY+MUwlYFpK5lALjPXlM9H4Ph/i0gLI0MDcNcpxdSCLs
c7RQeZigAXShF1dVfXQIiDvuDkzpB4n+0czk7yannvLCXpgJERr3mXl2pTWxVU34
nN7lg9DzlmeB5rl0JmSFsDUru6Ddd7eAckNWGN+k6g5QswlrSleP+4q8Vj1wyf3z
ssCE9+zaTzDc6LuEqmGgIlO/URHMfrWd27bFHwmubCyCPKpC1ICJZJdEXMNsiAQ2
UmkV8rt5nDeEz3QXD/a1JrTdZs2GoUzOYadLR+3dRETMxI123WLc+FDLQAellO4k
tax7N/PpOEbOuBh0G5KsVG0qX+rOagWP2R1KKoaKzK9EjL6sgk/ijoIwhYLybLiN
ZTDPZ865qO8kP+ubxb/gqGRZzz2zKpWeFgyBz+1gJkG/kFSr4MvTLeUa8F+046+e
JoPgeadlhoYZGCoUILzpeolzrK4CbNjJUE4TELf0P8m8OX6JVYTh/l2a6VS09aRi
ORS1tVJyMAHjye0cg3lnJlr6N30UnsONUxQLO+oW6fbFUQTwH9ZzTnsXQkQzKUDR
Z4s5TIA5uH173pZHZlLcNvLTQ3W3k+qL4XeBCMpKIoSLXGqeisOGPDvCl6yRPpne
Q9m0EN5k8NWe63ke8MpDSa4oe+peHThth/+nFs9V49cVfdBSagzQJmzI50Wy2TZz
4ey1RrawlyBbirlcJZtTfcOGmE8QNAWb+7F1lQIOOAKl9dxF/kFZ8B7PN/mHd/cQ
NJN9qSXIUITH9/eY4df/NWUlw8xhCRjVjut5ne++pii9LrCCy7IHiAXX4aAGSo3T
U3O2MJgaONQ35dtvM4UpoNWBBcbMy+SAAkT5/bVZynxMGP9m3aCW3NGw9MUElhWt
+PJeTNtzuBSgqj5kw1+cXN5KXp08ZVroqw8AkAJXCrH/HFj0UmqVwiVjXdn6Iqu7
KcaVxgfyiRd0QIm4lJO4FV3cawsn8iyLzLFgyKDKaVproFjg4Vs5NvIbhOj5fC6s
i+AmJnkz52Sx6Z3Gm7cACsHhh4iRO29dPdFJZ7RmjkDs1Av1+M+dVtEGNf32pLAP
FCFwPlTEagzBo2jZmif/OBVQrXuZvlGmlU/2iwNL9cvBMl3xWZjBO7uR+YR2+XD2
N8LC5teYJuUi/WqpUyt8CCJlMnwlq9XkQAgip/MgpCeA9tYKkskErAEZ0MuUa6kc
zDmGyGzR66+vj/tOh6w2F3BEQB3Mm2gaA/XemWLUSnBDCcUFyU9on2E3jVhVF7mx
hxmnLpVrITjGzSUIdQQ/RLQK/wEqGipSxFTdrJYauE+hm+Ltm0N8ZkAFrrtgbcWo
CIR+zGBVI6PASIq4SqOavAHBLmn4qXicAl4w99wtbd9TFqTA6n2g0qb8/rAlo3YT
GI+iD23mIgz1rxkTgJaA6JLrc70IvqQ8QcwnQMcvN2bp0vruOKq6UsIRHylGZkMc
WMJ0GBqbpgPWkGmup1HOk2GhZJr6v8s8bjhlXl7Z7sQ9xt17lwDDy9KfVaT+pdMO
WVcQFHszo+1hJrXQQzRWgxf6CNOwbf8qFmVQdFdAfmkoYAZieQZHoCx1pEP9sbLg
uoC/aTmk19z+K8zqQmDFUHdTrZRcm8KY3en5SnSMWMnl7OjAYcriIK7BCd+zfWC1
CZ3DnZoUhOrBbKF2NfOC9xY78QtpDC+nTF5kCs7qfKkElWKto1rF3AhMYywjUrU1
xpaUM06lQWzMSR1H0zoapUNEuSwLAhXQUW8iHC8pGLlZ9KnT7oUWqg7ZRe5UfK4M
cfVRbGzpihi4AimB2w/yYJDo1mzEXTYSDNpo51jGJjK30hKhRLtfD3AtrqXBzOmB
EPFA982JLF63f/H7NBvqG//T1yJtul7EXAWXqCQR31UFkvVRXMEBrnI2tkVdtmv+
vzbCEIZq/xap6APAavSWly6w91zZ3oF50k6zj6zKuZQI7jtnPzmXkq4ZoO9PQUuS
0wmQ+UK7lg/xz1VQJ+I3Wne9+ok4KM7cy955zNJUY4wdDbQ8JLiKkqrHYNIGZrtj
+1MqGbIEmdmHF3TNmmx11Lmpl3uphYX9kDswJpLzb6QFiRrqRaKHXvQhwyUCfZgm
pshqEOVZxz/n3Upsc1dUJDlFEW9yGbj4Rbw75c2isyWxLT7p9RkmhRymSt4ekml8
6GJaqJrLj2M8xz6sM5cWGEUpuanoSeLdTWR7C/K1BiG5D52lYCmsMxkpEvTuaw2L
v86cYxoeuEbf3SZb1Emzo5eq7e+9YnjVYlM18vI6FU53LhMBgimAbjc0oH/vg0WN
1I3TDXRUNGhlbH865yD5o6E9x5Mj6Zy70Ol/X3dOH3iacjBayT+ZMIBT5mJDVYlE
mS5IuU7gdNXCpCStSDCqR7gY6IBAxwKAWua6B2fvHmJlG3Hkug79arC2aqLViUpr
2PlDUPg09/glvUXyK7vv4NRW9uWp8Yt9Jjc8JLupdcPxwk+iH3vK3ikUuQkDGNyZ
1HtY0RYkgS68gpsOyFqulSmYhiA3XmLvJyGOM7NPnzegZFnB0pQiAeY4pDlFNk9S
tDhvZahsNB5VjRGLhE14r9C32E+yr8/yzpNRLBeh2jliYPMvDA74Iic+LLbtpsf2
k0tUnvOQ0juNnik1iYE+mX300CU1F5OaqIo220YTsTOVkPeyE4YwycKGWURbE3vg
4vYpE/tQRgg3tq0CFFulwU+J/yjlWsHzlVmYBNegF43bdrZo4v4O4tC5si95D3pE
VdatK6C9Bg2GYLFxTK6t2eNT4hu4VeD/pHDr4bXDUvjL2Sk8tECufv02F41xj2HG
UkcYNvhC1856smadNBGh87B2cfMGMZ3Zi7kPo0qh8R+WQkt1vU7HfBncozqkPf3v
CwwDk19hNp9BRcDQb40KWL7hEWVlvBiMwI13CM6GX+tVQJ91J86NQWh1jrZFj1TX
O2nSwAD6iLtL5IsiMfBGZrnleQqQB9/e5KUtAVnt5zCGOo99AXqSniQpPEM0IY8w
xholFgWhVs4wEPRdSDco7hY8l1HHTY1CIfIjpeopBT7hfzfFi0RoY7b/20MjE/Sx
UgVtQozgXKcnNZdud6XGjZj83JlaorZtcU4poAMTO0op4JNi6msxq6+TtEM6qukZ
elCatPAJgVA3xDMxbdBL/5awF+paDifFEU9v3cV2u03kGg/70CjyORml5AOfYjDP
ggVocbFq5pYG8Xz75A6HYbtiOy+vks1xSkRwoW8tY0vGFbu29vfVgMNbM9c/o/7U
LPY8t03MbY9jaPI5j8uiNZmA35LxxTNM75KftGmIYrSQDlfEsaBT0eE1o+Qqrd7g
9/WkvLO1J5EN9Mw5PsBuCzXGkk5/0ydSu+2zkj2Dp6yhtuEjuh+yJWMZKdAkKN5z
vJ+zEIU3SJxWmRhiq7PmViwtEiPoZuZdlhOtXBVP5+R29YIFQc6PaBQoRR2gV5sM
VKEZHTvO3INwT3sId6BLnSJTvd12Wu/tzCS9q75ETSIRZJgU+WlZdT8UG2lo+Oeh
7/yLaR2IBy8kg1K3Wm1Q+jg1FJvruBOctkum1bXeCHo+rJvx2H71fiUo1OHoIGsf
3NxYoE+AQkli3FH2FWxFqH2ssX/UiwOz+SZSRaMpPubxmxenmmbLK7lK2B8C0cdh
vmt0bHDw/rhLT4P/4NeVDFmV9zk+jM7GuXbjGBGlg0kgE4rwYZDbN5Vt3xpnl7pB
00v+7Pl4n0vYDbzvLbVwPvYNAJnLTBxd0CMajEbvO0P6MngIWa+H8qGZyhrGF+35
dH2qPGSkAnUL3r/X0xWyunASzwa8wiVoXdgfyHCYUfGvHQ/RBZwPktX60R8uN+FN
MJeXa3IgffqFKuTNDfwqDDIxpV3tB3zx+xbmzP7AkQUqv3He1DqNLeDB6JLn+DtO
bTYSZieM6gBtd7+uAZfMahoCqMZ1J1fEP8vr2wKAbVJEr+0IX/1bjhz7+bV0YqaZ
RCgO17cDqGlSyLy+Ubu7IxBm2w6H07lTcq9ma1DJ4XGouPIxTLaycvXL371X46lh
8YVP1fSHaCac5Khzu/VnCp2THG+19gzNqLm9bykPmCRXdx1NeJeGiCB8v0JDMLTA
MKMEZ5fdseRBwT5lU6Vqy6EFbKEQI1tn8u2jFnRLrFa3dZQyTqEndatJ3/qxGuAZ
jgSmfcHCuQFPKKiHeNqIyTI3kTVbFki8tiouyPcLk6iiLdWh6gDkrwwylpR2QqAX
FZULgv1HAnS0TwS2JCmleXDo6PQBvf0/QRxnambtvJVK0mSKbvDfT/jGvnXkBrDg
PGs2yt6r+r/mXAV7jNa3VzZa8zwxY/S0cfEDCOXWuPLH9W4xcmId0fhfCrtTRLEU
MRFpLF+6oL8hQSdyJC5dQ73yBaxpHhEUv6y8Lpf3O8GhgYPkdvnxcquDbdpSyzSN
/xEWyIkeA6II/3sy8yMRdRztD95K5raNyMWkzKjIre1Snm07EjfihkFrf/KCLukx
Kzm3cxkiURCSvVMKMqGBK5e3vM63h23UC6nPt7r57iRPYG108mU5OIA+sqQkj6uA
WWIfERzuIJ+a+BivLlnlTpBSssifPnfkRaMejc87VTkDLYDVVvwZBxr53JsCDoC2
UMGtMiQHJL6lA1ndw8qDyVUPrXIayxsG1GO6tOFO6wZaQxSIv5M0VayHYt4CAh6z
HlHkv9vJXbq2HHJSzlLBlf0ppHDoitFMCyXLIu0NtUg/PM9lcZj2JebfJLsmTV0p
35Ga8wbVRMNY3Pc6g6bk1khqiuxSVYTPeN9RuvdXCiibC3rVJ1h3Y+nuWX5FpGXK
+W8TbM+/GSR07KCE8og6fe+MEVoa0IKOFzQup1uHgWdJc5IG/8Yz8/cd+bbiey7D
UfGxrNO1a4nUvHrQGJwxylQ2AeFpYDpanNoSOZuNBG/tEOuG5Jgcc1tqhivg8U1Y
r8qkm9pUJp+uZcq8fUPvhF7V9UqVAdOoE3Z9dBvCln8sVQd3f9Bj7HJb6nABRsj6
C8+0Wnl2KF4mio5vgykSofdaZSzCU/MNlPdvohmnJyKRx+5WGA+RrlrpHF79Lc4H
Sg/zK/aOGLKknPM1WjZjAUpHVYjV6HTsuwbtnpiynyxCt7wv+3GWF96LyhmX3o2L
YboRbdHdkWNTQ8/0iPEY4otYO3WtykHwMuPWfF62ycGG9lKCn6w2X70F8kctEMDA
IjRIe1SFOHcdXGwIPu3IC6Kgh5XmwAODPOaXv1nD5aP995JCVKMqDI/0MGPNzYIm
21DxV1pRf84+f3Jb0Ia/Frhp0qBz0xQXueJFFjTkNW4O4JlhLdBfHOBTAuV6cQBc
NybKMJXrISKgYY3XP3ab5b/m33Q7zafeB2btilnrmsW7d2pdszgTEFWOlBO0MWFe
sbVMS8YSH9uARQd4U0phP3s6YDcoGYSa9BkwMhqFY0DKyRAR8MXlkQEbePLKLXik
E7/bG3qmvlEmrI+sE9XbmHCHZg9v4b642udeSMzuTCcLcizZdId143CE5uzUpiwt
2iAL45IHTPmz909dqOnnvkmh1ePhM5AgmcEILaYPScQ3w4G4zk5gb4gd8WuawU3C
F6YxfeffRiN3aZevVTZEKffQ4s/OiJLXm6G/1pI5Q678PzVNvaii9R4uO04QeLQn
nKMoAC+RF+3VwtDGYQFZgrhqQ8xeM9crFPI98kbxNBsIMAee/YDHttfXmf4rkp0o
Wq3mqwyh6ebLs5vHYzyLyw8pmxCYWx0A3CkET6xTFsJVYQbTLQv6+JYYvqMIUKVr
IQHZurKHnK9YazEkTsI4Z8VOmOEHhI1doi/RYsm53mFofnMSbKKNp561LOQ+6O+B
IDyQ+THt6h/a+XuQNxssGU7Woed/jOeT5ptVQLKWr3MncMGH3Irsd4ISLmiM11mr
IlIBHE4gl0jDMg2segXCbWcURbTnlYGooUzNwKA37LR7tB4LnAYcbSnYBLiipYJ6
0xq7GliNddTr401iPlIlOp7WCEDZK4h2iakAxNrICJ6Cd8/q+g/xrv46CwhL3MpW
mDR/W6pICHfAronZmdbz8D1zfBbA0laJPr1Pcb2/V6QorNPSh1mB+g/5b9sMKcHP
fhuguGRX9yuzIpdaUvWqZ2VtO09jMpKy/4uQw2XdR0yyC0hUQKPbKnnGT5ypLCNx
buuXAaNcukAcgrQruTzX4zFyitQFwmtbLzdjS2g/9n+wNyARdNo2vknJXuyAqCsF
JxC8NsFGxYmThQEyjj/eikygmlrZSeFUtWPDMI9Wu0vbWKi/GtmMInb9Ivg80YpW
MNQFiBHlTgIE0IE2r6i9zCvIw7j0hReJL+glHsFs/T6GLqDP2p7pC8y6XuXbyJu+
z3p6Ucy9I9bX99bDv9YpBhsox2P6CSzIcr6plfq2tC/AbEMHpNCvQaSkcVjcZBMp
03pmbHN4H3c6iSjcBwiDh7bK+jYJjwwpH4EzzpFwTUq8OO/I6u2XerQoxQjf/+XG
g32GJtRwqOZ++nJWWVzyb6D8GG2ZKUFN8cO6gXP0mnuBHcNCs5A/262fFqsNxvVS
6euhCPrGT+opoiFk8I3viObq+ff9RMwCfrBl9Y44TQZaGnBwlaNMwhIvnNtaOVYK
ts7jCoZbQjGLM+FGxk6EkfeIdn75nSIjz5RcNxzznzZ24u2ghqIaVAvgQIY5kLBN
PCXBL8rHlHZ7y0o20hnb6tOxJgGpCvcTJHPQJeJAq+T2eZ82Lv4Xe03FQQ0xvIax
wM93SU3Mg0uhOHfkt0GyMlDzPEipU3jQ/v6RWNvVDzlfJYBVI8cFmI/3tjdxj9YP
j0Tjve6khDzbjMcpEn3pJwK8ltYsfInKMPzDDKyaiCa8qs0Cc8cQfdHvjL4pJYn3
7R46h31zECRHjCGx8PeCW0f14aGEfK6LibV/KnqLGsnGrBLRC+iF+Y92rMWYB6DA
apuiF/dSpDGT2hGBp6j4voU6ndIqrIDYDbFQwBGf1sgdB1+4OUlK9zptnDZDHPEA
p7aj18ldoTxK2NtOKFgKMF7g4jLYSm02vmYyx5wBaXNwY1Ia9v9+3L321NLgSue8
A6xNrhIVBIIcIeptOQCwqPrO7adD3cl74WbJfWPMsrlGXORhBz9Qqp7gsWKvQNAg
eOSosYdpxnFj0BhjnrWBlC6zf53hn/gDoZVyNoS0uIVMGFB5Rn0uuy65UP7N148U
VRC3/OFfugLIgP4ukZq9yOwAvPBuGR5E349XVOvSgs6wLILFz/zq5zaVzOCe7+ih
XRBgWCpdrWg2ALQvBomOLj54q9LOunN397Ikegc9T9Ky+RgKt+1ab5lk4Sc4gvtP
B63215ko79frB+MkcLIjH0KAHzv1FGzmQYqoRo1Jt4hTkXGch8+QGrlBK0dCwEr3
1txjgXacc0IAE/BcR1Z12emL9SzkZyTD3r+mdENJkWMW6hJNBdXFC62C/3oN6t3x
lfboaUWU1veMbbNUjdB0pjPoYj13fNzgjk27d3usZ7DWv64NzamLEOOTZIm1qNLd
2UPlrh8DeaT2Rocb9UjiIV+uHaicGqNDh297zxNf9MvLo1mH6lcIgpuNfxNUZrCO
qiL4F/3UQN1D87pQCS//G1YjsgBEvZ0Pfp9lMJMT9/KVCtv6UPrRsjDtUqm0yYHL
mLyqtI06/Ctt029cF4ccNl+e7rKQkSztTHAL4a2HadkEOvkUrhdBSuPmXGDhs9NC
LxVmHYQTmM4KApRoQVdPBdIIs78RodyNzVVmXn78rs4Dtr7yzWw3J9au8shAln+/
8jZPW11vBF/txdq4bo9Eu+0m33KJAWmP4ROtBuKwXKzhUshY6k/T1+shZf+F61Gj
RAkohLuEhmTND/V4mC5Y5DtXMimcnuF1aWQY8vneSMiL6b4SsGHosZhw0A0QjEqc
KghtNQniEOFFVlOvUH1b7gDdnpZk/FYHUpyV0/ja/LZYUZf75d8Lls0/oPT+7hhu
AHITwYu1uB82lsIMFtObPTtuGJF7ssMjND09nspDAOdhfhC+ILrj4AS7ssHGAFbJ
rSnQchusGXDYU51s8sUsdl8MHHSkVpK4z+zoP3t0GMjrVDDW2kxgU4QC54nEVeSE
MKtR2F2QWyoG0aQuHHFyOKE8Aq7Pv/hGY+Dt3/unNXi9HBrf9KHs7Se3taZ7xMYr
YuwpYTSb6oPjD33YRU2eLpXdmsNyFSS1vuntVgl4aUB7QCYslWUiZOi8BaHajK4s
s9UQgoEyW+b/qUZoGR0Zb0KRNWAkQN8q9vZnfy/mVyWsFTtrScz4iPpK8fMWPClx
XQqGo3H21HSTrt19StyPsznAAe9P62tmaczd1vo5y0vtqdC0+aulAU0NBhAbHr/Z
QcUdifKTc1rvWt0QuOB7eTvRR0zNh5iMwgjmKzvbvi/ygccndfy0EPaxZrb3H1SH
QwSOC64YThy/ljxF3XqHVofeqFzCN+LO3yP05zc/xkQ3Z0KzzvfNydm9xbzlf81Y
rxYxSGR55HAmztDjK6vOCvvbasOZwvX69FdyDRzzaw9pS58cfOuhf0gx9YvSaWPj
PkFnirRcK6CzX3uKQ6ERzOCWsySclKL5iqTrFVl2vSCN1/mhtUg6GtYqDdp9gw0P
jMlqFdDrVHlSqtGB4nQJBNaAty7YsfnFfUNy34HH+k7hY3uVTeAqQog0nV9+ttPb
WyKvTIqlsM9jVmwzyp2K3oOlm1rQvQbuMPCVaGvNWponu+zj7tMBNRv+csaCuCJa
js6yt40L32VcJ4jhcQKvzvaWN1Iek+Mw14jRQ3Tu7d4D0Ab7cCRAthGU9DNdP/Rs
AG//YJOOgPoA5bAWoRubt7f39DUngkD6Nlu68dIKoW/SukSI77YgXproltAQ4uM/
SjxPoNzEm9QKjePtj8v5uVu/K9kEY2Snts9wnTntsfaq2V89bxZiwSt8LkFsTGma
aBWLnXeeH9fa6E76hkDvIGyl5+IxIHVD0pf9v3XszbUT+7z6kDws+fCevbWFL04e
juskZ8JsOn7jnI3rf1vmxZz0U07smv3jxSKAKVaYnWmDfz6Jb7wfkYQ7A1/WSiBf
jkE4U+IFrqLwuDPJv0SUn+/cq5P3KIAhbACEIvdQG8rm6SFzVqotItmgzfi2c7Dp
dqCiXVbgtgqXBHVPluUdv0sUNsBFh7Eq/S+mKaGQ7y9SQumcEdB6sjhRK9WDZ7C9
fwBfwHvzVZLVFU+FGQBpx/JuYUfOwQd6WUstzWGEMALFzfu85T87TlrozKiBfznz
f9AOMky88la+589WIFIyp3dbAYHOk7CZSP6PsoH4um4tPc4RC0iJj+BMUfqRiCN2
KiEIr4Dc6jLLk7CcZyX/jHYkMWqUb8wiTnE5HY0q1HOP0qY3a4v64Hme21TAFreN
YfOhUMmr5we6oo8k3YgDQ9pXj+90fo2dbmQml9qhpe47/KmXHU1tln65hBqTUVQP
GmcijJlZ1HzFBlmh2n2KZXyoMzpoPDG0whJhi0MlKudbSo9Y9wu1R9rurY23LxcF
Fh1tQZFE30CU34/tpuQoMenC58BfdN4oAAeDvcKd5Biqu70o4YD9YTmchB7Eb4pl
yLvSal2Gk09W+LhEJDtJcUFQ/8cXbWq43Bx1fEVnx8yAVzQMk8WC508Ds3cYfEKs
wQSCuvNfyWhGNGcSajwb3yC9XLZtMq6+qbIZCcIIxM46+dmaiuwvKF7yPlndtn5w
03n8w5J5EqSexZ+Dfsb2HTK0k6nOlstwdN1733sylYWTQn6vxOz2+F8/GhP4c5S9
2buhZ/M0TRF4oleUbq+wwmjhmnlE3SOz4e71I6lWawGnNr0Xh/SuzciaOVAYtPfA
JcFzYEf12aYRfWGgnCU0UdYCCKkmAkNPL1WIdPpRo7GodD4mlfBqIpGNB03f6YDP
oRIfq6594lUUoe4zNRJ5wYexC98f4nZUoVmzp5k6Us3K30nmBzLwn6RBSNCpTtL8
He15v66HFbPdnkiJP9yg1Bv6VWEeJsp4aRANmCh0cCID1TTIzqpjFHi1QSgGSo6r
TGNwSEGIMLI27O6Fyc3r+8suLkYhioIMZ6baGQuy3uM+aQQxlgZx6y5lyjIG7PNo
iiim3tmBiwjo/okm9XKk5IxVzLAlau7Tkw4zTDQrh4opH4AliFCEdyD45CVUn1cr
Ak4WtCqJ+9jubB1X3Kmog9Gb/zC8v+4EH0N0X9rgQ9gwi6GIhtFVUqlvL860A4uy
zK8veVoXuQDn57dP0vTyDXOKTQAw27tBKHBo/XmuUhzH859Oqk5d7DMfTAONk8df
tgUpwKIe8Z8JnYwOBYNhexF68S8uAhnJ2ftoPooGRh/BHS8UxK2E/+wkjX6RvMrs
n4RxRucGvmOkaHblTeugGGba3Dh1zlGZ7fbZ86wl2oh9MDNcAyz+SnaCppl1OJGb
QXN/AXohhq+N7M1pock6ELViL/3Vrj9Z8u3VOBTE3Bo+lxlJKHs6iPGUfdIy061i
1jx5xYTV1uv7qWDS8+a0WxMfk9zM7MjLoBMU9JSHuZZsiShSVVCZNVyP3HEoWb02
dZ1xUnBxi1gA0oq6HlNozYCFtIh7FrJnXOX0WolfZlYsXJrHBlvhgJGkty3N71hU
8AMbiAJUf80nFxD9F1P6asVCDGGblsc0P+CQuROIaHY/23lwIfEc7uYvgXJsHq3D
tPMto6Ts04AHraRIAGRGXD1VHPZgdQ/HhaVc0eObHSCjE6xnINFFaaaTiDVt191d
QnDjuubX2stP7AosrVtKPHh/ahr1xf3F/zbPe5SdsORI2v/2AtSvgQIRgERQNuuG
tCxok9h40dZMAFIZseQU4W1teoiSXP5/4ZKsIDxIjkc3t25mUrhaM/e2KJDY+AWG
KFz0eBR939BEgCyLGI7qeZy72SLFj0jBDgtXuKIUf68LA+M/sZHD6FeM6P9tsd6Q
/wX+liK4wXv8Fc9D7ND6mcz/irW3KEzd6P3UI9S8ThdNFrYbaiqSiKLLBduQJSYF
AS2yr6g3Jia3EuZi/d7o0hR7K7d6bsoM0DexZuKfVRVlSG2eCCe8Q49vsUZPI7AC
7Bg0OnbkZQjugEqBQ9JCwWe+bNIYoNb4d6TisKv2RtIXLXg54kXu5R+ds1+KSSEr
w226mSadFjYxcGYnt6NrMi2eXeJ5C3FSA3vG/iXlcQ5aGXGCCHZ6XTkfEFpZK5Z5
gWWj2lFxxm/NTi29MyAbo3Jq+UecdIgmTX33jm3Zy5lHJkXUbPt+b9pOKK5MZ/Ia
rnIUzCKEu2uXC4293UBX6f5jSzAtdP89RuN5RfqlM7EANHvn9HrneI2I0iWO0yf1
rC3nCMwQFfhXl/fvB1SXCaPSTpnH8YqSa0Pbn6N1h+G9Z18inlcuS0GmYAsWcTQ4
qdYpY1otfC6ouq32Ia8Cnc85XWUjG2B3sqnWeEb0i1YnxtPRWCrnanHJrSXj+20w
H0/GyR1+3sjTVeFgMUaJ2FRN9Uvg8/M3cg0HVw0QmAlYGb09qtdgsZjdwjlA1Wxw
jX++2hVMkdnMI56+/Dt1EYN4fBD/Y/Sre3aopliWeH1NnS4R35H4tOSwWn2QC/H+
AgsyiOnJFoKBK/rZWY/c+biLkFi82TDE3qGV4ASzcWTF+O4QzDNitE+HdjeZnzgf
plmzKrspf4enDlHnuc1qx9rGCegmujK/1eJJbf76Ri02itL13whBsydQ9oZE++Cu
vYT67sVw6OkTmxtydX967NQTPLLEZSPpd95VoTCAQfnTQzDlEmQO5PqAP9V4HBZ9
wnKiGNFPcH+ynSVmDwFO7RDX/VMWQOHOusUiRdJk33/3hs71rZcDQUWTMB8e/mhn
JjBB40d8BV+2KxrE0awB76DQAuWt4UdCj4v4D9xuk4+1tTwLsCqrtbBg7BWozGwj
x9DLDMKPGkwrAyoLUBWhJMnZRVwmvbakVQN2v8jGamFKnSz2kRix37Z+Vub1AAur
6peXOE3Cjc1BXIMeOKNhwMgQ1RJpDC2bHhGV45BlXSOhdExZM93ITPF7Kk6KU2wH
TbGHlOdkXKmPnPUBYlvF7ovuDZdeswx9Ne1f5oB0JMv4VDhU5rRQSagN3iHpRgEN
IRqwIKc0ad31ra9bQcp7UNnh6COzGciH0k23grd6RglKJ4zkMhoqpOsZhCA+febS
sKu7eKQI5Sn3W7hFzgwSc9Bqlp/T7uWGdVdJisEujVLwSfvOqht/NhZrnPIZ5eFC
maDd+zKaglyVCcpUhTgHq9U8aMu3WfsQEIhKQ0qYTBhoj/i15g+0FTOjZpqkeCEO
s1/zhx0nncrm8FM3CN4aN2GOL2DHFUZ7VJPqRLstmvm2uiuzQrJBv+CyayCFVaI2
c08UrWt7QfN7HFuCtvjG+1Fay+QcnpPxfkn8Q/1ZHZVd/Yem7lp1GQKx2lpmAGP4
2Rq0gZ4pMmvIVN0sJoO7wgDuc6Mdv2T+89ZmX7FlIDIRcvoA6AENStAvZM4an7SM
jP8u3tKMkTTfN5tTHJztXWcICkFjfDx63OpO71ehfJlCFqZgCWWvTQJqRO2kUnwW
IqBYvhbavvV/Ork7k14aOLQVHM44lBTc8ZOfd4PMz1zoqqBSuV/VSdgkn/Eoq8Oh
m2d4vw5+XPJ1mOGccQENl0wYSIu/ilKs4j0gvKpqw2coXPZVAYiByuRcAP5v/itd
5HDv+zLxt1oiL2Lp3klshVWUUJwIJ6CxhgsejLLgVX9lvWR5vAl5dMnpzkCi8W5J
VbC4bXsb3yMmT8f/HI4a2eTrHZMU5vPdu/Wx9pUIWiYhm/47jUC5gQ/AvBwaMdOd
wzOYrFYoqReCemF3iUcXHqBZQlB4h7K3dNQCsLQBvyNKEFScxCWePCEyCqcDdJ3b
UbXkvy8Q6B2B6NJttUMnzy1lFzwSJ01tD5+fowXGQLOiFuXjRcA6hKg5NHp4BeMS
EzIiKnatB9hJiQgexzd094TGUc8uN0gMvZWcG+9RsRwuGuUooY7/UjKgTEDmQIiW
O8QaAF7PzgMADS2LUl2Id23ANCcDoj5iQiwLaKvBpvPDdtsWeZ837Vg1K75nrGxs
TMA+A/riMfGtv4vk1qwe96FB4xdRGF/17JnjpNr/EpgHbT1P0cl9QYM5IW2kV+61
mZmgu4wMFy/aIjEzQWRGyI24vJSwkrTSqeM6RMlFWgosJ0O0ISxWiLtyBo46H2WC
vro1qbGxW+b6cdResZAkip3r1QmohXUIV7WoxyMoS5vj4ZOnO+vNqI5BdJAD2ARc
qIvD3QGI/7PwWnOL+c395hTooC8+SXFTgyC5xFef7dU1+NOKQKUVivqvVpGSuFQO
IGPjG9aV5u3lsla2MZT4cZrvrAPyVECITcLP3AeFMlLHFz39zQnNp7gg+LkTgttO
GUiuRoQ53EdjkBOgJGu3b+ahrpqOl4N6UPuPFBHKMVnNMJyhH6Kgv3bK7imZcHXy
O2T4VTr0Z5hWTAAUwAoRJVqHHETKATYFch3a3Nw9UirruDBSbCIrNzo3CRX3c88K
POw1JDewzpuRjPtU3ywr6WjMw5Nkmxw2pGY+HKsHV9F3bHJn6XgdoWVI7q3lwd37
xK0UBkZWSqKiUebCf5zpMRQD1g4Yj2k5D5ePrPGFA4TJcukJLSSi1QTiIIDbF2Pm
3oWY91WD7jtt/JPVoutqzAwG95FdmVJQJ910z4E/+omFlRPTPEIZqeKU+sscurB3
vL6HvCnWJlsuXXut+OyyCTgaLYGG6QZ6oMH0NVEPOYxPvSfG6BWd3Wk4HJsRHa06
v+yWqHuYgrZHNK4hSM6mlCyQOWlCgUlL6Vot9+LOl2bH/wPTlHMP4sBljjAZIpHl
AO6gSDfuShzCdgZPaMMOHDuIcj0oZx3N5hzYzUBVnPSYujmaE5CxVJcnZo6zbpc+
biLbbtA6HC0CDSp53yawYnExFyQj75pUr4fVjDDLJcVLNtpqHiYIvwCu3Q28Anbn
YkSZgy7gbrAfERNiNSHVKBo/pZCnOfbwjZytiOUcNWmxwg6FWOXB8VFw2ouJat3m
YLoeSldmh5UteDt3odK+/SSsuLJHk89lvrh2FzJ20us85G2z9ee4AIDO5u89C2UN
l9pVfBasTt2J4Vxb7/KFwU/4OvbCCf1DHYaOYwZOgowTN6Gf3ye0jI66bMVJDRjz
XQ3TpMuWzg9lYsK/qRN4AN3gMhhzfPgvsJus4QwFjAOazEkhPvwAYqiWIu/creUv
Q0UjAKpNXEi2yDT5euFUlQaC/syzerR7EcLKB206xy2nWLQc4uMcqctadGnGcCgo
AmQ1BYnIQM7X4hb1ErFS3fy3bgtOXJFUOftciOh316vlcep0YAl+q4ULiKgKdXdx
BZ/3vcmnAWbb7QxXw+Nx3EK2y85t9gJG1doKEh3TJwb5Lh+ON6OE7AskU55ZbOi1
Zhj1YgD/q42g3LZYjqUprgPbD3TxqUauC99OPd/yjL/kiaJ0PhLNY3pJX/8olVlH
naU5mVBZ09QYtaxyBbcER74XqRIPnxPleZNwcpDLgNa/7Kj+KVCPQXQXza+9Rm/2
DBUBSETIIONPHwJXhonFePAMh4YWpiYjzTFL9n2pqXzyT5LhQTKMGw8v+gAaVNPe
HwL7WYetnLUBX+P6tY55J0SD58FB2Wdxq3N1tOFAk2xjF5ZcmS96p5VnV7uVHC6C
K5zpUYKdZdeWykBjSTjd4J5qD+aD46c7sAGlR9JC/byEzdQdb1O0ZO1Grku+Jj9H
3cRjLdLhlWeixXY+Ria9Cbo34YEEGxi7BGncSl8Fxxpzbx21dkYYb6isID1fQZzc
QknplQAchraIgW+L1sJWY5nOKmh70KNcIH0mZAK83Hn7SYr2imvr+HnJY4UI7JNB
poe0QPr79DGnrJwYZyRJbIZ/z63x3tfTl5r/DQbpfRlkvGrMczGKSOaLquWyfMgZ
XX1ttWxYfuGia1dwiHe6fIqlw2rGCsSGRRkjM3t0UuECMcYnogqUMqTWDXnNbMyX
vtNrgXyGe6fycQTVWd+EEAdOAyA3tYrXt4a+qZw9pUa66hYIxcTmZDeVcWYmuIe4
wMhkqS8taxoMvTKaHlSHbVz+c9pzYppUcOU51tF/7jQlj+sPQArSkkoR2x+COKig
JzUSqnugZSTwPUFlfq+sxFDM/RqPdyXlhh5vwmqN7W9CenO3MNt9P874sHThPppv
H7ZseOjdGgP3C1Q8XBhKhmzWw+PVjiPqwmtU2V4DFFGt7BkbHbpk9TTVGM/uc2p9
Kv9vFc5VlA5tQfYAmcCrp3raY7etmqft1wXz02TBGp95uSlLuBNxsHJcFiQ9kudR
RrtMs10IpGz8cFqlgMyA0oybcY3gpoVpuHxT4GAu9IoQiVTbHMwiekciocUfjW6Y
qlOyl4avb+fwxlu8xcbR9S55gqu1YDrF6rv/P5ywuZv8A7/BcTgBPFxf9Zw9FcPX
CSXRhmHkOmEmFMhmcIJ6dEvC3YfIaB8QZju5114OSf3iPLuDqHQlgkAkNsXM/d/Y
OrNjC8Lbqqea+27L1h5NhXlpL8v9eSY4pBGqDS/e9NJgkGxIOa8ubFjwq0oekS6U
ib1waJa/vlu0BATRrUeGTaDhkze5cAc6rH5Nj5+e3F8eIOOSkgxEyWlHrWW+EnuT
4NZfFjW7Jov3pK1NEp1HK9lAnBkZXf5BfBmYDHT4OwSP+jom9FSyYcvAxk6M8G6e
BC9fF9OC3v48mqJSQyrLH1sEu3P7Q74T4UzI6MvOyY1IembrAUejCy2661UzFA52
x75vs/oQdxgVLKiGzQDOcsM+bguFNleQCXXIBp12rua1+2uv0biIqRF1JvL7wZgN
2zB20rKob/ovDEewGlrMFm0zjX9FAs4NvbZVHhTkL6GzBL8Vm+4Tt/riRrgFzgMB
7gzYjXCCgOrJSQvLB/JusE38Yc+otwWtaUa1+Go1HuhtqVsFBoOVXdWERQLvLJ4r
DZWK69STQfTRJGWlaedW3cDHvkkV5r900xSFDUzfkMivHC69nLEdwZDp3t91/Ng7
1AqlzKinwno3MjSCxxBzLrv1bxoAH/3hkCWuzbdntFTDPmWq6zj5unpgqw9prHQJ
TG+KhYc5qhPqLaQeZi+/tLQPc3JhzCiTzcSyTu5dt8y1AMy6P2H79xQfwWxu+cXM
xWv8EtpPL6zdkIrRBjz+5PPMkJiuVy+t/Yjs7yWm5KfSn7s6iMbWn5jqVU0vuDYJ
oB8Ha/CYLjNOkL3X7SvUsVz4myEYKibQQvEvZYNABSXL9L+ZXY5CsdqV4C4Jau4Y
Kg/wAvhpjdfnB7a5Kl5wQwiQ3NYPqPpdcn4aBYdbqFWVlvNhvBGhQMlmZ18nuLGx
mnWa4RFE3fLsSLvdwfsB49f3hZhRLHvSzLSD/2MN8F6mFPEIOptG/RRpgtoxpaqi
StS/WpLOlsEiKS4aoAvJNTI6adk4DpdrQENlWNfhMp3BjksiolVQQ8BgxfbRQF7z
/vVjp3/m/8TnHo006vWQnGdRT/0xwrEvVWr6u8u1vU/Z0MW2f1z++7JUwo0c8Hzt
4s7gwcFCubpVq0HR94yerstaywLDLxofADGW3qNKw47TJSHRclGGvnczweQsCkoK
2WHx6Vynn9NGiqt0l8zOh000t5ay2XPdl5Y6St/56x+iD0ecyWf+F8/55R3XFiVr
dQsYGKF0w4zg7qQeY18pzBUUsH9e9i6ZkUxS/q0KCnwtyaoXYlK0p9L13+4g3Fq+
14nz4vjTEmF5RlJgrlz/nB977oxZhn0r1NRDFUGXjW29YW+75HOCHO/1fEMRUeN7
q80eLY7103bddZCZ4Js93Ke5zjPIK58Pn5uldfcmbAdMGxnjnH8SdIwjwzgjpLZO
8yPeIeuehY5FzLt52HdirWhSAe+KhyLOpwUaVzqcoStK19UqSCnRo2l9ZZYHtbVk
Q7S1AlLGlFesqmXs+x5L2JpFmPN0JFo+gDELT0dJpISoI1D8PBsXBl8sJtNvzUBi
V47PG306GKtECLpNmvotSp3S9AHe+nNZGADr/ctsy8ZUJbbmtGERNO7YbEkJHdlU
o+MJ7BOxeSJR7iBIAap4t2toIsQwtcSfhvC3V1p4Gu7N6zqGe5x3iq9/SLeo1hjW
cOS3uAK2UCxU3+47EHzQmDrsX8r7GBkaOetsQReGdk2lo+m2ydMD6+Cartis9vNg
4fNP8D9zuyZGznqjhM7k6Dkd46y2yjkHLUKdbQ28SZXP0GSKIOvBbz7eaZVhcYO8
Mc+xA5RihnhJdMeKRRQoJ2PmEzuvDXDrRg1ahFOYp5oAsfOy++waWv+K/XrRSVis
XjhRbQ/eN1hLXqgSDt2vKQe5ArhBx3xQYoii3eJKiKgLvR20QEghSf4+YTPdxN4O
GVXawDbTYbIEEkvd0oiItPeJwtg4wTaDkMs75YtQMow8vLTaKizKMrzTKv5gRebq
+Dr8aRWf9wmB5MNEczwda9q3tARt/akMM9mTxKlU+46uF5I6cCaJGB7958hE7hH+
+tMzsvDJa3oH53rgQ0/opt5+mzjHvxO/QWbrlG1MFN6saHTYHoCTv0H0ktA0Tf0o
e0V2qOw2RbC6Ly/A9JH39SQJv+EAUJ96j9IXjjkWwnR5v066Eu6WDYW26G2XWYaT
1gQwAoOoJ63X6CiH/7Hf8AaUfkPsRYWLdZ4zPVc3EpO8nLARlTa+SZywNimZCjxr
qLaJyNvHA5IC+g1QV77LfxhgIJJsRHYTrpUqghMNYPFGyHwR0Rrv9jhIcTcWwr/e
GRxeTFjZ2HmzEb5KxdY9QSnVH+i24Ywbvc1pfayyzZ56Nq9WaNAOVSNdUnpvNFdh
74C64SZbLmpSqsjloXsEg7e8CROQ5vhaGY7YcSg75Y+qIE4QIQbhWmF9n/y6b/Mc
vXWR9FH5TuLqfuoB/1xrgxYXaZ7eQ/mzCaRjrq7ZA5YWyvl+g8QFzuT8drIZqOj2
E6Lq0VMBPl2DJeD3lKmm3ICH23EKxkCp458KKVPimfewgb7GaA2rv9rfA7ADT3ju
a8DV5cx3W1CpBwPe5lMNNZdigDcov6BfQVgZoQ92zAGXgMFjxywl6Netx76sy7VB
Ts3w+ZgCZeruJpS/4U80jN7hztDK1SR6XFZSXnZY8mywxm0jDujK4CTsb1GYb4qV
beu9uNJVJL/LFI66UNonU1S1PDu7eHWLFciH6TqTwgA46zLopILKsvZsDOxgklu5
xhRoNIhcwF4H21rJQosGe4dSZfcZBE92XuQ8nVE5l5IEDzS9JlchEWm2JEjzGmRt
3rKvwx7hZrVcphcKji+0tYf7cPPKoyd/BtIzhWsL+WFwXOi0+nzMEa3u0+Jm6Sv9
t8E2eSMC54cHV5ozLnIcOuRlELzOQ+B6zk2OL+UDd+V1Ej0nJhCucL3nDob5Ld/3
QCrPO3iPxp2cpxnTKujgwH/+QcaAe1uNmmiNchr9CeDq0Kd5npVD+eR0yltn2VnF
QFCjLcKvMDDPi62iHuGt+k0a6zYxbheYRyfoJJK+Yokp0Zm0yp+KG6o20Db61tjs
6FatqbA9CLMx0qmuRTHrGkS16Rg6z4xyiLlTC0HFSn1mhzeMigsBBa42R+tFx8Ld
pTtHtrgF0xMv7eOPFEWrhD6ScjNxn8j7wnb9CYBtNL0PS7SbxzSQufZ0YihZloCp
bzpIjnN6yXBmbiWJsiUT8pv65V6UeSSr8okn5Ys6R6CKZNmC/OU2S06Taary7UrQ
c85+xAcHt829k82Ohm2OZA3t3RbYYjaUOyWymoi/T56YaA12+qMr2ZK5RMuiIDfP
kOvBJGP9tLDY7UuN2eGuGXgYFTQe9GFY9jgUe/x54NVAhe7ZcXatbEPAtift99HI
CtHJBIxunCdSoUereV2uhqKiaEE6L4a5/a6b7kFLB4OvOgzuslf+h2sBo1flbRmq
Ll38FNWT4Gz31ZIXXO4Xr3xWeOlJEgU4AjBjAMuVl/mZBSt/lSrwZmphOL/Q4C2W
VUUVdUGdT8mENYGbJb3gilD2eX6T/9I4noCp3JbkLLnglIFAHJ2iCO3vEciqlwtB
2uVK6BiPnPrNHtnjx9DLkZWMGLyquK8SHJ+yFnPd2sjzGLgDgyvcvyJW2fma4B3r
ypK1rcScRX0jS7ww4/o54kboz0CzV1VyogMCc6RldAjaF1x3bovN2j5CKtjkren1
IvIUiTta9Cs1bIUfFaZcPUQyOew4Ukto8WSlF3OinfDeWZNlITb56KI1ykmQPhU2
BjaGYkkOfIygIMU8DQABbd2O1tnzmCjMKa521kv2DsizUELi5n7HV4+d7dnEF7BS
MkUfL+6PCYvjK2V+vi+nOD72B8gFNoDClUSadwPkrDFbaMXjtMryJUkZ8rdOID0h
Bt2V9tRJEwr+DK8DSVis7fsE0TF78HUangOni+6V3dbcZaxryT5T62xqDJp4V8+a
8FIPzHM3z55HTfBB/p/Rxb35kmSg0TVQGDbiL8hLZTL1Igl3WltpEx1IjRcvxenX
mgy11F3c5i3Om5gYsFvFkfSa0L+Wf6F4xC530KbCKwy6pcBro1evXYuFD2FiK3mT
nTQfGquHWY1T3KPZs7L597OjhfA/XyEA9s6ncYwfyT0LnE+XFiNkAdsTINmIMMME
O79/FvBFhz38xHuiR840gB8IqiNzLOoe+7mUXkeSnjKL8oaETTj9aVe4s1Ie8YSJ
r/jY1XXO+zC4fzeGcWiWIp0Dxw8i/O+/taNTd+IPrNkdqO6LGNg72SAUwiKVdanL
VRx6SlGf2ZzIXv+078H6+/FRPe7KjIcp2475L4RQvdED80SqdUokEoom042l4Ed+
FPpELZ9G2k1DiCaeollBiXJTcfY3vI+8+TQ5KDcYsrrrUpO/e3oDGMpO+jstaeyv
+ckdFrf6lQTXrZMjBeANYNU+njdzDpQmjxZkB69DaplgI8Jf7Yu4iUIqtATZNo2V
PLkZe9tcRdhG2KXmuVgTgZ/UWOE5YS7LdTgwwNpHIah5zgUcnY4QLpUdtPRY1q0Y
X/D9nRqYNDXpdf/SxdUpi6i0LuV6bW82wlTuYFRMsfO3luEUMXTbD0IBu1hPf30t
nnOV/K5jGSo/mGmse020ctSu4kOVYfWcRhTQE6pZdbGuJ9aP27TDB6n8W0JVH7n/
m5FLvKeXm6sSmTZzECxduM0DKIj24ou787m14+rTdJO+hC6cyVpD4+9auWTNAsUP
d9NMs8u8mRAt9XW5nDeheFfY9c8GSXzv/8U12z5BDtkK4OzGYr2/HAL6U+eMBgrj
nFqXtzfFuFcO7l/kuoLjD7CaNlf/s23fXBqtikZm8QDFPdq5gwkQnn0QYAExolLI
KXpni9TwN9SMaoaV1s+2yTPtvpVXJr+HQUGrZm+xXTnciLov/KGSlNGb9a36cMfz
3cinOE1VgqYLUPn7SarvZduTSMj/FDhAYEHg9G9i6S/b3pmYNxmJasg8Kx5AXUJQ
x02/w73UuqjQIMvguPlvgPlIHfkAh0frqO0y2RaPNdsZ0sHvfR5RBL44KRTP+pbv
9neFchG17GTAzVQnrQvWUUvm8didMEl6V2fTgs+Jmzuy1j808sAfmfMAhOYHRQ0B
FARaButTop+jRmbF2nU8ir3Pp8dQnbwH5BhGA5HnEGPlAHvI9S4M3uiE/wzBAI7L
Slx/mQpmtPfH6ikZL9CGxATD5Axb+xdGLJUZ5qbC8pLEZYq7aEPH0eoF0VI7kJ+1
VJAQXnPgEt6Q+IZ/l2aHHuPg/i4+xUhRQAVzmxeoRkMQzXNmILndaoiO1TB7brJJ
xW46oY/FCgyEuYtYOcoDmI/q7iPx+ZiLz8QU+rNPFTcZC5+1QL0PdB9Io7Xp5OiI
oP15YVat8gTTK+hDKwfg7BZa9hbVTK4VKkkr1mzSzYNXPUZ4xnLseBNt/si8tTfq
psk5L+wk45mzhbskUgQ7x2aNHkIElJrNH0yzreOM4NInLHekaCJmZ4JKGZYt7lru
LJtO6UIGfWYNiKHVKzBxkrWOFw4ifEyY6cPaG2OQQhbuuHanAEKUmjgMbMlt/FAL
EGHZqyKIqJMIigZYQnQuXYQg1dIbmuXqWMrcZO66rvo+RgAt10JrTj5UnbpBebri
IfG29AsZfI2DFoxBSQJo78MPBccsAembSydbTDWqcPGhYr1YGa/uAio8l2JyuuqZ
csYNNtAbxv9hcCLclmPoPlGaolS5m9MlE49HFVkbNz4NkuFJjzCD3hMbCV/frgoX
I2NGlTXOZzU5LteBaAa9mPAIe5WE/W9cnv0ECAmS5DmO6OANtmYvMDtUX2Q6cL2Q
vY4Q1oipc/+mkT23Z1Y+2mFGOOEeuJ5okQz9G1qbl6jWgw6VvRd24n4fvdkDXDA0
3gahAd3HV7C3k8bl+VbqPOfltDVcskIPPZcgwG3+LO87iSXq+bvf1Rsqv0IXYiyh
aCW+kJtu3x9XdKzslOeGDq+hHc+h5bROy9TDxT7uEMye3E0TV04HqaTKNju1y3Rt
OyHp2Pl9kgCvp22dP/dPJgLI4BpkObz3509f64OD8Y5yJSvIR/3D5jVZlwX1h98x
CiGyql+1z8K9Uhyol5+kWpzt1hLuBpallZf9H9MKj0i+wn5IbW9NTmWJXAuUjPYC
RvRp4RJMUcg884+k3dZ8hSFMxEQ37Ul5fGTI6Cz5crdawmHN7cg/idLporSkF5um
gH3jWffHHwXTAySln6C2VunCmkRaLJuDlGb7dycF43mERQJO2mAOP7ephQPoDJFB
Ed4to3bm2pJ4ab6N1QTDGu5+4xv0QQoDnfIgLCy2BVjX2HLa+y6Le+J6iuwYG7fH
4dLMSunOde2TezMUKIyV+B3o7rQRZGqUp+EOMOo7oQnqgCQpdBkkh/0snj05hwoX
YZaM4IYLHnaavpimw/JRWCQhPD6E6T8VFHn+ABy1UWtUnKsgtfIn+W2W0O0fr4FE
YNQwv/ZOpRiR6H5+N2PiXiEVMGSIUEAzwhQ6j7oFw8LlBRzEyzKBEKVGF61eB2RY
aXyd+g5H/C4KA+LJ6HJtCc8Fo5WavUubqpeNHiUQKYQimSvcUpWlwoRysqkTR/nh
7g+X2+xDpAKmwBFtcsKchT4xpbn5N4+uJFjuI78Nv34/jKclll4F0RMlKPFlkFYL
s1lL+DvrFio7FV6GoHYwOhdtF7BqFKFYGMtMnl4Too0TxcQVtSYm/+hYRLN26w7P
ZhF8zF//8XRLLOJ/5679Bj+jGgTzipFDUnxxcT3173+4zT9ZHb4/sGOCJ5mXhUOF
j1w99M7x2dJQ9ysVZtxisXHK627ltGtbE4IcXiqDlH17FIt7VwQmJQD4MiGTZvuW
dObww61k+MMHtzZxHSvK9EqEX2R45k6JkxRfpKLf68reMUDYHuPJDObZ+pKdtEo4
V3nu0rv/qcQbJRTMjvCAcLVini0zSIky1BoNCMMryc+PlhRVSJJV1gCcZh7KNbHN
C9i23hNWYU7YuFuzoX11mJ3+tAbpFrYS8w3xIBBkF8nvk/0hsNs17jus9NHYL8Xx
ZJmPGD7bz6optOBytxrUa5NL1FwW4MclWJit2hf+wyBdTHKhmjotn7lSIRpE8iWs
UiEi/va/vZwIT9yYnbcVLkJEhhvcnfXemGKDPMO3aZxjugk95B5k1COCP6AwomCL
Wz+ePV9cHkR7ewSUDg4ZR5cd8RlTlDyzKb5esKNIOnCvVH16VCD35ITBQ7oGWW0N
0mxHVRblvgcLIFAaA6nl5J2DONlDqQBDWgmxJ1afgOwwKNX58RBF+dZOGT+N39U/
YmRYLdpW1V4SyqPrLRuyCOr2P8kAMq5mkEccr5sBOsoItcZHkEoj0tE2Q7fE6Hcl
Ibone4SWZ3AwZwpD6FTJFHJTOXl84nfO+DU2vtGojkEphCrGchb2XCJ68uv513tD
cw9fjMfPA06c56YS9GkixaRwLrKTUMkuq1JPSUtQBCgFF0iM7GIEf/Ordh3D1zzG
h9vbN3eMmeDv3pb8SBomDJzz4NBP6qCXCNr5MkuX/BBdLdS6xVN+zxxF+XJcRLom
LrE7mFZbEzuCXwGOY7fZNXLBmG+4+64K/ekkh1INrElLPGZniFOARydl9P1Z2snT
BCm8HTo1srooZZP+6t/rrmqXs1CyYjBifRboDQ2XgK2elv6qY2gsyFbOmYtMOqMa
uhgBLuWONXjFKp8wTYOkhdTi4DR8ewlzRxkQtTL5X+Q4DWtzLyGF/7PuRqTDQ5wV
POpmNp/v4gAFSLZStN4RuE7tbMbEz0SyxqhMwq35WqWL1OwJWsVv0JUP2z2FjZCp
dlsg6GzAC59YCBfyTFHOdmVJyFgrv2wUvlMmY8JhBSdY557Pa4VxtSrFdNc+mpYL
FewdB07DywK/WLUT2euHXv7u85++FuJyHzKv+IZbhljLBy48npygsPJsoSjU17KW
GmBoA0FXZwQIClbDRU6ydtQ7Ft5HoqO1c9TOaYM1GvwRb/eii8hIwLB2u0NXp0xB
TqoKUNgFDmyTNhTqDzOYR74DN3v0t5sA0evVEX65AKGCLg6/mrX71i4dI4Xt+R2R
JA/vTCq7YYjGV+1LbOPs2bjK/dzf2PxoPGe6580SQQsViA/plcYpk/XOofEZ86xx
ULE4qJVhVBS+VYutmc/IezU/WsPPy9CdThBPxXOHDpPaHfbvl6QhdDfpBYuXqOh7
bJmBodzxOySl0pKoIza+vlgvyBgDT2nCtJsPjXu1kVo1I17vgEXPgYj4Hohl92VK
z8ImCjRfyq6lM1hCXzreLvTFSY0AEqVQtttj234goEEgNqcInNxdmlIZDQPS5blv
6bAVUXcpdow07xhz29aDYOIYSDeYucfYll6wLTwFYnIPeVzusqG/nGZuuGca8Yfg
Ne8Scx+HgzRUUQMjfapK2QDRRQOS6APtUjIl4wURaYdOntGPgXTNdGZyFUikKmUG
kTdKA956c14+M9VDuJ14HnkUByEyDz2qkKK/NYNHvET54UCo1pf1tDvwHpOHzLEE
+MzOvYPW8HJLEM04PnhcvNKZiKDes7ykqNG/nX/ERNm2cdALISiSFud9jZy+d4FH
UG/TeYlH2jyG2DHtAmofr1kqxGRie815n6/YNXVam6gCTPZlnSXrUE+2F+5UjmJK
VEmWvhHGn8ZABi8QwZOuD9GJkgt5LmP+pqEKxkdBxhLsUFIaSEk7199niFn/E71n
RRCYVzHJCTtOrW+2VHr5IXqnpfEuB3gsLxa6kcvcEg2XwetpjkGSpUto40S+lgJ2
3R8LFH6yXkEUfxjG1WRziKW3hrKv6R6rJ6nelnpTOlDfrsAXb5gLnkB7MDfBtb+K
m6CrItu3cf5yJEMpkwi5EZAIG0R8nKePuHA5QklDbAuudkVEYzbs9esdZmmAzTOy
6s5rxbf7kmo5JuzTAKUcZ8jvcCxFDwjWZ+3ntfpru64E3pPi2455aLDlMnuiryx1
H/+nrom1V0uiTAPl3nibl33cdWJFW9N5UJ2suFwz2ompWNF7Guu5EnRrWcDEGK+y
WoTmvQzia/wUWy9BDeg3W0mircWxODci/H0to8y+gD9QAxiTQbGcgJ5Z3gwCMXMn
1ivuY5LCIWhZPNI5hSC4EDD75idnSy2o61epNAE8nReblE6z9rt4EuR2Ma/9m9z+
tbU+48yRHsd2SVJKzIzdGQzMSEqhN1rLUsTqTb/Wb70oL/wHSHFd+t1n5yGeTg9L
bNeVPUSXSCYKVuqBPvu5gez40zekQ00r1MZugDSIlloJ52hwTDhGeTDo5XpsnaUy
NLsOevbqHZtgD3rj2PIziJQJ3W1WhZb2C4ykiuaxFXMqUI2iGO1ZOTup1LswDUFV
uWmF0urRLw9lkq5fDvT1qyTxvPeeV3/NqKRhYJM91lzTO3dMpZJIUya8ip6EUHZ7
BgSv+qN2q6zm+as+OoifmWACRLXXL2TjJDv8GkFHWXyA7ZWppzAx0W5vQ/D89R5p
BX9UDVPiNPTJKPZz/ATulomHBX9Vy2IhUovzbnDPXpacNaIcSKXgw92yCKblefpl
uW6vgnynVDRHjGc65RYWgJNXqgAqV86rSAuNCa5VVRl2IevNxfgjcC883vkuu4cH
kKEHlgJSLlSh3X2e+Ycf8dYjqI+ipYiOs53bnie5ExyOddx/1iGp5hHtHL0cK1L3
Z0CJ+a3osYUZo7EtHafAl42EYvkO5y5+ugfluNFgcUMz49mxW05hAJkHM4xp23Gy
oz4ikd3a77iC8jrB3gCPvQDxsPB7bBAL+gi/unVQbe4IBvOMPKr7OlKEgcRP7Unz
62QOYka5wRgfPKa3XeVNoD1qX2eErYP6NvB7tkrgu8QRl3Yo7tSsdmjHP+UHA34H
knyLlCxHyV+TUoIitEiPJXSBjZcRu4Tz3dOkKVWVTYP5ucxyrAokHtffzcszjSh9
DkRSTP8r5GQMLiEp5zOxqM+bPEDwcVxZ1VdpPvZtOaz92djRDjGIEwkaHiShs8ll
c7Zh0QQT4z121W2ngXpL/iWyb/xFWE7xg0jejA4rANtldRph/XqoqnhuCcjYrApB
mpH70y9Vjlcza6AWJW5yDUWDcjGsSpN238wyBNbwsNSqx+yEeWv/2Vdokv1EbkpF
MN4XIfIjN/hTMROGm/CpaOkVyP1V7aobaTNAplFrOGq/iM/vHI5Q/611EuzM9m79
8nTYbN0JCOXcvzoqLBhTatbPI6r2NYvQz+ZogkJP07l0uxOua36Wdr0qsIg/cFpf
gODA/x4X0rvBiYpFufkAxa2cd8ZfdO9106kbzh00qhAK3yKhpeJdzvTqQfTSYjo+
LKP3zJpwVSf1cxhaZOsWUjqJXRTfdR6ZwhduASpzODEk9DxRefS2pkO3cHkNHB9I
UVFXmWQwHckNAXVE5iC29ThmypxvQ0jdQM1S8ZjQJXDoP9N00SebqQ2AkshH5pTD
87DfCAJY9f3niw8Qd+9VFxNjG4xdd2xMnhiIG5BIBIyaTL8T+OmvdRFoZpzjEN4n
er0olNgSVAUDya1WurIQoUtN6hfLuJVy6Iz81EXfx7R0hHtT8WNTp+pSD/RJ1e3L
gdXgDb5P/5lKIQ17hfHjamQBEZQc2vgk7cBa3Dz8ZpUh02SAtkTqW+cNiajlD7d8
cL0dJzD7Z+sL3gbh794PJzKZjNPtwwDQ9UbQlO70VDXbGYGsXwesTmCelrm1WfMJ
/uQUbMovzJNcXhEwFHYpdcid6btgNSV3dFY03fNAHP2Z0tabdmWfgYvOAOcNskIi
VWM9uHgIoQ1q7+HOo9xdIpkZzOCOF0HhdjwaesgGoxwxWBlJmsK86JBCRHq1Kr7q
s3cmTdGbLZLKYXRtP/ooBB0IuWz9a4C39QBbN0LrNB6JnXvCCzyUd6bYWwI8o076
f0nntlpCvEQErjRfGqheHqXmY+hy05qsbx2X0BVOtYf1HI7e176AhDbNVINC4YAn
BFjQXYEoqy7M8FEdJqqBqPoDNPJuG4uIWcjXbYtYpbKmDGypA0obLW1X2Kx72VJh
Kk9jAbRMa0ei0GwxgtZQEN+pCeF8inp7PYF8Qb8pRrvu9hPBJDyB++pLd0ImykWo
s7TFiAP85S5ZsrdYn4MhbMcGCm418zl5GT22lkQpe7KouE18BSgw9TN8l8ybZqCy
42RewAxubcGaSAyjoQuvhZ3T4bbFq0jR097JgQ6bK4BsvUSJ5MqliPAl8wGClkvW
+IK5iMD6bJdHThyjE2rXi6L4gkJpHojOusUbmpGTo5dZtRxNdgPDbRf7ePbtk8AF
hiMWhUIwGAc8UzF/sUphrp3DQo0Jihbj9nQNXjk69C6XMOuYr3XbNOteM3lPdXUK
OA3yujrjclU/sJw2QHifUY5TBgMoUrebd6pK5agWXIyYf7rBWeawNDop9GalNmVA
Q/YMdRmxg8plegQ5eeFuzsAATtcmSz1GhOFtr+IkAOZ3HRPiU83pf/i3q+WFRhrG
R9hZyBw6GuuNU4uIvvtZ0Z0gJ6OwB8gt+oSd4nzbXkABxiMW/ll1aS3YXFs1Xy1h
GzOxHuhx16Lx0RHAB1EDnlQjKE+iB+E5XuxBTsEFSUkRgsSebd5wi1kQWlp9Su9V
cYp88Y+DL1G9MC+9hDv6PVsGw+ycPXyVSoQpfmwW1e8GLn0bjBL60tCycMSlEv+l
HpgC+PCNMZnZ9pyaw+jFriejXchC9oI2orSMWwoaMvy871gaOcnJ+nUH12ZCeh4p
zc5PfOWGNbgZ88TsgD1bFAq6h/CZa+1ML95AwoprK2Go4ONp4iCICCs56DUOFIny
C6Y/ipTco0bOQYHpnBbFza7DCzpSUJgHZ8w357lekrU9xrvyHMQ43AjpMDTAiXjY
U1uS/O2W92ge3cSEsSvLfdwIjbYkppGO7NLdpkrsQEaAAqNrHuP/S/A9/vgQno7J
e7dqwDHwMz4L9Cfb13vC6Y4tAJclTBDHT8mEQiTQSCFG4wN0NDqY4TMo1+D7NE5t
1y0cSa4dDuLFlqnGhnFZA1+B0n/34EY8FxoK9vM+6if7dhyw01mvHPhEyLU36ehZ
/HfQj5BvhsyaCAcm6jh2T6EoPsrlqSk5eAlwUC1ozx7Ro11kifuUIZRYNGdb0J3r
EqJdbSl/zhbRCrn1QZm4AHPYny1aML2iXAULJAnB8lFC0a6J49gg23VYNdnwqhX4
vQMvyoemIZ7hQ/mXeCmm+szecd6+3TWr5tvrYYYuxxXDJKcqHF2TFF3b8sAc+F/M
N2xD8TNRqF7T8pjL09NANzktZjvnkRncsmIaC38y7+g5gBEBdmiU8egoUp0SX2L4
CGUBHhjq45w09wSpsxtPrPmadrSGTLM8hrZ8Zy2agxhb+e1v1VGdqwPsVYyADY3k
n+ebU+5c2aHyeT/Yq3zx6HNZLg1O5XRIJEcsVRUkPgeFdo8edRgV2nXerhvSEg8m
ktyZWUblqD2WzL8wjZ1q5Yw19n2F5oGyhJkQWM4gp7cVtrFygfHDlQUtEWst7Fj2
B+aI6Sw6k0c2Ab9Ref70t+aeJEz7bWuvIE2Y/tKFyzpNlE7lV4uL5tIy2nkIFzGe
XJoKuHTmZtA8vBXmXWu07t2MQ1d9C22q2wsxu+MiLC6g8sjoovZlQpyDijUie+D2
T7/K5QT5pCjgBRmTQz1V6zTmydhM4Ilp2XI4KCISLiQyZGtT5Y6huaKUNx2bKhP9
aDajHrim9jGdn6vqfElqYLB2u8Nzl/KCbpf5tmQNtfsTmhh9/0nXbZlPxhc6BQ58
xjucwNKr2WYbztUNjP2JcWgid3TJrHzlab/58epeKU8E1aQFpzL7jtm2TqBns6f5
A5fFvBpVvf0Y/kN2sSbOkzB8VyV3Kk9VUUvvS6GRdI8/Gcj9HPCR113ZH9onUsSg
V9khViIDwePkZ6troK7Ct31dDUKcjp562Wl4fu1S9yWlNPLr9axdPMs6OJ+estcP
pDJrHe0nZWwEvca9jOilwfBn5lKaAZoqVBltN7Qvp9zHrMuXuQefouZ2Cm0EI4kz
JT2uMl9ZXrzdMCGJ5QInNDdV+8T4vbupHtVa0mnN5yNT52rj4zDPLpluCd+6dMPG
0oUuKi+8eQRBXm6OTquxnrynYF/AGFyvc1mU8Rli3RksmR5h8OYVUX/FFi19DlwS
OAdMA5/ltmXUWE1xvP8PDfST1s6OMXC4Pw2YnKHBXv9QJyQ2Tk9aCX10G3EDTfzr
uFLsbcutTEEXZk/3MsHYZfH5TJpmL9gC6TDQsVwJ/jUf1BFFw4NkN4QPLT/mKZCt
UfpOY/CMf9OI7RpMiTVJJgl095zquMma32x1spqyoew+QNdRSAhn1ydcHF2HJY9+
D2JRLSeFsKvyix+b8eJx/32Kn2ZrZHbYpU9+TfNHD/mhqH2dXpSzzp47Zy/avYox
9Rxlw5ZEPEz2rAhgjEtwW855ex6+Xw61XhvZL+kmIQzuKnRepEOC7STazsuMryNX
Na/5bXHje5wy3DFFHhFaFjCdl+NyyH/29XCNn8GvJ6SV6g99lqxCk/DDRcb6Wrul
AI39DuRcLDZ3Nz+v/L+3u1MkqJ4wJzqMssU2UV+56Q1iAFivKEOQEH+xoPEWe6di
2MFUI60cN4aQMbeVUY5w1qci3JQ2rndpEBIwulnoNJ5BPNLirlAHZHq4ZbWg917R
ae/8d1T3QNsQrHQU3SVIFkLoW18Bc1hZlw1eYRfqIj9lAGjlEizVlG0qoyzR3ed3
olz6YjefJZvrpLUqKGq3eS2LaOFPH5qkhUKIgRHB6Yepla/hgUZDqKigtLeEM/52
X/SYgmkkgbXkXPpHR9WTUK1C9b5I0fk06Mo5kcxpCsjhyOpghu6eq9XojrzP4wD7
r69W5Dvu00+E1KMOy7hC7fRMKvr5bdUZgcuCUyeLIqMEBXLkGDRHIvN3hZT8NVTS
TYcPS/9iiJTS4ouDoAJELkqbKxrfPov18hyBJCgezQMXvw6e5zfynQcpp9abxgJm
jzEIUtI5tTcKbbKg5zorj/wKJQf+vzEssQQ1yVUd6T9rtSQYuWPyo4AWTtyK5EVs
Pg8HJOmZbLmerVK53LKwWlq7qA39waFT+ErGkygQotsAgd8ueC3UsbrPlqzLRtXW
z+yOK3ku+ReWnbtgWEIOVF+zOY/XFCibUHYjUNsIH69h+6EN0RCJRecImECEVK6O
frJv0jSHtNmrDweLw/ZiYrnqe4ix41NxuxB/Pzd2BBqvJJet+mxgz+j4rqSHq+dx
DTtOLnlB/rXKVB7N2ToggF2AxAISp45a84ViHwDzMVfa17+5qglyoTG/xjT8w6jC
6O2NJX5Xmh4oG+CxkM3uZgkOLkaJ0qy7IavwR0R2gQoHzy2FfKrsSm3XBvRKoxDh
7pcwdZOAmtJefTj5Xnx2nrwn1kqzBToFsy5GgflIQ7k6aVSI178D9869fOF28k5J
4Gh0hydBPCM/5jh/ocO+VFbqyEyw8M3kcf3tDukr+znjvC21kOIbVUBK9QWk96x4
yvtNnTNzGIVPbt3B+4NveSKVqJkYu2C0nsaY9p1n4X9Qp8WzQtxxrX4deTMbKqej
G6MxuB+LHYBqfSfyYcWDmaDHzGM4aAuaiGIqAnuv9X0CGWcpryoq4L/SE3yQJZsn
FMW1x81oKX4TUvXMf2ITIUravyr5I/b2cZ270TffleUtAKucGKiFezMD92ftiGxP
2KvKwZ7wNpKTahzyTi4R0zNS+snbBQ/VFizUIqoV0iTtVBsru8N2W9FBgZabvZFz
zh0tukr1hdFMljF56vJl+EFMY0bBF5vhKE3FzMpVqwZDfpir9WkVbD04FW/iERyG
4VhqgY1bLGzvqrC2FbUZ21kI/5MjqH3loTaBxb6SEdoPKz2rXXtWqkz2/YCzTm4E
+T/V96e6e9M7DyOu6xStdIjJKzuerc69F5VxvEYJx/wXcFviZJ9FFW6Rv8TkDEzf
/oirx8E8ZstXnHhf7+V6cpW2gooOHAy0VL3tSrLb70zy8n8sTEIYYy5NGhs8ITCQ
D7lT5I20uWX3VFm3DpyLd1rJEMhee6cDOZGhjK0yxnG3dMX367a3Ic183Zzl6FW3
L6xUIGjpqP4RcC/CSlt5kQgmAHoT4WqsDzFpwmQpJMGJUtxNBi0eg1pptBJz1VGg
1NO655DGDkZKxmQc9L3TXCmmv5efGQNREF2wGdRLVAgk4WLWyHrfNCMySeeFzYC5
l7gEQ+cX37wOD0OsiP4iOXUWkK42M4h0ml7TXuJj+q/WPcEVl9yCXt0OgiM9ggxc
25VGvu5VBdMhm+vPjBOlJW0R5H/B4a94ka5yhaMhV3k3E/JrEG/WLuN8htS5Z6ds
exEMSIUxv02u2c2INzo+5cmxDRp/zWgidQ3iTzXROUFY3DJKBLKWkpvPt8HK4GoE
p7nDdf5LkJ4HRgfNX5hcoXHjJkj5Dv3cOlsVwZtw7ZvODRsgDX1+WDglr4TfFuAa
9B97mIWm+XYY9ezC4NDK10N8PqTg4MtG6TPKxaU3aZirM5O073RGYqsITgf/Klkc
+p34zgik83/NxcrKYccakOxTYWO8hO7xJcSRi1SLNg7LDq+uJtt7IMSHY6KfFTv9
oAdTtpSPLT8VDwEq9U+w7xVtqBGNKwDLkXmMX41DuJ67eVn6fxr+VXzbTLOMDlQG
O39qWO7bx+QioTN4sEQnKLoMEPZgKZIHCIxnH5cmSogjy3bh7xLv8/dsp//laCzF
wnL/lu6MXc3qqaVK+nRHuoXuc+jCK2OtStEk49TcRt+44DswrjjgpB7ue1b9eFcJ
8ucH/AupZFpX1UjX938NoB1CsE/PX4mZ3zQxb9SRo0eMIIHWaWEpVnfg8l8dBd4d
4/aclKZwFW0ppMP9x/PgGYKnQShAOXyxVUC/xM/VTZ45TzEBIoiqkoEll6KrW/41
S3u9TwGvKlUnJTraMuHouOeKX8Ib9dYzDr8sz5t1Z/5FIiDwK8Zv3MtZnWhrCVek
pyxJrGfMLRLa2Z5EthxD8k4Sn8vhsIL2NJCjYDAaDTfoMG+dkXuazZZtYD79GpW0
2/wYgup6jhaYCZRiVrBKSzj/5UFnLCAFKH3eUQAizoaVlEl1ngfVhFkOLWaZW9CC
2sdUndYXqCNcNFdgxfxX6f3ACCTRs2lJUmOJEuBKqGukReBExkFBCZj3UL2g0ass
Ma7jWZD+vSiDPqoVvl3r2crmzeXCYuGRBe4cOnJleIjBNPrHGNZLjrcOhw9zQyiA
pUiNjhl0k5uVJ4RUsSZjC93MGFrIPBkFVUip53NaJYm6MvlUzxHCpDH5qsaJ+8tR
yDxpRCeXhG07cCDqAPBZnqzUZcjhRTFlkOxN82U6PF9PecJ30s8B436s8/LOrvj7
eiVev8MlgtpIUlBdUDzmeffOmKMYw4sNLIH8k0+Do+qFe5vDZKFTRH4/lb6Myc2J
cS7TsQqOUnuvaY3ZrK9+KHkvmivzLyDsBMLuxvmteKcfRe7sKC4h5Xcc+bL4D6Sk
oCizTEbNORmIifGy94GZSoEv347mBh+eAqBPce/I7uaqbw2lwePb6AmQXCnFeMr/
qx0C8F12MJN0xkHMIZvLpqvoPD4b9NZd1CVKx9zau4fk1EzJYyRc5J93GVGzvPUb
eQ/4hrfx75P23+VJaGzjgtnVBqFFK5vaAz+nP4jthP/uTnu6RJ26SmuGfHNUUTXU
k5AKFZ/EgN+goOmobSrdgHKA0es/mRgRJ7f6RCnWCsKK5gv6KytqHDeXf6lpO1+M
TnXSrFzhaG3hH7+JH4UnH7vLV5K6TO4ep/lWL6Ezw+KvAiLlklgCfCNlwBnpfxAd
U1TRSyKc1nWiO3RV3FscH9zVJEe3LqU6oBFhyoeFRf1F5cHk+DzLGsJzesWybHkN
Qesdf/HArmAcN5Co4PoPFR4tVlG2MZWRPuh5Ksd/OeN+I94WzZ87rq70z2xi/cFB
OfGNOO2WGVI75Lcmz/S2xn3D/Mw9L7PQ33G/i+BNKU0a7J/zHjVx7I4wkhn3tydb
kwGTrLriNlzcPRmhkkjfeqrsAeyT4KBNpjRKcZ0binzPvUYJWKozhYk8PBAJADjS
X128L0BV2gwYdX9h1uZgB7+ITAGMAGcU6pyNA+QQB7WlkxmYLddV1lRc3Y2D72IH
DmXfPMIXsIr401x6eMkXhI34up5gH2x8TNEUE1/fLrpUSG0s7eFZXKSWjaumBzLW
m+7Dmnnw+60NBihsc2FWobwqxqfz//WXdKG9wg96eF2X5B+FKV3jBLG46UTURust
gr2z9hKhm2Xt2zMdw6vlSgzRWc/SJtsxPgsTbEZpNoMS7zbov0k3r9XsyJ7ywf1N
UDgE+5TZFIS6z5sz79VS/WmCbACyKYWV/8eEsVaAlMlY1nNms6ftp6nHierKfWZB
4m+kXM9e5a4YefQT3QDur1svOs51Nuihfs3dJUh/bBk0soWmY79xn1SOoxN93YbB
bQ2JKiVeWcBDJrkpwOH5tDAMghe8FacRS9A596fvOaoz6l3S9TRoSz6uf9of+D3o
xrJX8ckj1yXXyfouVcBq9y3vPWVAW2qGmnFwELIdOUo5G6OyeNP/0HqOvpM8j86G
7+2MIwUZfUMHj6Trdwx3YcTygYqYRxwPpG41lTotLP2nC3dqO+15y57Pb1vDi1gN
Dfthw+zk712jHcWIqqK3Wz9+tw81EregschdMAqsT61Q1ueM59YhdEWZaLoJma6u
WXIeiZafJA2SmvNjo9KybhEgCg+Rz3FCxaCpF2vsZlLJX0bqLLvaySa+MpaTpGXs
b7eVyn1QDAVCNLBmDngq7uRoJuI5n8flTspgUZjL+9PH6Dsy+G/bqCRk4PgquBJe
FVsouAnLYnJBAcqoyfwRqys5wJCvTMqQUqfBiiXFlScrmjhAVg4mWJpAlhD8WDLk
kFoLhgDaPxUNvSj6TYw35NnC0Ho9NCSJfQVHIhvabloDCvjCqZoO8Od97V9RyWa9
kpQ3YmmuKxk4GSonRLYz0GV8BM7FXXPvJPc443lAQpindGM5gKpQIEqhVkZp23me
KLyDZ8Q+D48Fr2VWriiK3SW/j7QPWyYbOC2rbcyr3jys5im4R748yVIsisub+XjA
n5V78MBAkPlwSwIsyst4ZFmHlu4uigvj/SRjSgFPdarHOWCNkyAR0vBVk+fWIg4i
luQJgTBPRC1XAZF2NEP1GFbnE0YwZ2xA6XTO9ZLjNqe9NgTx8p5MCZd3bqhUMt1m
tUg80H/NnZJ6IO/+YrXL8Q00KuwWyWhuXTn3vTzb6MFLAoBNTW7Q2xTrcuamvYxV
zyGxJL+oyshwdmHZ8xWnvGXlKsuOFErmRoonNd6pCZItwgVG0RJRZxDjTaySJKlC
uR2a2lRIxdqMriFdg5aeUKqmGwsqcvK+KT43NYuUZVg4diidv0FhMGY4AbqBkyIG
qZOBY7KduTv3vFRrM5BH2pZkpv56VAaRHXm/CSqaQ56h5BcQmJxVKdoGFmm2yDKl
fm/tsbI9OM4n3Zg+L5F9bF2S0E8fwfcj+6XN00lqsOe0Qc+VY69Ncb8PvsASjuW+
3iCzASr4Fzx9zmPWvwiIhFzrQqZCLGesJ3B7u3jmsQ3g7i5in40JF1xDQavXVSzw
iDNUUgQ88fziMfkP50oxav09MIFhPAgNnxSwsjREFWeQRIu6EAcJP828a6wumw4I
u8UX8WAN6PFxtn9QME3KnJSGIa+NNqvmTyECy/GCeBOaogkUxfbTzhEbFVc7/+xb
MNZUHbLr84VCXMSvdW9G5Ueky7zv0IR+J0Jih0hUcH91nX6ef8Y3+/XPib3sOw9P
9T+pPB7EvaBRhI9EZzupK933pu3aAvHLFy8BZ2HaAYFORklXLLe3i5lNVkXZaIoW
lFQ27AkrzccpNasfhA7KjXTQHShrPBqN/NiDYLMROsxCsWXtU91LghW2Zz4dNSSt
5LwI4+4KYp3ul/ea15KygKSLHGxNnia2eFr+AHAY/S0IIh+A4gOW+4g+YCTmaMAq
aOJI66ymansQ4S8iE2Kitj6NwX5hOCb8ba9uN5+AuyQqgr+rJfx9SVi2h8ZplCkN
mrsPZWKHneFQ0nk0Z13LWsbReFVSwnd/JNdLjJsFB+G3pkrPVHvlI+1QGyED1Rn5
Q53wFd8wHCboUJp5dUtuEXH/9GnKvQeEZemIFOZMLbGxTSDoNe+EJXYExgpVuJVL
kubQ231QJ8MaXVZx1sceuLsy9n/+rIyod5xtznSJW1agAd1JY5p0UgNIGwjWuNYG
AhbXyIRu2sfdbM9X6xms8fH6mwKFoJ4S0HexfV32p6KXwNM1Lo6BcDF7qQRuXTI0
KWDSK1/F1a1/Jkho89q5W2rksxLb8MZWl0uXSbFr7AyvEbv8eXNIv18dEStC5MYI
GXWYwVlc5r0V389gQ1pBnv1x604C1hwOjbzZT3mq0HEBjD9zKOxYn0/h4tZi6Lh7
c80lFD6ay8o7oJaMGTIB+GJs41PVy5Er66d/FRTI+mUsrvGpAuAUC7sllyqKx7RJ
s+IMR51JHw8Cnf9NSrRIkcdq3ZjeZC6mm1hBDWHAJeAf3TJvbWyj4F17fz9MQQOh
f1/0FSKJva9OB/UI78YjycytG77NLHGEHPtXE46PjkYIMKXArCrISSy9raUm1dEb
v6MWAGue8fZPU6beho9uGS0Aa8gXdelJsuFhjeBb6tdkHbQbv5JZG+uDo+dXyrIT
z0ufgZrjJz9Ow+tEvMifBuk5JFgSTEEsExYM8FkYQUgc8OuUD5ruM0D/10qHWEZ9
sCIStZpRhlpwwR7NUBjhvb8HOB9Ow59u47Wdf/oW572QwCbqit9aQC/URiu6H3l1
qcUW7MhaZI0ZdO1mps0xWshSnLv/elyw2StIo8Ivcm6yFqoV3AuTEFmgvpgGuGTa
5ZTwkv/25PPSOE2wff8+FJbx9yl1G1GrsVBbXdKuh6TJC8AgydCcP3CexXN36/Yv
GdOthA2LqC20SiqlrauZjYPt9u2G8HLksxg+VK5YaoLNNmpLNMU3K6sXbX6Xlw29
T/Ul7KbMFKfFl792qPhyfG5vL2uyqcrmgTNG/2DqDd+1ngwj8f+lEbT2cZ6N8xis
qf3ZTao3BIItJOXyL4quz0eSnjFvQUBSxFjVCf+7BN7E6w0ZBuhBGWlAIr6PfYk7
HnBk4DkoIxOZvOxLEJ1PuPztfTaKenZF0wlYJNkIg1uFZAiXUAXVCu9E3eAc2VmE
A4eaf10VBhTaZEaj4wBZ3/JURb4uFPYG70WRRtfjCP4vws8uY/DJ87b0fJyzlwPr
r8vkpt0ceXa5pmyldfzwAjjCfECaHt0X1TnGk0Fn6iCtSK4kji0nHBh+iOl9M4Rn
hoJgqZMIKcrwX5ZSETtojWukreq0atmlw0k06q/4vo6jfViklhkfzectwYGEPCkP
vkQRixeJD/evZAhKLoJOXOoSbLON6iTAqHQy2YJr9BQcl3IUl55plRLYXUeQWdWT
V/t2LuMGnH2T1POq7L1Awu5RguG/R7gTSQRun9ireMVG9ju+meuITndp0vcJss4x
yZuFZ+YFJc8oM67zd7KGWw4oY3frKTeVgmh6lqYDHipRaN/JId1jeSnTFyV8iGMr
E3vq+cjnGgh2tcyDF6m6MoNY86LRO2He0bA77AOrtUSskBHQ4atCXftNWK5pGG/8
2h4/GK37RjIWQxj5RmQASxdemwQB10S4Jb9w/fnq3DmTQ7WPQ2diUUn3Dg7uBj+d
BnLWYJ/NrLEWr0/w9EyLMMgfcZJp1+HrTUGzG015iPBzAdmL5wmNF2PyGfTj6Ne7
m+edPWBL1GdH98WcyqvKrJF+WWLInvOvbLX+/LXouDBF+R++O4D1SFnNTgAcMKt4
VSVxl2tGigGRyN0jxUJ2MJYUivmiMIy5iLgrjTlAHXjeAqRbHykU/f9zz3djewNI
ntXzZAvIqijIZwpnSHP1fMsI8R23Zl4KlLL8Y8Aru5xGciAD9ibjZw7T1WHn3VHY
RoP6O1svmry8BoSiWgwDjyt6VpB4ZKxmFPeruUL81xxYB3OUBXSiWVlPGPBzkEP7
ij8/aHJpGpsn4DTNHvZz6XGNPqUZ5C2UHrHL7UQNUkLe6O3KZIUEdLNsTgAF9Wz+
NLueojYIBJYJDCLqxAljjxr1wyx/t7t/31l6r8levJ6PA9kFRwpnlX2uqIuYAwUB
yXO3PvEMc5truqkkgPbGUNZejUjQf46ho/U8w9nsfPHXgP272XSc90nZYG5ZtS49
UBcOrIoWOhAI71PuLZYyS4lny2a29ZGMuEVwdpmYCkQW7OFhqwB8G/1gSZz23DS5
L9ckVodOQ1NvKjdjfXRWkQTd2Xt1Xmm3Q8IDetfxEHmMjd6xB1Fjh/5TCjqSdmy4
im9XTUEq0H49RZsO3yetpTpN8bFQeO+YxXe1tczqLB1A2axU7t5FezTPk4LGCYPY
XANZbMJ+H/E0XU/lAE+ckYBGVoIUPwO+o1kDqNUTJTq0fOctqS2POjrDJf1W5TL9
uPfON5NazWG2sLxHWKuwrs9N6Nt1iPEH3ABjUmHpEew1kcCZVbu6iZVUp/UNpmGl
10gyP6saeVyfrd0uQRDmk98Ek+mGLw84J073gLxSbA0YXqaKe4ln3qPhMcL08ILQ
BcZfN+VOOUKY0YTQVQhp0aLp6MqxGO8ja0SAIJv70unqKOTNsg2b5kzA9Z3JimHk
Te9Ku+xKueVgjTUSQcUoeoA6bWP3swAfYrvaHurLIOv3Ohhpp/fKPsnxXzQWcB8/
vm93vlq9zumX1EZvfbHxpc+ZbiKomuNOVNkIZdSE6CUEh7OiIkdxU1MXtVLoaqoW
WkcfAr6A+aV8O6aoINwO6esCfIRWnaBqr1na3ooZWc/952F17PW4DLQxbjFlU4HC
Gp9wGdk2Hbpq6totnuxgojNPIjOe/tRXdZ6838KCkIGmPmOm1d/ehMHKJ77C1bCa
KrSBOoACyS6U0TJ22H2+2JWG3f+c8mfyRm6xxLC0aDFE+B8RqDnsdFOBWAaQjTl2
vcUQkO6eWQoSmZLiZ7x/X6nLceK+E5umtbgLqNSLUSG7ljTb74N827sTHfoSen2/
G+go+7nPM0blG7tV6D9ayGBlTKToHiKrbeBbl5LEDDteuM8Dnt+LWYb945YmQxyB
1L59fFxp2IcRvI4irobE2VoB4ORHDfs8cVM9deJkxD5cnTFCgUcGQm3OgwzgmuCh
POYNeXs1Rxit+N9KMNpHvFvoZM8BSew9xZuanZlPuqOQMEDz0dHXxwgMACXu41JM
y4Jul4zsjRA42fjxOFgsqoMkO6SNA1GKLLWtRqSPTUNBKOORXlblPUatoPEhPXxq
EpbRzrTZVLoAOoVIb1+I3A9YE2HH0kfHYhdRIph8GIfGk3TN9zvGBjai2lsLfRGp
o+zui59kpy2IPdwac1lJXzZNCLuPNPHsk3KrUJ867LE8GdDgsxrNBPwVjKfDBvKH
OiY5pFgN1HShMkb2WbgKPZzSafT6EMwfW97CbVkGvcWA1koYmVkmzQngGkEpG1VU
DOtTXfDxRswPU4EZ7+BRZfuhVol7ItUJ4hgsKN6vV45SI0vALQwIv6CKdRTMn4Pi
x6Do7n+QqeDYXmhSjT57ljwiMwe2euYo5Tv67S2kkfR2OuWaBWGrZuUpPxqrIdeu
l7TpxFPpEP0h4RbQq2OijLy8IjJk8/4glWVBTmyrxDTh08FTQtoc966i2MhC3WYi
tNien6IM6AlJuE28bsACtzdheLMXeQgNf54F/eQMeVm6z56LeleqxABRHithZpK/
Hb6eDQ/cgAQn+Qh8guQ422fJLAeCOwGIUius1pztbDcaYTaC7UMpAu6xOCiCcEOH
Cp7msvQXd01xRgeG5lK8YUURxHz+idI5evJQqwBUaz1bgJa6hskMaH3DdVaVudeb
G0AfmkVD2pCp9rB5JbghIMtvEw9R7B1OV+Mz/ZjeprNvWYv1risky0QdFsgR7Zcu
rceG45u8ez9ozeN2NMvfnTMnVx1V9gKrynd4/5luFnkUpiIkU19jWS845C3mbqmG
5rw5bbrR2s5GLCZdtr65SF/vMK/Hmpb3zSUY6txKz6hcLNF/kjaSFYbrHi1n8wEK
DH2vBQZSj+Ma/bxARrasgotFw+RfGP6RKL4pY+WQ3Hu5lv3MlnejwB+0sQLxS5ff
WhTMy5HLaLfracqvrMNtExBiGoiRsITXxOvyDwfd4/T/umNelD62eQD2cEoJuTKx
dL+mF1KvGMD7FPE93P1m/pcD4FhQKAhwE2vgTsRu26I29BbijfoEXoT9AIVTfVhm
KHyDQqUA/+A2Rzy/1FD3A9Zj4vxV0sC1Lii7t0OOMC0iPIr7UI/AaarkWmqbG+Re
18qoMXO0/F7cJcYvkRkt5SFFRFLEm+cR0/cVPapzf+6Q3QOupB48rNfb1qJop3sa
SlgpfwcPPDjpKhc3f++8tskk2ZrMwNM3VCv4idZ8jLjw+tz/kebl2bLhWw0qBBHU
misLicM5RNkTrFnpNRHAJH7kgM2x7E2Nwp+8Xa2wPwyWSUtcVQUnSGxNWb7DKrMb
Q3t54Fs0XTPY36X7M5PNgQgi8BsBJ37firk9rtKwjW5gnxrt0bSkT1MYaldZPCV8
031XZ+L21P0hVGpOS1c2ZkLeNpv7hSTrEdg2bEbQmY+v1ozOO7qWW0R6tWxHi+7X
iyeCBirrbRRi5zb1dfNFSg49/K+1JSDN6Q9bVclEWS6gfNujwpl6GKzBetCJVXvu
xhigWJxMy1sDYoRKsnzv8HgGZb29HNQBn0WMea44lRXf9/zO08l4j0u1gzTjqrGH
jZ8u5MiFmeGjJ9r0t4x2pUZ159wWEmUpdfl8yKlgmvHbv3yA9woYeCu9xIC1wWzc
1f1rhz4KgFC+Aejg7hVVKmHz+FufV1s173+7eYehDH4v5kOpYca1eDFvf55npjmF
3/frOpvlb+bEIhl0I7UaTKpp0I0hBSaASjWAlA/05M3P0WTcU2nVM55jts4yut1Z
gGi78anx/gbdzEmS87Vp1291/EcixY73XQxvJoKy9aUuApnET89JPGFfiXFOmO22
PHEO4GFtz3aoEUT//+aQIlX6jhG+rAgMrJUSHelxXWqWoSHr2oLpdBvhn1t9HU+2
44IyXL3NHUmZf8fv3NJhFeEC5cM9EvFnLfJ4fwrc/CUSLw+xBYCpGSlA9nN+PEZV
mYB+3X8fXt3mCdE+agpxaO+RVRb6bXAx5Pq6ZKHx+e+jGBqCWlYQsjwFT2Az5OcB
YAQjakGhap3NqT6NK5KBhSn5Pz68nkh/G3ajt2TSgYDCDqCJxFl7YvOBra/Uiufz
TVq9gK9myokvZnUuhD7RrlHtj0eYhkqYwdHyk2iORzFVi/BhRT46q+eLQ+T0kunw
8E5QrIgTtt7vhju+FoK75JlUsilLfoJn4P0Kdt76XjWwnXLrL4qBDIqskurASnL8
3dxYKkufPVNJ4Zvc6RLxKk7xdhsqrVKxBDdNNUvRFZSR7O8Fa9EIRhgT4V/8GlSD
GjGTMS6rphH8c+Tfjn10JhSFnQDK+OjeiBxhBKhvL9t4w1yzn5ZjUNmNIsX98pC3
4GudXvtivTSozx29uYQ8xlOTreUKr4Ow9I6s0obblT4Fdyqm1pEXBHt4RpiPUdJA
+bdeXo/80oHiBUR8wLSE+5Nu+Da7ykl7cPYbvhU4zZwpPficlUNGUAqpZTex3adA
cb+mbCtW3clFEJdZ2KH4UPLGLquHt+8T9cxdr8iewl60Xp8bntKo6qDoXb4/JYIx
xX1SMGg0leXZCtQgQMyGhLHsvbqyAk6XTYKgHUeJJFu0xtCGnLZcCaPF3s5ftqtA
Xln4CYhjtxpcUdeY7/7xfH5CSPuWj8gj+LS+EsGWzUF0XcCViLMSgqy8y9I5kniS
DSxSYAbUv1HOafi2KzXfnrGoDRUyThJBt8xOiPO+ncwDuqHX2I00pDdBVf6F7xwG
af1kp2iNhr6761oijLZivFnRCeAz0sKqtb4wuUVQ3+fA3WeGaLzUcK0nXFHsjSqs
vUcb6z38QS0why6ZlwMnY2iBnBv8uHaKLSJHqFWI4UveILzTIB+r1EbgLe6Qr0v6
oeCg+et+0Pt/fPQaibWXEOHNg3lk9qt9aPTSG84XHwzitpTwlqWz/NFhB287fyBp
veEak5Um0D/DBNS4Lpjc51rIxj2XYZ1zQp1/7dQ0uhySnFFR7tV3O0RFWf/Klcvq
SiyoUYMyfuUxZ5VpdOMXvgjN6tkunLGn7OLpXJEVdWZ7suyy0l7MTerYnttEImsg
PZY3T0SQHHq7os3NcRCKx0lytsculwEJj+ibSsMVqgKskaGHZ6snLiKr5PSKrKIS
X70zhV7O8RzuYGnJENiehypB5uSWzZFbx/MEH9A7Xyq/GCSoTvTloABBkM909Qxm
5wWug1IYFS5Kn5bxL/YGvI2H4UyHOn0YkPMVOnr5ssUAQ5oyvf7SLItG6kAPigFt
ER3SjL/LqdiRkYHutlNqtAvuTcxCiT8/lg++1QxX+jkNXWCjI/wwrgW2Lau9Fur3
v1k7OScuLcPWB5GoQFsAFjVw2OSnL4BEBlznPZikxzBkvKWwLPHs1Y3FlrBCepg/
FLvPTa55i5EdGOf9zPRuwlpf8FriPO+V4kRFPgim1/NPssKKf135ODcDJwnkX13m
hEfxGPTFN+mv6jt64DHGAR23ekipDEc2zYk11+jCrLAm4x5mJ72XWz6nG9HT+r+l
4QrtBeJh9CzYWIcZSNY1gRitj2Jo0RinIr+4f4Uyv0Og81CIR99dPuYrAK0ZFAbZ
PIt1rkN3AdoOZW6WjNZK8PGMhR/wIQf+MsYq9oq47AeL84dkzEPjM4ja0/A2TqjG
1muM7wsQztqZNZ/z+8qEBnn9bDe+6mVkBT5DlObEkZrCTF4jD59qgvR5T8Jc1HzH
JGqrDsebX1gSe6bvVJVAF5Sg1JJpUfbRucZv4lnA2cSYRNZjUJK5NVgh4aQ7ZO/c
CYnniwD7zYR1IEsiZe4Id59WQPTQ9mczIBmRUBBVAbUY+B4StinUD6M4dtu+55mi
hAkCyxuQN2EMa5l5SirN177/8OpiViYUlHBhYDW/F005RdX78ODofAxrckc7yD0m
jEF8jKDbAFxUsd3S05GasfPZFe7C9XQQb6L4sXiPGK6MrHrMIM2pjzUCK3V/Gt8H
79HGvqUD1ONWfTRPI4HcmJYuO3keA5V40I7+b4yz97TPd6J5mJ6cI0w5PM9qxIga
ew0n1rOPqOTNWLBn+L0U+L54SUl08/hPxaDpGrx7LqEX7LfLOz0kxxX2533Dv+vl
r7CVUb0tliKAyIv+tjkAc+T5LcSrMljulke9xGLHYzekE6pDn7mfOAhPpGZv7f8x
T3Q9y5P/smQpNnUb6Al6dJwF60BrQEFaNjBudyE9u05QtlZQevTTjNEs5JVP7srG
2kt6PI/UzqHV/iuEKU5biJZrSwjPCm9Ts+eCgnfd58CfBXbkbA4uia/GZhdbFQxp
g3AXGNfivNI/AX7XejUdGHMuQHloc/wb9LD3ID1mCtgvzf5wnla/4qDJwO37XuQx
kBhZk9cqF/+kTmUc/gknezrYl/OIlUvunu6T0WamYGJ7Ipj267GHGz6zW42EYr2m
EWbFNCL4BqJhM3B+VjNfFy85MV1l5nUDwd+E/2U3nbqBORbTLFF2l8CN0UvkwmpM
KgT6Zvd8sxjEd2molGirRL1s8epmTxijgDOwH3QDEWxeYZETp36B6r+mdp6R0XGz
pbYAABEHRn1wWJ+zYtoTvo870fQpfEF4xPEJs4evvTamKEWM077h3p+zSix6dUn3
BW00mYupl9SOCZS4lSbh/81yDUbT7LTWPFc/ZByRgh46h6r+CyLdzOx0NNt7hvHn
LZ/Zzj+fwf+yc0Xb25VH93mFfsgEYicgI0uWAclikWY5SiLBIR0lvxANjTi/3hOL
FH0Ne5cWT30ee1JmPIdN0EQuYbrj8C90jJ7XYHUxAkK9PFW/2Wmp9evNkirCWhJn
zQoonMlkxergC+6wFh2rLyYeJ+IZ73sjYxgvfhQetH07GiRdY62x734sFKxnQm8H
pypEupg9DLhTsW74uaU8n4FPNIdSUJ+gXLKAUcPXkT2qtjfSzalI7TInOcVAx4/n
B4eu+JM879sJhvPdLq97q1WmSC2pGChHiEUkIZ699h1tbF7nVRLIlA+tp29pOkSP
xfrC6EeL+pU6h5FavsnQYHbXkn0vpHgKwAlLYgsWIx0VtqEI52obj/jzGWIbOYuh
v3LM+sePJSVL4E2E0f4j8vqXKo1vzWaP7crhk/X0PE49KQRFbumNt3j458YHZ2L7
y/I3yASy/DafWEO1X5zFrOISBgWALrnD+SxGEwZQ6xsfK+PAeSzTpRvTyTxngsOy
t2Paecgux9v+mYF+wTFeA0HV8SmxL3y7eGRQ7A/aE7NA5MJ0CQOGdmzB3EmI6bRp
SfDEpXqoW4bgFrcOL0Vg2kn52tS/VfioH0LwAL7QZ7G8j5GjnNP4BdNvc0/Etm/O
VypjhLKoWTJ/xEkDfOcgj/qYGfLSnHCq9oMHuoBIixk8WPaKBVXofTmuKqbrPWcZ
/fsZVM+kNO5xn+U5+lt76H2TahZ2Rjrp4LaefUGNPL0nHd+mVGLkUCsDzpu+Z6JA
ER22jA24rna+Rnl30zrE+mBY21PgCxaZ01HKOwoT3VgiiIpnZ0hyRCP7l21gPFK/
jkHaP6URHAmzY1MQl4Wv0QdN/klS3RTJ/P4jtgFiC1C6E9iQqqzCx+kh2v2iHMCV
SBi8MRNLiau8qw54qfdvcS74k7ZyE+dZdY1FmGEEkZyN245sIhgaHcedT+J6Yqt6
jrRPx/aM+MYgCkgsOiMX1ClStgSmRzffXuNqVOdJb6jnVgn63sjOit6UOmDQolFA
VIJd1Lu1HDqh0w+EJlvFpWnJBb+ALTcGtpSKgWIYFDAArcFFsQEnNajJzdfvINU5
9yzmOl1gj/QKhZ4uD0a5E4qhjNR2VsGlkcfVseiWXxpV7Hs0BQweVyWGfKPkkkG2
FqwV4nh/wr9jcIsx3RhRuKia8jZ/9cG/V35GeCWHPh0U1lVOMi+iIuh1Hn3ynP84
H5AHDw9MxLsRq9o7TLLVwMfVSh+zihxwhVo/pXQKiEt4K8eGdpYfmKafUbDxcTfN
ujErGqHQNtSMa4NFLwbJWVEBayz/MszsaynLCjbZA8boV2ZwtqSbvduxultsMoGf
5BnK7CXUeUNaK50zNzOKONnI9cPTOdhl9oMDku/eYEMSQMJS1OPqq3ZVjOVj7jYP
6xYIHfUbdphr5aTDhs+OzAR0tMgI5jzfYkjL23acxZ9ZpbWcbD9SdISMKhxhux0b
KVCR6SyP87P9HYETPpsL7Jn40OjLERLGQmKuF3bv0ZRFYvXkUkjgTPwYs9keaQKl
x1ARPAaNRQu5iCZaBeMRZztZngtaYnT8qboZWojao+cdxPNuSuiJ7QWDXscv6FUw
e+8JmBsiqkKJ+hw072hm5932Q9nKPWfzqHE/dcm0VlG4MIbI3avpSlurdQHy3reV
gRZzGWMWgd5w7wZtnC4Rhtvw5f7Gp7KiTDZcMuJnArkdD4dySKArewbQXBlr8Nk/
vEk2OYN8Wvz4h0O7BBLbXhbGIG4wjgNZfC+yUy1NDAzRHbKOPhcmGzfRsSYx6BJ9
Dn5mnnahVj6zy7nSUD2rk9GTxbcOVEpWSg+wqAsF+d9oXI4yZ75+F8AoT4++s978
BTQpNHpWYTx5eCZvvS7CrLkLcLZAE7m59KALwIK95qJmzKge7IWEduaat7tj3wto
EtSW2GQ+tQG4st7o5gd/GivI/FgrchUe6k3wau1flB84vWb5grnMfXjA/gWRS1kf
2wQuL/EzzPMX0zvpN5bxu40FOPUZTl4Q8AFAhZtE7sp6u78CcP2IvmCjHkiTFaTg
D7AUQ19PGoziJ4Gb5ZfLUl1mpS/ApqvFlEzsBNKdEN27nEe2R8/Osp+cxEgo0fga
aD4rVnjj3GpxRugmV6YXG80yxgeW3FPtGfao5+3lmz0XZmuMpKXOqNbdwWyYI7KV
YzLowSTiEL46XMZWgerlreZCOGmgsvDRflNusoQp1LXdhVN/6zOXetd81A4l5QJ0
QXF3xf2ehDGlZu2JPI9TKkX5etwms9HTAMp9R85NHXXKakSleaKHmZwazxSF9hGm
hmua/W/SHyCMT93bkXT3+ggbygGRpZrrqUJ0aGU8W8fm6BzWrRMeslhRUPFrj86L
KcRap2SFeNeK+Fj4PROIab7masy+KnSDnUM8x7zh6kG4D5a+zKYwvcO8GG2uTgS1
hYD8lcQ04wq2R1P8oaxFlUjZp9SNhIeNBc2c21zD23wvb2vrZ1Z2DQJd+zF4FoCs
cKbKoSnXzZ9PmWDFStuwdURRnUejEhBHed/CwFcAieDJwWF7YI0PSQLMqrESHgGK
ieMqhnFLDD/h565rPViWidOzRWB570PuWuJquo2SBhCaOiZxDJLbiw/znSE0gpDw
vsp72GM9XLXr18D+IWiLq4z37yHneC5PKHwkq9AnUo2Ifg2T6K4ADhtv/pXpxNyF
oAwz/jJj2Jpi5h4m383l/i2kKYAMgVbxLFv2jBwcn6SPNl3aQ7m1ZRzLEabpng1v
GClLhd1BSlWYdHmc9Mr+NET5Nd7hZCNmjQBgyhVQ4Lc/SdjlGlxmK3LVJ6J6M+i6
VxaSv3OxMUCKyPwyrlPNsysG6q/mDIaycQ/EbCLHzQPR+7X9kl9T9qmrv6Kx9j3o
oBxYaV02UOibASmPgEnHkgOB5gABQ/91VhovEtG/TdVoyOiAG1j/tiGCfz7FYTGz
/tdjxAXGcyce/HHZEaAKoeHrUMIxfV5KY0K2p4HoO84znpl5U5kKXYzeDqKBiOZR
Thmsm7pBFOhhOEq/gDp66nGBfOzjNTwr3x3f4DJLhIIkm3/BBHG2I3Zie6k5h7dZ
PsNMzsQQ5fwl0CUJmxWmZgtV7Tk4M2AqcTGi+CJ33GWm4wgo50M22z180v7X5CvU
YIDDm5kj8BMHeP7n8Qt1MOm/Pl6V+DZG52ck2FW/WHUw4dSrVyNw75S1QVdG9CtD
lmlbSCgb3mloJO3hKdZ8q27gmK64qVG+xr6JGIT2rIPp4qvY5PtCj605o+cpMV0u
6XozrWp5X2oOvPy/7HauXl8kVph4X6rQbUmeyul6AgKia+thJA2us/Lod3JenrEE
nOjV5eaJYt8bECklvoJqSGNDdA9XVFy0evbXvR8Nvg/xiN1iZMl+j0UWBsyae3/Z
XRQ45ZZWc+Me2QdfHoTvUf/zVKdxaXushC5/KhNQOxOGf5eEI+BWj/AX4rTZIfMk
CpmaG8QeNsd/4O22ksfPIwF7UG7ZMIuay3SLkz8e8Tc/3E/1hhXOXZGWQ6Jj06rf
4cE57Rg2ZKNdYEelOqclaLRTiKXx+mFTE1DRYKltpZefmBUkQjmDW/Tp/+WyWqvV
qxkTWEALrRn2t348Fj4klwYw5XVqDW/Eyet3fWEivXiZ/IF3u1d+lPAu9zWW63B5
20DQEme19X/BU8/6mXIsmvKPrHfJKQuzqtpE4LevES9oNKbAse/PlO4nbYWCrJvW
+0qDNf4P/n+Bv8MPTk2EPr9OrCqWD49UfvS5VPvrjT3IEfYbh196mpr1aND0cyy8
BLyO4wHhfYD6tUrr0MWo0l6eyw2gihihzC5HUwUltV1908Z+nB1J/I4ShPnb84dh
2sI4kkL3Oo5+OPyhPpGVTyyWjKtJgSeHS//CKT/zC4k2FtOKAmVtpOQ0OZKw08Tz
QpDSH8vgZsFrGb++P0SV9p+gZZDOs+jEI9Ze4H9u2d+bNPEKerDMKPGYkXCsKTeg
e5ePQB4BSb9qeBatTd4EkMVG62sup9lDOa7XCP3ZEV1KgzujxeOAj/lxGewckix4
iXogHQ4XvP6l5mL2oZwmDWHtIqOuU4YQ/X04WPKpZyV90gCOqL/na17tqSGIIuTx
Lb9DYrtnTE0PH64JkKpeAgxFXGyYDCCPU5xF7a9UDcEgHgv2gxsfCKRu+P8ttfH+
dnZ2xJi6xj8RueOC4tfaM0y2ExVRMLjSQSuKTYHa1TN/oIm2bTRXw2b1jAl8jlJo
yejc1dRpwq92ESxme+PLvGZcy+0fuqsDOWtj563ChcShEMw1uumD89tDFwJtY5hS
JZ8Yb1HoDbI2t+ug79+nUVlL1LxMpwmoif/plvVHLsKxWphe1P3xHneUGq4UgZGW
2x418RgnarHbLejQPWagve+ieHcsZpY13m791krT3y7url4eDujMiu4lGfUMf1tP
n3plFRi8/F99J14LROzkruA3RpfwOtKMiuJFRTb3d5Geq24dI7QKwqK6VvwD1MBp
7ar18U5Y7WO+2w55HSec08GVgFqJaP4ia3/oJUO6gD+8Q61QnCQ1kCu7dINMYU9h
3MXiPrLqB2bLq38fNyXa81jVG04haLilC2FSNR9NsHXtXg7MLmtT8C6gKgefq2i5
XVaPYSHqd9+F/UfhWJRjGNGELBDkqn9s2ni5OPVQHGpUu1KTF/UrnceiCaxxTykn
y0vV4ssbQDkW3kqHZkgTfwsha2PX5B+M7ZtLBMB16sdcgS/S5TbjzlTXPmAmFoGN
8o4HJ8X7AvlwDh54Dwicb0DRiRvvNJKa943umuWZ1bcQpZG99YvTjN/KEE/RXexe
W40EZv1OJKqDbfwJ8/2i3PHBzX/9Ynd6CqAB5Nx0ThX+vyziOFQNl/cYcM6SonoQ
K8F6Gt7fl3PKhMn5X4hWSJmKKphgMu+w+EWFqTxxGw7Yuuszmn1Kqv7tVto54xbP
81kcfUB0tFm+Kk8z0GjHqmAgGwPH+GhHyoiFDXvjyHyrLcuNkSN9AkdobSUoYCjY
oigVGTzY78bDs/E0nV+3j7lW4cFF0zcV6XdbFlJvyxf8IS8E/8LcWFcoiDUxRvEN
/cags3vaZXoCwzbwxbVsATUWCuw1TCeDcUdzgcRgB7AcTdnirvu+aVexrw/779Tx
7dbm559jg3TA/CZCGlPFfW+td5SP0vsFi0xT7NhOJ0Hrv92WbjBTwTST2oKmEl+n
wuJWmhn8YDYr3ds36sLzgVCysi23JeDrrZvCmhnJ5alii0bPZ28ngwLOIozf9xaO
Zcv6GMmcNI3M2T6LaLs/GGqqdixb8r1gM5QPp8B2AL9fNTa6K9LfFzkFIElM9Vwr
0wvkMS2vAVD2onSGVXEH59U2pJc71nFsiev40HeV2IP1NlFizkuLYWX9hjvnvg+r
ZIF4YxHkus0jPuaU1InHPAWKYmqQx99SC/B45W/In6KH0XTEhxOb4P6z5CWIXaM0
VB78DI9PZg00euQyHWbayr+chF3pbZ7RBxFUF1yMQDwbi2OB2wbXMlq+miJ5Xim0
EE6fzXmp6g1tQd/2LweZOtz8qynSMcoPixbOrcx5TBgvhzlFKBEDOUr1g7q3jMIk
J32z+tAmKIssgCXJU8thOZXT8Q7Xjoi0oiOEIi0oMZmZnFmmmJQGkmxaM4dH/W0q
FYAD4l8Q6ui+go4+2mSEesxt38Zw1N0z5hxhnKoWRDm9TS4G1NRpwpiVDGUts2E5
/uBKyJu6grxYmrOqI8TnxDC6A8P+laiqETS/XEAxmjCVRk07o/PuKcefX25k9Q3x
ncYWomQkcQokFSPNCcH+2TVzFpZ2ajggUaC27P2DEbNV7lh1X1yUftJIX3EqVZZG
RhQTFlB38Bh4e/tkQhJzFE6sXw27D/mE7FIitPb04yxpCWCL4ckRzJ60ri+TAbAf
PfEwzPf1U8tci+Trp8OdyUxfUYJRw8tHRIXiu+oAvOH93dCrQuxGe2RlWgDedBF4
3d9abUZKUbcTfyjL8pKOyno30zfmXax01neju57CFnQ9IuwBE8mqrLjUQ3cxucPZ
g+I8aIVal/9fSt7bg3Grp+kh8I6m2rwI32qRkA/cnJBpOVeH2OuAOzMBeCTMP0NO
CX74uGwlHFN02M+qs69f9gjgz6S9Z+MTheetXH6W4BKSJ+nKVjtOO4PBxvqM8KR1
psuFzF2o+TVGuenWfrnBjIwhhz98Xosg+g0lcPmu9xaf4bLjJkCu6CTz/zbUhnuj
CJ3z7GeXpJqvBg9g8s3/0XtR1D5xXs2gWJBTPmNYMQFUqD3LGcYTAWmSUUlaX8XG
Bpf2cs6UeYYVuHgtGwlArGWRRPNiJN1huotZtcS7noligV1Z1CU+Bav84vlMQjmR
3VXSBakbVY/GaVbmVgD+5REyIxIH6i9C1QPe1llIJDHKW3ZrIS21mUp2+bY0PhS/
aBj7+/54ZIdxW4kHk4q7nIwbrJ4Wg3GEV8Fn+N49grNe60h+fPFKvWKxTZ73d5bZ
hWoElEMDAjUBX9E2p1UO4eScguhiIDC+g0nTfBiT8Zk+4tOkPBxUFwG1b4Sgyn+Z
HxY59UXtnrUbfEU74rwRDz3+Suyi0a8q+VybYq+WZ4oSiYWs9eNuYMzEd68l8cy7
Sd4ilANMHdMUL/ZAkswszEcq389XdBJ+h7d5nTZlkQUE+XiD0vIdSoI5M5lpq5ch
c9itTBmsEasSdS8urgBArYlm5nyFSAgywS1lrScXVmg042Z43F/nVmvpdgMrR/Se
ZfrxzvDzM2JNVq0NxnQAQrjGq6kL7LyZxO9i1VEfpBvOsjVZZ2Dxf9myYG4c5H6A
DNkUWYHGFrSM8EjK0tI3FYePtp1KEOtXii/Xj5LXVLrcJtZ/Sxi6OtYO7RnH966M
JlL2KU4xDLdQ+8ac7DJz1Y9LAhGKk0IvEJ/od7moQ62yf8Y3KK/43Od7cniv7UaK
IkwvnOJi2BFYpXiti44gAkF09GymOKDrfCSVqANsif2DX8E7OvdXjrea/H0fdCMF
e0zrUTxvkXz9TLdxzWX91z0Fh/yUX1Tck2edr+K1V/J1WnU/W8U3MAcWKRk7rw8t
ZHgrCdgTUI604gjSE5Bc7EnOcVu662q+S5aAWdpx/hehhKrVYOmgHwVIqAjeRG00
XV5pmewTSimiNWFfLeb0/DFZXO+XER2YkIr01NaH4qYj8DQ3ymaZNAIFhSN6AlSM
CgniBw/WX+RYFQED7DaS1LQl8S+pxqdyD2HAmGIX6oS4jv0Wws81RsGAVcucNCOb
Az2yX2BqdyG+V3Jf/TGRTkXOHBedY4gDwu4MS4YUi0vUp2ea60qQAIrEEKx5lw8q
NQsb1omgYe1FyMft7aGCUsjWOWCkOZ1uDdQben1yS+Saii5KASOXUVoPZ57NX992
R6ZssXOL2SewBAfgC5Qz2c8hUokCC5OOhTeOhRXPSsCJnHTixvo6Znh/2noGihwH
k493pylBgMIyx8GErvH6nF9QEwkxCwxakO2KYvm5mZMKAzSA9POew5U+f+tA9D/Q
RXv32acMBLgmZZqnMfZKwQQCj6C3Lli2sR86cTOgQ0/qhvxooFShzMqDR6+PoXuf
UPRzAh5RpixpzuO7O3kZ8G7IulMgmz52KnTBm7gl9B8VnBiVMUbxWs2F/3UZHEOi
t8v9rKlLZ9ISyJOgq6M6gEY/a9/xrpefj/q1IBo6Zr6oUh13qyywNZIp7y4bK9My
tgsevwCz0ZZY55WXuapKbTU5gp1uC6FEOET/tQETyl2ySayZbfgdTCnIQiPBd9fR
zn75i0m0xzPOdyvwmMAOtyrbVdOR8srqVy6cGsJ45FStGx5jipqqerHuRp5aTwcB
9ecnCd16qHMw5+pKwbmUpkOqtvBHEm2NeDB/ISVHEaKHjR3Nh45my5a0eGXVNcEF
ByYrQ0TPaiMfKhPXWDeIBR1QO0k3/hdUCHntYcYwE/EzBqTwXcF+Tv2YuDQAllvh
XqGe/0rAHbqLARiv0j4Uov2xjcw5yYovP8l+hfRpVlL043AhAEHXtFMrFTAZnfIc
7KI3NVfvQvNufeKIyijvnr2LZxrwBBaydxSdGVCaVr34fBK/NvwTVd4do0g8gOjU
x+yTj/Sj+fGBD6OfyLhZJqUsDvJAB8us29n1EM2khYxxSoS+nMT0Ox/DrgpQ5OXq
yA+671iCg2sxfsA7vMUMCq2NueB00d1N3xRnYs4PCMosT1mgsZF5xlQ/8Et6YEV9
CBptQKIw69Q2swCXg/wOLcpIL3K9/qCSmbG3/2Y7SbNcjqoJzE+BAS6ljNLCIA6f
5pnXF3dC4XY2xZLKEwjkDkhONCrQehRA0czX02yzGaWo/JJJT92EDSa/A3U5CnzL
KKBcuDzVCu0QK6d27QF5df0OXLHmfu53Xe2AJuIaMDMlloC3PDLgZBWMXcAmfwRo
70QqLMK9TEyLJWxl7y0oVtGxfT2crz384TpDmzNZWFjbRhrbpOcoIWpb8jTpOuAG
sC1uwD6MLAhjQdYG3zOrxRorYvETeRdfsEQ5fZjqtVbeMvhKWuqx35sH2gch+b7h
pD7OARZD0aueLt7UNt3K9TYSmNO14DnVJg6NbFuwL+Xl6ik5jg/9ATo44HQlMzYl
GAikMBmPzzOoTpYPPrA8bAXLNwX3ewReAZAtpy5X9mgfJhZ77Bc0jiPAbCsHcuYP
wMz65tg0gN/r9A18MTI8eFzqsUVAjV1ikbjtc89up0bpZdO4B96tWtyleljXxpuo
PF4UPQ3ea+Ex0RP7AzcuKfqYxsz56lKelOtUcADXuJck+5WuIF0HQiIEQbjrBV/h
S9jzVsR6Sj+vPQOwJR4VWKvfOIJB8hDugd5fJ/0uo83lYcVpdlXW8lm06G/xfbJd
XZvnBiivHzs3ixxuaTzVmsis98+eIoUdGdDWUVDeADSiT0eGuJj0RxsQgD2StWWa
326U6IN9fYT66XRWZ3tYWDv8zMii/SGI1+xG2BV51OOlTZx0KVeM7H/TsKEkRtSE
1HH1LLtrouc7HnB37Gj1Wf27QCAVrzOvQOHBUcZJ2QUB90TogwtEKu/k1ZUM74Vo
9yEwhjQccCVfY/O8XJoDccpFDxdVA50YIO4T9VP8hy5OiKiV8LQzBX1ShIf9UULh
YExWlrwhtP2xvRtg/P3sLQZGKzTAp2CpJFiZmpuNP4A+I4dFLCTdGJzy3KqI96sk
Lz0HeqWloKbzwF/BrZ7vusXlKXZlf/muJ3QN3kuTxCTmOULz6AzFl8F8baaxT/Qp
xZiJnfgXeGQ4s5a0pBuQhHvPXyKrmFpU2SwkpPlS4qNc56GTGQNYL7eDUlaHk6ey
g1dFbhwtJgN/uPRZHqZ6itfGX4mCf0P/mcebfgEKf+DIsF8SnL7bQCPk+YgZXmhw
cf9ei8+ZaJ+OBqCMSpqrWO9vK19ia/m15jk5DTjj/A4+QRFcOfJ/6Zxm8NdbX3Hv
4NV7vxo+K0KGLaqFsJ7qabvQj6nl099oHjbsgu26hAQizTJtfjacj1jHzOyPML7O
L8ak59MtaIO7sAQPWbnopjh1TdGps2p0mKmx2NYvEs+D6nn3w4CId+dUTWVhkSCM
XvJYA3M6ADc/HhI0C824B51ril2KJIOemEgf9eP1p6Pcprcu6e7w3A4kwQfSQYp6
uO46Xm2msSocFG4cOWdXjkyRmOFZjcPO5+1vXTfE/2qUPa9n/4vt1xt3PRG8zGRI
/7Zf3I2Wwiv8MB3hvENvTJ/2m3dfAdw1VSozernFuk3u7AfzyK24iy47uc2ANhBM
YtzZC8OV9brpajDr4psQErYOvVvsF55xkqpm+zK7biuK00dIRLB0IPHs+coLnuHB
BuQqEpICSVAiubLuD7ZG6sWafUUcy0IXJzAwGN2Lrvo/tfIGm0YTBUt+EGHyiJZI
4Il0IfBpcrPQUYhPPxl3Z5Nzk8upOW/IYzCcgl+dTQ+ZnkpnocwEn9AQoz9fxnUf
nT8cXfACNPNU4YDb0mKfRts1q0VDTQYb0Y9rBB576KAbbfITKRqqVrad1cGiY4O3
sNpGyDItuo75b6gLkcYja16kECyjAUTIOyf0klHAd2GBBtIBQ8UcKAvl42+fhX/n
7F0lni3aJvNruEUREU2l4KyUno7xLfSUQErITBNAjHQU2x7bF8zTSkALIxo2IkEr
BA8MabBgleEdPEMlBRZrZe9aZRpjfzDQb0sgLbzUbNvWkBdJdLDXIWPPoW+3lH0n
jvM5kjkDJv3BXLvt4U6sRjsizxHnR8eHwOnRPExF1Qpz30XAM5TDJ79j6rbulPKE
+Vt97EnnMZ1V5FPiMWutqv+Nd9I4kejjf3SsgauIIcGKEt7RSUlncD+ML6g52zfE
V24P+ykHe8iKwbv8Ia9bnGyEGUMEuk4KTCYsua8qAns8C0MvSaBf97HLR0Vmd0u3
v3Vem8G6HvnN9OfpubvkoVdNlJO1rCErcg4idn2KPUrxai4r8xOjVOyA1dZ0eKYW
6PjZPHuXIDXWJbbqByzZ0bPcRDRLff0Iwkmoy6a+KjeyXKsLgwEHpPSdw5NPvNNw
i6fFOIBtpeEDJNXwZKP9U9ryLi+g4nmgQzX6QhbstOwTBLRpEggUtmH6C63mvN2u
V7eD88suNyUmG1+We/n8R8tD9PMWEvchtAysEA/SR9JZmWx8GEDhrbBbAJfvAoac
U1iT+/Kq2iBw4YtDz2FDAQBwb3zBIz0dE3+O6BZsM8wffsSmkyYY2q6zDWJRMZ2B
qOY1eSPlgE9wZVByWdb4JnZY+RdiLHzY4P7wofk+6m4cuseKD0iJdG34lzo+u9qe
ezVIrgWMYvQpGvr0LNCrHGPbrwW73RSa92GekVrgFY4NLx4SErJnfA/Lbo77hoir
SEzURQy5eEcm6cGjef2nCdbFZiTi2YK35RhVH08Qzm0pmmYR1qE0AF8iqItgoaLR
vnFUhftJhkiQ7Tww0LOuojzUjgwHS40nZuJUSJmumBdnBCQkGchENfbN3FfkrZ/i
mwsAS5PwsIwFDknQwtUHg1662Tw+eGlgbfVCAINt++vxYDijLHFjZZGySDZjhCJN
C1Xlf1IzozmfILwK158mZaf33IqEOmaQQa5+9zKnsKhb/U4sSa/7Zp1Kz/vY7hzx
wKBmF7yF7l0klNgOqBJ8iV4CWiFzH8wkFgpCBKvmZXBz4QbmKusiRjdWWBzxLH1Y
IAmoesh8t+FQlFYkIGxySEYnKkDfKeOSFEPyVaraCfIpPeoc6nF33g//iA9CndLe
a5elUYokK1vEJPNTonapbKUfsS8XS4pvQvEl8mrPTFQyqGF/8mpcGyzz/YnyOujS
3Xlbsia1pE9KfgiAfa9QtjWa2d5mAWx7B0ERhbwT4IDrzPiEueCejcJHOPJ7Ca4m
ZXw6co37pRIf1gVl3+AEdxpiXJfLQ1W7+L4RTezgLMDVhTxe34cUAw7+yPI/1CNP
8T+gDJjhoIS+l0LCLvl5WPdwVkrUX8cENfmssaX58+foiA9wrd7B9CxAMkdMcFFN
UQx9g23ARAcf1XsQxMvHG6H+PrHfjnWcxuW+08/Bb/vWvMqlsce79yDaOIvlcBuw
WAoxB6AL09qJqJ0nhWSqbL+roQe1UPsWqHqbYWyOhS90NN7uw0foQNTEY7mdyBI3
jI1kcOgwcPihD+0rC/Y3jzEoDhhrFpy4V5cBcn2vnWFaOmpKTkfPjl8BzXCh/H+n
JFM4tVvSPmInQ/8w4hn9Zvhr3hW025HqLieTaoXQwepeJ/rpYr2Dm5ZbLRMAZXPg
QSNVeTliTIAj7IqTtC1PGHmDt3lW/EsHECSNUjzdEQ0wFsM6od6/6cUADH+ez9jU
SWGEsSrcpq2eyoKxBoEvxvogJT0MlagC97MrZrEddvCZAcUBR7WeJ9RmGla31yeV
zV+U5a7hTilxg5Cx3L6niHxN63VYTm+c6ieJwjFRIVODIdK7cvsXygPRNJKDr/xU
dHEuMM1Bhk5uO0eBmh65OKyP3AbTTM8BevUSNz3DbwmSZXW10EvsmWTXqReiQUmp
JKmSGEYOnZ+refAoUdRUOHDlocmpbJ9YJxAy/yMj14NoYjDj/+NzozpSbMbq/Gpr
7ZCgCRkoK/+3ljK6RTi78frC1D8e8+8fZ/hnt17ZzRY3E4vzwuo4kJHQGbs0FF6y
Bwvy0j0xQ07jCOrlcnR+SWlepDR9JI/qwKNHj8ixYNF117QDDbxKZGl4iJWIkDbV
1qs5ZT5H99uWkITaAUF5TQIlcYDtsN8JmPtzHBAOdqOBykOg4NOfaXQwWRYrsQuX
pdMLYstZuZpVpXG0ugj3oZA+FARYUzm+dK1T/p63GM/pfxR7wf9pFglXMbtYN2/k
mXZ0ztqwIVx4XEFCD9cyNdVKYmk95wHEiPe0XBopEMFLmWIJVnC+9XVTNgqqJlmu
N78bstWLllbdXMiUx8qNsTKq5capwkS6ETUsDuqwGED0Mr6wRBu1KI40mCO7BYEn
uv+AJS1DoznlF/L6nEFDSRUjMl+lvLnUTOFP69JDgeKsL36p+RmZuIcx2gdap+43
h/6gBApJ4uzsFgM363w7+Bm2jkDfmxQ54JMYMYOoTaKcE/WZNIghsXil3xbWcZBx
FdN67dSfHFkYdMRtjsNdY8W2UHvOPZ3QRXCNtbr3O9xTTsDqAbaVJEfKUoUEc7b1
jQec6cbBWyyAAH7qP8uBG9M0ZcoyGiWofnKtDPbZmYO7WSmpL7fXieCXsejArQtw
z9Qj7oglYKbym8Ujjdj1v38j29RUMBUbU6GiFistfcVu0SP5x8EnpB+QOzem/769
HJhV85+/Q1hzRecgxCSDX3yKBSJbiSob39Ron2Wvc3ws8crJSC+6EQiTJ2fPVWb1
7sxwQ2Jm2cLwmhc8KVbd1iHBh+smOPugkq7WszcrIWgsh7LmuDYqJ+4r1XG3B/Y5
dvWA1vMVNZXUUJmK0kC4jMjjefHkgVBBlPWPOAyJK+qfiUxApVPjR7TX+b5a6Yo3
6lhs2NbPOPRCbQJMNubKjayoR1lT6EGuLnm/j1+kekeJpx8IyXw/Ism+MlBgGn7y
1Ly1QPaBFcSRN/OLnqdEYXCajN8JsBX0+8YYHzf2CtT6SAX/vNDZPzZqaUEOuHVs
+dvcJpm/ABDvUclZeeiizsa4bZEjV0nrgeUJ8u2pKj49KZQPHu4IUHTQkfRsO7QH
oJWCVKAcghe8mE+8XP7VQPl2VDZKfIEewKUH/lcJNucMIB4RtAMJsj4vLrF08AES
q1wcgSaCdGBxxpyEOZsaBmakfwWbZO+VhpE6HhG75v9f+i1tlChnhqn6hQdCVXxY
AXeHM2PJN2/Oxn+5g/1UpgAca9wvhJp4sniNqndomhsgzTyennnUznbPrjka8ouq
hEz6z0gHUOLW4apTfkxrute39EB2x47Gjl/m3tcxiqMOCJU79H89YKCWR96qSR8B
3pveFafPTx0FvT0Js7tEt/Y5jGBaAU8lEbZO7PYkCW3KTG1JdY4k9Gu1RAMVxeCV
pfcXxr5Hi7+9Kzy65wsvcpUZ4sAh+uX8VloggnhcbAh5oF84QJ3M08nW7gCvPTd5
5CJfgVbyDdgFiiq9p0Np/B8hmRgLwvPJRQTODtcevJuPfdnHICyeRgZMlmPUl8RC
jvjOuD+r1IWnpVUK+lphc7X7hVzFvp4n2pDb+J22makRGirEbznQXzOtSJRtSCL0
8P9GFLwBCf8t93YcYEygTB6RG+RrYglGY2gqX1aScUfCVaT0YYaxFkpSkRxMImE2
mzdHDXhM6+ytPUT0uJzLKQPHu1z5ySCuRVfI+NAmrbjZTs0I3MIhVG4/Wj1mRuby
5UU+o9fN7+ecczgenXmc8jmMr/wsFDJpsBFFFni1Bg9vk0dkt3HsBDShgbF/2PNU
CSyZZ4XF6kNYYZR7RtcgSwOHmA04WNDvM4aWB9oC3Um7/yjJGLQj7Q6tjLCnhUT3
IrcI1o9ds/IYIT5NUZ0jWZrIo/CxYPt1T4EhcB+07EVdHEPlzJD9nEiToHUySsDy
GMXQKPWyyRSAdEixm/jub4/w6kIWNzTXWRyIS575G8VI35GW+3SQEUFnSTWlCWO3
CnxMC5qaucsM4uFRFhuntRzXWdx0hRJI/1J9jyxDkq8CRb/Lxuva3oStjo3NqzVU
JyzBKqW6OLm9knaIaEV4vCit8040WoBwJX4jg3pHqs7wZnlTWEdJAqNRMV3uEfDv
hVjFa9ylJyDEf5Bw3xa2zi6hEQp39v+DVGFAuUFv0eMkBcN8gjEa4VTwbIP214gx
G8a2lYs1N+aTnOpm1gFcTNEsdEgcK9RdvH91+Y+/pfcfwMXgY+4P0qXkuHXfwCLK
+4OK/X/D0b3V7Uy31H0R1r7SD8EWaZjGU4G/sqfSmVUx/wK8nW3Ga83hjjkaZq6N
O+re04jcaRaBsAMmXXsVLu28sFkPj0z6VnXnQv9AK4kyiEA/TthGM5qQXSD4ULxt
xdEH8z3nlXHoqVWUxoHdJ3iOmx/hVn4yNq/e0pW2c2iSKpxHT+8ROdFNfiVeN7iV
Wz0C+zHigqHmyDfVB+CoXt1D7ghdVGerHVc2jWB/lZHBLFXZ2SouujxrWeIw/VSn
r8fcBuojTPrBQwaLLt9fL6lWMoBWV5JGTfh+OoA6RVHKpYafWCxkmnRKf7PMtKY0
MJrdhj4pYWB+m0XA9qQ7e5irEtLlNiR2DjqFM+gRny6FhrOTqJdzVB/Fwu6Zvrze
oM9hbd/uegrxkBKzRX7rbXu6a4UX5eEAN2Oia36EEYRwIKsulKzvZsJJWYBRBsJe
IOZ0DPcDjyp9XD265EyeFcb/e3XhvdT4Ofnrm+UCKOCr9i9ZT4iwz2fvQHHp7Ya2
lhEYaWyyQRZXCjoWbq5Y07Fg1fx6NMuH5s/A700Fxd2v1A0Pel+64jlU96RelP16
s/DUYJdGLXw7bCCRSTIm8VpFCcCl+DGa8MSGe+a29FQ1KdpjXbxAD8jUA9fog3TX
aOSf5frnCaH/cqZSZih+b0ntoVAQrEupwVzNlgOyljKv+biTd8V3JAQQmJdi2wT5
ilvMp6TsRPlLCyTvv8mT3MEBIq1TMevivjxPhtoLR8LyzkaWJer0IJQZIc1EM/uZ
MMKmXKl0clTHy0B/iGLQaz3b/H7+rPbodYhUlsZum6kHtiWeKH3p1jsPDg3J+Vd0
50vhv6L9RWD4EKOA+JIxo0GvZhQxZZs+QCuaPks4g+JeqWXqzxuZNJr3Vx6FOlSy
iYqSA/di1hKNcdEb2yNs/YO9H5HgSmP2cbTC88o11blKY4cC9B+IctySRW18xdlm
8+Urn1BaKpOkI1aceCThJAUBpHQwA68imwkUw1XQ74Dtr3Xtv49dzB9uWd5H9Pro
9r3jn+VrwyXSDVXni7BJrkCtMw4Gpu1GLRTnJAu1lMYLpVsJ5WRf+hA5ScZ6uQYm
1+YB9Mn3ckvO8mqv99B68kUjW4CyVhoKcIB/bfIc8lvLwKml/7ywWFPYhvaNDC4t
qMQuHl0H5Zhc6thOhTvwy4ZCDLnUND7B1FPSZ3S962C2dKUkKDnKtHnv55mRc7Nm
VmK+pvRjt1NKJiEoY2pXXFlBYYzSXM3aN91GHEAFSNk4Ll4TFOoQAgPt8ZMyX4bd
QrymeeDAnpqSSgqN/x+Axdv8c6xD3OAbWsjCOHI0OOsvrRJvFkCgGKr2d54E+pGv
d4foqJ/CX2PIFhlQUuxgjgIIQjUR9nONjWLiDKRbb7bmF2tP9ZPASlE7Yjz2/UHB
HuIX1sy/gZg9XOw3hoqUxLnv5Ndr/NXJPXXciST1zUkl+ekVD8wYCv19iwffvZzB
K44wr2Ij46HTwJdM5Uu1rgNIzSHWv9MTM30hzVShu3OfmjLe5nlMmySxMz5ZGuN7
u9Z+pPZwKZ47GT2HDRSYr4V9mFaUsi2y7IdBlRbHsnLnHHvOzIRCI7BIAUDDPoVI
bXgH6F/Ka9THFDsBYXn47iCbEudd8wFu1u1z+vFKqOhUuc2kRrKVC9YoIpdQm7LI
TOXbfwGN40WwThXDXiNOaJhsr7sBhlfwtB9Tl4tKTtUyBwjmm2Kk67eIAEWVZFR7
IGlkyYgFsXB4ke8pFnzcDSjPpma3oZUVDpGBIZsdV2izu3cxixIm8b5/xk/b+oxT
21qjL+GiT6qUgEVoVDe34N8Ru1TRIdRJonDpHw9m+YVt/wHmtIEols9fMXjReYmo
MnlJroDWgDVRoXk7pJeDIndmsnDnTz3pcGZ5JX4v16ebC61XyYd/cojnJ8ddXL+d
6nS635ytBczwclp5lRgQJy/KhXIjd28sjsRuEQWRY81xHCiU0nmFfLxwpYI2u/8H
h0NWPzxFgb88vIMBW63IUcjK+S8v1EPulCjKV71Y5dX5WS1vQcb3Qu5RebpSKKIe
pcgWPms+r4Nz/y6qgZ+e6FzMQrpo37EqFZwwMwRvf65qO65zA7f1qtLBXPChWUx7
BxLanPF7zQ+VhHoB0aXxPgh1x2rXRSm58KlH8TBYIZrXsKSoXedIUhaoReOtn+3E
K3xh/1JtXQpd2QO+cJS+YnsVgFfktxF+hpcSnfD7gjBo0+33YGV2MnXdvBpjf2k1
NraqMEpEKRU6SRe60CbjGXPJ62tM1LuI8Z3qCeJwVkzrHPuC5WbC9R0ctlg1dUVx
l2Z8agQc++pi9keUIQQbdrcCG2TaXbSEiqZTlyFU61Cjw+s776dVAhoADReNkeIK
sb1/Il4kuxq55SY0mskgGkZ+3HmPjq31GtwADLZjfDDzB0C69z/lCLXphf0I407G
9aT8U8jVLdu6kQe4D/TwVgVqJYpmEa0RyfDQqfiZpq+JRl014bIzcWsN+e0zFr/h
4dFAjXHTXUdqNiR+3ISLHnIJ3cOhtqjnA8/GwfwQgenpOyLR1VBJOAIXo+YfOWas
pbt3KSSSyP4lf22lvar+DZ3dB/5+ZxejkhP+DM2tVMZAY8rRyESmj93Y8euBsIo2
xVSidSPa+ZVuiSKCKBRUIefT5ZVnZtTqWUCIo8WW7N7aopRmayfwsR/yl5/Qqt9X
azilGMXsAthgq+RC+9Ob96jYhszBb7gplfU/27gJlCP9hjXKn0vbWsSN44cA05tr
bq14iE+1d4MB74wZk1SD0d9PcOXWEbxdNbiqVoh2Gel6rGJGaUuT7rYjHGw1M8MU
5VxJlxVZHZrMzXILDNK8OlxDt4xjFBCOlJbb1oFWkPKVUuyC73reTh0NTR4t5ddE
3WZS+tIquwd+/4axoHw4mAFE1tqjL+G5neVU+HaiqIf5E7yEVIxWc7QUV2by4yxP
778IlY2V8FIAFixO5tLraAsM+kk4SmilOBY8yp4lxzPWkIGX0ZiTKPhszv0Odxuk
3R0MG8XWyEmtjwPhrYZ95dFKnh95f/CKOiRqHiC5GdJkZgXh30/3Fr7T/8n+MgEb
uGYIWBz0bWL6uuuOo9Pq5DN2VdihFPAbZDaQj0OmI8Y2qjpekiVqDrrq1PLiupBi
u+miJdWv8v7zzqbLujbERQxACCJ+T/qf4hFTy/XgcZ/ayvvEI0w5sObvbepbAOH6
UwggZitR5aohLeYpWlQNleytUubQ7uuFCZsGIaaXxqmVAaGovr+YwqIeiEa9tK5Q
VhtAbX6y6LVPKJvLWjpseTf5qaki7RUe8qx2aX/+hHRZVXfleWmFZXpLZ3suTyv+
WAuJFpQOVB7C2jnSDQMK006grYRAHT8e8Yf93IRiPxGAyOQdCWd0sNW/oGfPQYN6
yDtPh5y2oca9gRR8ZSIEHIC+D5t9cSbYOh2KHe82fYt4T/+4djO3FNmuTZGCH9bX
JbbqlGusnP9j/pdYQ/nYWoNjIe3OFweyQSIbfk8REDwjKITEZ6pBVgm3Jjs7pWTk
W6qcIHEJJ+buF+xgicyQ7knAt96c1kMQkdfqLNjuyJvgguuP6sdw50JPRM1SJtZA
28JEj+0mR2wNTtUZ7OMoykwgdjyTSqe+XaTK5o7SKzsrgewEv+BvTxsnpXA2fD0L
vNRxujWHs73uPa7MGhfCa+EqpmxAvuuKE9pi6/G/JRA/eBc2bSADWzxfcuH56kWF
CbWi+BB5mZ7noWCBVq5LjqVMD5xdfnC6fXbNZaOXkwxmBtebSsXa4RWU89aHj2lU
Xh4aYxYyYBHgxDvZvcpqmpe0PxGnQ+P2bsFR0VBIKY7cmPfZnIbODcePFIStCAUb
q4TmESxHNtxhg4PLxNsvaAObPlpiQ8hzWkREVAwOxmv9b2pwEKDjisqXtHF6JVuY
IuA0O3JKoAFFmaLpFy/x4H/Nugg2M7xOWX/J+ErdB/4RXylNCCKy5vGj+dogC9nm
QMLp69HYG1HnMyyX2Rbq34Yon8s2irJCRPjpk3AUvPw52MUo1XyHsrdX/HE+AYxY
q+3O1Ue490YK5aSoN4u3XO8ogZOdEEub+MnFH1DHcC0G6zMgl83Q3t264h32UlKo
zZR10Y7+vKbKtN6zYMzrg5RSpDSCbf7FONWKvc86mgnHyVf2qz47jDyt6IISTpos
S38lrp4YHZv0IqWiBIJq2SbIXfq7kelzKe7Ouc7zALrsAa9/bYv6NavxF1z10DcY
3rjXarptkKSy9STClbpUMSo53N7x6U0O2ZlHluveh1r1fVdVHywSrX67e+K7nQ9A
pzChVE43pHzBDe4VeJ+cAJIiSoJyPV0rHC/eAkkojJ8s9bR73l00czFZg9grZJNG
jy2UJQb9WaAYA3UOfTl95ysYn0x78HT6rNYlQI+JQ+ZatH/cWlOm9SrIRN7qqIhy
TrGdhZmgX+Oj9ZBI7yb/pNXIjQAIOST2UAFsU/iG5GQc1oV2mhZddg3xI+UmYTdg
DPyNjEGmpbJjvh7Zz/Q8+GD5BrHNBZdbmYbp5vbENc+to+swxABOtr7HOFQVJwD4
oF0rKnDyvBmrw74bPSdMB+VugozPJTnEoRzPL0+Dn2ql7l2FAm/Q8JsCo2PgC7yK
Y0a8vVGYCFj6lmRVnqPoE80zB8H61adE9Ho/PejsXlBSYh4ENQWFhCCzmZMzgix2
oD1nM1IYU4Peq/4SEwdyLnnHe9G7D4UJx2vv9ewvLQLScU1dzftww/ZPMbTitU7s
qYcVlAaQzh6WjaGaJKYtn71IZ5a2vulIbg83rGje3LOlFC3BuIc3U/GjrW0vhiad
/2tej+e9W2OecnEb0RVZP2QUAbYlkIW6MGqREY68HlG2L6+Rg8YKfc2QXGRP4kpO
MG5Bo4UzG2/juhvvlpzRpznQKRMytAH0XKj94QStahBRtnINqS8boEsgySRNIo6J
LBf2ZRLC0Maj5cJAAyv8A8dSNGEB0/HtroU8HPKqBLNswTD09wOigS+8lGBV6zeh
ql0EldHpv4PU4Ut0cEoBoEB4kkFg+bHePT6eDMnGL88OKl+l7ja3Mw0ubdbjVjFq
OcuShkL7fVEbHWFuSRtKiP9vzLOjZ/uqyxYLjyWrXB6x2DaD9dyIaB47gVr/+3p5
RxB4PlcFGlp39j+IoCDr/thPK5GpYz5FAiVqy8iZaU0a+mxGNrWj0OzcdcHo4KYr
91Ftrxvjp50ryrcVsq2zdJEam/YA2iSDs/rKxF6Ov6Wp0yiwffkqOETXdOFbptoB
4duAy7FYbqtbk/+s1MCfl9+V1hcHT6vmS08GuRCEcCBbykXLqafrowMfH6nRCte1
mN4gwfc0YK5kYUzaWQ6Vuj27DnXoOAoUTxcCFh43JCYi8U44qN0VYddVrymcsbI8
ZmJAdK7iefrjsAIHV40b9ts5v7T04+fYmtTZRFQQfmcfY6d5MFLNgLynXB2vJRP5
MsEMBc91xCRfF4RVJ0iCwcGZEQEFad1bR2YoQz8Y0oeQRIaUm1JXw/pALsfvPbXq
tCfo8TfmMLKIjhd0kzjFivw/vjF5gnxHK+Af0pNGhS6SKLx5pWacIfasVK6ShyHV
FGY19/LEBuht/Mo/x7GfbmNzgVRKIlE/zpk+xQQoLHVYRuP6j4Muwc4z/i3bOQx6
Da6DjxZZj+jIqGg4gytrySjAhOkeaY334Fbpyc3ZOnbGxy3Dne6bpKUueHOqrlrr
uJkhDsR88650EBwoEWWiu015tuZdTeoQTGRmuZ7SEZ/QzgB43OtueLV4G1qTBGjW
D+W3z+CB8gZPxMLtn6RRTRdSVWzfebYVCNC4jWd1femg4AD1rRmY1STL3S9mOpwN
aKFakWrMYLP/PAELvjD76H7LMCJyW7+IbsZjWjvkMI7cl++Xz5c7GVF90uLY3JtS
6ENfltdYttHnbiOi9IVPGauYSA+GIZnL5LetnFDrFqymlFKA20I/lZaX6ZysjZl7
7TXvH0iReyif0+OsafWVLW9JXyScpnGt40u+ZNDBCZ6y0zlXy8/nAjG/VwOL2Lfy
FlDEaRlqfFZJT9vTkwW158IGqICOgBPH0Y6yxppd7HYrDJ3r4B4x4hPxB+JFjKlo
8atqhN6pJ1Jpw7gh1B/b51JcjjkOhxT6NkWeYe3X0ilVUNvpvI2vdfvddS4siSf7
ufJ2OOc1TToT2rqUP2zyWcFJn7AyZrKLCdJFvWH9qJ5HkaxllaJXeqUIzOu8rtD9
x/8V7hZzDt/liN4nzyg3wppN95DhhteI4uS79Hr7Kow3+BO/Z3eCwAiHdEUnz7yz
CBMRPCHAuS4VT8SpkkKrR3dRiIpwYWFMoyOoaT2KJdMaX7F3imlVGrvSz2jkF+5v
Y6SKCoL7PQ1RtL2jPkPelfqjMAviDBYSt+ul2+3wTqnCoEND+FwjdyUQ4Xo7dH48
lf2HTBHuyx6N3K2YfJuvDtCv6OaT5IIRYKgOncyz9T/8/vu8+4eKPD0fOLnR9ePW
fhjVNhBH3keGIslhpekzk/VXpmd/dwKyk2iWmw2exgoYaA3uodW8LmJuDeyoQyEo
X7Mg5ps20xeioDbUU4amjGVDTzpAIyHQC8E2Xe2EFozVrLXCF/MxZCj3i7pGDPso
kof3bdiN4TXuTsXsq0A4lAk0ydP6ZSN63l9++2HcSvrOCpWfJBe9Pf8mWxahWry3
n0lSBDaoOXV9y/7E1/RPs6zmWGnTOruqNSWRJsdpmNXTw3UOzM7cOQ9ck1iRgsXH
vvSPOilI9/XAYyYeX12XiTwzGg5WOMGaT8AV5mwAUpAykzZq5WxmFreM9pqmCW4L
Tx3uT+9NzIomuizjA0CC3GUYwTSn7aRtPnlZZdMAMWxeZTpQAPXgpimvl35rijcY
tcojkrdd2EfyLqX6KCpBI8asLDm1UTe42uAMN70klW7uC0Huc6pFN/PQTYviErnX
yvuhGUWJ28tQG9Qhl0sG25zKiF/QF0GZlyPojEnysnqKHW1Bo2Loq4q+qmz9d0QO
neEVcXmVNnSlJ6w3RDD/cjeKiSDTTRQZSkZk3fvTcuXfxElCEgjq5JabwGgc+G57
GBAzRws2iEs2Wa0PifxE3g2uIrEgsM0RCFRMsQ7rtjtWoIm7G4Ha7H6dftUw1YwN
b6pLhu/hb9rinteBmR5e00KPqRizYSnsv+IUPbtTxVmbV8XFZ/b5H0S9HWdXCyFx
nYXasRMpSE6JYm6awwMmAhnHw3UwOzQAzqp1wVDdYWSF/r9sVLPrYKD/l7tsTfVy
b0UKrRFoAPf0x80ez/Cf3ffjJ5Ftt2ZsWWd16gF/dT/ktyt+J/1mbZYm8iC+DQw+
3HivO1PFXJWaGIWDKDvSHa8WRxort0sIP1o9PnL18PRgKSWPo8QbmXI3RY3gAbTE
ZoPDhUL1Ff/48zrWcS9Ou66Bc8zsKeqpI93h/SeNyH0g7aCAsEyQINuwAIhvp5Rx
fKBXJdW8LfkoKMe7q/cQf6ZbZmM5jHA+fOm4ZqcIV2OWeT2eSV54yr1cYFPrHM7n
GktON0p+cWAihXM1MBATi+PmBQmX+XSKX5rLH58IG6t+3xGkecXVpcE1zKLSejYC
iAojti2oPuUxHA0Rr+55KhaSysFW120hQbvJ3PimXSz/JNRoxdcQ+8LIDS2v/hVs
16q/ogrxBWQePnzss+NLmhpx2z0AJb2qXSzJwdGl0rTe35gYxWbVNdhzQNVsRcce
0t4i3n3Wzh1wz17QY4bf/3EOjlsdPZHEBL5kgiCcTWv+IkazWxtTADU4McJEUPu0
lUyq1nhfkDgq8q27YE0lRwwgtZjEMLjrLbPWamCm2NswWfdiuRUsFw3Ka3kiQBQJ
SCMTP/nrzKT38bPu7HNWmrEBlZhfX5sNCwj+Dp/71fPkPyhL7p/+bFqj7+wI+UvQ
x8n0RFCzC4+Aa0Dptmg1MVEd0O96Vr5QTrBVYc3RciNPRuvVi8CAxLviwl50yK4g
lMj5XiDHiQ80q88gTlmm/vF6PJJHmAcvXnkUiNbgM4BswJIVLnkigLOc3XpDiSnn
g4BrM0eslIJ5q2VPyVI7nD655WkM1wyXonzIjf83r50HzlXZg3tTNEERW1uf9PxJ
/O7IqDHz/yEOnH69cvDFrLkjUnsfGPRbZQl3CruKVDOeTNmeJYCtmDTtklMXtzs3
oUV5oedpibG70l1TAAvkBkhXt9n11xgxLbOP249hYOHVfBTPSw/ryLnGQDL8hXYT
X0/KvWwM3C0ncZ7j4sQSKXDtXWqEMHcw+6Sn7Nv0/m5I/rHhfbFq3xjmilMHrDcC
/wcnwq4zcmAF+7bChjS+M8g8BEJ/xuTPQCom5aBjgPO2lPCGotJ2WRINxY1CTnIq
URWGyOQz8W+8mJixPnwB+ZQaKX3BX1+IuNBcFXbYm3FT7K/TsTcbqfwwxXP1W1sI
tM5k4ZUuzftQb47F+sc8/5PBGj/pPFB2PtbRItCn1XAz6cvJBt396ppvO8Sh7LEG
zuA41MhH+u9xMGdt+tR+EcmLJuhCXcuQi0b1l1e0IKmRhUMJniuJxU437ftBMVI2
i1nHpLc3Hd5fOK6/POLv5Vn9xy0iWZLGhjHsZ27zRTksoDRYFvrWkFRsjiP5ahvR
7dgrgJmHEJ7TVD62x2QweReZ87B4sE7pHCYLDzWtUXpBBZbkbc+WUhtli/USLiwn
gvPlUl65oElr3+6o843NTIg0PpXIpjoZllvPmiJz4AWToSYmP75jpHgHzPCkOvGS
U+fQaSZz7LD6K2acnsYKClISvFa0lc4xgimQMrIx/VX2LIp/NgR0UeVwRL2k9fR7
kDAAruL5oiGc7QCyCoKqjcHT3NBNx+uBfdDctw2qTafUsogjwOqYbWUvburSW4O8
TlJstkj0QH2gOxl7Xn2GKR49MOySW+itSZFsS3+qutgwZjaOXu4Vhe1U6Lo5+gBv
KoHlUMyRyR68y1ODTiI7chajDwpnhPMzoOj7lJu3kjM6RvtTdGmXa5ovCJwCk+2G
+efxfkl70sv8/KhPtjn6gX1PmZah+I8bb162ro/T42oA1mqFT3DrDYZsXC/Ubu07
Fmqs48AKpnWQIqiqBcmE7rnameBtMxi5pJVxv7jMAdX7gnQsT+rlJ0VmmbaSfa9z
iL89YrI/BHrMfgGO7/9yvPkE70Qqc6o3cHyb03ZcVgfbTKIf1XFdJwZ+3zkVk8Jh
qjI3dMc8bU8xsKjiAPkzVwYb9OgijIEPhLJc7zrpgvzvtwowyiquzLIH481nAdB7
W7NZzWp40P6qk3mAbRhKqM8rry963tQ27+Fgyr8HQghGA8hBWDwJmnBxbHwziZUH
K9zF8UW/njU6qQc3Nmn4/hxTvmXkKPjqxXLCKB96AuPCqdkkGDnG8zO5cZGXEwoW
knWLS1g379VZnv/Tk2hWi8UlIuzmD6SwpI3r/UAZbrvRpF6gxxuZ/ydOVCgjYXGZ
+P2UFm0GXxlrRs0aSkcR1j0/iybp9l7RzSXZds64TJCNPPoN3kEN6j0VBZNwop6c
BYydQdzL6k/njq0R9DAadLBvutp8ag0GazXO1qzrs8C1ZzPu+09a2r2HoLI+TcIq
tWeJp5NognDn2aDhKfOgnTrm9nKMsiG9TJVgnc+pt7dS7J8JauYW0qftnc3+tzm/
J/MsNumC7Vv8EWyoROtASoKfaEg6FJuYcIUAAH/QlLYBXW6sj8XLayyxwlqVZsxJ
XcSFF58W19PPy/+4saiUs4RhH0teQZM0lo3SauBIodtAuQQ+5q6tjhgWtbFst6yO
b2NvMo01D687pzypFlMkbVcDMwM51xSfG2uJ/m4QHB3c9PZk7nkklzVoEF1CN9Wo
FTgnqg6xuwLAPNSx6IyIeRAjEM6WwjoLuP8R6E98tn3KaAb9l0FhWBTWxwPxfD4r
u6l++9nPU1qHoTyzumGBZNGde+F6vEFJCeuZvwNKkVk7ELDBUXWp1GdG10anlssu
M3wkxBRpq33tNiMxiWePB2PXCa4dma3jXafaUYP1IfT7HXcGmjco9qjjw34IhD8w
qbVOHPb80kwP9YH1VtcloSDrIVzztJjGB22wWStCMX2D2vMvlpypHbzQC/3iRwhH
gyCaG76XS7GH8+S4kqf57CKfCUwPw3pjS7QDSbjdPXGB30TXfZ759Rq5IwXUZWOV
+vtLXkboklLjV03FhmqSTS7HM+V+wrhd8uWkV1jVGjmrsx60FLYxzp5noO2mrKIm
FXyJC94dbhmNBIuoAmV61/u+co/nb308x9W5Ql6+MyadBJDBrgDJpTuo+LJhQoFO
AsRJDwJuOJq/63iTxvFQdSpDXsEjxeAY++OxBkrBa6Mx4rkOFTotOFNfJxo0KW3r
uU/pohn43sM2S5uz1YFj/A/c1CRo9kgXjP/uy9fYMiH8poLdL0HHlObcM3hzhU3n
txiczT9jrUqjLqsdwMMOtB0jTSoGFeFytbIXmBxJoGxfETk3k9a0AzNMpKD+p7gE
0ClJHy0dGLFKqcvdb8atD7OWeap1UyQf1h4AsF0XAWANqlZta7zbjrrZAS2++oIx
KPOmBgEbgKVLtwkc6QkMNpjcBlBNyz/V1hSx7bhIlFeUTnBTjpoQHy9muOp9I/vX
YgnOLRVM5JPF6JcpxphehWqIbICRU5VzM9PfwYx704H9bl+rOvneOLBsNi+3PF37
W+cuV5f3rbinjvmSBSmdEEBgvpLfPnK6im9tXFP3rvRjdEWF2EGqnvuuKyxoH/TQ
W5fq5eswnQjKNsElqvXwtNQIv/z+CelBwVMZPlhjfRMSf4RC1LNhRj/O4JoYcWY6
t8ixZ6Qw5vJR9hGJ1E8eiHYS0qFgeRqcbu5CTeAYIEZs8eGlR2i6f6qkx2fiotmG
Fp22wMfORKxqkzAbfaxmnfIji8hqaI4xXStlFxR1wvdP/0rIc5jNKrHhTRcmJhYi
fw5QtoVusP/R/RehfibmdGuPEG+5pTcoY5OZjxhzwZnNHGrB98bFDx5EACSEvWNU
/gUCcvTEWu4J1YlxiYvcw6+jmTDeeLZQZ566cnHMVslzyRj4o0RVlG5lvP8jlkD/
oXNc3U47HmI3mD/cm6csXHyTGOKsOM096GMpwYkIW/wzriAOJkddH2gLDG2Qzii0
SDzCoNTv6bpvQ6fKPEoKy8Iofainj0bpIZNOn12QLoaUTisv6kT+p4ErFQTcen7r
8/+uhE0NuWGmu4Ez87YFq+YNcZtjDMYullbOOIwmBxM6Lz67aoeX7NleVnkv79EN
h/gPInbQk3yWFKs0L6WmMkfo8duTWTVFckHFhqA2aCRvzqD+UxQBITUMvw08pdXO
nXPX7AONxFQxnXgYR4X3cElkoBkVFLSMvkcZ9f6/qjORsHjasFqobcSUS2Si7eMe
qdqe5j8NaG8DFmnCO62/8G9YxNeC0IgUgYjHjU1QK9lIsKDFh5HVZti0Ni0tbB6T
A90Tjr+nf0UKj6Qb7OVHgqZ4asaTR+2dIAqtVSPdLiifICYqH6oJXUdhb/fxkoBL
hFXYYw6aRNCQ8sT6I7ronUznllGQBReil1TOMpmn2jKbzMovyCA0fjdTOuVHubDa
hj1VYvZLDivxFqFoUr/3kQ0sOTdNyxlhump8Eb/a2JEV1PjzenLODXI02r9LOQU8
siTgscEg10Mme5htKwlrIpe9vebz+KFgRJ/5WeYnXnaAE48tZym8jMn/hYqDhqPh
OD0xD1Qivh8QnNPVW8M8M4dK5lpmzJqPxSHUAkGGRFUzVfWUZ2u9w2/Z5xiWkpZY
j8RPzDEl31OVxwu9BdG/OEwK6/4EVN1Y3g4H2bSMvvBmJxWAue/RaVwm4NiGSw/a
oCOdVRQcs5+AXAHDA8GOHfpnYOGk4MuP0TG6gGsNqVsLyGG+SJNie4wtKmTjTW3z
T3XcnZjvO+V9QKfzD7JQDl/oz5aqC2cEinQFbof15wBOozhmMkl3tagp4z+QOLtC
osIHoFHdc0nmgYCRPiiort5AIpkCjgzOCBx8RBUuSdDWXNskjyKe3oPKYNUFie2R
bFHGGc6+JxOHx3w0MjV6dmldKSl8m/WhnhniRciZMQ5e8HX/O6159f1oMU3J+rAj
RSp8lXZK0Z1WtEW4Dw5OJVZj7vojda4+yddCVNKB8EachaILwh3x+wQ7wS+lZdWV
MnKvxhhTJqry9ELQxwNFVmpuk0yt5mrSqNFik5OVZ7wl4iEuEoOrelnPnvsELzqY
SxnDIDk246Nu8NKbLAbuPwnbsMgqbdnYBGb7OcSknuyyOh6vo+KPh6dmjc87WrG1
nhoiP5KJeD9a5+kF7adYiY0R0jjU568EXTPTCB+KFcKf7d+dqoTb1sx22NgpU4o0
JpgTe2KeSWJy+PTygOtCkd3teRxshdHeatPfg0TK6N5OUCGh9Vv0K2J/LGNKpzm3
Eh/HI609yEBMe1WHrEajdWB3BO2O0cEflhzcdrAIysFPMZPGFyBJUbsISJcoRUH6
e9cCIVgR+vvUzyUOtlvTmX/5QcrmHy+RGYOgRXTRlOIn3RDs9OLWekX+7xM+fDzw
C80La/SIsXZULFi5uaY2YcN7wljr5r3dEZicKVo9FNWR3ORcjugcDYzmio3gSftc
VQjNnHIysISOk734AfTIix47ln8ZfsJOPYTK2pTU03xbF9+acPshtbTCKXFPB9I9
Vm2Lr/JthoXuD1ldVVb/m2gFx5CCa9D/sSgo1MRL0E3dkrefcZxewoocTh1H9eXr
3N4DxYKFzBQ2vMT5ov9ZBqbTQdVsB4n4HSQttjmQ1lw+/tBVNfJlQ7/F+CY1Jv6P
HK9Hsx+Ihuu35XdVQP6yraAXdySGoowpxe39Ajn6fZrjzQ5Ph4LEba1g9Cddovcx
4en5d/rhS/TZoGnXq7rwzPvGXttuRLIca1al0OcaMO0d+2nn2ly2tUsEtF82zgW+
Hx8X4sL1Bad1sbwnvEhDcHMqNhHGqiNwmOpqldaAOp1whHAXX4fr7fevDwl/ltwd
zBU7INHOeBk4Xq0xmfj4kikHjI5jrGbU1LY8Q67XJSitHXkHY3DsnZNCG9qFoOdr
MfbNTAuATpDG7mSO0saqg0UN0sclnTZhM1ZN+AO48nWhpXtjolEwcGE2EkOQbev/
uXblkH5cT+ADpnYFV88FPXcBgq7i2SqYg08/ejyLzNM/204OBioRsBhJZz5/ASXz
SDIZwKEXeB91WNA47BJC/TYemBclFIhytqp+AOndqnhBtCxepEkH5vz8NX+YX0Qo
qx2CKOWf2P8cXn/cxXtUBdCEPVL/q12WigG9ICgdWX+VpjoD0i0mRTrznd3gPmT+
aAzfXZ5rKehigRCnrk4jk70viD/DMruZksiEcm3gSRgM4HztDaoDesavWyYa3UJF
QmnitwQd2FhekxU3jBQUAuQxSrEGpD/yfoGC//u3l/5TMDKNvQ9xFR4C6sxyuF22
42TbG2vRaDoH5IXCWbo/sCgC1fndRdZb/pyDQgNa42qwLTROCCvVGjh95EEi9fmF
JThXtE12x4jXCf6g3HpOItZf6wZZCgnffxsMd+ZB8Qt6tEDvg26YlkU+66nDEOVX
/MulPn+XHr23jksWam/e+Le/BveyDIjV0cCbv53HJGVBb160FetMdLXhaFK38OWE
2MwRM1HUxglL4TStSGVyj9tK6B9Rdqi6pP48SBEvM+ts6+BMNYjG653RE24oeTGP
58tPwIEweT3/BNOKFZZhxilVUO1Up1Ug5mO4QzKH1Z5yO82fokiXPMinwrXkpWrd
7Zu39WBveKd4sSi/jqDbrU56MZPeZEYG4OAsLK6CoEtGURVZugYkqaNE3kb2DsnI
msh4HW5BD42yKdpYzM72KA8EUpFNcVPN1EPzRMGF0G8Cuxu6fY5RA51WOZgfC8J1
T+V5sl19MyuXJeWdDXCho7OxCHEri8jdco2JTW8ja5r4V/t9t4l35QKilBvj63Mt
nH3XdIThVScOcePvWNRHMWbR0TWZQe7FHCpQebQ+luPujCABGg40KnNpe+A1Ex5M
JcWeCk1L1a43nHLgfpqczFJjwcTfX/JXwzmUE37B28XyjJbil0NqC1WvnwgQ3o0r
vkpAEoeh59bhzg0fRjwUHTv0e45SFKvv4jyaWLDVei1czxixiZnabtZMuPGySbD/
ZkMY3TO3qkABgpOtBV6bYzyd2ArvVM5rE04KvXBhv4Ax2d8z2j48vfI9JmQYjkhB
zY6sAkA9V+jPf8Czde8VDwt6JJ5vQVYWK/yYlolylIeUL50MS2fErqFiLhAs0xbv
o9Nw9TSS90au3joyJ0jNhcDq6bGrqfainpMVCZImC7IPl+4KvBzDDOGvp7ffiZkg
RaJPAo+JG5e/UNnA/xHxRFCWjBmXRL71ZaHDo4xYlk78CZXx9NqsJ2GbM9FeA5Pl
tc8cld7XvBBRQg6jQg/SlBBVyMBWRj9EACeTWvs11hxmYnnkfcz51w69DzNiD5Wv
u3vbBjlEaOQ8E0S3Mi4N9fs0ACeXq+KGK6wArqhRynWSnig/W8c0Zbp05dA2muV1
5q9bUcVTfUTzLA93/ipkOqrZ2vyQ2jzig7jJOzl6KcR+1uc7ZwN2vewo6FX+to80
/ujqmHM2eRvDZ/Rmip+WzVtAg62ktQKHkkMZ5TxPITbb54af8LPtJ26RTS0G5lUC
vSrlla3CNiR6WbGki7m+z+owKIX48TsDMBJHAcxeIHJ+obEH7/24HI/EIYcrnX6m
SrTxx14dc5ri+7EhWz169XoBAGdasGoTpyjtOIE3UCiviC+AIUzfpTQ7L0ErwxYC
+qAWBZ/B+riAdGzRFia/+rbRztvapEMt0vID+rC/AhNYQLRwGeXoYEdPnQNkGpT4
Fl42QcQ8FCirXxuivJQT1lmMm3Wcp1zuzck2tiy0DUuYw7TyorWdt0QUHDwxgRjH
c+SK5K1J8X/KfCvi70zcQa97I19CoomjqeUGjPoTwlbVSNe5BqV4lgnWZkXgkvwt
SDK3ZH0mZEmYNItJ9AxXoko6w0wDv1WCDY8F084XXaVXLrMRw0LW/4daieyL/Dnp
S8AD5LYDUUHABt0941DMHA/GvXH/HjhxhinwfAR1Qe6UjAK0S7XKZh2MYuz0wMZp
4W7k5OYDduhEShCHAFWooBsSmXT+RoqkwkGlEAlgvHWx8OsrGgC+J8q6Oq0PzFEg
t4F4Z5OZGE9kKIOYQYme7iHKqz8p/zSWWk+hnVzdw7xwDuZ5GqqGWfvSd6qZ2Iep
E9edcydxddnvPuhEivgTEdZPggO7kPEywpV02ULgA296imhgRhuIb2rNJ8IRTB2z
iAbYxdOZhUQet8Iaz5yhfy5fm4/PR0Tfc1t3N+/+k9/A589sxEvuR0DeU/TL56IE
gbFXk/wAbGRTRzjGiLJz5iDC62op+n60uO0IlLaJCiayP0MdVSjNZRrmawwt11QP
gz/Si6S0gKPQ5hIKMGa5wVojqpBxZM0nOyxhvdRMVLbNyljimnlb1bcQtiH1Gn/l
imV/fkEgdeklFLEfPvk/C41HWwDpHP8lG/AoW6xSHegBjS000SMVwry7UerjsEro
TuH6egHBZdvjQLq+Us8RD+pDQlzWhJBMDQmLSUlwY2sBXRSAviJhGbyefMovODQM
eEwIjwlkP3brDuilo7Dya4rYpG75sJhnipPMXa9duGlIlLCqXGWNrWgEzDsf6Xld
3CRcikiuV52joCruoLjjMB8CvZHJWmq4twdZIwlyEYyY1v93Gjma1MWP/stmQt36
EAS+QZkOT9tJg+4/ku8+7hXSdm4LjCIuAC1yQd1TPWjJEF4AsAwTlkhXLwdmnRkS
65tmpuooAdvqVOvEfhCcE2Ca0/mnAzorbfAouWvyG5CCO8+ZEnyv95bMlGf0vBBU
/kTAJpXT0cnD2ufvOIkfAWLgzOgEbFhFWDUEgSCWcNPaBPImXwtg4vWAoJ86j3KF
fPZwScvDsLmEPG9V7OqygfF3Q0uzVA4iWH0W+1m2f9DiSJUynXN6AICTrQNaXRXc
1VGXDqllepzYl6IRLzevmV2VMCNK3jIZy+e6stCsJqG0/a35AdvcMNvGq4JwyQAp
dKniF3V+XrgqrZ/4RXrkEjjLRYlpIPoqBdSRbr7EKr4AYF53ARTjAOPFfIKq1CsA
oRKH9xODIGghsEpSLfHdOXyVSVqmMrShsoAHP/2vcI9kiATFFQI2YtlCNHmhx4bs
48OpMfOcleozjhNd7+l8KwNzrVCQxLQdH30xgfmrzJTu5yZjUBiFeGlO2zYgY23s
FIXR6tjhuEt6Z5jQCQxBzHTd/VElvaPwD0WDgplnEAY8YbMduFutTlx0frdvaQYD
r3LWH5Q5sfmjx5DuwXnPKl1OMvh44vdQm9MLJcG0W8cUFsmFa5X06c4pZC97f1iZ
qu5g8sW3bJg7VNakrCl8x5nNrFkq51JaknUyW8uf7Z8gVqUlONONnj8hINC+a/yS
MOkkRvKsnyDgeMY/YQIKOIW/4Zq5CzRVQuv+uYAhxnxPRxM8TqWCz3tNE8n1JMRo
HczuKQjiK6x135S+eJsWhMqFnXiOtZwMfQ2ubXffO7jikmtp6qJ93pIacoz+aYQn
RB5HuX7l3Vw5wEy0gB+a095YJwxeKOjsyR/WKs0E3ztPo8hvSIfOHjG4OQ52TNZE
OZcu86aunIYCVe7AajVhzc4+M9IAtxMZr1sIUiSv25KjdQ2XiqI7iQRpohj670nw
KiBureXD23hxnzbYLBAlk8aVUtY25S1K+P+O4Eh9LtM7CkZVwEsF6XrI5vg7K5nX
Q2m4T4bwbA60Lka9spQife9j/7GkCbz0BJ1gq/pHWSTvGGdYQX/Wsc05l9Mbh4q+
TQOF7XzEf4bRkjd4v6hq61y43Tm92zSZpxUQwsZ7Y1iXn8TFRjfKCX9/3J8WJmHG
7DILmV1x7AbVLRMZuil1NQnfB+b60q3XJ1OdsGkWKPdFKzPXVLviR/YI7Wzibdh9
nLRsHQvxYOEjY7xEpf7cTyU7BxYyc/njpCQHag8dNZhi0uBAlfTMv4JC5Dmn2ehu
2BXBwvRLG300g7nJd5AIoVyvE01BUHUFxUN7PX2SGDWkMRa35G0aJfsGWQPXemyC
s5YIEmjMe7y4cdcI4X3R8LiYpT30rR5QroesqUs+15k4Mu6W+2FPPNK4B1Znoa2g
YtUU89K7LNNQYAH5GCB/XHBtUoo9xR9PcRCDGge9BE/alHfDdh97oHbTb/AiGQlg
VqMqROWo42NjPakk/VAciTHVczUai2gR6i/KrBr2H/vZ/3reC26p8VWDTk1kf88h
UzYXSHrnZs4Cxl+AKIFjPymE1FSc4pQC76BUiUz3TUmV8Z4Z/U3VjZM6b1loouOK
EW5Cv0aesaS7HMeZXA06ScdJpYviOlTSQ9FuXtuCaxMGJcOOc+EOzx5DWwX0lhjN
D0R9IVMWlDebTRcK1sXo3U8wxkf8Nt0BEW0o6XivGiLLn8DU0Lc0nA7//K3SEtJk
iWuh9IfChE43rVYtC65oFS3QoqI7O5YXFTnS0VxZWvVXsXy5otPFDY5hWMKUPaS9
dnz/o2DBjHpw6HRUjaafznKCZCVSunTSLpRdqFOQ3DjHMjEf5i6eNL1R/i0Toub0
4TJBY2VVQAJ9BQ7Jfwl8HFzgo4NnBVihJOL/R+n6ZmNWQLbZ/OoZxct8V2s0gRl+
kwzxmr6w9I8rzOa8NLzUopovnmf5skiChP6KFveY9QgxaIMpyU7ws865qNYg+FhY
zk4Ufd3tBhKDDRORuWSOs0jaB9xC2TGfab9/fgtWirt2iYnK/afH89HmesE5jo2l
DguhLAGmwinng8nqPl8LXldsEVfPj7iqHU0SeabpukNfeORPaxLOcShYjIzwOdgI
humTaxlQ/qYMbzOO2rMSFG6/FBCtd95Ff/wsVHt1A34Cu2XX7pk732YX4SqFkaRg
FF+JoGAYUK2pLjxKTfu1w6hZ6VAhrmoC1wtcLaHPqaZ3Gc+gaworrVtXKnla44ZQ
xuuwO8mBmKqIhOrxvKEJtlusVzvWhykzJKzofZ4eLsrhQgxpaVgeEvHpkOGjYIEy
uOqiJuYpFvjSzha4lPy08AkNTQw/rz/wcjBqGX4HbUYXLvzL2nz5TOPWIiyI/wzA
nPXx206Fr0LT6LUp2+rwAymD28rTtj6U3Yoptx7jGqjBjrQT+Rp2/d6/oAd4U6VF
LlOFvUZKWsiBsG02kHsVZLw6EiOae8tlW2woDD+CN5biMH8pgsVrGK6zUGwkcCeM
4WTZoLu11+c1r8ukftzU75hFYDC1lu6QwjyOR2Oy9v1Ofd/kwhfH0amNQQFFWVXr
+kTwDuyGSK/wwJV4BS6p73xbUvJSSdVp5Zugv/cTvKq+sLkEx3iNOctYXGHnIjw8
G+bUhac3tvWvvWOXBSu8a8HJeQUpfPA8wvnHf/PNTPeH8YAmo1NgDAKEGTcC74dI
mBGFlP/G6kQvEOj5glq4rUh6GRaTkrfzF+HPq+rFcydrosmm2Qw/pvNGOsqlaYUZ
0j6eEIPHA9FWK0MajVJcCqYKHEg3fjnnRcLdCw8UVgM+HZ0yiRGn7EPp76mErhV0
TOoxLqodqBJ+cxAvy9bOCagGS8nSXadQckPLv36XUUsO6/h91479hfdn1lCgFKXP
bcAwb41a5FdUVnjno7Hiy37w5B7f1I8WN8FjnKd5RtSttmChQwed6tETdsv9pl0Q
e9svP2JuX71FaaX8nJHDQoh/IZsnHXRrXgg+4plwW6/eiEF7OSf20kqLI352um3T
x9WuJH3ZmtOuCePdLddG9cxaFiw0bB8/gFzGZt9gliteZZN0n220/7q4MI15/ATP
a3uCje33gBY/u02zFM6i08A46Dnq2xlxyjNEDPStTUwizaQnRehPo3FeiDiAuE+C
g0jx9nwS1SiQKVd3szyoede4DxT+3UwzOQsMy0lvJ5eO6fDmK1blrx6sTxnLG7pK
Za85gMj1yl1iAUQ0Ac4OftW/LYkt/1v47uvvxugO0nB6jAtXdJEZaNWRu6JhHJsp
XHxm1OARayGp+i7isw0UaSY0ZRNDBGKZQENFrs/kmTdksDbOcLLPVE03+gDHdCzU
6p5R9bfv/Y2WGwpXvKTOOpQI3QjmG2IDtlOrxNtW0B7t6cQP1QU2pzfkQorFfY91
R6WzWMLdTS+OE3cM+FxCUoaUJAviUSUyh3En8LXW5tl38eXQug9TyZ6vaqD66riK
QeZA02XEMoMNaOIQHIlOO7rv5758WHAwt9BEUfXN1KuHOjKFAOOjFcij9FzGjN4k
50uoG1ADcEDV/Tdz3wh22vDZK0EGut99WMgluXsHeg1KcEkNq9hNBTZUAYXvObth
Z0ERkkQEpqnfCLG6/Td7gojO43Hk88W9LqilkKkIuANlBxFv7s2kVWfifhxVmviZ
O9CxwLFDJzo7D00ax9UKZ7xsGVJDCS2JRz3viY0Gp5M8IxFr9CUObSUj+EFedC8U
aF37iLJ53x/27/oshMFSn9/cNhR7O8lkbr+5Xa72vW9o2E6/JhXsxLc+UnMPRz+S
3+T8s7XaT+WAuWr1jx0h8JMFNzWz0mtlXeAa6bsQdjWOYeruJYvitXX2S32Klj2z
owT2VrUdhdXKPa76iWtCACryzQTZCfXHU06bDtzz6SG3ZiSHShHca6tVEG0u4G2K
CMID/wbezCuru/WV3jw3CU916OYdhv4KFQRGaj3gwPcdwzPPf9VJ6L/1ICQT16cI
rklljiUH8kOsNZXMVfWE7sLtnghEP7X4tUU3HhhQ1/bneFpierXhvB1Hxu3Z3dsA
GQBXeyz6XXpsDZeRFMh/oyhnzaeKZipq1G6dQltbBfpqmlEPpAcUsPFFAnlOlk3b
5jwXGD+ayj70FkkN2WiiVtmMhC0qhYUbkoB6xPEvt8ResstqUMmF3ZNN4UgGkDRt
Vh6FicXVbUtq0LVa2BMoy1/rTmYt65sg0LpbByBxuk21V4SN4OLBC1ajTt3/SrO4
sHOMNjuQxpu/X9vhDLSg6+kMYC/wkfoAp1n9ms7JMVFvmVFuxNVFZ0k+CaLCDD9r
DuCoJxIZtYVzppZvdPUCAlriyKV5iHB07Enp89AGYUFFNa4I7B0eS3uzK18hn2/0
5adSQDYTkxWbTWgpD2kjObHdtDtXwMtBPXh5ptgd8zm963+Tor/Vd7Beo1PxyiAY
kn1AlYlRAiMg9zY85xZPCnIGHOR5VHYoMv6sEysGL0+OlqaEELV5l1/4CjRr+X/Z
tvq0nJSg/F2gbC7EeVcHU9BJ9255CRLRIU8wGYZplirFb6J8qA+9X7yo6UpxmoFh
5MHUk+GiASuyCYQGz/7DFV6jRCHfc7WDGJNzy3SvoaPRjM6EzCdSSv8M3JXkLF16
0z6rcvtY91zscM9gD8Kb6a0T3007+m4gKYnzc96gGDgJa26+4i/5Huz7yUz2mX6T
8Q98tG23n1jW3N1H9WelS0oqdkTBeeWYS97849ZP1BCwQC5djvHrasr8sAS9vKjy
sSgwj+Ky4NKWezcUnh89JUTzkN9uSIR2kLsMu6/X9iutGeIsRxjwietgwiiT++B6
LGiDgq2ZE78E0gFdRBYwuFGvaKARapbq8gRsXm/WUAgEY8u8CG34AFf+bZf40wLU
IbeP28dY6trVuCpbSZ/IhutCE+hKvIoeaz5uqrVoWWVbfL2wX4MjYbbTTAp7anD/
6Ydd12CN5xbgzKIeYnmcj0Iv2bMXZOFULPtoUXT8lfTSF0Yh3Y7dxwSViOzCI+JL
ot6xJJvy3a0yOB/8g7NjqT9llWCz6U13FtFIxhOXT1FlAAl+LguAovEkbfgjKyFL
Pn/iDvHZxKKPp00mxccnBbiqyu7tVrz/1F0/pENE44I2Mq84mf/jXvzb0v+TLWPv
wTRa0fEWigTfzmbBLdYTh+/jBvokY5XTMh6Pu9MDeRn/mC7gxHmBc3tO6/VTV92c
m7j3zrjIC6smloFGsmkwq5Pbg+GKaBOqhb58Y/SCQi/sBZa672wsgYWG+ZphTJiF
QQThxlV24mjYukIHGurbFrb0NTF48pBjeJvOLQjPd3g3GiR4iuSIUU1CcNLMH7wS
I8KB/3zDIXXEIchagNoQGDexAICVbOZinNZWafd/3G65pAKvW7FfC69oLGfHxvs/
nOSlzJsUiIRcfWpRVD4if9mpt0LBOQPMCpcLjuNG0R0zD2QeF6CaPq8rVy2Aos2c
reTlMcgAlOPxrkBbRHfZJsechCai+cLueUhaXGLlVADuLHK0hWeE8XvyyvAsv2n5
pk9rjY20rI/iwM7k3cVH90rUE2cCzrPRHSJjtgkEGbGmYpybsdn2VNfsocR3y+DS
jfjfC/P/0qtVCzoe/iIYeJU+5DCBuCQGMDZMcaGguV/RB/HePk0FTAgGNRjc2/0I
A8PFbUtmkjVqH/YLXjfVaeO6L24SCWHR3iWDDTmq1aIuj+WMKJMwzNiWvNfsnpKt
psfF10nrK2WAkP5fzu6d67quC36J1/E6v33BG+Dk37uh9mMQOZkXQ/OWq+nv65AJ
bbmXV2283mnkyNmXdiX5hrUNVM/9p1aKrD0/eIkm+mycvmfy5ZxVLQRzz7Bn4w+r
xUSvhf0X59Fck0+PNfb9Pjzr5I7PI0OzcJxGqd1MNaSw0i1gPI6d1myQHUf8z0Kd
kzpWSlOg+5PgKgSVAXxiPZ7cOuJxUQbMw0a+Nqd8LVipKIUF8tzBLvBO1iri1v38
13XOoJQG2oWuWQKJtKrydDF38X9YG8VKX3sweG365MR3Wb6/ZkYhyXzYc8pGBJWT
Mf1/Dcc4fO+ZPqAbsYwxgnFyojENWXIzd6GblOxzb/pU5QA2RtmfmHy7xcjg701S
qdC0nKG9eBIKhgcQ3B7o0TxOUJn8LkU/5EN3rg7IxGnKMpoGxVkvqpjmY0wkapCN
uoFGNk2TgJ24HpJ/JJL9xcfvsl5lLdxph0Ih6DtwH55dGCN3tWPODfx0j/3lxTKX
WLnr5Y1TWlL0el4enDC/CXWKkliPAbGKjCMP/msvMkY5tZuvLM8keWyg4xfRu59B
ZH8adM6aUCAyqtPYruLGt+EH2pT7014lvzC6FifwlsQZCZ/5srkPU56F8ulvQ+Q0
nu661SGk+V5GSIhEgk+UsBc9K2f5foqEo45jej0j//emW9FyQTGPMgTD0RlN28in
+hHmP/kgaFMetAE9i06fvfspM8E05p4PvDixYglLiRDp1mPx/wnWYU4NGpvBGAZc
6f8QSPQNrILwWry37BpVmXojUIvD4scw13oAVE4+oVf7vEkA7jogttYx2TwoWrRo
DVO/UqXbWV8NuY6LQPE8Kfp7Jb7NsrAqonRUkcvq8HSSHdecFrBYQ/aZOUJ8ua8c
Y02V0bSQfqlXAHKI+bVRlvemMFD1KPlyBOqJdFKnB9rHWyrXKyuf99GtsShWFb9m
n2ZvjDSfryxgnqrvzo+YFXsrICyi0xvjzIragxoSiSbmy08AId+ylK7HQVIQDTVy
ll8r0WHqX8JLJjP0BlvMYfGmogFjvsZprljcQqUNX6UT1ca/G9/Ea8AbTqsFlyPC
k6i0sdtp05evPb+sqvLujQKAE1SvMNM2xn8zSCC6X81nIn70w2/0zc+56wU1KeYJ
Iql4tROdiKA7I5VEMHtqIqtNCscidIMyPRMok+/+Dc4mRcEAPQe0nX7Kxkneg5HT
fj3A6grENNJ5CATllf1c9NO1GXgMqsbM9n/snvYDfAzK7gYtMkXDUl3whc3IfKag
tQuarXwUZ2hycpXyZVWu2uxjDmK+DKFZ39xLG7e6E4RQZazW0Bu2jldGNhnmKYGp
Vdj/OMF9f3y/QkZs3qRDSRVF55Of34xFKdyM5URnssVSNaOfaPVTWv5+lqdckmpd
en+sUUutm3omSTbX7Wh7k6ClT/NOKUYboK3I1gQ9PqXCrna5LISa2AusOgZHIZWP
5uEUOFjoNk4tbhROcMKAHNNcCN4HvL4b1+sSco3Ma6pFpL/HEBqDtuL/HM4gdVSj
oOyACYFqbjfnH+lbvtnKWmpgbxkPanGGcr8eOwzHdeGaoyZZZFmm1nMRt7GeisZR
3dS0aLSHMtZZz3Me/O5gRrwq5jb8WjvAMPLJrNeWZmlUFsNSmZWlAJfRsP7uY5fX
MR+yfYox5P4GBcodlsrzz4dea4tLQeiTCdwPa4jB9QzvCXyAzSP++opAZqF6Fe3j
vdx781BluXiXS7OEpK/ivzW5JzgsgGjzFtouM98UBIUdQJbvenx0fM4e1R1gg7I4
yGK39OCjfJf4H6vtKHmr5tWJAtc9k0hMCMsYoDaUvTdaq0bRHtItqVo48Y79KBgI
K8IiQjnHHMwjF6HIIgR1jqZM1rx5iCOk/mcnLTHeR+bxb+lT6zC36jhngIM0vOsH
/8khIEh1sv7OPslcIkNnmCl9M72Wl6DRrThF7O35XBwFuygbP9En/REJznvAyuoX
AYCPHv+BtAgegFbKE6N9W5RxZgiW9EGDSB3bgQq6ZeRYNb/y5j2ghDWnhdOmVwjN
Fa5HE2WlVoIamqG9DoqACFQIX0WI1uvYSgbj766SG1v+sBdbuuTJ6fpIEQqspU4R
Oqiq4u5uaGdwKnfrRilsjuXh6Vo4oSfW6g6hiMDSuaq2Z74RORf+OUlIbhtnH2GM
sPNmqkQW/tk+QgyIWxCSZTu45teTptfUV3JNBjWlG3PSf1UrooXqra2u9VkZ1s2X
qE9sqaFq9fs5bTkMOwjI4+BWqXZkGd/A1wN2ILRE6UpZ03/tQGrwPu4cVpAVHNzn
SafJwoKHprBqalYPtXFC3FXq0LPmckYivIoNXmJIGQ3eAFloIXnqNEiFFj8WyBcm
gVkzMlPVMAbUT/KhT5VlHMsQ0fyYoepQa9u2t8mh95AK9WtJdnfczrGhvMT1x4yE
K70W3v6Q2fEFcdLk1qzBaRXtZ2uDwyZEtXs8wN2+qLQZWz+D+nVKVRm0pvmN/MZr
CYQHBeMB6HMkO0fCoD4Gv5d/RAC+xc64dc9Nwinc2u2QzSOj1fzlesaZzx/sAPHs
ylhk+REVhjMjgaGhPZm2ttUxR5J/nP5Hf2+jEItmzvoArO+ve2li0rGna8gNHcxC
yOiWOojRbfqqdRhsnMvqAwdRjZzzhUFUOXUTiCU/2+cFxih702ozqIXbxZp0jzUd
4Gn40q9+ICmIXI0UBMsH81fuDe+/pYfwS8da0ln3F83A+9m1h5Vjv5AFCcphOeAp
2H1uKeKEdO5k0gsgo0+AIVleq0We7bZ8Mrlu/2eXlXsSyWzVKoMN62AnnEwfRFS4
Jz2kpLZGTB5nOWvllZCtheTXTMHBunNxWYBproGUCWtveNsd/Vm6Xn2XJIZOfPiA
aKH4JcDEgtV+vW47lIX5pdaCZ/6dSwz7JoYwavwkuYNNmlArd7bORvkBjvtd2TC9
30JbEo4OgTC6Ev8PvnhdXGXvRX5Em4UIkwnU4ngzPw/rqpTlr2QGUN71wPwHgBsZ
x477IokbYGvkLqg07RoAshNniCUDOZoeuAnycIwzS9z2N4ughYALpWXPhdSC1e8n
0Q2TRl5VQum4Ni32opLqfjq7UYF3Ike3XDgRAFrOKMfekBPWAeBZlgdU2XGFIF1/
UIwawF+NJ0OsgvE8cGATX/MshPf6zU4olcxeCICZspZDyvDhQWVq5f6Ry6Zy33F8
rXISoXa2xf3Aecx8u5Xqys17yDG+YZWRMAQ3AibbOf2+zuXyFjQdhWoEhU8qJiGZ
hGZ2PnDiEfMwTZ6aUPDr3PJ/LcHIYcb3bgFZetoP1UUS6M2f/ldj5ovRaVfPK4yo
juaJ2XYA5GCZ7ccN6xw/yAjVo3xz2G1arQS1reUG4gQDRBZwP3AXSGu5m7B94gWt
SScl1+Ou2iSHtYu3BbaJjr0i9hWteKwZz4wGgalh5A46WARUJeGCAdMLh8QsEo84
F33J3xq0Xxaostcsm0PZdLjR+yj4CoeHybEEiW9JtsdHFnqVchKmiau48Xy64eDd
gUnrEH6ymFOP1bTLPhQNtG1LUzQKXt4bPfKqAc3BAijjm375sTEavNLHU3kprWJK
2z0Yag+Y9mZYjOLNyjNLOjwZG/AALwzoJgWWAEc/lhFUt5gHeYoFGrLHcf+yvUYB
G0RIVIGqYj1gF6S5TpZdd++vv3lwqCtJthfityf3GtIFPjmUcsVodzetl73uMTwO
80IWS0Tvyq8O+dC3OTisKVJkrRa0dF/DMiP81wZCqLRE7MeND/A7IYs8vs4Jh4fx
W0IXVpOr7Q6eJ29pf1cO1liMeq7AKxWZ1QqLDkBmzCHXdlSN78ivix/Zc1EeqrTR
o5W1b9CN+mzBJ6SqBtb2D/2oa5LoHMJuFCISck3RqlHsm3fZ9/8ty1DeJab88hdJ
OR/jAAULmW9LHstngf2LZdrqowWBC1djnPgfqeZxpvg83soUn/7DbOgyVNJ0cerD
x5386YVZrnOCoC3/C859zAG6czFI9sx0NSZfSy/d8PAsfcA+8BfDMJRXkqFgbRYh
eWtOBGwHk+kkXSHsdn8rJarRJZNZQKY37HNqDW/+tZr/hEZMKJrkkdPjAjP11wsr
Ve8oIivDHD7lH5h4BzA7vt121bXfPxJyqj5zEhV8ZtBb9vePXbiSIfqlLZvy0che
VwQDg/uc+XthJoJMbClLA6/YDm2/W2eqreorSqqqb7K6+pcpFMZx5sCNwLHqeaMI
Dhoqn1PEoTSCgyj5j4nwDuvEMyJB66pDqhKz1BB7RurBM+gp5T0NTRufNojn7m0M
fhMDqsFMWXZOnMAsdj/kpA4hSlefeUltDU3Z0vv13LCh7xhnUfYwWtZdaWyejFo+
/ev5d6EkFiiwZ2TG4Z/31LFP5RoANXtXHuEe8GzmKojEEzEUcmzlQUf2octdke8w
xaPR0/aiyohLkE/WL4z+P6BfCPJp8fqeAAfvJbbAtL2QBH+O61Zo7cufl2cUIlFw
a5+zhAUMC/RaWEMqUjmoC8G5VDARcp2YilXX2uKRir2u8/e0UgDOr0qOKdwIQ0Qc
uBGjJ2OjRYVRAo4qbGoTedZBDdHLzNhxPfEEuu76cwuU/yrUsCtHwMlGQ+ACwiMw
rI7Qt6B7DgsBlz9HuU3g3L37L/ajAsfiSyWkH91NZL2VwuGUpeOa1zTkw0Ly6IXF
mryFiNotT2jth4MnXylGz4u6PYYiz9LhSCpg1gRmjm0BjmDokzMeELmA9fWeksA3
8Sk0XY42Ur03S+3dWxZF1G9UaDflOR0uQt9f4WijWeX3wl4vBJrkDZz8ofPQ0a3n
KqR9Mn3Jb233+xa7WC4gbUgEHNs28DJkCCBLe7xwkvh9TftcOXiPuqf2SMoI7MCb
7OlbuOwh3HwYYZDFI/+TqGgpK+/MJBLzzkj0eVgEo428jl8Lc0JfMCIXlOWz+c93
pk7proUI2RWhdWeBDF3Hmm0sb9Xc4X987pYXLj3U50bSpdWOP7WNKDlvtVmvbwnS
2R127ZzWbRYdh+NRli8D5ypTA94XVsAh4uincKaa2XPC1uNzDX3JvpWcZv0kP2rh
0LLjnvelujFnM9znJrc/m7UYTL0liAlChWRSSWeO1nZ2EtZdWqzD/JHWGnn+58gc
DHlg4CYpLeG+SjNCzyuJslNn8C4TOVyZjSdTtJTlgpFcKFgU54K3NI4N86oVhc0Z
4uRvj6l0BrpzGATtkvAJ/lNFeLpvzbWU63Y3CKP+JqijGEOiR5v/OBu/wwJ95Wlt
sfKSFJw5gFUB4rgBUdZTkwRQiM8Ve120AXj7p8dw2E5xDYM4aO2tWQePdrVVOeZs
1kGe9MYyAqA7wE4NXkSmrQIm8JARR80cKnULqq2D9VEJs0bTIZx0njoPEBZUjXzO
W3uxl6QypoSmtw4QYmJ7I+QPuYrbPLLhCXNnGhdoCdgr4jxshqVMAq4XkRMPre2n
QSxbV5vqKCT976pOxESHzUT5Od3BDyatrjAZpfFOdyUMmld+g4XTlg8Vu9yJIN4C
UT0u8ypqMaoH/f/51kO2U54RVW5pw5CCmv8a5i4Ch+6r+FZ3t830sL0g3YOA31tm
PwWjAmd20ufBDDRTluN1EwC4e9kyZwbYJl/KCf513C1yFj5R9012pGeadYIH72wY
k7YQZ5h7uBVNwqq1h0BwRJJpRAuTXhQPhumo7gKuyQqVEsH2lzWhsd91uo2A/Ec1
mYo8/yBV8xLI5qcVEAoYeLfbakWzYtLRlIcRqIskJtsgN3NpHwRO5aqk9BOY10tu
w6uAjmZ+UK+d1rmGwrDUuruTC8BXCyalApvtP9gfiK4tgh2+eHME6HJZQfXnEDKU
C3RO5zYmQPHhcGk/0otif0MsTlO/184gGkwmSpZe3wnlXRhKPpN2sUdHMMPvc0q/
eAVNPFKisAUItl+fPr2XcqPs/x0nzmNKMYq6usoy/tBO7f28bCOAvjdYg8fnlch/
CcLYYKCycCLCXy4kQEUxL4HEIJLIhn7rKd7TrBug3kTm3rWvvmqbcdvQJafbWovu
FcIHVEWS1BZDAqMsrBC/t2NLfYLwQkQwQhGimAWY3Ed2nTeR+IXlURAa02zIdu1q
INU917a5wjuOJ3OndBdaKtjNJ/KXqBRh5Vu2NugkpEx8EEUXFpmBM4D4hyZwQ/Eb
HdBUvXVGgLlEAJo50cczr0MNhWOxvYPb5dSYwCYY9GGwdW9DVGkcG9Aj075sR25a
URpOT2raUJJKfbVWP4+9fZ0wA7d9hp8PSBQTez5cFxdpCfqvVEIU4lOP94wJkrYn
1hlfVrRYoB0Gm9VPR4n2Fn3GDgUwS/UNQyS9SZXYN1Ywve3tl7jrZMYmjgaVOwxh
8yiLcdW1ew8oeLj+xibUhL20imYUYsypohT+qEDTMpmwqmdD+C9FkOfGrZE/W00Y
e851DkrZQAAzp54TgHpyw8hzCE2lEJlFybPIqndxsPqo4rjd/9VLCnAxLohIbBxB
iwcEQqckFtXNazlNQD2wdT/jinPDvJOoKxjexoolJ8iVRB2gZHlLKH35OgnrSop4
Z5BO9T9ETJvZaYx4nttBz1sJDIDkDpjjILr/SKORG4KynY84r9Q5HNpy7c7Ta9EG
tE+swhVmrFoZsaywEuR5oLrYUVXSKhNTe0HJ1inzjdZfmuX6FiK6G4hx25kDPw/J
lJB4Hl/LqlbwGtUAp+E7n9wszm62fUgHIoodoNDNOTNb98IyFiuNcMuJ5kFzIeb/
Om7Wf3GuRFI1WCf0p+mywLvVP6R3nJsviKiCbQ+YzPbbhO7LdPzfdJ6gugIEaSp3
qDJy/QklilghXOCpdSkXeGUp/5ZyHvGwQJdY6eIMiUDIPTKjQ1GtqDu4EoYZSzO/
Lsg2mLcelQfZ4w+gJ6gr5oTrkqQM3PHI1wUxwxLetuWijW5oyg3P+vTfdoe5NoXI
KYcVc//PsEYcRpKqNXvBQzoEvDzoutmPUB5QkU3GBPtUPTxe9/s/ESxtF2jmUoZS
xq8jyL/qDJVnP6tX9MXT+ZbxqQS+/Mx7H+rTN6+RuxpdJEEXEvR997DnRU4KcuDV
QFTJdVn51n2lnasu99PgJ5NEheorsGCG6WrqsaakaBEW2kZ/AiCO5GVvwdSop5/4
wTQbVfRD70O7EKJl02yR9Pa+S+kZqVFvjigRg38oU2vPVLkVxbEz9kGll42pq29+
/aGqJ36odvQS9EuT7gskHB30wKnW7OIpZVgSERupQqOb69BU4AZqHXmmFvlVjD4O
540C1yq3EvgSNPekT3NyT+Ugx9mu9Ur18FlcMyOPR18POdLyIPUyKbipOCjuaANG
dXZCC2/5eUgGPIpAth+blqODerrjDR/TRxNl4A26w7LPG3rtsvspo4/NOFwSUfJx
kgB73quiXD/rJsPCefEJ/n8xWXnUjt/0QrQq/QyK6QkFaiDGwFTuFeywdpy2v2zu
ttrTo6O8ijG2jkVk/2oOJSDZd5gpqHg4XXV957/TdDvyDxP1u1TZdO/YtEG8FfMH
nvjYQUqlEe+DlZ2hglLizdrNf+r+MWkuC4o8RuDEBpGcSN0HMsWFShF/bhaU4Auz
Hthg7v7Nu6gyr4Y8gnKE0M5pMRBxFfyB50uwiYo/mcdq0g4ZyyBsKCono2BnkK1E
jVRvWVVb9YSd9Whw2mJuVlfW2TmsaplUdKypCioxYQQIVo+NMbu7Cu6frzemrxJD
rgWmRMALLHAWXlhnUm/ifmuEbCVyOWz1ykiqjTrK6SB8dgKN6tk8eFrA/IPJH3QB
g1bsvqsuvjCVtEKpvunDDXHw17sBaSRJqNnCAyCIIofKdiuayKHfP2zr6WdGF8w9
zGZplnHdjhgwrEn1bWdodeh+W1Z9Ks42RSz5MFhz25nTGI3+yppwYTF75ExUtrkE
CXzIh3Hhy2fGvYJHxSXIzRpYAYdKj/pR9h+6nQ9T+5Hq3aMHxzTzH0DIiVcB4dyT
Tc6O8zue3v3xsbbyNJSTLNsD1r33+pxCA41usMT0bzjtE4LhAjI4DdaCUa0vyM30
lPwicJ6eZpHLFlV+4FY0Vg6L5hT5mr4dBDdu+qQWiBQou37mSqKHlQ4OTh1oyfWZ
v+5ofD6GCj0+w417fxGwLnCodaKgQiE7cYfxGAedCO1YZ2F2CfLFJFz6+izk4Mcy
uf0YyE6JQlw/KL97BV9kj4CD63SMRWHPQHKZ8TzvP4jcFG4b02E6BD1a8JhehQMb
xoijYZRMCY79hG1tc+mkAOheje9dZPspj9XaUak54FR82yDnqonMYD7O/EmHTQEc
FTbj6pnPCKY3PxGPAEyaAVyhkUdUSttCn8tfPSazDWM+rlOLhlP7sh1gMrlAzTGJ
zxJl5qJ3ADAY9vt+eFvJf/yEZUcIjD1XcC5vafFJO7BViSDdR5wyZydhKSXBb7ls
LamOQZq2ivRL0etaTJD094OVC/OUS9ElNCkzPw2VOUkeV8R4fXu9G6lh6bPqwVax
720l+LcJEj+KpG0+yziBhRElMvaMFvbniEQ2Cv0iP1jM1Pr9AX2i1jsssBWFzXcZ
PMDtZSFsjuzO+XcaITP4404xYl48YsXqKfVYHfKFqlznF3coC4ziiH5o/jiHYgoh
0vnV/sKVq8iNfUGoWlqF71I4VvY50Ry56KfaTfVW02MKQxihEOTXtgXLbxpUDBIi
dN5qoQ6gqKkIQgvJrkVQ7YneChZia6nfZDVxfQHhN85C1YqDkt2vTAVHiezegH/D
7jSibi85MFnJYT5qEduHCA3d4C3kFBMA+mvz+gqO3W1mFJ5qdQUJ/svWhGnKhCJA
oVR/qEMuUW5x3e2AHuUiyFwVdCLKlhAK1a2I99VUi2c4wyeXtyPm04ilfa/VgU7r
pE6yjzToeW/FWWOCJH68WaFwUyeKG8c/VNtXDxVUUnJt75V5NLGHG2JDQ6WoyLDV
euQnZ9Bhl0AvmNHkAXjSjgUtaxDTzcq0sKsCvvCvFkatYLHr72igndSpsFjdzGua
k9lBl3jRrus9u5xIQbq1dgCBu2YHcsh+4LMTOnN4VaCfhmS9WiuDf/03Oc0foH10
mMYDn8viKR84tGBXfryWIFeYpfh8TnnGG96Q11tOLffhDjX4tWwrIg7Oe+Jwx4i+
fvVY4zSrGXFut2jFAIGgluzMZg8wXW0ZUsiu4o6yxmYy8RKE8pW95MregI94EQT2
6r0Fo4Oznvu0vN3QeEas7Rk+ZwUQrRkYZFw2wYZy0hhhaEMk1MfE6K1gXdCxw5/H
xZkwdHQTMbWjFQ5UjSvqgyCVHp6P2ve4wOeSzPfsiAx+2nyym7Yzn9A9Rlel3IOX
gFn+poS+ZsV+lVL5RHZPfF6cZVwW7F+ipsGUQgFVLFrrM4/aRHY2tkm+3AbhJiPA
slEOcGP65eu/Db3Z2Ng76XQFXb/j/4sf6rgrsBx8BgXRRFNcyAwk91ipz6GVX0D8
ReBjqoLiv2k3Tqw5VIlkmB1HE0zLZNXRhUra1428pevJW54+Moz1eXIu6bepdChd
7Vb9YSUn5QzMD/BuIgz7guLXjvnOauo0HURDi7g0hwc/ZdQvJ9IZVKtOyKTtSxNX
1KX925P7nskGyiYH2CIVgbjwVt74f+T7RPEHsaIJ37cD8fc7YVY2rQGFQwlTsAtk
6r5kLyoW1NyxuvEIQbn3tIrai5aZEPEXRbjhy/1s8qH+HtQV+0LlPXIMklpoLWei
nmRpEdczb9nS9Rcml5vncCqiAvMsgGC73E7hGGzSi2+9t7H+grNHkq+EKZpWmKSr
m9H37qPkjly3RJlEg40AhV37Yi4rY13kw8tm0D9yqrsb6D9j13/IKZ8aoVJctU4D
LvvPcRm5YDhakPNWRIuTqp6z9OJS+MyCOTSLvBdRnwFGEnTi871QtMh8JwELzveG
cNeK35GM/tT58wqq8PExnop7IHYfLvkVwOF9VvGbLy5FG+4df6XndwDsDu/EwEyu
0lsABAgifysfpJvmFQyTOjAWyZ13EWJgev421lsI6Yn6dYCKPjY1vrtCYsyWLp5O
2Z/HBS4XzigdO//+SJIRK0ApEURpwP161KwJWhjLBt9TnO5TPTsM8qv4roZ9Uw7I
8v8mGHBXIruxyHLdovTl62uJOIW359Rjls6qf+gz2rqfR6cBlHxYQlKlXVQOsijo
kWaiBlQjEL6gu63xLPYAF4dV5sYkTukL1g7h8/EchpOdcxceQL26exDxy/omy8ZQ
b4suA9XOuTrTS95Rs0jpDKyKwNO+K0Y6xJiGu790ZO/X+R29W93uGo/4jDYvHqVY
wTC8LiTrrkvsP6sf0V7qMOqiffWhclRMDvrb8ygCpAjyrJtAaQGLuawKMHFqhBg3
N4emTGc5TGa3PFdzbzC8pSfnD8EkqT5y+JwiQQECM3gj8FYooBaNj3nI27EKvISE
jid8c4NetkM7aKd1WKb1cS/N5HvebiI9WHaGI1EYijBYyZrkB+wUfqCjNMMBSIrc
QWAphMWRPwXQh+KG4EbvfqvzOKfTO8+J1QZBqlhAYr3CMX98y940wJleSu4xqX1c
HDILtn4UObaA9B/K3KamTHNR9C3Wl5oWHou+eya7OqL6Rd+zs8pp6//DMZRzlPqR
ySbaJi92MkowCSDBvmORK49nw9O+0LHzWuSlfZkZeYSHb8t8qfoutdjNEt2z89QM
eEdvBJUCZt48ZdixP5L3KnIM3Sorrk7PyBL+8zChzZJGmqrP40AZlRLgE3lBTey5
pC2djFw2vrd6+rUuaCcRJ9aizvmtoMm9HJ94oWJhdPeL1kGumdfXuM9BwdmNFIY2
Z96Zg9FyZxGv7cCEgQ2tX+likuVH5KDII2TEIC+bkJJuZ24x7aqG3vp5fUn4Js6g
Z53IuCS0TqLZiI4M9spDObSYMr21Q9GAwXQla56FzXLnwrxvL7blsa1uRZKRK5Ei
6C16TBbKoxHsXdVsUjt4jpmleqhtVWEhnsOg0cxxyRVWHnMs7EK8llU4PVdv90kG
YO0OiJy3STUAwy/rcieGGoL7NYSTRcepGDF9kMbqh5qxarK6vNqkgBvbp9v92e75
HdxNp0ZpHJ6H4gL+4UD80Ixdiq0ZYTJQz4KfIhozrUUrlKTKm1q1qZjdFrmxEz0Z
3VgGhisv0v3FC26BYmypSr46ymikV2P/86gQAA+kMIwNaWgBXXWGV5YPCuMC+ZVd
laZs3iajc9M+5FDaqwJBiSynyf5QnL1GyzKhpaR3AyDQLfFctKFbcLlx0cEP3Zf4
m78oNJ1410NmnzUHlcJCRA/38QjFimCO9ai0O9VtZppn6ua/zy3IeyjxI4Al1r26
95iceqbgGDiTzwlj0/5bw8vSnHUXc32nALuzEZeCR23ufdqCumGQnziYnYh98amQ
F3qH44PdTqpq4mTEkjRuA6oKKtnYk7RXy/vpI3j2sKSozHA51uc+Yeje81CvA+6K
qooQ/o4v0BshNqwAGoUY91I3HWMYI38QqVvsX/xrZ7FO4CirVwXjMNU0BAgHaKci
D/VR7a2wVsk6O317NQGBZvilJPpJ015ooRKsgcX/mCwHdkCf/A3tsYkCFAwLgHr0
B345Vc4JqbPgd8w65SIjfaPCqlWR6LmdRYMOcIyiwa50fB6rjSINDG5wNbxNGHLr
wMxekGA1IuUZ8X41EenxwviVL7SUD0n6C0SJ0L3MJ0Ch+vujNCw7DxWkF4ldDAHg
2aiPNxz8bUak8xiFcGJ22ssjoeNgG5MYzKEeWS9h9vjdN3lC1TOpCdWQkKwSNEmk
R4Ukw5s5dEcen49cAVqgeS88jKE3JEYYaJH0KHLi2Hwbgm3ngcjjDk+cBCAHVMxn
jvEVzaVLWv8lb7LDuf8tgTBxKZVgKVgekdWP4JtTTkvMflW7E3p7PBgq3dwUonDS
5848jHSwMXb8p2/4d3FWH0K5a2wqPC1yid6sYJeO1oZZiQIS+Ig56+0aLsNitrmP
hr4tN9RDfcmG1XG+3MnH7jcd+Ds8YVKnPC8n7UvWQS8aWX49ML+Lcp2h4+z4FME0
U9mnSl4LxSk7cICiQLeV9KWc7QMAb7IaHVnUAsU3trHtc5s6JZtOcHUPNXChJeRw
jPzp+1Z6e7OYAWsaaLkCjZxu9MqL+AKvrd1oe3AdC4dRhYl5Smsfswh83FeHUa36
cK6Tm1pEswVTAdYcIVmSJu6Nxvh1y4+l5fI753ZKrx9qaaa488NfBtszDtCnzSnl
7q1jurBdfFsT1JSfst3EVQ1sQcB4tdnMUc8+a7b7Xv55A63mYJlxX6u9mS9/sE8Z
935eZAv0QELUq7Su+GjI19rvhBSCsN7qcaXgwc5PRijShkmvuQXBOtq98VWAWmav
X1ilGBjtCskxOSAawV1dVvwVSA7ZDF/7CvOFGskRPk1pmMD5QUZ/XDKolVOb02a3
XyO5YlVwxmyQ+w+oZnNDtmFcpUWJ5bU4N80Co+UGSEslVnTW7cdiNHRQKQiSxmrd
TB54QHNSwcW9cDu3DIJ30yhhPki2CXzWS+gjjtIruGy8u5wrPidu9RgP5Xv3TtZ6
dtyUO4/LNJsFi+kUdKqP7QUVy360XYTeeT24wwo23DtYpJpJLVKVSUaQeNb2zWvs
KkQDlrj2E46wdZpCYlIhBsp1dXgeFFzWpLdfcW69jVNLgt3fH+FneNFlkUxXwWeK
rwt5HRo4HycryiAptpXWf5X+Wzo8ly2TSbBCZxZEFlN5jyRm5mQx1JsHDFSHZaZd
Y2C4qvXySDoDZiPnr67OvURqxUr2s3kAi5H7SkeVnWZgPZfWSAfDvSzcNn5JhbO3
/Qc+hQtjqhxJPsbm5xyZM/DYb3V3bKG7NzJQ4MzVcePLbzZfU1r4et/GlenKt2Ys
U+0CVilMiJmvTdz0hvEg0ms4wq8+qZwxwESqyujgnI6VzJRdEx2pfS9O2ZLi61Wr
+XX0peFl2AEeEnBrEeFLH2osGBfgn5Y523kabg7FoMDn+EKPehFGErJwfx2rXRVI
+Xs2ulIWBSvjbx0Vo757VGXmtVeDWAJ20Kf+r90XF3NSIyWoX4KF8P4z/y/nwlTg
XsLZ6dYo6jEwNY3QcWS9lTbrPBq1Dhr9r2FQ6i3Itw6j4Sy/eWZ6WuK8BJ6YDz3y
Xbe8sUs3rQ2ABYXOw/j/9Zg5BXrNhtlGg1jDwYay3H68jmh3vtPGHlGioOWTXgwh
52NEtiXaPaSnIklmM1x70j7PkKa0rjK7JcP/Znp5szdFhtBXzK9Ay3Y8onSDK3zg
M6KOf+2nwd5yTLyrPaFKe7VPNueZU7wbHnKhoB7yq9QKR/fe3AapXNpMe0U9qC0J
qZ46RCsGcXfufZtVk+9ZmiviDZu0mKMYiBMGwFMg0mgQw5pdzfwDLpeNKgiTZAR5
lvcr9ZzWyd4drrJ3j8AnD9Gco3OagiXqwvE0vNNR6OoQ1IQb26oVdn2Lnwum/zd2
q8NrJ5h31JQhDJeKHCNuuNivkdIVphDrjeDWpOu+lOYQqk4LpVg5eLkCkYfA0y8z
b2v+QDjdHzr2p+89Af++sh8AVa1EJQeMVaFF8NYxHg7MZIpOKATwycdv5H6P9bLC
tcCvImzyBEW4I5AlLAAg76oZ+nIrqqxihkIicYtAs3FwzJN30dNaMlWVH47EmVGN
DMtk5Pd36Y1HIQTrj7qHkoL6T3M2cONjA0QbDw3T8Aqw1ts/7dBEKE/PlD3tV4tk
XbNra4qA9Fzv9tqloEl1JKByznOt47h2yAXfFodsx4wB0a1KulgzOhY50uwhmLUc
u0oY769RF7krpClYNG3bgkiBDgpk8VJWL5Hgaomjr+172pRqgAsgW6GbK9dPhc2V
4B3Lf5F5h0/sU3/k2342GzC7+IIl3H7XXVMVX/TDTZ0S//+eKtzGHeM/5EhukGgf
R5ZJZskJddPRCGiYK9Gl19X21lT9lTCZPFrwF3goNT37QyTBZXXFwrV4GtVjjG2B
c28x3ELrrrbuP8EsyPnt6G+dSWttRQbxPobGNVxDbpneHCunTDLRbWH/RjTjDxJ2
JfS7mCieBfgCv0r0cm2+OwutaEMZJAFjRITNI0DSwzuiLNP4eNxCQPmQ/jvgl/fJ
5CwPMcoHipGtVQzd6wXrg9sXhRAt7hqHO8t3JZoCTxXQwjUE1JMjkLR8Sj0vgRMi
WN9xNRlNWcfYNU3GjL5AsBdApcmQc/SF3our5kVJa67S4/qIb8KnTZUY5LaNXaBo
KOKyxinafTdJgsKo+X9dw6kBV0fMX6PU0A1wLILN6vU2KQKv2/Ws0EJv1aR5239D
xGwel9/ZcOY5osZWWzYXrgV7sx8r799p/L9ffZEta8eIjlPuJbVBWDHiYczs2SkJ
Ugy1Xp3N6R2o+TOPgLzkW6YIjifRNl270+hFUCiHVpJ2K4bcLmilxEb6jWnwhTqt
bk2QECfOUXcWju4eS6/UNsZiHTenk+vzdoKkRUE73QhzkTt5x/oL2Muq4lG90uvw
Gxlr9UWFZguEgPiZ0KaZwqr9mypmTCwAHY86CJOAbqhW7t3Ino3TZ911/PmVl2oy
cXmO5jhCxfBXhQXO8oEKOlNcEAxavSWLVm2HacRKqx9505Gx4qqVfYss6bpEN0aL
pT6+FTMblId4Mh7WxsT4b8oDbOpWn33Of1pjk4Ije0VDBLHkXsr2AMKq2YbrmllD
Qas1IP8GiHLq8993OiQ5gBesXG1gUkZACPYkGy5eGuE4SziTXrlHb9sRfgNpvjsw
z3fbJVAAaXvXp2nJcOJbDr3UP/Tcyb27uMdxFuGU3a0jsFwOm+8DMYZpd9NXxSUZ
3sDgfC6iIHWVmZvJHSyJFQ9/kM+ntZmvoENOTfmrqvGv2ORpA4UszVB3tbgylQvM
xBoRcjhbG+dvbZmnlWw6tNfpTbxC/ZqvWhZhmlUZzNxVLDorNq3DSUsmdbtLskGE
peupSXmjU3VubzUhtSB0Ex/8dO1wjLbLkubDEfDVIF9Ph2iQTSmnX74IYatbPFq1
9pYrW0AgA7/M5WBVAixy+qPy/PPSt6/Zbc+m1u3prlR/4r2DumevnogN3b6/6bnn
yxCF6exJ1UKktYbGRlB0uzbT9kgg/DxViDZ3VvST2OE/YzIFjchD6a3msKFDA2SD
Jsw505fk8urR6gN4MNAr3AYLRw6DfSVEBxxOWDWEQDHN0gVdpUtBc7pOkwTnVkl0
1whSOvy5JtsyxC2iAl/qBsd7ToRU/Gz1Ii6xVqVvuI8zEJpNPG9VgLj1ggYOrol4
nONK3oROmCSQl5gPn6D0koyo6S1ycAhqi6ebQpVQEVjbBzsMTwHnl7Z+/F+d0kSL
+6nUj90vipOZ6msbWs2HfhxDGU6TysMS4aRV+TTUi6hKdQPkseZX2PWEYX17XufO
hjoajB4dzC6KUANE6qSBiI685DBsaaDdhnwP9Vm59qwFUNDKF8ZIp0FbqeHlXzqy
RFOi1Fo9pQnXlBTrl3EL+CWwa/SERjWLS4pvwFOvO6OZvZLpYMlWrpVdOFEP0+R5
U1b4EVGtHWMNY7uqLesfNwhOpaND88uDcZLzCjN6FVOlGU1o0vL0Adb7d3CE3hLB
myczNpl8HYwSAu1B7sK1cSVH6tOzLGNkymNioyRKcOZWwvEgY6Ga9F794suDPvHm
vgsy9e0ky9zmQsAUCbJ6If1iJr1DlOxWQ4VB42sZbJ19qLAz5thhgTA1nFbhP16l
zxdDR8z81/59k5u/pK+wPuJ9H+CnmRaie1fr1QdJuz4NGOJT2F1g/TiSrJp8gSJS
Y0sHFt5PuI3hnUtPWqJIujhFxXc+G64FFZ8teQ//Znc4VGJkF6SwQue5DCFdBXE9
EG3KFsNsprKOWj7PNF1pB91/JYvWWNHSG+iC5SHgCo1Rvwe6LNX1ro61GS9Iy3/E
xWD+OV9LSeVodoyv7uSJW43B3AO6Wrk4dnGRrklBbLSpeJaMzcvOaI0h4xy32gPA
J3eRTJD45JRo1aYY3NfV0CwpOh65Q9foggwH1PXf4Lm6t3mh0GMNIsJ+aluQixxu
eS5muk6hU3Ka93J4OhFu+yb/sgrbn/JnmaC27IZ3iB5oUd4xve/UsYGRyDr+q9Sz
n5hCqWb7tZ25mtiH1R+/DQcu59r0rluxWpIV5OgWtRlxxuWPsx+fIuL5bxo/Dlsd
YAZqMjYw0UurXr0LS0jct4IHAYowAi9fMFxPkFgrehsADVKrszFu6sofTJ2yOb4G
1KfA3Ht6Qq9wFJ+YXMDtkHb5/gTJnwpXygqaz6/cdKBLB60bLBcOTD5mbRbdv1sw
/WkZnGlsmjZMzHHWslP3yVyKkoikDL4und/GL/3AejJsaAo9fw1P0xS4HkFfmgWv
AaMjKwGBj/2DIpX0/SNfBOYrUmhE/0IXJjU4A8KSJYtrwebvzOLmQT1b8SKnSrGk
aNjZNZarhqyBup1zsDeEF9P8HtJRwkmN95S5naLz8jMQbhYMOF07RzIVcp0MYomq
sHtm961gRdaDGOF7DHBbym0HRD9v4kX1DooU7gH1mCwcb9IhefpN33lrNCQxPPDs
+LE3vtYP4nyNfSdv0Mvr59jrnyuni1TKr61PIoHkh/u+D/Ifi7Mqr0rHAbB076P1
GQe3Uet8KzjHn+wLz5E/p2euEH0n47v5spXbMNcPRudy3CwZ9knCbfnzl6x3NG2o
dYorNXPIkVvi+SfKam4yMUyXf6QPTKDzOFLHzXK7EoWy1IVZRdL5lpw9p7XCk25E
TOpYHKtzZRFSCTpyZf1WQCDQHe0FehtvBiis8B4uSJL+4FQTl5h6HKmo9vUygatk
Z62YlBo+0HNP49lB4KtmJwefvVkljFiGVVRdvzyViALSqq33FT8HEAlvYHaduMBm
F1/2oHLqQJ6znOXRD6ZHKfFl/bbQPsqoY8b/ftt0BidmjfOeE6JRcwgxxXun14wU
wrxIFzOlq6NXHHbZKAkw8/1uz0nEj0rn3n1kN0RZMdVrl/X9XQXSrNmMQ7/AhacX
paBnhyEOoIj16eSWtWqowlh7BejHnzT/aAJ2ULPNaC5WRW0MMNnl3p+TjnLsqFHr
v6e0QjjGhKUXTOUX1KDvmdkCQOVnGZ8VhxT8E70wQcrDqZBD/O+81JvQbw6J3HSD
0BaJoFR1v/rvVBKg+KpfU2WQmlGl8fZe8cdM1OgMcQMp1wHS2MgOiHV6gTtnqStH
BLQFxa4fzDtSW5NWjCvFXWTivMJBivB7BGWmK5xOts9soFyEPy0rh2VSJ7AEnGIE
fbT2uuk2uq13OrfT+IB42aSYnByuqQnqXzV6HLo0LNIZE7z2XhabF0YBx5kJScJy
pu5VNnmzdNNmNT7P07SGMJIvFcApxHYt+JVK/7eY4KdP7cxCROJ7a33VGGZ96Kxf
kP4Cm7o18OIgxMnbOWD2oydM1CU7T8k7H1a0xmlAI9s9hFe8qscKuaU70hbxwMoE
WUbi35VwH4nCnJ8+PE9xpTd8E6/S6yCxMgtbsn3KoHayxo5lEjMPRhmHT4wWZyPf
/g2pkaEn4rdtnVBV847YH7rDWhZBo/46g+DEFeK3HRrhSXoev49TW232dyRQDsS5
748hvhbnWT5HroWZb844u5H5WxKCmFMFyVigE/ajFNkOb4wIbxjAlpBfIImAGfWR
YqssVDvj4zE9A7Pzkjna8rUSLA4rOX8qedguCLyu7d0tRfHDNb4b66DiFfZV7yXe
UHw+9Ebus9x1PFj7fvtDonSg4IV1tLGybT3EVthvZJxvBzfT7y350N3PDQCtZ+IF
jSrc6RBCRdchVFilR1uaw/PfHMRutBJPuWyF/1NKc3KaQAGhO6g261mvy53Ob3dv
ZNV1vwIGu3WubsUpT9PJpGL0oZQV/PKFirmgoC+/Rwvf/5DuSZIMIhQB8CVxX7jd
rPgqjGLYoKOAvmOszXKn0O7YD/ghJjpjkEK2z+vCUJFMUuXSLX30GNwIe4bi38cH
sPTyGD53N9sEDDZJgrA1QVJ9kkNlLL8JbEM8LtY29ecSQx7p5+BHDG+37nFEtHtn
+djSq5D+jOH7BCdrDovnMLud5PTCn12XheXgoNDKVgb+XuGVgfpL5Naq2fss8S7e
Rk7l0aXHPtsIr1+9030pnBvohpxDE+K5+mHfe9LfAqAB4wIEljKiGm90Olv1Voxo
WVeYXGCo3SOt0ZAwaZvcmR27CLZnkA4koyvjDMkq9KWlriXxQrZQ9u9zoT148L/g
BSdujbIVuH1qG4Es4mNtO8JKnQUkKcLKsQzFF6BafDlTy9Hu20wVahlvgjBkwFl2
Bwr5vlq21PMIzBV/DhWeWezbWsUtdA4ogzFsyYTACg9EIFeppDlcM9Lrn2qWsCrF
6HZdJZ9IbTJOMQGfapsxegPlAST8WlXCD5/rxudeRaIM55B/zfAr1b/eEyIUkDhO
oyfWokGxlTqHcvTvxqZ8Dy9TCdceoXwDlhO505wA+27GipzLiBjI3nc1N9lTdRuN
wuTrxeNbqDtT5sy0H979vSr/uK49rE8P189kaJHqU6cr6C+b3O/pAaNWIwYK4IcY
v5XzaK1w1cfQlF1G146i1kMSIYSgiyMMp21oeg+54Oy394Ok4QmZduXSGOfKTHAE
RqG75Lgt2byBvAHCT42jdc+E6kzi9X8pC9tO6C87cmhcD3O1G9HbzY5oHPd4mzC7
a9e5E/oCLhqNA4ObEYUbjKeF/KGkfUgEUVQTsxvWjm0De36CFtu0S4Ggq+zyQsb3
Rvi/BMGHQb2PjZEyemQjL3mZ6+jz/pzE88a4GUTM9V4PYDrsMcVwa9GzzzU8KrDz
/Xqddiu7MM1f86/1/mzkfhBZbI1SM2y99h6+SYEHLVbiLG0dn8g5pvg/fhqaRiZq
Sug8DCidroi8pJWqkhdDhMVTLex2RYQXuRgIOOl8rQ/Q482W58LNucvQ5THS93ZP
VtHvXtWZTjSa7h5RhraNq878OLX9NXkRK0zf4tnWzrkyHjWLYGYqq4/tYxP9e3Zh
uCaHcSWgSRpdIGJN5ofTiU4ccX1vid3v3HMxccW5GZ03YDqlnDM9xZhf62oV9WFA
OIdqQOlSibwf1YHJYyyb270rlwzrzHednSAdbdfRHeevkYv7QqJN8Di+5pvB5CF6
sh90N1cGeBssA7/B6mHkNpbXNRJX64FSySE3o1VQEMjOMxZiAKI+RjBsOCDWnCK+
1y+7yf/JXvO5CwGQ0dlbWeCjjdr+dKjFZn6ixmqGfFDm5Oq+OKqzk6cwRot1H4sq
Plct+EepQlfRjzXdNwbqDmJmcoqIWkTtbOs2/2tyqb6LTQ6C8ly/ZJ0NSD+h05D0
TxCtizSFUxyKXNPcbuyDx8cgLcLZhqSDYU/2d0ufrD1ARg62Hb7TPxAwBiBRBga8
iHQokkNgOuEWFAM/gO9olzbcartTZ7zNo1K6RS2F1NSsQ+dnZ8LtxkY32as19t0e
J31H4IDWig6ZtSkjWiGuIRZZ18QMp5qgSXCD7Kky86UjJPwQZOnKNXvPycuZLDTF
N0EkCj9Hv/DmeppsopR9MgElxKeIVuThoTqUL+bX9LcgWhP8QhWctTbOyyboAflf
IHnml2tddx/WHTOsjbAbLtg2Iu7cCXsqyDWihjOoHrg+8Bs2gn8KeCpucDRtmyQd
hkchwojbrqV6YMOyLzZkYLtiAEwkNB0+A8P1DdygNyOBlSkmxjzbLgnG50CCd5G3
fJOO/mT6RdP4Ie8kmaQ94PkpH3IlUQX2FlxeVOfSbGl8EDR8GCxBwI9ynhxGwXX1
q3U7vAY3VJEp3VPIhzbpIuye4Y0yR0C9ZqeynL7P7ves0fbLOwNsNf6NSeIbBR0Z
28NfFr7YFWfomXZVgV0dR+w//xAD1SEuS8G4Rl0sxkN86m3xPs5WGLmiljhG5TE8
jVuqG91f15Wq+AQxZLfTH9t2YghJvvcJ8pNZB+ZQfmq6sDAEHiGLoBP6+Ju4RRsY
5RRFZYbyJdsagiXPGeY/XexBwpoyP15vye4DX9e3I1NGjpC5btFnymwHtAI144LB
z3bJtDv2bQ5S7UzhboHgN8+OaSBuBrRfeqkVgbr0VgbHrJmRl1sypQkOzorK/GLC
zvbgIPvd10JCBzHKJky31mbsIBGEqXDN7rSDYQBd64GyIPyYQMYX91v1Q53NFwcF
TqDy5LP3HdxJ8lHwUWL1cqfUP+g1FB3E2cMTOCEFfUQezFuqArRgA2KTht5J+khy
+u9LXEGkN2IyLwjP5lPNYMoAxoW0Xi5SdWVAjXd6VaRPVMHcPZwNrT58ZOylrJ5m
wgy9g2ctZXBY01EARL+fanonG8P8rSHvJA1quOYH7G6UnWD1/uwtKh5XxR7oV634
xio8mgbqOrJFcqNX6bz76NpjL0HWM57qrD1i3WM7i56B8iBOUM/9BK3fWShuip29
9Ji2nZqSMHdR2l47hq/kbo7bfIe9dSiwtgiPNzhUzI2i1gjuj0D7iD+7se17oUpZ
56/g9GO8hSdnyXL1uZ2g8IAAfNeSdo4R+3qSKIthuLc4YzsJoYdh1jO57KS416lj
ozxIARbqSn+4XjwOWi3eX92KNL08PhXNna6R47udOapJN9YghaK5Vyw2Dgph425u
QwNgH/zfjnn/QA7LcpxTGmTjtxvadd/fjsoSd5SEEF3Ga9mV0/G/EBcF9HpGRDwY
N9agBMcRV5pdmU7gSrqGIyZ2vkH0OSsnVsopAmrZYq86fuyHi3OkSVNi7WKHaT8j
a6lrUNYfjSDvcNrfwfBWwuQTt1IKiTekUT3xJfvf1sj0HJyZBCdKnWgcNJQ77/nW
HnnLb+Yz5kxyxQzY9TPtCB1U25xeTFx/dM/+8s2K8NBZa/+jqWmxO2ZYJ43g2OeV
+iyG6xhjje2wCe33FFclPxWsIIKk1DtTAftg5hGaep2daJsf+hp/dCDq6pSCEmc4
gybSgBZsWFRhafdPBTDGgykaR7U5AbzaDuYU5Mz7kSM7M4y+zu1Li5AUghE/mPom
oxdX/yo0cP6K37DKP/ZA15AQS4NLwBhYmcprgeZDdERkLWwXFd86ErdqrymHk2eK
PcSLFsx3XdCcRzaf/WlKwGm7rpJmQaXhFU/ffPLZbXGZAVHuUF4IyPed6mzkNl/k
5khEI8RAbeS8W+YNX6npoXznuM71CYTCkGxUc6tBFwhHG1BA0wmg6DItR2Qb2Slu
OoyYSc41I99RvPKqtcjgcWxWO1p58ClLzCAmFmhP9z6mkoIiHhqXc3cgyfqCEhUV
E0wQ+IGi6/76ZskRcEsMpwaCmLWHvKEYSyH7yfXJVMKEmUXfBQYs+53Mcbf9/oKB
b0ulEnnk6aexIpr+90JcqnG12ck8XRpUN3AwOHp59lVIkDbf7SyqTIQhHBsHvV4s
I9hjXAUCTTQCmpWK0tC5WQ/Zk4RMMna7OaeeFTl/p+nC4WZ1V23vNLjcdLom3MqD
6nwz+cc4KGXhY2uacnaDe9Xb7mKXmeeYc2ZP35dssjamWnwnJZna25x7U+ZwCXbH
UMPqBgBEI5ggmOVBHqdkq1de9J4QQhjQSTGXG4auvhxVCbRJylRhaI4Sk48N7T3R
6WFN11qXxSON6I/ClGXK3oud8l1xHtcfDbPSdAVlEg9zarOQUOzgpRVMVHab56oo
2ot5NlZZFFaadXNLYEsbNWNQDdPpGqhTDFgf2VBWrvf0VPW9hWk2mKUDzPgkuzbF
zAY3Ny1PS+THn8AeN8IMIUhNKieQquSulLwSKQ/2ClG4x2mMRLaedz7xQHFdtsIJ
rpaCDT84IBt5ouS1TFzRNPdK5gS2AT9ftp6zlcObqJTZaSowKKuwG2zz/xJifjZQ
EJ9LQwmsTLCFMpGwxo6wxp1N6zOftjf8LA5oM9+1JQOsovW6ORcZ/bQn7WK/IkPg
SrB7lZKFRnSD84X3r2uKgWtk1GAp4q2DnQR6lHkKMbTTffpmaB//qoUY/U0YQ6OX
/2b88Zl5KG0CsSji2bck4fKDgZxPTdpAgw9WebG2M4Zu21HXAgJlF0VIuX0mejZB
6PXl49WABzLChhyKXg1f1N6c3W1YclNZSBthc8xYMxj3VKLID15EE26PXqtLIKcU
0dBygyiHmnkQtA3EHuGX88IKZHqdIzicJSsTzbUOSX2mGtAe9IuLdLjOW6N2BKS7
/6uGerqXIVxidcZoqzMvLCh/lldtjyOyCEAxxCDgu/NqeCSrwThOza5cRcVNvEL/
lmGWqRWffLzR0OCDKiyYbcDzwGWo/tXptvjLN20sDglHEeBZPmlIapRXdjUELh78
RlyFR4teBbDLCyoTTOBRRWbDAiErbPw56OmPzVdEb9J5AgFCUmzPTObg/Okwbwlc
Xiqon0YVV0TGUgMqpzuNI04Zugu6BIAx940AsrNYVkr4BsEyKgScew/4SVcELr6C
l2XoDrd/4cROxsLRph5FzC4W7XiiIWPBpcamYbi6qdZYumwUmgtEgjcWhbDXYgSe
EyI/pQzfJkruqEi0SJljmr5GGlkLpkWehGDt/7vM+dBhNGfWRcPb8PTAYO9CVsLI
VMhpXntnEdklFtUkIx5vzSNTchagFd0Fvi0OldSeM4Q4Wkk2JSCB3d97XVuyjhSY
Et1Hy8DXg0WClFN6F7mk2R/YA94TcDr4jEyWkwWEvbLlN5GTfT+zoPjnRotqipqN
71aF2zbcWZGjG1evseuGJcD+Wg7A74IFvR2L6Bqyf3M26ZU2COoPnp9WaOsXVuec
bTR0cTqXrCCyJs4DKZEL/4vua4TDwzgLFuBhx9nZ7wVnFeYP4Day7YZy76nsA+aT
t+yFkTQ0YhZW7Gb2g0GURy718ZphhwlBkS+JNHlkXXzwacwnPuFB6aIJPEoat6hB
Zm7YReTf1j/7pNNxRjvkqpEK8yyDP25GkCIUAoqdPHeaVi2enqnsNuJ/uTznoeGT
IuY0N0/AcTnXDAAqVbZ5XiZA+1H5m1QrqdGIj/Y3r35BWziyvsW8/BhqIIDw9OHP
V7CwomiroJP20iqdhCkh7aqQl3vu9Uc+6eRaFeh+NbgZgKq8HrdedMkmRXTNgQBA
rXYbM9AMJ6el17IFXroE+i0RAiLjWCzZ3Gnbg2IYax9NgNkJvuvWk5zjx5JHJi3j
Hep3VJPcB54icCBMJDYUG7y3U5NkODUMJUKGeJ0ivpUaCuHYE7WHV9TY2hnzOQse
G5o9zfXggmHkH573P5iqphsa6/rSeu/+W5GKs2hZkAriaY86cR0NX7uCEpDs7lEg
GYzZQ/rSzsMqj/qVqu5wIy5/iQqnLbfGf9cNvmdNOxRgX10Ri3X3YCRnaZGbDGKF
r0biwuUzETUAvhOfc9ljXRLY/8pjUrpyuQzxsYBpvD8famrfWjygfK0bTFfezzQP
qiBImCasQVUTQjacvcLVutyj9ZlU0ltPokuCSaQhX2Om0+Yv520p9QypAYBcmXtC
ewkVXUdiVh2aUgp9oJtOSCF7qtjVn5LJDYoW8kIKiG98aTW1HPXjLNbOpM+xbBee
MjiqbEndYBmdDzR6oARPZQGWT70zTSaPUOyPhGWYA86rc6hcNRFtOyIVRR6GwJsB
siwqYezZA03uLLCMOEzmyEDeJVwnpeuWcEg2TUOhlYJRtxYosJqIkkWlElaequvK
Nv9JtRcZQ4QCbXYRHSxx0tK5BgZaa3gBuhpJdujDGz7XAbikfO1nyBujOmToHpFj
1h5e/gNkq0MfXc+DMBfywuaBDxMGpl7s127ZqwWJopWX7s/tTcvtlCist7yb7wt0
LQMrnmLo/dNpz9aXDPpvZlRjhmkFqKXdRYo1WxdTuygZmqcbeyRB7PFfxWuZ9UwV
6z2kv1gScsQCeCMups9PyYnw25jUoCSwBqcsSnQ6jt5TkAowSJd5+G9sRcNIqbHA
vbLpGVgzEwH1C5dL6qX27V96RNoDzqWLJoMew6PyQTT2YC+4V5impnHWHjvUerVh
CmTZcoCMQNBmCi+3ijq/uN2QJFnitKaM6rVvDqhcNWKhK+SeXMLEl6NXj4gYTctI
LEFQZy3Y2KCbxftrMWFSTcB35BSQif+UYICejK0K/VsxxknLlTztHa7QmEbEqRYX
tnvU89bLUKZJ6EDwzXIvt3vWHOOisLra1cBKHoxn1GprFi4Er20VVIO4SNbt0DFD
OsIOOaHiUNH+a7fcyrChehC6jQsQbd7ooHs+1605Uf8ZouCpfG6XZ0xSiuh6zmVF
DlhOBC4wFqm/nBIJ5ASWyXCnwDuDYtexibIYT/30fJojvyQc9SjhE/aN680T08CP
Xs1blu2s8/h46Nyr3sJC08A7Sh1dQbgCH69DWkDUuThFALT9J7YY27/IHyCmXh5i
i77kS8qtI29K39pEWTxRHFrJdWGcu+mxLPBTGuMt3pqjwkh65vMlVgyT1Je4bu9F
yHub7Uqsfcha5CbcMLWcOo8+t4OPDhG3jF8tPzqaIgxhJVVYAoErFEnovXb+NO1p
JoryWa/d5BtewNsbN48IirX9pgKjui3pUEU6/r3nJ2k3mrQqE0yP/Hfi/YznvzrW
yq4QyRfV0XIIhq+nnomCUK1l6cr1aULY7ozjJ5rNhEeDfxDculid2s2r+JsANtNE
7fd31IEuz6gQomF1rlYWchXXGlO50titlyZllnkzzDGA7fwpagSwe8sT1lfJwZYg
rCU32wQ89/6DjgD9bbHHCHfAPuImnjSSvyEKblPxIAoDj6wU0w20/8IcE6dkQdDd
HEsRErUyFDUOugZc+L+mWcG78UklAWXU/mnV0lMU9QWdBV9gCqEM5kiTdWd95OLn
WEgZZRAkIU0EkKs2eQEdSnMNFdkwOqzKV2w2ltAyphTJbSLOofDYCzKxIPY+mn8D
S+GqI/jw9xCu3IIhNdNky+eQZPCs7DOWEnwZH8AElkdae//jPzjm99KWRC4FBhjq
3ezRXUScqIbEOOuzUWtdj9E4m6O0r+eMhz3A7SY8Qe1aIsyctEymSFm3omgLpaYK
ylmcQBsLyoaAo0+z8OODMmgc26NUxcU+j3d9olswmBaHwd4uMBBYkdKFl01hSvqY
0pZ8P+sTSYMLEpUBYpkrJgg8hE9ifkGAHFmrmzqPzpNeV6kM72Ohv/9f6BVjkx8s
9tUekU91SchdWBD+Z5Y+Zg/ZoBMmMUj4tKTifKu4jYjnMGsc9nHoN8hpiB7iSt57
vPCs5dZI4Kdv88M+iz0nmiujYwka8hFYxNZeGjBfZzL0J+RORXBepU99NJsWIX23
XXBoUr5JAR5K4ZiMNI93aqw/0i602y0jKJHtmNnx3Z4+abeXI4NBwlyxTHV4RjnP
TxiEI/71Kx57jYIm6H/4xmAJW0Vhfdx8wCeLfWTgWMrsqzb9o1OHDlVPmV1fTG2N
xnS8HfACegQJigUZQT4WvBQAO/uDlm+e092kwwQFL7bt5TyBjZB7hHSHh3f6mhwM
gKX/OLbznZKvaW0rqhNlpnnC2C+viJXc/08x9/Cf3jb6ulSC+5iPTzUwE3W5s/Y/
jRwdzGKZncDmF1+7KcWutCY2DJtvPu4Scc2uP7F4YgoqQPGoUxGRlvDNBI3cYzzK
tD4SuRxEdY440m4DRGj4njcdc8IuARfikgPYdVSitxQ19Ta3XXV8zeF7ouadQ7Xo
qecVOU//Qjrw16ShT2GlhGXPeWBkxP/unYZliNXP0LbQvPh+V0vaaWP9+WmiQBn3
jJEsS8hhPOpbSjG3UiNsL1RTYJ8TOc4POu0Y7zLnPD01/JGlMNFlhV8Pfwdk+lx2
INyGnYAgsZ673IX3mIusdShNuE/EFMqHrC33kcjY04qP0lTrUcVqzSFrsE48svUc
JMYvn2H988eN7OtJQ+kGSP6M7K5zaj5zedf6Uylw5AhmUNbFrxbF6AMxHTD8SDAJ
8d7HHjeJ8WxdIDnI0ARrpyMn8Ze2qu2ryr4XH6nB7GzNXuSpcbRgxbffmR3CRxH8
uYTLtG58ETQtDwGWHe9zwe5U32nFgmeBMCCYkjrzebLHfiq+CcLhrLqah1FxXCQ7
bGJzfULQOf+tTz9ryDHZCceTVaXK4pGodHjnha+SBzIbsdnvE943S2B6lJU9WMhC
DTMZs+XhpDQnxjGpFx15jMTD06vtJ2WlB5RGbljx9vzbJ/N+RSykCLF6afMtjXAj
JKTPP1VzATX/JuRpNOjrzGrv8RsU8nHeds+4xsS5x+QMo1h0kuKQG0SsJHxgf+Rn
UnTuhyoktoG9SuxbxzesPq1slCzKIeLy22bjODmNPGao2kwG37LbGTO4Z1k4YMRE
Pxkde6hx0TlfclnnDwSuy0gFcOyts4NuoHnevSmOXqqSz1I36T8jn3CmThciFrIW
9ADO/uJnKnWhUsR00jeEt3HOcEN9V2RFcRVa3wXS7vAd6UnCx/01XesQ9B3+1uhN
MTGCJLyjRdrz3ddj19ut4f/pyocR7ctQy3Ib4MzLu+G+0vwf775YJ+EXZzeCtpq9
+u7XyGu9qayMxoyXyO2ao0qeKMF3hfkVIC50s2p8SHdkIJ1R8iuKXX/zjvC4i7r6
3X5FaPSZwi3MrGe40mxWvEMbhqSd/xcdy+YvWFyAN7ium9+tGs03tl5y2xjhQ3JM
9EY3uO9lnqgALsywHzDaQYynhAGPmNbzR87gHh+jNE2HMGVW/cmBerj8xQTXcnfe
7TTX5MKquPpxWVMrrD8GF473U05mH7xFZaPU4PKWF6EPPgBBLtuCRe+gkUO2MYUx
yt43WI0lt+ZvXENsLeFTBVHhj1XyXsMsjUs6D4H6towq8NE9JH04bra4uW4Al4KJ
N7lPWtaUAgwlUaVoO+Kp53V+ObKeR/h92d/ZBuyzqLKCQcC0V8xbetr7uNJsfBTY
omF+G8CLB+73olAZn7aq7YsdvJcciUn4JiE22bL0J8XvG4Ezb0Q2/is7IKNICtlC
slwtCIVs6LzXtuA8bbn8s3hO7a0r4k33HwOt4V56hED1FPMkEYD9YAUJYu7er5ZM
lyHEUCs22S3mI2WnxKoycZm7h/MtUy0as9lPpt7F+2jbzgY5EQpmLzH7eis/rb4Y
ZUU85VO2/XG2U9WGIePwGniXuhIpvsCt26WeopIhhthjlxyKsAr4a7nOrB68pte4
Y7F7y7OyoSHOsMOoDDEmlNcmVCCb3Fba5wecr9OemgRHXGi/D3aqKnSeRLRFHT2E
KuQzxx9TgncQqcEUjm7fDcMpabp/pFGAaZ6ZdgKCdLkM+rO7yqkxDEx1FZwMw/JJ
4QMkhu57IAIo+RHTrWH658sFdwI7twa+QQKgCD3NlQX7o7NIOLwnD8MtiwV242vG
gG+3l0Jc9yEoHnGdZQMd/yf7MWDzHiD8JZVXk1BirbV6Vf+QwLF2PbWQpmQ7Xs7r
+XR1xAMyeFExh9tIbw9ezi/E5cIcFcLf/gvUeZ+OwOh//8zarmUfkqvT/XD3aWNd
AO9PCA9meByAPqzzfKlAhGqmk9mKue3GiNQvSS/drk3460TiNtwQ3wsLKENwhaMJ
vsLtKfaxn/xKvErsmyKQyyFz8k6ChXeRLqqmKUfWP1uaQphzxiVZiUOjPs2wWXJq
IysJvIKRfL2LryZkRgioOFKxgSN3FQ4YSq4Haba90r3Jwie2uDoEgtjioSv4h7bo
LCVGGHhnubSKCjkeTxofUMFuISS1hXSewbM2qxtSODe+YPZeaRjrV3VFM4tRfOvv
xVyi8bHAeA6TCOx3M3sDt+ioHRvOn5okzUoycLJMGlXLU099FNuaGZNEteZZV0vq
ArU3AoGz9gWqZNQVV0H8H5oJvtMKOlmeypTqPk+N24pOYyvtBEMbdMQekas+OmhD
qw3uQydHniXJ00UeRk06Sn8z9nOY+PpUufAF4aJhtTC1J2zIVxf8Hpix2fcVS11Y
kXYsGMmWxfIus0WIEjdAaSpQnKx93XMFaG3M49nrQlHAirmjDV93OaUn2VIMs2x/
HkfZmyszUEGEgZ9a2BXjVtbga5Pk/4hNidgZq8zYi2N8QXtQLUgA2woWF+GSp2hi
PCVVvCZmucNYNydAPwXkXTBg+MGY4jHlz685ZFmiDC/PaD9qPvjUf8h0Bmkq6rmn
q1bjhjcVGOPh9hnEL7jhmz14SJp/uOGTYoO/DqtTqdoRN+uxYDxL5YImZwooeHHJ
86k0HH51MzAm9iqzL7dYqJrg5idXJF/yk6YxK9AS/Etp+5o711lTgCZ5NQsvzOBJ
WU3Lq+YfB54FV75j2I4HYdbjADuqumHRkJ+T3mC0l7kjtSY4GGopVzsFvYXPIcuq
WX1o4g/z4HTwNkTfTPbMw/kquO1kQ4Bn06iqS5rLdJPLB9TnUlHKcx1Fr5Wj34M3
oMo+27AtQ7Sbn9A6d+ezrnbjweqm44AIZf5Nl0BMJe2WLui6fGnSPVpJASC7448E
6WekCbli8TKei2a6KqGu5dxuJf3QyAYiAmepDEiZhAoq5nAvyGBAHM9r0dKwMdmp
qR8i9bZ5UGnJWZjMIVCSb8h1SJsJrbG5QfeEnOYVe5qclrE0j12i0Q5g5t5oABZO
lqh/OScloM92MWbFh9TTQYAc57kxzlPmRZegCNc5DsUsYU3SSvJIhEo3Vrn1hgDg
2Vl0ouMGofBAIOMwzSTuEYexHAa4BHXMUOZzwaNtzMVP/qKnAo5pTQlD9o3mNIB5
b2/ybGTezq7xG7kDTf+zPI0F97ggKMKbPs65my2F7G7EgbqOqiPzuMCG+MdAQWgA
8FJVWd5lETB451u+HgxDh5gQdygRe3tJoGn66appRJR94oPsrzw+wnczAqSMCqUQ
B4g/5gesHgU1RmmBtxuLnM9FbadezjrnTys8o1dNlUHNKBYbiw6FHQ0WRx4zmFkg
aEU73yq+YbSJo1x1y8/3+qBSErs2xVM7PRB4iSAT26GdfchH1qAG6IRThWiimHD0
v/jk13Vhh9Yr5f3b6mrlbPjdqkz6SRSnL7RrQGdsZzIDKuItOtzzryoSYyCpDboO
1K2MqmeoMnK9d3A8L5D/Kya9E5IS3xXJYa/Fds1ixCWel/u4d/Bs9zCYdlzIbeGi
sI4eEl0yuxCtg/F1cgOCQPQ6r3oGHw5+Y/3xSxB/VbUsB2avL2E5D0mHZueCmn7B
7Fzlfj/69VXl1aut2LWvXparoFjJ2wANzyW1ZwqIa0oNO/EpJ/8bt/EBvLHmyoQz
2fd1M+5WOfFz82KtRY0drA/9tHfSIQK/F6efmoepwiYC5Y6c3qhwebnNtscl+tOz
tmYHz6IWxjvW5QZ1WfJin4SAAWwfqrsvzbsdgHxxitCOln2hmTOtHl8PcHWetnfY
cOCc+kzXShfRt6herEq0C1X9h0JE/bwA2zUpqCd+OqJsrU0CEYvAmK0KUeNDvx0Z
NtEVRHoMrhwGw+0Sp1FWDP3fwzD34TBw+ItB+BsVbr68j+mCG0Zf8ahW5cFkcgwo
GC1KNCDi0mdAfTXpApFEp8HjJ0l838ZLXhqR0XWFKV4YikZsW+3P/5y9PyLGr+RC
IRQ6Cjrp4bG8YtGUDK35AvRNdThdS8Vxagt7+lQ0bC8083Zutat3XQUKksxNn0D+
U+SgyVQu+BFArggMlHPUu+zepZUA+BbnTCwHwYxJDrt53VtbGNXAqO65qSyPX8sI
5bvPr/I09LGsBrufZWAuNYDN7Ne0PH9JzDeTeFXyBz7imoypvx2G2OSQn+x+06on
gkcfSLfHpJEHjizvQJaDrGRohyZ+tccElE4z1HIXvPJ6iUuP5Wr4gYV2kn9osBbw
BApnfw2wxL6ThPnqgQgj5hCXjuik6TwNqMQW75sGJv4SyTMCBanSYJB12gO/Bs2f
DBhag4Ds0ag5EM5TJ4TQNRcAg+vjFkn2d7feui1vb8z/R/JHKD4LtckfY82M5zsT
M+eHQrDnFy4KSJ+13bxpLVgKQFe7Agi+fpbYC9P1R6cSBY1hOTdltIilRNB1/ep8
cQDBdfbRoNogAYcJk1IKCYScxRJceGRTbNeVsDKQSoNNd8gUg/UcwXYamJ2GD3jf
4Fn2XAx23JTVFVxD0OZ8J31HZr1Hnu3iu38776zzSiG43wRDBsSQPSxkC0nqagPK
wm1LPUC1Fm0hlSMh/E0OcrL3dSwwRy85sNh/WICHSJTOEmUY8VCa9lkyLPT+f5ar
bEKEojNGVDN3FMO1Bg0S8+GFEJ2isXXWn8y+oZb2tUUh9HZ/K3uwNBeceEFJ6NB3
Q0iRbZ9umrBLFjhMoK+gE0FtOO9oE0sacb75JNfC0qxM37U50HDFwk/mwUhaH/bn
HVVaAcwnAyAI7902S6T06S9M/OxwN9KVvIrPUrYlnmIZN4YJXE+VAVvBpUwyMV5v
yDfivIvg3Mvtn/IPOsjVwUQqHhTP0qi2oR16z5BK9ewJlmPDwXuz6ftYyGcCqZal
dvqtJARE+xORDAmdni2/REyKxsxT4Aj3W5076K+Ep2DgsXPEmd0h70C06ZbDjYPR
QI+EZqhuqGTDKkiIaUSlbG8iQzfOBpkgFB7MwJrIMR2STtolhWsi3++Cv94TgkGS
B8DjHVMk+b8tnCeolbLBObRTcFJ5LmyIdqoviNWxG799Telz4nDFONf7PP3HoWDO
e+IZu8CMEBAiSY+cQpWqclm3TETdJrlYFfG8kkxDmNK+q7zt+Ds7d507Vl7cJKx8
F4x+S7z5SaYM5Ab/wVNX/B2ND+M8WH41rExkMMOsJ/vKf8xiVkn5FrCrjAc0Vm1M
bjTEU32+I4/qGEiCLWOcB559BAI9azn4K4OECSUGPeYR95ODW+xIRO0P6A/QWnoS
8dAgkHAfEQuzEGHQDZFrwSqXANyscPuqF6lhcKLtjVLgCkH3pZ3ZTnZtBSdj7t5U
/Wujyg93z7oWLzz3TR7FID0rlE0UyJ8gZKhk+cNsOBHnu4hmHenDXmnlAJnHuNdP
zjSnZzTjF+bMvvcQQfxhXN09jFmqVlKCaSJ6+oNAP/8JvIy0pH9hN2/8pFH1/OcL
1fTTdd4FxFyVR8/y2ByAQVwMhsbg24Ts2ERAPfdbIDuyMJZkEeqX98D7VIQJo1TH
FOeK3MddeQmbJtTKRry3EcTcbs8updaVoawMKrY93vuj5CZvbbRyILhn39HvLUOx
TVs6plkFIn5nVpSHjhHEKZfOR27NyubWx/QEzML0+56FyHR2ddEa7BZJQHzgjiTJ
8t/oXEHWPjTQgMWmBLcGME26Ek4MJMaC4JNVdmFcUQx7zyTHpRM3jKuF8Q+bqJPi
eRZFU+dg4RHawxOjH3wcKi35Hy2xJJIEbrO0pYmF2kQ2VDRvbhODKzOg4jx3gJ+E
Dl7ESSr3oH4F8wmQwVKUxdhDMJlCmESFXiuS9I+Wl/tAux9ldBTrZhZBXRi/f9qJ
QFPOOimh8LWsu5JthgIHWZXzKsWreTnnkSGRvZYLuRWEWpyUYbrdgD8eDv4bHVWh
caZ+QOemt85MQcyj4WkK+MTEb5cEbvIGQSNGRuIxoBm2OvzGxAyVrCsXRLuDgEJY
dBGjHjvY+nrMFisa/WzggQbcCj8hSob38RMGXSVFgHdmDLj7vG8h2xdO+XB3r8kc
STv24rFBC6Qk2vIk9xjDNi9FtW7PxUb9dfBhhRsMoKi2tYndWugdN2mS3SbWu3sJ
MYB0RUYNurzRHrkCj4vY/53fs2Y7kmeIWd7IR+MKpuaV3/lZOfXATmvR/TcF+ebC
Ki/f77QVOLP0QKraOvgBh1J+6ZzEz1DWCM+dUrEne+PBVLosjYuEcWhHOCXHUZtq
k9RaLtQef5OEbR3Xsczkby4K9m8xphauzlPGQ5+kCBAWGSUK0zPpu13L0bzKY1nO
Hr2QTRGibMSxk6d7A5VXuZ2EiFBVnqzaqBtFMdg+F9MFXK/tcKZ+QXTU0gQcSP6n
tgUVhnEJekPGMLM1wIWpzUpaqjeLbDl4GNehd3dGQTDxLmSOvb8e5EOrP1dPiPMG
jkS5/D920V/6si1Jii69byNpxxv0z1o8O8kq1mJJuGgi9zJOy74+cFXDxoLqY13x
UHAIFTFKUU8le4udZnwq5JaaaOUIlO935AmksihINUIHMPiOQmf0oPh+SnhNdOKh
VWSYVQZfSF080OynynuiEyn09dRl8e/a8tp/SAzdPlhflQ0fZqG+uYXUK1ylbvEC
BOtHQ7vh8OprH2Ph1YHRaCYFDS+dAYTAYTvzTiSQ3E5N0Jx7GdxoxKa4eNmTiaCT
fkn/riTGhiIMTtzGc0OHDkK6bM91V2ehMZh2fTaiRiX6DX2YDD5tDcu2i+GWcFo2
MXDDjMrryMeK/sNCIbLqTGsNWVcKSA9P/lDmLuCjAPVsH0UN+e89qeqFnKQMlZ8w
TtrMNou1Veb4xLIbGaivF7BZNTyFyez5KBXOzFLbZVYa4XMqxhecBP/Zeq1nZKO/
1utkbxxoo+Y9UATEhP7Ym4OJ2vSTnxF523vqqrn8LfQig3YUTXkG8h1jUaJOVPN+
/ivqM/WDN69V1DvkFaKnAauUIRbv2bNATx7nQy21Rfe4Kvm1EA9+jglGESLgzv0n
UzDeLAW/+tKmve3DK7XJ9kef2Il+Qaai++2QEiJ3LcZrNwJ7g4D8HsR1uITuCOoj
+ETZXVd2v+wk9Gn0FYr0yuWRJbbMAAinAFvf1uQdOFOYXu5jd9ZsiR09sCPPajuU
V4qNhgqhJ9gIg3hhOxL6pFakHEfAj19+q4p9mrCU9qbsPaIbXbSkgs7jSYYVYv8d
O+q3qDfaOANXkkddOAIqVG2WIVVOBKL3f5sogvf2WN1HM73Srm5uqGrFzTxeCj6G
j59hs9Ulvz/X3GcFIpZoou38I8uN4LdnSUvKaMxBAj2N9yeWS0GzFN81JGErXh23
YWDrWjyzsS8jRWNXVA5CPMwbuKwfOC6taGUJ19YwcqEvBOuRqLi+7B0ZbJCL7o1y
IHDiPQ0zP0H8EtqARjs7HuOIugUoHSwBQeA0y32IDM8r1Covc+pd9S5Z4i0/KlmX
Kmdy/1byzx+ndnG+2k+rudgpOYdgPA3GMaITm1qFiRw8Q/LIkmAEPd8laS8sLKHt
O4flH84RSy/2sWxuKWlBlcIdXqEy/SFTuZ4eYYXifCkxSahbrURrLIZPrw9cVyGb
6TfkobFVHSnc9zQ83ONhmtsalDafAT8lgNtFjYkemXgDS6mGWJz7dLyWUiuiuiQP
NCzWmLnO5ok88kh5JQqT6EpJAA0VR8+foOyIfbwVTe/mKfVtMfNNvW5/zVg3WaWT
oH66AdAhuKHBk6eaocAjVgnMYFBcfKI4Wl1uRlEWG1iVwKc7crRVQrnNtbnItq8P
RVuL+O8vs2EV7HAtlfdXVha8GbI8ASpDKpcQrTYbrCZQ2KWCShjZqzTk9svUCqua
pfXWdWP9Kfsra0EBqMnsT4ln3cap5kQsp/3TO3zMB78wGzgPh0dg1Sw8A48Kyjhx
4J2zw651bWusw5l8Uw0JFmUS3VgC+tJwoqAPL78o35QAVsIazKxnVGXYdKGodSqc
Rf5P5lOjkI/6pEUPlc6w7ycGR/d+tVkVu45s0kuMYc4WMVBaTnlk5X8EYAZ5of+x
T2rZXqCwnxb+4Y6XckUY9WVZ9+MbYS2uqmE8+U4ytHbZn1VVQGZ1Dl3ZexEJ2V/8
JtbdCkgpGqA2iwvPcVXxGN86i68igWPq8NQiUeIH/PDL9uhU6HSXHYXPToveqpbc
IxSQPjKmh4ZqEIg6MfXJPsTpLHfLizQO1fZWNlUyL+k8gX1tG6J9PLvJrFR+gl0Z
tcVWfFj4JxopfRD4c65c2tqZ3GBpleIStZQABSCKUd7wjZtCsXDKN9KjO6vZ/QTi
Ffiyqf0fADlcMjnCF8MSDzMNE+N+AjHnLDOilCKaXS8LWAW+ayz7DOsto3Vaeg8s
YICtIX8myn4XE5U1QdA7JFPSz4SbUD7cKo104ir0IcciDANks98DOPWHJoMwZXCP
uyrxU+Iw2/wj/2SOKLvUaYXSaeFWsHV2f0vcNggyatMzNLkLlVPtLr5u+dxw/BOf
4aT2fpkjIlIY/TyHsLEIpHoEbmPRCsgSY6w/UWzfEIGS5sel+g3IUvMyLXd5J0zL
n36QA6wqU/2+idLzznEsp+azTayb8E+gC1HUBygWm9DEGmwPXXvK6qPN86xZE32H
WUWD8/GopJ7wcQqiflDZ3+STvfpC6XoOPI4KZcb5e1ypvjsXGA26nQfZhDnIYU/o
rrh4rLWAZSnopaZeSyiEtyylbG9fwpTvhyfP6/vMH54HAWOzKejGzRiZriiK61Vx
xZWRth5ttlYMK2xwVrQ/9gWHm+OIw2KDKdUg0iiJ3vEqqWyCyiAG/AweZDrQ7orE
Rq092BiSdG+m52p+11iHxtR2KZEW85N60bVQwAKXvdaixfPBbD9h1yFOOgtQINro
CzmLc4p+hU/n4DHWGJCCL/YTyFzX6UIeKouqgAaJgTMc+bRZ920Ccmh4j8I0SHTo
rq1K1RQ5MJ0c0HKdMLmrzo1NX7RSzueJzaJtbCTBXFD4sE3Da1Y+sSvZGRZwCK6h
b1dSHKXh08PfUuTQfHGkob5+bn07NHDAaUzB54lFbbihjoMuPQWattH+Vx7tQx1S
VCjFLwN7B/xa9R8lifnjsEHzL9j9e8y4Lrn5arIqm8qlp3T6Sai2eNFTq04hldlO
TkWsICgIUD9uwYZm5DycQWuaVak2MxQOQs/WrdrjgTGEke0G8fxp6QohF6Bn7EcW
AD2ZpSOTYcJPtObjzr6KMLXNDPF+sL0x6oe8whUKOJTnttpBuXEt+P9h96/bIN+e
+OuI8GIX/qp0+K6pXqLpy7v4fWeiiTbaCT530nkFO1URY2ou8+h2WX9JpoqPcGCn
ZzTfoXw3C+H4Cy9YGUCuUCWum2w45wAPwgnH5BexAq6ioU25bfTwu3R1jxJ/YH2h
hcfHKfPtnHnaB/5uJNJ16hBoFzDVS7p4nfrdE6MCFZV0tdEZTMpo261lZKnn8tn+
6MNgOLMPF7P8IvCHLq8arQdJURrwBcbhdiVGOza59hFO3YMEKtZDymnSGuA4KZZG
5nq2QRKBVmuC+cVLgugoVePrX3JPe9VEQtgxbpD1l8D+PXE3lLTJenElncMIIOU7
OckLgvrTuULGGNMSKKDENwPjmzvsagA/br457YNF3CE9oUnSD9BnPh+E+gn5fQ6S
BoInHr2UJ94rPBVuaXiyrXzajB3jhI5BP98EiWDW6hNl4nba2C/1KYChRTsE0+Gk
hSEFXvE2B8QRBNpqNDGPnv9T2/ugwdWssjvXAuTskez51aTQZBsba+UWmbm8iCOn
qnj5GQ4h2SWe6QxzFZAuooojN416YiWiq7YrqTvNvb6AzReL6GGTkx38VXJ0kUSB
BuLT6FwMzUWs3lewKE75HTY3eeZ0NXFhvU2hqm4oqr/DRscHV7KHYGOuMqDkPbMA
JLIYBna9aRo2f6+JiVvfZPbSJYmW1Mp1j8CWStN+q3kipjKAgdrlbZBV5yeyTfWS
orEzV93l/r0vJ54r8wkA+6e6ve3UFN3XZLaHU8KfkximV3IKnpX2h/fMzVaGn8nk
vqiqOrT+9waGETmr18RwCHL8hUDs6pXWuwqxfZG2nYct4nwhxQdEP2beoNk6FK2u
jNrAhwmEcUkCxGEFWmUXELdB41zoMUbuZgwfaHd4J05b7J0gwz6YA0OUbEFpTA5/
p5wkeKTr6RlYxPqLCd8KgvHiO3D7P7EpehTo6TnSjqRI6Hk/QF6yoZFp9FHGE+ev
4cYiGLp20eOVuf5Lkbe4l15FXfyytNNCehGcek+KYIfBtUzL0CM7Tn6YRWDHf1ey
oazmKlr+XhR2V6AU3bZ2CDTzeNfigsTnHbs8kzAl5Mo+Xt9kqkom5swjGi8fOMui
Noozy4Jog/DRUev2GIM0TcXWe+s6h04lrNtuymftUQLE6BLavag04ld6H/RD4Bg5
uwKnl2mVspzghwYz6qSVlNApDLJiSFgZvMJvhTM8hfHPCvXhFW7MO05tb+9IDUFB
hrvB1ad3GMRtwrh4osaQJviApnD2SbjDtrH0mPMaiX685GetOpksZ0S8uqjzN9DF
5ZmLrHdmLYf4zEiKvxfpKhrkgdX6pGrYHQA3Rqj7aEzM4aDcbdbN3qFIGluXv1LW
skstc7g0a31BzlKwSZFY+F45UywTrhX+LKX6z44vM9NsOIqHDPP+/bdGEQam1r8A
gRzxymmy13/I4vADOLUsKIR2S3aE1h3AuqRwapqUYLOxKJRkGQ5TzxlriFPRYP19
G6UFny7PsHP0tzd1URSxY3XoBPMXQp0tC5bAYlDxsafOO25sg7p45SFs4Z6KS7Cf
qXnop8JVJGDlnSUOvbKZkkNamQ8k8jpR57KjD9x3ga8yFgUCyJHcKkZGC+JK8tDb
QN/c7IIw9DCM43p+5+xmcnxJduWA4rr24j4jIGeb6AwEfeXKogGtY5k3VhJ5EPvG
mn8+ZVOcJthjtQ5cDcnc/kU44PPE7qBFS+EkATqdq2ZVIIiXQTRwXc7iOoMH79BY
V1zIzF0nRQU4ODbg/XN6YWoxu6HvOFPnP6kPMjbK7e1sPlJw+xSgnLcNmMhTmjZa
Rts5OJ4Jfiu6AFJcVWdolyJvpTpzOilGqDDlgMCzKvHGE/TXhJzj/ACSEwQKcR1u
b7Ysd1IJ/XPVrk8pRBvcm/Tmg1yKObRlbpA1xuzJDkWw40h+Vtzg8HvtcMfUr4xV
ZJVvWD+Mu8pCb4MJm2uVxHHw5LhZvLBRD9bFija+wSUkp6/RkBHZGFZ0nxguPgsW
ZV6tVbSZTwwjBlnlV7HfeNavpjoq/znH9aXdaSG02BddKWjXlBuyNtAcaNLxi6KT
fHvdgvp+t4o+EO8x46ydSmhEzpTmmiFW3bN37tHdXdNVMlSt/7PUCwkbDfBsdgrw
2l65Hy0gHmGJLHPTE/WQ/7QkWfC+CLbGN4lioCPL5jkWabwJ9XbEdeK2CiPXtBwY
31Tc4Wq6XoLpu/HOduV4D13GletY1FDTS1ue4nxrDkMngLq63P2mSAoAf4A1IvT3
TtX302kEQGGo4VjdwLUXUiNdPGBmneVkaEEgInkm0zUoBVFd9IRZOHvLWT4nOKS2
bNhfWH96qy7/+MUp3yfjK6HgnRRZETialvnd0xua75hB5fbvODXZ9MhY6K1O9FB3
ZBmFAAJjXJMpB0wM+iDwMfXxDWz58G2B18gxM4yCzrbyOM/fW0XG0U1t/spReuo7
WXYKtSopCevdyY7/wRw3SlzIItnyP5i+7P7h56zEXE+bjtuHMBTP2PMU5+v/iN5s
TNhOSzodYg/VkEK+Way7cmZJq9wVzZJ1WC1b8ChuILY/N+oNBeTwYSEiiOaa4KHU
qsSJnbiJrgEwQ6rH80NBod2CEvp+w6tbcaSPkAkyR5p7QcH/c+TX4ZzzsGnFpUr3
EKSdHS2qgCM5poFaNLCauyTWDN4R58WdccCIArz0DlLL/cRbbyrPrqGzyfvZ63p4
voAfOkPuPkK8cFF2dlteZe8f/bbHnnIqGQ2tacS4sx4rbBWeZWTMerNDIlvuiUqH
2AeCM+FXop+niynvwP7WGi7hF0E2GTU4uBHyaSSn3lt7ppHut7iqCeSR3R3pv0Et
nHhcRXI+0tB+deyfX9I6LKcyhIHRF03/6tE22RcaSILETKhcBSaELQxgW6vTWdqt
vXOeqJpjYj147q9fN6tmTptezm0JXQs9H1guG9oWPeQDM7rpMl1vyjhHf4Ohli0N
lihUMNpwrANjqNihUFPKepWHrSG7Eh+E7A1WL+RLYUKdCtKP04Ry3VvS7W5x4n1u
my/+n9iIsnAMJn3XSRfH56ST+tn7a/35t54F0fvFa4gcnWyQCrdFs2SrH2A8rJ3H
bgyVEwxWyAboHwkTnfIfQR5dls/rRvTBPoZng+Kx/XGsIrFCkc1xuOUQPf37+TtP
i42ybjRVtBeDd1x2uYVVLDLvUWjf1ZuuI8adyX1kBYWFeHRu90pun0xmliAXipVo
qV4+YoBGaxtf75gABbfXpmcq8R+HNKk2dpiInhrd6v2CWMbSVvsEvzhn5N+msPoT
l2e4SOG/SLHD+wnXS9YsozzULHFvPMW031cny9+KzmHr1m6uEaWtZ6kLD8T82sjA
Emi0zTxtCVcmnmuKUZeUj4esRbtULAL8fLRYKaqrURxvu+sFkd1FmjigGXUzho3j
Isid70Bf7MoUtd4z8h4JvxC5BPIUQaiLYYgS2BdeeG86V726lYgm6XE8+i9S134c
v0WcjwpX5Nm0vgOxAzv0BftDyBeDxpMyVs7DP86UDslxw9z5W2UB+BlIsRfhbkcr
NDoRbaWxeSnI9cxXffTFztiuylpyCXWrkwzvl07ZIst2iksbn+E7VAQXSW986Gxl
6P0a8WeL4dJUWdAJZ6N1fnQRC4n+wRqZrPE0loyYVLMgGJHmn70heptBw7eZBT1v
H+HYAoQ2Nutnh1/HBQuuhCQ9tCMh88swxcC2C48t6YmqULTo5THGO1n1TfRWs09N
GiW7MWiygyA8P2tEAUQ21tP0VUBbHWLE8XSKS4QbL/OekX9Si2DUIzCkJpFFKXxY
Jt8ZJGGMqIJ8Otv94RUKT2eqoDP+MxoXFW1IhcFgVYFcfoiyiEkXxGc/y76VkjWX
UZPpnmr9E1yIflFS3Bde8j7dlZtHs9tA0G3DXwWpRiDhk8YTbCIGCiupQrFTBlQX
JngdNL5JbpnKPegBXeLXJfNzsRxXqt/KHNOK0yt5lrMm9kv6FzvIkyNnAV03Wsp8
Lt1klV6TT+DX180M6lCZ0XaBXfjJFD/Hm3nSFme6sBwsS8ZL/De49/rXTuljI7Ml
wqIwJ0GbV3WrfFXNGsUBEbKNg43VmFKCCbwY1egAFflFudGgm420z8QAt6BNScHf
uXE3NZ5ZsLE0oc+UgyQDWJrLRPKYQqziwiMArYottJVhvtP22f41WLOtIx1rD+O6
sKoVjFslm4PCyyFb2k1plu6ScuyMOHxC7ir+zn33CYlyAR9kRA04/X6Bi0jlU9fk
eYldEkGf+uLslarnQJKD7lkFcgJkIfFlQL9Inen5uglHGbZYS5LpeimUZV1Tkef1
C6GOr1N8HUun25JAdys36Kiajg0HvKHRPyeeFk13QHzHj5NfP7FTT/tGtLKCusFa
h3vZ9T/MD2hi/svJQ4DFIp9Qg9psYOSCKthGe9iBK4bRFRHcNU7yssbYqZz3uuME
+EzGSz39oT25zfhFMC7aWeRuO30DcjFpOLbWTgO8WrBAq7cVh7WyfKxbc9YfvNrI
d3PVzxmNUzzOO9KFRcRgn85hdum0kFmBM2/PgXQvsjxLnMiZiiSHsZcyKkYXY3l8
sVMn/HSE6OS/F6YcGekz3c9gQ2Yg0KNHdSdF1b6ULuTsE44UiuVY28Q2BXpWpbVq
IyJrn6cGrCWQ1Hgc0XdAlEWuk7lkqvfDtWaZ26RAnuXD8l1A3KOwCso92E9WBCuP
XufTJ1LwEpZ7gtV6N2oIacGtL2A23jLMZv5eptgzo0/BUPp3C+gVvZzlCLDMKu5z
RjHitvihyqvHilVwL0YUXS/SjL94+YV82tHz9vexfkhe2KA8QPmGtVwcsdmGNWom
pSHtOgX+lUiurrMBVtbzEDJLH10g4TiRCTcRuaEDp52OWfvxZbzE6Gumze/KBjgH
gGtj/q0F+gePeJzShIC6AUcw4NQjDxTKYMj9jSyXc8hm8kDN53qx65xm//cokQeF
B8TsfnEqY1HeIHxOXDRAijelcklWiA7HCzMMFVek1QsBVAU9CVnmtr4F7osf22Fu
wWzHZ4WFbpmJacjMg7bxi5VsQHMrMbXLbM/MsfEsegTVQahxs/eGTJidH9YBpcmv
xy6eThCjzzOAVA/E1je/RZTqE6MB9LzxnINamcaGIjuPskwppRF+LeBo5HxnWtMx
SGv7flAdpAY6JDmhu9v+fm1pxjSY80YWlnlh0WjaZn/7AEYhOtsUcOQ2NtxIQssK
q3haIJBeIGbKWdjR4Fl7hO8l0EDS6NxFckb76AjqNPtkEM8jc3oBkGyRxUTawQLV
NXT/XcceurMZ1j7+r9r/6XZsePQnJnLlORFgC6D6RBvRjHLcfe4GcJGc1u7vsW9J
+zDxPpb2PokAJ9ARWPQZgo2iTeCnTUXTVJEMQPC3bGoL0hWJXTaZrshNQphuBVnq
mJxIxrB2niS3VYaBwWAiAQqVeEZSREjPhUaAI2jvIG0qREO64VPkWvSBI2cp+Vek
gxRLrbkzUNIkg4/WDsl2dNgICaHgdLBRoa1QrY+trAGXF4NyAR1FFNIFfFThRuTR
nL+dscug6OIkere8wEvZdn53eMY+Bj7kuHBeAoIwwMucL+M3iwaStRx9KY+MxeFz
1gPgN6q0pyS7pe8u+AA6v6iIA3uoGWqPmxbc8EW29sGf6w1I/mQKhZzt5k2YCA6d
1m5KEVJ6tDOwyUMKjZlla2wntwg3RpR/c08W7y7nYLj07Y/MzQENh8FAA0KX8B8g
jw+HihrwbLq8G0mczxZfamGZU4ktg3+5LTA4QSPcyQ4kcaV+p9/d96RIaSnLwVB9
6/aKE76npljRmEvtMTzJ/5RQQbMz6VLZtRnzyrUrcDp3lW3SPKuKqeT+hctxyw4x
w9YUQ+V6bnd/QEGhgDZMBJ03B/esvQHFqNDhHOBBgYjo7JzPmZ5op/2QBvJf3m8p
1EIICRaRQCWLIIc7qAAlMEVuOVaRGdvrBU2RhSMTOVHaY3fLGq3hLq3XwBrVEY1A
SfSbO+rKxOTaurH/Oa4aNN9jIS/TqVATORfsunlQqEfGgieXwYVoY1E/OcxQGZpF
JVkyhWwGiF4YtaO2aVAcOm+A+1NVwsZyjYD3TJFF7ETpmvW/ENtGzuubGxziEc2w
oXJ3d+sEeVtA7XNKc45DGfmvA/x9gLw4kTgxLERQ5mUGOlHylWSXRNIuPC0IBt1S
b0w/Tg2UICfNVtA5K3JPWKvGOhDz6A6WXDlR2UWrv9zMmNj9Q+JLvYRDJSYva9Xz
R3CUbSmexf0p8N9f2wcF8beO9+uns+UyYdPCMcsD7D0p6/HZvt0H/CG2z+R4PxDq
byTkyF1qUNM/J34tJtrat0iLgbE5jiwnXBUnOUr5GNjFj9qH3WKINZbqn0LSq4FN
jYuG1N7A44DlRYFqTC59ayzq0LUrfSq8Gkvin2ZTsT4meFBygL4g1EaDFr2iOQLd
5pAg4hYPjSoEpq23npWvQ60QSayXYnkq5nQWETKntQ9ehvrI9TUfSssSM6PANKrX
4al0WATqfWfZAiBhw+nipbKxY3nLU+2oDW02w3vsgyZ+MltXypSF18XhP9ZD1Bmw
c37mAUYX02sGuon32M+KJl8FrWLG/CUnTyd1Huk0t9hGjd5vF6hfAxsVJSDSk0wV
Wc9vxKku6FQ9acCph+/kZqxZVw8mZg7rK6R5BDFlAMyZxQODR7oBBBifeC7UrgRy
nhME5d7UuvA4sy0wc1x2CSEhdzygXE4NGxYZfUsn+3c9U/fBcSdJHfmAVIL218YX
paEqSKpYrgmWY+OQhXbBK1YhDYJioGFZ3P17AMGkQYTF9yunV7WXjLw1I2JUNLXR
PXuCfC91xNulWBKaWEkyh5q6/8ceGp0Oeg1hnSrIAe17dNdRFSefQiTooOsLw68Y
cKm8jNfWOnH/sGENe3tJa5rQUdSoyh0B2UNpfGimmYqhGEwqv99UvSbwyDenDoYk
M/9k903lq8igatCSkWAGM2QRjlRj+qZwENfW2DJX9CU5zNgkoYu+8UbGOuMhjM2R
yAFXb6lDfJDggM3TL/xCnG/C5G/z73I0kEQV/9v6/4ViR/fdsQVCramkQv/I0O4J
VwE6Dx0mLoD0DwdZTFz+NWWw2tG24Vg7dWpvV6ri9cqjiFsv90GkTO4CfIBySNLX
nxauIgl8dW2zF8X0v4eoGolVBVxsOTc+j6YNhNKfwWugwS2d656PJTdJfoHw+TgM
/C6mXhRVLoXfxsPioTe1/NO0jgr8beZZ2poUzJ22bEsDaiip1p8ZNvLt8tbfB20u
Rf3f025ONFWf4b2AoiXl/IhaHEeSMBYWhRBGjRABF2T7Oj8VwBdNxRnAqZvvwqRD
S28l4O9HM5ImLpDc7ZIVto2b3B3YMDS5Xcm+3Cl9JWPUiqSwFDpAnrCrWUjFd5Uu
IHsAHYo1PQ/6W3t6tYMHt4346Q+OFTEqWwg2GBqsVbhy9une0+PyycjAKO56av3U
QZN40z8GoMheXFaeMgLTgbYq8TB6vGjBPEoVb6LwDNbp5Mr3ylCHZ2VJqZ2WWZCD
ULxydGACRjyJW0vkurmMTgV1aXA9oRbsiSG0prz2yxrOlbpwHrGR8q4lcW5q3OyK
U3C7xanUpB1zVR89ckAvFp4gyxlFFbK+trGwH0k946KK4/E9r2tEY52drdSS/2yp
w2i29agmfqV5MBFV0S31ws670Z70o4M9PYTXOzk+AI4dSVFGZOOKLXrkkP50gDn7
+E78Zyh3wEy3vdUYuShgP72ratvOubyX7x+Z4LtWaVZqCL20LY4PVzFCHK1tOYQ0
9e0QgSJ7KlUffyqlbiH8GmcJkXlLK7+OGelZ/TWXw3KOi2PbZuAkNMNulSv+C253
RgM8vyRlt44FruKrekVNcnfHuvfSNHf5OA9FCWCdt1s/4VWAbUcZOft4NFBOO2/7
wPzwNpjn6lpUy4dKyWGbcT/TDwPs8zHVv7qLcX3rgup5CAalsaF00OEoX1H375Sv
0m6rIwxkeiNvRGpGNPt/9/jsbGJbY4ULNXL5GcHO4dYAI2SNpfBrGZ4WaJt0jZZS
WguBfkx1izV01fX5DW7kX7hgrJasruXnbENK5MC+xxesfbaJhmBQERe8JHOFGu6T
OciKaXwQYGltX22wGpxdnbn2t9K3RPdUGoDHyFJEUF/3s1q7Oj294PHnN6lRdfRr
SsU1HoEulBFEVVi0Gnwm+C40WvFYgS8GuC770cgSaMXXlcfISru24GbistjpNURA
cl9dPYXlwu3o1ljFIuQf3wDgt6kD3ZhOEI06ioC9EvjAjxTzkWCwFDquPgphc/p1
rpNBXuUaZ0qMYT792zYe2uD0nUQxv9KaKik9dS8Yiu0qUveWCxfxRemfHBNL/mnI
DO1fxQo/bdZFyiljNYPGKUz2NhxmpKvnVIDPZOT5FxYkgLIqBEBElpoWYLPfpcvh
2GnmR+3q6VrOXImxz+86GIzOeBDB2SPTuFFW1U+5X/RSBYT145Js+WbVMS4Qm7xq
XVdvX58OA39jGnT/P3ItxBb/9+SdREr5x5+vwZJVQpNeKlhOeedpAxA3MJYXVNFY
uRKXwXpXEpishObSmx8kXHDsjDel9ii6MtvDzs5uIBQBHaAyNRVZVpqF6SdRUrJ+
QrJ7zqj4kdpiCVsGdnjKCsYQe0WWkSd64P3jGdvvHXFrXx5QAskrGVT5WKN3QxLS
/jqSlngpEK3E+co9VB12Z+38d1oOtlAv+W3ZXUor4XbqdsICDki1sUY2Ayka189I
1cv0YXyjz/X75qGk4RuaMEqIDuJSdk0HQzyZkSZZhm9rHFsh1RJOTh54Xu7UD3hZ
FuOp4MOL1og9ySimMel4SyX3RADMd/GHSVi11c2Od6n5CmllMQBJ7Jk+G1faL0yY
SYPpqAdc8ifobV+96YH9mmivQdrJd1OVHu1f6IchPIVAx8NFw0XnTVcu4s1ykO/5
DaIOHOt0+ccme775cvkdMr9o7DMgBv0AaKrcxeWsfi4Q+Eb4OQ5A3phUsIeFND3q
K2S737L2Xh/9avno5B244+wrmFq9NHouHM48fivAZQgl1479CwTt//bMOq2OHfn8
lT9o6xTDm9eb8cqPXsX3qqjnIgN3KxDs2KsW7oWfJnwNSLq4faicX43RO6YuE416
i9Q4MsSiZAv+hNVYPofhIpSovse3jRemYlPhp2qDheYwNQ2DmLpKypZHVGq2L551
U5sqmKWKWHMAwr+6Z6mYj2BBKQ75DQPgLYxiyHf4x9d8dTRXaa4wSJ2lS39SkNRp
2NjNGXAj2yRGQjqOdr0kQrmq86/wijorrFBKHRhxKRRrXCTYZWhItfrmMJ0vaSQd
2Tdz924iBvKGLW8eyqwIuIM0MX/Q1qARxOIXlQchOcHjz9OAwa7UgagbMSKXkhHS
PqGcfzmoD3bmx6CML/AnNvMBC8cclDpoWZOwSmC2DQn1sUk92jJ0JkN91rY46vQe
+BylXV2r95bE4dz/nT8BP+zF76fbL8Bao7Vyn/itMM9EyWbH96tZ4wfC5nPSx4ej
84LNS9tLrGlGcwmFNkX9I4PwYtd6kIFVWOPOxFkGfP0XTOAe0k/mIZYWvTUQTiwu
59Cs+uCcTbwvE6MkoS0ERuIcNiv/GFC0pFE6dmw6SpuSrX42F156zFXzDBfastUB
iSu+aw5dOmwgEMDtBLEk0LrLiVUAnmnExo+A+wmRQcEwFoIQYPZ7HdYoEyquK1Oc
6nPjXJJR0cQhqkba1XK6/newuQgLW79cNA2KGdWejnNKM5fZfFGsKWFHjqLr8MZm
85Mrgghdlqbz5vIY52p8CZ1JfsrJDu1c0QK0LDc6gjx/FKahTlqI7ud79f8ruYpQ
RUzOsFOY74DFthKrc+9R560gPgBwgsSMOfsu26m5g9+hwzuZQrlCZE4AJPgHYyRr
wpQRwAAjVIxi9t8PjeuqbTZNLJFUEENyVbYuv6uTR8KultxbCjumlWKaGlI4UYT+
PUIArbwBD+DuDRa0+B79HJKqlwq6HGy6PjSJOpylKVbWPDenutFtuxycC0wsjkwF
i0I1HOhuM0iXeSW5bD41P2/tx24dzwPoULuavLmAb7daN5eoCje4uouao5I1OoDY
wrLA6Zj+aZO1cMiiZDaDAVyAyAyFM7rqnySkBlkvi6pVdj9yZjG0lMHIE4GLr+MU
MqwrWKDfS1u3QEBqN+hmUAZNGiySbReersjjMzQeI5wvSuBF1H8UOI0bYvH5cejW
Y1OZ+G48N1L/9io9kmFjdPZWjFKUSqnRgICP4kBGu1asXnlhDhcg1P11Tb7akKaJ
mmOD0aY3ELjVdjKOJXbTFheX9F1tZqI++xly87w0ibgmJ9lE7vZTG8e/SuSUfrkN
gjx5OwFPJSida8T4/zJ0JJC+BHolMzOVro2Hw+hbKr90VToAlffz8yubMb8Hd12y
S/sguSa3ayZD35WWiiniP0zzn1gn1WiebkNYaxCRep27t/ufT1YfAfBkQy2M6w3a
wr61C20Prd0Wyi7R5y6RqjTY2+/l2hdkwIaQjMVVC0yUyAEY9zt4niFi2S7Hdnsi
Plwc02a96Gwg2a5IWiGYlfV0z+XVqayZ35hvbpMgFrUiLTCbp8Q1NBNiBrknjqtu
Lcw0Gv/xMksF0jo1s/p/6oqHYQN+jMvjCNw0FHIUi1tBr+EYOrkEgPMdJbg9R36b
3ALpT1gfoFWRrM6jCRBvmPJd18/UN662xhPXizMyqLyCRCx3eDseJd0jNst07bSG
hJRmNCM3S3sbNet38w+ZEr5UxsDD7l6jUMolGd0fhKouCS3bgma7H2DyY9moT54v
zn1/1zjl5Uz18sLqeRj4RImhDx+njKCK+2eAGK8/MijyOgeXZCymjJp3YOeR3ntR
Mmb6uFX0QZA0Fy2Hxkc4fp4for3CKw/Q2xF5IJUVxP7bIZT8ijVjV99s4szSgXVM
8PYDPkewFcTLfw15G203VSxuZN1TYiw2OQzOtA/tJKPPe/VrfaJkWyyaYU/Y2Wxx
PEw+KzgkA2nRcPBhmZgSKMtIIyo5stBLDBAgkc1souNEMhB4sfRWjCgi/CY+36ZS
8usglzML3AOFLeWmlCspnwgz6kiBYIkn/9BcjsOhY5mVhb3VrLtYyZWrJOD3dfDo
DW2pj+lzNUeMy4vA1AIZSubwsS0K99SqG4K5h42ljXbINGeQnAUiv7RX1XIYKvOY
spwVjD3/6/GSlz9bL4QEgH2/LxPSlVm5mE9x+r9Eg6QfeLZKIhmc8PrDe38MVI+i
qLr13DWWiPeRFw3g1eSMRZ/Q0x9nx8FEX4Rio9dOwMD4J7vAuHKEQz/owhsP02xm
jVP5nsBRxNP8AqpdXzXUjyK+xOLfVU9OVgBjWkMaRMnZMA7riA9r69wXu2YOVDwb
gDwk7JN0BZgQUVUOV37qlwHmoaKDqUynfDyBieeUkBoyluLvDx17OXL0QFPqUjN8
4TOsExXCCFvbkPphzKnCvjzaM59B786RJnH1zjtL9w4Zny81dq48I/OGJ0XJKYnv
PODAYRcJfR8j5xvzjV3v42o4PKUEneXXZSaDvS4gh4tqguZgWVdzSGWTClHmJOQz
ZqZM9IVJ5BoHChqw08+rE44DyOQ1W38MDqSf/f1NYUeSBH5CzlTf4bNYXVuH9Hs6
/cvAynB8t9lLwX3RK2Rx0BDPDjhUTBQ2cS4JtFcuJv3zCCZDvKXW9H1o2nGILZve
7FdEaDkUWYDtRjA6GMBdP33vWRa7GGnjMXNj7F39TWfOmKKtE3+0NvyDfBFTJNHI
KnH5DCyEoSK6lt0uPi3tB9gDumUVbkQvkCodabFoSrsyTKgZCRtcMfaqH4KOJ02q
EFpK7Ty5O/gH6aVk6VWZrViHSg+MAXaOBNBqCvC+sgmTda9jePHGc6MhYfZw76ir
SFTwlXP9h6mD8TOTpy69X47ppyfuBzg05KAfu6/VWuCYwYKKsk7ETTeGhwniMjpm
tITuBLbIx5PIQ2yZzzU+4ElPKf33GNf0njkjTWwbRvhYs0zErqRg03XirkUaX+cd
9AYdsILTzYF/ojY3DFOmeMNOBdokZS+1tCGGip4OlG4IDvEv31KS0mj9C/lqqVyz
PHuYH799BohVFr37ZKIHqJi6RwdaGfeSZd+QxpeZZ9ZfJ9SihhBjv22HoK/fJxs4
W2OKvmdptAmhu20GRKzb97mBhZJEhqaeArwJIe9KEIRnf7u1ji4DOh7VMqLJfA69
oxrBnh4TeYo5J5/HyHAJAncGQNXcqIbX7bC8bkw0BMqZb/tVkmyIKGHyqZ9ZIRd9
vq3OK+CK1cdv2WnCtgOp1JFIl/vyMMcKPgJ6InpUNcs1fBuq6XVmooujeAK8MBqa
lWvinXEJxynYEBWNF7dqk86XNXYPR3xyFsjnq2YeYPpvKnNXLrOSkfS4iPtI7bnY
hsnk8knzs+tU1UzW1uvzVLEsEWJ1FAdc8JPix6FGBA0OXuEfmwhuZHVeMiA9Cije
uFul5LOUsxJa1sXkXdXy34RLmdPG0msizGJll6h2KrydMhcOZthk8bWJV5MAaR+U
5kuh7jnSJNdLjb5eGIVbRCY3z4OK4I6yV6SPQfJew8HrXmTk4sX93yf99cxfe8B7
1/585dcbM9PyEKxvTOLFMd/bFT/jw3ojvBp53dEwbyad/fG6VCXQVt1aLNOEuUx5
IrsXjgaBe4vVB3FQS8SbknZWs0r5EHnaAkfFoqrGvs/PrUlUZcrMKewqsRZI/2aq
kDziYA0Tg/e1K/OtFiC66dMwHVHZG0fG71hqqArUDwGDfXkeTfh7EyzCSyPBOCF5
K67MSb6P555fMFkfR3cNhKyHcZ/zmdBFyZrc/Y4lm7AdeBVd515Hurw6ZyOgzQYJ
nnDFNlGh95dPirxF4Od077ZOY7Poc9Vy3rvI1oFdJtbJeIuvxGHJ30fF9hLSIo3p
sY4tPwMD49DAH6N5o5IeLGYKGdM9qfhAuady8xmmPvcG1zlbZx7GgUiW1/Sc1Dpb
0kOse8MUjktBy13Uy5pjDvij5BEurAqOthtc2pwayUS7kYd3T9TnSSTzT3OkBydk
pey6imCzkvUoYm7k1nhW2914KEx3dsnAqQBQzkp1Ta76fSShpNhVay/cc7GsZmjt
stzQplegxgl8GwZq85HDgfUWJsOiTGFogIJ4l3Gfhlj3uiNnDIPm+6mWiA14Pa3m
s8HIGIzqL0+sS0W77r2/aUHsyGCaq7/REF0v4Fg7qlmD1Fiz5qacoPlrWCTC/w1U
WSKi/a3PG+A2x3KGRAsqBT0bvQvSDHMz5JPGGV2mmPWVLDDSIjNOWOJUlm/l/la3
VkxBC7QNcFtboULU5KkmHJxNFlazSLsN/oMKX+p2flq8tjnASOZ3Kmc1tvLs21Y3
Soy8Aa6/6Ov3UQl7YQzUEkrUqjEdBB9nyDvi/HtYqviQi0f2xuNk8/dpzUHviMTR
Yym3rfKX67fWjmJFQL/O526eioN+V3PB6llYaRSowk3FAG90n9BXUwaaKYRF+q4n
Ijz0uAQ67fLFZ9LF+4Nnv0V4DJnC2WhxxPgDH2EqGvcPctslK3Y/+S7fMmebwqs9
WDSLOaM5RTNwfibddlJAGOJdKz6LoK/lbvd6e3lgWqI2ivQkblpji0iBhCTDct5D
hePhr25i2JGtXya6Oy7FahGOWyv/lcZEzCu2lsXXeXdy1Mq5DhQmgRcFtFP2sTO7
n+qGvs79QAkOqXlRCXL5mrOcLAQAVC2o5Ev5JWWsstYe6RoCwGgQoxI8dXWTVsk5
+d8ZcnWRbMz9BJjX6IQngQkGS0i7XLxJYtHBbwr1QvzJR2/jNJRQCrPxAhy3N1RY
x6c6F1Jn5m4clRbW7TmPSgQaVIb0Q/z7QjDXaqSeKDDZpnjZBgW8HyzZ4kQy8n1A
dVayCySj8H6Rz/ozJu2amE/AxlQWb2UXsE/BpYhz1bC35RiEf3WMMCWjJ7j+ksW7
rTdPYtUQzyxwJmDpUDiT9rDnAKqRy7LAA8u4ej+YEIJLP+MArJXfKkoJspBdZDUD
xHEUyYbBuBfn/8Erc3kV+TeDbQ6fXCY/3IKUOem2+fvf848oCU3X5qEx5JfMsGK4
Tn7kX/9pMarThWaU8wvXhZKNDwQARCI1zmzmxLC9LsYaDLh73gtqUGXUrVQAzS6T
2yaLrRDANoSNIEuCynk1h7gRBcx7ZzQ12/LH/zy0eUI31q2R5IfJVd6tmCPfshfm
RmW8jC4+QMCroYwV4FGs3J6qshf25GHOzOR43KGwJeFgGgUgWzznEU1T++iWSaCy
fsHZEa7ZOgB8rEIv5eevXeyqrR1ES8EFq4A9Q9NM9GsKbppKF/Cq+e+o6BSKAs3n
xmnkghBuWFODSRuTEyWsIwOqgaEZO22LHDScVYi7aNKMULJMa0G1B5E6aGDATjpt
3BTbG+vaacFqll+wmYmETP4uJaUxFdKCiybLvjclM/I5B1kIIWHfMldlPsTniIwD
VyMHGw4zYjK0pBA5khApqq7T3NxfIcWAGfIVCmP1pD3rkey7NRNe2tEjbI6QF+mY
BBVHZoCZKuVMrvWpU30d3iQ2gKdX+uQCTJHwcnPFcN7Aur5VnmtiKsuFAlwqNrBB
MX3s1Ha0K8bjqQOs1FZNsX/5/kC6VUha3VgSMwz7vfM9SPv2zsiXsDMg/WO9e1jW
JgprNy24KGykd30+bNOm2DvTfKoBSvwd8rbJKOW1duGjBBg1s5rgsMmXa4qW9Rr9
gQQkzReJMad/r630n2AEIKVzxWN3gamH5UvAgEmcrshzcT+Cj5x7dGaTCICE4wsx
ueH/QJKgivIVa/1gz+6Fgw+aMlirrGXTU4g6HFtpHDD/ceZz54+mShQhegoa2PqJ
zbwENpztF46uH2BSeEj6NTftdIjAezemQ7AISmWKeJ3a6D09J8AMMnoIH9v0dZfi
jpoplVCfISaMeOIOE81YzB4fq4oBo/wPOVZ6F/dEt+g3vzmFXPYlBxIRHPInzMY/
UqeUAZ+z2cBJvjBLzu/szgg9FB9YpNBuFhzN6eXMVBrY+wIqyiZLEuqk00ytfXYV
CQBGQa7DWoP7CWcnycm+djRJyyYf+SxGkwiPRhS/pvAMMsaAJ5vAGRSoL87mSanT
bnxXUTwZQRRDS5kViydaMLRqhemL0ENoVGm0TB4wIjZ1n/y4c0ePJ6G99IqW5QfM
AqZNynWwFKNl6bB4UBxfL86jyPW6WhK1+vpHNOgiGB1+aODmVBWRpNziCeN3UVvf
0tLxlR72YfRWmbR1M/qpVO9z2bjGlYWXLfVaJsKMWYmIfF9RCU02oSuoPgIXXGOc
Qo1+/Hym7LHRlKqC9sMMZ9wKT4sXERz7pdCjxWTHGGqjH4/B2ll1YyaN5EpIjTiY
3MXFyDXGt8iNVdH3aRUlW/vQ9meLpCZpewhve4j0FZv6ydcWEHMF5Yk5UCO+iMdy
sLrMaEtlHTh8nEtK/tpRT7DkVYmWqcUTg+jHKwOXc9MufhRfIMg9Y5k6SfC0Vi+b
2/Y/3MEfO1MUsGhRGChNenvIJTNJCgnsmV+J9bz58majuZijkxv1qt0fvqwH+HCJ
390++UZgEAEBqqrrsuvWKRCH+ozm1sY+M9wWlP6UocYbt8wxUBg5OF4fdcX0Xqrr
BV3hlHzjCvVtDHZrVfM9Bzq/DTw6iVYiNOJvacTfaU2xgNglXnQQkJS+j4U/s6JW
n61z7KNuW4y5ZfeMLFeSZgjtsbTfwfXEhGqMuUlBxj9/0kuaiTXhCV4UYa3hsAw7
DPfNDuEzV6/6uXbTHniSmAa4k8dVHsA2ESpA46s3+UY3ZOfi0r/yzF5pKhR0Ac+v
yIBLl6qtzONdwr2eyYEEnWB8fpmSOoV2Z0j2dzyMacsYP7TfuJPZMoTt0zJICZ4r
s6i/eD6bvgGzs9IBiqqnIqa/CcYGN9wo1LogFxCMhO1UpvGoyC6hWVwtJYb21oC5
Pcw8bfb2NBF1XkiBdqfn9ZGTuTj8khawKMrZsa9ARu8WK5nIlwFglZdBW7WWiOgp
5BRobt1WJpqkzKA5MvXy77CxC6QJM1qRkKiScnuO7faCmrCpveRY4ZLhsGJHhJzY
vDavxysOVvypKnG88dr9PHLt4qSOjpWTw9Hl+Sm0M3RCG+fNMrth9xx477HXJMqZ
liCrW7UoZNaZMN7cEDBGgrq65Mf52jIDwwh+/b0ikbgwRdAqHLBooaBK4fEeKBUS
ximObqR0ci0nDs4OM9v+yiD9UQI60rdkBet5bfPCuVUYqllfPYviYaoFyTC2gT4r
SL/ifV+JYJC1wwx8fCDV3lVhcHe/MhLdLKTwmZHX4rf6oPTiXjg8gNk54qM9UR3a
B/NK6/RSGWxSdX0OwNsS/rR7qwSk5TSVf1Bj8GSD/Mhgv+JXF0Ifb5ZtQ90LS9r2
GNJG5bxq/fqfH1SiZhMkcQ19g3uq35wMzmgyYA5T6HbUNJTIACA0IVvm3bq9PKdD
4y0QEHJzRXij5QtjebUcyoEsY4OfqrWGHsfWH9O1gu+Xqz1LYxppnsQvtbXU9139
k2RwEXso9EDfPkSa0maaNYgIoBUDsP3dmWDP6VhS0GFw9TB57qOaobmvwLyLwAgh
L1aWCpIX18G4909n5+sutJk8/avN7/TSpdvZ/AtQ4v3MmHrR0N8vGLSDJvzTutfU
BZ8CRs4JQQ78aplpdOXezTjCF+2FPjmT5Bk0+ZsYQFjRiASBHLxVc8FgOh4iyKZk
+gZqpxlNv2Bf6h+iKG3DoF2OpBnosHLTv2V9hPT0RvMNSap1VYO28lUXAKzOABUu
PDYP7tfNCzwBYYB9yT579FXbnQ4WZvK9APTDhZlXXU7/hYAqgjAObRJw4Jo+d8a0
7DQpqWBhzLY7tf+lKo6F7MD0lLR+3Pg/9Lj2tqylCd+hpLYhIcdikO5EqOYkCxmp
NnpRxJqkGnq3LcZEcF9oYpL+N0OVoxQ4k6+jvQlU12G21WbCnnxEuCZ7BAP2kuRH
zvhAIYOnOGPW37W5ODTpDU1w7VppCmQIuFjOPkMFGW+qMrysaXNkOJV5hF2H7LqV
pC/DHTx4nksbiKTYgan07b+9Db/FJUgYsCZZpfFWEzCCdUP74LpYKj/DD4goy/lA
Kd5kghkMWoB4jPmOmnBuleAoLF7WZrE8475/Qfgjcm9xesoF4uNCgl/S5N3J/URN
+igkqxkvYoGAPEAIzVjB5dailEzvNapbp1q3CDgQpmm3JWifgKed+9YizCWGgkN1
1KCdacOaarcbZpWI1Ymf+NXpUQwI9zE4E1I6hk9fYRJ7fP9XKXF7GOtNawgZhibJ
US+x5fqi0YL8JqcaEE+vxuEANDmB6nKwR2aLMRMBE8BECd9FGUy+kL/JKctgs1CH
lfGF0BGXD/mwDCMCcE/i2SI6IUUlwXiqfv6q7BRQ/kL4lyWrSJWO78/eq7W/6L6j
CzGIKvEI767Em46NcAWX2zDtxuccv4HSu226s4rHQTc9zx0jvmp2EnVGQtMZQ0Ho
6euXABz5neC4aBpy5F+w+nt1bRpAxTY3wSLNMw6+vHu/RHWJZ51QL0KkFwUhETbq
uJbmUoHvCbWmqWcF8BID5XctYHLzVesNPxtrG/klOziOt/rmUgCvnn0LZHVw9ANt
BBxUy5JtfrPIk6R4yt9GTnVSzX/Uqt7AC0VJDNv06NVg5mcvN0/6vQV9veLrR+vj
C738DoXxbY14PYuzzvMPU27mtwNyXBpMU0gaJPXaY0IphP5qzI4v4M/hVu3RyRS0
rrIXHdnqHRtsvYZhUpuSm03/Z/VrsAGgxoLtg0vNViIIqdsG1yZnHcUiJxOrGith
2TrrK/LMXJYzzPYzALXDxF9feTgpECdI22Nw5QisA6ovcpz+xXYUKexOzmZCeeBY
CWgeKDnIOfcmN/Zch1MKwfw6njxZVP1slnTIBVgYBU201pvGQalEoaploiM6znQh
XNmNrFwydxkk7Pv+15uDEUAtgJaZ7trGihCE1YBD3D5utOy6+YbmQ+S7if3plJ3d
M2dXMBFkqk499sy0U6M0Pzp8LA5tp4/ICgTPqnMmtIkic09LGGEqigBtf2qT+dvg
E5zlTjXIq/FCpMAxmiU1hC+lvsY68qpdl+tjOL20MyDuFVSNAVYo3K7ZD1umHF9b
g0WXPdXrM7LYeiXWu7JxACrEcBWTUle8XCgKMWkxsnHgUUZlpvqkCcZKMGCcwkuk
llmTfOrJQK74Q8JgXUttJwWp53bBgNZbcAhLnbkqf+C10M/8dU6We0ppoid44pzY
jnG8Tqwmj6s0Ykh1PbS+uddbdMiG1Kq6RZ017KHdS/L2j1HQFDTsJePeLCJ1ZrFo
oXaK2AKO/UOuXMcCZ81POVks2pfQ/jni11v2gv5Ah9bqtKq/OD/aosuGgfrQTay0
i7dKJSsvjaBrWSEfk1BYI/5EjkzI4/jfPIJUAmT5hZVIOu4EGeK7fqmqFx4T1iN3
vOKMX/muH+67+obHh9lN5KNohLcarJVRUzlXTT6ZAGzNLV/SQTP4FzFMlfoYj81e
YKGQIJJc9TiZMPTXqkHHqbVpiHJH4P3UsJSXtEi5OuLv+990uWr6VCRArD8hMVwT
2EKcZgq/JJJypYgNnRj0eLKlNrIci5VZqPS27lOa5oFx2gwsEugFCqQcekvpriUJ
p/zWqm4xWn6VYrdhhtfewMdWPmeDcsbQ17k3jAEDtt4yLj1cXwWyei4RQqH4xgHX
y9Dr8FEhTa1I7c3QZsXfc0Hskdacuf07SqTWhCpIFp2zNvV8RFE3w6h/NM6D25Ya
nEa9E4pm1LmsaG31AQbsRQE3N+f8Rn2To2XQlpKrIYVhR1qylvKOjkNJHz/TAE3D
lXC8jS3Lj+8kpNJxWOsglOu9QjYYSr3qArLrSHXDZEjlmYa47zI3JVk3KcCBS4YA
PGOHQtG6u1gMctleFnXH681rEUb9dnMeQWVIoMMHV7M/+SjSTGF9sqUaEZNDolYq
wfMiiqQo4MyoOX1njbdeBpukyC+aeRnlnt13PY3XJNkQuIWr2hJGfuou2CiuNKZt
DVMUSnEHc0bHp88fLQlKTfgl9dKyPVzBYAb0u/KzoLGhMgTPxuOhOJqiETGsxCcf
7II3M4mJs7jDNhnme1ZM28C+1ol2FPNqhPRJMqrZi8QVtnFOSjcUNSfOx3unBlYb
3yk66tfrhfK/IM9u5d56ExrYrP6e2o4+0zC8QdyLLYBbYq9xzGfFQvHBGjVRD6Qi
M+tGN+yQ4HWY27fEBcho3BPxzxA2h2yFIjujek3o2vlP0Pls9gdYIWc5fuYcAWU7
EEt5GjehzTqVgqWPV4o137ESJzNh2ehuF1hD9hTyVZHiQu1ayp0ZCET/zdwDbR0J
bhzU/6yocXRANClycIylmJrh4up2G0AebSnjGYhU35orj5b1Xmck5po+755nxL96
WaHE7/DsBqjR8Oghp/VoTfrP+1kppzEFF9h5MZI7vBSst2skNRDKpdmDI1+FKhwc
MM4AuEuVLJhlbLlO5sWX8WNZrqaLsQ8bguVoVr28uDQNe3TMChq+6xzdJQds7UIc
Uir9SvzzwD6GbOhxcNjumJ5k5sms/IO96Gv8CWOKzxYTb4zE2WSSLV+sAoPpamqB
dodkvD4F6GNZ7SZkCAy2Bm80ZmJHWVwL87i8k1WCMdznSe0REPZQd+zjG3QXiFgw
99BOwUjyWd8WO4ILJFmhhpl0CSXtrmLwQ5ab2ILvaHkX+/5MUOz0GfRNzkje7UWZ
h6Oja1RjZjnxA/olCrruiF6vgfwrUGmudX4Z9qjbCvOkLKMuzxFjeyMIZN1w0ojF
EnBflYgjMqK0znHN9vF3kaWBx9ar8Yxo0iOtFKBau4E+pMQyqN83/eKFDzibazqB
E889PmxXq2eEF/JXuRBk9O10X7IS5GHuoskqek9Rg8xssArTlkKNtdXHrTxq6zi3
Bw1dRgaeNZ3/yVRRI083txHPAeP+iBsutf3n1Vseps1c5QbWLO5xLEFJhCaTzVDO
vY/is5hUK33VbwGTtYsQtb/wSA0qwPoVWwR7cuWX9cJS4GpmEp6cT76H8FP9kZx+
Gj/Q2ecPqSgxa/6QAbUL5QLXPTV4w5D7fdGBFf7XiRtujrQBjqc+oe9anBUy2/rH
6DFj14zrP0b9fNbNx8+oKGM1y1BuOeOtXUXXXlVEfIczw7t+ptpzP7WZlirCDX/8
ybI3yYD+8aQ94twGCcyHgJz1Qyaiq/lKSh/Z9hBYRpZh4Q938JPqLDyJYrous9nA
5LDvbavmeN/56pmID1sNZM7M6frEBvwnVN5gYuhizX8rPPr0NfcRsjWUK9MtuDfk
n5UXQKUqL7/C44EaFS+o1LezorrQFLXO+4eflFYsiCBgsQrNinWD6PvylKL2dcIa
s/7z5NRnkhhcc+03b5bTUkKEfoSd2bGcjGZ9pvrzrouAMgME5zlrT8yYGavF7Bte
v3RvuvM8+ibeZvlmkLEkE9MOozEG6CHuZRci1t96NzIWDZIeLnwBXz9EBkbhACbH
XCUsbVMG3i9+W7JLne5ppPMVLyFdyta7kEZadOECWOlap6I3kaA0CHrl5NXh4Y8l
Tmx+UxwvLD/VSrPs17q2lK1Soqbm57QgJFkidxk/cW7TaIISj4/dwRnedBG5RR20
0FlUO6LB+aYAeoL5X4+vicfmuFWWSo05Wj8te/at9Pn8oyV7BiMPtjzawfVAuHCd
IEHr9lgPL8BGw7FrNMsmcITLbvWzVXKc7vnanwg6YNMqMH8TldI98b9K7zLQq+Bf
1bRAwbDAJ/82u8slWjf65smaYcHTYRVh0K/txrB3dlZjk+Shw85UZKH/ya4VruO/
M9zDYLsXiDXfrqpC7kX2Wj0WxCvnl5LVQj/nj2o8YrXQ8C1VAb+aDyAIz10Qp+aV
062Ra5d9suRKUHpO7wOBMF496UBoijIVQ8+vm3g0GzgdiWLrTBVStaIiyEUtslFU
Wtp4K0mr6wCzozZRk743UqL/AN1XwwP4F51qL+BTeX/794MkYYzDHY2dLUlD/jD4
cc+9aunEgHdb5dIhOckx7RzxeQ9uu82qnyhxGcqHqIOGGVOuSDDpeKnncY6wwA0r
jyjSN9NbXHaNJ/X7V4KsFPJ3/Fo0TgMaNd0a+NYXUe//UqCPiTnU0bRjEEQquOUH
omk49zXZt6MKCsQ+hUeHytdLbXHqYeAQBwFQWhhr1SDYQEElhKckJjsXcVVODsyQ
f7k8thzN3fl6XgMhjmkzHwMgjoqxs7zU8TkgW3A1qTMbUBNykJPML1ZVeMqPj+Qt
Us4a/YvGKgVUabm+sh3mDcfKhzK215A3UoprBuFFuP2P5BP93Jk4LDEoZWp7quDl
EPnGbGVLv0TYjuK4q+/cWGebl6SoFivU4m9w8KMVkbFc8qdHKcykw/wDS2L+Xd+Z
wJrVs/m3325YiQkCouClbV1zOW3av7Nb4K1ICccvX/U9UUPPmd7LKrp8Dcoffm2g
GprcycQQHtKV8JvozFgskm7Gm+mRbRQx+iXRyz3DEKkFHlJUmO79pJ1FFmmJEmyn
l6/MWaGZhQPkWzSESDNTpF8gAabuSmkGoqQU00gwGFMYIMeetf6nIV+kASp5NWFk
F2QouqD5Bp01GR5AxyGtAmL0dmtsO8NyvQ8fp8jIq0YxZ5iPoMrt9Xbi3oFML5Y0
xZVBsNKQ9Hpo802zcSVaY6lMYAd+PPYIB1xHoWEQByNDjaLrCWt07ES920fbkWry
DfpqixTzXsyxu4WTFrJPe0SdCCmcj80BSjOGvSH8hYZCC95Xl2fRj+rSxRDEXVAR
HYz7CTYuIGx1hJEunoFCTEOdF2AJ52IjGTJC47Qh066ggk11k1KgRMkaQDIU4hUY
aQv9CFScaqcPhC9uoeh2dkmvzs1ZufYat9sV34zvJMmsh2ViVydagEm317j40ByN
Q10AnajyYu+7e/nvi5ylMicIDy2Ay5n5t/J4/sWSQTHhENzmdYmKecxI380cu+xx
LF0oM8fEfYOuD0PIRiuU+gMbxqrGvFW1bUeapff/gj1naDUCQkMYGWV/28w/uJ4Y
sRDxWCt/l8DNPX3WLQb8Oa4P44WaacqZKqogupyRYKQZBdrTrJBvbDv/IC/uB4nt
wKQZfkfbqf8QtBjTVS4QWfBIhTx/SC159mCg/JEpIwmg9v5EqAFnAmz5jr2cACVN
8QMOKxU7bAxiUkjPURf2LvxrTk79RKICkQ4H2NShusnwUj1VZpefb2kTZlBstGpo
vKy7o2aVRk1i7zbMYQKLDMNY6ouPkqrerliucr+xuf1Q/ewP9ZLAVqtWymMruUHC
nDJJ01qzBEdd6yh7TqklDg6nCr0idIALQ3FYvc2f2uIr+qwoyeatsyO5JeiASuTk
4WV9BW72gn6YuG9HaOqRvpVHoY2NSXS/w/SIXg7JOoCQZC5QMYdDV90rHfnJfVP4
/rgOLBvWLw2Wrwxo8jnvG8u39pGx3UNFzYSZ3ro7YaNMSecD+aRwN1Ww3BUDw1li
qaBIgd4BK2T7QD46e5tZRAQY6YBnWLHOhKazjOKBVffr6nLb8D3XfVkqm3e0EtTf
O09eL1UUhLNa4cRmCa1mL3Qdlb7zfXMVKiBNp9xZmB9bhPRP0VA1oOX+b7LFAXJx
IeVjc8b+mtocTXdDbIoiTGcHM3PtB03a9BOgMLYr+gKSfgbK8/sNTCXXJeZ2TacF
eE8+70rdYcblgfv7TKH56kTHHyzkXJenSEwzlUJtDqIRVgbhpzkrSuuq3rps7KUI
gL7GVl/bqSKTePiE4N0Z7gIo7SnKpDJyQ+ygMdbD7dXeFCk/6z6M+FGlm7cWkfdG
QePegMvJcygmbz8w093xOtggByoS3rRzMbEHdTT0ulcX9g0stSoeahZ3Tuysxa39
dl4VFJ/c81+1L90RQNq+2q/TEO1s/VOU4f8sHmnZruQnO6e1OjxBO1J1UKVpVXJB
cXxDdVMGto5RU3C2q3K1K6VFdwY27IA43/xJLWhQcP0/5kPzRkcxYBtBBn01Ps7S
kEWkiSRLyjS4GD/g5saIgBlqEr+scqU1ew7m3eUAoNHs9dvpqYqg/1RX/Vg8l1Zs
fORiwMUoOw3Tncw2Cw4gwS3QTsFUjQ8hbmVW4Bz21STdIwvInIVxvvxAMGEMYL8d
wUdp8Fr0Fl361ZHyC4DiDnW0YGahuLvPoQNb8l5pFiT0OY7GwD9I3hJx/Uz3KxNk
suqV1DdhGqlmXSn8glIziCuJhCPAT6iRevs3aL/l2TWRHTK4JDhJegq83cLWM5MS
xSyojFmPK9iXLQ8etOEeiv4aUzD83OQu9DQ8wwQ7Tlyd+dgjetbD4egYxr/te6M9
dKKGm3Pz9l6290ierQ3JtFNB9XJERuvT3FW2v7dSiCs/qCN5AOjO1DnPYRYxH3q6
a7luZ8XBSqIeBKxHKDe0eJxy305bfETFLJDk+3ybyybDOCSIZbUlxwP1dqsjrVL3
fl/Tc5Vdd4w2BZIVrvby3UqejarB7nIWl9xSrd0S6t/Nbl/zSzo8REty1Wvf6f3a
q81486OSu76Tx71ZFuXVTekfk3aw73R0wS1hU0mN73/F2dlMK5EIQZiHb+hRXCPe
Mdz6vqoD6a7arbiGD57/zd7Ltnl0IOs5LWxJU++EQ+iu+Ch/hRnfqVKu0U9PTE1x
82ktq1e7s62VlOliqobPGiuDy7Ylne1Pfe50Ayh8I2fH2Ffl/1FJjs/wXe5H2TDv
/ldV5T2+cammW8MfW/97Yx0i7mCg27F1bUqyUshRasynQyE4oBTkGWS1polCYn3C
Q5piTAnswoIXWUj4bFkMRBrqEvBz118VkX+51TyRcs+3KYQeaX1YTMNYSpvrtMp/
WySdBqmrLgjPopCuqIsJU3TNWaRRbHGgRe2WIwUA/l+6OXGUoXtCH+ZcNrO1Es2M
V9xZMirFXuRQS8X58j2nSYuVo5Ca/rCVYKOcbaVmr0IlnFUAWtHW7Rnu5HiH08q/
usoYBcRvkiL5FddjAgp9Y86fShfxMpxtqe+SQZT70bDBdi21eTO2gYRp9kQnduXs
8TL/rZQdV9bqCLMQ1NFOPS7L4EdPfmTueeU1GGUXfrwoxFYiCH6L/46upIdEvTmv
ZC8Drl4tot0t+onXa5BLU9V6PdatZr7uurabNLvGdadGzSfdPrcWlLVxiV1EICRQ
axAi6WFnA0m+F+C0PgEsJOpngGxFWxDOn3AiKJu5OXiQ+CDmXVSVPsjvawtdYMQE
pIOisVi01K1j+QdRC8LhK+WYg5yJcax7tK+6jfHt67VZ8dqN8G9FJo0BUuq/wpA3
rBIrLUJZJt8x0h1eecbegYt5k0gC2Zkv5QnwnHdqunyZG0deJSa6nI81FB6qI/10
dCFbbaJ/0cbT36arJGy+FwmM+moZmMay+DT6sDaareaxx6MscQTe9wMZtuZywmnY
ZqM/i3RbZGoj+5727WOW4U1h5kSyWbTGem7H0hyFBfi+X4Pts1/0Sy4bQ1TCINy5
IdD7TnynOM4pchl7T10eJVImx7R1GDe5rajrrSzgyebM0GTWFo1xXBM2jWjbD+PQ
n57Eld43AbLA5inC25yU9YDSGTg0tVanWDQBrCWN2Zk9EehWAF6SWBEMlgGSxPvM
mWBQ0DEq6mqAEzr66Pcov7I/o4/p1FB6mavBHb6afXAsPtYH+dLIOjBHvYYKShzA
+2Moe2ZbpFt4uomYgM8F7Ac7+guiCJkrpqDEJaa7uR+g+394TCBMcbCaTwIc3khy
USW9E0CZHYfEQ4/QNRLVQlUz3TAC1nkfmX3s2FW9vXHYA3OgqBVBpJcytox4zvDj
ZrtQT/mc6c4oB1M3jNNefTwP0ox+ag7q9Tjt6ksnQ5hHgG28qaM2+zN1C3rgmUiC
dg05pC89KFrCm3UJ3i167kqFlX+FWz7EBn92UwL8g9WdmJZKElZ2/8kJJY0NoiB4
GRDdgJa/FuUYRSAkvcDfd4GiyKz1H7FOi2naFSJcK7TwB8McSITdv6bn6Ncfxmw4
mf6XYaxcwppXfhRMUkq3fZ0qjad8zcw5vY/tz+X3+pJnnDCYteQFxz0bfwmOrfMw
jSMi7QOgITgXBxTRhMU0oscj2jgwGUdF3JXzrwNCbGt5OnaqW+j7B3rJ0aJ20764
MBUuIDH9l5+bWGyH1hajyGOIs9NrVxThmHr7MlOyzCG7qtOmIx0RChkqnvRF1kKD
NuwtXJXZtV87SWkAZ4mEupfutn611g6S9bk/+3DY6K/0d93PLMUJABVRaFZQxhFG
XWacupwLQhXF7QwFq7t0WtZzS+D76+hAIvQkx5JCiNgAjFSADGoqBMRqVCIKEQRl
XklhlsWJJJhXyGvFElHaG2pVuPH/EcbtALd2uSwQ/Yy6UG1jA/+Cs/hU82b7HmRW
eVPLqw5fWnNHi2OGV0TBcVo6y7kKZRWAm0JGMoqnjJJD4yNwNC0JqNDnRRClICYd
zhIvy+N/Tq8YfvSKkb33GIpXKmPrZcr/MiagACL6OGEEInr6Ba4I2/jGVCJU4vP8
L4D6BNSk+NVTmVKapzRrj+XEnEj88oUBGwXvT8VXdiGWvBAO49b3ALBQUBJgf9jX
CrDcnOi62RaNfQD0U/2KuB4Y0hQXFnhMN1QTF1f1AdBOrpDslpTAyaytacgiUtae
HaFQ0ezAebbejkjXemE4rfx+11yL5xhUtM2YNKhQTdXBf5JWTQXhP+q8d7vuz16N
yJ50jpUsf6w8LPdOSmr/gpnT2HilCB97L7gnVtYABTfAI1eyp9UeFpKH80mbfnpb
foMZli8CvetlSZD6yg0dVDK0EAjrJptsN+boWNs9TF8Fg4qCiA28b+pvzBKKfFOi
aQ4TQZhpGQ6fcrJLUKkKto+rIbK/GfD5Fu02hd0BchOwfhqBLhl+4+1D6OZBqDZ3
xwFfNMvEqEtozQAzJw99qDnTkt65eJ8ZfLLGN3/Eb732jWxznMClQZiqI8e4GPjg
wf5UuL9PRzD1PxVBt49ONPuud9mQP9FKfiFnGPKOXAqG6ijCjAXv9Q+7TKo5zmth
JnLso2D2IyMECw/UTod8/Oyt1XgjXuzGNQfUJ4BqQHt0iTfvEGJU2j62/w41s4p2
8VN1wSMV2gh2M9SRcX5I8S3H2Npwv7lQ3W22rvDypFtiJHIO0gqxBDCziiznut86
WerJzYGiUkxlPvEM0DhA3oJdNgDJi1pGaM7CuKRrdYP6ph5HiRQiEaBm1B93zdRo
HE7DTeGO1yt6cvekKOh1JajOIp4ypt3y9PJkOLlFOt/6zlelLerL4s0He+iF8fNj
/PRdldhs1GBsDYB0bifoC5P1uZ4epox+PoJ01yXzDV4IOaGlExYa5DF/5LcWr05U
SmGhWlMjJYvdKW1jdum4shQo3Up8zj1vcYscFGZkrAkcb+P3+5SfO4I7r98u0M4T
4e2Jffp0sfqt405ZAbxDj2x+yEk00spn0EYSmGE47KgTNAM/wIGtDnx3+P2fPmWW
vFYllc+2c+WM9exLXi+LdhfpxJ4b7Ybh3wFpj78htKE0/YV3OKqr5gguzn0+MU5y
ObmejfvaGGeO2EIH8gxLe2B4KL3v61nGfTdKd9XAX+tJTijDIt2yM309GfLMbS4f
gConHKe7DylOIqH2zDgKWxckcHh/Whlly1n/vG9+NumH63FWhvB/lp3EPNAQgS16
jUVUoDumeQJwfvwS3aSeFlsj+nAMfAtuT6wWEEV94Mq48CmcwIzAb0sxeiyMGfs5
k7H3ttsPVRkkdZ0Ni2AHArRdtVUq/CyNcKC3xJ1nn93Ij04UYpofYT61nSAWtj5B
pP+cdNot9Y09ns2MUXXE5zjAB6eULb0jQk3ttn8FMWzpAJ44STttu4LTmFVMU1NP
4pgKCpEYl81Oz5XsMiQ2jR6wh8MeFgvoyrI43cX5pGa0M5gLs4oWewhFenMfwScg
/UQ79U6ABB6qtpam1g3OCOBqsI2A/DnufVwvLjvd6gPAaF5/27JOoC8JKeOxVM/F
rn7IweJipeEz9EWUGITqVcDJ31AbZSaJRrKy93q3gAQnj5kIHi9GWAwnqA1pbMH/
hw8u9h7wUGzLSC5aZuek5H0/hsPmkHmJ2f8cFFrSS1k9rpOzcKfCBoZFd96b6R1J
ic7R8ztjL9qyf6lAO2sL2ul9i3C2PZdJzFg5Rrc2mgOwcdzAjeTaYIf4HJy6+oVm
761LEvU+f7N91TihRUx0v4+quFMZ8IYM7vZFcxqi9YWxcJPuV8jxN6UjzvTmsZvX
xCEu+IKmDBu74MP0RSTDQjjajxDKPIcFgCGsHU7gE2zhu1/kT49ifdtXjyZgcJwh
TnK8tZ+i5Yy41ABtTZlK9pWG3HrhW/eisHHgWcnaF4l2jP8YdkE5PLRcDGpqEla/
KbzyGrOg/BQaZVpUYuDR3Q1l2ZeIHddwcrg30VJVT0PT9cgba3RVt0hTvnBynQiq
TnOlUBmB0hCBYSCXEfKQDLoewuioFWJYCxrRWjRgAl0+5eiera7HjSWvvFf58+DI
T0/z/JnQwtMzAMviF55PCA1urwUGXmoP6cz1ILjAhC9QC+z6MNTDjL2umYRrWUpO
yH66LRyVH0l2NRasxCwy6XkwxrHxHSzonADA7QQJhv8ge0I4tFe8NPPZw55SAfTI
HpOBoEhSH0yTawwtxoDaTkF3npavDjX3Ph2QQXYvGZivtFJagu56/JMSABIMsFAp
vm9LytvJ01CEscbyiqRV/hzooqESUFb8/kgyYg9TArg88IwuK3Ny5km5CL3slvL6
GFuej9y/tx0EDh865ET4Rf9zaCt/1ZaCaS6Y0BTTJWmabrv+SE1nWWpIj/wmryHd
25u5NFaN5HhlG+iVzfmSKQDaON/G+wczbgDDjIdeR78cXB2QdL6gsdUnWOuozAFp
4NLweTCdqBydvjzhYN908pwnmKPAb0oC0+lBTBS1BgtIXLffQuT+e5lG+Z9W0J+q
zheL8ATwle3aEXybjhf7lmfXHCTRi7t9Xr0OxRtPd+0Mfwl4teqiPEDOV7wmqvc/
IoE+GNVAMvq3exCfiHiKxmrtcc3r1myu/l7o2sCJdZEJ95wMiMvkzKysFQidbcuK
VL1o1FVdU5zp1IsDUv3/r+T6ABcqpJ8kTQn7CiTa9gj3/tRLtGaC5GFLUgm9dXC2
pkaGqiIo900fmRISNejR+sw0b6dBzK4ybsRKhda2vPOoJY3ha/AOPAD7IRGWhR5D
O34IfGR90I/83/o20AHGGb8rsY+uv3/wP+rfvRm0jOZXZDUVtx9OXWMS9z67vHEo
ZByT4b8HfDomLBoDndClR6ZM0FqExtKZRqp9d92yptXA3WLH5N7mWuQjxpNRDIhm
DdDzEBUTbLTZnBs/70iNmSXmGC/cC7LdOXxZfNvLWofTsrzzT9Yg2nveQV90ewsQ
uc361H7wl6CT2sOcHZaWy3rsNGfRI6Nko15KFuug0ZDf9TsnEM2wAKkKFcfqrgBX
1PuiWStOZcURy0NUpS+MmJVcZ/PdgTRy4cEKWh1OwfF07eycaynMbBwndb043qGs
0QuSGoCXpGv4kQc8Po1uXYMLAtAddmPUnUd/m95IuudatFLdomWiJfio+pb7gLem
O9UieKv4/O1LgfxwKJugu/aKhEA3JP1vcBTGYs8+ICVoaY19XzUaytS0Y44d+ibs
UL2Waun28BC1Yaff/G6FUvh1rBHl8SYmX5BS4DH2hyTydnmHfMgfbzqom5bbKu3q
Vg9osVuB/a47bYSWDqF1Mlv6sEgFb/aIjP5je6nI3BHQOMHD4U0o+dB5aDAOt/aI
ntB1CqtlVe5UuYmFB5OcxhZ7SfBqRA6P2TeVAmboQNY1boTXWHr24yYwcdVIMgtz
XAwpXPhPNx2WyHhBY8oHcu6MlskyUbBiQjq2Ubwj3swCNXa7XngMX5V7dQ7hcGou
4RE7ySSjz2vgRkLBLo6JRSSDixGC//ihrUqbU4Yuzl6gvNkYxc8PiXBtHiy+gqAW
uwu/2fXmicaSfnoVreQHj6+6OsepXC3L1PWGwsqcU7f4FEU+9wB2CZERKfn7gHVi
8t9z69Z3zVrqrWwh9G8+Y6Hm2gLltWD4xTqfANY7w7Z24Z5uEMapcSlYz0SfSXB+
0ojAlvJTWqNlvm4RuweAc79G2Bj8nCXpND2fZl7i4NinboK7P9a3pYpkko3LczBA
MoUorP02E31+AfN5ICM8QgfnVnmqPAqs49AYOxuYM7A/GT0GBMTzQgAZxuzA44oQ
KIWDWUH2JqtkgTLcrENzk3UEUt6gK7v1LNa839PCNg8ax9YElGuUhStw0KSp+dWx
/p9WKF6nFKE6ingHoaq/wH/Yxhs7zXSvfT2aVfLdSqR5Vy4NaqFSRwOsQX42QzYr
R6Bc+2/FZGdORJGsERpvys5oZxxslkdE185WaENH1qbzNgL4TzmSUVF47QkWdEx7
joulexkgTnVhEyl6bCD0/ETFVbXr26MQJTDg+txFyjd02k5vQ509mxY1cBrQZVw8
hDmu1WfU8BOn4OiIVhRuo0bJ6/lHVvhqBKHo6th6BCDYKl2GaEkBgbzfIwvRwgv4
8wE95XyWvYseZNWPtU6EPGfuy8j7OETP33fcD8CKHn0kP1M9cbTHrEBuwq84zX9Q
0GTMMe9P68h8RAgmU32SSk1HjzLR8ElZeod/+ZkMr2GGBjYuskrrTlsDSJwhDHIA
xAyc08SLEfCXNnyS4GustYbFSHSNF4KiFBYYrBAaKQSFYkJi6BqhmYgpiehld66c
vJoH+ojJqdMMlD8aoGw8DEf1tq7VGJXg6VgIcqBhN3UHRFtUQwokL1kZ0AwB1zZi
oP++uCsUPwdD9J+iRjsnamJrycl95ivncwA5IBGSwXFeOx2y1dtOXybLmWpIBEqd
9OKCZAcNuG6M+Xby2ClBbDDhQd3eOJqSw16ro2HwLgoV5cUg5kMbiFusia7hz875
SbmIy4/yUfTnStHnXV0NpQHMvoE2uZuFI6qgGps11ASHLKf58IZlg5vAAdp494oR
rZdQGof1Ne3B8iLgGoInCjlI8qx1Lt7yfavlavu1CtGSGRTguIYrMEa3aJFeSALc
cJSJEu8f8PoR3e1FwuD0fmwSxKxlMfWQha6ILVdTvVMhcolGJY37io5i4iAfcY8U
dshyQ1LhdOkfXFUpku2ldb4DGhdyDL8DoTePPZ7e1j0ojWqIPZyZiFsXto4+Nafn
LQOYH3WI8XXAhCWziJLcvtTnOzzlsRR2ujYkdkepO+DY0PIhq+oW+EmeGDl/yNNt
de3JreGRB6lU13IdlVRUzo7nRLpHqEG9m7alf5t5oLpLZi2OeOK+RkjRVUGK5HpN
6Q53sZyIlYSdCD7ZC5cTKrC/O8OBMnsMkx5r4wpNddL9m+DSRH0EWbDvJW8edrp/
+TPFLzKMhl+zySHBKo0d4BOCdZhY7yqpLXUlnuFblDhUfzOAf5rO3S11t6sPuwxG
kpdQfJzz6y3fohOySJ/5veFKRAyq98xz7VC6xJ4ZKHyFEdcvwud0gWnFM0dzU4eK
gDt3oWoT0ci0eKBvw4WR4iSGn2s77AnLBxA8p9DyWqJOY8bgaD9VhvdN8G3HPmsm
FBPKlPhFxVIry3LWzbww0eNZGyTG1RGhR0wLgVK2WXIJofojr9MGxAlHk9LV4n1O
ZnoliJ540owvXZAO5a31cVgxlvZAA7z6AJEY+viIlGa8DgVCPhShLB8+AjUyvpbg
Ek0Z9FOo0H1vbUMvgYnhl5HqAdkhaoYoAjB6SmLMQs9qoScDlht8WsDL/6tcfhze
VphkdAblQGnAEflCnau0/0CPagbU0Is+o8IURzAAS2YzJ3c7vmwsHu7nEjRBeqDW
leq0TOYSnAU2hlNI/RLfjbjEo4LcGxJIMUX8gD+iCuCLVbftiAvpVEqGuoQ/NDtL
MXR9w2pzZOrmAZjGMn6qyxjLBZrhwwMHi9/Zf9bC+8jpwkPXftWZ3RUolsWSEzGB
JBKvbyD0zRY8VHRGJNC3lJBIjiAPS3+9pBnPof7oh40PoKTBiLFJwdp6VrIFhjax
CXexnMZU5CohQAYL0j9s/IVw7e1BUMisRXu8q8/MEEn6vJ+QQ4osnhyQGq8QHEQi
9sVE1/d6FayjCOHu84Lputck/I/3CBkSlRWwHaBsl0t8L39Itd8EY/60VBz1OGwT
7cTGPlURSSEaNpLKuvR2/WZIPEqc3+WRbANnfEy4sQQIO2yTArhK0z8lsv4hw1KO
nFYsTDRF38jT1gtLRWPt5MW6bHpGOW525xuhzqeRWi0lyNI87yS1dxhaHxDinXLH
1XiOzupj7p8iKNq37lUts/Jce+sJpw++Onz5464XDHsuUSKEFWWDEE26+2KAkHEn
9kWhTDw6C9ifAjQ6qyBCOrCfXACIYxy+f2iiH9r40tuauP5zFBYAkuSInv1IvyVE
wx//13W8K42Ht1WE6c18iZ2pAHl1M4Rw5KYN6yG5QT0Xsy0OBmFk9TO5hyFs/5WL
6aL8pUDSFmYR8T3obi39xpdR13jURtmfSuEB9vmcOuPF3PvuigBcM5tRs4OeYLZ/
vfuGP3CbtMe53O1BkQ3ISUp5eqiPxWmLzdfvenFyo4OYfg81urIYLpNNH11RkDpi
V/eWKOdrtiszHNmm4kdubuBMM+U8FYSuSGFRTVGPuc2+CfwRj+iO1g+vD5912Pqh
uJ3ucJol9jTq4P5bTCuSd8yDLfc2lgWh3D8snnVxBEbU5gWqn9zGdiysEWR7E17X
qcqjUW9CMM/1U+1pjQSN1oOs1cA+fDodsW2OuFgZBG/APId0O9h3cUPfpADFi3c1
yIkCg0OdAaWAG52nhJcJK13Am8ayy8MVtCQ9sYfY5+0/Pc3JzaN9JPdWEoACoA2Y
OALyKvdS4DKWv58HYC54Y0nPm/YMbAAj4IjX4QR0YQPEp7Y95qwYZ0lPpA+rnPvS
qS3yJHnkWrooSZ/2FdYwvuVs/DA5NvtvBGERQcwykOnbjmuiWgSskQrz5JtSe6ej
tAkWza+6BEwYVPM/HJNqQ4+HYw8gXUwVn167MRsy21V/IiT6tJL10AGc52w+dedc
1AkX7tn5dC2JkbGMWjZl/08vZ37ij9YNIUn6Z541MV8//bJEm9gWSiVpvND2IZGb
A6JKz3W4b/N0NhrI9QLp0JfR1EZjXbsxWxsrhDIwfwAe0+eCCT0Onwr34pMR3w+Z
Qq0Bt4YwVmRIyEneVjHnQwtOETp7K4/fV73jrVlroclRrhEOHOpP8vODVbtyyffd
m0VUQMPdPh2e2oE/uKXbM8P9EmToZUUCj1vnQSnVB7h67zVDUSNBOOIT/G5+U8PQ
qD8pkoexXY+JyMf0VNgDewBPhoi8Aoy86I5YQ1R/s1rIc++zz/Z5nZOTfYXM/1r3
tSOEL/36/Qb6X04uTWfPK/kywYEejhTxrhPpd1ANbnsKdWa4SM3JXGyiEylSQ2cK
wvthZ7NX4QqCwYBNllzkEJH7/p3Yh2YB6C6rn66Hcs6BlFx5+A23CQbvT3rd20UW
Ewfv9k8QIqYs6dZ3sb/1g9PNzUBa8bnIzygTNDvwWU3ksnxFpoz0UL8VYUNQdfG6
fq8itcGLxnOgTCrNN7H3aVzG8K6uL4/fIXX9vuxXlqW49vr3jcS2be+JmOK/ZNlm
Evr06OJfcM/JpxUfYcASmLEbJ4jdy8fHjjKLTBTVN8QRb+RT1u2JEdmMAsf9iNrk
rkUDCuIWmdW34IZFv0qk+a0Dbcx3/0Sd8vfdqFH9mVWlGqLjZh/K6RGpHSTvpMb0
QUw9WTajTouMAYIvUd+2UkHjVAW1fij9/vqlGOzd9wQGpMsmbmkK+vkPF2D+yREe
5TqnJu7MJQqxF+kdWjNmK+/ZS7fa5zqMPVNSBynmPihXJXTAhBVXcHYWwluD28LK
hKlWtJtTmCPLWwJgeV1L0oFHViraI1fT+JK7THoWp9ABR/nXau5l4ldaLCjI8ZJS
hKKxyXzs31isjU33Dt3GzbHaG9D5mV0omna0pvbX563FnbQ60PVq5PQC1f6Rds49
kQv0WBQVfDXGP8rTluI5ilX4oIBCXUu55tUBkVZ84x+ba5F8jB6xjGs2BzR6Joh2
FRwmiIbW0DvF33urPBKvNUyRuiPM85wctSUKgAGhRSaMTZV7X50hFuPIo6VgXnC3
eIGYoFijTxSgNAKvBUfy94yRESB6nxIBHBXdksYDYogl/tTj6kbzVzW8l0J5946Z
dEjHg1TKzKnqFexcCD4Q43LpVfvn6iAmXr0x8y0fAosQf9tLd7r6hOIfuG7e5xYU
h5NoHSSW/shsvEa8TgUvBjmS/biJUD3xOSzAqD0kv7TE1tVPdfyCasyugyESN5uA
vFVYSIdTRmqmha8G85uwr8qG50u2w3VHhNV14dgFKKrPjrPLRCPW3FnmBFtjqUZ/
jG62HJ3HpkmJ1f+A3uWBn6pPI3GICpZrr9Jw5QEMYoi7u622jg9HiMrdql03zP0+
hlhLToqqmzPmO+Wruh0JOJW0WdtEn305YOkTIn1YIgOt6UMOSHCiouNvjVJiCeIT
3fpfAj/nFUCtV9WHqeSp4emknQa/ZjaNaeDD+3Dh8ZQT0OgOjCqDk/gsCysmNx1O
Bs2MI9yWGKQJlcl28K2gPHu413ea6dv4/1ILDuBOsmxEYR3lhsQUX2Cy1eHV9r5Q
HAY/iNo8HS5WuS1LCg7VkNxNN+9v48R8hl5H17yPt5o2VzMy4CHyotFGng9v/38S
4SWFH8wSVCvkNmQv4aqbuwRVEUDj6AI7K73tDFdJpL0ss7YumpVbFnu4zRSPGj39
iKXzSS9DZkEk2VQu54+nzbfthmJknIXpOerYT7avJp1gmQXu0WsfYKA8NfQznmog
cMy5qyaXwPNJqiht/klds7mSnf3w2EqPm0/+GpagV3ywBWnQqiR5+eQso4YI0kYm
wkpiZ4ntyVv6NHiGcdKn2Bo5XuE9LTHXoMG7kqZ59T3BdzT3JqaKWA/LGyGCa2OF
U7TiijUWRvBMUtpyebQ7V288slRGlx0hE2mdnzJi1QrWoyJqSo796y/ICpVTqw99
mx4tnRFR0xYaAn4TbgsQ9lg/sAELHl1vzAt0WCpNLhReOcut7N5F9XRmqYEN74RZ
ANMbRy1lDvWmnZyOYQOdjg8ev/5PezwR5idQ9++d9qb6E8/kp3rHmQOBVydUFTKC
4dNjeylncmSz8SjKLj/NVn6meTmpvDF2r/j5EgMPWgTXHLYQskAHYvanYBNlEGJZ
GntXsohet0U8dXI6u/7MiSk4KcJyOQajITYDCQeB0OCA7dk8XJ4ZUQoGTHcgILGS
3BXkCQJvV7+10YC1OWg0yFtQ7HrHC8GYc4UJ7rGXCAARRawfgGF2X/qjfxV9Oyyj
jGlWQMHDwNYBSNOQjw5/KW+QCc3yQf0vPw0VtzFJ+P1yNkTWDrvb3uWX6/haVLcB
B6OOVA0x4GmzUkfH1yhS4L5dVHLaYyWiF1j+ENkItIV0kysf/nG4QAYGBkaLoxIW
WNNEHiup5obeObHmC1I4s+KZratNKNcBir8LewoesGWs2fz2cBNUfsLoWcy3hxuI
89vAgAGaR7Doy6HWMdd558pKk3tLzZmHpJ0Q1t5O1QsczhHkAV30GO2ZKxSUzuzW
5JXxM7qmziOwVFIUEDHzSK53Pczp15onSD/mV79TslMUazsP3GzAo1Hkilal1Bra
/qM6JyZ7AD6DFByN9SfrusWJVZEKYR5cZ0+zezEwbpr1hgT4ZkTX5xIB7DpIK3d9
cZF7jfaAarTJ0ZGj7iT0yU/TmgjP4zrmLWqZcN8MIYRZAypIToQnKuRUwl68TqGd
B9bmyY2i/FY/9+cCVq87EzHwKWaEG1Wmu7O7/cb+/rOXqY3OnA+TEDtodlOqoeKa
m+88X7vP0nUnEZBwf+RUtRdbr0+IzPUVnMxH5PpbbiwmARjStUXyIKKT+9AslUzk
wbR4MmzxGUeANxGahpvAWSIGXGpX3rZ5Obg2vr4IdPsRFTg2RZbApV1yj9iPel/x
P6CRqjTGmDs9TTeSXEeNGJ7QNvtf15Ulka2QKwet/oVoaRifVXqy9U36vxpZrR0j
xbvtXc4HmIaAUqrUJMjGIfHvYfAJ8aWhJOMjoB9mQcZ+sbeTDRF4BqC2ANE+tMAG
iJCF0FMHqO5lNDEcc+ACa50j267LsBxzb2GMeR0uNl/Wk3Ex1eRAS7Kbm8IVKD15
s1hrmySbOopxZdTbbLyTqZbYPXdtR+BG94y1LFdX3Sg/ypJyKaxl5F4++H0/XxZa
grNZSBa6hzs2ZYoRuJhuDAoiALoVDBd7vTBEszcACBMXkb3RcHPVBO1pkAe8kkJX
pozui5RB3jN7WoQIe8gRIgE+Wk5tBR7T5shzYr2RtLoDnfMA6GevwV9BWwPahIbT
xiF0ahc5DrAix7otA2/uJKo8dBDwr6BXbNV/9YWNDME2L/SXRv8aHfBoz49DFzez
Ins5m6txiuCjJjvrD8yVyS2F+ysj/81LUutJEfwupU6iYVuPcJpXA9QchxoV7/MN
ts+KDYibDxj5Al5Bjv2zMuYd9bFwhMerwgOLuwTWWASg8HF3RXNYX4GRsGZGFUJn
9cP3ba7AxQd20dABcsEpV8Ys0mxXAhQHj/kLNJJCIDcx6lJuu/KCCeID1f0JxDEL
T4ppzbqgXbv73Yq6LaoJln0jueDYV3RC9pB4TcoV0CF3MAlPpzwNgRigmDWTI4iY
7cDKfodZ9GBEwJUGUcPG3PH+v0Yi+lgDxD4Y69MqBhK/0PQWOwb3I1Ik7cA+kjRF
nNB1tnLkAv9LyCA6EsIRvrjDIUfLU4UOMXjGtngF0yRdagE/9y7mbr6ELY6Plhkl
159PsSqwDypDYcEC6w2GoYRU0SmMycZ2UEjPPKgk9TiwA4uw6TB3ZI3u6chXzBmi
bRShztigduF73vHJ5pE8L5MtuEVUrrWGc5dk4iQRi0zPlYiQLFmXPJk9Ax9q9o9y
nl0TTmLkMsYidlDI6JLyg9L8zSh7CqQiQf6kNnHKvzgDlHh4X8imNhvPgD+g4lpD
0iIF2/2DOZGvG+t4dbe5ONN6xp/eUVdh1T9M2l9HUXQtSI/anoac1DH+LLnlJnOW
14tVZ/BDP2/G4LfAwzo+Ppbh7EndLTavuus87LprpJ2hDqKsnc9A+IeauxJmqvQ0
bG+z/kFFCQ4/YYtlhVC2ARztrgVcTDC9YT7ZKrWub5C6gRtNJgvTjqY9MhDw4d2P
zjmDfssqzzvwCo+iRkBw65MI7RfN3KMQtyOqUwD0UMhLnZoqJ3VZxQ3wXtGRM3Xt
0kpvanYTXD67+daCZFtzhDsn0kRNCAJIL0p+bPFMAuaZRkY0bgLDmxkXLpIC+fDs
qA9+ZzHVOuXv+0m+fm+FBO9Lq1mZRGIxnvZbn7p9mG1kSXWq0rldG1gg90BVGD4x
EbDP0Fh32FSlxcVBwkHpg2I+2PfV/Mtc2/CMrw8aG2fKhSjAzW0cb2RPo6ZAAa9Q
zyj/ZMml6oeSpVMSP8qsSPZp7QqZW+4vym5w08nd3KYf/7FHATuJLJq3aoXwB3Xb
C1PnS36j0M8qUTvejsLzC/u30FqbMOgu1MARcRxPSXzgMnJ2WvVQBhCFTOlTiYjk
0iJLbhTa7cw/QpdZJxw6FeVCokLMn67iQG8wUojBxhg11ZeonAWDW5DlZ2DYdWQh
/US0reNBPy/sHWWYh2cyCKt9mEnAdwCOTypKUMuIXKc1O6bSM5bAMmCilnvy1I5T
JjeZM0v/3pgE8Bisp4/y9pYoVi3bFTujH4IghWYkwimXu2rzxdkECPnzaPZ6vMoQ
6/F9m7PucaeBBNdK3/UL5ZMkcErp2tPN+xr6eFfItT6geEovtc03BcQiYNvzJhg+
dAVM4vzJZAm0ejIMk0+QoDF9PIIi8yuv4mR7HkNjaK9mUTi0RvYbrb7VDTfVhbfU
q4WZsc4NPQUqo130PF9sQbWXJLhz1Mqj5+pLTp+pQB6tJ7gGi77nfEAulft5VSBo
K5Fq6Uu7iJrkA83SdzQfLj7f2G3NEF8Tr4qjZ6k2B94BRnSBvAYNy64KojQj24g7
9wRPexbTTMLPBInpV1ob7nzZw/ADOViVGli1bCrndF1hNRCFxi5+DuZ4fDH3UBE3
3AeyZszcuZOBpAOctaKpp5RRIk/Nd3Og7r7PoQNJoA02ImuPrD3BgKs1fI7cw3s3
mZyU8TPFblqgTzFrfhTTEFBiuq0KPDvZKEfUWxCLN+RpTe97wGn1OR5m2ZFDzYw1
OFAHtzvQnz2NetnQk+9ceSl977Q6D0vfLTAs7EOf9AJcJZUfx1Uqn48G7koBYTKo
qXPtHadDZi1SVzauwhsP048bWhKPnH9WpRASKQgmGF1jSm9dlnPMS+mSGrslDqtw
EC73rsq7c4ougcgCJXBaUnv7w1EtluhEjGC3G1W63S2Vt3O6dBjpe0QfHB2kaPaD
HGVVCr+WR4zSU7w3XQkQRvLDzSHRIj41gp8/DRiCjpL/FEY7xzS/WWjMj9ji7rcM
PzQlwOO4JL3MoLK/IK35uC13Pp8UxGgOAJT+ybPWsxnAsEs4ZpQbc0xGzXMCqHiI
tKL4k4rC9Kl2YO2sd5jcuGcijQ4y5SNBL4b/9Tydosrs9IJv9N9hlyTiIGcIX95b
vwGvERUH6WZNS8Un20hZKE7aQw0lL5xNeuvGDYjv+Mdo/8VritnIXGfsRqOjGsNZ
kQCP/qsDcWZsY1WTIdTve6s2dt4194yQM1+T/HxnD+I3O0DBB18Bjergd4Sm6Wx8
5KjDiMYXgj+bMGttAIm+GwFWWftKsPVo0NtJHHHW/SCqkGNCr7/aV5HKMRv+aFdo
VOO2CznDyETZyqhbZSk5YgWcFq0GWN5P2taEr/Pa3a+vA4RotshtKdP/BIizHQeP
VuxzTwndXn32bPFNnYwdihfBp/HPcRuq4qZNkDpREGPHgRY6u+4nC4RxMsI1SS9e
3i7JwnyGKFosM/Fj4TdpX6WeSbLK0ZePSIoNNDc7YDIbmv0DsvgQYIdU5y3rxwuy
ghmHUgaQrkEckHekuz+Xdyk3sDXNj494e6T8o38U/j+B9D8m9dfhhaWSVgTd5u1D
poZi2l6MZMadlNHTINEjmcUQgX4/9lN99STOLzgueGjYSVS1WXTcOEX6l1/QrPgK
30Li63ImLWew6+61RyZVol5+kuiiNXaLUtk++mgE59v+D1/YxsJcUpKRBhTNMz/d
eicAfEFqbMRJQVE8WcJOI7OsbgEjWGwEio5fk61NiQAFJkVbZ7TJsOHhavmx1lxU
yYq0h4ZSMlnq5JG6LnmHnfiuaFY7ELni/gELQ+VPu4kpDW93afFB/Y3dffcTIK71
mwSZypl/V8GRUbeFuynZBXp8jUWTA03WRXiPDfUEjiEuuiTdjSN3ivEYQkZAkmWh
mrAiVnrG1yyyr5cVaSYRgVHCKl+SOGYrFl0m65SrI72XnFAtKveaVEogp5bAgKkx
o3829WgPA0E+sY8NDYqcmy1a0HyUUtfTAXiKpu6oOEeK3Fl8fDThLRCc37FHA38C
Hb5At50ZdcQTSPIeNquOQX9dumDoX6kZxfTZejWMX4PFwhS/wTObkGiXO51GN40g
Ea8/D/h0i9QjyEPPw9BW6YHc6kkKAa9ZcDXeRy+tjSbE9Gd1uPWLXljZPaI7fDwR
1Qpg4XUQxGGjdhSD2PKfPF6Gl0/LSjBsB6aqyervt0LIn6LO/k2rsmdSBAtwJBg4
kk8vZnrpddOSIDAXuvQda6x6bMwCbqel2Gmk364y2HcPGazlRnOLaKfjiYIOziWB
GhD9oZhmxXCIUDTNoy5zoPBWbfp+QAoq7wXeNXPhX/gIRupkjD6QOPwZ2IYk0ofW
hxhD3wiZykMQGloQmSIhUUOmx+iJAUZgxklX5g3QLImnvvEgeueeUFuwP3VoQoH+
ZKJo8PH57+joVg6xCJfPEge80bsmecxij8wRwoRgG4M8UqGcY3sQn+FzM4GjY1fR
0UPsdvDk7SAzOt4yWf/9q+NfFFSNJeH6xfFwgtDhDkavRv02YqR4Y2laNpehU02a
MU0s2sxmEzgwm8Gan6cP2BhlCjq9swRdsvc5GLVNCrO0DXsYNrRna3NvGKrDOcFD
h/rexXUzzOeuOzEnBHQrowRE9qQsngt6ybd+yukshdJUpdnpq/oLV+WiCFsAdLva
F+FOhVHMeqOFfkXb8nStPuB6fluGXx3NCcHa7+/l1RKO6iqEC9Z6bB0BKp45G2NK
8eB1UppgEbkFcB+SDx0Yev/GDzSUEkjJyiUsfm22fEtygtCkhwb/bwHSerGjcROz
fJiCjDrEhFFG5alIgr4JZVrHLTmEvEdpLciEviZmuXfwe2R2YhiNbNDG4ki+j+T7
KgPpWPCscRA+vtSTw5/hHiPkbZGFyx51VAdMhxtZIAJGQ7ezULTBwMQOdSWXFmS0
wJ5FT3N2oEWHfZs47o7xNzXTuoWzwLYkYM1OR26LV+HvUu+7dnapQa9r6koD+/qv
cBj3UvlTx/h1lLg2sSdFRYtFsnT4tnHOXgtHS0U4BAfzxjp0Dhe+g4rPaBbjLoE2
tZ3BE5rKZb/QMP/3q7tB/J2HGmyR4MPw9I5rqyCl0dW2RBD1vZR/kL0OD0P4CZop
iPh0DqZas6INqh7TdPyI7wiEviBagYm/2EindmZismbb5VileIRFj3ixKwLBnXd7
826J1TNb1/5ANk8yD2dA1A75lh4Le4RdxP8oeHWOh1tS9AgdqkFAb4H8Rf1Rl8r3
aJuIjCgg8Vz+yL0ufKN+yXRT5yUmF6X5dXoINTwbSQI12F+Vo3UxvBFgRb6Z1O+E
cpXp4LLbksuXj5C5xkZFgFMcUU5SWS3Vh/UaQI46VTjzmi/MiQNhM7DoYAjQVERS
yYsmgQc2aOavF/tnpIjWj3WsIbo38TpRiAWRHCyhAoLHngtyLUcdbevjlrNJpAjw
qqrtx5YUqoiCST4Nqx5jIeobPjNPryFhGMv02nRuhw8Ga1h7N7IFH40TBJtIe+gP
QQ1uUcGT7WShIagah8ulABI38J2m+9xXA4vbjJvUQTxSGHsrBiEJmAhrqYU4VvVd
m9YvqmxoRM9Ga0jmcEH3DtFhVdQ11nnID8q823qOLRg5Yp4++rbDAt8cY9VYPSl+
nZBBiRPKYGedWndOTMB2h3Cru5UQYGjkiwjnih571rBuUhMDuhxWN5TqZdDpw08Y
An7so2flm//hd+CDOQFsDdwXWOC2IxNsWmsAolhmVzv8eXOIzQlNeph9pwR1daHx
RhXrKYLA+utGmu/Gx92fOZUi7eg80lOuubnLCRtXNC43SDN+7up6z4GcbYY+4EZ1
RlFbFTZ9NjzM8I/FOHY9NLpAmlue6aMLssuPvWpRwiVRvtRNyQtUPuGs4xJu5XBw
2rSc1SdKZnqiOR9O12oQAjTqACJ0s2EWv1Kt1gC+v6U6smK1AFEJMSFQ5L53e6lw
PEkhxmr58gui4ckEVQadNsuR0rXzJt88ugIEgaLOyzTe5asryVRObeM9V9Iw39OB
5sCGZ4tX3NoXWkI7NdcnZ2i4w/qoN4DgkSH/2VoOd1pXYdWum4BtIr3zbuHoY0B4
+IoS688Qw2/1ikR1aTypOV/sUeadJoH+4N7XmwndMPLdRd01zgyCLGBa5L00LadE
OCsvsC5WJIEbYuQe/iw032dF72cG25UFqGxDlDHRTq4Nm1www+Y/pCfSMv9tS4Lj
cD2M1oEnQDk5QI5Iez/U0VgM0TfxAiGYISWoXPnJXUFpfuZoX32bRfJQgNu7Swoe
/2X0qRBHFfDnHyjq9g5uavYLATp4IeqtATPgVeSegyBmeMtNXUbMc+kg/DCnXPJD
+CfvuOXT16h3p3prQs+OavWHAHAbkZWM0F1ii6WUP/Ud0eT+kUiZZGNYUwUW/1N2
6mF2YYd1ewTET8D8CpdLMvtMTIldHp1bsG3nQh0u3til4L7CIN+yttMycaEBQFf+
qZVuSmGXr+VQzMhkFi3GMILthtf54PtCnUj+SQsMDaDUj5vbcSYYAOc8W5OOSKl3
F6tkXJReGi2pQx+R9X6lBDHRr4wIe6SnpzIEoSWBuNhZEMbF45pL2z2Kemi3tpaL
gA1TiMWg0phf2MMmKpKMVw04feQX3XiT9MgbzyYOuZpRBFqgRiAQuHWddkoAEto6
PewZ8g9Y5qhFpjVdRwptfJlf4/IilSMVZJzeiq0WKbkAG+iSaEDkaIjANmdqJpsF
tz7bbpl9SdgAmX4x+WAjJGAg4bqBeH3nGhqDQP//c/RMdQQroeSK3p7iaT3/MBAx
+XU66UP6Xz/g7krNm0TcwUDSVAhbjIzY3/4KjQIwPXK/cv99P9lo8F4VyaZP9OGv
UdN98TesjYLUFThB01OotMvs6j0C9nSw05v7Jf5a2eB34JlElIAnBP9XZbf6NQ92
MHKqhlGKgPruUDmLDK6gAiQXmEKh81GmMA4Izoi8NYj9v0eXKK0w7UdolyPQyGA3
hLl+Z5d/vwJ1P6halOma6PMIGT+2XSyRi/va3S7gdpdPP0ub+9B2T9YxqpC43eu0
DJZdp3UEFAl1nfHuJU93hw7boMfQ13faYo/PrD73gOs3Vqe18EuMO0OniSBNmkf1
W1lMCl+CRcP19US0BvTTUWbxU3Yh5uIT6uE3z6VB2RHOqqLIy1rWwPkY0XudrKJ7
Xs+lwJiBSkgl5TIBdxZ9M+XNxJjRupZg3DVcFun19aUa3SpMIE1MVej8daqj9mUA
tOtul1B/WYcn3BXqryk9kwJPwqUX9vOxRLoVQ11exljwbQp0hFoEfTgqTE3HOLsU
XFGtUa3wubRyjMwtDxGiQj2FnA1tYXv6yPdiExctubAeMS7AKvAM+9U1OHE2k4+7
6TYYnpd7teBFvbjd4smpSIo84/mVZyXDlrrJ7p5m6rumtJHUVmOdAht79aYfmEEj
BA5KB1gP7gk1EwdkiIXCVnDPOzWvT11CcvuLnVMVOmR1VjHmbdcfyCV3ayBQdwmy
u5qq9zEP3ACNaakXaLCVmp+FWVkCrswjrNhz7XtHtjQOfbyTOB7AvKTPCpcmXoSE
NMSeh6jpWQGpXhc0RZAbz7Xh0RohfT6+7khhCi4kliX1UBzJaKXqd9bR0jvKp4yH
eMb9Q9UzKaEGhJn9zJEg1hxppPm1NOZmiU0UufKPx6ur6i8PDTm3VcqxCGZEGKjH
hj+d/IoOsW1OqBEVkUoxUxObIOjfVpQvcNZ85pgPBYEesrEquu0hJnI5UINBr0JR
253ZBur8pnpukoa/KtMwEdftW2iK0dC7oNJia73toqmB1V5FVb+olOwbVo6MY6Xk
TMil89WgUx3t2BuaRZKEf92BS5MT5gRHr8f7AgvDPi/zuuSUQV29tnAB4pCcvSEU
vcCSVt90+FZ/Fdw9nb/AD6scr+BkPZ868gzv4W99x6zvQvzRkXCiSWoZtmfg5g6r
H82qsUiKVkUE/1mFdclmhHBeGylmb1OKkayTAH6vW3kutRpt3PQJpDL+ws2OGmu/
AhorcPYVUEjyMeqWJEx2p2pK8y5aejCZE6hT0Xrz9ucXS/V6Lf0U6Z06rUkKfwIJ
uUUexNL1YoGZuj37UutxT8kX6Hwl5qHh/e1rK3ISQj2XEqv9J9p26cetV6DFOdf7
gdj0KQPa+i/aobnpU/92SLUCRilXWqrq5qA7vNpKnfHTYjvzCIsAKTUsKNSdyfEj
9s4j1CQF06Ian/jqsLI7LwDekNu41WTp4Ma9fGi+cQ2uvQFPRhV5ynK6pAFwkOMa
jUCdsiiuZRI2g01uRu7Cn9iD0aqTsOanBN261olaoQJMABoJY9cSt6few8x+d7PX
MV7Yp5q2d/fUrUxtSUsjcPIS+IVGTquQeDBxGOfJYocwgjxWCiD3AynjHKjWr3An
VjeRpmtBiMNq/tBtvhkp6G9NYmWyhayvad4GiJGUvFR5zkVD3oi1ADYMzp1KrjIN
C1yxdXvk6Q8JTuCMUHWY5V9dIf8HH3DOz1tcXc853RRfZevZhlR80BnL4DWo0hnW
ftcZYm2g8cQeX1BUq+m03nmippYAlh2NenbXsg3rt2mWq37sEfHRXPQc+K/XwvIv
wTrI5Ie6SlD88HkNhNBa7nklia44N4GTWYQk7aKCUNEGB5ElBy+NtBqd1/MVC+WQ
o+rGLIMp8aD+gGX0DD1+Ll43YKwQVkw5l4qwFfePG/Lzbr1rk8k0QNxM6BRgPmq9
RTj9hW0zrfWQd3vITDb+FGaGx2SSGLmt/Hv4FD55op5/EO0O2VOFZfVadG/AZ4y3
UxYpWkLNIcE4vl4mClIpIggQKaLaimmA9VlK1qpcKT9NCQ9UZv2IChL2toQg5bjC
3s3sGqCz3qwOqMDT95HfqYDzg8EigNk5ze9/3W+MfZ8dywzqzX9wGt4caTUbnnu4
HyoDsbGMzCt7O71PvNaVFPwCS3/ekj/amBXAWT7BsSehMqSznGL0y2+JSnsNgHV0
E1EJcZsNxRfuMgNtOUvLjFpapKeSDINse+qTQby2cm6k6h7E63f3/fgoNv66/5kp
S4r88aInk/sNhUC2qOCAMaMnvvBMyBwRjkAqv+N/WSwnlNottat81aYbAAYK8yVi
r2MTenqELKmkT72cctCjr4GyHCDpMK3Sv31XYh6q8HjW3xwD2awDURaR/7UOQ20a
4+XiuOwCtPtPpHGkToHnw84/D6umGl8qQ5O/ss7fYytxBzPmR10nl/N1+ATGWeID
sDxxiSy5eb1x22iTbNf5a4XefBM1Em9VuI50wHff84e8jiQxFYDW92iYRT8qkigs
2SwF872KHi/qInjyhUjAwwpUGWK5RltGbbWJ96ol7PA8X0a/QbFtp8XCp87VIW+M
qjqJZSJTxBxvUVN04fchLjGL5GSYjyEYNoWQ5L+tGSl3Rag6xRkdzELJNCkYnBRa
I2UjCtdPQeBWT5Nzip0V88vFLT21rLYd0KTqn3kI90sszP4EVRb9/OF/Q3/KX6jX
F0JK1OMQ49BlqhqVMiciEpQ00sdy5z2nlg6OvEZJhd6CappPq9AWF+Ub6mOwPpWT
fTQG96+ESoRnzIwW/JCXEN5vf77JGhjz759CbSUtOhNiWOfOo4cQzF7NYf/Cj0b0
lPEjaE6wfFGZNgUxxDY4QyT8SAizsO7ObmcCZ6+DhPBBff3z9Ccbb9TYc9cRn1Ri
iGLX9xKr9GSg34ZUKe5kLf4gwf/gBHg+h2fuV1dBCeir+WwI9XsSFmuc/P87oS9K
VcuuL0FV/iZMJgn9SZ+Ujk7doNZMrs3WTTxY32M+BwephvPVwn3KkbsP1nhNcXfN
TpfUhsgFq2/lgio3q+08X9A6dN44r0XO4hk+XkOk1WMB5HvA8+hrh8HUsqwtL9+l
8pCgGg4mJjI+x7RMJZz4Iur7rcxp8Ctrr4o5ZSEA2tp3Nih0oiVwibMTV88s7ZS5
X8mmb3HQSiEt6WlXVPNaj9OL0P1HrWRoPC4D8PclZTQAIauRDoex0CtAra3OrKzP
Dm8cT/zPoU74S5ZhfGnVcS4rPMJLu1V7uWO08Regr5w2gNZgd4pCTUE18d5nJMXZ
eqk6GXmLk9KVO8ZMgqAMncnsUyePuPgx1u9mfhfALe/yeQteaqCs7mmYgVPN1zfP
SXBg5TqSOC9GENVC/RMRImULd5FmCBfkdIGRi3ohuE52hMLV9WWrbwgh0S2GEcV6
l/SfJWPL7yW9VmkZEmMW6FSc1TceIQXQdQ93Y3rnimh5XJDcXjOK15EaVAl7TlFV
tDGOr9fgY1hMyszJRtUVYlFFFKopbiB6K5fUBRuEvr+7rh80N0ZH4p5TB0y2/UUH
UALAAnviCKUfaaxzVKX+Q/sJESJDDpMg0Tz1RS6SxlULefOKHN0h24Y/mLGBQtPD
U5/gu50eNANJOd2Eko+/xc584U2HVY6yqeuIZWhKhBaEYx6XZ3C7ABWodyxenG/k
4RTh2xBne5saQGSBK+gCIExck7XI7JuGb7/YnAcDz1RqJyRexH8n8gsMaA7pKT8x
uigwrJiVnVVIiUkkHUoFHBXwUxNX8x0ucFY9u3cb+npZedF84eCpm6gMEk8vtKwo
Ukbgtm0PzeILGk28RKAb1fUEmwRtca70Tvi8j//532toCqSVitLWLkiD6/uvS4jK
YAp6p5j7/5EE8ku0HTdjKLYW32pAoNeDQEiegoeHwpq2hysHch8xW9rD70CzIpGL
Mc9EqEC1ctv7/w1qlPk1YoyojBAreT0FDQiW7yIgXnOvlMWs1xzO/xLrtyjaZad7
Xvross1Y/LNt9mXNV7/W5MrzmFGXQKAWEo0gRBbUuP9z5upn8Bu+uSM5FDqOT3T8
JS8dSwwjw9jIN0SK/MLiZzkuhGiIjDTWoWKNLHd0FmFIJAmQOJgb96DxKxZHsnwW
JQ8EM1qixoCRm+NvMlZjG4JCyrZMeIfbmcOPFUlJsd/RORUFvHVV/ckujcl/Z22I
ZL13VKx69+x0WQ2OmszN+pcBsTDvfDYiWyM/i53OXHBeJ6NiOFHalw6FnS/makOr
hDfTUY7G2qGztVW4Fn7XPof5vSNke2pZtGlBk5rw6B1mDsze18D4wcr4ZFuB3COC
7Bq4BaqSyjYfU8g9z7HROEVlV5ltcoF5/DAcmqXbRdP8H4UnnNBl3FpA8Iy9yoW3
FURS8DxhMYEceFgdZ0fm32BWgitZ+PSx/MkCq+xVSBOcKFrAxRPEN4B8vTWHvM3N
jVI8+Dan3AH2EEedundnge7sCd8O9bs0DDuhNGhfoRgLN/JjR2JkNsJiQsZuL/tI
emiXwnWJdftbtUvGhU7ujD6NyRNoGTOy8tZ4sK3xThjehS968jP7YwjACphZmQ9r
IQb/18gybv4WyY/+pl/GXHzPzWsKCSM4VYToeWgJ8ZEKDkNabGRT4nVAzXCINzZV
LllbmZP8faBFpp1gjUwgaJgzdDZDl0NOoBT1z3jJp7AORqCgcAecChaT/PDse3rV
VeBv3rTmWFhG/dHqG5mK+bmtBe4MQxTxtknJw5Yalx71EKpIfev9FzJPKc4B6cFs
LU9aSWE2oiTCnRFmHaIgoxtBHjgqZBrW/0A6uZFsCshsKes1q5rX3lx9GAmizpLP
/7ZdVf4a0mlU5ladJWv3d+LKGkzmShDJGps9t+XiH3h6Va0nUdFDQ5OCbNq6TW7O
w2nF3jL5L81tQd4wE7S36doGv+5mE4ns77TAAM139wX6RmJg8gNcVQ8wEslSPqEI
3U/PgIUn9GIkc2bQ0gJLhHU5bBj5wYAC/M4Q/TjL4vsN8sT8u6dywhLg6oaNzdgh
MCYCJveATZDADgq7/wYTTyVOm2GKcMXY6AqxEMNjQ6KuQdnyIx5jOM2hzhL2Z/4R
U+Se6Pk950tVKLtmesRSR8dv0eX7I0JRg1YwYWjackeGwu5QzxyrDW53413rpHbk
YwGCc0M6phveYG7qOgWY0zDn8tsPYK2MBgpHW2kaCOuj372f5Aular+sr9EleHwm
TFQMCbKfyjL0rWyAZHfUqkxZtm/uGPx6dMF5zO82j3ssP0ncGJoNfiqcI59dXPGf
GWGc6XL6m6bgo61WotDhC+A6rD05p07vJMhxRvjVzIsHmRW5dDPX491AA8dIMon1
eROISrSjGEZCbkvroj01MlEbYGEvQOCpAAPgGd/aAGotUWHz+2YETypCsDANv/2y
9XjHKE0039AXoHxlamAro7F8+p6arO5McqjIo6zhSPr+Tn3JiwkXFwBcoJNd8nom
+H19omyiKzEosD2QBjWZS5XZoo2NXyQ/yGqZIQQf2iv4Jty4evAB74S1U5PMsuwZ
YSFCxDDo03Q6bvRvyDNqYuT1d610HEUc5DDOqqWw5Um834VJI5dphgLZrvcbXags
ZjfI3dBmbLD0wY9be1jMCJjnrrLCzyENkmDLItUm5kcJmt1OX9mgUqNBWfsb4lxy
ypa0Tmivivcup1ZoWiC+LD7xlVn/+xm1Bz7Pg3hEI6ZutBniFfTCuaH03oIs7VXa
pSd0nh910M+My500+7ryPwY96OL1gc3ZhKVkV1x09zkz8UVstHrbODoYdCnLzuxl
AxAgaWyRIpV5uKH/8iVdxRJZU7iQnLiILfNsRhYRBEIYPwBnc6w5TU4wAtpfzLBY
VD4Y7RFfRq5B/jHkcQpQpUemaHYcSV796CCt7j2ddn8yJlsU8T5ZsMXU1xUu9ESB
6dBz7tShZj+hiNLAbXbkTMoXHLr+/Nkd4R44Ci3wcWSsFpFJuZ42/oitHHQILcix
F1qm6iYb+nk4DJDB7aUbkexPkomv1Np1CiitJxQdF7SSc/6xPt922QpWQS9KHV3L
Iw+EyZB+5BANoBcsF3MoF2om4O3huBhNmg0CyQ6rh7Hjjdeqm9GIsAJq0kd0/GNM
XaT55mKc57MLeLTDbFakMiAIlaFgl2I/BqwhE6Fcc2qLH0I4Ig7/EL+6m61lG943
oPvEbGtAQeRQz30Y6tE94kBUtFTsiIzf/xs22P1Xc1k6R/d66fdIGVdwupiNKGvn
lbZpiYO3s7H3fGBSgllDiSi/NKPIPkoYTyhSIvPdO+M26StwylKlQRBCtm6OQV5w
1wVSxIUhStpf7AXjaW+m8eWmaVk8vR+LFlB9dt4j1/yau9p3/oJYRahTzfs/79Sp
0JSDCXC7bpjUr8LyWI9t6N1UeHAegcxpw4jwx1CJRf6hjLjzIQVs9mpBlSnx4osk
0gYOGZBFDJM96ZWl8Rr2brBYDP7OdSH6oGRKuKgNeBgY/KsO5XtoqfEfEmWUF2y/
2VMLQZ+1akCyOws1EcaWgxZNwnO98mFNfxEVl1n9OTgpUp0qtu1AhnEI4v+S41Ur
WGcc+Giz/LjwZ0b0aKP8j5mJZ9/1QVFJCtWHO+/UX2pPQujMSUF5wsoToUZUQ0KU
0cx9BEN+31LyyssoGR9K4IlX8dU4ffbfoGzuF9lBr21YccIvmay+y0X8zlzvALcw
/istk4+mWEyE1wv4Sfgw8gNadWQgCWUfHLXwUrH3A27t8H5TYTxwCl6ewG9yMo3p
wGqpFjRTMMC3fs4+RbBRA8isapUkLoEOTSV96rUel90QwE5ogwE2Md2cppxYfDO4
+5EMBQLHUl7v1Y0whZQff7wLC98UjsBuqYbt+KcEmQj4vgYPq4j1F6ERRR0fiUpL
UsMlqWJSjTs7TKclekBzSq+5uL7z8KOXTrG5y4DApGoXCe185VdbbWwdJ1+uBc+/
WlafVSCAQ2WrLLrVLnuIjsa1Dhg8Mv6uXJUZwIaHOFQ/DT7/qD7LJJ01meO7oPEV
DHCWikbOJ/ZFIpr+p0ctFUmyeeYBq6gT6MUO7lezvV07Gb4IqL7ScwrVKfMRk/dF
fZVnI7r1SnxcpI5LMEwZPdSurLK6A2PtIlUdrWL0DalAcIevxIw8L57hZxc/vMK6
LBvDm3bO0xqR2tLjlBIPOAibVuqYLTwU9Bo6dW4hmvi20f4NsjJm0IwkbjqDn7hV
kBaWbkbyXdseAkuNEmHHuYIdFA9Cp8IFG9dCPLhm+2Lmoc07ZD98rfr1Px6m9VXL
+w+jTK5sdsmOgWvUQInPA73DZdqFsCf1Lld6vE+OCIkXPs4ABg8GugO+Lz/lBsIr
zOqC7y7pGmRf/iE5erZxhsyW2ZuXjD8+/54FRF6wm1Zsq+gsX+k4bxwcWveT2HZI
ZsrYmrYQRdBALh9Pm2mXDhXQ5e8fFBdPf+aTar/7T4QcriHNiCaesKmRa8egvEOV
YLdFzLnpO836Wt4rwbdAAxnMmN+qQIiZbOpXGGLlGy6gr3t348fLh6xBzRyn3n03
0pSwJjPPWs/0ezPFLeXLCLFO6peMpQwAp3fyahwmehmRhD5O+sI5yKS1dSLgHFW5
T0OB+wLhvWyQnZyq73bJ2UAcXYNinUpP46rCzrTiin9LTYwvm4IGqhzrkeSxNCX8
r1iRvP25QnHT1E5SqcftvKjg0M/PZ8ryJpFV8V5Xst14mHMWAyJOSvFqY0S1aNa/
Yueuhqlq+MHx4wkjTrQt5jCV0yT5E4odVEa77m4dGXNJ0AXN29EyYy9QtytXB2Du
WHNrU7AhGQNd5mf5s/CnF8svKePFe9be+OVjo8ZYF6ncp57x6FqnagKGIb/cG5lf
WsCJb88Y0V2yA6T+AlIqDFeuek3BEsAOo+V7ZzPWjyKtJQ62xa4OI62F/mL9w3rf
fYgQjg4c6qGz4TaDqiqDn2ju3WB6mAaPE7a4ijIcrKlMukGVjhUd5Q202o1b9WTD
NtDLZNboIrULD4Gz/R5dNMBnyQW+1Pxc5uZt2eVU9Umr0JtFIWLipNpTrqto6BAj
xqvEqquwEQ7Q+BvKE/nZDrOyfrXR8e0+AVIwknfnXZADrSX2uPSD7siTU1QGUkdP
XSUo5DAQR/CpjHPhe6by46DH3tqiS+IgkV9X1bE5Q7v603NrLbxSVhtB02JN9SuN
yO2YDJ9D6RRJzj0mIoCvk6FnJh0vqIvIngfOfDWE+myd7hYZ3O1eSDo9guPo6SN7
BFS/vV56DquewC3GpW1Ksv+ToCcVUeAVZHcePA1SeTTtbInUGm4vPJBub4BLtHfk
ugBXlMibMo4gRsNMQ7p0+HyIVDu3YusG0TxMESr7vX0vMYyPjRGQlIemZq7E8teU
W84KduzfPUVmla+SuP1xdhClGXh9DLsAWzeBMCOeGt2WeaC0ZYSIBuYAFnsbtmGH
8B3LsRR/QcpIQfB5jqumWK0ZEJnwckmnebG7rpkHojvdTob1679Z8yQHQuMsYPF6
XyYRtSPfwFRKXHwsFC0wa72yt9s7ffjdQlAnSMCsJXGKAkytQgnBk7RI6nHGELw3
WO5yqrp+5vpmBnKOgtxTflOYSc6OmkyoYXm505DrNaWv9NevTBswI4IhJcng3hPo
VnlCVZWcnplVd3oQLgRC1E7UExheH8bjn9JwqHH+Rp32MO2er5+YER/t05SgMKIf
8iQroM208BL2T5JlE+8E6zzjiPrfF07J2TQty3NHUV3Zc/8HkBN1yrN9ls2sH0la
vZBt9xuPAH953MRwSAczNW3VNAUCsAxZCKbaiRdKVjMAgh+N/AF9yaiHHqUi96c4
rH9W2bwasfWhByMrZuCBci4S+twpim6qZGWJWZiiJYY53baJiCzWjYJC/e/d0boh
/NJe8S/h/d6FcAAiWs8dhaYSu/Vi1qPIkqHdhe0qBLr14LmguCH1Fw/H0kFIi2tk
wr2rRsJTYkBsuy9Mv5FAFI5RYQ1R21F45D8v8h/eQWEOqg5N9egDfTfpVYfSERPj
tPDgxi6CSEAq5Cf0eLjbC4kNexsG/grso6BgGMHiJuLeq5u1Kh34MtY0FLPvmCUc
dS80EgVAZjnOoTeudZJoJtsm+//QQDmnqHErSUsMjn6kq3xu313E2AGD61/Zap4Q
JkmgBj/GdchJnECS2ObLXNNlvDE3ZepPzSGppbiyQrKUWu8iMeUxFFMYWZXMJJ4p
aHLsR2Js3JBoULsTIfM56u8RYKSTEQFAm9TxId4c0jklqojP5qIPGLTpTCNFuAHL
un4t7hg8n9EvC29KlYeIevoco04bGc4eNVw/EHUPeLDsONkHOPw+xA2BtuXDYEhG
SztqkD8vldFcXbEMzEmoKKKCM/4aNFAQORsd7/M/0F1nQHEyaUMv8OgAfR2u2DEa
RGR0u6lzDKeCyaP4iz8FgC5f9Eq1b/0oe5PjNbrD0mGCOk2FzFQFSz5fhQZqoZlc
LvPeE7r+0OYNDRc0lvXiO898H63hltaj8oTJ8Um1M1lP8PFhiuwE3oIzdzyHTLJL
X4VFJ9lYakVcb/9qsNI7iDjHMDgyR9soltfc70ikl+UhnX94geb3HJEprHWinxeZ
TME8fqk7oIf2MJjr+aL/WSLAxId1IH/1HL04yn6+cE2s1OUk2Lb8xE+NcoJJVMfO
U/oAuqkeiZHxulakZgNOuUuQgzcfmI3pCEY18GAT/6FT/Nhllmh/2tENP09ow7/J
mnu7gZ3MOhbOHv1prYT6qc5G4Zu2L7Jo9X6kmzXgVO1WUpPdLjCtsT2DoQPxFdI/
WRXXqJz4+NwZ++KIzEaapXpbq5mPBn8/0gdiCRaktAVd+E998DukhBMNloeKXphZ
lJAQMCHMJafVpxr4YO4j7Lwcizhj+LxiqAY04AocjM0Hcpvc9UaQVzEG/m43aYFI
PMCZfT9ntPp+Qo+G2Bz657k9WIxPuq9S/QSUu3XuTtUvFeenW6x62VKfQc/uXLC9
k8/nPFV7VM0yfu2QJBWe796oPHfqCXcm0o6ymSxxLOCAsCpXMlMx/AbXySecPuas
fEuzkjxhWzEBeeoW1sS4+xInqke39vhMQsakyqYIyFcbKYm17nOis8Macutq0v9u
/2s8m1KQNUlAljyEhw5x2GWrCXVRo/2Ft1ANC0UArflvcm88B1jHr3xmNv/pkqnl
WM0Hbc644Q1ytPAheej26dGJn+pobcitFqHo0ZGFY8EExSc+oQYHaVtGUMqiIGu9
fp7t6QV97Vd/9Xo5ER8owP50hmjrqJgWa7UyIbjA1BD6NuZMSw3wguiayMdtFKyR
sX+XbVSVA0Hw7iCGR4myFWcmlG24pCRtldaiMP7cL7E1omjhHsmiYW7pmZneYwj4
NVTLf9DFr5yxIDdq+HpUuCmXh3CZvg2rUq2NLr4PpQEPtvf9GMonC4s0FefFzRdz
eWS5tKjrSPAiJXLvvCxHPJhDlnE3NULyLEProFe+lQq8MlodA8vEvzX3GJzVS5L4
j+uLNyZYkttGOrWtfyGnpQ18x7DpE6lZultoKUGrirRepW80nPftzMbrRrQHTYPY
ArU4Hn3RQ6ICXEAnh1oJxpTc8oP5Rn8D6yU2ljBkON1bUuQTUxo7waBLWMdl5DKk
G5kGuCj4MWjaWCkYuWSapHsjz+RluBa3mEq2pfaUmnYPI6FPfzEfNYFB3gyasiMB
yyX+ztZQroZeIVS8seZhm6Yyeg1XC6Avc7OWf5EASzmQI7ijLc/GIwxIezuAEZnY
Ldu7u4a2kk/cTt5NA7x0Ybs92A/mUmecFV4XFIcvAbQXIsRbngRtRB15Vx1yfPHW
lwjVrBa5hJs7qNHIKUz6F7CkcqqDxhKkRSKsb0jOuI8UTj7lxww85quLuRPgx8QI
H3TLKDiG5+BUIXAJEqjZHvFz3HpN2Qkq5sr+rZrPAmPtdmsUFHcMxsQe25CUmfwa
zyo66HD6WQgLP8vlmT8uah/2wLEHsbESbsnH0IqHqXXoacK/kEPRN4s8EiPWqmXe
czKh8+8efrqehJiiOh7mo9oHlRL3ijY0zRyMp25crmFEcNJa2hnPR94ayLMb894G
F3xnf1YmoEn6eZqFYrj+HQjdtOz+NkfDmT22Jo+fZhwxURO4w+Ixb0tnmMaUS/bb
H9gLXKJLkGn7JDxqAU3v0X5vhSpvbshRKymZo/G/GvHZNaA5f1gL/ExuTlQf5GUJ
EAGQObwFU0KXH/sWooiFexxypRZOZCfXX9p7InsLuVvw1XKMY44kGRq9CZNbS5GB
BfHk/XVuAY5Hzwv9D+WxlPe6SCuX/MrPKKkPaefyIuDs7h4QH6ipkmR5jUD4NqHp
vMd5vji8pzYzcFlpBH7utzWdISnU9xQ325mKMLTcO9sa3MX32sCFuslxGWgFmdeP
Qfo7mFFu6fMtJH6335pmdvSF2+hFzX5iwUktj6pm/QGhqDFqxemcjGWFTzxcN70E
AhTpBjA3r7FbPk3ar74UWB1T9JKja4Sjtyqe6S/IbgvP3/7pwPLkZh87Ylwy4Xnm
MFFfRi2pgZ9AW/jP5Rz5eN8KFfasrrmRp9cqVI3WKRj5lAFoDg2icfbst+6eT5lo
G5ZgbZQENIGchClkf+34ExcRru54XPgOVn2hbiiMFFZtLiuLxvo4tIqQTC9RVFye
okiJ5EuAfI5U1IdNJ+DFVSqbdi/T0DFak+52y/iYqK8VEwkFWA9B4UBvz6/r/ILN
sWGjXG56ZUevzS22FPjwB4CnlX6Rw6f6vWNnJtFXTfAMC8YL0feb35lRcNitwJHs
FimFLnPsbT3Icklz3JTO74TSSDJjPLgL9H8BHx0SUTD9f39BJcOCIwpM4NqDo+Qi
H+FcdclJDIjlUa0Ir7zTDsvdoM0jx8vhdOpcByMkMBOt6sbXThCya2SSeIwWaJGM
rL6OMXD12lLFRoY8umWLPuyfEcAWSwd7EWS0ADKzmgzry70jLI/bLXWxXlXATjMd
JH9hHWPJ1PY9NCrrOytSdgCmfjQB/Sjo/YaftxpMc1LM8Brp/0K0iZ5qHxrXfW5a
55jRiu0VW8N3+Ukeo+Vo0prCS41x65I+fOMrz/gamcGMNu9EbX676wDi+lKcezLR
ih1pYKLpMkysIw1FhGL9DO2y11z2S0DtbLHi9rukEGtqOHA4G1/kFQtkM76rdIXl
6DIRwajqS3OpCa05NmSqjv1k6ibQW/cr9hg9F68EUEAcrgcNSsteGNQ7vI7IaSE7
3GdZ9P30k1AQ9t2Gbx/alk9d8KjQgmahEveaZjY7Hz1UX03HYVRUByPpygUIIb3I
9emS1TNivH4IoNFaSdMGdMK2iuc4adnDc7bIfaXRbBPL6Nx6+8y3vxTKIBLMPTle
5cyNZsajR17tTqGPB6Niwj2LEFxWKYpan5fm83DH5FGj9J6/sPvR/qEqmZXb65XN
R22EvCrbi8BZPZicro5Wt/qbuVfWnDSvWpGM+crUAiyM+GjF1NQoz29tJIoSrVU3
0iby1bnAI3DMEwHk4RjP+1ELRuzp9NwfGiSSgbcQW9vj+vmVQjxzryL12anEWSb+
jHevogcNBcqrYoTTJHJA43iGGh3G3OsrVWZdMWuF+Nl06iUtIWRiieeIqPGsVyYs
H4V6NlvSCcIi3uAufbjoBSdcqr/qz+o5skFs0Ckg/Ycbf4Hw0EYIA56zdejE5OM5
wTZKKHDCdUi0VS+16LoolL8xkMj7REWbAHU7gTp+w6m9MeNZUE3C9j0fSHJ82DUq
kmMFBd2eSlCrSGLvXqryemLZQlGlDxJXwpxDY7peoMs9Z2kdI4Oq6YHt/NfRgeNK
wwusYFJ6iKzgqNJSjHkfGMjWKFdadRj4dhOCUXme9hC3Y8a384HjrlRgexje562B
W3R+CgoKaqQ7QQdO0OwyK+Bn6N+z6SYnCuc8Vm+1UlKOiDsNOyZ6DEP01GSLIaYh
zhvsqHj3LCMYKxsWvuL40eK1mhJDLA7U6N9AGPJzrbGgjpW5kkzZq9Y6QoYWTN10
b+LPYBlpZ1SyJtUAhUDI5qc+L9bO6qYfM6uGVDKCRq956LktZfyy25KhkE+fYAPg
34GLUSNFcF/pqhvVmWXXrwIa6itWe7KyuNbjr0YG38ajP/vnyujafYPcDDtPdLeL
EVQ9u79SwK/YwnsndRjTgYLDYR3x0ETxogNkTD4QnedOE77UDFLo+6f5Qywo93fp
OzIs2F9lGpq86b0JHNSjBBDT6ZyiaHM1LUHqjAUV8BRrcLakTFdDFMPayRyPc8Dl
yy/10bTY+VSEVYLrDDbOocqRJ0sJMn5ZidWZDSSqcDLfUiBC/NTwPK5CKE0226qF
hafrkhp+ekJYWms5PcBZyyKWK1mEx3HeyV1sUEwv89Wc/rPDFH+83KWvLAMn/N4g
z7r8NN1AFjx8YTHJ9HFOS/ElhOjkyQy4fsYHuUh8OOEeLjIvkm/VnPVX1ye/Ugxi
z7Gl3L1Jz7B0EAqdTzrjKPcmwaw+QAHrVLoLxVaYruD/xgMkHS77ENL3zTJjGX+B
ndbQJ3nn3SMmFhn8p45ZoR6J1hSsEsfggCfJiwyruyKnTEb3/dMvx2t8KFbWlpsn
99k+j1yaaUm0BH9gtL/LwEsBbuPVgZVvMuCIJ44V5KAF+88JXIFUnr8POdiva2ik
nSMdcCZ3EPoxJd6zZrux+PXZJhQ57F5A2ynI4AbZA3cKmLTlH2BSI4G7S0q3jFST
v4WgjvGMxJ5xyuTACcyGMv5jYO9VHS5YRygK8Ru+mLveYnRneksf0TA9FWl8z92O
n/W6YWju0L+CyGhMhzMKUwVWNUWywkfFB1ZkUls39n8D1EfrjI1hu1adzA6eRvBa
jkubReL81jZgcph7AeUKQM+nL1JZnS++NhhxgOs49gcF3ajyi7+CxF0WoH5LfYK2
UIRIlJkgAt9gaO7eRnY8dBH+DqEtNPUr8Wy/QX/S5MNVjHsuNEG6kZ/p+7gzukbr
6ad4eF8pCJULbK25ShwbmUjbNYNFJW3t+YIp7JE9f8Qoxj/5FbvgpNMItG7U5Kow
x5H9bX03MxDmH8EWUUZqGBSQK6Qf04lnlgZY4o/hjvzBCnTmcBlexzzmdSN7/T08
9StWIQfjVEke9AiNPXWIMlHS2DQsqvP/2Ui3cFvjKwg3Ix5Hl8cPix2OQSAdjVW/
TjmTW0GU2XEtyVxmqXLo59lxkroUcg2NHHOCOA1zhtxdXzhRBXeyaT3SWliEmosO
E4hQ3wOIkDUjDAyl82wdMQMPA1jtb/Vm1TL1CjrWF3RSybnKxiqYWJYLApgQeAQD
JH24JaVTzZ94AtFQAk6JVNw3885B6f/vKOKeRJ2JhsApQxUvrh5/2zrZYJWOzSOQ
O9L6Y8D6y+qrKW9+NS/Dk+OIN5SB1vVEfMIIDzCDFjIK46UjbtEYf4ixNjtDjxQo
outVDhuLguzG9j4GckR9qLuanl+qFXOCUIhSpj7cUtPJW/O/i2t7pJTkR4AF6UZY
JJ3pnppFRML7VO1HI6Ktev2h5gUqsMqCK+uiSwip7hwIv7E97ZpLk5NaUfddZrNk
R1GRn3dci4E+7Z/h9Syzy5XaNQI9yUHmXWY2osr2dV67avI+T7adG/6jYFcdTWIC
dx2Jk7K2VtEGdvpWQEsCpwSuxup7hOIV5kP5E7//qfI1q0pygeJdu5Jci48Px+FX
g1dzREQ+d/G+GWLXlk4z0Frc11UaAKjMeZE+XFkIC+qLoY8ONR+CYnjzUS05Zz/I
yfegfG1NQNA0lEnZlcQhQIsvP3aM4byZUwr0/x6doRg1VX0XGmUHmoKxXFDk1cVH
Tc1M9U11hBkmq5F5C17A8ook1c22/vzo8nk5wmwsOAGv4+HhdvSEujUxUttxJv3b
exyCiSNBQd5uWMmouLjl6CUQEWXPcsQGyFBO3TMSkGM7SKF1qSCJF2Ju2O3KUhrM
/UGWXEwvNrgOCn6dANq+1WiNe/+Tjuazqfa6pIMyv3pbvdjRJdvzNOJzJ2E2dZC1
zhkplLOPL+fnS39b3oe6OJaEzaoJj1KEK7MK7OVCqzaoJ6LZN10RuBvOn2k8XSHx
gKz8DZ/Ome79LBslcacuU8QXRnUt2mXW045JFFsa3JVtEtoKxAHtyBM5lvuoJJDB
VLLs24QAMucA3xlthj6/H4aw0ALeJN1WDtgcZ0VmF5NguhdohVXGYCdBcJK22Qpg
8aseEUtl/CISePyAo7EanADzzNUDvAZg+JeXvLqg4oEMYJJ1NXpLoqOr6wvEcGi4
VzA9h8Ndpqse8vghXQTzc6cVx9zZKxeolyrLKASlu3n+4H/DmjSLcqPI0PA8Tn4l
UDZoZebHnVcLnhMv/+SqWgMCLYpkZX4QsrXO5wrIUy00D7PBQYTT19kHwr7UlOLW
5gMayfC+ooo9d3CpXyXjED7bxv1RKzJko52cA0NtSvmIMDiFCkIJc5oKqpzeQXVw
bAW/qTrEseyHgBr13h9Fv4N2WNki710panytgwZ3eg6Q6d+ZM/qoTlZA6O69ijnd
aTWMYPse7DkbG5Jd2Flmk2tLNNLOMyGEQpAB/KYpq8l9RaRl6sEqms7OfR0/R8VC
HfI+ZrV6GcWXU47FpICC/xbwHL+tQrUwGorAGVeWIE6jhzKQNjL9A6/kG0c6Md93
bw/IcNBnr4EWtPPjDs32+S0hQGJeirRxJeh6R0yxh3qstf7RKaiYtnfpKMLci7Qu
4ng0AMyc/Qw6kYQ/fIOeLf1Z6pdteSzeFkaQNJqsoVsWEDZyNms6bItpPvClMrHJ
1AeXtPqqUu4jbrrfum8xVRM2UeLUcumX61GV49Odej5rIudiFJ3xQUQV1ymhZqNm
6pbivSEkPDnDd8gQKzuvdQoidssbRRHQabWWutRW5TA/NEjN8Ibl1ExDvL+zl6gj
WCxblqSHG4bZxCXFzGsJFkIznF+icPbHDhYMkHzOcMDkFqH0cl5L+P/Fnuf0L5fl
CUjosJXTplE2y4oWSQFLMvd9yocfOP6qsC1SzqsmzGYdPUVqNXNWTyuocMw3CtHe
KlowbhCV/tsFeqQnA+QeyggNCRJ7ZfhY0cWYmHJVufWO1hq36FeaM8Q+5Rpbl9ds
yXsQngRwtr1fssbWchw4gfv/bYs+FY8WFITfpypvYv8dNR5vGWMF7VgB0dshGt14
0BFec58CeoQlMS2ex9DfwJPJisPIXSNQ9F7W1q0pdL2mIyHeEeshfOdguzeovogL
UI6w83tG0HUDXNy1vzASTga9NfR+vhCW1yjgblyUNoG0SO7MqmBTA5MLzhpSNZmc
yNhQpAgzkHbJApUZQ8Zbwle8inlMr43eoywACD5pDSDIXIkoZdGiMnnEKcSBppNn
TYQBCZ73QLRQ64AZkM3tNEpGewjL0hggoA33UTbItKkSq4Zm5QRijYmiJeNDhAIV
vG0rWG5hqEHX5NQr1cmIwnbO2AckB/nPslUV6M4r0BGW41ryM4SynAzRlWGmraQ8
gjznJ6oaMFispGbCFy1Ikv+5Xlw0k1cxk5GmpGqPJ50DZNQBsGOED+GXjOEBUPWO
BgE4cMdXUxnhFlaPbujcydoslBOH0fQQ4mdUiRlfuy2akWB1uiAdW/PUsv10v9Fy
K7TchAxeS5bU+1km2nuZl4dkSXbwXIvYPkb5LqaEzxh6osdWeup9BzndeM8aZ4Sw
ihpkdmbb7/QvXzr1icyA/tz+PaPusV3qCZN5EfATEZUqbVsCBiXKR+4DHPC0ja7H
3JaeHLJnZc0DLDBn+FDjupnnKFRi6Cx+E8cxUzpacgYK+iwBGYDUmRdQ+41E2ru7
oGnrDmE9YWfb6bCyaRvCY1ualCd8xNS/XIE7/znfOgdHZoEu61oh16zKOOPPVVen
7VJQnYpTiVBg/Do2OxkE1klGD7WS4ZVaSNttGo2Rqo6RVqFyrh5ifwAqg8lv0/Nj
hmO3Ue19AICHsAEhMRT5hFgZHVJulq5/VZroalXdSBJq//MlfpeJTDRehlrpGPy/
Yt20wXbeYOxXeTUwx8ZN3uZJ3IxmAlq2wPg0yRhJra+cQ29dyzscKdvtcsLx+VC8
ZRut+PZ1hDuAQpwegOt4ZqFD/N6wNTYRrWyPs7cZjtsydH+ERQ1q7iZU90tetFoh
9x0ew5sTSjstC9FBtB6wD8xgwJJHr9NW2oXlylNx4ys9yecl42fGVe4DuO+2Ehd/
FTNz5vihQ7n7vb+7rlrGzAt7i4lwjQEQSycrv4xFTjaobFg14BK2mBx3zyo+xZqy
KS1hu975/J2AdqyJLBb2VU4x+UX365/YxpigdZbuqS66BDwwztmuBJZOs9yhduY5
U86PVeD0BRRa732NPtBvpIOJ2upM+mQgi/z/KN8Tu3k8SntqTaUAkExWf/ZPJhnE
cfsOLdFJLj3m/ior4teN0cG/ih/WO5H2XCbejL12pA6mVCeNHcx3Iyj030iZjb1r
wn1E7sS+Tq9w7iJjxVKi2hrZGekaUO1+nuuYHLKXCwf2IYGs4hJqvglOxDDIyg1t
FK7vEGKHKp4vUAHO1kGcQUz57oZFoBF7zili5O+Fnft/qe+I6pJ6qmAWYTjD8sUG
VbsSxxEotGObY2ibzuRc8/VWFsKS+us+YaXPuDE028FtXjabQ7lDJQiNflKY6s0y
zpylbrx8ll8po7ho7KRXPCdqKSYDRMaBGCoHBydWo25c00IKKFmG0nT6aEOLjFGc
SJN+WJw7qFqmbM0e5xemDZm+l8iC5ImUvLHdS6mZVS8Sd8l43w96zPohZdGR59Un
G7wrYiPZsUhFPvbBwfyId+4ZQoRyC7CLpiWZa2akfM0eu2gEHlKRi31iCDeV8mH+
ciL/2RuUUQoSUs+myXY4CFTc/AXzedpslbc+MvmjZQCZIfmDZL6b2JN8Zw0MMf4X
W2C3aPnVRl8BFkgH1f70tYmXuZG1eUSTOd7TmZmbN5ggPA4A2F8QRORqjaAfsfkh
vVd4OAybuKnFNlAiGrOIAr0TXyROslXfFkvRs5MfhBtB0qhWaDQvaGJcKuGK9ase
i0+K9Sx8Bjfm48jRq1TVSXaOFCaIFmxHdy1FkEV/Vhy8x0pSf+nmOjtaMKkb/z6S
WnCHW5HGR/k2gDfL4KLP8a8nk8NK8lbEPQpz9odZpGdbbpj/DBpTvbUGUop6RFk8
yPiiEoIccNMu7nq1nPSrmI3CIQ7gt5M8/sK7cAHdkFArXpQTQuFUgyXtzcY3BzPe
KuNhIQ3GqFMR/OLbkGObGEfv7xC3Sb1TwCsiW6dRw2+26997iL7gjdHcOfMYj+Id
IQogRAAUXwH8ln4mmDUmYndRZZBqW0327ooSuvdl0aZGfSziyefqaqqJrtuz4eHs
757G1AhQ7N8uCPaRbSnXWAGiSNnzB2XJngyaxmLMmX4kQFD+/0NbJ3J5VKHlGOtV
cuiy+ReTfg2rrUllWtXKqpou9HrxMDFNCNsOU9+ZderpJj1uYRY8jpfHprHsljiC
X3yHqAsVbyfPCZQF5B2iuMbA8jxcphrOanZRMQ4ZbpSmAm/tF08hD8Q23BAF+qPn
NLj2G5d06RCSJr6HBZ07rd25oYxo31lzWl70aKTf0ZBTAs+aebT+QM7cxc/LR+Rh
TbAo477/BFTrNtsFzZ6wJAKFLcCODF8RQZn8NAWzwa2n2vlBYJ6rbwH9VFbWmDcJ
zcWR3/IWguclElOVtzg5LOTCOKP7u3C07/vvcUA/9Q8lr5QZsvsVr+npibwGOjJo
9EzGCr9BiMSO95Mwlel1Z0qzN6KZ8bvqDECz7qdPlDR3sKo9UFhJEXIrKtY/xuKq
y0BvEnb/aolH/66iTBukGR6O7Y7bL0HEo5rxdUPQNW4GLvQTA5u2JjA/HOneno7o
GJJiZiAoypfKcZDnaBEPLqHs1t7LAa0aQZdGWxk/bJ4419plIm1knQcMSage7NBu
ydV8ELP5+K0AlDMuMVW0n2SN2p4fXtcPiG0ZV3sh3KHi4PyBYChATzK1M2zPTCp+
C32BdV0B/Ml+j+BzTCUHjJ2D/2rd3gkFruyLEUnumCBvSCHRdtHQHsq9+WcXzLaA
qA330asNl5De16R9epWTI5+CVdkxK9CMNY99NG+wHtmGu8X/QUt/YF7+JsDgMWWn
rGrYRBFi/QAR/c2tdSVLcm7MWWUMI957ddCrWdMjL3zZZUKUm5Wl2I+WWpgHPqI6
BXvEDx0QV5CH88XU8/TdyU4y45PMBMC+6OKdYZ0uQnlpGs19hF8GI6yn1qVv/9dN
ggcuCrVBVsfq/wkyn8gvt3v0LWBN4oazMNO9C8xZ7nAXuYn4HCd2uRpg68kPepT1
a9yEfjXb24g5XU5rWD/smH3PDWg88eSFiHcxMn7htOItwVoyHQ+Tix7s8Q6Z9q5d
fy/DqIJKDfAxlJxTOKR+NSZt2sPZ4tR8p/gWU2yLbMitHPqTAW2tpHTif/JRO7Yc
ZiTFbLocVeOPVJAKWRXnHQfb8EDQ1hGzE7jxw2tpUXZCaSAQ93qNk+Yn8YkHSa+L
mGEpluJQ7/OF/RB3yzr5mFrPDulDLk0+aQVwyU1ls5KXZ5w3rcMvik+suHamkITg
2FerViTkRHucMdPZu3w7VMrSnyCiAdWzueLMkxFBmBxt5GiHuk/DgAQZ9CPACIUr
hAaCmKmfOjL+Jkf91jx5ptUQLuL9tRH1+b5tGyVMpdV5rZk6T7LFybtTnE1YP6fX
waHAyCJ1McHB642PX9ALJg60rSQOoRmWE5ePU6TEEWVU4R1rdH+US0lNiVDyZxsV
AbDfR4e0tB1ujvhqghQKcqcQKK3MAjn95706NeUrDsYlq5fuwr1vhuHF8xFSMpk0
Az5PRh+DCqS7j8/322zaub7ZzuK8R9l6l7XDdaosXqKN0EhWwNGStbCE/5RAOo+l
og+5/mb4uEaQ8evzelrIgHnv60L8bN3lajcfeKKabEiV9xlPFlyDpF5fOmkjFhLF
0Qv9bHYhiEBjex/nDU3CUAIAHdxu4JrI4Rx0BnXH7xbQXOp0hFtNn4jvE4WKUGVK
7UewM8RicnRRxbZGCaGZtTMM2/H9hHE2sL37FDjXonrpHuymikbAZztscCxVEmDA
rGB+ZRIAJJzeND68TFTXRQfI9hi+0sOFPcznJRkGYLQnrHoaWQqVFnjt55znRn+U
xbTlMkK0xEGCvjGXYe1xraMWR5xwMcormIPO8YzLg8cBupawS6kGQH1dusXjYG/a
BMyMyvm+vp9hgkXNWCBGcc25G9UW0rbqniKhE5260K626TsQwQHrQJkLhmeEEtXn
EQzX8d8zo+ysMw6auuerNQ8fCdUAn1JIOJJqFJ3JnU1TQu+cQvedFvUVVpCFjAKU
ox4rT9CgA6RIiBY5B6RmSZ/KcBC43Ma0VMHFflZsvUPo5PnNVjqp+Qme8d/pt8RW
BWGHQiAHh676d7Nlgc2XsO2KJBWa4kzCOQJ4/WSRKjLCppSLTh6GoH/beiSR2SPU
4uTCpj+TReoC88xXsZgFw3FUkB6bBn/LxSFOcRirh8hTTnrYsIRh/GrW0CMk3SHe
dxCoTH0cTnIE73A1PYx8jCC8rYpoDk1gA6h/vmwXc48LnLDmEBngFFdDhpoGegFp
bUojoUARk7AV3PsUdkdbjwnpnNLT4jPNB8+qZ0Nh+XNilDOz9tRJXeXNHHPcTXiH
NSqulyrvoekA0WpMxMZXRonrsilUDfRDFGaIuk9xdG7nwbH1QAVkK1DH9jb7bNeR
2bfWNDKptI4r66uVbZY/lYt8eCCUCO/tiSW5eHELUELGAddoa75SlTjwOxr4u+Ko
/0BtPhg1JZJUgowk1Q9p+Qagif1Z3ATB+cOff+QXovX8Iu6S4CY07UxC6KhH1682
1YQsZ/tlqr7hwSIhIAXOwZWrP0TdmPK+q1wY9CnIE6qNhEwmTnDr1pGh0S26j1Ps
ukA8QhVtOk9QvK/3MgST4snulknNzE7iVy7mzdZifZqUBgto4JaK5z5xtBlwDUab
Hqf97P2SnplS5Y1pmho45J+K7HJuVQiTzIaBoiBjHxcCJjmz9U62n8e/I9b70g55
DMHa9+a2/ZFlreDA4Lvs2ZDHHDfW9GSWeXigkCQYDr/kyvuMkL0NtJUqrUKVf+cr
4lG22X/QQ1hBpMN6K5JwakSXGgaqpcRwFfJv9z92BJfsCmBwZo5JA3aWfsD1/XKZ
sQ5xq4VlaVYPlfQm01ELfKv618Y6nP5WS1neYRJQ5W5KSFuJOD+WFseZUYveHfdj
UFb1x53Ro/A6bNSMYOgLw/TjQo4na8xbU/KbYXkiqGkLo52tKKT5GZsLMi3PdHds
sCUfSRW6mosSw60/sWDm3WNI4VS2rUIocaLjj34MJHvWcFOahEViGWcj2iQFEr8t
w7CFxzVpUvgWc6ZrCMCiPqwDdRLbS5vUlWqRgysDjiEltsmPTEQIH2PgmIRKCulN
LPXdcC2XRk46xTZXz5uiWLedGvd3hrsjyTbQbEfvYoQuoF7GDp2RTi11sVkzX+qy
PMThCD+H1J9JVc2QBF0eIsG+Bg5IqH9FOCfJKhmHj6gidyZUNxD3twC1B1zLj9O9
3gB8ZrJO7y5zTw70e49bBOWip/aXE4x3IrnOxZj/siDjVd7iAUpWy0n/OjXAv9hU
Dt7bCrE9O1bA8raTTYQkvfaBSa3gOH/PUztyfghCStVTc24nQCVU0OQKzwOIFrqz
dArznjNr9zMNj6Je/EcYfphBateWi8pPkcn+kbTmvTn0EfCBYdV7pBfYiHISLX3V
fc3r7zj2mp8orJ1lzWa7UtXaw7Mc+Oj1IjCTOyXfVWrGTg+hv+2okfrvAgFF6WNx
tF+YTKkcZcyIy0ijctdAov0GcFm5UBLJXRC2lsJdQeQiUVUxdIOs+5vG6GYMS50K
XBHPNNomJXgZnaX31xbxFwMyoNshGVJgNvJbwkOKQT6rPUsxXLZwmRuw5qo/DqHW
vqhLibvyn5LdNCpf1y5KXYdUGQZa/NM2xyqPO0OiJAbhSofG1DE8jENCTGl9GEC8
zuShX7QZcnrMqZFiEEI9GgsbQV702rsddm2aA4S/2qqEmSG7NS7FY4oxf15sZfir
U3+pSI+L5D6zOokMoMtIKTGXUEud9x9S8n9vLVRWQuQtblCXtwCUN1/LFm9wwfZJ
mjaJzugvq6jlFqZDRjdmeBNp7Nxky77mq1JllO83C75IZFgMBdd+OY93HiRogMBt
E0bgnWEoUPnP5fCITs5oTYI1U9Y/7csJZkjfha2S9gMQXkUtKTus9fHFUndPhS7O
P2AcgA0jMS419ZIVx+VTtC2qRsyfgVMdEQ/PEaj7Ll3ZYDRRDRj4o1vyHKFcR0l0
w5tJmwBW1Sh1Y7YOgxahe6yUErUbAP5/B7208rO12F0ENoXcMEg3rpI9OxZOYn9l
jSQ+aII1nKGdse06LA7WPG1xOZ1WrryVu8OD8yg3vLqjxZhoYdYvjD47PdVBvjF2
O14SnAAJBUdlKEl/4ywP4ZhTHSdEsi+dMv3SBfYJC7jyFU6ASdlE5epaFj9Qf/zd
H/kVnf1Jwq51S+IYUjTFi+boOtkX2SYPE131j1Oyvkq6T6qgjP5+XPue7vds14C4
/c9yM5kj5fV/NRXRk06220HvhNVcdxyhlwIobvV/+ss5Gi0ZQL1NxxLMheWN1911
mbejO7wmX66wlI4roz+cFn+UyXJ6nf1lrsb7qOFxgE9DI8gb7nAKaoRn3lNpZMrB
mFI5pPcYud9jC5+QzhIVHOMpg2C2f7gRHBt/jMIlV/d6MKUfxJRQwiK+RE4UJuDb
rqFVDdgCDn5IhCb9tkHDEpebfwQd0Nlu7V+ljJq3BVTpflkAgJL3ubslDMH1THKi
KLtuNj8CUS7llRsyjaBlRnXCquzrKahRtiB0R33VpdUiKeaxjyQJBPFkKf3MDjrl
STuXlcd5FCh4FjYoQK8++wRjr2YLVGO9I/zTQ3BU+4V3UmK6savJaR9L977e91S5
HI9GnTCdMQs68AsrH+glbtzSwmJyNhNEsckbJPPnARwXZQNkwQIde7XYRhc60vUz
cQz5l4Haq0LKVIsFxrO8U7OpllhPgMxcPGagOQZTpAmvowlyxrhoDlqHtqx7LSbz
NGyaJ7nu4mcC1WW00uGL7ORx44gwil2aW4Yh0GlIyfvipJ3xWqNsd6Xm7g8O1Dk2
gbNzFYhcb4AeGp7hCy54nxZjw4/TWgEg3QRp/Qv0FQgNHdqLru4J3B04JN7q/lY5
2R3+kMEYl12maVv0MrmT+4GjFO9WsPHTL4+Z4GWbYOJssb8abz4WLb6okjikmnxL
29jj3cQpU5x6xG8uYnUQ/YgRXpmdobcdZ5ZZ4Jpd57Qi2X4WzRT4DTIUNhcYgs3Z
+66zYka3aP+P/bGvVrnzDStb6+h8E+R2ynsV3cLXsKfjDvLTJ0t6Q4zjO1CtTMVI
dFjDs5OikV/jo6W639UDnkPM/d/pr4bV1DGKkcdLESwyXC5iLgcZfSP/wK7kbZKr
ybo7D+xEiFG1blW4uIXYKhjDnmTMnJc2iHV/CefbUVP4tcMPezkhaAGmbih29ttP
VXuHkF/Pbt23646f2788MOJl0gZfvm2Fz/XABHDBidsfnyqyYnybXWnsXJ23rKkg
+HswRERtzphHnNodm6RallE2OIIfhN2R2TEzlLeZomIWYQ8L/LAdtg3w766++27R
vYTutt1v1VlhPSPx5h7BlLZxp5aTunE+j9rjqxlL1VenYLf/msISym+OFQiM8Yo0
sjPDv6OWsIeRSLU9D4WWQnQxlOSNRTvFFckj5JUKt/1PaKIlTqbzh0zzQj5lV93n
WSN8csVRrcnytyI0M7SpZyClMBidgVnyDCX8OzUSpIf5f8EwGjDjj0QpOFuGILft
MtWtg2Sw1LRcsHefcxknCSTsz0snqD+3HqCrA31cVQpA7alHuC7uTheokEdgcM2M
mmXI7GrBJacQtHtV8+gWVU5i4VfwNuoK7tyMGAtAJtZedajC4bvkSyjm9CCg3tmQ
ajWGx1sfl2QRYcCI44TQAWq2SKLi93fzde9vV1W2Hn4CUc8Jc5yAFbLT8bzFFHUx
FK2Uprlqs/2J9WEec7N0ID7SqBP7qURN7l+gBDVHF9OLOfy/GOGH2xx/jTkKEF9v
QcZt94oAlXwyXZ0gOHO1HXjw3I4zya+dUtOP6C35dqkDgR5/QTjLk/CsbjPSIIuh
F3T4MJ1Ag/aqxJEbYuZp7WqcqskV5Jh4xctC0EsGc5N/eWvryupXVpeZWMhZJ8me
4uHBpZfkf2LRdZWdWCDFsmSWIVwit8g7zzMs9gR9bUnK9frCDNMC0210WGbcUUIZ
nazwFRLizLoOotk6WCbK79jGdYSl2IWF0jfyN9sUdikz8HIZi11w8KjAksGrK57b
K0TQ59sVw/HGXRvRxnuXsYmL20MpiHES1JDj5TzGTbj3CzWDsCXvMb1Da0BgD+Qw
KSvxT8AlY2Sxzbx0RWc4KF3Bwq/ul52c+LbM+TQq1NM+t0juf0/kwp6fxQHVULZV
cKHrr/CvoZGrW7mOcQsrtoQeEXuCKupZDMM/1G4YPIkEkPjh60duOLUr3NDgYFr7
r/wYbBEENbI5wETv0MSzd6dtSraJlz3R8R7kciiEYBkGTz/qpZzMxBl5mYxSR1k1
vM/5HEVs/ZxLEchK9HcbNFKvJxeAk8JNzV8JbQyASzFVaHauLwa7gtA8ccHDnViT
KIkgDr0Vg81H2AkzeaF+/pU/hsQMANHMKWdsUG9doDHRb4vmPTINqmzN+l5vloJA
a1Rk5iAUdUKPf/sy1Dn4vifIInxICXZzD/qd6gZiPOvm5e6b+1bR1wljcNj6LyxH
EjCqLysPNM9GNmYyvB+hpaSH80KE2haiUxPebYpaBGRdvontFBPYOGFNjlIxLh/D
5yc53f0LxjJPmpieVUf86IKIlC9UJMYp03+RBc7qDMw055gywb05l7sYMONR90d5
zOYSXvSSIWssXyYEnf01p0g5x0zD/QlMdO/x/WbEF2ycVG63zzl9TzAqx3s8ZzWs
XIQoXd7C2HHHx6R8Bhoqs92rarcw/XjXsCBhL+lcTiz7iJYEgzHV1Zj0JrAbbuJy
EvulkD5WAa6AYWd7AwX3EmWyGbibW1M9oU6YAn3VFJ6+rJ/at6zINe2qKZ+Pei8c
5767E0eJAmJOUR2X53Vwf9vh8xiC6BHOLB7krDIzY1ZRURUz5nP+agsX0HsxVSsB
bQnOfp7uJJ5v8oiODs9NHYxtxsVpTL93uOo+rtdAr8Ofuy5XMAlKitp1DUdrgGqQ
eeybzRDDToYVvVTl1NnMK35h7tgx35FB7IcxWnAA7EbRaAFyP7eZFAC/MqfTnLfp
baouaS4s4c25B3OzeVBu0lCTmiV+Ur2CBfSGH0TL/1i4bcAzrPQSVTpa9PSbE8hi
r/n3/PxlO2Zqc7wbab9s+avdvp52XPs2vrxD0VFsmJ4H+trLp9TeLWQul24Ux1bC
SqhKiNBCCxA/bOGv2TdwUK6dwjpSVQVtdhhKg+LUqWbOVhpTkLr7pScfGZmo+Zzg
9p+v1x7q41iXNE9i8XbjxzcijFTA8XdSexkvscQ7ozkIojYi+wmmCoG1Z3pJO601
NwUdudbUyNuNlHRrda/FpeBHmxer41ZBnwBR2eRNRiLmgJpfVFWXrXj0egIrwafh
9NZN4jkpUn7OOmaoruMrI2gjvSVvCLvAWzzFhGgIb3apfGeVEys35YvhNxYGCUf7
8MaGhSxrt1OVlNKZUHiBK3X/V5NM1TTVZ5B5yi5sitsSsRbXI3+V4oU7rnEGERd1
q7ebdbB4tHo/fKRR7xER1a2e5JS7H34+S+9c3Ahc34HUGrTCZrsk/nIKHUnRbDDR
/mdMNQ/M/JTvlqK72ufC6cCIdyZyC6om1dFYdjS07KNyWUtrr5DXjZqHGwxhk1U3
/WKvQhliO7AUgFlR4dU8W/P0MrEfhaFWdZ7q7BgzJehYZ046ENPkOEg1+yMBnpBH
524Wup44eHPqSaeXPdhc1aKCQt7/tc3F30Svmjcn4F1ylFWg9D6reFd74Fb5UffM
pEFZUotXXv3SJBDkR9lg8baPZzGEx423VP3X53XnRbmadA1fVv9aRsmPSIbPuwRb
SnGR+ezml1dHT9z6frk1VGcpSQJJHz2CFmsg8sDsiWg6btjdizZXr3bP6a1c5IdQ
jxl2KdJog7vEEa51yeOQoA9NIJUiDB+X1R4vNslVzOkIc7zbc477L4Vro6K1XzYA
651B4FfyW2EbuEqin5q2d/eCDlhq/Au23ZzxRYErrJAgZq4KymIFpiKI5b5msT5C
kSMPjUFeAwmIokTsT4N9PwK1xoryiUZuEVsnBK5K/mTtE7yyK3lEFzxNO52lNxu1
zMGRJA7W+EnwYzJQn+clbHimfgY0pxL2SqFtNHLAZUv1plmDcJojepAbcDwyHKex
XRO7YBg9GHy7piwTvEpL5OUYg9laqEgXErfTtwDYZ2GI3e1Y0jrSPqlBlRYuII2f
UXcBJ6y8O9GRmaOMCdWsus9vbZE+PGC0dFKdAneKlvNY04kiYrxOjs8jFVNOMgEW
7H3Rljev5v/Ku6GmHEbEfvaVMEWcdBfB1ovQVUF3KiVmNLTmDChoGnFKQoLyCK77
dWwADg4uvE+9fkR3Tcu68xi05I82kOD+FYOsb0cP8TCrq0nS8eJLCQ0Xt3L4XV+x
iQkN9dV5REetoWnQ/QTZQhjt87Pt3ayI4P1UaBR8BPFYa0eIxXdIcvFapuNibN1o
8lCqnLN7cZZcjNiLJwHhrefwuL4r2Zx6y3tExLLIgN8lBRUcthTbrmVfte3j3kz4
nl8S08xH8FfVeMy2vVUCmZRa62PZp0tVU5vYL4f72FSD1jgUmNyLaGsO28hHiHyF
bJLPvBNiWaJ2wof0P02/SxOehRqUMbFc79kBILv8YCZG7t/4cxpUE0v9nEGDa7AW
ugpq3GLYvdMJCwPy0QJElfGOEBXAqmAh6CUXCEBGLDkRqqSQSDyRmBJIOLThpc0h
zbzAXvUZ9wjIDXUXuXqZ6x/gYzp/MwQG1UD8LakYdjaVYVa3OdeLf6znk6glQ4DX
MS+kmkryIrLAqse43Mq9QMJ6F62hppTGvuc/5m9Lw5DanD+dKrjphDFnAztSwgMX
aBdGZDPyCXxavwLF3Q1mMj+wWutaU9IwC0jvQg8jzszulVxzCzoaysuv5ZcHk2Nt
EL+6r2/zzK7LlHfWGXscoRk+fpjHhFp0SSHAVCriq7sjmgSL9THYIKYDORN8K8BS
8GNbGJ6rUJXgV7SIQZoFISzeCAaGPDuJcmPqCLiQtc+MdICMO7fHtpTJegG4r5M8
EO6H1Ixt5WR1O/ccIBbaOyTeP+916F+wyc7fWHaSStfjGxRmp+0AxLuWPBGBax4g
722yqsPCbXuuVHgsyUe6elGZ+mj6D0MqKvpi7KNthC3IidFMyyGcGw0PP6nQsqyL
RDDf5b5paWFMgSBgZxWm0Ri30LFmfcebhNFJU7vINEUBt8WfmLoRfB6WPunkBXGx
Oq/RJjMSYn61WlMUvoiDWT6+eBe38d0cs5Jc411vBZh7OZ6Ih2UJfLV5J3PklhNS
hBJgCIWb7QOY5298fL+q4Zs3xrNwj9nmWRBAaBp9Vkj5GY5m9mqT22+ZrVZqFMXN
ETAxPvjE6TYmeNrfKBIVxvWVmQqcGqqeXnVE1d+ANrHQQxKwJ11wIK4Y8OTLGZNo
Ik0qbUOJUTd2FbbRQlVmkLCv2Twlgkxw9JVMabP/DftE9KTNweeNXsMF+wb80VPL
29kRDb5NCNF4pzZoj9hRMu8rMJV4APvKslqCK43xUoSR19NOoiCHlUrEmOGZaAHU
3Iocbu5smeKR+vPKOgGBZdjlIAX2SFiWf/4yz9GM/bAHP+DxqjL2mBf/dyn3BjHt
IHZMdfSWcuwPDfNq7CTSfkUBBOtmVD6RNEVxBOO2vvbyknwv+KaokwCxPDHXfm1u
CsI75u0vS5dDn64bO618re+1vyWKcWInkB/rpmzF+CpdIacZJIPsG3n6xe//6WR5
iGWuQ6/0O6fEUn2OawZ2QiRR/GJ0fMY+Ipb8hJ+UssLRT5aZiv/i837JXIRHrOzK
QPJQkN6qbz5ZKHDwQhiCq/MuDb3CAyOr/z7QeGOTSG5gVD8AQjYeJthacGFFAFeW
wwLfTaqs6/xAV0svmHCEf8dXMQFw01jCw7oI4w+/BVYey7rS4CLM7vyCQCB4juhZ
DV89AJPTIckPAzyJiuNDdvJUdYn3btK5UkrLWWuxfnCCYMNbMAPfbLULrzzB0Znf
jwUMt2mAcKgGRcQKCT8pDsYEICASpv4Dn0ZvSjKekUaQ0VXi+lOvhdtDCjwZO5OV
KV4Yd5wWYzd/NIc91xfVYBWRV8LU+3lC4WKOQM+lMHEdDC/rlbQv21qbD4Gz3fKQ
xdcr3vfGPtvZMY4Nr4C+FrAdipJwzzo3oaA6/aI+Hw5FxYtbcmoKcML693PmHxha
nsB25B6HxdUBDBr3vIWF+M0pu5lBu628B2bb1syT1aJbFLEmObMGSUbKIG8FOa6m
o1KYagnuglA9kS2ctxCJidp4kMxJ0nLbL5sRYYGO/QyWe0BBWRccKB3rs8cRURZK
3re/LDN3EVrrkk+QLbBBRAfbpfutgr4F0RqR0QFH7osxaicbiHDMSUmCjFsnhGwq
a3Y1r//ohInOhw7trSstiYKPnvDhE2hdl6IoCc1qGypNJvnZZ5XpN+vVqX6xiGf1
AGe6r05loOeB0/U7ZFhVTFIf7t/tCeovbFxeoqMXDDQad1SXwLSdfGgZwf5+nP3Z
w5X4Uheufzzru56zAEw43LdoR0jCkOJofiyAPl3hiHDbtUkUWaSp1UxewARHaN2n
kli356yFPR24DaBfx+qnU1YTai0FohkrCvpX8xAqI69d1abGeq6/CJXGV/0JskgG
417jlyjMXpaeRJX2mfaG+yulYNKu+ak5i6PwoFyDv62w2BiqwVV4SRJEPlMRXprX
PSmjdUeRJ2+VsIGUiZW9EUdp3zHChv29wcsNy+BUbQBEufOib1dSlBBxDSvEEhAB
rqzEuD01wCh6HPuHumvD5QbnbQgFF6Pxl17oyiYM3hSDw7oi6z6hyOLNC+hZQDAw
8xaFjiaq4G3AMktAxDqWXdMMAakQxutVW8grxEDiJi7tlx6Jx01bWOZAgH4cgpzZ
0ZohJ12lzcZ2AxdtmHMKRyqE6vO8RSFO4qBe7P50ydilSxCQN1haJnEkkfnyWqWC
mS5HWm3O0he0M390j0FYvOxwidnoeVvhbA+xnURI6VWSN/5ZHCxlxadZEGQqt8vF
UM841zz5Xu9OHF9C30WIoN3g78aW+xMpSmh+KLMYlt8G9ZNPsGclMGmn2VT7LAY0
7TrKTEJHkzDN8i/dKl3c1DHL2VmPbAwFMWX7uDy5dqEGal2E8VbLGWXer1YdTKjN
55lEBwdEiahwWFH792zmkOZW5V5fWWky666HXQ38TpgulWkpY7P6y+ntIFmk5eSM
6uvafpmj7EglGu6/KLGNRNltuwDDKntsIlwjpFgyMn8uS1eusHgNXsUwP+9voA/z
DRI/Pfks+cE8TwMnk5VT/Q7gQEB3I/q10EEp3xmnsS1SRmcbKLQqTbzUGeaGUQNU
Bh85QLaWj0IMut+lomtQKm5VtZ0Cqt08bcxEXNin0YrqMG8R0vtaCQpPQ57ID/e4
HInRt+NKSwRBufQGnSnoFyvKBxAAZ9UF8c7Grs6iSU8/F/wfBurly9FWVT87cGIR
IZzag5jTHnZJWGLscFYo8AAcLoCAp9+4SdrMShH9u0fCiV77a9FBTNn7lFQrlgVE
J1DFluXLTOSL0Iqrn23YZcBUEnt/G2rtOIyqSd53k0F7TnCWPQxCBmD2AD07n7sw
3TocE5AluafrsduUPnLnKbmnjplZwDbRrLbtE8ybJolOeAENF7kEijkmRvl2aYOI
eEpN1Q217kYHdRIfjt79LrOcQxHvRT9r7wTKaxOt8SgOYuoZHTEA5ONLcSBg25mj
IZO4V5YLqpTGvuXCA851WCFeDGy9gs5q8GO9ENMB33Mmd9YlGlrWsjRlmoYpJjK2
xSJEtgChpqUsen5AcjWP6N6kCZM3uwT0TwjfM9IrP7vdBRfvrDeo3eTjytk3VaTr
5jlbI+TWe/EV3S6M2F4WdM+Os4i7w0T9VnCOHa4xTvzmRx4yWidOCo7x3qQH2H+G
jcB+l3HEK3bxS0D0riY42b7Ip+OrwkdWrjjFBLfZ6NtslJkGBDB0tmB/r0RFoA8n
wtgtcPPUm1uQL9fyEM2DjMftx9WGyg4gvLwfx4FP4cmJ8yOEgow5QGK5h4rem7IL
8fduhZz7lOkPACYEAL7VfQP1EEWqVgS3puimww6khhiKX99bj1+cnkrafMEtwSDz
EGZ1i/7mVnL5HsyQ7hTztU8R2ZjV66qnQWgTIJ3abEIbzNSEoIPPI+2mlLb3k7yo
M+Lk3Mo4Pgq8SYavePVs1LWiGkgfulvSJpE34DYbEO17JFxWgWVPEN+Yx07/eh54
IxBldfqWGGEGVqVrcafe6f19OTdWPIysizOv8CzN2zLjoSI2iQVzHLW0bLzjHBe7
ws68VyRz9RjwHBeFr6e6819DJPKgnhga11GlBnU7ZyMOxT/wWaM3pXKfS7vYGgL0
hFWcjJzlRkxe8s5ZzlD2zXzfJXmn6y5bKtFkQirVF3Bm6n1miHVVDz+kp55hxPSo
t2H3vl4CaDhOUvSnQERob0w/SSe4Y/fYEIZT43UIzV83bzmas4GvNpfM/5NrrbOR
frp1pE4HBoNfH74DNCSft9feiUJUCS+3uqZ6stecC1sWi30PE7nRhoKnxHYyiJn/
Jz263CY+/6hqPOo+C0vFL9qk0tu0YaJWZKt69R5EXQYyOONPwoT34hwJpvSYi+h8
10WgO3YiGD0BsvG/5h7OjTEwC/abKOZeg1bVI/qMj0XMb6uvsYti8bR5+veSADhU
MJupirhBUYur3bI8Nv4WCbFB3Evdr1WsQGS8cEjmtIdnOU/t9uHzu74i7EOUfe9F
dLYvGrmw53YPOFQZcUZfLBsn3NYiiF9zp6Qr971sln47h5aFXsDcbVqyGd2ZilNM
MmhE/YuMrB22Sh59o1ECH6QW4yfp1j0w5fmZxyjrGQ9/8MMLZhUNk/tlIA2aOrj0
+8ESFBNaSlWu6Uvb+XMLP/8x/GVnu5ZRazyAyOyo9pJCEa5qrokDOHr7QHx8f+mv
ZtcLJyaRyZUF2MISqFSKQI/yZ0NrTtk3sTSN6/BVHxp0v9UvrpNLT5fW2wFsCeFj
dGg1PjGGoYVnMo6xWSHAD4xuPsOsfV/W3YBWDEKXdAyYPxoQmc5Y3OzOWPmH2/hu
bsx6eK/MDHIFaBV7I3S4XIxbUU5YxNlkw5h9p5VErHSKwKihCxURkdLsL330OLYB
94aYUItc/PXn69Z0IMjiSgh4RZGwM777xpuxITjKCDG7J00Gmsy7zlTqO6TRCQYP
JeBvb2ND6xgXL6SIqPTxSj7orJRwCak1oYGSLyR8SZeo00dv5eyqGgUONW3oKPzP
EmclLakzzwPzfwb4SufYYRKAgLEzi+LDS5CaU4qMAw7JBxDSRwYQ0jA5+4dQHpkb
jzPUWxkVefoTB/B86Drj8PLnVLV+B2FpEE4e6a3ZAe7pO0cg1jwlPr2OANh9+iat
SMDNomTYYGCWx+9nAzwn1gntzwIU4LwpnpTDeqvVxK3OiZPRfNBUMM2TqrluZGCQ
1inYDufIftXxYvg3vywkxtkmu0cJyWBPg9xPc1MeJWX5XH2mN+YEm3P0c5A3+Sl9
KINApqGIYWBC0FCnAMTY2d2e0IVdjcfHTFQYYfNplmitgor8KENj2sRBvgzDOxxZ
phJ06wSku1sr7KaFAdTyXSFXA9I4GDQ98/sQJk58tGCMWiLMEo9ZldUQApo9MUfi
FSLeXvtSabCSE8bmKvDVegqOg6KwYdgA1MiQQvxn9P5KttVBqHcernoamsk/3fBG
ZktFWzAvCjAFhL24xRGHTLTzFifa9Dia3hoPjsey/w1kYMifjwv2kwpE5tUKWU+r
t7bFkri+AURlgI6hnmxwvnI4lTPDU9VE1T/8uJ95x/Z5+BW+NTxm4y+gkfyWFedT
ae1DMiRvbH6ZPp7+bW1CvgzMUlqlUYup9Etxq6QqDFh4XnaYwC5U9Lx3dIZoF88n
HVWXFGhPkCFR6PRbFjbqy4l2jBKfyu/cSPO5udhl174Pb9OQtvLB8v1Y8AMc6AjD
EDwLF3HqEI4bqOWWcPvvOg+hJpE3fbKlIv9MATzvRg1TewaY7mZhhp7TP9k90MLI
BQxB8uRxd37FqXSxKeb54hqGIIj99QpvW7VlMzMrWYJrbip+R2fO80UXlwVU0TPK
lmTs7R4dNCHft1GVrm0s6gNLhDE2phq0tVaZKrcchekw77IMDQuP8bc7qNB1juLj
LByNM5wBglZR/RaeXmuDzV+GfQo8lCqi7zCUYEW5bwKGUIqbL9ZlsmXtbX6Npsyb
WZPXMsB4l0vs98rmID1XVaz78JOg8ZHI9jSFN200fI/9UMdVDpe4HnN/UQSumRsa
X9bq/YZjfc4EJTwg9zb75RGvN0ODruj+vD0atPk2pzUzsLnECZmYRY7+kURtS+fJ
hmoRlhLacWP13lCmlNGTK7a7pqN4PerdcS9FltCV0/jmfCaVsc/M2QjWMtJV6qke
Iul3N4wSMG5M+IxJ6e++awrzSqELQw+RYTLR0SgQUimxU7Bz8IRKlkq30UxEVIPa
7on4omRvqvXWOIkzQqfc5/l8xTetzubF+hupUvnYUwGgyoQAyi5j72fl4SCP4+VR
k5WvEZ+BlGpK07qy2zMETZZd9KaIkXSCHCLh50oF5+mdlhlGO+4iyZalZLGfFWsO
j8vdTi5MhOCVFh7srfCpgvVx+6p6RNMkcmV4tCUZVB9QCcREj+TFXewvnNTIzORz
otlpqTzrHuuHpaizJmWjnvkjm8TPTUfVpSkSlpVNBnDHLZBqKzmfYF7ej5kZepX4
806lBmvI+FZHmchRHrampYOsqbXY1PEArfPsvIHb9Zaxncp/NOqE3D84k5Y7d0Fs
JgjYzqX71yKtf9hyHjksKdtCctMNx9bshLrKZrNcYixe38CbKgHY7wKuh49clj3Y
+wDtIStJSeryu/fzrH6Kgw3ZSbqOJrUk0wOEOD0/JSi5RVEjXqrhHta7EPgl2jOU
L7asv2UrWeEBTsm5r0rwXShPLeHb5EupQ0iiuuSsAQ0VRjHdCpU6jmUVa7Nxhu+M
f6j0w99MHhLma1Hj4XwcOODYAwlLSiy8s2L96QdQh5SCOH0K8otXNu4YvFec8sc8
ohJuMkA+bMoxjzIVHdzcU2nL5iMTxUguRmPwmFsGaBlhC0UcWts+u/6jRGYN9+Tt
tdeXKWCVwO8yr4QMx9eYaS/MqYRciqK5n7xddomBnOQ1gPgWoW4rsFBnFEFwr/Nh
QoQetDvwQb0OeKi3BXXDfzL0KwMvf9hVBkAWs+9iOmm7Ef8k54R8tNvrKxXg68vh
4OISXQyJoFyZBJufhrsy086eJe11dBYwZLjq170+uTBm2zPKEKP6cHFed1769pA0
KoAWTuH6nbeuAIMNG4etV0UzYiiFwqUchSZ+uCKGIzBpg7SnGBSD74AeOiQ8nEqr
qsTqHhjvmdYbyZnSTZPrMq9URwC7BKQ09FYT2Lq18nW7WcGuzzAJuYa48v05wd7F
xoEcICENNolxq6UIaj2IrI1JhTYCIDdjdcb5WPbuoMqi1sn5FWpUQ8rTZmIticUX
bJQuUqpM4O3OU/TY+Bde8SOv5c21U86dv7dvUFX1Hu5NBz/lzguxMiZHEVi7DyKX
7TjqRLNdJYRL+/GQ/QW+isIGJFFcFOp8qdqh6o6RfMnFUsp4b19+7Ivt+KXZct8x
ItrmNdtBeKx7Fe9u3htSY4dIDpkiz8VYBgvmI04P6kScUEKOJMxN3/sC/hhok78D
JY39gz9xB9kzMZ6qBYa5Ya4U60mpQ6J4uhSgeUTLUIavXoM1qUbYqqos3mU4cmgm
sspE/oKnWorGC3QRpvgnlc/eHidybdCUF7qpWqSuyoXEhptmbVyYzPWtIeZmBfaF
LkynOJ+FP1bHfkt65rwAvm/ef2qik4kdMwJ/DbusFr6voFifW+sHwTZQQ0v4FTgx
sUV8CQV98GlH7cQMcxI5d5sDzWgzRrsFojhC4UdbXOWcLr+mvkZ80tFnVjhx5LwF
V5mvnfPCUR1GICUWPK/R8jWUtV0sgwes1sNOkfjFVlQPhBhSHGD73R3IKpmJaahA
sYmIOKSElST1+NjBVTNt+ILTPQ1llnOGVLSCMIIPLg0Tkx1XaBtDpJ6Wp+97DMDv
LvRaBSsZXWtXUVipBVBMfX6HgVooitzI5ONKX+18gtOIMoyn0N2UipxZx8/uEYFE
bvXi9L+oet++bV9TXX04lMt53+ZutM++od9Hjw3ZXoo7dvu/vAKwI/9YueQzPdY5
OHapg3ZqVSjLNeIURUwp9oHUmeqkWRuseLIiXXAMEz/z51R2JHxEYnlA5Mly79u+
B3e/nDDHrbWZm5DHRYgCLKCRvU7vghCMO05mnM1E643p6kBfoRVmMqZ0Nu7WLFC4
nMIfGH7IpySuDq4C/RYfy83n77UtGJc1mkaQ4WUtZjbYGUN9o+WmB7FfW84Gqh6D
SbTs7edthIl1DJ7upW9vT/SeF40RRQKkFhkhqlsgfihGTFrOn5vMzXD1kIQ9+Aj5
OpGCd232mDaCUVkyWvr4mC/TieSqjUtbNTJJMOH1hZ7BSElgCYLtVLvUxlt1VQh3
Nd6qqNdBdxKKVhY/t+pN7xppgbe4YHtmlnIANgfb2IirDtTmyCaf3JdnrV8r0uux
uBZzZ4+6VoH99kjvDMUG4nYz/4kN1FKYnYxBqlEkfoIKwtWote9Y4CmfrGT780Q4
c11YlxXi4I4yKvqDoFbizxIerjQ05F31WBn6nwNx0pvhna2wHoiu3MtkFyd7OaSk
Zi7uMTLeNEx9JDjSlXYLAO3VDqsyOD82itBDhgXqGjIqFC0Oxc+Fm+/Iu07qsa4F
jEXYoJ0uJudBjRW29oVi+Kz8iujGJKzAMKDNsApKxRuf6ycq4UPg8MklKyjtGYjc
0dJsC7sS3Xj1wWucDUDgtUA3z0OXCAJS60jzrHG8LeP6v3kG5WBYb5mO7ndsIkkv
x8TEO10yplnkjojWr1AgRRM1Tm/XWOJe6Ybb5gcIAZYOQ6G4NY+p3o+GCTnjiA5A
0bgUJjm543Ups1jYLkX4ApiHMfmx404ghH2OsobBPwcbkWPxtILUNT5Otxgg5NnQ
Lcf/efrJJMUiV4hzEtOjxzOZrv/EIA344n/uELwpDwQjLahpx4tUaE5yuzZ2QJ94
+/BbrQWizLo7aL9kA7SaTRHxiTtsV0WX9X7DefjtemxlrpAqpYmth15YIgAdpTPj
GgRewvtYitMiR4EcUBbrSQu7jRqFvsMueeOsuy+tzrGlyy+X7nKvAtRLBxI8ah+i
UsUaPMBA2p8lHkLowKa3Q1aJtBT7m7bV3R322ppECoLKKw8XSuBVWgrpQqZlm+Q2
PFzk8XCGgxrGYyGwk0DVHSY71Hfvl5yzlwxfg7jkiF67tGsMy6sy3vFiQJhZDZHR
ejQNMtHKJO36MBAstFuvb0TMKjttLk24fhklI9Z4FRXr+WJ++MtuQ5QHRUyU9wok
Ea/XIaos6JcXbVSgJ70QquoK/sgX7Vwp9K5+OguZIHcIeziXn5SxkjWn87VDSQ8i
v7NdVrUz3TsAjcLosMQcELpF7qLYvCNjYuFfE3Rp49otC0nN+G9ObFfOiDhpwlgc
YHJJwEZNZvUJJXKByHUUkVNljNFmv5MRWWGz1ExKOGevUzQbHWkuHf9LKtjRA8Qz
JB3nEn29rretS9NxYuQu1D2jA/JfaP6raMqoGt87u32gHRf0/mXkQmA/Xz/g2xaD
bSYzq1LZ6mJgDgIoAJ5BzBNs30huj4FAjl7Fbc0Vkv5SP8apf3cgZ69KyUoiJMlY
5xjq464BUAJPlDzCmMgNimSS4UBoqYd15DHUCEr+83IzpEs+j2azJFStbx3kvmho
oMX1rS4V6uPHa6HAdYlp3UEHPPSBJLT1U9pwKNwX20YxAu+PzLhkrLJzIFpg/Rfr
FdL4Twrj8C3i9H/V2q+yzR+SAxwNIWLEaFOpxEnJ+vpHVYdsBOUlUmJQNQV2TYwJ
hcFe2W1BdgujGuMrmmWqMdkWv7YaKERj+Kr3jHCfCCfeQj39TRcuKXbUKMIBEtpA
aPLwE4wlHRQ+GX7Z8RPxULOvZzS0AFWCTx2uiY+AxT1TJczd1l+JDDpGn907EEqB
ysFgUufICagJcPh+UzNl090jB+ErpOhjJSEf/KhwPfJDtAe115XOAcPjTl+xAIXY
h6JQ9O10jaT7eM/M1S/wRye/iGeDrA50UE2gxk7AAFZbxVnSYT4g5JsqNE3m9GkO
dT97JYbaxMwP36xSY7jPFV5AE3+heoWZLg0X10Wb8mAgGwCDAZbi4SH07d1gh/ql
y/5NR0HDDq+IxM81vs48b3mLxbKPLP/CFWULn7ojKVfTNhNCBZ0Cjb0tjLctq0oS
edfOJIudY04H3Wl2QAvcN6SdCq2s0iH/DM/Bp6ce8Ujr1W56b3ZIrXj46qPBuS+c
TbLlZql7NR1nA1B5Hrga9PJgz49WoK6szwVmNJFC2x6kFOFyy8eWhGz8aeG1Z3JG
p4H8nNnikVfpzdIv//oZju7ZQHWgdcScHBsyWJ2mauqJw5nz8ooT0rBkF8yBya4T
zxDFpv4Ohl0DJ8XuIkxoGceaX57SCI8Qd3kuXTS3EQl5rHKz0WGyf/1F4Jpl6tlx
n/fxICmXI80fCSxKAl7ioUGIyb9fW6Hy/S0e6ASDUEbvdeMAM+hqL6lJmSdYlmMT
aflUfQRRIqjW1OW3hvOEQ9aN85429woNzYtKpxFePkJJ7wHPxMxD+o1thLXvznx1
yZHm0ks98bfNI3P/NXVwJjDI14A/f/xZt4h8GrIC+rDf707L9JdgazBFEhk+hFjQ
4vrBv541hDY24x0H/CXPq368FXEXeWKeaYs25vYOWb+zTZ/0B+ZltmWQhJum9hwi
F+udwdq5/XJH7k41h3MCyVe/KG9vve+X+eVYwfkQro43yWgShm6s2VRwoLQPHXmo
+s6s8PZ5Xm7VQplEXt5RcRPD1+KLCKZ+FKpoAByvHf3HEfdkWBwpWnjHWqnpH2bQ
7RoPAcQ/ppLC0NEU1zqCoA9WhDuILvknSEY/NeL0bUvG3J63CnIqz8nkFb+qqKv+
doHXKj6nfyU5m2DVuGhFzGFkK/OOCNvuTMhZDDuRUtHYTDpqYueJFcK/Alkb5Aq/
lWQ2OGwHtdbCp21qxV+TAUNq4xOmHZQCeEE/VlcCyTDWJBYGbKxtdaGXJbbqBdaE
jpqGRT0fzsO3eV1OL4WsKx6agh18zDkatNh+RASlk7HBUP69lBAFvOK4tpCMw32c
XBfRO1VuWA+Y5OgWu1wsmVZouH8zYYGMOkdlnrLcogo/Z/mVRtpNk0syevvCsD4E
YCfz11J6H22EFAupYFP2GrNCHukrj3sE7ZZ93l2FYEQ4T/MRGB/NevZImVjwOYtA
8S5lgIF+3lXfCMzjInUsiPdpow0/JHpQ7SsqOEsOcxbZVq2LOG8h+lM3Y3N8xxbE
OwQ1Y1NEJMaGGdqLvmesCSKu/Qlpit+r/laEjHyKCseuE8rQer9xrXPtLmHfOhqJ
kZlCsdxM1b0jYDTiVl3lD1IQby3OJEAuRSXnDhlq6I9ZskMXa2aaEvNdO4KFElcD
Q4PgHlhjcruSecYgH0bMzloTh37BWwTlec+39T2lu+x/n+IGw3S+VzFlKsT4kvqg
mm3NmkHdNd6U+aYdQw4C1IuI8g29kldu9dPgBIwzSj+j3Q6T2RK3czrnO64UwDBH
NaTd9Pzh1tp+7e0ovcdBQ2fjhG6RE6cj3MUtWD7aVkmr/M88QUg+34FXuRDmjBa1
MKO+X1DMicKa+zXQ+hQ85I80xWtJ+7a+zedVB0bvnqFGmzdFCZh/VudmU1VO0dsB
CpdEG1pf0lpMfYlzWiC3G/Dpd1K297Hbw9fKuDSc9RKamxboRtZkcY3A7t7Jmb1i
ZA2VbUBIlSNXNQ6ga9vzsIbddJiqKh4IFoj1c4BVi/uEPYEEVMReqbHk9OsymNcy
qLFnWNxs1uqq8n3E0JAHJernV827yE6t6HiV/T7BI11Fx3s3W3Kp/0vM2vIYOPop
6GvQCBp4pQcuuDPAWA0CtNqWCnumflCfXyfNEJw7Ap/avoVfdf9O0cLSxjBGxtSg
/6oUpE0F7cPTY0ARGvIcH6gpkmv89xKYhFQpha3dVXENBWo48WNyzOhRzKU/N3pj
fKuSBg+Z6/XfwI/db1NVkGxbHcOkdEJ7vb+p1gJtRmKKac6GcDwSypLu2fu2CXiS
gb9gIsEZfxzzkOyQ5UwoGRMtiHD7/HWsSOl89TyiGQupqfMHjhtvFEuL+xeNjty0
QUJtSrVsf8wAe9Ong9XYxNn+qgHhKFBv9bM5fIvP3g3hs+8y179SHhWQH4rZx7ok
233YGYZ/yUP7ipobhR7HuHmYa75faYDOTUS2K7rA2BNYt1ghutB6maIF03oS87R7
xdNjtpXsRb7qNrPXXyO3Su1Klltg4ScPzs07IYUYeJI9p6LF+tEbOZ3ycU+xFWSe
8eQ69kF/dUswEDtOY28wouL0jBYMEgtmLkhBrZLmNka7YU612b48fu7l0PSNrOK2
LLOpT3x2o15d6rr2lqPiC6zUXZluWQB3bHWiQazA5IUyuyHVIR8atg0dag5GL4P0
Vwho0iTF0q7z79b0xWsCYluJTBsS2Vz390f3gYRKgUWCZ3okONdAiR3lXr/yN+Pi
69Y3ngRK3pWhInt94tpzgpF9yGrgwf0AvubZ3AXAmBHyzzHBSQruh7fAydE8g/zw
L91R7TMw+eAo78dD2+6B8mCfSKTVZvIZxiy4S2q7fha4Bm846qjfnKZrkzDkp+sy
Qzb9eQDldmapPmW56SCDvKFAC3VS3U4pn3qOpuVHACP6rIG+V/UrRvyuJcmdZVSu
IUQvMJR7dUnXuLITNKD6d+gldATc/aX/hpFiH0HbPvWjuuGkrOjcXzQppOgBnA3O
zwTw92xmKDthbuUxuI+INghlOkx5kKOlBcn05nAaQ639RxV9YZDmDv7TDhi8QWz8
HhYQzIjh5ocLs/Z+q6aioqGX5kD0DJLbIXDhE4Vu3lN1/MW9QG/lBiEJInlZkhAi
p++bEwCrSXhG6z2uP7V/haIVjJhZu//Ks1AfZSoWkWhxfSrWYfu4a6bHkKQXot5H
s8RzKUHxKyixcL8EnY+9oal1g8EZ8swGnKiijklbHEonVF5BY2GRn++sZD7sOIjR
iXZtlv8AsiEjd/nWofVey4I3FsEJodlNlxnk39R7/UqHrfkbJ/iAGGen4KtcC6Xf
5GtLfOyOk0JqQqn3AFY7lZYnTIy8Gvx5/swdBiIQzU9aXfADurbwbSAUsD0V8LDH
DlIetxoqY2wekUHe2bX3fZSuIDXCV052W7+loieuemKM96mcbVHciHubOpq9Uhch
wiX+0kAWOVbaAuLlGslMPhh1MBbpeF+fDn8DnbxihXmn/M1+KHeUHYV9QhLxzX9n
tOax7xgSIrGO6hJcq4tm1fg+/6Qxtz0+xT/433PRQiGExcl+l3Fie3OC3+2UgfSW
wBK+WedVm9UuhVO+6z6kh07itvXYuajSq4oqTgb5ASKCDJ5ozNxeUkH6y1Xs9BMc
5YHsJ0lGqRKxcm23kZAFfOKIXzzx+DLGlt6gHbgCGEDBbx61d6uTlLTgchIKGQhS
iDhYTQ6EHMm18DKOLOH/EszekHV4O7M3idn0nxHulZefoD7g4BvGMHqdVLbxpfiS
QZdMKS3I68LkVZ6sVps8/m9xOaS6ne3rGBbuaEzKU3zvIhpe3L5aINjx+S9hXnoX
vgt7JS4SEWdj89CTYgvQ9PZG/10ZZ2otFXbikLrVkgXUQbd010mj87k4chuTTlyF
e/GJTWiIBQ3+TiEK6dLbvDfdhOGL/iRNv5EPytLZpnhn7wJ2TXvjHauz1qqW3cXf
2C7K+FRFyOlGkD+Egby+MBMf3/peKDVtij5WJ5eFzEXOTugm9D59y8a34XR7tPTM
gqeuO4YFWM62vhy1+FZz8ZUuGZdEYzyVZmoULVXtSRhg/855IYOxsrdipTwb1EKq
92iw8j7U7PIe9lTVdMwPTrH03gXQ2Vmhhzvw7ZJmNbaeaHb0zBNICAp6sOPJ8qmw
cOlCiP5xN0/X1YUD7dTLToqw8rIyQmycZCuAfXQadm674m6301GnOmdQW/VIZCa5
ybrJ6lVEXhNQq2CjqP4yD5jcZbzEQ7z/nNXw8yT0PTtjMUU5J4nNydSDtxXsB7xP
JaDv/QGx80FsB2wDmrHZD4uuARUpR1FrhhKQBdN+c0QFo3VQgCqOUN33tj7hUAyw
R/T3oqG31fZ/dT7/6u4vo7gjMezJDtnWHyYIVHMySVW9bsmSS9zauewoZGmD5psJ
RyFP/v0zfxB73Pt182lV8jpVWmZZbqPQX5LuexPRY+uYQtGQ1p74LRyB+UxTL6m9
LWKbAZ347glsfv1wl/3d87rdzDkVkAhwQJ9+7iwIRqEN8KcGsN4SdtlVPZ+cArBw
nvEQw670GNuPN5eDZwLhDgM8J8gsMb/QmxCc9qcJo/Rjvf4zERQ7a+DP9MonJtMa
2WxnOvsIqwD5LnDuu6InUYHfr/1JESoZGP3ustewIBOKOp3KKXnykDrHlVz+zStw
bI5gcUZkxbLjg5B2aX74j+jxVxHFxQ8CD+gRHDvPI0xOwsWP3XnXMInwAIzZNUoG
H6Yn66Rn9IltRAVDBaGSUZ1gJ3VmQQGEbDCoQok17ZJzyMTZaifK+cKIfjmRfFp2
BCF1YWjz3jBTrPhYgby83J6Jqz28j7bn0YhO6ho9PYfMspZR5r31HDlYKlDQ2dcV
JWWMo20qpiGFQlRaMDKah+J4P5FxICZQPSSr1IfHAW/P8YoLyvSUVYz+95WLsBBM
6/VmRRn+pabeA6FVIHjgVRQW6zytcCJyhg2LcaJMG/dpClnMaPsdwwt5MyvYrwC5
x2ccxGDFskiLD6X6T7etZz5Y4vV8hjy2OpNPakUhfK7htvuWXG45cE7DIWRxGwty
hSKi7TV40XCJpbNCzQsRccm4weMM0WEtX0/07/7hWhVAFXsagPEc3rSZbhzibqaG
j31RvzqKXxgWrwTnSfbKAljnSPf/askpHvsNlvCYZlx03OlEtHoFomAVbPctihhF
HO3W9AgSUM9G5/j2moyhYzcvghKod5v1lQnHbsM/046LXjLFifbhfYCTTJTlt3iv
BcyJ2cOeJi1iAPhyKp7w5E1t6OVqzQcAka63EF4GjT/raMMrzlLnWR00NFvdh0J+
qEmNbuJcRvpcB3p6qkY4udM1rI9z4NatFVBWySs5n9droW7ldxuFm4HoyhnfBJaR
yDoi1PvFIlZH6k7F//BbgOfp4zFwl3cT0OYa5ZHd7eMFIkbC102KIpaauiFneJv5
d2YTLI7GEAGWPXCMQuO8Z0uSLSN+jPZBrbbB3R+2ygnN3+tNEV22kZdT0rI0rJ+9
JwUIYTAmqvdff5pTCh5ZG//VKnJMB/V7Bumsnt0YV0PEqFltrCr0eqOqKl7pQVgL
e1cwG+hRPzOL7Lfcqgh4bTV69ryivkTopq+mBLx0ZCxEY2omNTmr2UiEcRTPSLly
wPoDMUmdxzbKZIYeCHBZbur3dC9FRqqk17mv3XUzlYIuf+HhCS2nFFYIizZsr+vX
NSTe9Hm/70GQUOhKOMP/EWmsOwLqaFcNWpnz9E2gXfcNDXreasdYqK7Hq+jXtYkN
Jinun+qKDtKkRWBzeSUinYmYbYk2RKxlWD0DGBtb6hlwyHPmvES+nL3aas2YnBx2
1o8H8rNmJgz2noVuFXf6AfiTShD8Ycfg7hL0lXDAyJINagepcbm8UAS/T1R7/AN+
KMA/5moWQ/bs2tzPZbqnWRtGuSqGiweoyhUdndj9yZpz2M7npnXbSIDVgVMBbLVt
vprSsedm1wriE1V0ArJ7vsRrDhJbwuglPWom8AxJNlPGA7uCOBlYxx5M8VctdpB/
7c4Ze0yDMkOwMRc/mQOBkDchlQU0LFlJitH3Qwc6cmoHp4iT+/Kn6jaCdP3+47kV
eGiKAYtYBR4pmpWAxIx9Ef2QNbtGdaE5KZh++oW3nBU5K4PcTh+FYx+uXeitq7rt
LYbeAq2X+GPkfsr1Lwy6fUFem/wO7jZOjmtxAUTls4JFBS8WMU1eJa6agmZ7vh7z
OCUKLS9+JucN30DZIx2jxLtJdDMxJUneoKv/qEhgD3MhVastQSupH8E5rVzARgqz
neqYjALq0PAJYXqx//7ZtZV2qAroNJ7Ukhjk2uqby2c7QmPHc2nj3gNV3nNVDxC4
DoJ2jStFgl1nTeUHWqu9xr8fqjrqdv35EX4q7qKAytIm7QB3xXtxRf65X1WPJtcz
zL4NERTwMs68wDDU0ssWi1Qti/ZWRtYGApM77Xd92JsFLxSy+/WNQQCiId169kdd
37k5agAxOy+uYxQOlt0N8Cdb5YQgkVk1P5mS2gkFwGOyO0/X4BG6OozoDajmhYGn
gHUJKFhsiLOf8ADis3qrpRqD9hN7VXXL63rcqP7HMxaj55MxaOIojSfTEzsoIlWM
UUte1sKoGVNGg6OnHScivGDF+hp+Bk7oC67Pk7S7uw7x8XI1Gpfr4immP22YFws3
5czeFgsUXUBqjdeg2/Tqk9PKBnX/RxKKP3yrzm8uL9XSV+wdJrkTkaqo+hCcqRZ/
uBDU4hXxCgII6Oh5S7DfBTF99lra0E7XxgNSyev5LtyvJC9orx5lS5VGJ2TA0esI
iyd7aQqtSgcnJoew7sCdw6GNp203+uaflgniI9IKzbIG9FQkExFkDlJSYqs5TY9w
FQ5pxa29yDBlKm83Rp8VLu/B6SIFHt5NwV2qNP2mdI0k1VXqKOmOeK9LHAWbHEMb
dWvfIEgZi13YXWufOddIq6m3rELlIhVFwZiTanpbnfWr28VAT+mvAmll9AbfnVxA
Td5hTfBqMJtfXtuLPiuNfTklL2J/Ssl8kCcDtSQo0+xhZOl++oytq+EudaYCliMp
goUA9XC5OzVwTbeg/pPa/tkt9qDH3XMe1hMYgWBdWVt9/6MrQt+w77Li2F8oj6JU
8lfSHleljBhuQN2EV4HsHzn3fkdTGkUszNrBT0YaqekuUQDWcohPOospcOuLU3Ax
jjQWZdYDcMBeu9+nN6l3oKOkRh1CNLry1Ik5LMgX7NKHwoiatmztbST2Q0Ws0eUi
Py9Ag3r53YiBuOSP2QPWGHgXv0AnHNSB1ASyUzwT0erfXs89a7Q2RNXQgifVPvUa
Ey+vojxv4OtA1FqDJgE+mRNZSoSzogKfthnbRgaufGsKmhQeMHWx7vosmi1OhPKT
oTQpbOZZ64oL2RoTyR/2si+UywxcG7kX1ScgLGV5MwkMHOvbbQoyPn/99dkBIO6B
kXHDDuofcOna/KjGLJutwjSw0fE81zvO8KLAyZi29QhkTahoG/+huDxSPFxDNQf4
ij519ySOL327zSg56TGBHk6WEZUUtGA9tLQpyfk/pG6OS18VvVv1VzXgW7mDtn9K
laUBUbAU4Gejgof6kc7EpzYhlNUdArm9ChV8pCYKI0SBAtE0mczJ4KRYKX8U9cU5
7QDfxLo9hUhcXQtM89YDf0GRyGh/efVmvX45d2GGGOnagHlAlk+ivZ0r0HHh3/eB
ge0gkEPUAH2KuToHPfqkdCzl5NWlqqiyc+I1SUVkAVn8BKcNSAXtZ/p9UjGv1sxU
K9E1ItEgm+sr88TZWikmgsrzizomsBDMjaS+TotylbJwk/+48U6qMwl8ZZfSkMD9
Phh309MT/hug2hDEg06TTQcap5JZFWebfJ8e6978oUueE+DiDox7K3SoO95neOpX
AL9UxiLa1WfGqnrbyy17s/DfKuaW+kOxzB/fMFA4DlXHnkA9mbKBYa4J6qL/ZsHM
ts7vkqUZzAN48rO/iRxNQEoBPZTepbqMrOkusZJmMGAkl23qg/wueT7j2cf5ip9E
npCP3hVv5UlWNxDNwhVVQo0j+8As+UnVZdFnEwCkt4EKz/Elo5JNQTwgOsrSQHvI
wtq7GT411ikTE+EppGPAcbhGZjFF9tuJ72qBaN4Gtb6oOpF9QlQe3m68ZK67sG/u
FaZdl828PVCYx2GiEQj5yoRFUajrcZJTa/xPseo2+pbbBminRM6L7PVQkvVVM8zy
/C3olVwDG96PrM3WhxAOvuHInN93oUsuMQj1v2rLJNUDtaBk2bOa5tJNkKXXx0Zi
ymf9wHTSm4iDCxjj+CVbJyDZTmjutPJVl5BOD7wC8AwrxDl1cb51Y0Abg6PIpm3B
l4Sio/G1quAtdFHtPHjtrfvRPgmN3B8BGYRazrxdsJ0DozAbYbN+cR1JrCarHDvt
sXmU/2Z2y3tRC0ZEHjVJJ97YrJ9ieY0b/E5A+QvHpkrdND5tYVl9SCvJ5G/+e3K9
82D+wmn4ocnKBU52f1neMISHQvsnbBc3MEYc4K9jFXRo+R/1v0dPBt/O5ENtCtbj
k216OxlgE+ZRkeiROscm7EzLw/n8j/6Hu7vwAyLefeGoPK4fTcZljrgFuuWaL4ZB
D936b79ZFEDd29i9ARj1K73yrSQ/Bs3lyF6nehrUjDhqPcpaEJJ8TQQ6dP/3J1zO
4B02uKP7dojt5Wsab8Xzp5YNiSqS/tlsdlcP5unrMwCyW3jk64m+/BEIk+44Rgej
enRddwRYVbCpPz0cOEFmAnuQMVHBK9L1cVJIwfdwvGMhm/x7uWDb84P9JQ3tW/VQ
y9yoHzFg8xKXsxS8Nz0iqa90WwOPiSj5y7b5E0BS27W7h0EWBScm0JLUPN7Q172J
JgSkepZ83WV0ZmOAgJBRj6/DbVeDkXnx7df387vt3L3+jnZTaF/J6Y5n1DcmT1qu
YTordopL564YC+Z5oeiv2psQDpiMOh1lboNMyX7xWHzFaiRsLDDucwGYgRj30QLI
2S7SvAOPAFJAlR+yDHlFPySaR3bVhlaO4jX7L2S9s7Fxv3V1kAdM7mIapIXeV1nH
1UY1y3SHW7lMmTbRKPY6Zcg3lBxXgS3TCTKLZvwdDDwUs8YHCSa+2esvZTiOgRqR
6DIlK+Qn88+AuVy+gGmLIzOTtDgknM1EsmV2r2eAqCtlbgOJGx2+oj3Ax+vNA0P9
QmlcbrN4A6Edlc1XPGBpFx7dKLPR+fkQSKuFfpqIF4qrbjd+fxdKP9KxDXN+Q6Rt
4UeoQBebA7E+zi/lzKgkJIMCMgblwuxMQ3UnrtwmQ9albj+8+DDBA4hv/wYDoXew
hPqd8AnXaTQDQWFbYmXviRdTfLNyHlLmAObOp89wQHVBnMEkxJGeM/HZcg//nGpC
0CVP7MQJJN3Z39alEuQ3bwPvhth1BD3/6cYqP5uCNJD6/HUiVKPNsbV8fhfQMS4I
CTV1auT0DnXgE4HHMiwukjtRKZi6IWoYpYOkV5qFZo3NKUVLUy698MLxOyyDqxf0
HMJqYlWB+GLSPWdyEUWgYwc/+o+RIdqh2wR51/KOJN9JTeC1PkFgaP9xwD2SPLok
euTh6Su9daf6LklyPEtJAEHBZFhCAj6xmausO/BKP4LceDFllZx4oUZVIAYakRNf
KMY3uQdVSF+afrFwhShFLgfpa4eFi9UPJZGKCRAPrV2bT7ofHXwTooS8NdIXpDat
VVdJxVaeAepiUkRo2UBfsGUVJWHF+aNBRiPmF774leKOZX6TyHMh3Q8eLLI2tLfb
XiwugqAYjl/XxwFca2ahg3r5SJP2KxLFdUqYCXME8F4M0somRa/vwog0huYLYyZO
tPHFRD/LKbezrTeCPtM15BYlpQC4yB068e5ZZ1GDvFHHkltVeDaWLuPoeXbbNrzP
JsHBqyXiFmQUCBe0HXBF88fK3tIA6FSpQVC5WLkbzBZ6sDD4j6JE9yAwURbAEhBT
2G+WgPzg5erHieUeHW2BTM9KGwC7MVObkOmnYNVWo8Eu9ArkevanMPrYZVq4pjnc
zfvzNBgs1zru6z3XN6ayQUUfSu7/auGekhTyCX7Zp7eqICMkz5i5RM1N95mFYrYV
f0Yd1dc7+jLs+OnRJTTGbYeMaW2X+DY7MaPG9uEKz2+emTROuAfepnaYc7eWapQO
SHFC3fsBGCklNZWzk9y5Duwcv86fsy59JGp2/DpVihi4h2rCr9CN+QnuF4Z3Ja37
xUlcJ/ArbD5f3Txyc8QDTBB/h3V5rUspmsChEjf7bAdT7XdkIyGirjt1K2YO59Zz
Q7GWTrkg9pe9thR+5qow55A3BYrzJBdRJcxZaqXC5JVtr14tV3LtBlPqvoC2GaZ2
5SWTuL+vNQKSynCyK7kdAwQYCzefIYy31iC61ffr51NVhSRKrMH8xQ2zFXY0FfhK
jt7aE6FGq4yegHJDMgaX10rrUnbBJxn9MYEpoM+tDTZclX3hQqU2THeNOIl1HU9J
DJahCp9PdM12Ilw0fFyiASyP+AzcNrIAF6aVtDSHzbGxtwR8XUrzxxqLtZ3Nw/+k
RYrmLgBRlfgpB66MIDEUnBF1LIdQuDGahFHhlGyN0Tv7cgw3D+hJ8zVrqZr4S+wk
zApW9FmO168NI17WtUYj5QBz41ZleMGAGg5sdsQGpP4uKxo/7xJ2XNwtp1CKr14G
V8ws5aEpCacgCGUv3zeKM8NFuYB8c8w+trkqdWZ+Gusm5hlXVCAUfUBRZ9OhZaI1
EgV97Dt4jXK9rzNxLPRnb5VipLG8rmiB9xr+eNHgbLHfeniyG36Jfh//5You0B4V
YMYXE6isMU/Kuk0WlPYGKk0B707L2t8Y/PY7TYLEkJtyyQp+jWXkrT34+Xy51jLm
t3hzEpxPtNDXKf7FaRe53zQkBMx23W4+LhDflU/ymXJRd5UqkPj213rroG3l6oZi
JBiimj0ptq6wkp/hGOZbqqu52CxvlW0VII+7NSRhDuHsLWe7xVGoWPLC/LIbGodJ
HoecrzmjKj/F2SLuC1Q+wVu1zP88g2/0ZECNDk5py3EF/XiBbSaRbTvJB2hyyhKr
yTiRkCLn0hLsAmwL8VmIhRR2EbNIwFcGl3r1YUu54n4l09ebkttJtbQ/fox0xAg5
m8A+Dvg36ItDmM1itNNT3Xeztec6lvioSgWGg1qKVXWBHgyLoZv+JpAlSTBvpFOz
Ko/du4JudG0Soe9GsgsDIcHOXDSoyHRK1ydkPrt47qzZhj3YGgYbCRGzl/OGMBKm
/Dm0ohEAxgAJNwh8DhizX63HCLHGQ3Kk+fxuWRE0PIl/IkP8LylsOrpQPrsY2NOw
4EstwXSSBfvBLe9ZB9fnDTnqZn34gqwlpnfGSEeXafar/Dh2nxi835W1lsdzie/b
K5sI2QSVdnZVwdigJ+//GcIGjZNcSOiyAM4yQ7K6I+BDtnPGwouPz8Cc8EL3bwFo
1nmrHCXvj5EKv99JpPZnTIiPm/zq0NLBQyp8qWQQXDhedI5NP5lhc4UcZG6usQ0v
CnANShdL9VmMH6fby6ByPjEUF0l8xjnu6p56l4m/+dXGrBUUlNfUDCQToZtX1Gvs
blBQEqIz0OJEaDMV1ufCAXqhQSxUkfiyKdmktYJe8x2ni2rA4x3c9sOstBF2eew9
FkYVPlINLHB9JY+HuEy2sx9qC1qmNhfC8rExszv/ICY9CRDdU9fRE0v9oT9js2D7
Q1d15vrEkqqdJxH0xGpp+x5hX9Ger9GtVAM3xHOiIxewRI6sSbd+nUnqDyELIqlG
nR44leTe7aX7rT30TPW/mKAYvTAbKS1Gus35SzFfhN8dDoMtYUIrtze+lr8JucXe
nKfHetFRlY34FyVvy381lmhbfMfyASfoyXfzFWL5gnvDkvyJsKKkF3zjRpkOLMJk
8ntFzW3wBQV1KY5o9Ovm5XStjPmQQcu0UFA5W5gKp+tBu/41SvdWMHrUinkJvriL
WagXFn+louSb8FrBuYjiNUN3FLUg2CY3Ed1W7sLpnzjRC4SDU8fxtKYtBIH2Hxrs
htlHNkO7jvXYlxP3O6CrspbyosNVtQAqPrV5VbBAtZwo+mH0vjvjU3X/vi4J2dz8
whLboBXT8aaLk0n+iFs2XeugzkrQBuuaPVT1aPqIXbJpIONusE1QJpHpakHDkmzS
9cVMVpqlrKsSPgNOQxRijiY8SaYNSWBH7l6+tVoWoumRoIkIUBmBzlKNVCUiz+kQ
DyshavMgAFMRU6FvmOAaLibSOOkuNP4spUG3SOt83SoRpiouOFnmu4DR8cjK27QI
vU2F68/PNq8P312e+pFMXTW42/BY+cHMwpY9oil20OwxOBYSFIWTdQ1BLoGSXnut
AkXI+Ss/L5SV+fl3+R5FCX+CY1CKn1MrtCxRxRfhH2zK5bHBFmhv+zqQgj1VWh8Y
2vYB4eCAVc3YoFzXRebJd/DH3TCNtZym5rVDx4uPOhHhStNBOr8gxAFLccQPWB6A
AIlUN8O2ozCueZEtKJzOXWodZetZTE9XpW8hejpx1O6R2bMUswwRhB9CkCVo3jW8
eD373fLAw++qbK6b4U5Bje/8e0QTI+sc/Oq9FDgU1xwoZoh3EQaVfZiFJqy3IMGy
9JGIJGTKToYnhIOTcMN+c7U5TzRuCfguxNwGHNb5l7zHEP/IhubXbNK5EmYHCwN7
ObjN83ysTSuYNQhvcnxBt6xisIyN7WO4gSdc/jTch8IGLZRWHoe68n/xFFxe3j70
KztxeJrSZjInWSSNpmjChtvEsdxCMQiSddOe9tza47rrChhOXQ+YTkhYXFMpgQjC
Uxd8iolyZ4+yKqAqP4V5QpSkriSCVSiOwrfJjjE9xVleD3NYBdYBM2gk6V41gqkG
V56ACBowa8cTfnEIY2wSaM9LlDMFGmzZvhBRbTreRoL9NXtntcPzq90txe7mdQ89
YH59k1b9WtjzEu+dEr738Tt3j7O787aa5oSvfYwOJtJglTjFStiZCzDSFJg7U6HD
/ZpAALKhsL2ABF8CsiZOMOMZOp5FV0BenQGKblpYRo8WQNSHWowTCk5tPnmmLXf2
M/2saKHcUeQpmLR7avysnS0fCAUGhuA6D+29HQBwAnHOQQOe2c+mN5rgA7a2WUxa
qi8mFheuOt9o92pwJTxDI0j/phi0Cd5bo6ZUL6qFLiDLAW8epdRNgRsyumw1lgX4
fpVgx7HC0md5ayQ/kQqpuZNsedQ+z8OnDzpRpytPPvM+19dWgli06Ne643kx980E
pt7bEMICWZ+6IMM5ebh3XgTE4wIRllTAyaBXd5rZ6VzsitXPQ8aPgeNivxvfigga
C/4e+vaIoPae91Qj1Ty45kSeovEGCw+B6KVzV8mJjVM8SNKKd8dEJKLswollAD7G
qCEVk5S9hFcigOPZEvnrWC0hO9DpMtW1U0E0lQI5bE8AK5o7lQNPm6m/26I3jY4+
b3EP7YXd/9KyaSoTWRWFCO4BWxRaqqUpqG5w181n+CCmirYfJzAMNA/ihxCygp00
UqxOAvTosrrmhDs2mNdeIIo6JuwINo268ElKHrPHPxZcYidy0aYBNoXgHtvNshnN
nBUjut/7tkYnRJ33xoIPKuSti9068tR6LNBcmvrhGVrQo7Wrrm8Wziay1kgt7W+a
vG+que1BP7cebqIsa4XG16kO8CZ91pAP4vkBLnj1zh68363TZC9hFzBGhP+gCfoq
uySdO69put/4MAGnse+kf+fNfJcdK/g8zPvtYbrzZ3wlyNSyx5FRLPyfu0cs7pNB
yDzLcm43eyzELZAR1imGXAakKH1Ze63Ej3kkCF0yID7mNMmYRp4XVtnO8uhtKdw8
uBKyjYICXwslfdac7+bJZpyVclKeA3+M1y57QCBReiNoHWIhCe5y7YmQx3KqRg3I
v8D6jjGjIeRpeJW5Rx9uNQYS8NXEXxFr4FctGE+Y9e24s6+u6bg4lZwNEiSy45IF
/hHcVF3fWiyXM4WX4I7/OBWuteIyKiaeZJ0clvgsNuERmmQdTwqxxLRro/p3xd54
GRlRMSYBiirJWWbWPQbn7xM3Np7ihpYJd93DT89teXLR+bxQL/HB0zuyjfL/vGf2
ZmJxCj94/7GlmPpY1LdviV7y1bHPtY8aYeUvOLP+qpX4rKZ1m4Vp0+IyhkxTPCHa
7mhfOuSIoa5XjhoiXCPD6ZQgIhJrgooJ9EbYBVBexToxTJKi/66g8G4gvDjKNjbV
VRTtUnTUgVXagcTk0ts11Ld8BtqpkpYLtMrAVZyoVUUSGMFa5yEVNU7Nn5eT9yxB
K9wk6OLD+YPOk9oPavtNBo1bOae7jzz4vsoeExJfVrB1FLdSPvgwCK+lfiOTeBt6
C7JhPjLJUfoFRgZzlv868/1lamFmLoz6SGOzUcInYVDPR9nuW9FGkQWd2ovT1QGM
eb9knqogI0uPxsenky5WM45OdinntZdTd2669BEeK+T8VgDIhGuTP0iq9Lh92XqQ
3I/7k+o8JxjGaxR+0JxWLZQT3dVdC8Mbp8V75AFRYokO6CqVNY+tKyqilC65xZ3l
Z+LiNHHBRUjIspXad37mEt9iuCy8cbjSiJMVxC+eP3WNkmxRw/cXauFZGj00AD4c
bN+UA+LWRhcPrr9kb0IEldXy2LQFLWvx4IQUJdGdsrojrR03cdBSDYXNfTqgBlEZ
v9T49Nl3giRSpe7MzVRl1rbV9hce/iCiZMseIGcKpaHQC6vVQJTF5xeaflUHgivj
OjgHoplU0qwQn20ZndBh0aJtf2KlkX6T+FtnIRv8BLwv+josQEJNoG0PfMUnVKhc
kyeHXlqXqLhGW3hfJ0KVlZhbUZNgGj/l9XRkm0HzhbOOvIv9bIIacPbX2/Mqzabt
yzD4rX/cY06GFn6P14hQJ8BdrurAigLcaE1jBAlpEtdBRFxXx1tJ48Qo1y35sA5q
NEZe/lhvk9ZcjYg1DM8ksGeErmJ/BpLByv7SmHs+WEVS7HwLlc7IDBbbf1idmKlG
61l9x5h/XJ/7JgsaeAfrz6o9ppyfkTZ/V5aL77t0dQWNVFrBDvTinFFZgdFa+tDV
jCFgqg+lWcM6nRV51uNKR3Lb1mYisxNnA/+0fkVpktZUFsRqHG2o1Wam4UYMAsxm
3grlxLMHCvLJLB6Vx4RULITXIChdO9P7RSKOWoheusdZbnWWiyuw53ZXy7RMNpdZ
8pCZ4mUdID+aFSulZwRsVXfVG9eph2c2Lke7r9RWoOIFNoYPO2VjAww3wOVZp2Rq
Lbk76t+rSgvQoKNsEtUdcsYdz138MZpbjqWt1GI7+oPePMVFkNtmAQlNn9qY8tze
BYSI44BnhlCYxU2AFw4d+iY+BWcMNCGfFMfFOpppqpvgI0p2sTSF/CkJfA9j88u4
ntyBufBH2T/a/dQ4ZO6M9BPyDg8Ir6lRdAEcLhv2jYslZNfOWfLwZfJzjFkld4We
dmPUXG4q7a73L9LWCjEVcxo4QnfvSJwO5rm5kzzL63b2Nz52Y/i+dhoFDzcl/Ybh
OoZuwcWHG3UYkr1m9wddq8juopEDkUvmVLKfCkEk07RnMhQK+BUmZxONdiY0oiro
d30QemuEOA1tSRyfTQsmgav1N6xhEWEn3RSFu0aPxhBQa14MbpqcWgleNA2dRcs7
d34R4Gimm4dQO3N3ammudu4iZHY+A5fazFmj1orZJpQrdxe7Y2vSJFtbWg6HsMZZ
Yf6dTMklkITrOgMtQ1Rm+JaMwQl8C+w6RFTXHCMvfBHugLSOm1IrUBLSkMA4BREt
62HNf/g7AWfzUsy8vDhB41tpP5v0KeAoVg+1EKC5znX4yP0+Dgx+9mGTV3BPVOYH
w2vJAAf2gpq7JJpd9FoPLM/Qy8SPd7FXjioEPN2w2LNo3pVJ32oz2Sd02vudYdFF
W4AqjnoL66I28i9MQVcvbgE3fwu7JGXY7MLiinNM8uhbtn7JgVg95j8ft0OVKjxK
dOfdvp09PCvpZjXsYIx18WlRa0iojgxxFjemMjNIlTWA2mUbSNetbxOJPH543X6M
5okGi9Z/DoNAFTljk3YzVaJfJPAFixeO6S6Iwp2jF281PcWFZxgWMTA8ztv7A8Lr
fT45EyG7hGE9mGrYiDscu8yOYfq9dKL3nrQ5NmyuCm4K2MSgRVC6iBi0Xm5T/6sZ
xuZY+WX01P8d0Bi2TRWRVQ7kLN0oixdlNnWdImypfmgu3zomTAobPIUrgCfwUmi/
dvQpZPlFRqdYxNBrWwMEGsDQs7+MbCTFeQRoeAm1CrppitcaJIkwxhS9RSTTujPw
38XPcnsxXfyPBNQalL6xZITDaodnFhkekLYXR5nvtrpqzJbx2k8UlufxDy2DFmiz
bFmS1zjuluA1wT7SfIb3fbNyWvq3l4UHhM+HfQfk6jLPYWkYgc52dcnb+LnC9/TL
g748nd/9GZ5l5jtPOOgFMkgzewS468Mf63VMoqDJTlCDOv/PUlvur6p7TxtGrmVh
p2+EfdxgIJUEQZWwefUg7jiEHGDotibo7ETkRum1Y+Tc4RHu2JbdtnEXk+agtCre
Y8F4xnwwmCUl4mWilDKOA90M/kSTRamMOBN6ko2+X8KpP3alCIy7JKB21i8LfiOP
EiOOJOCqJlMiw2wQzjr1CijtLI+jnvpeQNevKOcnWslAKxhhF81GgMdszpiy2Ni1
gXjc+HnTa0RjC8AHVYdARedEt+VSHoByyR/N/2JKQRvL6CSvRYTftYBGqvOkAuvR
KCduDemB7aSz8kmFi0yACp8Y71HLXKnCiG3Chs+m36v5n+nLlE9TZTpsYRE5NRJc
SKE8casPSlM+WUIZXTKk4C1Xj/bJMHRq2ao4X8UuENuA1lDHyni0DOpPWlTgn/TQ
isBfVyPyFjuvAyRYpW/9xiO+Ne+GfwTWpb4ah5XUXGOVbUyVDX7x0Sa4ESrGQq/k
c4e5sb0WtxVOrs2UtuadCPYzfRfZcVgEG97QkdAuf088qvRIzarniGpCVkckE34w
9/9KnYx7YtBVijZK8XOS27VQomCYJuUEKpCb9tNXW7yj4OjnU8+JqL7JUSVFkH54
jtaFBrrrq+f10gWWIbLb4HPbSSyvGj/EpPHsnParsMjHGC7OKd/okxyPyyk3Ch5r
MmM6WQYE8IHW8gV+FDOY2XPcBOkuSCK/Z/j1lu5w2XoTO17mZ6RJRcmPdii/Z9en
KuoGS/pA3rxw9EafkQQ1kY6jwRDelHagebMdCApzYGRhWuV7vM4Rd2Wy7iUKt4D7
pHzW7iZl9aWryK4p6M6Nhx9MsZW+AWTYBFxqOqYXvNKk5IACaLRkSb2As7BNq6PS
mkVr8j63OVKoBDWZiDbicbFBcK9CzSa/fYWp51zByLKmvlh8Gm1SqvP5EWTPoyBH
lybfcRNIgjWGI8AVg5ovv5Ozga3kcMsHfj0k9iALZSUt0MBlBKARnm4Xv9FO5em4
SuTWmsoZJ/KH4VDg6s6QVS3xGRS3TQgNyMcfvGxBOx7fbfL35K4LV7P4eWGBd+fv
6Z/iODe8GnVqnbSIGMUIBVOESWdB1Gboe0ZgzHxktHGt2bIJp+F96VgTo3JfGdEc
oJH0sGbC4KH5OihwDA6utXidNX8B9rH4/Fs26Uj0dX/DtEDfcFGIOvsSHayDwO5W
LXYro36UCZTAlympshGrIUSG2n/uzQ7xWWdwV3pmrRgxuM+m6cVFHUVvflsKQTDg
sVlNpSM+rkGzdI/7kb0bfFfe18oR7FSH16qQdMOLUYlBAGsvGS7idm/HKe8juZdm
6T02QWEBYq06QPUiKESRDBMJUgrjOTsF6oqaDAmbc/1xt1+IFLGoOiNYOJMnL4JD
cZABTFTpDlcQ7kgK7ESR69T1JvuWIqleQZxlboBAkPu2p+rhbOBJD4QRDdk1kRyr
vG4A7VV7xqY06QcYoaDncYdxPHgt2Fpjx1rJXJfL4A/j2Asxz30ojvQ1EZj50F4U
tja9uwSFMbuPHyHXWQJhhqTUlF3zCTDpmEK4K3663VTfka1BdNEa/sWgTlMuDMlt
gon5r9bguEYGptW8u2yIaozPnshjmmk6w3u+kBa0UY3ZNP+Cf/QrLHWlaz3ShJEg
sjr51PSTVf7c5xhIBsysXD4JMMCevZDfbzwt0A8E7WQGOxL9i03XrIyY+SW/6gCW
r+SEvRE0J0nexmcd2g7QPerTOhmLVjgT4/rvUoPRPuG8z3Q60gYodP2BWGxwq3xF
2UpkPA/USBQL03GYzpYdNmVc9j8yGFaao4lnarrtNe+G5ujaCqbe0YQTRHjMGbaw
AlUsl+Sq3nd2n2Fnv26Jmh+h+TDXDweD34iFYQUj+jGymLeY+m/uXv/FzKhtU5b5
NhBoKkjqTWQlGnjZU7ltIVPc3vcCDj9HGbod+U2SdxKG/XoYHWs8vzs8QEBzSYpN
YEQm6yAXjpgSTuseaaPaPstTQW2+flJlxOBCW7VdQeBhehhmYuuRVJTN1iOBPDJI
6uXsqkgrv8Zua8Od2igDqZkJUilCVe8Eq4Ezy5ryyxmVODqVzyQeHNwt0CzBEAzG
E41AydgrnTOSY57Qe/MBCSxVB0HSjWOWP0lmE+Apv7wQKHb/7/pC9vol/BmPBfit
STsh/SXQbqqWa10ybS+CcTPssUxaTfcNyw3yriA9qHOmCWa2tZ9Zbl8WrejDQ0Fd
BTuiO6NU/qAzs667LZg2G/vXof8awjBUYGhG5szzwMPkJelO/h2qdE+fQnYNeSm0
r5n4I24CoUvLDNH2MSEK+I/+XONQ6a53pK3Ut62S9f6OE6qrb6kZb//yiDLQEiSf
RUm8VrHgGVcPYaehBJPNsqAj+TuHuZIGIV5faoDYNeTh93wr4887wEg5GdUvJ8Xq
ZDlNkihc5WelTBkZJGQI1CBeliSZLfelRpNdMW9PRsxLU2uvXaC5UfCa9GWi4MY7
a4y3OMWeI8Srr7ParDVDdvN9IWJxMipYi9onkj6sle16iuh5Vjfec/Tn9w+BtVl7
Ad8nngB2+sjVuWfpV99p0GUDgfAm7tNi8d8fHBw3U1ZN0dVzHOTO6Ehw0JgzvKCo
eM5tBDr0dtg5iyrMB+V4DYjUOU4JQPaRI7WLBfg9X5p7ytD5ZXzDE8nnKROT0Zel
kd2TvtnB6UbIU6JndheoasOIUnop+1z+ZqCMhPPo+0mKDxapAplrPfqlci446/+l
AWVDw/rmT6fzODtVpAYdNl/RyFR3qpWSw+OHMTCYjJ7e0ZSzmZVr4FAhHTQBSndB
EtweJ6aFq6pooW+TNCg1oey0Gdha36uvXP+xY4sOvacDd17uzE5sFN3bEAnnkCZK
/RPxtQ9dPt+LYtR/UMcWtWkhj1pPe1aIiK2UgURMsE8cSq10JVpLsceEuziJIrhm
AeYckHPZ6Vzu9XeipFq3UDUBwoXOkloR4MGc/rw563O9eN8Z6nq51O16P4ERLul0
OMUIrEfjJKy9Gatxb9ZA8rXMnWY0WKeukFwglOrG7scsCOKDK56YGPjSUAn1JOoC
oJCELDbthcwD/XHhRDl0oqx42v0O1q63ikSttXrUxFntMx/xgo7qK66yn+3GBJV2
ZN+rh0rtU9EBsWkHVDEXFw3bnEH8EYWlfywJFArdjcZNyVerhzLyd75IhM6ilSGd
jaI/UDNYRJE6rsgDKRhU5iuz7bImeMc8iIGbtOBk9vfm5MVdoZnRiT+rdJDNPr5N
MipJIXhEsSKGJYocnmXJ17P2meH+lG0r3nHtgS6Xbcaw+oozoGw1LVvkpw3Y5FqY
9USC5JGRbQJupJH1FIBiR/X6ZZ2GHbjyowMtgLg8D602AQWVVTpe1h36pdBhJG+3
hpOwOCi4PD13fSbq2AtYniB/reLrfeA+M7gQTasdoEECAOSDvz+r0CCvBfxDnzQQ
zI6+Vl2oop4gARX8KSops+mFvTp0i8OxnBglir7txgo+9PEXyDD2jUyKJDbfZWmp
otAW0XR0zdTxvtPT62njDvyuKy2AiL/CEseysStzqT5C/qBqS2KMO7ONPZU6Zjq4
q5EYcye3AgeDrCmNi+HkL1gh8nAEI9OzKy0UP2RPXx5hr9nBl9HAQYIRQQOwRXuv
f6VOoGrQRm2Mbv6S9voCz0s0iTbNbtn/ZX8HZr5mOEVaoKffax4Uw/WOm0cuWbJD
C3OpacLLVB9NWSuq7Nl2qnQqR9943LJk5h40DaAx2qndvWS7nD/sCiCeScL6k48B
51MWvKiY1tqs0XBR+2FkpyYluvJVh5HQcxw4rrY1xSkE2q92zu71gdcz+XsmqqDn
InxZmcWmsLR/nwYoyRLAT6Z+PQj4YT/QlMy2LtyoA8KErSWDPhNTbguelgcHw+qs
AfXtIIt61DfvW4+tdNx0PxbwH446clvVE2abChYDfVVpJ+t3nQA+2cVQTc9l8/FM
i/MWwhk80VzrrSqG4IX1do6++6gmyhu9qQaA88t7q/v1M506CyIQcXebeoMPrZZ3
gOErLuTxSgGgs6CtEwu874hZHNONX9gh2NCQCkFXnh7sPC9UAIqD2VYoHhQaHwC4
tnfZmGxUbvcbAQzggJD4GZ/tyTVx5sLBZDyM8Hys1BLiG3+Oz8I5/tAMHfl2onMt
PRQ77xE6Ha5wtumCp9/ooTFlWAypfPPrK7CvruzXYYr/SLMnkA/gmMQZNySDvxjL
x5kWR3x6WQT9+3WcQysJlv3kQL4N7A6KQS56Bx9BcaOueU8GRGXH8qBEXfUFdhge
70dmJllmLzkkjbn9vI7VOIi3qXvKUpvXX+9s5WJ91yBg2PXr/5lUsfvdhXwm7aeH
ECZW5g8UMXQPqPzaSAmZQecqhyAvuE2DEVbcbZ7v1KzZKQ1ATw+pusLdxIzmGGOu
6ZD832Mp3FaLjjCrI3JoZHbD0+bYQ6gBGBFX2+bUhkXUh4YNI5LGsixRxbxfDljH
LQS5R8vef5knJniYgXVkKrqp0Wf07N5P5B+QY3oSejF5cr47S2Vr83Hmw3k/MLIa
ASl/fEVr5RAIOmBsho1Mphg9YchGutDT6OIQnctkHhDUMLEGmuIypLnycbAsoXBl
Dye9gAwmHU6slTaHMpTuJJeqzpJF3jod6CXE++ANxZqlzLH1pXRV21bIsTIpmhFb
iaRQPlJciCCZiRFl15FK+uH30DSvwE0ia1qKajsB08eRLaIMN2rCJGkh1oWA9Gip
iFClk3EAfSxUhWSukiQOSXr3guLtLRL+US0UcAe9Za6Rdtg/OSSF2KnLrV9ujmne
QDeIWUtGQLY0Iczx3XoXmDFsjFzaSXQ06XgOMawBIk9HJm5KV/UjK0ICEEUdRjot
hDxSQP6v0v6kqqbEXvr8tf83DoQjz+vCMnkKW69vLSfvdh7Q2dARdPtWX8sADnKS
ZAXg/qeSAPMNSduJovjIZOT9ATk1wjPvjAaSLBLzBMwZTpmSAWQFMCGaodYONRb0
4WAYGZd2xMVCql2QrX7CKZNWfxyb73EyJXDxOISJ0BNoqhjAprkKKmPsTgiao56U
pP76zDUmvpwSAWs27kadhtkT3CNh1mNFai4o5LdkHMtC0+AWrZnug1SSXPUiYlXx
FPUp2kHnnTd45ffY+Nf7LMceLszBv60X+8d/us+W2NDCZ+8uwdjti4lnUL5jG8T1
Bri8N9kOwzcfuXFAjE3E3hYeWf8STDQm4KuzAWLoiNdW526dSNsQom0HxjgcBpUl
hlWrKw5YThdq9KVuewdiBzj9LM8Yhv/P6cpOitkAQLAZ8WhPSC/3uBVTNws3u/Iu
ZAjHSxkfJU3sR6HJH5zPCKBWx36zqyZdmYQsCp3Z5dnej7LJaULtJmgaWL3CK3xN
EKt47+auOZgpHFxPy4p+3snBl+m91EK7VELcFfCbC8sv9ZgR8DbKSA9H3D9xCmyj
PTcPahMwKWFf40t1GVQAiqGMPpSGYDNMl46Y37DZxVIDLto4lmJXYXms59nHHRrc
YTzT6vwol/+0CEe9zspZxvl1O+79746v5G4mHcGudxSMa/SOcbA4yit0MovGy5P1
f8oHLR9yTkk2XAYwv1fo3IITeN9USZ9zUheMNAa0JNkyWGqFQKReBEDWdijIA/Y0
R66Z4VkXu/UN5mdwqj/oOyNvxvPei6tSQnCXelQ77DPlATgxR8c8UHJ7NECDh3eP
Vykfnbz37I3WrCCKsbmq0qdwX6WnfnaWKrm65sYZTXmtl+bP16r0ZCOLbe3SmviS
md3DJae10F6r9lkOE84xYGGzmll/IknMXEpGVvXRejyP9a8F8deiSrz8z5ULSX/Y
P+uvWRNpTI+QZmlF/L1PzcD5zIHbNHNLbJSeoOnWmYlVvdvzXntSVDluEI4sFJEt
h8bEvKpsTjuV/3c8895wThiA/sxFCZI3Hhw7frmWFANbq0IZCH2DkQQ/gV4pqJxe
lWk4hgEG/5umEI/oIik+B7ZMm/keX+XTRaiuxPpEYW1O8KWyJfuFvm+uvLcwaG+z
/ov4L8yYFhlECuN9mpyRhgk2rWb56gvErcaL1W+iPbDD9VIYQih0/fzW1CZG1Bvx
toFd4gvLjcN4MfkPNgHJ7iF2NS9212TOJoVpCfHkoW/ppc2Xdf+IcMLU4P8BRQTL
CGA3oKKf7zIuNceiS1yVloYT2IDjYWC/rpsRd7joQV3s73gpwev+Fc+oEwZgBsiX
96SkTw39xl+mm5ri7v0eDm0HjGDyZCuI1Am1VSBopy3q/1l1gYkXYUdTIzpnupct
Wy2UKVNP30E0bFNh+2Wope0KFJkDe0P2LfSOULVoV7rH4f1759SIIpXR1q5mYJZE
B+OFQ+6A2kqguxEUAKEnvlhqumJc6WyIaJE+BDm4aqSanpnTw5x2gbJbmumOpc3T
eymNsBNBzvTn87PvBGD7KK0OjlmSiZCQaQUHNDkjoIfoPUHptks61K6wrbb7nSl8
RxAIXp3jlkvzAQSVajSFuXSxeHfmCwAwE+UpR1Mw0B7P9IGbi2pONHSkyVBiFgFX
NI21GUCXL7LCWd14q6Rv+g7XSpKP8QUTaYrqezcWj39MXMufsR2RoMWUw2KS4217
EsWW6oSKsxrPpi9J0OzcB2MxKR5aQCncMQfWvYx9RwZCRFKfaJnWcM6jMox3xzC1
NRsaFUKqGXYYJpw0tldNi51fVwajoUOkl+2DyY5e5ke1gi/kJpS5e0iLOIqKn9Wg
SJWLFfg40YHppg29t8dxSyJcDGu0nsmMDSUGEUKqSsTIS+Cn7aoBT/n7tWeaE4Ms
qYBpUvSCgaNu8/1ULzp27BKzBScpHj6D2Jkaxf0OfpAB3axCgFwm8ooHIlmNruij
cM8u6dNCWH7zI6laePce9WaEdWBqWeqvfUqaEJr6L4uqe4K8j4dWEWmmuUzzXSCH
gpErB9S3JCvbWBsRtH0FtW0Xzx1pc/tlrEcASbdCY8DNs+0wfZuOITBGL81xmvl6
8GKwCecv4NmaKLg7iK7tPcyLdcvRDzvwGnaLNzjGm6bMzWqgh0emJtQVjKzBS60V
cp5Gzu69CFnIXUdzbdm08KFY+i7QWp0ZyBID84qS8oxDOlTZOyfPdn11OgJ8FSUW
wBaB6lsz7Gh/DAxFxOAKJWBaSIx8tlEpP2wVXSf+7xa8NGX/DXbyBZlHgo+J4TyX
K+EiFOCqU0xeQ03E2VQfrJDXEV53hYeGY71miEsCL9sWqjprodIZzW8ZI/lTHeWv
yIJc8lqGDoaSBhSuJCzaj4pmTDzQRHwsGJ1M7f1gn1jXEAUnROd/7osogUOZfzlD
8xjVnmbAOkWhYBbDclJkDAIFwUsOuyedeazsR4lXhGPhtZGoOLdEjx5CSzktsqVn
/qm3VaOJ2Bw2lm0j0B4r5aJoxHU8u7m35DLGGgnxECh4fUN53c28vTDbT4wxufis
jp83cyNfGHXVLIv1A6BHC9QmiirB91I1hUVVmkaQnbQGInI+yptnmGti50efu5wj
U7QHpsB7ANMm6xzgxApn/L/gRlEiomQuCktgY4M3BECZIdj5E3qgJg0n+7YnkSUH
IvbUl0FGFlpGMgRleO567Dcxk4rm6GqdJfHokF2qvncsjadccb+beiIOQ6YCvgmx
KTUQiNZdJ+7WSk1MNbe8RN1nEglEIaXaU+OfxcAM6UiuWEqTizEoyoN3tQh/Ftcx
00xLicbgUVTk8fPmkbTbntxl36xcQOWNMRadFosKzAx8nluGioUctLn5gh5/cBQH
rTXk0YIvxdvC5UBp8geIqqh9vASCNtppQDlM9/fX71dcPMIGLKPQ81I/DAhDG75w
K+xqi7ES9cedpXoWktVaMPw4flH14y143i5Oqo6ku3Zas5xzEvfv9kcXF1VvF03q
0E9xnOw0sA7o3xkwfWxSHFlUxhcUCGhA/fdCJ3FnFfQcbQXmcC3tumwaTTURqgnz
ZZFLUU+j9pTLVG03+BD0vw0l5iBdvA81c/n9xvsf9ggao6JH1p70NaWyTXfA1i/P
s5HKby1AuQkoLRrRkWNTulerLhgErHqyzDpkGNwHzeRIVC0bgNjwhYSYUC2w8f8+
Zk9GLBlKYxKPDdEpqxQv+ql6gSbf2XtbjRXOdwoXH90Nplkz4VLZdJo3K4SVLqbc
lcISslGytEBW2Xipt1MQEtTpXWWHJ2KZHgmvLZDPaedanmPbyZnNxHO5it4SjGjE
ii1dmh3PS6yWy88sBBhl5otZFx+jeWh4zMKHWOVxMC4ydQrzRbt87Asg61b9izPy
SNXrz9aAKTYSA14oCCKEDN0Hz420eMPI88xyyfyObsGs3sqy/d+C85TYbwgh4wws
m0WVxDLvviLvCR9CroP6gLBN8mgUmYIz5pmwlVXFnsLm8aK2XmKELwGpKo5aPGkU
fHhmc48KTrd9NiF3oVwelMjEufXSciM4O1Kz3hQ9FMr09eCOLo10eHWauTAf3TVe
Pg05lKKbCErTT51oYC0TsKVgOZShQ6RlSFzJcKXcDLUm4UJET5VkmgIq9kO8pEGR
Cl5kv1spsDc7todYdyaGXk1XCbMwJqLty3rkz88Z7vDjOQ46aHoNGJ6n2N4rEIrE
QEdZQdgxdINs7bOz1kZoaDaErIzWcRWMYwIPgk6i09QxzXXcLn7UOLgyIAvB4ksp
mMvF+0VA6su/lX2cPLxgT0gLY9rb2sZZdRFjegsJYVwKxTZSEnJ4fbLChIKUhGGV
ezzcWgNwhksVS1HPCDqYhgw1/RWXa+rpPStKXOzfaNReG95EHbA9wu6AkHwA4lIT
2cjrILWd8V/to8TkC3DGGR7iNrDwKj8suEYScFjbrZkkHIIRzbiBT3AaHUW6iL8e
mOi0ti15luKMbvIRksyxxaYcGS+U9Si7jmOMmfBBVDxoUrPIBK1ifqek+ZQJk8sI
j7R6Z3mFsWRe7pcFmLyBJrarpMC3EkyMzsfh2feBFH9nQ+uwaui+EhX/TvoD+f/c
2zwuIn0lD/2zxKnD22lv4qhBO8XDzJvLKn0jA/xodffdNUzw4ZCPgi7gbcuWBA8n
PzPDQNpltogt2BMrFbK+0msYn0hm2vkYins0yCRsvGqcEJfRTO0ChzBnzTqWg2Ba
2wFPrJJfZaFbYsd4MgSt1qCw5TVeY/o1oCPynflPLYhTgaEcBINvqlMaY+vEPH3w
rcIk82Vo0LL9/JZkpyu4zAYqJ6WOXw6aKvEO7l/s3//Jidnw31L7CJRnkMbjnavh
H4ER3eSgcQBBRuMrgYD1nug+zVxkmLqE3wsdbYawku1zITQHdHUQFv3SEZ0uQmgM
HDW9ZaurMGnoJseZtIC+2muSz/8JNWZBVsc8mO0CveMGzv4UzX9fyLCtDnNrClRB
429TiaNluFcPguoy2OPuz9wMKwCMQiIQvA59pxorsvSfnaDoSXbgcQLcPJjMDxpB
lD4yC4ww6FVo19f5Hkj6NzsnOUK5SnLKcDiknVz4ZlR3AJEXHlS9zVoj/cqWHQHL
GAis6n93OWtOwP5b4pi+SDgCArPYa78qU9m19Mxmxy7HtBjurtPkUP5EEYpa0FR1
SJ5/cnOQUbPEbPi5bZ0dNMde49M8ieawfyJbqwF9akhTwtyEMwxpg6gGxyTJr/fm
u3h76SWbBQBOUYeVMhIIxq6xAbsahCsFDflwblkKxbY3g7bIol3Tj9L6WeLb8uqK
W89+P+yWnTL64yA9s/KdwvSet3GG+VPv9XXt81uk3ebuA7hDZy4M4XYLakpIB8UZ
uVRvEUhw9WDvCZ3pgO9YuIox1miii9ORgUGWtAhKvjYBp1fKHcLpnoO3kkSpsIi6
qTwXi+N8Wd1iqBzcz3V9Y+7+lHN1aMmxROvFzCpZC4j170kBUABwVk0VCDRDKr2W
9kly2tCFQIpKNJ9XFX9Dv0J2iWyXqXkD3mM04ZNzeBsDGxXAZVLTZ9B+daDwv3uG
IXVQoSV8ySvQ8u/QygWYnBTNV70fMomQ72mfU0KOyz95EioSlOrbtYSYxi9bRB2E
AtMEhd/3vLRHgHJqzOD+5Mk2paGMqY7IlM1XafYUjFigiERLNLBbo5Q7FgvDe3Qh
80Z2sgRr2zzO97VFCyQkQHJ2gC2/1beIkLM5mCYtbgsJj7uSbR7My8qrdj4479PP
eME+h3gz5dfdSQgrXi6l2DXs8NvE1abO5uy8j0Ej3HeWC85zdVki1lcUbD5UZo75
uiFxbrnKTU87ZSuVQTXHiXiuidTCMMo7iPrivEXV5kBj08e3oU0+sh4TRMXTR1zI
i1mXHm1wJHKIP1FyjlGypn2QqiNZLv2lXruII949NUCLmxSulgd6ynTJdHg7xst7
mx03AVS3lZljQfcVzivRM5//yYeOJt7POZRKjh3AZFAH7qz7B+ry2BpQp6G0DXBJ
/jlGMd5pxV9whHEwp+K3aIfDl5PRXsMDUj3m3cmDIoamF0snmoMRZ+rduwrW8G0R
n0q/2H1Is6mNrPZX88Niq6ljPF4z5qnftnBh0v6XlfjRje92NixGgem6pOBbzjVj
VslLShJf3et5yYBZy7HaHKapTzWSqWvxJe/sEog2sGQrD2HeGEkeojjhLJzALaaZ
G4Frte2R3Fkoy22T5qwyLAJ2yARE2sp63wxzOFUjbWqPSXswil5VsKdxeLHa9b3T
8U7LXurYAyqfdvgljp7FpX3hSV0/x1FxcUZovVqZWksBeYnpE7BAyE8muA2M7CgJ
CXp5f3YLcYwin/R8Riy5ycyl6DM9aP1DONSI/+6118ouqi9xVwx0CtYGiRDh6X1e
QyNqfkIVLXypOhfr3ukKvw/4SOiZ1URPx5Z+BlMBHxhRCCZveE9B7hm/W31Mmv/b
cSy3DjCmonP0wNfJ5bEI3z0nobFr4J3GF1RUgK3i4q3fNtt/eIaHulHzbqCJLdN3
MDb3T0DhJgH+AgBT0gVjRY3eruiCfLlCRSesKWsi7v3vcrIqgDgOLZyyYfbFoSDl
LAos9GYNY8SL1obIz9GdYWRxawYU9ygrbX/2B1O8AkfH4R/fINh+WCJzJm3puXFj
cI+JAwYhtZewsXs/3xvZYZPoMhcAqn2pG+n45MUl3Ft9Y2oD6SzPMf5+VJDdZ6bT
dpxWYayyeaiAfhVCUgYBHXXBFuaTq5BCBTXX+gNPYUqrXui2u00l5mz9a5tMhaig
nlYSE3NacE2OCYBarqwojbL3TTVNpxzEb3d04Jrz46DojstcpKXXdvVE+63VwKnm
imJS33+rs/DDQYMV9kveJWLQfsCBNkUv8+xKhgc8EEia1iSZW/4g5SuXtWOjoQQI
kj4Ja155CxJED0xXBT4Zj3E9jZfFkYQ9RJZSxsaTSi229i3cVgP7oNZJ1WDRT2Ln
OXCCBsW9aOpTwKfkO3xlRu3d3wGcY6m6x4S/5fNbB0QnjxOS6pOEnFeRdkpoI2JM
we/A6izu4nEHeZUOASRcCPt2u5G44arZi2aL5GEouX5aYaZ371e/btOk68nIC8Tt
G4OZ8OoFZ9C0ai/2CoBlnSemovjPKd9Qg/8ey8KIi67pVR2mcm5A+WppEvTpMim2
zQo1TVE2q6tPxhIHU1XNMxkPsjTnv7ipXUc6mVE2G+b9wRzebtE7MgXhxDypXMUN
nxawc6GzlZukmet3zdlBCB515Rd1lCCpCYG43Q+aoT+IFPxpM3JzJLEJMVhpBE6V
sP6ODrtV/I5mQ8gkVfLIvh3U1oqhBiUzcgta6gHQYSznSlEEC9YmltaklJFg2IsA
Ty/K9dOeWaE8UmKOVROaaxNq5V4Dn3AXw7hJsT+jQ9r/OotyrExtGZLaHoUZhTdG
FrPX1rNWof49nDXJIcia/SwefOCbkf/yN2IiuKJsX20DsJcTwCH1z4FM5Oj2IZuO
YEROlUOZacxmfgCztPvWtl+AsPZME9LXFXIP9OWmRy6CXx893+kGTVfz6Td/C97N
IUZxZqHPJGI4imN/nRh+0BuZkcIZZ5/Vb1k8Kyk8JAMqjaoDsq0O3ONK6QtLNqax
8NM22Bq/fiuP3YZdw73+eiO38JJsHoJXjIFub42rWVAWg1CdFUdtJfZ3wgf7MtRk
/ALT9226hAjTtrbB+Y7uDLME5vJzjlCylp+rjX1hgYw+6zbI3hJwSC9Hr187NZiL
g1Xzc61FHgZjNWxVLEwgMjhK7iWR85xyb0W6N8AGnU6p0jbFwMutRhzMlKzL/wvh
w8Cy3zJLWKIoVAuNfuxOjeapKsCOvSB9cj8WMkbQ44GZOCFctEyrwFr7/j0frDnv
lvkhJlbfX5aM8R6fu7qit9xbtaz0yoC7sWtABfwK5O+18Z5CsDg96gds5IbSxcoE
YS46CqFxHDxq9gL4tlIiMoqu4IEbjww6VrTTQcAQ4TpVMm9V9m25uybykSbOjieN
TR3ki/RDkOpqYfsfcTd/JmDVxWBHGSmed/1RCLg8ZwsfN3ekCDqgxXv1cXrjPB1+
NQD4zHC3GCT2DAqFUN3rVYaO7PZ8krC1eIUpsiY1U6YOFaq2CMYykLmtKh0YcVJp
hmAtiZKbelunGqNqJgXKKgyW7PMWWkKaxABC+fqI234RpMIiWHtUylal8Zyr+Lmg
RiwlKY9OT8smvBrPvRwDEhdktzzDLFtusGuvPMT+SqpRqTA7WYsHjQhzZAFQNGZD
hv+Nr6EkLsoq/XKYZLieOs8Qe1mp1E85GYVH7eaggyYgKsua/BFRYFRdX8Ftnqa1
36bbwCpezF4mnmba6fpUsmVqeDqFGUxBK54PKmXt16tZDwmLrJ4UrgTTHCzXEcIP
EVn+RJALEtDYUioWmG/85uqd5ZSwtz/lheYWhQUh73q11s9DeH9LTK6VKWRNOWNp
CFk1gA0wCvcjnCqGV4yXDxx2+37rlsm/ZMI9t5EwaStALskl8hvPLlT+q7iR1L5c
e8YF95LoKyyUwfF6RcIcxbfgJ+uEnSttpoZvqajs8i9hP3AjSUVPkvnTB7+hvcHi
3mT4oyhIWbJyG6+L4jX6YckawfvWExibUw5yWTT8ur/x9NY+4qIdAJGKaItKbyKQ
vRnIr/WH3+M6yHYBnq8P22kJv/ECwBlD59gbPZPGvbYtg/ge3qofdbR2X9+M5W2O
LdR22dnSZGtiaeW+2KpVyuMKfXeVIbT5ycdsFCsejVv4gOO2yaXQR2YQvoXKwvEF
KCoPHjod0Vw0SBP1+HU/3zJEcRRbNZcjdqsO0IWSjTXE2zCHM9Pz2fVtHB6UouPy
g44438s59dscLIlkAY5juCCn4EH13O74R49ezTYumEFtMM4PQmpMGuQfjZPRExQz
CZJLbTNxZ3sMctMYf4YWbzTaiyOpWQmOcQvRbgRQbOYnq9IvCNtTXcZVg6pwUgyX
6EegTXs+eHdYk/a7rejxXvPQb8pkRyhbvsU1QnDpnrkEbw8Tn7JaP6iIx9eehMOG
wATTa2oX95SruBxv0Bb3uYzJO+4IAAcnrZjnNSGpS4KQORncivwouGAMfKrOmG7j
mV/VIv35iRPStXjUyGhYMTqDeuob1yiBVDmDYbFrODDrUgnRZTPC6MQOgRyTA5IJ
9TmswjXY86K0qv4+w0m/knWxmoBuVlLoXSBVLGSBLrVVoZLv/N60qhW4w7Y76m8q
kYT6LKjUBgAyhZcvaC3PhKO+jdVvqAGnAwQwv0snUop7cNaRy38QbPijKGYutLjH
HDP2yYjTeY1fh67ncJiSXVti9p8bRJF03OHAcCGjmLQODZoOAxduAJiYFxAPY4tb
RnBifLfkDppU2xsYDD5nW9/8jWFXpp296C2L+fRGwvz0r61qGoKonteEk3R3NCwq
3RG+v1ckg8CYRo291C+hDS6knYWNpG68m/S4Lf3WysYR8gSnbz+R7E9S5SkWEIeN
1yn9MTU3Vm3E7R0hHTI0981pONiXJzN9qKJYCrwadzBBIqC08xG3MJaql2wiLfw/
sRqoHKS2aYTNE21KIviseJmmpmWOodgamgNaqTKHXrRnhMfKPWX5HMye+50VHEvE
ryt05Klxea3vUXYGih2kbCRQMwRyRpQbRm5VsPurRedK8OvI5OIwdnF+lgcYeVSN
/9Iv/X+fT7sp+bWMORviHnASJYF6apRefVKEneEshWZliWOA6O2DHtONIhjcsSwK
BH8r2YUXmzW0Tq0J9vXdRXfPklE2ylDBHBeBmN18/UPZ8nwNPpqMJN3wYmSVY9/r
mCjFh6zaV3KoAEAZo6cQX5LGeJSSctFapBBY/+uKRQlekafx2Pl7YGxQvVRmy6wW
4IPYSowy65ntQjZnO66M7sg5yWa18dEfvqNEoO60jbzDmRi79MlLQsOE8o5vAaVX
CV0HPtnHU+SrNp/83wLEfdt+B+nyC/qKaFHH25VZNXAPmYYLlaDL95c6DIuCOxFm
sdAGjdgJl2ma5jLTJsGVRHy6d2kzUjB/NyWfHBr5ZzfA68ZdWjIx7bZomw797eE3
vHJGza1rP3BjBzkgwgQKr7/0xoyiTecLMrQY+184cWD4+ojn3ECaytXKtU0qEaJz
nq+zoSuCWSOlQeSth3vHcOof8Hb+mi6zGmeMZ23t4PflIaUSGKFSx98MJfqpHp+W
zrOkIM0vcq7e4DMdXZOjRNcMCTWtDzfoO2jZRu2tvD9ZZ8s633sZHYlQMOLn1ZaF
Ot9eFjC0JMmn65QOY7HWgqqzq+gYqsZqJlJOP9yDq9bRrDvAcVMOijMV3ju9wj4o
l97FY8GKlOeQSjVA5Y35w9qgmxvjFLetfQaJDZKH55XnnHPmGo3EgcobDYLk7t28
oYLmS6Bb9J6u49fyn4allR4rzEmJcMXyQkyCqHujz7JcUuyPVIOnYX7Ek2VwexuQ
95CxZaror/287l0QSgiHOlnKxpktM03nWw98Ii+J5wvH5cBvtts9QcSWek4jIwXr
j6qTM/XB4XFMh5MOqJNHtuxlkTIY08PAhqs+RU41YyLjVvAXTSCAnHPzIVwV+vYa
75NB8kJ2luwS/6Hr+n3B7T2PNKBLgtZKB9VTc5RfB8P0sNZXDc/C7WSwPDzDzO86
raIfGf8tb8ohKqBLVIue2RE4IjIBsFAjjlrocWgjnWQzKQZSlchp9H+7ntaRkihz
NN06xwsRnnfJHfNC9VttcQk3hZbRzI20GFlfHU6RjGQrQCvFQTeG7gE9eT/N3Cm9
1Yn0N/+be1WSXot6j/SCYjZUzOgnXifWyiLvBNOGoMlFQruCbAJgvBtcFLQ+rOHY
lJAy5Ey9bSjRNlsOfhb6IPb0GASNid/U6cVkJYOWrUiNjKgLJM4FYEFoM4ixRNzu
YE5dogAzL2lRV/qcFEet8UEbvTi0H7CfMNmR3xOnbybH6CWIS+79vHEchsgq4ctB
QLkQkHAbAPDmoQvG0XlZNHLe1Bzckuu1K7od4yP+8o7pKnAnD3Ov6vxK6ZtIDFOq
52adFs9rsTW/WKj7ih1wpBvnmuW0VrYAZysQSY64eFz/S+y3UsTWlESS+IiS1QmQ
SqI9AHdZWDiAZolE+4YLRAdbSkd6ND5w02K/9Oa2lbq+8owsWez4WikvM+xBQvW9
Xp7FRTN6kab1SRqlU5+UAlAERObxVW9Nkr/UVlmBLDSFmFyOqz7o5fjiYZF/yEkL
iaPGu/3wFGr4iKo2sp6LlVeCSrDPUgoRC5eyaVMQPqw6i23lkxagiEbeORFveYHJ
+Qrr1gOEFfuAVnHRJMrTh8JBeAHqPJT6v5kr+HOTkICGSdKiuKjKlhU21e54INja
ouJOQnplv+DN8qqAx6MjAsY90440nbcpOGgB6eisWZdRhrvj2bimq3PjkX0KQnXU
BeF4Db/tuuYCiLo4XjMLw9TV3wsFwULyj4lhSl4Otv12VW4DmC+1vlZ+2eGKwVng
VsL3WMg9qzyYzNPmqbl7a9laAfFs/u8PtgftT9Au+/Ea/edyM/YXsZ+1WF4fPVsD
KXKNyuBXyQwXxxDfoB+qVVw9IzqoR4J7MGEMLXx9ziQUB9F4liW8e5AXDVAWdegl
Mu6jw7DO7rC2RMn/ZLtn+VyApbI2c5SiOe9R2A/1AKfaigy8yMRst1XZKYk5jVaR
3Po89LVhA0ZPbwGzLiHCG3sJEi2B9JNEk6yun5gmcRmpYIUJVtoNYr8t/7ysiskB
gHbxf0pmUVQSOE+QZ/Y2kkSAC5AzPivvXvoBkBe1JmXOxcOAvHpRI5DzLcA1S3KC
dp5+o3nGhDpun7kT5qvJyDg7bww365L6gObbZEgK09GR+PyiwgkRdWWgi+jVQE6h
qYCwjQGWk1BlwH5frRy24GodDdnnveSfzbA/s5b2rbLXAlNYCi2Z4VsU6d+CeAo3
9aO3C/nGaWhvUCZGoHC5kdk84S00XPZaCf2JQ7Aje2kEoqTG1M7VLvZsSq0wJ+Kc
tSSwOyN98sCbpTnARk501BDLbVLH3G9CzWLw+v71QKBKz3TalAsmuNZ3yZFcUYAg
v7ZLbJD3C/PXDbHWAV510RIHU3/WKKuxHM9l6god6wgXZrcSCAJhfZyOmEc2lA0F
sLHYNVTRjVofAGQbdo4oSHB1NxhxKkiyCpg1Eq3n9N6I1tHvIObShi4VsHDyuPI5
BPR/SCCc+CNC1YiVB4gC8OzXhtbAXdtIJHwaA8j0vLcLuHy2rRJYZk2ewfZlpKsa
su0G1BbvpxIRNDud9WPF8cjXwZfi1V9YgRD0KCixlZnObCis7p2rKnN5/y89+BOl
JxlNFrJDLmFZwDFPdqPA80TS7WqjPPOWS0QvmaqBl0oGI8+4DAmVgqJj32J+jRy9
6UtRpd/98RRfC4t1lxdbU0i9+hgHPYFcQtfYZwterQlNKD/lCnsR4tvUCuREtgR/
zpuOXkyNythcrh5MxxDCA74vL0fwn0N48fFehUbxZlLd62QOAWl+u36LCJoRhjjF
jEu8ebZwx7O/OexU8I0Uk6pcTY3QkSyAYFtIuyWck0PvqcJuLEiIT2MzCikX0JJI
a1Mr9FduJ2jyW9zeM7PwYhrB+uvIrQ4cTd3GkDL0XPW0y7g7PllNmixc+zZDIv0R
wGHJrvmcTchZKME2SphLntCNNJ5QMnsm8ErowfigwHQTLskziFg+j2yTJrS2TtD/
7pbkoB9xycLzl/2GoiP9ZdSfoEJIyjmLKnsVmq8J9SKz7yX9v0yM6wiM5T5taQmv
/rg1guMsXD7SMXv3skoCO+fFt6nP6JAwdiwUFe5PnpY6JPPNw/+XeZ3jo2qckYcG
o203rdPjxfALR4pA3ifBL/nPuBwsoP03Nfoqv1MLXF8rHrwWyAjx0bUc69UyqSQr
16Vg5m8GJiMIJzhKyNUBHRkQNGVW9xz6EcfLw+I1LGYznkS29x9zBqRGUZVkkZaf
D8illWYh4+2XXUsOXtjPdGV06gIs9+mbYVQ2b2rwLuRjLi66hh8cUXeiBjcZAVkt
nhfq/36lu1ehjGSuxFljfrFKJECafU/ftMp1xj8YuhS3yglM2QhG4EQ7BPLKzmpT
ZQaTILuP4TlQNrpy5Si7tvQfQ8f/RsiLtvfgiCDHewyEVwcDliTVxkI2rx5C9mXU
CjOTIEaxhXqeX8Bnb6K0X7CFbHCLINzUQvXxV6d/EqHTGyZO5iDKy47yO8rhbtEV
CCr/l1cRlyj12ft5vjziUt7nvNt63X9LVMtZbG/qzfIW5MBW7b/jh7U9YOjammAP
tKvlTb5yviNqa6HCkWF3ZB14Jwxlb1VEZglO/u8lXmYEm6dxwVlp9tjNPXCOlcRY
SQsyZHYqmqAlD21hoKUPWftekEpclrwCG8wWIliFG4fQFZem1sZBbnHyu+ttui/D
jOc4nSU+uHzzBFZGU26lS25rxYsIViKKBjTevl/G5vc2Vw1/wcZtG3sEFFH/sdXJ
0fvnFdGRzvv2bqTQGa0is23Ik4XkWceAycvJwdGCW+EZ4PRs6M/AbzPwL7dIXUWe
rJy4IjiaaZFas5J/wljyJ0fPQZrobKyWorUYMiq2eSF+lkN5YUZk2KLDuV6nMogK
MOeT3Oh/DM+ojVOu55QCr0MwTTcMiI9nx9IUo6RogIZTaFUMH6brPT3TmCNdfbvV
/+wXJ5pCBnsDG30VcBbEkpehwvHB2Lm/zgS8m/u9ppjLUNLZxnkgGG5U3am43n0X
qEag6BFaUkei5VMr/LZiQowTrUH5Og5VhM6gfT8B0S5yGQ8KFP7rbjfjcfkHAAE4
CAGKJbUrqjHskpEC1yEXEuLuKtgzDWxnM65CHVbMYtSoZ5nZETP1vPtMO3El5BzF
HFW8e8z+B/zYqrckd2wTFoxgkF8ldp+eDZDeuQSkofMVvImfnBB//NnXDFtWo4sR
rdVKPwUJQQFQKarhrYDOi3GDwv6Ppk+FUik0DLd2jZPY1V4aSEKawwYF20FZca0/
7MSuwkI4Lnpoj0MwpEdsLIFIsIBuz0nNmyByjUKIz5jNfC/vA5tSWsIprnJW0cpv
kgZqTlEStivHwpLXh9OaD4jq4P8IAp0m94eSDj+6SBPdWYBlFoUTIENttjGod/xe
fNYHzMEtFXbu+6OvkL1zOwFP7RQXwfw9cOzqlSSSutF2qVSihwxbriKZF0pLLh/5
WcmQiHcT5qAtKrF7OhmeJYuhNan8X/T5uDmzkuq1MsdfOucqQug7cGOTuywADcLz
OrF59vxB7dU4FLHtKqWsRRC1tdyI2j3VZeOCia89p0wVZyzXpSBSxSXo8irXYxqr
unSkXwEpeN+FaKbEGPF3VJN0y36cqxB/09IhuKEC5yR4F/PxRkAPl+rSvIhiMBFh
ZU7e/AeiVGCQKSSbueKWUD75agSaGK/ih2V78W5Z+83jkSsyGWIzcPQvf1KZOzoC
ozkuL7k+5uAn8o0DiMpuFTVmbxT0EpaBCM5QY0xaqjLKYYyrpDBGgSlegcW3zzKx
5BVk5xkE4UBR8MXOtBHzbDBJCYo1CFiPlH4yZ5lFox5iiZPBl/Hv9SSVfgTyg4GF
/BEyFmFK6Ral3f/5fVWYJ5PnA1SBEMpx3ML41uTg6X8aXfftoHfDtZ0mQXw1VLWV
0NMRoTI3fJ83ebQDnjSfWZ2d/Gk/OYi9JO795maXaBlM5e2Qra6dplu7x11T/TZu
GhpgJO4pQ7U2IdquePdzhM3VZhQEAQJdnMOvoLmI3xfCPEAIXhd+3Irf2qMWOVYJ
z7Evyn0ywxysDx7IanskIBkDbd7ljNDUr1oVPikDnTSiJ/4fZyfo0ptn/1XLtaf5
sf9Ehw6L4fEFg5SjeuOG5Ts5Vi8PGJbe67CUX1ci5gybtrv2wnFhH01isrbgFL+C
DGm03i9O5ynS9QofR/eQcjc/U5zmg4O1r5QO95U1kk0c+nHTfBr/+q1KQtIN/Fsn
9E4LiOM9txhP8LJmtds2qrsOc4jI2aeK8hpWOqaaO/MZLOBGBGsYH0kzQo/Ka3tC
mByhAqLzlaVfzwZ9x4muFQ0hKf64b9mdLXXANtj9FpO3k0xr9+zAF6n+O23Rfbnv
RaeAWqwKMKaI7ZtX507fImt+TipkvpVq8Vl+geKZyca1bu+UuHBOT9Gd4hlF61mN
1FXdZ6ZCrf4QbCOdYRbiLIx8hPmmSLR1TDQ2qKe/6q+lqJliTSHZ3fnFrkK5l9Ww
WFf3+ptbxSt3PFd5ckPQBJN7H5sxb5B16lon0ALsFHNRa6YM+VwpzJoKzoIapSZD
lBBbRG7KYxJm7brmvMF6DP3Fq2cdAbU7QEq3zNZ/B6xp06EccbtGGn2IwkijRHkx
UVDHS4ECzJtMokiYSBzJ3FawhmYded+LBwVHwl+xNKt+YTxDuVDIWN95oXMAM5zS
+yPNVw0ZQRtVGacf0DkVHSVaHEgS3nspThdn0XIfG/ok5ercK0ttii673W92XgXa
fTqwJk9Rlrz+9wDqicN9eg3ddxn4qMnMzOcbTOQFJxrYiIBLfZbKT+foD0fb94Fo
y8YDpF+WIMOzvqD7Uxb2usuWeNl1s581+TNv6hED1IoUNW4d+N3nMu14ne90w48f
eJfWpu/8EpTsOs44JCD5kA5t/ZcbqVhrhkSSoKEzTauTCouBnXv3hxh70acwKei9
EZUpHbpjyuAALfSS4ds2Hk+tJhfh1JgmTA/pkBZpr4xPGF8U0L9kp9ZSxN6KA+0y
6IIH7+luvcTxapwEzwnoQ9T7pqPthJpoboxQKTd1JdqDqtQ/wp1FzFK+mh0+I3Mi
/gJRbbmQK/ZstwXybXJvs/Hy3J/M7ZcVrVcP5K3beEA1sAiD8ynq5HNyMO/BLwpj
egPb2ulIlX6ipG5mug8W36UfvN6m2eoU2Y9LI5hZWzwTqfRR+3ZEtcLA+ed6cgPq
Siy9ov8n0twTzzb8Q0ngfyj1mH3GwzofOkWqoy94X6mA7A7Jev4Su6ifVK5Vsa1G
cp/KYRvBnE7o06UVax8V2boQoE4cGrEpVsiX7cfe6IBFQZyq+dacFx1cAS8MGjXO
975nC78fRpsoAS+/uCVHdJB8W4KmOVzbbVmRYs0ZOnUMEMfkp6NN9CgNHJzXkw/Y
SNSAP6XPe3NvA0CJe3T7nqO/kvR33ZTv8NWpbVCsnb0d7uVVRaViND/bZkaRbLfC
Fcnne0uUJ30fCPt24yjg0/VCweMkjlaDBg0ce4SaQP3LZJyhV7tLFmPqfvP+dGs9
M650bAyFYw25hqH1BET4goz9nOkmrxVRqCvjdAwiKdhg2rIHLvHVauP3vkB3RPY0
rSwcK2VER2rNhbQUrjUbIivLt5GpyXk2Io+1DZ75Yf7ByJVf0Uml4Nt4p9N6GfdI
t4aEHKvK2ShJwf5wKNrJN9YvXiiSk7XOO/gSePvo6GXtruzQHB4cITbZjCcBVhTa
PEEnlCMB2QoYNRgyphhTiFVrGyTjDiAP07MGEHKIetgszRBpa0XSgSwK2AgqZFyI
1J/MYyJRyeKrl4z9jye9E54P8sXYyuyfTof+R5/z41RsUssa17gSnCZ+fpRKgIh/
aV649xKghAheWrkJQQFo+hjpHMib5hqFe70Tp1RQpqB8dR8ihBZym1/F02kMhyqW
ql9e7v2xcEGv8RxhkUYEu4x9wl0uRqsWbUSfmFO+J2ycweyAlci+GtPNq8nHrGxO
rPmjow6KF7oywNDquSIU4wGamwxtOBbRoy9LMULY83aKWwgzxLb/u5/oSdqAXJPU
HTBjF9ls//+rKYr7uIKq8fY9R/mVn7uwlfOWNZNa2xL0kuVq/3/b89hpfTF18x5N
whiX2iTGom1ZB1XjTSuhzGXpabZOu9N8/AjXFoSjTtgpJOQbEpwX6jgcP8KELkCC
pXEygYCmwxVLtMF/NfppcsoTY6F/4N7oAEI3ckCqNixgPAVFlXp0qQsBZHAFFUsf
Mzp2ZPQdt0xL25EfYSitiALoydHO+AeRL3UoZDksFfvuTgL50BQuASmf5hlWCriB
HXot6QF44+onMmInGwqnvGhBKy2jgfg60GqUN3w6y3rXDcw0q/ureG9/tE0P7fLR
ya3MMwdmjgD99auj6QaLT26d023zFu+M2zXYaujKHJhxeKOjpIzkyO3XCeDi28ny
CHmSH1ZZzpzy6CsthcD/t52e0UDDvKgQ6+JLwpmT6nSi5IOe1DyPh7ZdfdDTBYuv
Sus2iePYPlIzW9s3fIn/kL97hVLm38XTbYQYBejoGpvE4FXfEvQniZL6E8ptmSRq
g8kQgiWEOIIN+M6RpXmpuIxUMsnWSaZKR7HV4QXkeb/UnUValLB9BtdSImCcs5oo
zJKl7qc0Lsk1QVgmbeMJbDyOzj/A/fF5qtk+mh8vb5WuSH+6Tc3rtntcesNevnoX
UOXLBlVjvHmG0B5u4cXGoompGUHeEf5ckCvlf042AXvCwLedgNgDo9w+VZwJu2p6
Fp0MPIrwJegKYKCYHLFz5T1mnJM12RTvAYlZDMO+vM2hBRjVuxj+AVP852iU0qPI
csWHQSIjJWidqiophbffCBRjwy09vYbawgqj4JykBQuMr/Be5gZmtk505nG5D59X
70byFUmmMs6lSyjfabsmEEeMn7OETiGL5GJpPok74jsgpMA52E6Ib7I1RjJ33QvN
EgvEar8D9MpOCMJZjoLPVG6nKJC3+neOLnxHcgl8MZlzjiWAXtLxHkjbm52IxAn8
Nzr4xyP5JlZ6hS1ZfQ7PJInlJMKg3VdsliWgRUZqJPAsqo30Fo7oj01GcIRPhvOT
Sn4tAqruitulISmEWfTfDqyfWUcutMFLIfRbyxqoUuH2bE7AjVOQoCtO+/5BS2rx
hTqYz8l2gE46I04RE+4Reak2WRM3y9RjSF6jfT22C98/5i+zEZ99DpZTRHd7aF/t
WTcZdXtwnnNXH3/NT6OLwcbvv+AjPk1qPRZ2An8HWmiRAcfIU5KtU9SasPee1Wir
i6qNHj2rlxfP75HiWaSbdxhxUdNo8v+iZzIK4m7Rp/CZDJF6+ImL9vjG7cY8K2Rd
t47Zd/GlqZlRvimcdWGujLVF/BK0peZTYyRb5fc5Pnt75Qhea51HLM2Iv9jMN8LK
xaN55hMmj/ZtGnJ9bKDMJfd8sPRM1wSWKDf3vqiQUFAp0/B+yMsV/xM4B0HHgQfI
jqJ9LF4/jCxzOgYp5Htt9vZAUwVuiaDHJyY0I7ystcRpkjwwopEhYZPJ9fdL662K
j6RNwseyfKYaYruDAAYkkS5A/u9fFryUPLsqU1ZsFHSUJI8AZXfdGFASLKikB6ka
u7E9WZipS7DXGIag0SIiod2j5vlxpikq142FFzRcOYLcWFIsGowCa2XR0dZ2etpi
nDIuQ72B/DrMb/tsEJ6dhmb6xuUvZyU4BR/DaOkIkAqFr/kzdRqYpf1eKhpqG9iM
QjzCTCsipB9ScbUoEsbx/w+QiKjowAdwga95FCu2mwISnd1eRwIi1ART8Psz+oFT
/UwbuNU9uk69GpeHzv/PDufIp4yMH5sYKeGmzGbJPv8CXggpMYiXOI2BYKfxvYtP
oZa90ng88R/ZvLZQ3wG9vRfKWBEFRweXcLUfO2Zs9EVU1WSfOm2HcD+Yy9QqFwnM
8tUIcvBA8lOX/jo/45b7EFh/2GAmlHD2bfJlTY702WGLQvcho6W9dt1QX3TVYkO0
YiTL8G7bTjH0w2BZu5Pa/FRltDywMYHXCM28ieXaBMlsTuGsAle5GQ0y2xSgYNFY
Lga6qvEWRRd48NxNmGD0jMd/nkXjqlUppa3fPyc7VU0gVJKjwW0d/tjWwxTadO1v
ABx4jpEJo9mv7QW7z5wT3NQPW4hnV4p8FZ37XOJyT80Hz7gw7EHmM5krYVSnve5Q
LuOw3y0BqJpkBt674S9LA1ZLjUiCBgSyOBQCj9omerolxSzRHmuLAQ/NQmAaRJ0Q
1ExFX0EwvwJwTSfsyYsv1jQ7r7Dw8zXC3ffljiMt9sEVxtZP4Fh9j/yq7ErAuitK
Aob3Ro9aUIcbQdG+IlslVLeq2hOyPZJ/XaPJcVDrvlanFYfhUFn2OOXDOJhK8vw7
4bBnUyVeXLjcJ3BvI1SMWeRak+ppFkT6gSBqy0tLoGSwr2X2k5gfTTy7MHQWfvB2
Rw+QCYcHI4JDp76ztStSAXlXZCBXIoYoyhe+2p/nLlWf+XnI81HaZcjX3w/rGwHo
RCDgT82RqQtXYUxAl+EDJyz00B/aWApuNwGOQcF9uw1zpp2juXU7jag2ZPXBF7kl
NUPXXPINvqkoHN7gUCR/eXIkFUsm+Id+3HxB8YM4RaqekKRr+hdICgkPxUsgfCd2
Fv5cfQB+grQsVRa21C61oSFp/CG6zeS8eQg75VPliDSsDoR5AjFLV2noUD+uJbgo
5pyg1++ZM6LIZxCdXYVTWppSmYodHBArdyStY3TPrHo74UrnQWMslgmXr2LIpsU4
aqDC1S7XlKz5chvBLauR/AKLZENiSPE2+aJVmTi4Lhc4gtybNzFfQsKl5cQP9xB4
e+u/GnA7gQ82SQNAGVY7bsyZgtfH9Rcv+xxpqYMbLseMZDzL+looHCN3Inq1hcnp
7LIySXTtx3YID8eKt0BNt01tLojqlJEttTMFMpJPsPSNS3dYAnr9XqV8EaOMy9mE
/NxFkVKz2+QSsJHH4Ysv2PKH6NhU33CZ6DSMk5DEJcH3wHONlMYstqKwKD1YFXXb
p2lV/GTBS9O7qHYuuRDn9oA0Bj77N+sknzwvedrzXKrRVLpVzPHk1eatWnHdzIVx
9DsgyWJxptzMHr+Z0JagsPKYJz2PjeNZlQQHq184L9HvHUrJu0AFC/ItMq4fjrEE
UUrndhyCOkFkVxmWUaEKfcSuNeuUQth8EBtYzi+wx3LFO0ZaLTfLgO5llWX1mvZy
/8NcMfabptMY2yTk6uI4ISAdCLd0XTbgIo+AX4wCgnHxEqciXB77tvpSp9E3LT+e
WBoI0fP3/zDc79jCoLfZy8mpf5/AYkzMM/Gqwl7JW4fwvtzbWl5/JJal/EoiEvxK
36uRfYGkvXn8d7AuVIPSdQdARI6MEiW0SMy/WeJzYoeVmwQv7UWE4sYHwM9NhWcV
nZCQKgR4pchmYpG4zmDYc+zxdNaXcsEosvewPS8KF5VqBA7CEZsjTPB+TsoHQeCe
idCfoTSBt198PH4mOsgNIGBebmFpGWDY2gkcKL40yYTn3FoUE4AuSvByzXVlKjFP
6lujnkoUzmmBIN75KCR3yxiZ1vr2RinPsA4AGGWZqPf3dgHBRGRJpQXC3IC87LR3
DzeeAJidFyJyVQHZYBxK9sYRVQ1WKEY5G4m1SG/eoqukRHJJpn3QXWlCuzpR9IbP
odygLlSQ1J1PbdjlrWNjSOgyBF6PjkYK6ePNyNPI9kj1QkI10IueOqEFbJqVt9I0
q8B/g1aFC+rEKglkX2GSqL7PacYSj4zgkamcp55jE6umPmibKUSMQFVkNouNgeYq
qOZminqc1pk3AwrK1HCAB5KRcLmVsBOGfoWNAQf8CR7utDkkALgqQjqZhrhJ3nsg
Bjyf5+aeEb8ZWIt4I0p0WLBWmp4RgMExCdl56dfRfx5U79V9dFWamrUQ/usd3yoY
BZ4UzjLmwGrjzdqoF4Rgt3dDqzjSoQHdznzEqKzAVF6qbctiHYzprrw3a/58//67
6aVyRXepkGfWBm7dPdoEmbJ2N8kyMxIzv1BKvjWbcdQpac7rUljflE4GTKWE4KGl
GMSj6w96tOfOfhOb0sa4NajOjzxWIJ6YpWKe8kyjuFyZ/2ZQ9hUi/cKXCcWQp8qj
Cnhq/OSXxDCap+gGYZ1WpumlMcNSO477Z/hT93nyv+FsvzVzL+JEfHXR1+6AFaH7
7Jout/qpochjxzUXYaMSBKLP+8kh54pBHfRb8pgp8tkPtLxF1j2mU5VhpQEngKkV
b8jZ2ZZ9RIhD0E6OO06iTh/meUC9aX0qtQogZZuj02f05d+etvEpoB+rIzkfjXDx
/MuJW2okrPZkVvAzWQZ57MMis3jJ+P9JIocsKftin+uq1LuxprOLrSpfZnKZQJZ/
uDg52V7JQ2y3tqWSt6M1EinCHhRxBWX6O7fwxwiYyXl73COSjptPWkOvrBG3fpVn
T9ZszeZ4/SjQS82l0gDWyf436I7vKKbHVlPzlSyilwug3uqm+/yfjuFKhxIQ+OqR
71xZ7PCJ4vT5b+D4cQqSfjyv8jG7qAW2EFoAZkH+uwUqHmZ2KlYvsjpP9Y2Skc72
16hLHRbI3b8K+q9yAll6Xi+9QbcYm+ljYr1qeTk86pMw2XR2EcgRbe1py3NfItVz
D7rmqfNG72hKSLMzxkHgX77Yxds62U0lsw2uQvk9p3DYI49VX9fsLD4NZNI+C2c8
7Molmx3bWEUoXc2JtUco98PQGr681d/GFUQHVEopZgwBPBcf0yQnsdMYVOGjlyJI
7AJRIkeEP5ztFoEeCMfkmua3iA523PbCUKj6JCrNlmIiG0c3pLXxLr2APRMYPygm
qo84KBGPlQzZBpBTVUIEfv/Rqzf92pIzH4z5yL4Ft5FF9vsdfinOJ2f5lFWHpml1
eK6QqrEWKkI+dLFJ/3kpGtT4+XS04M4EE9VB9Wkhxeaw2mWt7rbfvEJ+M7pERH4W
dkASqK8GKvWSqUO0OS++6mgR8AO94bkbqadB81gw+DvrPZBRhRxhLB/r1/Nb2h8E
A5h5ODc477Sp9Nnr3Jnm1su2iXaRdaJnB+m3BXKM66+fDggaGOGjRhBkPyjK1doV
CI7Smaw9FgljzpVKlfa/pSSTferhvExlzPGWW70bFnOu9+feVaA3wuKyzMZKv0/4
CDKHXuozJRTug6p/X7eCAXKFfMHeqrL40b6+HiA+89ShB/fweqvwMXCs5vJnCS+x
j2HOufQEL3/7MpHdRh4AEEeKMSPp85MSLdWJjfePcl3KZbM9lhU9SpHHbhosPrk9
x/tQyLoczuN2eFDcrnVk6Ek+TX6+Uqldd5TbXntMogYtnFdmzn+NNR7+Ylc63Bif
iM/zLyqgfxHxmyGoPf1ye/6tfmMIamlUm1avrTkWRVPEPIOmoJH8jbDSb+wzoy/B
zehS6+j5U+Fac3K3Z8LTn3rWcsfR8sQuqApZKT9avKHCpKUCtv0woXcOgzc/D4Ps
macnjaPAARAKtxoP77BZxq+I9XyPin/ufraoxCKQOLgqugz6XOmVMYqVyF4q0z3K
5X0XAY0awGfYq5ofDhCI+iOG2iRn8iD89/X/6Xact7GS8EbEr4omQS2WWcIZBTeL
KAgfdgWRX359git1/k6XhtbaO7czOxMzZn4Jsqd5WgTzqhuUaf1zo21ujHzc6nqi
eSrEQj2dwexUutKYQ6nUYShNpByRqd2Hvqm4Zxao3DcszvNQ4q09QcfltIVlFEDc
mfo7+2pRKt5qbwLFk4yfpHDAHrHNb2c/pyp0STvFQPMSD0E2f3wcPkkcF4UZuDGR
uVOQtuqctgx6Z0sg8gMgfIkiO6yrDZVLZNR3U2ci9t7fEPc0c15E2LXu6KOAscQO
hOuBvCHy80KUBxlmAHgBYS/L3gpPjPPgqBPl5qVu5LLVg/Wz27YpdI26266A8M36
+IHZVPNx3iIqIF+Xj32LJl2pCo23fEq/7uMs//n+0LnL693KlCyq+ChxRvkNYTkU
7UIqAD3xJ0s8mwZRsUceSOorm7wXuklo6Qb+2ZTWgsnD3ZVqbIBGpXHlTYzLI0Yf
dBsBrotP2EiFzmRUcznO+mbMnjA9FD3OGnXL9eWFC55//vZ5nO2l/9bHG9qRvqOm
cGTZxBMn4nmQ5vm8q7VV6NumHbBScF6mqH25ryPm/vwSMdY4NhJ5RI8QddvuqEiz
i+G11YSdLP3ToipZUMPrw4ema+uthOkhgE/M+qCsgBazkEwTrlt9Y91e+efV0M5u
y9LHEje3Q0AoXDYhAIpkUHnJuuDEdQtXBGzoJXTN27AWhlyqwS2CLZc6hhxVoOvz
XFrpfQxzhsAHwCabEn6e6TOOdnk1lk7NIbaPOI2ht2PoJSUrLK+uraX3aFq76CLT
U3rWSGIOJBiV/ACkEpN+3VWtxjRZm2E++fx5pMuPOlPWWNmc56UrA+n2EZVQZJC8
JSH2oJIUlFea3NMR+kuPbT+AsEGYF/PcLPoPknfWR+owLOVWnW+drNx2zIk7zdBM
F96LqktHz4iTdxAq+L1H5+FnY8bOpb5Yo1s9HcIDd3t0CVuIR3z66lU8j+Yws096
0ClplrNfzhBM5GcU3iGPBGRl306BdeqhK8c0VgzHH2FNwQP8S+LS5AlbgVkagkCk
7G1ryIFMTPhk5keihX4oPfZEwxjaZALyqQJGmOR7pj/nO2ZiHKlCpF5Z6e/PjBvP
qvFPZhMC31J/7ONa1TF0Ns1dZESukOix7zZmDLAcny36Z3lW/MuFslKnhJR8DnUu
GlqvpBRXmDN6dfLFrbuuVeebrXiLvlLenLymTobG1CgZTLpSSqp/4tWygjwf9tEG
KX+GLlBxI3ZN90KuL1QcWODgOTrww38tPNuv4rBtCnvLMaeXgcE22A5gLFqGZrsl
EZ/Yr89rQ/39alY/w3eSj2+DD/8lFCl8RgjzX4fg7QpUB34qMeEsJoUgSatubyUo
+bKE38dabyGkF+qfDU+7SpqSnyjGKnXMmgxFw0hNpVfGa9KuEhEaALWp/GL1cy2Y
MPC747UYP6+aJ9B1MldvkihQdNogZCh6Kp1AXdTsxB1QWelXPo2yRhhZJwHMZicT
EVhmPPPsGb6EkYHw7P5C92k2WIqY40i5NiBENlUXsZyQUapGzlMB6J0odXXyv33t
W6qAshUVGb7Yh6wndXJUpmIgLoNQrUzIlEaNRm+pO5pTvcA9AmLDoIfbtDlo3bT6
a0x8XHmYd2H2bgh7IMkgW3QWGSnxjzHeZjGaN6xHx3gGY80v6bQ59PLT/zbCz5dP
lXDl5o8nOHqvntVh7Njg9W0zmWAf4sneEh8ckw6hpAW13Pc6kyWPe5HLeDvLBZQo
wjKKljeJT3URMNy25bhHl27M9JRvHkz/KdeUnnZEBxjXlWd9rW6hGaTBm0aastfq
L8L0Ao7lLfnOZYIFLZQojf1QK/vqtZwQUy+4ImH80DvZciDfjmSS1HeDsGKHYuQH
zkSGVi+uGi7nkhrs+no4lWmAy2hRu/UokdqiD4GQxTYtYP/8gNDEBouvxq5AQTPU
XfUABi3w2t39H4VlUQTsvsoeBrvzxjnm2G1KLUNEF+U6k10zlAlRLmcLkYzZZBFu
bPpkWMG4lMbkm+42WJttsBRqzNNIoU58vzS2MjuvBz07lIbn3S3UKAcK4mdeZuRo
lOsX8Qs5IjI4E2+ViI6UK+87AJwJKevbkVx1IYfSBd6xTkZoj7UY/5xL7na3StpQ
t4XpLlWYV4H66NUzNLhTARSatlW4h/iV9MllzWbmPuEFdfLif1qqm3yBvDW8rxTL
ZKp9amPzvvcKKD/qnNAJ8DEl6leIvI4yQSamrB08f2fMta2/Fl0R6Czy+UxGHjde
rvZlPLbN8mSDL0I6uylOY+J3MkiYlaW3IfZL5FQ6kI4eqVHIjqvOj7lPcR8xu8Zc
WzeLH4bztBqNqOz3xDYCHZjVVFVD81qoN5TKSIE9lp+2sheUA0fFoIaxlvLgEgS9
JZGbEaZPC24myvt1UmD+TtewyyyE82mSsgMlAR+zOkyu3e9U5x/UxfoSJBIjhcA3
Y3C2ljN+vIZEiILgouFZqr19dv43u+v0r8vCQ/Ji6OEv+JCNtvbd89cVub0DLKXp
0640tnx5ACZrhiQqB0pfhaAW6DcevLqE9YC8xMniNElRPi4FOd4QiluGaZDB1neQ
aFbPuKjWTScWJuiJBnh+xleLSK/mQeLw5GsGZYkSMBuaP2logxUQHtUlit8+o1N/
S9MOhDZiXW1jq3HZOLaKw6lnnEe4aIDCOoc2fEtitFxYnqkflLV69ymJLYszNTXs
dxLOFGYjhH7NgSx+OMdj6SYCppxinnmC/RawJ6YAdnim8xSiplImRHK/qQXGf4Pj
qCFx3DAaUkwH7UJpDx9R4OzPC9D8Nnk+M0bJ95V1/Q5BSdBiuc7AMaiyn+R7xRB2
wcuJ+9UsFXj2B+lZXiwkWNA+vLjhuh67Nf9bTbH+vsLqL3MQq/ZOksrWlyNRtDnl
HV8QB+F2qxCi2L8jc1QMln/jeLkYDXmipAw6uBToh63IvqR7ZijUKlq0Pp6BvZuZ
kq1cKaOLNguH6Lyva32hGWzfvdy71HTBNjdv5Bc4WXpQLT+xEkSVeHu/twJRoIPP
2e/GXChPr3SW7SS+PlXV9cAaM97oYKUUkldaLFuN0S3hIxRh4MUFw8AqGLThCsGk
nT5ihgJsX0FmPgNFp+O79IQ+o34Hqk5ST4f1P9CQUbsng9AFdezGaP3fh/3DHX6T
ZuqBTLuxjrcIISJ7+6DB0efxSEdJR+2smOJtD58h4rmHl3hpD6jzCOrdiX20lJF5
3oadilTVFii3EWqoSVtXSyZc5pBTzbrOI3dY3cZM2Yp8xs5yJc2YipqT2uIT3i11
CrI7P1lGFndPgDIgGPrK3OTNdWEPxQe6SewnEx6oc6btRndsfaJxOm45r7nS9jzn
JpT4zfJMw5j+ZmRtbXCoT+6M9Hx7/cmgAG8Arag2KP2DAXIcdzkY3Ohs1iI5oNLu
yPzoP9/UPAn20ZESfrRfDP7ze4jNyxhuxJMrdL/DDm9NMnZfdSVYRID/G4YzUlYU
2LnKNCUUdEckiyc8ODQyv4dCzvPrIjciH3ptquZIYmHjQ0PYXIJQUe4wHuQjTE2J
VLlGz9hNTAz/HXrZ7MoqgkSD8O5qw9iS8R5uadi/FzSMAaoqluhFuX2YGHprlIbH
NmKNxSZ5eAZjlwA7lpQoSn76b/KV7gbmlQR67EQmaW/7Kji5l9F1JJqmaBR2SZXl
55LfANgSD8fd986R0VyJPuwr+dMf/ZOLhE2xu0ACXy3KA5Up0DXbb+BND33kLhdy
qo6lX0Mqa0JwnRhj3XrPXrMNE1rIstxWih42zioH13lErS/bBGYbVVa/vCv21X7m
PTJETSwqtrJ98+C8toAwxhkAXiFCUrQfL2De+IBG2CHryA6lgDF1TvELsPfWqhIM
zZscO6ltMiZ+AU5eBt3FwS+eUn2aaGT3pizsa8Sdwah8/DAFtUVSoFdeeg+Hor/P
2QCdnJT5PhFI+KvSkb/xRBbk5fwlmF1KBue7KegfG9xrZqWOh7+cGAkQBJnPpHQ7
uKcHOeNQCR2MnG8SB87Scq8ev46HgFFXHK4unebFENKrF3izapQrUd+UNKcqzXCr
NxemKm6TlM+fk3aDZBnhM2K3mQXotIOLYONTduiZlQDeSHODP6c3OODBeTAy9r8W
r6YP0UkQQPBzy+25TjvNX6wpuB5F82KVjmNnoxR9TBCKk+KPaJZvr3x8JgQo4Zzd
XolOim2UOMXireSAZGz0Lyxufs5onU+TwJS2/oh7inWlysRZ4RexU3gTKHBrz3li
UsS5WtyHq+vTrfF74ako0F7VrgP6jc0Lre00OfH3Rx9gkuoYVgTbm5y5KLCnqy6O
zg4HYiobMykTHaOGTVV/QNjks9YLXxYL46CmIk2bfj1gu62c9AOVxRfU6ef4SVve
93NCDvgqwkot3WXwKfUd6V4C8pZSWpO2igo7AsLiCAVi9dAuULOLg1ennNuMJs0s
UVBgan7iApUJXP1oZgHgPpHjyDggFz0UeIducM/qF/mZQPe6V/Ye7rFxTHBeMupt
NE+9w2QimMcwxmuGFgukLuCLt+ZeXTr78ZiX2VkotrWOza6yQIm5+TEAaHleGxqm
PQ1lEeH1ksqvDEPaXlA71+65FDBS+BK91UUNdRCp1AmQJLxm2djJcbs3pm5/AcMF
KKonLo8OOn8ojoziyojo+mNOLTbLWseVvuWD/yQ10hbFsLENYfVVCgJV+xlG4vcw
+0VgbIBBLThy5PrqX7EUebF0gxWsePvi+zTm5YyX2CzvMf57IldfrYFcggCNZ50A
0zAgZ2WlEsSDJjYg7q4Eepzu+9eetqd6C1xCb6HKziihHZPYmNa++f6MLhr969r7
8R3qlGS45Yycl/LR6BjUOYwGsTPu382sSCNcGO69+WUGGwatGXg/0ohRP+XB3bew
FPmxrPsZ29P4x2N1SXm4rxFxWFvOdVQ7vHE9zU4b1SzNZGp51Gr/Ux9dzLT0kVp8
rJLZHG6yNsOvQoPyQU6g+ma9aPHVNIIieuwV3xZJocDo0SBNmss0QCV4xcHkK/nO
ifY/SJ77sf/FatNPJ7iWntHukjlBjnNn/mqhm4gJ6LWVJ7jyS3jbPbfWKz/wJTix
5ev/z/80uWjPqmqv+2hgT37EeirR43T0ursTsDUSDRN4UZh2uevCrrNkdZnhD7uy
yB7nNcW6ypDSP4KswN2bTSfgsn7n9+Aa2V0j1tVsdZCl4bofpIk7qe8U0QO3EQgL
b6MEdY+Cg+kI0zRlI3W/9++hTJzcSKluVc2WvjCwrjGRwtSCkuC8MzYl/3HuyfIK
FqbMX4TaNjNpYOsoZGtyfwTkZVx9usYstLcLlv4jm3/Jie6ZFPMtbrMEjMFMS83E
R4IPm/rUCB06cfYsL6FG1kYG77qMKI5VohWuFi8tCLFmsYlEghK8d/RW8DKhIA1T
t7QpM3Y7jDp+cwxanXmxZMSiRWp2wJwFJ9fqQfOsQfMKRxYejCi9Bke6VoK9srfh
7r8F/YGoowBsZtFgDkpWmB7jzgKWARucIDFgK5PQqlae8neYWOwuWFZSNYp5/9Sm
9iWrG3XDP6GPZO9b68IX9zu9/S0hwcF/++2eiZ0fYdkIuINMWQx7/DxGXA0ocbf4
aF9yIwOgfbs0IocIQi+iag7n+4lHxfZ5ik6rTKLMzjKi6SJbjDUBRi1w1KB1Jxeo
3ld/71E+UGLP5wVx34K0dbo6JXGFjvwuQYe79B8vOKtiHdvq5HUnhQovuHkqTPcd
DhyzW4T+RTELPPWlxY0wf9sweGXepPGwv0+butnJ+dQTQNKD6k4jrE0k1GyC3kHC
/PjZvB6VgC/K88ttj/TfEc5p9bdSV5U9sn0FQeOfZpiJFcMIq8N+vLe82rHU132R
zEA5q1zC/2c09w/zHdQJh3C9cPSBXLR8uEFmR+eA7YLeVUh2q4v2iv5YpGxF7BIc
u91yvnzzyedrLUZqgxdsrv+R5/XpVrbA2wGNX04XAkUgdOF9qxJMWb/TU8FgdH5Q
W9471CFUck59NBNkq0GFkIQkHjsstrbX3Byhjq7U4nyaTUjk40PhWomLRWk+V46m
WUVvRcKejpsCXKetcnCJWYHnAngsQm/35b/ZHBxqX5HSCxUqSQgSYA4RtgEfy1Av
SBbgd8JuwA5bKkSuJgCKeWgAFUqTmEH8OBVuBJcrP7I9qeginiRuLxXJIjV24sgR
ymGIeH5cuFuVo4I5G0SU1jJ6HxqPHhA8ae0ZFI71YZ4i79lUB8tnBr75qLR4qbrM
Ial3bjFHcvbgD65pT8UhzT/Q5Xyy01pa/WVNoDoAqX8ycb9l7ulmF4TulNKEk/uG
Gvt3Mt9L5jx+4uZVxrg/SGbU4Xw3eI8tYm7TRKI2Wt4U8C1VnTns/xwKwpjrD1xl
Nur1ycAP8hmnaV+35OWY3Blr//X/f8/NwfcK4FdhyQhHTGyqB1GLTWZ6H/F1gxQM
7irwtN633OXf2k7/yhSCvZ+NgCr9Lm+AIfYejkCke8/W33aG5P3LTjnptgDW9Xb0
/id+eR/BVa+YxEgsEUr5wxV2CxNjdnAOpRFFJ8Et8wJ2uRVXO0RBo7S/Ry7uiuL1
2eN+/4/W+WmVNVaxY2X+aJguz29t/UHYywfe8+SDYsTf4s3z4VOlPxDBP8g6bfQy
p5BlffUa5tFBwKv/II7vU2Fy7zzhmeQC8i1EPMJcHJn2Gey5RUclIOeXdBi0AUt0
jPBYKuH1Yq5rvOKH9LqTfoLe3pWFDIMGFFeNKfic1ApGedNBQUw8oIJPXBKyRN1u
Rwju8TTYej738rEfeuiCzF3NQBoO75Xt8GvPidA3ZW93/tEymciWH6WXeTj3AG1v
s744yqi4+pZUWEIkV3CGwX6iIJl8BT2C8eX3oX8wBkKb7iSVamRxIu0cGOFW9vz7
BB/YNiet9wtmXkqWLGMcP52/NSRCzQNrzfBsVQzTzsyZALLjbNBhIqoe7V6kBzNA
tNV0dKjM/I4ig7UigGhTR6LtH/rTL9NctHWBMw9TJ3lmZelp9mxmUHDClOBGdHza
0GQmqg93diaoZIRncWnvtoWveSvH/cWo7y0oHo62gJ2bCxbP4ac4sNLLuT/Iago/
kqZTMVrJWEGdTorl7oECQQn+fAXXH8DVRFTL+M+u1jt4vfmK0OCabBRYHXCfds9f
kmCee90Q1sovfTh9CEQeCfiSut7bGxeRT0gn08tISFsUJWPkoFKCPwDAdjzWh+8T
ew/F9qzIuKEH01nlZ3sKeFtFdJyWAVJtAbX8BkP5eySEU+o6w9X4TbFANzWV6m3R
peLO4IzpJTfMjrd7p8go76d/TZYl2aF1ZXvD4L6SJF30GwNU6T77nea2NkifqU3m
OmKYF2E7ICLwGx4HCPbvcX29oVOz57c2NNArr4p3xRqiDFHAmX2SjuicnFsVEs3X
H/7kvCcnYuXrNgmKtycUoMuXqc7XUgWJQPwQhj9OgKz+J99vLAWoFaD6TmubP3vM
oHLYnDCIGfiU+Ci9bqid5r6GF8LRL1e5/q70mI76Ig9j9t342O58qc+LxO+eoWHe
ABZUWOus2n9PJrRn1rLcyFpKBACUCK6yb+BYrAdcAkkNktHlE2Bi/NNX4iGz3j9a
CblrV7Zlgp41NwaLLVyD9p8CutfR4ZESlJ5xgyq7ISFWJTKq+GlKqUBSSX7brC+0
daAdqroLo0IotVkULct89uxXjbjc6gX/M5vHYXNemf/1RFB9zf0raxZyI76XgkyZ
7ZLng9JODOlTieY9F8Y7lA+E1aAyOcVUIPj9FLa0JE4Gdf+23u6Z5tGvNxEBLGr3
1ZeVg/yvAirY2cHp/zg1df4fiGiyous3MfEXBRIgH7cB1VIURmRKAKwICW8gZnzQ
LSMKcRm330uFv9otajHPq8I1cu1V0G6hj2Vv/nmyittQgQSzwGOfY7uy9S4Gdo9r
6klDbNN1rgvXRmRbILiOJ0NZxem3jamlF9rgx7rH8I80RDkCfPyFKw+UaCsnzQEO
R9FgzZVOPEBB6JGRFGVRWDpoMdF9PznnaWJ/+kG/1fuO2a83Ye3k2Yosesqdx0Ta
xzOF8pnp0jd3OmmzAbQlx8iChdQ9QlWD/HhZTNdTfTy0qL8JuF8hOqeSY4u/Bh3c
WvWZL+xshPzCw+1YM4yXWK2WXMErZvVGIRK5KidrpoZnlahGBAHLF3UdGMbKVfom
KEKqFNARfoFoaCRofCl9rgDS54Bw+ongoE8mrirZKz/uXqq20JTFKZS9KYH79OHs
s57wJMNa989Gio8e3/fym++sBUlQKJ+JnQabLTXPGHuOhr+rW+yFP87SU78FybI+
xLHOsrf7Pc7atjgBquTLXubAZRPUEBPkWw+/5c4n7gfXh218kCJ2Nc38K7ZbTLwi
IbB4fhpN+DlwONuHyRP7qBXyiIazR1jcdZ5F4Vc5JEhvbXPU9ba6zASXY6p/YNP9
zHJ8w3IUJpAwYBABORK+COOfU18FsGrbomLfizlKvOb1FSMzJX3nTsaSaWlbWzd5
0FtRSCLSkDNLmS+Mw6WLDnA7tSi+zc/AFXml8qWcM0vZp3ON2rijBppvJE+P9hyY
+IU9BiikEoFI9tZugOOjVyQs1/1AnosUh6KsSEJIxpBWlSaX0j8Z7wWUivQtMQ6u
8crMfA8DrzbfeqPueDJFYqR1Bt8OW+WmULMBpxdNO0lrk+xl+AE4e58vWa32bg4Z
ne0ZSzwabgT5Rbr7ivMB55Yjj4s0xXeWFIzFn64W71khAhRA4noEQs/TpaEzPBQr
pl736E89lZ6ynhH99+/6g/yKjXHTJcrv09hIh/96Fn7J87uBJ51htXhRrRywYuPM
K5Zxnzk9bEoIcw1NJmSHDegpUKz05qkqWM2akBV2SaDe97fjFGNLnFIDvvo9zrkb
p6k4rInCw/RNThhrKGvMitgtxmYiZTXaagpuRF1rl0jCBvr9Dv+Ej/fJuksZQmY9
J2IkGrzmjKrPChoxrVo+/DsqXBDFwkAbl5vgkaOpA68Rhw+AmYV6XO60ukKGGgbr
di64N3Unuje+hLeHY1GIxirCz94cmDSy6LhuQw28LFAVTJw029di3S1QlugG3FOx
tW+FnoJRlUNm2Rv4LR35JJnuWK2OJLqH9tstiM7YS4kpRjB2h4NlIjSbVVUfreMV
q4nrAd8if0FuR7G3Cro58Qapzf2gdcQrDueKdeJNGm+5M9m3wG3/qK1sON5AaQTx
w6TckS7cPkAEjwzAB4LFg+8z9iCHcn7Csc53dvI4SLoWdb/XnREgLKONihD9u47+
Z4g4P+qLpNH8+gm6gw+ygAoDClrwBe2zPy2aNaG3HV8O8S3EH15tD2vkjRcjG9xQ
DPiYF4fFNGpR+Ko7XI0PkG4jzRz+eOCk0M50z4DeiipDKTMuj7q1G6MA38w8+hP4
pozdm0ho6fEvgpZ6bjutBkHeVqPPDOLKt9bddKv7iBFCCRR25gt3pOWNhY5HvzZ+
iLf7LEHuueaNhBXxeRSGHlpTM7l0WJkT8+OQVPQY0mpD7Aq89jItuw0xZhXXMRSW
7x2MVZFclVKsuKibpn+W6ZUmcz0+hIPlrAAK6m5dZDl2hQSpj3CFsUSFWfpkWUaW
g3l8W2Nem6SCaIIopBW6uc4C1Ynic9dWUTWA9F7MF0pOYpaLwrHFFdiQk9nSJSTA
aw2G22GdK70pPF54sPQ3tsSrW6eSGBmG6NZNXJNcnfs3qcIehBInKxSFscmil0YP
FxPjUmAA/PjYFTukrW08qzW5PIGer128cbPPpnuoQn0IMstCeUpFzQpJqPL00/Sm
fVpZxZBLQwNAzBHutBDGAOpCJVZjYMCg2VjRj/exphqkS41JYNF0YIA/hg95+uPB
qc/l1YZMoJEbWhtWfVkbilfD+M6bm6V6zr5g5zavEjL+V3izhuNMkTESHH/Gi26v
XO6x5uqAl/tUcUxQgUlsMQPSjJywXkXvYzNUSk00LF+DJWWd7L+1tGXIhXPOwVLK
LgX5AO2t3fbeZM6a7Nb8aHWsYtCqXFcJms/h/PduOgtWhCaQox6PW9EsBz92iwKy
IHX3WpLdMiEf+OGa4St/ghuP0OroXkN7R9lqhSDnYaSF8w9U+w6XzbCREGcN8A9b
MzF7ZMDGndCjcBxwT432hdLYqvIvVAw/aWFerqEWTdgNCO5Ipt7mU9DYdo4G+ZHI
0jQRtMG7tMMJYw4qNc7tLj5pXT6hRmt/W0XPyZMPfszCIpb3LKx4rTrQhwMA36H3
4p/6OE/S6+Zcenl8s0XBEhttyKa+xviQD/hr/UrmEqD3GyGd86TUw8CxBwfaNvy5
mZt4rKVYtxT5qed9z/a4+/4B3vHcHVJuM+gnoBTPn8TswaORZqOZT29pjf9MoIzI
0ZKujfnCWEel25n1rDPz2nkYaLgwMzbQxasZtAqIHhhbRZGXgQDZ3e7PsfEddMr/
44vky4jT/PYe6+f7xsdFiETJQ1IuoKsxb8ewJwGYPXNl/k6fccNWUWuW6o86Ivtu
TD7BdgOcH040ojVwpwbBGjg5QsrLyNBZbYWA/X0BGoOaGDMWw03v0jVJ4TUgM5dG
kndahJ7+TSYZ20q1gLRFzR546rNV2I/yF25Vw+pwexhpHzOXD6Jo0RKeJoKH4tkJ
WDnpZkiU59iAvIuCy2APZaDceNPIrUklCDINDCxcVdRtly0MaK98o5X3Y1VLwN5q
AJfwWVo8gZ28UT0VkJfCmdfm5u1AUCerBDXV3il5kfiwZYcMzkp+6eldz6+dRxtV
LbXtD/PsKTlkyj2AM+zxvrjG/WA0iv3qexB2/DveLJvNjvnumIRRV6FbF+oES2qq
++n//YNUsqZt+pERl94lk0VfFLB8Fdg/ynx3Hc/nDklH/z+bkBu9Q6plLSiQ6Gvg
DGI7cBTFkbbERood/Mz6VNQlaOU4BCh2qcRbzB2rN+OnZICP56TiCX2EewZDQj6c
RQS7HXLb5lLM+JluquW8CocJ9R+CL/94NKUmnHVnyZ2jokQWC+2tSdWtVf5NLdvi
2yo/7YC0FU3VBQ1t1MxfAV5DH+nfrHWKziq2vNsIjeWjF9l/mS5Xo92Jo6S4D+qK
EBrTD4tsypTNtstcjFlpKZKSQ6CDNh4tWkf95+V7K/E4D+NcJ0QyYvvY2p4dI28V
Mq9e+7QQ1zgi4nuyOaPQw6DFIi/v70eotNcDnRxEDcoIiEWDkc9UHMRU/Y+T88PZ
TiEoUeqw0M/KwZN/tLfbHdRK7YPJJInuw9/p6aEPCvoiwIQ14SAhwqegsoe3zGiH
SNTsEcD1xzjU98QEWavdrali5NtkJ+57wV8thr1NumS++u/uy90s/l0QivZRUM0F
70lk2OHhlo8lx5USllNORPXiuRXASSWukAdeKwvOQaPH63ZkDCb6ezDSOf/XNkBX
Wb1r8F23FKqBwc5xsLUZ4/wapPpWzcjn5MrrqTX/0/JnaO5gKQfLJp1iJgWYw/Dp
FoUa208Px+e3Fbr0IzvavV9h6esl5gAh6sYfOHWYaYlBqOH0p2Z4QioRdNKsLo4t
c9LUgkp+q6HNYlzku14wDdVTvmsJAxgOwRNhaY3TsUwzZXw2Dl4hjVZIqWgjzzdc
a9HDyNuFhcWWoRGHUYq1zEvdK/ROzcpyVxAfgPaBdvj8mljwvZ/ex0Iz0WLsdq9V
5vyYB7Qu9UPga+wXEr2RXCaqJOVwfpxM73zWzo+JgSSzaXHNppI/8WqqFudysh/P
mFfRrVIl3I0bS5uhC17iGxin5wF0u8oWVDIHDRPIroHpo+yIGDgp5bipICra8TZM
axASBrBBwVIN2FGcZP3/NZaEGkYh5fxh2o0WbIhXgokwL4SxMOMW/MbKSOd1lnfw
i422MipIsF6t37/M5utNrvPiA1sD5MFSJLPqyiUILSLcKMWx3vJPWvvxMfZ3/gNC
1MhtMRZpGt1ENwNX0FlJK+Z4/cPPOPuc80FRHuQiCUUHsXFyBPGpwGYwKW+yj++u
pc2pdx8bguFZGZmkDTBRtMUDrm6TkGtzT2bHFOVqTa3qPThpmruPZ3/+bxOB7zM1
p7qW73CINYmpOLH0RBCv7ZEeKAnF7Go8xgt0ipxxWWrTeQp8TsH9bcnGM1lnp8Ei
uHAy51SwISKGecVBO7XF9atqxDtlaibCXwEIZzkVmj7+gnDTk6MbrQIFjt/4X+TC
inCjBL+VYjw4ya85uCI2fDvvjxR4XhG/wylczcglijRTGNq4HdtB65Bg7ywYmvbV
ABG6WIRvPtCj51vJ6JRUxjs+4UdGg/QDt8Ft5Xy/QT7gcie9R8wzkRq4AnUNrdax
mvUNtmEwYXINhrzi75y46GDMpcIr4FR0V0nctGOF4hOLjgf59uwfBGdDe+sDeMLq
WJy2GjvCoKIT5gGeTuLf8izGOdKeKxCu8YArMMwVSzn3A5PtbO6+RQNKkYxNPHZP
Z+SzP0sBA8ZnFcyTllHzsL2y9ik0ZlwWqYVEF7ysZkCs8MjkNgNwJg/QFtanMTKS
HMJ1HUjUqkFZ0zh2GWTcS13NpLwlJfQNR5X/t6QEuRPYBEtpf2PID8aEYN7K9FoJ
4vaSq54r90rPWqVGpAHlwLKg2LqmfYD4pSogi5/yLjhCjOAbpWjyjcjm360jvEfb
Idt5rlKHiFvDk42jaSvWnrfX0gDxt6u9tdG3vKqelTryAUco2Mf/K9rAzPHUmkFU
4lHbQNOoHFjpug/FjCQDVZ061UWv8f/GMDSN+Jbug4x5agC4Axtx/k62RmhTkGSk
Ttx85+0xuoCoNIzUAkbnR2C686wqdloE3KEsrPFfJUjfOt7hfGpDkc4AVXIV858m
zpMKX0rhGAVQ89zCFj0LVRIibb8psufp1+lvefvPcSdmkO9/WvCZsxTxWMCYOP/U
Lm5sbbLk4jbhzXQ76Tf9yA5Yjwv45h7XJg1bxLHUEqGa1bQS/e6NmvZaRGuVC8cs
wcFbwprRy+OLEKq2Y1sKt+Mq1P6aL8EwOAPPz5rN2jgQaUZ7tp2aHsrqEVRPGfSf
OdNiFsAuGOCMOQTtY/lRjRfdf7QWRufVa1jG4RviUAGjaokd7vWlSSbh/CP7dPhM
ypuuk6jo5U1n+TgbKXq+0hSpdutC3QNb0lFoEhXCFIDN9z0FU3GQ+blVSF7y9QWw
QuxyPaAoSW4oI+n5r71f2hYYwFJVhDi4jOX+GiCk+8m1xjSA+Ui/4/JAhk+tKc7t
kLCzovOZclE8D6rCtpetSWalFsf/6j3+8RbnGMtW2Nc6c/cefSiYg3cIJDP8fAd1
OKa6Dung9UAYZkoO1Qvl4KBk7mwGIZbkobLdoQ0e7nQCKBspoLhoCWf+KDuJjAcc
SAfp0GmhmPtno3vhGJMF1ZMrvlAacPq2m/pm9dH+Fq4pA50WBEg41Jb9LRtY8gQL
L8CFwRjC+DOVsJ0VSnYbVJmbwRgwaZdCfXYQl+/oXLdwwVICRHHI95QF8ILww/9m
IXsIKRPV5Ts5u6foMqC50qWAPBWiEjhXGSXxgg3ORgHyGpuGivHMMFCETMnVuMoR
bOQ+kT9+OLDVcxzc7OGiylm7PZi/fGIYj4VrraZsnHFCeYMGSr936yaOHgW3g3Gv
E+HEuZcyDnmmvoRtPE+YUFUEXWEJfJL9oX9YvMeiyUCUmxmPVreaknhe4P+rsaeH
zQLEvdYpEWDbCqOK6JI6O7horB/O1DnhBc97Q0oybYJeUwlWI0yuNxlf7vM183wx
O5Witlw1KpVxRB6SHdaDYbh8LYDcjd5MinR1ANC4bPDgJpFD+sXv740fmFJzI+Vu
0kG503yQhAs9r/7MihabOfhIjMGP7nhbO7EEcxiv+a1jzqmr+/PCMvkcJuh0ql/j
+spx0i1mAPB02rgxPLpCtUbvqR1ro5byjhxL9zEx2QAPnxZYi/JlxLTM0IwuRPB0
mYFGInNFIi2izPgmvJjNoCnMw85grulgnGpZD67toTjSR+aAcKzqlVFOCVVubBN6
ygdtqzrMCYnuVS3F7gGUemF4IBESWjLkgFHJPmSJxshGlDLsXtVsMO722Xpysru7
0S97UvCUEJ0TXQDjBlketuaxRGdPsK+6UUcnMkPIwWgXFaCqp3TjYdp3olhgOKqs
0uWBlLst0Sam55rULWjM72ZwuX4v7Ey1kN9yV0MQ4rSDfhFfbIyVBlX7mrAF8KRH
+a1DS5mgxueqKpVXsZ2pUdo4t1cKHMhO9cwlCIyJOFdNldP4ODZkUMW/qB/31C/q
+MxCn6/QFD9cvQy/8qATKv97o/rkwT9wvDDs6Yc8Zn2EqLokinS4Lt3k2p4ka9IO
kPWDnIY9KMMjKRXOyOd6KX9++Xmyeo55SJozWSqpHPM3EmvArdZiFmSBliG+jls7
YLEqOJOIO19R057OvXBFI6NiI6OpDX2Ya1Xa0nES6lsnqeGKTAlIaQi8lBxFKSg3
2f+VaQS0eGudS/sGAziBG/K7xPai8dISrLRESkJNdrEhc6BOQ+MaP+Yy2kEMoNM4
+geE9SdNboWWiPEgVpntQpSjyv0CSPWpzq+Vl4o5ylse3a9bI9qiEthHHJzRX4W7
1vYHmBsesl3loLNJaiFWG87HiWwkBc0F+LqbPBgC6rxv9+NlNebjDuuNmFn0SB77
1EBa6W2Uo29qka8FD86P4lUsNZaFOWvEnJstTmbJd5fAOzXfLdK0wnuUXbGK++XW
5YGdFdsjsPn4jArssKv2bbV1RRj53ZIy1VDP2gCh5eMC9TrCl9VSA9LWwzchA9qd
LOnACY+ipLlwbjqEXI5Q8xqnM4pe5nt8MDuu5bia21MDmfTFYyuQzcQ0XvDCm0k5
Tc0aUq/gDKYgsrLJvz9GEWAzfqmxEFIaHIJPqLsdXjVGIB9cms/NrVR71t2QU4JK
4UKoRiHBi81iZjSFt9D2MRSamj1TnWwEimsLiGp9Wp8nnygJ+Nenn/My8HkVTRMi
NoV35/HKCrwlM+u67JIMzSgJDJDrm7bCmReBj+b2Z2xEBg0gfWteM1W7dDpkrfa4
R3p5vl407FvEwuphJ7YJjuhkvJvLp6YAH9WfAK2+ru6YQHRRANpl1TTslPWOC086
1U9Ya/XNiu5J/FZVebKBqRrHyzMnhp7mlQdTEijqiCQrp1brNGmwv7WRqfVsu6LZ
jZYZLre4U2gKFFJnj31nItzLH9gu1G+q8E4UBBx+AieB7a5As9mvvTSp+k0Tu6ga
hfLNdaKPsfDV4VkgKD5V5SXmforDmzXZAcaYbuwbc4n2hml1UGPIWSRDbGC7G095
kUHJCCY8G4XnAeTog/4OhJQb5cJ8DHzV6Wd5JJMpvsVmRX1hr8La1r6GjKYh0Erh
s0YZLTJzOLEIjpNMUFFFfRvQHFqLEH0SYw7pW1gU7jROSUF6y/0nQhinS8pPbYEF
lS28C9kcwX6A2MCCiVlI8ziX4pd/V/3KxOxto7135RKsNkmoraXstqqkqLWyWbPq
4Jp54HCHCJ+0GGH0Ckdmz4v7K9oP/clfBIho0NlV/z0IiEpnGkrqKRvHLK8dldaG
5ZSQ7mv3wGUykIlDx9eGgpFOzUuWbR8WGL+EzQR57QO3pcrrDouW/TOkyeeB+IWN
ot/w84phVduMhGW1bHaUXClpEKpDUoYtyU5Fu75+GWlpf3akUZ5YwuDWRD2DhRnr
LdDbbBIoWNpA6ZBKlttu04spVdwWJ7kJ3xc4cemCVlr/5z0l/NhyrA/umpPFAzNt
PThVnH11f8YetseqZD3WaYbNKAop8Jf0ZUKf0ORED5KqfAKYOQ9oD9O0PEjSINa1
mSDSfUm1iQiQST6/6no7P1qqm9H77wSBoQuAL3NenR9XesYiiJcc/ArhSQ4Kktu1
RmhRcxM2JjhnRTgJrE4bynkNFVlb8TsFrP82s7Iy60VlwtNNeyPZC3Lu+fZmFi6J
3wbVa2i+WEs29JerAnPDF0jVY057UoaEG7RMcvRWM3szQf/noVo2Y20ErKO+01gY
Y4wwcCORhVozQBu+Bq5B3zvvES0H/e9uP2+UzehDBxon5EacEeICyx1EVLy660jY
xZuWM1UD8cG/zZUxDBay+GR0cLhX3UrohhegABuaAs9l0mtXjtZKFDk6JXBOprVK
S9wmigxt60AMXNeriz7vTMyf17j0FJ9vWmiy16Y9Yd9YB0HvZUw3uurtG8IcU68c
dyuva1limXPdUq/MLRcq/Ui04NKVjcdgUryI63a0f4b1FQul+KNKSvZut+68/ze/
nlsSDfHEEc8TJMTz9p7+IvaWB9HkLcmm+jw8Xlhd2fqoWx4I/1EXjoJi78RKWHJv
khpju7XJLlSvswac72LLbPgbCsbPOp49r2y+fafH+JvyqK9CBekNRO7zpK5bKJ+d
shNh5BvJuekigveVIHVfJ11C9X+YwoDPSjOrv87TI4ZLbwZklbUDpCzoralgIuY7
KxCbyYE917EJSMiDeyjrsY5YwNbNNNLG6i8WdrdkTTyJc6JpSqe1cS6jxO733ciN
DPbsjjasVErfBGp+l2bWVaAkLpiaq2bJ+Ix0R2fFjKvJb3NroLyPV/B94fQqtQ0H
CTiEU9QEsRHxn9I666pk3r48js67H3LrOR81JKq9QcChXhq9mqgQsZE47rq9NRRD
3qvsJtD1e6IKBG7SmldrDFuhdzMt6miT3VIZG9I/r/cokJPLhRLdzEPgSszZzsm2
97OLNvg8KdIZnPCcB7ionn63rs8uAmC6loGs3fG4/bRd9CeKmQIV0WsVhH6q6bFL
28WSreOdywp3/FFeS7cDROVRTvqHl0t/z/qkYsqQFuu5c4aSCtpYEUEHhCu7IHGR
8kK/PQqrlL6D5WS9wIEaWOHKEap0uHXW6QPvaeidoeuHokgZbzAMXna+qA/rx2AJ
Lew6TyW/bOBqZR5EwfvrSluzr+Er8Bsh8S8gmKe7/Oap4k0qm8B2/DvCbOGBndXO
hSN8cdiP+0saHmLALJ/vTFamR3Vy3cVwX6xXaNFef07rLPhpn1vcNTzad/jM/yku
5+rPtEX+ehwpBZ6CKj/7O4xvbCMfzo4BTfeX0MPNosF/EddeaeEnbgDQ262LesO/
aZHiZbvI82BP6G7t4NIcpDAXpGtnrdATXcZixpd4FKLlU/cOYb5vfUFGzpAbi7is
jBRhVKlOMWfUiCjSH+nqaIoqBzAsfrJcCFCBwN5SRBBlX7HVg3P/1yI0i+KEODqh
B4LsTUlAETIUlcosZsRNMuY7tsbLNNsmIIfwNXdU+MKu4Tzv7qMUNv/DcWHjaMkG
5pptPRbGfVOMxwwQElPLIi29/CXviJRigiWka2FEU4HC8oIIdgZBQy/1oICKRCti
TVivc6qm+FloadJSvWj7AcGJ3oU8dEV8WzWMXeRi4RwVTPxYEYOXlNJGMUwZl1mR
rD/URw9AErS6N8OrZOP4dvG9JrCsqI078JFTr4KHfW5cfNkyAlYe6NZ8Mr4OOJbd
AqMZ1dvsNdKbbwUpbHKQLY+WTqBtASs2hgWjuZMgtHZKhPRVFz6YukqL4c2cQCSe
UxI0vM6SG4QMmsfRBBWM+yEI+sy3Wb6SB+P4UV/e+P/eIOyt3uSaY2MS33YF5TuJ
EN/iSHEt2r9OFor9oGjh6VUIusHEesuXx8nDG3AH1U/WG2aZjQlsIvLvbHbzR8LU
NMV0rZGYXYeHmmZI2IkHhO1A8+ftqN6HtomieCY+Jjz5Lt6lj0RP42XiYYHSgBM9
tyII2nbKdIWKf5qbDF4hF4r7irkgp3InkdwIRoxdVrHCjeB1TvKF70ccBeCgV57v
BWeVvozqhJjB1XLwn0mul/PS2lb4cEIeaIJqxLC/0kNAfkiXxjEHFAQXwoiuvvGe
U2giKDKqja5zr2Hl/X/vZWgY665FOeG4rOF8LhGUHYkSaQnqSagE+jGdewys04Pa
ChETf0u+hdXWj1+IS9v7aqGp+HycCA/Ye+NTF2Uae1UKk6igidpVn9ThrnEB78yR
YTmX4a/dMXAFrcJpYNH8XryNq0Y40c9ZB5xPAggYhRWvhL5HCPpWfHG8mjU7ab9Z
IDkEdj0K+PQ5r7t6zOdygqEkVNxeE67ClHc9H3yzNoptqEBem0veKXg2hLf4FaOI
oM7pUknV+OI7IwI+tFc7NOq2aGJUK/jqNU5hyQrV85x4wQFkBITjSDM8wkR7CgEF
O5tYLi963Ici58MrT/9YvicP/UKhofwhVkI/Hg7lp7myKGCoZSDHBc5cvl44WMYN
/slU0DFgaPWTiXcWsBwiawhrJldvxXJKJwL12cO8ikuONvegmFHF+WopMSQ+FtEA
GMHheg2fUoaZ5Oel5/HvaaMJU/U3qIfZYKgMLwVKycSkst8GG2fUvc5CmUMC5ZlQ
5qZAMCgXQp+b0N20j31SZjT+DxxHAikbxRYX0Vts7B/rLPA04UaOCgXgn+ZsOf8X
bOAP0UvRE6Sj3ETlJIRjAUlOk/maHLBZ6T+uFjAB2z7NIGNxxWcylXpH8NjQdfC1
nfAQrmv27o6nbvelxRl/yvjkqsALqj03CiK9BXpdFA7pNa5Bif/RM4G+2cQLdXYu
eNXlF4n3Cn5jCYcpkrJpvIxBk0MoW3xne+bpNlKvdO0MUZnJpMBic5rosO2ukO42
Hz70RqbrLD7sDxcKQ8cypQmx9KK6J54QEU12997fnABAmAxr2hqWbiDx02fVDny2
dBq8iQifT6Eon0ufP40QPBi86hN+zyF7r/lmUFGIoKzVCFv8twsIdKZ49G17ZDko
F9ZswxdUnKWBbIv9aoOag/xbfwZY+UBZO+1w1LTkmdEzvDM0CM88k/VDA/uaHTE/
nNI/ZYyz/kOTdsXT4IlqFFSDYU9wv8hXQ9UqQXUyGVwKuEe04BLzgzlBSQIy4tBY
rH84NKcQkof8dyDAELhIvOEkNvvRy7gb4viRaqZ4cQxnCHV7QG1MisbkaeHrUC3k
WdrH4HHPMcPulX11yN32a+uLGNqtUV3QMMLrXJvKivwWqnKaXfSE8QV/hurrv3vi
LM3x4g5MyELiA6YPdqDyxwYTk/9dTmyhACeEayHn1SARfH1STO0EobhjsQKJcuvx
3RhgVyB74pbvo1AZ5wBZUBHZcG3RZUUkK+P1djJRUZCduNoqYEaSsLTIK36k1z7A
k5mhznt7Cqw/GQPkOjH8xX7hMD+7TDwKj0TtbBihuREn31w//fc58vKxCsYvGMu7
dwOUUChYPERb6At12ic9SHo4XD9XDN+zSjyPJPuhiMaqU+pA9MLbOFxXbK/9Jgyf
eoLHexsWUTl1bhIW5VKC1BnIUUD7l5tqsTBpwUyGQiHNF1ocSnOxt4bz/lc/Xm3y
I6VL5fVVJ4Zd9P3U9A2ZYIa+rwUhc4pLSzdD9GaJjEf0vaNutv5xTNRfsBe4jU8Y
G8OWwPXbQu8gvV757FtMl+hUYOC61gMJujsopN2dlmeFD4C4nhf/4nff/G0ufhL4
RzPplyMNR6NsSeDloiB0yIp8PlbHWiz6PbU4zXYnOrocK8QHw/ZPZTjdw4ELgxCl
dv38Nvvix8yvvyNsSvCJynM0UBxZc2xVqp9Ll6fMb1HyDenXhCICpYIZir6mLE8A
KseRQoEoZY1YZTNQkO6Nm0Lxyztg0QiQlECnOS3yjG6pZSxwYdLlzrjvP6hj8zbT
Gljpl2CzkSieI4nFClaG2yHPFmArSS9ZQkttIqDfeMgO386BvctNZMLc+AzhKoZr
mB00S3MY4ouFgc2bMwYqVgQo/K9Hy35rGG6RpmOm4Ul+y/ceHTuIa6qfF8zPml9b
Y/4GA5xXJyLnWMZLDcQSiEPCbXEJVwlvTX00j/sUvLH2kgRonsCs8jzmGUk+UBUj
ZrIHQo0kRJ0/sQDgdK0bBzG0uBtM9EZiRYzH2rpCu9iySyoiX5wR0TM9lbslT4cK
ZuydOs78jCAqXurodSCO8gAExCCL4IgbXR70G+cuepojyrPXGupcZLZD10GjWh4i
8jTb3aFrwgPbD9h3/6CCWuQzMJROo9fgKcH3sP3JpAx5AAMXBJYLZGgjrwTZ4hUK
0ILrtKUqWf5YFMG4extIXL8qgrXk65bl9CztvdyLbESl2/RPdPRaq+JaO4dMC1iY
tPvSAW2ViMLXPiU/lxaH+cdfq1wEkej8deM3oxIUErdINws4dxWK4tUlxSggjiWh
hGZd5+AZSwrH3iWmWVEbiRmDytEbdVhMB/YGypGdTlwzTeKV6C1hXU0+uWNgERtP
rz7rl5vZF4o5xsdG/fuZqHLVmy58qHfK9RMR5HSe+gzC80Vwt/tPGLCHuoLfMdso
fh2s58LCQ+jK1SKSEaQ2tIq+M6B0ao1gdWO4BfSXhEyMiFYLxYgq7rhZ7GpQQPvr
O2iMB8z+ezNNf1dl7X7JRDN0j8D265kV7l6bTZMVyuqg2zaNS7gD3X1xkdhNE1tj
rz3X9+QnyQNYvj7mLc0naToHgfFbo9L2NKgCODg80g7gpSFRoPYalql2AxQaSLty
mdbUQWJiWZa4AxqMiQM6SvGP2IMvHTIjFu7N1z+e+Wutnsk3tR9ulFXx8QPFTAwo
ORiaFVDA7eZOROue2RGsEB1FyCBAB/C+ZS0FP2/jTWyoTvKHaXzi17RNuZ/7mqyy
M5NxbYyDzfWcdxF828xCylhEWsZP3ZKqZ5W84X6KqqceMxIH33J/RztpCPxqQbjY
FIxfdSW+jnB46ZhSYDdJY4d6ZJ7PNjQfdr87Hx5tLttQD17f1ccO1Wa9JoAFFlCj
o48zQmqPu3sszBhbmMfB7oTuQTRijKrraIthZLnJqCM2rDdwrefD2JlnJOMhdcrd
vjJ6DOppmtZD/FpMcgXJChT6IHCDhivNGU175Lmyc7osus0c/q415YWcAwk8k3r0
X7RMWkPpYQn4Cj9NXA06JDUGdKMXPZxEuh4yf0uas3Iw54esxkxfMumgWlny77ou
S67VrsrylP+ZbxfMqZH8uQ52KqbZHUDKzCIiID7nw0Gd7aZ87d0TJq06ZedcptTZ
BFY3JHkUJd9si2UdoCD5Ufy9XDxm8cq0VtAIzHCPO5FUsSanuHdauy1Za0Rpqc4Q
qNSGaPggH5PN0FEBeU4TX6hs1hKml6wmS34uWG/fb2W08gFd5dRfZGs/DGgc431U
PguilDfIZJZC/iaNFHp1Pnkh/2H7LVPxYEaeyVzq3SS2tUtsSNk3CUXTcS7QL/5J
01ZztiO5/Z1EMjZNFDLawAjlPkzhc1b6sBDOyQFqx/36tbmNe05GJW4xc6vkcN8c
r3l4ZY1Em5YRT7oABORrsRZbZbIiJ6hgbPh7pJgYqYS3BZmGn1AYv2OyPYFfeJ8x
afBY0LuJipLnrhrgWb2cVmKNw08rYsYamLCi8IumQhe/ALYob4YxK4ONgeZh4kYC
caJtPjUFFvcTFNBkASGr8lQeYuyYYMD+brXg2n3e3R0S+uCUXUoAu+vFcRIgY/ib
qHMzSz2DdoqGS8Fdb6oLNiNwsp/wkVCa8ORrmwodliFUytNfJaB8UhxxCGZMY+Jy
89oeC/BQWsHkckuXlRU5O8smZcv/Ekcsh6I24JPiuXbQocrgDjFkQ/e4vg59Lkw8
n5fEw3vj+nGWndyr+ndwj00U8Q5Y4WkWbDVLr0A+MXlDz9/z/maQInuHWz8JknNd
mWvXXVkrNbCKBAznn27NmqC8N6Rvs/GvcdKFyaEZyE/Q5wNLTtf00vGk2hw2OLXq
GIEknD0YLlZEVybFOgOemKZUJgMyXvyrj/fqSOt3nAXjmHOJ3OamShiFpEmdAxmh
47x3KkDGub2GNEdukJExWS2rZ985Fvs8UzTaO4BUTXtbzd9DR+puWNkmqOLb5NYb
XsgQOrXCzyMYQkSdpOa8elvseBbHOSMJQoU/novcC+Dr7U57Bsg2qK0IymSiWFct
RIdnvU1yYJiBjOibyhmlgTxTcore8SlNtQ7dHYr2WqjQII2RDEpFlwylUzQFy05N
pZvvLgTnEG5fTJbY+SMock+AwcXli9pgy1AkjvWUN+10OCrIxhL3cOFIbJf8nWpn
AlBWSq0njOtElf/VkLqOEF9DpagbxN27ByE4y+gCFCEFP2fRZrS0CPjyo9RnOwyx
BL4kIaLGoIEzwQkw1axmnGEXusNAbXSnHH4eMq3cleu3GAZcFlrWeLoNJr7e57W1
8J/JjzRGOBQoBlARqxx06dSZCU5R2iySPUP30o0SMW4fa6C2Z1Lr5C+Viw295Y8t
LygpcJbzfJ+bK1ejbpuNjjiLv5Tald2KJxXur7PCZQWlwBE1qgzO1FiWCFzDdFyo
AxLK6OGUBC5k74K83RRDcnhBjyEgg0OveC4fK6NJjhikhD4k0AWsdh56EsPGIMn7
P3zrQFTm79CyRDCvyWPBalB2Wf5SyYO1AUVCM9BpqJwvyYSidI8Yr+jrOtScN/l2
wyRBmZEHnh7uDbfR6pb77HjfVfMTqYmoaiw6xfgDoWPmjixA3rd2Zx8eTrxBf6u4
Tdzw5b0XiK/kscbkJCCDq2IP3ue2o7doOkB1oe7pPya8TxmxzTc90LMjWuD4S3UO
UjLTOqRg487IH0PcMIwWYg9GpM4vuIy3I8QobJdHLPw+uEXpIPExk103Fm9SlZ+Z
UN2itfsryB5CLbkln/QbqaGEiDuqX1wrAMxKlIdXflqM1ZcG+7O76X0pEz76ZTBW
R9nHkjPX4CQ3VLZngh3Sz8UOXyVRZgWmQTROz/lntGLKmX3VEkmUbZf02pbH8e5/
Xo3zPUs6mS1ZbSBqw726NdRmB1YKQaE7pN3I93Zvis8659+FT4G0xTkLgTL5mdku
ENMCuc1E0qVKE3N96NHy3HGgN+tLORtDhjsMJyEE4YN5svylweRzjSp3DKuvbDC5
AxSH8x+QQOayXQp/HpMsvpIzW7em5DfkRhelk6CplNoJ+sN19796+lzEqT9jYaSs
Ea2aWvo/vz35qf3LICLsS4nwW2jxrU2Qh5e9/NlSVylDkGVX2eS5tVk38Zr/WSJA
khH9mtI4nLSrAVhvKVOLB+0FWPI8W+zUBsrSKfBHd+db1HjQozp80vDSSSWh3M3b
WFZJChWVJWgLsKg9UAmiZsAtwFiyrXUsMH5CAnK74f3b8UFtuBm4ux0TU/MntI0y
NZXYqKTS1tjovuqgL6xVZz+4SkERyDY++hGb8boWxH7Cuq0JpB7xOFEXVORfZseW
nXg/QrtVT36yghUWV0xhTC+bQeFHahxJUauDYuxqhTzpT3dAU14a1FUb4vUEsN7Q
H20RW3vtG3ZUehD1zzDXCCKOvtTATG768nepReXnF+7ESbLAD1bMZzLe0LdzYWVg
pjsvh86QDa+MCNgsjeJGFwvinVBe8guH+KyAtDLPJ8HRcwT3gE6hJ0hL0ODJmrOH
pey29Z60uoL40WNbY87+dLJGDZdnF4jlwIXxBJmEzkhawwOjhtm18Or9g9Np6kDg
7sKs9mOcQGbHKy2eXdTpoDuX+vRCCZTEkSJsqaDZVNKRDgnpCB87mIe8dgP5qzti
3hi/IGvlrEZytKqNKcJrJt2figSt7vYFTw2R87jc6cfhbKOo+3ByrIfxQfv3yg5V
OeWHIug+pydHiep56lQUwEts1oMnlQ/g2NmOjNpR5sa9i0lKQ7GGNCDtbGUSpYtU
hlajW0RXw8WBkDCLFYzPpiuwmk1YBtTC0fUIBWQomu8ryBTC30O8GNCDL8VHtfOp
6AvURnP4GjSHh9KZvFk8cF7oQ9mNXhwWgZ4QvAdZUxjTndywIzpWZ8U0nvAwZuBx
rUmFglZTFDHBsM6etJOPOYm7kYpo3wvZ7/un3dvidNnbHR4PBi+xC96r8CZ052lo
mrjJYgwGG2RWnaLylcV5sEfyCiR1GBUCcBdLIJGFRcvyLtKq1F+Ynb3/xkCcKH0Z
ZIw7Tu95Kpu9F2rCFxHtFx3eqaWEFKxPK4o+L+3kUqqd3olzQMDdT9wtTC3dwv9R
yfkHg5ov4xOCx+ma4ZjFhfijXWuI0luXpd1pBqTjD4KHb+/6lSYAvYYmZc6rJBjR
n8JTsoVgytLUw/zIdk4hBr3WIbxPKGb00/h7JSEXGTbJVogrt5TF4okbr5Jd9dw7
+wUHN7s2yGJaSBnqqPHxB/Do4ikoV6DfbWw7Xy/l0EyNw3/cy7mdrTWm/TCaNgFb
/oIDOk0lbqcXOWweNTeHMJx0bRsMilFtU1/uy6dkkVoUzb/PEfTRjhTcfTKv9mqy
iVabXiuPthKCy+ImhA+YsWqhlj+9jhhMCDlCPItpiLgsrdWKMeg1BiTdeLMQdGZh
2fX0avF4KxV8J7TJ7q+CgrC+IU8uUzp2FcTJ+H+l34iUkUIG+1ztQol6EXwfg17r
ZR+dMCIjs2ph6VnvL6gAmGbuJI63tdSzqCaAruE8IbS+GBImNU4AVfS5CWbJl6Ac
EMDNC9C41vDfEvJsOZwwPmrmiVORXh6wv/dJuPqzTRoXcdpm9rTHsU/tDTRPI7Sd
f2eGfp/Tc6BRx0qli4s9XIvt7DnRpUlC5EYcbQqsR9UgLVYgu9VS3VOLgEwWhYlT
HfwTJMW0LYccH1u8SwzQupo+0n87I3da9V3XtqjfFNENArwNaEuOynjfPELVa8sk
HZFovzpzylt+xoYPiMtsqEe6e+7E8zyOel8JJmExVTwOJHp5lw0e6lGN6+9XP1AC
t+8UrJT5JZ9B/uq1a88mW2kQLpqjAPGcyWFzZMvEZni19XCZKfZq3pZegLlaSCXs
jMYQCI7RgbcrOt8VOBI3Nm/pNivZa8baGmZairDd+UKcojO8622S/55QPUzrS6Zp
BcAsdjDrE24C7oEu8j7snkzXX293dxZA0Oy8wRPe9LNG68gWXsbLMJZOAbqQcsqi
S6wjZsfdVcl11bbvlqmYMpmXFPjqy6eNPZa8MxNL3IuLDssBaAf3Y75ETwIRTRze
AEwyG+aU8NGXEbvejLs9kc1nuXSj74Jh64wKOV90CUcIt4+3U6gMMNolzPXua/NV
rKzCbA/eiL1/5Wwsd3rmjtlSI1t60IKgHg8G9DjDbsi6Xc1yIhatbylAwABhRvP8
sI8B9ZzwsAjgnUfojtKJ9iEH6YcwrcuxIGyt3d6He2ZPMKOnaO7mpw5pTk0yI6Kg
hFGCI2/UV7FFpHM9pnflh0fTgXHosJ3CEBNxcWPkRk7123Yuetz7tq65rNuayOkf
sLlZUQW9sBFYvkPxNKD2eqdy57LApzn/1eEC6I6buzI+P6Jrw0IFzwG7mgmS4bpA
V7eeGVBB/5OpG/pVxsFdo12E0S2fV4bHQuSeR4bN9kNCW284hkgGkRfIqCqp04ZE
pEbERP6ZoxcS+E+iqcTr2zVJhz/JmRdC3rU32itP8gtL5h6GhS6YM296DsaXuDrK
PU8C+fqoGY+jraTpGnjEKpHR4/bGln8T+lGm+ZRtLIcG7bUwUzWr34trBzjGjeQv
NrEoPpgGGYyFUBOiBbj+rUM3vtOeite30NoL2R1tnIFVSHM+GIvGd3tbDhKJEC/I
MO2hhNAwgnTGG+GPZWsNYtYuuWZvCnRdPBMT5AhUJXdveqTjb3agpcKyBcVjwiWB
HQVPUxxsTZgPVOG6FjcZ6uc8dWAtDe0mQ+Ve2tDxDN/EPl8XX8q1Uftq0ZhCyRKn
oU3KLA5M2GUOokQdzKsxzkOCdklP79gmsUApyUTsgC0t3PG69cqZIGz5yrYLNYls
zp4idzKg7OKvu/BrjeFLuCyeBDbE8Uzf6r7yAYWsP+W4Cq0Lj/5+3Eaxl8Qc0kPi
XEsX2bxNa14+i8HQHQkBpNDpjqV6ocBANzo4w7QvYV1raHO2i417Ghev46guF4nN
AuAJWSpH3KWvF6ue9mojEQgO0G6FuEmQC3+P3oegGhknr4cmSL92AaXrzxecEu4h
PwKzlnQI2dP39hTDvSakyCwhBuGHKt31k8NdpehSBZPUJ+O9CUajrGxIwWIcJP2C
+gLqhJijxFmFyBLHzsqeeoH7HIbeB8AdnXuWeLpL7/i5htxR/FL3uvJYiOUGLoXa
oMb/9KN1MYZWUw6s7KCO78W6SyqlFJEXbTR5SR56guW+QYLkyf9tbhgnM6g7V5eS
lsBQreEJEPQPmT7lqsGz5iv2F38n/JhgdKbt4RTuM9sjdn1ocnLWkESM+oP5sSsk
6zAzF0qGuo/2ABGVQ+vc/iWQJiUuyW7AdDEkayyQo/rrOdZkEgPlXon43y9mbom+
gTJprdR29s/dAsAdTZQeU19M2zfp1sSf9bjfuiAguRflYf+tlbwje5kaenOZY468
4vihtSiwYoR9hwvbVBstwi9Cx1dW8jP4tviZgno09wsdWwAajLG4Qz+hrIAU5knC
CEmmVTnm87EoIAoP+Qo7Y9wT4NJ2auqi2gfN2Bq/cycHHk4M1lu7HjeOMc0STx0H
6OyoT0/KqVLNKWnP5RmTFvrRIqnFW+PHl2nGpfmF7HVr2Sl3dZQYMOv8ABhF2vFp
jR0MM0DsYuHJtc3ya7U/JKn2IRhR/OA1kNYqpWoLQj373VkmcEBqR9d0dpukPTUy
LUMXbhnGLnviEUxmLzLwFIu2niTi3sRW41Sdz7DvcOzQJutImMbhe7pJQDkEYdJ5
+dnDcDq6fH9smxRrURD4x5OpdCNXxf+xRwt0TEZm5uM9xO+JOHVqgBWntPFgISP2
jYWl8h5arc5WuaXC9HBqaNHllsoBPvz8/SvIyDTCdLqQI6cZMztjG4gzveNS7xcU
zlsLx6ePjThO/YK/7kPwaow95T4Fnb0xg8Ymgq8bfS8TysEHv1lntZghSKxaMoBI
7Xtn7yshJDDyDSizi8bMS/wADKIC9YngD85Qz7JYFjLAoJ1UuRdP+gGPsCZVnFpv
rDuhj5AjWak0Alr2XYiFc1aUKiBOMtSmPghoPbwU12Jj8IxV003iEbVzYAHXpuvm
Tt9KXLUkxzvXzsBbtvy0SFAa9/WpAewizUn6gWAfqe40djDqL2/6OM0edaCpBTn+
qB4diuwRw5xhAFJQJK9vbS4YJAw056JdFau/IGqqeoxn3DYZXh85hdAZfprmY0AY
P7Re1quyTe+3i0gLk+iNtyk/S/FE3A9Qki3QZBN1BtJMyPwY/ALqNb9CgfzuWnzG
gFX2au5kWceNFIgfLjCvP2pygArWIyEe9Tub7Gy8ASILaE30QhYf7fcMbZqrXYrD
GpofJKxfVjD1huyF5Ez7TwfZva16+cymyGQaYqdyTKeluHIj3epVp+iSWjEuc0bA
AlyAgGjLl9GLF9FMFF4Zb9vrvuG2IFVLVB1VpbR7ULQgRSdMPbY4wVidNfLJkS2K
ZurfWQqXDp9nKcnVo8kte6QiXlMp96GMA1h61loKbO3gNAk9gqPQkJ8oNeUQv8Mu
jfuPF8hEBNiOnDe8PB0+x0DoR5dogdx1WnM7WIm035V0S6g/aztVd//FPp1LNV9d
AnznJF+eFo4KkSqaucZyfzvUWuCg84kfFcyELsKPHi2gyZ8wbM5WhRBdx4EoZqKp
9bTBEwUrH2vwDqbWfeURDIL/vT0RpMoiF4H5Lyk4/cR16SF2ABws9IynH5LFNJ+z
eLlsh8ANg9cUFM7HTsrJkyGcYALmoiKp0eMLLCVdPIeJ0RabUwijBJ0nAQdFvso3
3lpG76yVbpFDdCkfJdeXGDb2xI6qpXtD/OVsK6bVyycUG5QYUbUZ/cPvW9S1N1RG
Utw0OujGZ6dzyPAFOq8PB9C/UC5+I8T8VyEMe0WB70bORXI2QpGI+ZHWlZa4njQI
58wDQFvV3xByASmYkC6EJP8OUzS/aziW3FUecCN2adRNHldKMic95fU4dzFDTOxq
DB4dNEhQ1oqsqR9jm5OCmfxXvywMzgMHpFC7BXhkeVLhJmEBNkpBdHRUbbTUgsqv
igfEGINRbh2XUBxWawmygh0HvJqD2PN7C/NBko07OEjLl6+u0i+fxeLon6VtoMRp
MVOboQYvL/Zzu7kkEuCyhzYkUq58AgnXPlSDgJBKBkVgg9D6+lBv5MGuiYIKOw+U
5An11NbQM3lXlc2ij4EJiYg0u8zj6+UGVQ9zvWyEGjyRw11Po8PZ5p0E6oiDCSF4
gCa25Zg/8HrPm+Kcgf4a4iRXHclUkhmeIbYo4vRE2+ERvRjoku0uGFIXsg9ZydvA
1rKJrL8Z9ApCH1dPA+Ik/NqTxQri7W+5+oR3IRR+lBhfXued8Z84MtSqQCgvqVx8
bxs2ZKv5AfNt8cKNKk3RNIz5hleXNOkkVayBHxzDeljt8PCIUxUMUjHm2FvOd8o9
+bG9zT6ySYN6LY61gz2KElooq/inz+ut3wk46zHXOmcbUiRWU2LCrtdn9+8005Ql
y50H8ryCcJx2/S/wktKIpPITuVmzdFZ3y57j5nCd7YjRKE45ZXPJNS7oRs4bqEUl
YmVnVehCqGcbRekzABnZTQMjnOdYEdIYFowaKwLC/T5/igh1a4uZfusQwOet9szC
ofRN8hgcTaQ5TQqp4F3xvcDiH0L/sMyUO0iz5rWtj80hRXhalh67TeSCoggikIek
rFGn5PWuzMwRSYd3NiB2fymu8X9CnVyqNGVwk8/2NTYp0qeX4XHQYqi9yrDV03gN
jkoqKPu07A/SMW64exBp62qcie2mU1xDVyfeF12o3vDtHvVww64hXPUw7sXtnQZn
4vF+liKzVGE3EE3XL4h9yHZ9RShP9pQ+ovg5K5h7c/FNGbysR5f6oRxwKsID9vh5
Mg4/5wV0zAztRDNiWzDc2ugPwcNYG//cd2bNV8hyX89a2O8Hq7x+wHNox1II9p9Y
3jDwkbcuY7jh9L4A578uO/mIhGUTy8Ei8wPjAKHhAkwfYCaCmjeyF5rZ49OhAIRp
y2iqPGU/h1UNayLw4Gp5qBrl49neKmWS1M6K8nZLWHzEObYdX62H63k4XfWho6mR
GIywWdeR+nax4iJhyipTogl4pfxkTmqbXCW5ct4b3KIHRlrVVE9Ke5EJLPzwceF4
pDDrViIuRVnxnzgKri6v0yj4x3QAezgd2rPhW0SmnTJtpet7CA9xmWX4o40WRjfS
r9H5EvaBE7sWxu8kR6zhl2UM5qrnbAaFbgPiwGcPGw6DjsLRmsy3ju3jyQN/RxZ8
klD1dgTLkIrg96fDzaJoykuLsKzTC2PQJAZo3R/NMsE43AeUPo8diq2i9E95mFcL
2qplx5nxThfVEPFoLPb5uFHkpoTo8av73VKyv6jWonIxSsr83UeSOkTxRgO/9FJH
P4n4OkgVU9Dqzja54BF8/ot6xCM2/5RJPLQ0wLXigcWVHTwj6RjwuMcU5UEChx0f
qy8OC5ki1IZBY02v9EUY12vj6GXw5n5rlbZtDNx6SZm8pFQIpD89pb/3tkhjgRsg
5aEoE8imOvSAiU6NO37c+MB8X+hxN8oPwLtjT3qsxhp7eCB2AiAtwfXXUSD2vdDg
lx9W3KryHtd5iKMyOokRO6ConXVi4qVVOYzvH7IZyjjfWoE9TCJSnHJkmfn2j/YV
l0/JiAVjpdFLOw9mAMbIIHW/8Yz9W83XCiTKeeYU4/ofhNmjjisuQshCcTKoojaL
BemkS+xsg8g45173EFyrE9rBEzgxgfD/CLUc24glWyxBhk7rgZKdZGZS0cwbz7xY
koTmDBFbAAbswbrvZkJ3t91np2S4DpJBrKUU+pS0+lUX+6/Jy+g+U6IO9LHlTG/4
qx13J+KL0QTemTaA11ymxN85TxuoxwAD4kq+a1Sp5GCzf5jdlPdRzmvc6Zmt279f
7BKlpQX3G2dnRszhsln4I+LKa1fdo7MB31Mp2+k43T09Ef1KUrUDFpL4kS/Ij5Ew
rksE3ImzhhGz3Vv8suEoGTK3QhvFMhvTLsQ0VnHso+EdB3aMHd3j1Hn9YQ/3X1ff
sdWgpnXta1KnhFea99cxSZeBAB3K5AnQMmi5VHd1ROKsZsUBV06XABF/0UTBibgK
V8IQa+Jrje/ROXyvmw9yMEgCfFOH+K+KA3It0LVD9TPxkvnI0DQ9o/zB4BuccHNl
vh6P1rCQTxAV4MzTX0LWm2EsAaULD4oeg9wQAKdpQNrGNsY1BQHZ0XGN/zx5FBN5
SNH83NiSPI7FAswDzqy5EhQAaXqO4mLGHGEeaofsTGbsIOGfjDIg/69RzhKnuDUM
DYQr2ooIuphyDJcsh4EGEzSZoZwGBLz7N9gCx8z/hqXTmcSflA8aA7JXA7AhemCk
4LPvghUB06YO7rC10tLbAOB5/l1juLRme5neFcJd6EIGskREYfmtlp6puL0UXnHY
6Ele6MbEtu75oHW3ZyR/jiPEepIRJ6k0hkfGtrSrqiEGIPiX7+K+C10GHX8Bq8gM
hqv5/vJDu45awtpnCvFZ912UL/qvbBpT+P5xXZU+gPflYxvU8QWGeDUFo4FqRQvL
HJDrApUrmi9nX9uXksoiiaEKvPgofevkI0HU0tqasoTkAwjBr628Zz6Wc1hbcf8M
TDarjnCY7PMVs73DCMnmRV1WcQC+MP/trTmmmpPZDsidcElIVgDLcP1HfG86G42o
9ToV3QRWmTkw1Tv/tW6pmHcopkjY8O2NZT2SWHL4V7e9gCHfAgv0rB8jPW+saBA0
3tj/hqa6rIvkaWX4kplu4jBGKGd+gWfz7tR16wjF0JoRrTd1UyaGBFrFGIAuYo9f
FiyZJRTlJJtsoS9EkCoPHfLWd6ti6iiB8LwJWV1dQPhUp6JjL1Nv7dP1mFkb7Ydo
HAMBbFrQtb9j7vukTwRjN1m9wOm17KDK/pguf0VmMrGXl502nywwwN4pojPMQ9kZ
L84N1SqfeTAO2W/gd8un0qyDA3eZtbjuUs7nGb28mcPgPlmDcLtzuxsmYJcG/Q9p
PLdBlmTKoxDtfDoEvalybRZrGfoqqcA/QLHKeNfHc0WbwtOt5J27r4BQE0VubTib
50wpfybKniQxPvMSTTFUaUpNaX7rRcTuYGQlairbcta61TFPspqiBRktsL/r3ERH
ns5UHbX43zfS5h0YOrJh7rUy9XwP9T90OmOv8sgWmOg5jKPS6A4A/HUGXMD2xPy/
TAdRnZLuQy6UY8kBDM34n8+IAw9tqutbb+/jttbAXoT19lLgpjZnMp0MPtlFce4h
wNRfp2NLLbEGkD19Sut+y/jG8/4wxluV2WlyL3LsTm05IPjSMXPkmCnpcEN9AcTa
ArdpVyU0hnBM08V6a19G25zH7hGFKMYDxZAP+wkwI91qzOPCRzh0kW1oup5fvoDt
duSLnGRg3kp2tFsJqwgFoG8u0KYYRYlYzwwscNeUhiigQtV/Np3mMOyv3Qlus3lt
GTFvgVNIde0/VCU4+zp19iXPnR0o53Kt1GQ/7X8J+7NLW0pMibSgG1UQotQcbIQr
g0TtgQQqSTDs4NtYh69m45PeluLgiLRIrylOUSaZnkGwWWbR0Gyt9ohBxrU9IH/5
eq0fQkxC+o4T1+SMl0QGnGrnXCUjcbvZ6LnpuBhDxo6DSIWkKs7egNaIbS+zDzpl
jDET1vU3xanEFrz1jsPwVgCDw0p4qeCzIsaRrwHiey7Xvi+OnID3cPa1tOYCjh9q
V8jnpM9IVNAFsMfef4Cv2lIp/gyyCiE+E6hN2xn//sItt6ZFyEgcYGlQtmbOtmM6
nu2MKekJYjX291CMXLGkJUuUXU0hT38vhRY2QnkGXJbNrX90vQSGl0wTdrzOHaeQ
EgWyK/XhhR0YSmGfkufy1zHCVOnlpQugrzsADRVS4p0lmBKY1BtQVG/Q9MzPFzfL
ysCVjzNoN+9Wn8K/bxwH8YTQk2dUYyObRhDUVXoJw2Ohe+RqCH/Jxs3SkkocXm9m
P1cyRIk7cqFacOoNgdw9U/4z2cYNhK7igQpVMkP0pwcNRZeuwyQBI3AyaY4E9NLL
GjBi8xgkkFni5+XMPf5n4xnusocZx3SNMUM0ebeyXHuIbL3r+9uj+lHFDQPlOFuh
En7exjv8O7r/8prpdS2Wg05rwT9sd+4gZRTw1tAmwQX6amhlLnd5irDiB53qjLfo
MWLPoZbw6PzchrgMD9vySffgsx1i4Hw4BvLRjdRQwJQyeiiaV/4behZ8fEe4xVgK
uN7Aph4cmLmfeMRrzp6TOzpnYUoXAy7dRNjX1RGJKFzlk44yON+bBCaw009DJC0k
Nh3RvwUTbgKRfkpv+2eiiHpbrOywVClZY3LIBVY0vu1P4wA3EWERxS/qcm8c7z79
szP07yZKXzCEhDSZfOC1MFm+10BB2HsuCuvxlr/+5lEYQe5VubRvH21RRmqXIXmT
ui5yV8ceXTLx+koay1aNvdje0/Q6Ibhp6+eMM/14wjmvmPab4nXLjednoA6W0IAX
E2qT+OvkFEJOlJGfYaTDZ6w++5Wk+oPRrJ/SDKNesH0lDcx0E8zYOUrorcU28U0g
v8V7TuWLV9FjhHZVz4y4qk/M8RpdHhv8HQ1RrmBIDc83bR96xV4u6Xxk6l3BchBu
ZhCX3NmB8ArJKq0eUluXP1+LYKECT9l7+O36Yugqa+orMA8+ClCq8bL9A2eM25Rb
V9YfneGHlWx9Cmj65cTv1W0t+Nta58HU+yQ333XCb5ck6JebsgoI5DvbDCW91pBS
yYHlykc2WeaHTChHxFOmhxtMcaSVQE0VGBVew5Q6+aIYnsccg1YKp2wv9f8j/kaO
txEKyPbe99ndsaGF6puVH6p5gHOhvBJOykMB0ZTSPgwyNye1aWXnIbVFyVjjipDu
fbWuyJPrFFBdGr2YQ5Vpfk9HNFi4zT5XjYOGoneXU4HDJcmKreaZeMh63HbEvmgu
D2L4UtlRx36bdN/LvAX0GgNd6isb1mOhLBd4qbPlYlNzyc2X1rX2RX5Ylg0nCE+E
ZbRlJ2c8ZE6C6JjHMhjrE7t4rA6Yl9THVrlbRwlbEcMo/6eT5gSUFvUdYaJGsFcy
/Zk3jYUwrKdtzj7043X7uxuVcVTNpBvo5FFODJw9iMCS+BIjDaAYo1Lf02S/W1q5
glv3t2GTKgQE7PdGxTJQM2ke2EEJ6bGL8qz7dBryouKZBG4DcLb7MfrzJ77VqCAL
7MoOrEPHBi9iofYTQcke/OHTZfrjdiE97pwyZeReiyeJWnER214bA+c2F9l+S0Fv
Qv8Vv1d5VfLrj4KEpCqLR03KYctRLh3lyIBsXUNUlBdjpmVzzZTa3aXhw8mjthuv
a5i+LiaDiFRvINs82tLJKMOtwT51CQoR84wNt7GQABG63pZxowq33XIgHUhkGhGr
I2EYHcsh0CEVZZvQtkntJrfgtUZSZm6DCpdkZ7YQtj/Aaw7x0uRBCDsjNSGjtx+t
1BrwGM+Qc+DK6Xq78t+aZJczgFDq5/eM78kUM9a4MzR5XmKQuoZKZiVwmPoC5saB
FIqINzIZqjMCScPJgc5NsxtEDr70Bfi0ZIlR724BqNkm1heYbLg/64reUNXmTsAz
snpq27ikg2kv/GGDCMTPOgOvvKA6ivSAKV0ewkRwI+Q/OKNksCZYepYvFGrmtE33
gRQz8C9p4aDRHnAzryH+SypsHaGhjYL5V6QXCzHzQIpO3WpoFx7NnW5IDKs1jgDQ
oR+dLlEJfct9nrUnChLGWCg8VCs8a434nazkK2/Bz5nxDrwMg+8mf2kq8L5bf9yk
l0j33W9+OD+Ti45GdBrp8ofdtm6n/tUDdT14VPTZ1p8zxHxi/OoztYklslIHe88+
IJk6usXrXH9cJLD46H3pSfiJYvCZoOITzVJtQ/Rs9aqdfNFtwReazNZq9RhCHHII
IJxmLLq400va6AlSl7kilDHZ8dLTlsnIYidC5Bn//lZcEKvj5auGtJ+pY/XjLmKb
JXs4ykMBqfG3aTptmtT8B/NuwBdgqMayJMJXzyNU/LX9lVt1rqpq6iyAzmDAQWoj
qPNV7Ojue7EjyHeS7tCUNSyUhH8mtgFlRF8rQ3FQVhjwjuxN+SE3L9GYTw2ygXpr
ZLE3tgr+8ytP4PRvBxUlTIcqM5qZ8ZugDd2k7mhmXQbTJ9N7fwms8jixnHOG7R7C
o+PWtwPFYPIk1ebIOdxbz5iI+ZCA24wGyEJpOLiDu0XZ+PupS6lvnTaPrV3anxXc
sjm6WBqjAepJOy1+s4AMje4m0+5J/3IAmv3LzRGusRRlnSbsXAe+ERUh2wyVuCG4
L88vZ0th+EaXCl17spcokAAIIVPhRXsh7DFGbbYLxzIXfRPdJbwu/BBkFLe1zyUJ
T/woyBtzQPYSrUNR/Of8QETY+VwfyEyd0ZgEsGEtJz9Fl4dOyba1T/Jq4ePS6Dje
yMTbrDhGeECZl2eb2KaxUEemyVsmzPJmcmeFpQK5HqvhXaV2uneFQRR13q1qtFR9
+NbqwRC83uj1sVnglY8mmpXedZ+0LQ/1f2WoEBOBQl5MlD9746lAwg0CSbeKQTLq
BmHu6GRv8xCyDhzqNvMtV3ZDnccGmA9Uc8TtBu1nfG177kaLTpdYNeRqz4sHAa8w
Ce/ur62N2Id8gDhrz6hio6mTZxwVQncjRuRbFMAXsG3kT8n3is6nMIc36VEhhSTd
HncVpkA3OMc1X5S+Z4+gpl2RRqDy3St4QPkc22ctoDvcHGBH94B0/xC2SKPX3Qj5
/+Uy1nEMzFPnWB8fx/7T//EeAUMBqtElBd7jE5CqqM7eubpafQq0WREc7Goszcap
dlSL4hzJ6N1cNLhfFYGrOU4kZj2LwXWFPPXEC7yI9+WRODu1em/R/AHI6t2UTgOx
ji+JyBdpEXWo6mbHCyW0oyzu/YgeoDTHJ2DMrKqVH1OblOLS5xcT6Y09oj6Leyub
5vmcLRKTAbzwKnmua91PW9roQeI1zSB3dJ4OgiKgY9wBExl+akVWEAUMn6jqoDge
skh7WedNBh5aNzcXhtG3Lbv4p387xatnRCFpWx1nXAHH559bTlMDwEuSH9QsgQ13
Xm+jeLLFpHpnaq+hKNy2pEP8XvQ6TYdVohyg7mlEVaj79W1jQ04SuGYVjkOvGj2J
XsgN/RccM0WeD/MsaKfKWQZLe+d+SdS0f80UPX3eyXoV+JpgnxpsI2PrmA0lVS/K
VtsmiSYHTg/Hdy3rbDT6EnibMisDY0XdWynKbwQGDUiIik760eo9KsSrOaqdnZrR
+HH4LrWjJwR6FhoYigSYPO3GvGji28nER1olrZNvyuvOHnvXGlE4Y/2gP+Kj3aqe
ULh9mj0VU0IfaAB5eK79qIDD+J/6JHAjP5QhMw/VFHLDeV9ohZfbwvWxJGvjbCBy
AASvExRWa5d0VtdhzJUlEawBxicDFSI5DGk/gjXiyEmv1EgZjBB7tjqyTOXtGHPj
NCwO1NdTK9NdL2TOf2Z782puENUaLFGJnJu8jMUTB+GWdv8SEwccmqSF8lBmGlXo
G6x398YyHnNoQvsHvzcT3GLpY4aVaH+GpGXsKZu6h0AOECYjSm6Lft44Gk/G6eBv
9C5qB4RLUCnkKPisZVfuaiUcqvOUFnLRIIf+zncGiLgl//z5+joKdX9FAfOKeCIe
8ujdpJtwtkLoyZ3cy5ADuZZ0niWFQC0VRuOQzrXBj30t0EJrn4H1iDd/OVsBHo1k
pTOU1kqCP6iOlDJcmR1kXTIkMcSAgAGYgBLoWA11jF/UzzpVA/9qpnzIY07FVNkE
UEGhMFlV1wYUJkex2Rcxm5aSNcLgljLj73mGF0NUi7RleqJ8T84BCAScEE5/M+u/
pIL+WBtOP7wQlK+9UuwY1ruw+YlbMfZnTB+Ej1QUnOEYqfMLtv2Qyg3F1E4dlDxx
aElEo1EqqQO6BTQth44Bg8mhf9aKzKflXxbNWDMxXoS+2xCjK0WW+80waps3Vs1E
fgH5NDqBFqDKyxD9kWYaaIfjUwev4tZKaNCCGJfOfMlU61awWA8fTwYJLLdxOpyT
OEQ5oDYyShRxZ/jsHgB7SfZZCtb0zsfRryzi5UuvHVTe72XTRqoOH+6Og34GXv+e
qgwmTBDGPUtlcEuicb+/CpK/+NS0vgAzrnLQ5tHLkcziEOoYxDRnoRpcN9aPT5LH
WB73JNRT4744MC13/oo8bsdWPXfEYJw1lvwX5v5+WqeGli1JBsJejuVmmOiI7dFx
Qt4IlFLbMTVs5hi0F69Ft/B0vRGrHTosLYcLLqwCZa9403ph45DT8fT++OI57SKr
GM1ahdhxj4KKOpz5Cd7Lily0nQy76PDDQqkmk2q4/19JvOebT0/GS1p+PZzsbFv0
U53srIHE5Uvx8QEPx7mu7Gf+coJd2xO+d3CWSv68/vnB4RZmx2C15Y5MscVx2Krz
qdlpJ+v5H8mT1Zl9tca0JoaU7udBLqCMe9LQo7VaE29xYJMySb5hq5iGLHXkcDqj
IMNIWsxFPEeZqyPTvncYkZSjFVb8Qvr5MDEqfbXAZoyjuz6O7np4HCeKMfKqeVhp
ECCmVoxyTsffLB3zgrxixaKR3AkVhFTaz2+tXIcWZXAyTyN48IBjyj5oe3yGFsXG
jJ9unKYcKcOy2XUtxpFJTmkwIEvGxrSfwdxo9BPDyuTzDsQbZ2LZaJPiOWDbvlrf
JGjdM6T4+CBP7il42Ppmw3hjnOZGQkSNpWmwrpTclvnVJyhHG2l+83sI47hHnoPm
7SpVbQ+ufl3TOYLvk39KjTPJpnhg06T4QaRJzsJkEyLZTWzB0vNw1AirBeYqSSfs
Ruxeoj1f6mmO5QLSWioMKXOLQDa82azAKMb9qZI0sqFKydcP5qNjdWcEpMLJx/IG
Zxw71ryb8A70OCRKwEPuKXWqpqj22UMtrlmnlYYaMtAzHJLkrJ8MiKwIuDLNnxfQ
OJwGAIG1UHCXpcXdncKzIf7OZ88vGxDcSIsaQHy5Yv/RnHT+aUbXEyX5Q23BVshY
e5FyCqX1bGhqRA99SNwj4Ui8Cr1XPL8ADWjrC3ZPlzs9dWeqLLQ6anWO0jbHdY4h
Wc35R7fTVnVfsxNcezAnD2RnWGmkdyqR8GrwBnP+EP7nHNbticEnf5MnV5wIJ5wE
C5CH9szlbJ8KoMhk6jsByxny94DvfQa0tonTS4luAqW91uBD5yydgSM8NCqeA9xq
Vn9FBH2cS3EX9eYIG1NAHo8fZOqAoXL7/YCu8tCqiNdkMzYNz2Q/toTSdfLuIOWN
/dvqhhPadeB06IpX7hDaB31AafGRVIDPZpa40n2BNc+Olqf612m6Fvs0ZPvtol3k
bEDPjOy/ggrJZf15vfi62ALE15evnQb+Qm53xuoadx2Zso8zMP/cZMXRpdLGZdsT
Bypk8Azaf7/XwZ7boIn6ngOkZNE04ZWKYo4Myz+lIpdM3qxPnDmdHoxY5ZA/kM+y
SOqcT5Spw55Tcv32OgZpdi1dQnppNUzO0XCiw+v8vsH25cqKg5tl0fGpDVA9LVVJ
bIMThiElN93S8due+YoAQd0/dyslw5XCZl02FJGuJbHZi6MdBjfAJE1mcvHpMCmU
SgN4Z+DgkOvXvYoSWOS4o3HZw/5T3CqL4z4yfAjIe81gewdEGJzolqvOUjvnueaF
drINm4Y0mfWvuc8tTYSzFcWsZkfJZm1xoNdaLok2sdwdVQ9GZFcdryagkLpM/Igy
NrP8g1PPqSB5+Y52H+adBiyRJ4+eEXWI5vse2X0XQyxDdPU2EzX7B7x5Xn86P+xz
SjqVBbOVbm8y4jAm4xktBGf/kqY+HnDqOWysSp+Wr3+nk43DWscKTQC3K/bTtajt
CWwNc9Da6A9imzPFY/n/nhcfjHEq3haBG37Zd8okSmvEBGIN7Ccp5yGokqoG+vEH
0fJ+k0kd1fFoQ9SD8cVDUDT5gRL7ZZEKMjbDy/O2cA6/7tAOoZAR2sd1TEUA0qU+
surs8fFDRdh16dlNejKE/1iIFGc6sS5gTnVf/37N2eKRgs/WwZ/F+yKHr+FFZJNC
wyIs13efCZq2sCe5AWkrIftaXZ79S/XNXtLnLqdS0W12U4OGdHpZ1xOi0FALrxHF
RRgom0SxYFfc5IrOdEeU8CzC5lDqkd1Dn3E1piqymLxlqnT3MCbEWUuPbrXn9klQ
orkKtVnPH6t75CEXVu81530yJ6PIno1b8u/bvzRuZ7P/0oltEDCIwKKGAmmdTwyx
arw4tkB+fpkLk5qo2AVaIBY5LTAmBcxc/pxxxU/CA/SsWcVlWtYp0QNRXRaxJMDE
ZkViEmvapL0UEvTLpsgwt1V/0k5jUf1KWi7DcgP8xkCQCz52fFY7+GOXsrXFHuC7
YOyYOfMvL8NlxL6797541VcSA0LLFWhvSghTZbg5/wJ3Y21Sr0EI1y30rpMqk0+i
z6ibb+oW1ZOu3FvnWKWvIggqeds17QSW4+MT+GuinX6X7tBm0NTHDrmY2gabk3Gc
dNA/qf9hbLXyQvbxNHtHgrdMbag7T+aW0sSLGphB92sdcrXvORZzTSp73Yhc8gmJ
lO6Vvc1YyuX/s4yTfZkRo4fln1NMVLDsTwGt/GioW74QrNn2hjRrtQ9X5L6I04ZL
VWoIaXQNjTOro9CCFDbp7/MuUDQumdtPiP4eeXQxkoNUd1VIe4r2zZP5aYPu0ZHE
KwnDIHCE0OrwoXTmLARS30VJsHpV5X0Pd9Hh638EyvhbHTbwCenaVKVkecoOTLdI
GBkTv7oZdx8PG+bHY54/OBKrlTkbYy41WngFK6UAoAheZhFrqsv8YWuruaeV/3ag
Ab1LWjMCpoUrTde6whaHSFnZH+lwMfxaCqZmTv1atpQNrLmvsa1ad+1Vfx/qo25q
eXfJ0GrxAyJ06D9n2j9fLsP+mz0g02GTWEFe+16gLCMxPg0a18ozbBSAbvYvTvPA
sOfkgKw1rxL5DwvjtyInWyil4WEfM8x/JnjNthvM4vwFcDjAhQfnRiKXffizTqgm
vzKlXSh1eOJvGTSRYX7Cya2tZ4PL/alF45hC9Ie267CDDTjURlAMnKkFWbAqZNua
zWA7cn7K6wV17anjZ36MCDYwfa5JpW7EUczIVIUCHKpRGpbUtwvF4zdxZGz4dUyY
5kSzVe7tOQzHuvdZ/CRqAgFR2VcXiV3ue/VnLFPPfOz0fV0Jcsl9uV42f8UOQCpH
CjQlb73xcpFKIsm4LbmF2nelQzIZinmFOU/nNU6dPRp3RBhSOJTCtop31EaxzrSe
5kuh4hudxcHrm4j4EZxiladhvLc8Ts3C2swULsd0QgIltIhBnwVM29UJ2bh2c7G8
E3ylal1Z6G4KkgnVlDnbpatsHm8O8HWzvNumrtbx/zKUS8yaoNFIywVnyWV++KLT
RLNANxFV5OLYr/JVZk0sorTsFhsw4QtB8kVwvTRF4uob3DJMrJQV0VL1Swso0Zru
8aJglDVmNjWh26TPmRhjeNIhQHzeaOQ81mLMGqv00nnRA6EAxkMvL5LSHmh5HTnK
UoYmWnUfKRvTLjx9pFAyqlr67AT7/KFWMkHIYTwTK2cQfoP5vb9bruyIepSZ4ucf
ppKoKsQe91O0EI0qGcadUZh41xXH27i0clY5xqF/RRog8dgptJcndrrq+YQ23u04
KIoq3dPLQhwvIaHT/JHuI9yXFWYaqiRqBKFuTcYdF8ZiAEXfcjarsLwLDnyDqmhv
U1lt5YMllW7P0LEduscPCpQsC3lUTBiIZOpvpl9UbaKyooTosEuOuvp2d/aDTx83
50QQVVCd8KPKW0opLLLDYDRjr66Ic1QqoaQ3y9KU/OCiZDE3aiyNVRbBUv/qGHb6
7/NrFY7uW1499uG4VzQALmlqL8ztHNUVFC56P2J/d0rKwipcn9zsmyd1/0xqh2O3
IZVow6hc2RYXJaKi2/jcnvSdoTSDx9qCfe3rYJxt9dYv6ce+n3Hnf5QltrU2BPsq
qAaax7RbgFB71K1QzLOz+WU3/2RM21tZIASlQ2tH2CHVg1auKnLCgUPGZJD5c4kX
Uw8s3q8u7ELr5iCCjZlR35cIfcTdcR64boPSkH35+IBeN+kFf3WPGPjl30cn+YJh
yRdxgtX6vxRatJvt5E5piNS8zrRN0zckLm/zz/pibdMeGMC3hMcTz98SOBXNKjxQ
0vydBBpSDEuWblPpVm5D2L2F/Lg7CuFdscP05vE2FB5RQ7rks8QrzR3+YFAknoK3
VmJ4aZsW2/i4OShU0wL2dV3K+fam9dyQ+8yNGPaLOoISOt/JJM+vt/GoAnxY6BdU
YUxyRimik3zHPre4y1no5iiW9DRVkF5gJ8Bs2zhC06olldkftM43pjX69sFOF2J/
/GG4oDl4OKsToItAJvlWdiPj35Gb0GxGY5xst13ar1QQTk6+WTEEf/ZJWVFUm1fv
/RNDdi1a4BqUMUe2xdqVe6XXE22tSDxBK6yspgThzD60ZlSc0Dw/FiamcqIqln9H
8TOg76uUf5nKcE40WLmYI8TicLKmVCgkxFwDjBgugrWs0nemzLzNHXzPFbqXjuif
cj5i7uDVuzc8hKuMA3zru4wjf5ONelt1WZ5jLkOH0EOpldV1n5sM82Gb7MBEmAyP
54L6+GsTQostWy5Ru69V4Al8lFSWZ2WCuWn0DjKzgT/77bz/78FQijWbpi4MupQ4
WQxyNbSnOEbx4gVua50xZ/t4MTMkoC8kgrj10liHDiGgQMQ0hYRYrtPDDKRUpn4R
sOIUq4emzCl5qNX/lCuoqjjfSpeR+LeiBJgX5W+5+AZY7bq7PZgCFC4UKHqkPDJJ
q2hzfmsU39i9ZSlqw4jkWOXjHn3U/MdL3UzrWeLjQhdF4HnGKCBD/ZqhupcZ+pvJ
YkeOXZIfS3hbxBGNFIB7xhNmyp/8NG9pkoDNoHU4B4NmthHakOrsqRiJqdJvgkKW
XYu1hIzRInb6Nt+x7/7uvSWySn4Nk0nXJeEStBtZ479jK9fE/EqvV1X9g9ruqTOK
M7BsEL/7q0L5B8y3LdaQP/1XSV7pX2A60CVwciAYFpgPiySErUcTKzTuaMudpgS5
3CpEKPrpGHiBs6J3J/Pkro31iorUahfMc2Q9ywa/oK76GNwh6EL5mfqH8P3QywFj
H62Ryk981rOnyjuf85vjMrXKMgYnXnDEx9VpjKoj4YdE45D8sOrzM5Ci+9xoCP3r
dQ+VPaE4M38x3CZRITTX0HhPK6VGqHEVvkrxXAAmRr71/ebCTFntwA4v8sTxzLeQ
cggN2ZnKBCYFtSPhPbZbYQDmuAXWSx2lQJwPWPF3Wq8gfU40/rMAmknXl9EUiQ/O
TAJkdt5Q1uRHCzPGR8cJemX0+rkQYMLQVsRWmYtGaVPx7pXI5DWk5rzj3WaR5T3m
zm23Yn3zzqv7MGiHYe4UTXsgJzxuBawOKbz7FhQ2Pab6RDDMRcZHo7szjqgmfQ2H
uqojg7rme9mq8qb6r6dihxlg/vNRgP84jsFHhTtdSv32uR2cpgze0WcwBczIsMpw
qxJkOeoEisnCg0jXtHkeCsXnzIC0Nh05e1KxkQHNOOU6EAE/PJ++pmh8gVXFe/3n
lu6YXjpvo+VR9x7UEhxFphLMz4jTyMw+UOdC5jiekUH+1SxWPGJS5bUR3cXVJrSm
20/v2NcYINGFeN/2s1VsoIHroQi1nWahupb7IJUw6p723V4QMddcArxYO3uP+k9i
yC4mrqcCYa1tD4jNoQAVFo2nF1+4JgrTNbf50inMeqiitwihp8tIB8LmZvBXFKf/
VRtySCByWEohWzhAUbyvwhq2xje5PhiD/KthrkEwHbEG/HuVKEuPUfnBN5MwKfgA
RdHbqDJ4Q9bNtmLCfyHeILAm5vlbnUVmihTDLKPU2JouY0AWA/UjcL8/vBZ1aKEc
SzEdH/RXhqLZk3YCYlsZNCg382WmxCyIMb16flojFRAeBd5mUY/f30/g4Jea1jNP
QfamxRzVeOrYCAa6qia1Mb7una9ahPAq/IE3eb2RFOo7KjoyAt0CNpUmZhQ9sb+w
QsaxftRLCLmnThrEQTRGqf4px3gg30/SdKnm2GFzwug3PdQeYPIHfYQVdArbEOTI
65iQBAsBGRDNE9KiqsUj/G5P7kD8FNXsbShxmPBNi+tAJjz6rllNg7J4Z0jU9+jc
yezxmpRqwa/4kWYovNeK0iGwYa5oEiR39eBqeEkPIghyGWLqbnVpvQzI5QRhYVD0
9JQmTOf7CVIL4EkwmwgvTjYBJ/G+9nzvsYtdqkgKgqzY4bKcbPLNgCu9LydRZY80
rrVUsb9cJlyoM2Bdb7ggY7J44nmZ6reAa2nVy4U+rQQqEZDthHmuwFLzIWwcMwzD
ZiLXvEcikCsDuaLf2TD2tk7g9ydWzAttJNrn5z8oc2cXEbsslrgd70ZZGHmlu1Op
kFBVNHKJTQH35TpVAx+K+d3SWyKemwrbZzuMVxwSbQSsWX7TGL7X8Mi22QzunvvU
cM7icukLGQoYY1Tlp47bdmzwdo9+N+nonVyR34h3cgepontBmmRQeJZtThwA9sM4
4Ki1aWdeOsynYVvynorV1jAQt09ml6Y/+b4ieebQ7oTB/seCN2FyYZSzUIj8mA/L
WR91mFoUNSvCIHoVvfwVfXcmwQYl6iHUco0dPUF7IMZsq9ucpbh9Dx8OCqu6DNOZ
pVQcGBObO3au+G+9bdiQaRk4c/bql5PDsYYeR2DzmgqEVq5WHz8ooJVAOPWzlQdX
UFFAPoo/UCpO9QaVNTJReBMyj7FnM9hhebzXcuq+LOdnWH73Lo0dak2empux1ES5
Nq+yuycnSgN0xntWqdaQNwSmYiSVoh3SAJm3nrZNElS2dwZtlBwli6hqLb0paeQp
g/yBBk7z8Uf70Alz/dveAb25FFirMAzgnRDeZwlBy1PHkFvl0BUl9m/0BfCaZCh9
x25Pbwvh7KtYnR6FwUTD3YcGnTBzuFByhgI7fmWxpNxcyJL8OmEmX/PGFry+3bJt
exID2Hh6i8cZe6c/Lh7ET0i9b0lPWbNjR0i9b8H8xo5DPDoHnUFwCU0aG17qobsM
hH3R0EJIE2SjuvcFjr7N5OiRR1EJJmx0N7NEWUo9PSWNybQE7rB7c2OTBR3IaLjS
YKIEfbFcLAUr2dAELiwr+eqNthhqNOIpbc1ESQ23jBMeNkrs2ynfwNXym6TRlcEh
ScS2+OsD1BqB/PC/RdRTuO7sx8RfNhrNvszkIQHaqkXu43Hopffa72BTprG5Q9J6
d1mWpcQWMPlDblKvBk8kPGoNlhG64V7DzX3EPLZbE/35oUvPgWQ8dw9F2pv0lDZQ
ZCXQLRUrTvNRNQqFMxcy4kLLe/Xtr1pgApQzMLxle3JwPOX9zRjYavCJNR4hyP+u
+AQFuRfsDI1QOjK+vkIhadrWWaxYbF7qi8tD7oAB4F8NJNRO+bd5cps0TjkA+41j
kTQtYi7XhlEd1GcKYR5uuub0ZXoFoD4MFDXycU2Ri99F9Oj4jpjY+qw8u4sL/Zpx
GjH+XnG+h6D5nqTu/ZqKRpe9smFpLYA4N0R3A5A3+/MgM+uVQ+O6wZW6U0Kzv17V
iPefYNdiHihiS6/0irGViRt1/hX/rHwojmJzB9GRDyu/8jrdC5HmBIt9HA570bGJ
+ylZkPOTDWF6iI2deID5uN6x1cjH+xSv58tdq2hRH3ntvClM0J82Viv4jf+7wAki
oFeAo5ZF/cDVsO6RJ2pzNae6jNktO2k+Y1kBCDLQsHzV/vY8FvEB2RWVm41SqMBR
Cfv2GZ2LchMsEFBOERF+u86Kw5dR7iLEb+41/FvC139+gy+4ggbZY973rtuaIjIQ
AlLxT1g666NxpY+NkD6+vvxLF+7LXBE0cobfBIqX2F/8AHZq5hVhU4qdcs7+nJGi
5PefE+6j+MurBwouMnNmZb6VmTQpspG6vDLooewcr9kMvcRgH8/xrT/4VECzodaK
jJlOvMdp00gAB7BMD8LqPb4/oDpGq0jH7ooe7nDay7VeVvEb1w/eHbn6Jmhu/EX9
pee9RP0fDEncHzcTTkjHjcpk6bz6yv55wPhHuGrjFlAxi3rk3TSQjhIgbmuasPkm
SxToc3MlVc82A+bgRFoWCoq/osP7FQQR6d/Sy18zmLUOiNCoihcHFdHU1yrh+erW
anJJM2kDlf4IQKociy0VPKYK+j2w7fIVGMxPHrTcZ584fe3DDROlXwcvIkdZ+pXo
5jn91JECctLHNxdooyw5vnEJvDMD8nMzKk7CGVL/J+cL/9iMwuC5YpVcK1CLCNi5
/Ac3OWdrMr2jVSY2rnyYRewlEwE5pZn0EnGmtVSNbKx8FsNP4haAMfYl/bcOOC76
O1gLk6/wM/M0Wxzlg2HkenY16al80pFr7L63DIQGiZoQ/U92RyOtD6ms9/PHAh6U
jcJ+m1lI9gLPbXskh0INijVRCNNyHUuy+fV07Jz9ep4ut/xz6IxoJHJwTFciXYdi
ZwyB8Tplv9rSY59BWe1Lkhvz39KAHy/xk/TSZQgXJm/1/SG1CE3+WacuPTy/KZwj
vM5+F+4diQr1hSq2qyvG5nHWi+w1OnOyke1unfY0s28/l4dRxHG5Yv4kluZWurfp
o+kvRROQq3Q0piSVlsEggvNBfICghgbiGQ09cPjpWUZXaLmkKUM+LOLqTPRD5THO
RuK+0W7+DtA2Sqm8ymbbCZnpVVhuh1Y2SMk92f74zr3pZu2cmnBB8xGc0safWEsJ
1I1S1tuLl9TwWpGok2JZc9vlE8QzWMeKjQHsGqll8M3AFvfQ4iEBno07rJM+v9Ms
sgkzVEgYkntEoz4Y5Zhq128NYqT3hbQEbdAHq6ZpAvL7cQZY58l9KR46Hd7gaCNv
NfhfSzJi7f/BA73c35UJULoOwU+vpYkxp7h2UJgfLdN67YVLQ5RmzCGZGBksCXVF
NK/BAuYDvvACDm+vBmXRqMg7GtgvEp5JC8vDehDS68+xLQTNc5rzk5A2ZrWgia+M
ViO9dB4ehDniwNF/TNoOQ3RV0XTiCpSy3C9gxBmtnCQ9rYwSRTi7RZjDO/35HgIN
XU149PnZsp+DisSeIp9WEwvsAOFfQoevM2wTMveJ5YhGTGUvHg7dzK04FwoU13tg
IjF9YBPC9IOZ3zguV4buel4m6+El0LiujT/+PdLdEwRnup3ARuxBJwmp2k5vmnwp
S/7HXw0p0DInNYUdWIHq1/UaaTGMOi/xEd2QDKYDKnc1VNdPD7IvLOQUw49mfA5u
NjQyMdnMGTUYwhr3/B3VjMdqhwCE7gGbGRb8R1aRQk/Kb0LUXA1Pgm7p9KX/+dND
zeKIxmBSBRnpUb5aILbbQZwWgJrW+rtHqREGSmQwngmJGRQBASE2oNCunoX43tCq
0ilS81fo9ao17C0Oi5pTvG5vKCcUCmX72DKRSQdsnVU8RUYsUsyH+jUudW5+vWlp
g1bcfARQs4xLz8SwiadXzHmyjoVmCCWb+R4U/DKl/C890AOXSIDyJvsnSsB9BPOM
//vj9kIhClgW9MfY3TmwvROYJw9kDegot/AiZjv6DMzD2jm54hmpfrzvuHwLTIje
uF8nUFPkfCwPT0FdixcAhLnztn8kbINwY/+XWhk9Lt7O2Ds5Zsfg7sQika5hy7pe
uVu0jmOeqsbK2XueeYKzPAsQdXZ3GIMc7u7GBp2FHaFVlz9xxTZELx5rPFFt4Y8H
piULZboiptftK25FUaRWKXxZa19CLR+PvTCDnUKpD6+JYWielWuEO6Fs3HVwuNPn
k0T91GWIO0YLI1keMvIpMQCbuuqLceiW5mlRCzmn6HftS4kCn/Rji2Wsmxuo5BEn
YGAnXyAoRERzknvS8WjQkbvYV9d9FYTICQYFhwEnRQRz18vReDGcAohT5ZuhptcC
+i2VkvX7HCA+TT1KzMWzp0Do7djFHiMS8BjMPA8+hOdB1KqDsQNq1h1tCEdRay1K
/jdSqG82XRrRyH1h8AnCF6nz5/68lmtD3D0dktSwoJXp7UNaXoGGOon+osPZU5bz
rhbxOESC/k82ZJhxcwl3Txvkg7JMbnqgfhjXHUq1GSBDiZLv/UElofAaBrBmxDLP
IBiU59k61lxcPz/FN7xbLvCMoIucy4QbvO3ht4fYhxVKRD1nWjk5Cqtb05Z0ft38
NgGeVbEVCQZM733fuhWcSbr8gPEh+EGUKXg22oFaWoAENka1EGeq6gU3q973umgX
JPzLN8sESVCjJHfE8CMNBZ/XD5XeqwagoHH0HRL8yWuhMeCeFR1e6cam4vn2XXyS
JeYG4bk1if3yCETN29FVkVIsc7S4j4PK6bmIWZmTMhcyGTHvMivpf0a+RCooxwlb
3/zO8bqAJAb/yzowArWnsFlqVxlK10j4AyQ8hhjnjbgMO1qQ+NN70SjPevthp2Af
vJFlg+UUgHaZYlifCDYMgRBZEo1TzKzoMaxQFBghNHjIsD1Gbv2N/Si+xDPTa7df
aKHExCDMrFp1cA1F2xW2KRE2GS4CUwpdppIQjKjlaAMdu/QddUdrBYYyvsrqzh+Y
rc6qIIgQop17DtXOuoxcnkbDB42how6qcbpyTeX3JlFXpuZchtz8/5s7BIAx7J6E
e9UA+uagn76CAZftUy04nnAs7ZfqHcjCV9xN9TUY/J5stV791oyNDlvQ4PCIr0eW
siVR5nOkaCPEL6wO+sNLKJhauls/ccO9/vHx21H75nGGd72tRd971p7KiTqrutN7
CvWBX6ybxYLELM6X9BdSYL3B8M1G0RE96cXIseuWMRWkcgA5zHQ8yDBWVzVjcnsx
nIzCE6k75SUzxCZJ1aFKcVoSM88CrAgxIkMV/66OQ3bbU5NE2xax9pnfuXgN8qnQ
F+a2HtB6IwcN3rlguu3I0+d73iysp5l5Mwzfpai5lJ870WmpKgbm1SbEzzvElCfo
iXmAe/54eZBskv7AH5znYPIB4kx+fchIRggfc3Z4nuyguI8DC5el3OSC1D972dFX
nMtQcMbQnOdAxtJ+v4e3Nemh7tFoUJG/k6lDgzCnB2ZdMr+DK/G/WDHzFj7WSIwt
BgwZu6qnm+5W1h5zGLEZUCEXKvgmELN8Bbm6JDD8uz8VpCxGyYCDWN09pEZfqqwA
dzTFWOjX/zORfjtwYhwdeRv0hh1mYijS8QKVzv/3yOWZkZS5HX8X49hhW6Ojxgei
SdSqJAU6+O509tPYeu+3HwI/9pcysKVbsLLN1ldR+Yfa+o9YB4gUmaeC4aLP7+uX
lh7PF4uKsaKK9zubhKs7uQgB8pAUh8ozoB4czFbQxRRHaMoMKR0k/QhEyn9oBenU
GylI0AkSEC2CXJgrl3a5sni7LbM/QIbEdGiQ8I8tyxRME8XtCeVX+6tH7fIztlw+
3wvZztCydbKIQRf4onj97mzMJPqghAN2bDswC7apZUDKwAogqhKv+tQToFaIIi/K
eOebblKN6gTevvrkVn8kiTnJp9WrH1hJbDv4NqSkzUsTUpFrQP28udlTF9mKXsRH
1OUkGjFQ98Yfj2RQ+T7aKTgdiNUiEy6LSgCRWmf9wuVbNI6m5DMjMJXtWs2bUnlu
wKwwpBFJAAkgQAV5PHzDjEoi9xdVMp1Ao8v/2T+8mvroUdO0UNDbFIjarKkb0Pe5
Q3ga851J7aNcvqrJj/exMzmUMYStEaUoFV//4fYwMCJw73wIHKWFkf8hcqzsoob+
yU9eflfq+gESJnG4aLWbVtQUYhkSTWCSP2w5IvkhX1+CxrKQj1DOH73pi2m/xef8
zi71zN4UCFi9vy1YqIuoRbq4F9qF+0DoCzFn0Q28LgE/hmEKL5k3fRpmsQw2FPnM
pewIyzrUZ482md0NYQ0/y9tUgeQsTVDXEy/o2HYHW0/dVulPI3W6w+z9C45OThnr
gt/aiMin8PntRbC4FnfNthQMTGAxdWOI6v/cBSkijSw1h5HaNxdtKcKoYkpV34JJ
loBQPFarO0LMCJV5e9Pa5HffPN6bDFgn9BPaapoL6ALuVlXlHA15seQsc9s1mieC
7UOjeKKy/T5gw7jhKFn8uvcoUg6TlP27AeIRGYTMCHIXEUXrgJzXzKD0r1jFhOdL
D4PX+QFUfCEc10WKcpAGZDlc1sKJHoKDGO0L3/4xJa4/nvqWgBnHPAaJLLKR5B5P
jVa4JJaGZ7XaKUo7C9mEwJWedEUQfH7we/ECyh24GdfxdZcd4myrOCrkAOXmQhz3
U4hNreiHLloOGilVM6ifWNCp5LCSAyaB7EaAZo0tqcYI+k8A7QPW2q89YJbYcDdt
63DabFPVqxf7WlnjBlHXet6GXnssr0x9WMgX+l2mL6GvgJdxTiLTKivMr+MZBIn/
IaVENHmHKx0+BCKPJEwXu3D77b0nnMRO6APd1wZ7zCz9FG5gsqt4+pjP6HcQno8L
2xnmJqGPgov/5XUbWXQMCUg1bem3WkUc01sXXj78BpjyzUf65pabndxpQTGFrDSJ
wYfeynCHrJpKgxTWLT8ob5EKcXaVLW5KktmU30+X6OHTh5QeJzM7+yK02Dm76tI6
6NqExfNHmEo2wlPFB5jiRo8yatS02Vwd45/G8i1+NYalVuv7sKzIVybl5CfHt7mJ
lSQE22pDNmbOk983ZDddinZseqwBPUjGu8NnG/TPEbdwaQlvgt8Et9xBVksySO1O
+HQEe7a/gXf6m0V93l+E7xmMHERRIoUHRkx4cDYPsmx3DPgArB9rtUCQP77dbweU
3B4yVB9n5wzjnY+yGP+63/DFPdVxqV6/7V2shPjizB2L+0usFLcnZ7gES97GtofR
/fQekHMYBu45DnsZWSjhG6nqPEjqqWmYtJ5Mkz6C/E38N7b2mNQnSZLZidCae8iB
OojFQW7NocmVR4z7vdBaeFhgwqi/mrWCY3m/gCisPJO33Gr2gOYcHZyg+PMq9ief
m0UvcINm3wNrAgdZWsXDncLK4/o8D08iOL7Q/fR0H1yJJGDpzKL87+TmoR7+lZ4j
nnuy6EHeOFLxdeASEzwQxbiwP7Eduv/eogJ7WwvI/XTcJzOKSJFNf1pI3hv+HHet
NWgePzVhh73hGWGtE3fv1+BzrjdG8p6hOY0y/0WeYz00+zUF7GDVGTySf8/L41im
qML7WoHq/l0/c1HjWrMEYWY39jJIr1FGV0xOJ/2LYOb3mOqQ/N0pN0fnTCFfufRY
jA+mFfzVc35BF3+rkN3MyA1DTwBF8265p+GM3pOhi2qrCm+qj1CW2A7DNmYSUP6n
rw1er68AGjZb+g0d26VarPv3jnfFt9C93pciid+lcjTwcJFCay47qzwbhcE09kZr
I9vWnGeTUSclshMqXYCIC55+C9VGOt80/wACvSi2eP7mxVFohct/IbszlCvZNlw5
bt1cvmmCBSpUriFlQ/1l/BIpXFHASIGnsJ706ipAWgX3tBEvikTV7W8aMSQB0w08
aXwb5HM6H4XnXiji9M4kMqyQYiwPUmYPA+t/s/INhfubzDhSnP23RATD8TwbFRxM
it5kGGldMHrpitlii4fTvdecI2u6ykFxHnPF6N9v/pI1KITpPCmxRSogsTOnEycU
TOIOqsckyLYVj4D2A0HgRkTJsxadbB0RvTfzSgF/EadN/6U+BUvYCUJHI3nKkr1x
wmvnHJq3eaLD7ODkd1FckU07CkVvTLMQqHUFVV1bgBrIMudUKBkG+gmoF+fJETYP
vFus5Nn0FMu+JYZACQ7yU1Ku/HDUwqCKBD0TfGA1Q9T285/C62FR2vpHq9UPUE4i
nIRnN5Fq/gQ6GQBmX9F4O3WAr5eQiYcUEN5HCSiHze82IAAV/KZg0YaJRluNCubW
Q+23FggbzKnaBHuVhH2tqpqS9RkJtsvwIUH96eu0muQ5Smx6vEYNLhTjJclXkPIF
YpgOZve6L6N0hCKV1NZ9E/j783Qp3MSOJOuPboecoLM/bZ+ebUCtyA2jtQ+3XJgF
ncNJj+jK3HCxPD27EbTs4Uj3FLA5PKHuVwkiKRp+p5oKK083ebA3h+D9ju7xSWtN
XGYhbKkI2fpKFQPPsThv3AnTvBdwDCw2K3CjA3eLmUBWTpWzMVhakiuPBoGPCqrG
QQTCWN8f4SU6R0u/V6RF06QmS2lLWKGYg/1M8R7K3DoFyWfydosu0QehnePH2HF0
oMVsnmm1xju100m3GxpokSoJW5dWDInX5I3SWaHd5igxF3v6A8/AFotzoKHpYZPm
3AuhWH4ndl1Y0mvvby0OstStH09UwiT/HExT3S7fQfs/ylTClvUwqOp847PJnceN
coPYiGI+iIby2nQ1uo3m1yKn5VhH6kZENncOQDdh7frABga858P4+PexFT0myAOX
k6zCQGWxmaz1yRN4+nRPcD9JEjocdoxm6RNeEdYdw1IJGXg8pZrx2WH7a1PxjYDg
J4GsQjWDGfYPem05H1vKeUmnrz1XQ3dMZA40930ncx/X/8VGmxy4V7GQi2x+MYRM
OsgrLHsu0ASFyVDA2/8yoZ0qhef9M77nrK2B7DxwwEGEjSpVeO6njpmXLwUmTMUA
SRly3NXJNk4rqd6/KdhgT5OCelFOTzVhIL+Y9GJ/Qcgi05Q9hXxbu3vkYHatFoEA
v9hjAo42rbrPJzn9d8E1dYR/zsQAKPVJEdXEp5aG0E/EWAL/bFNhhZy1z2FKkb1d
67yXkleM+zgSmpdBMVTjfF7Bzq6U8keKXE8HZhWFOKkppC3KwaZXYuEwTqsfcogZ
iRkados7oOGtWNms5JkVgzUK1NPJaEuiXSIhSZJLa5wAx2x2Oi4DCj+3IIZL+cKs
BbR2Yaucj2MmNg867hBmlLW+fE3XCLNchqR3aek0tBx0KM25WD9sMjzwW1/dCCG6
/rMB0T87pOL7tic5Lqzo3B0/12s2wcjYCa0w+0rko/05g6s6fdy0D3IKPHbbQhvH
7z4+SVkjkBu656MBtlGoHIKmaZw6Bp5v9m6yPOeykqCKox9q9qWt/M7KAtfd2aHt
66v5o/FWszTyR7Pol6IcRP10PZmfCroYAqqB0QVfB0149P7yQC8eQ/ax/EB7YGiH
Az2ly2CuFL/+PiBCC2rddMzlsfzhaecfSF44ESn7egftI6STIDWml21ZxwvgQ7Dz
8RXHTrdMEozp0s1/NyZyvCdGTEyUbxvywBrUJ1xz5cXSEBqs6YoTIU0WAyymGrdl
Ppz2fJzy4+Shw2jJUVo9H4w6rZq6PPLMOz4+8D5xeyIZTBsMrdDxZYzdOdQMiD+x
YT6h2gRfx09wgMemFKeIhy0THWic/ugTlJwuwfOFIJAeyRszt/z2VWRytmL8fnKW
AzygTgEikn4HSVPsCD5bwHiMqY6m6YUctDI5Ur5oU0ZyFiTe6R2+2+7zm42kJK4x
I7Eu1Agi6/5Zjrbdy69u+XN7pUMe71HJpH4VE2fRA4ZWtB+0iLFEIJfScl6YoRew
xHn0jK5OoWHOh52desN/a8PS5oQmb3ckA3EG8Px0BActMaMJk2O7WIXPAy4wY6hf
Khfoa3GlphpEYIX4Y7j60jIV/twYbucwdcDZz4nhZAhDI9fO/HWc24fNEUPmnKsO
5ImdudTLVDyMuHVItNoQRttybzRvRLmHTFYYr/6BRv6GOFULOqR0qisfqVfy92je
erYHfxf0nXSoqahfBL02mZ2LrvAuvVWpUXPyV6McBsnehoIxzic8BGQ84Osf+Czi
zYwVUJZ8C1q732Hw5zYz/O+RtzZ7xsYBv8BBQtYmaWLqix/sEMZVLyuphuIe/XKj
WFXXnrduCSpzARQGZcYfmgrZ4DAOE86mFE2vPAds8T0F295RAl2ebbF9yhVYqFlL
LV80tdN43YkFQOsQcOxeInGOCk5HZBOTlagTwSrlC7oJn29L6SE7gCGnhPbc+WzD
OxwJR+JnqymLCBULbEgS600SH6y1KE9Sln4Eryb+42VxEenlS1W/oFpE87kB8bZ2
aeFCy/DFJg12hMoFo7H2pDFEhDJl4e0xseudRiEZyI9KSTaFGxw8M1M4NMX6Qgwg
HOg+n0JCvJ1T7JWmwTVRQI5SPC5hq35rSGIkdx5uSZNny766/vfZcwn+mZeSid6Q
pFui7HzJsIzxWdAnRY5xfygdMrxk5UvpWuiin9aYfIqbu3zTlNPwANzLNUdXL/mV
1NNZ4FOslDxSmXBGANAPDRjkunG/I6EmRXV/rBU0BGAbiGuULRksUiGHpNVFVG9u
7dffQJgV4cUdZBPEZ9YecFKLXh1hxeL9detgL4I7YbSHJhFUTO0yEV+7vZZTPcUc
otmnoTqHNnqaBjqGEDxvPByyFgoTmeMRodu0eWjRegxFuTK/Y0v3NKyalD58zQGj
5mL1HtFBGvAf8nqYF6CJ4RTFTpvunYIQLyixFnHrk1e0OH9bNEq3F+LksbWD4iw8
oQKRqhAYbTBb8OJkx2897vU94xPaHKlbdqTWKUhl9jS0OSeJ7N+6O/zJsFd8uTKI
tpROObaS4tv7Au0aqiJUvfVZrvAeAoolzH4hAsAK9iGeun/MHpTS3aCKcozoyq05
IBSKguYKLwAnI/XYeQZAhOK8S7wSa+o659eI6FKGnMBtOq2X5gKyE94YK8hLj6Oy
efE0+orXSqjZZ7YdFgwGJohVuMTYRnRUEyP05AHyxPMFzYqzzuOGcpXFz18mt3d0
sNj6V5tFNmR2hJerRYQwGLsvfrKsn4u3BS/atAON7TUt2nZPlRAYpDRfPrCaiTdQ
+fpcoA/8ffG2GT60bypbCq7ZmZpvzDeMI6HakU9RESD7uvwFZePxaDiu/VWCF4D8
2osYn0zUJEERWYzOvRkATJIZ0FJWWP5PGspF+mrRNg0/ISbLNXc2o+KrB2dxg81x
Ypw+2l/c72SDuKHazcs6t9H6/t7/HFr5Th3Lvo6br0KuV1q88kv5hcwoxs5///Av
vY57yxtQrION+NRfQDSVs1DmSOwL2SxLrFtjaQYq6OQoQzPMsvIPvx+Uqff2LOxQ
00G2XKy0ordEkFC9cg0FS83qZ8g09cviHOKMVsyLDWC2gORV7oHDpY6QTkPCYtED
+xwO3u4eni01agJ5xzY9QhU3aX9tQwte4bof5owBmySZvzSSxU0nqVuFLZtTvnsY
4mULSxRub4jBy+yyTTns69F0VjNfQ70PcFqwuA8q1N8KZsxwsiA/WlgSdoFt1ldV
Hfl+hGW3w/CQa8+HG5uj1XOkIhsU7yQl5oe3kxdDTrAbr5bn9T4ioiCgz7N2ltqP
rnlgRM08VYfZf/ijj02F+2ccew3Hb1P91dV1GOq3vdH0xYW0EkvQSbQGSp4FL7yn
t54H8LfbUT7UoRrrhxD9DFi4lsz3bZ1ejGsEYIMbti+DjZHxzmZgIJ/sMxkEXxsr
SZXJzclToXLudJgYz0ifPS8mTLRLp1ZC7Uf7wXqUuUZVlxsVO+bOiJyLxvvngzZN
+u3rr9oj1T1r2hAO5gBqrai9OZw5vppRSOsNgE/b/elegAhXtwrVZNBtaAv391xl
Kzum0cIVSNQ7gS9daOj3315eZOG9ZRqPGyLBFyVqQsuHPSwZjdZylHY3j2TmZCtk
xr2X3g3BiSB0FcLyov06PBx581yQx1nf9YwQ67CtzPWsA1zK0mH7gFoEYGPscEgL
QADxR6qpcW4lrN6uM0E8v8RyGnZjq2pwE6J6m1OZc4IN+8jCyTpEyh1L1fh7Lwpb
AMkVUZyMqRLON+J8pJY4ch0M2RCWq3wtSZxosPCG33CzRkkyK3cQCN6q8n2T0uCo
uypVV7hvAFh5HhWiTV0//ycJCtXwE92m9u+tHWD3UlLRLoR8v4bsG+8BH6P0X6NR
aaCVju3u+bx4v7gsKdVhIQiCF6g/nHJsHtYXedStsr92ErGDT60LC2zpGHmpeTRc
jyA9pMsbYsvcBw66WylZ04XbiMtdJ+rNLZRtA2gWtGEdJxLkHPkPoJ/MzSZjqpEp
g0ENRsgsGPrcjQlHQKXujPEaZxiAXI1TOoBXSx6QVmDtSTpl0H41u3M0UezaHUQ1
+ZLhOEyRBQ8Je+TSq/JezjYQquQdhYdWWwPBdO2u5sEZw6e2t4GaZJFKRjBRIAJa
lxHrzULqQkHa63reUkL9nSgd3mXgCu68FQkJLR7GcUkn7/XoFunNdNv5vQ7Z1pUF
eGmcZHQwn6Xf3ZnIBch79qtryFfB0RNVaNFqW2G7OHC2ZFN9J0f8dcXXfvGtWMtV
/r2e0iV4Qgwaik84fdjRSBYx0bwMWPl9MNDgHn7RMJZmUDnA1l6DnLgQKI1AMYpn
ABUE0SMRlMA9PfoDYh1D4zvI7QcmOsClByjgY+140QQxwQX0Q5Th891SAdLUpy4i
eYiB+M4jkmuy0s5oJpGIJ9VzTS0A5/cUQtcHU0xqM6JLQD0hDO2cgCuMYNoQT0hi
866lu9EjnBzyZsBJNkq7MM5zy/30tIqWgmuHeiaqn465eYT1F97Om1NBhUFsrWrn
Vt0r94FW/Qw+71bigu6qXlB2Ti1k+6plSWtRUeZzONzq04S+tVLIGf05Iiw23bzQ
tdEr9R1CsdKCeG4Z5VhI1on9ralCiC/AZDYw4iLV8745UlexPK55UewIrBicEMmJ
2+yjJZ0xUPMWSsz2CRiY2HR5/Nv4iKh+6Ywel96XexcWQa/0oEtvGb1bslYKaSa7
WL5kYcET3mkm5PAOzbJ81dkWVkMBFGjE49jWAIo1jfvNEHkV08d1ZjxwDJknl0eK
GLF/6M7P+uascm+kCZl7OptTTz51DkPr8jwkwGjwsb7Vq05VwEaXsM5cW2HAlZ3R
4FLGhCYHL3AqzHSWErNYSZIMJxla1pCirgMFSthBmM2cgOkfO8kRe2+s0BP9ugRs
vvzl7eP3mZ7cpH6wej/NbusKW0umr/dLhq7LygXR4XBM5uSjMJU1Pa2/uiC4alTl
1vQXPOo7ucLwI7TxGAWXz4YOAuvbwpUj+ZWez4KNvvNXwXlxirRwav8mM/iavjO1
Doj06G0FGHMu6HEYuXQGwGVtPlRoeZmkLxqyisfHBg4rTf1ZwJMaIdHQ6ao+U3i7
6C+kizeNGo1jJXrdaFjbYMxFAQ+F2gbyugJ1cimIvJ3DgwTBi/NLXIM8WAl+VFzm
XbayqPe1xhrI1Fc14t9DKAZhkIYpCSAszhdUcOXPZA50ufiO4+FGnaVrGJbEC9uI
pDdsWfKLc0y8XjVMkDs3sGqTin6tkrFbUrTTw7spcTVr9UAIKfu4OlJLyxDZLnLR
d3Oe2iCVQ3Wjl1N0rzG+6TY2JPoj09dEFHDCxu1YHxSIin3zwyE0BFT5M7pELv1Q
oIrHGQCgORPq4u3DqblotQmT2WyJJ/8BZF+y5DbMEMpOWZx/JwXIsJPPIcJBOnhE
qSOB4sP7hSjA6KW8zhRb5YyB+wTxs+M/ez3yyRyhZ9SWqoFqb6NHLQyGgdi+QAeI
3C9lXVek5lSpD8Is9JHU4tZMyhuNrnUML28ebpVR9YI5RAvPym6t9fLeoz/nhPzi
7LyckA6lccDjH39Aq9NpRykfJCSYsmxbmZqvvnOd8D+btt8GCv1TbRBeILgrFx0d
FLeWYWBql3FhcLcpeun3qNwV9532QU+MQZCZsTn3625FgJqraZq1fpmh9gYNJmi2
bK5X4bqOsOM7mD780z9acC2YN7EdNI2GCw2Pk6DgdNEb/pdXjJYIdOYLTfo6N1Ep
zTjOgWAoYsztC5EPAXntbwb2Eszt9HGXxNA2pq16wdrhYmNGNOZ50Kmw5/mYDoi9
ZIZDG7PAaGs7dZirUJ3tpGUIK9vj8M/wUitT5R7zXOYSmHNbTLxQjXOM0bHDdsBg
7WNerHWx0AkZFyYl4e151GjXjha3Q0M61Z35ra6vkF22V8RLbfEfBZ6D3tdEprJA
jd6AI5hS+txLEkNBBNtva/yYOAb4gwUdszjPu4DUVZbdVuijcmGCwCNBBO2DQuhx
o/JADsefdJomQ6EE2r0YGkwEAncqviHdJ9LjqNtbOG0f4e/cAh+nigdVh1h2lq/h
kActVcRUDe9Cvg58OA4VVvCdi2d+tKUP4tZZ3rGujJzTAMyOwfT2S0jTdQK+6DIT
L4oYjSb+QftzAthmxG5hyBFQJHe3RsvKnL+4A4Ve+1lgsOBoTZja+UwAfKZyYfEf
DENuI/hO8SROB6KZrJpCSK6fVyMaWX/PointHB3dUbDK+fXBxvKquCXibYzmSND+
QJpf3iSBy2kE2lD6k8Wh/3CYKrm3TfvgcspmeBfaVfYVddhN1SNjGTRusRiBu6Vp
6es97SYPwOFI1R8wiITq2oYw/MvIkjJM6AzhTVf+ouzmOg23oDLYZ24hgCbW4TD8
gpgZxYXldbxjfDHHL9p/v3q32zFIKbj7NIZyAgtmN/xofixhdN3q+OakEUdWE4Am
p464of861nzxM5CADXrqlSmbtXslIdDNiR3oKtMI1HVA4uc5wIhMBpB5up+un7D8
9CQbX0bEDGzGU2XDJu1+QODg7u1RjV0M1m3yH/IJuPJ6ZCWgFZ0dqM26+117FfeS
J+tnoc14vJT8dqsPvs/rxepDkPVJfG7cXobrb/O07S2miSwnv0UD/nqRPKLRnnFR
eEfUBL1Ll6mrTgqgmpe1ilP842CyQMWo0DIr2K7tcyAnCoYf4rHJZXqeOaOLCncs
xnp1GgrKeeBJqoWpEnr5DBgFxbs5eFBF07HGjzAfOaGWUfeTJ6hpRwYCH7ToXXwt
0mjnjO+f8b/SMl/evaaFgXLGQmLTcfKeLaP8V4UiLIz+QiWwhReMmLATkFTTGdyg
NDviPlMNPPTt/FyI8AVkZ2p64Reo+lVTXG2ThGupvisUWcuY4qbOgylZ2UIOeVHM
GrbQKuWkHsq+naMBIIIZqj65+zmY5LGRBdaiAh2BYiG2TbJHFPoHjPwyyBHpbquq
MZo0zoehQ4/l0JW6r2tVZs+iRADmQer4KVxuUBL1IeZgROJ0W/ef1yqu0+SK0NzB
ogx3PTvCMzJ9zZij7XZU9Q1oyKEER7rTukMWMGQhHc80U3y+BLZb0HiVcYk8Y1qr
IwBHzqUHjvmXaAehHOJolv2MsGESt6pQNQzSVDmVyqkcoreboakyKImtbG6258gG
PluCEC6mx6jUOFrO4emrZBkMMTet106hG9Va5lgOUCQhTXryMSIn8TkSN7jnQL5e
H/6PFTMkqlccPvNwYHDPapxlWZgxqXaOZCNNdTIE4Y5zjksTNQh2gLgpzy61DuFd
HGiFY/iGcZpHKiQvSu4wF6qzYhc/RRyl9sCRm1/uqC4Da9+3YumJgl9eZmrPpCzF
zxjn6q8SqUlm84r7U+/+LjZYSx3v2WbkhPW2DEed7hbjNMKhWFJmvz0cSPTIctwD
y6wyaLWfhb5q5SF7QM7Zo7EmHIHXndVEUXvDbcRmQGy1IbeGCFPfauoeeLGa0S09
AeVL8mZSuV7gMfEIwpHJjd6zY5Rx4B2rNMo3e0t8CcCG7KgBbbZXvwX/SYUGD3Ru
tncIy5RST61E3NT9hdtmdQjcUGR0U8FV2lvsWPvMGpLjXtU3T2D+PFl9lfN13UuV
xKH6h+KN9CqJ1zDz05k7GFh1VXSPTXMvxJv0gjbHILFxLAHw7jJBdkej7NUsUDMa
hamAFN80+2WezSOjXJFbvlFKrcprO3W9wQMv7mp/cOBIaz+ExW/qaklEulhk9g03
oHrc+tjWLCn4rhaxkX4SvLQGDCxW5yVz7CS7ak8W9H0Pvz+/MGKebZSFAMF0qIdQ
PEl/eTS+TkPcr7kZgUujTt3uu5pMVbroqlk23ofLfBKEmhTbfRcQFHc6MkO7nS+i
8udiC8EQKbhqDx6vhUEslwH3p5dOOW0R5Sonj/wypKDnaZHrNYltoidCo55oy4ej
C2BA843jcbcxi1Uw2McU3cIQMqCeY+QXRKXZyz5bSrOwAxVNJjp8d3caBhqs0ve9
YNuw7eLrPYKpGiVPCgtvL+naaEH/iwAFsbxXmNVUe+q6X1GQRbr9Zdl/jx76pNHs
2GXrAEft/WKx0wkSj/Yc8ZOgpg/Eg1bltCpfrjHnKFPkZ2ukx6qBJfvmFOi/Yk0y
mGUYLkXh/A4v+AWeRcehEP/Ou0lhqXvNKR3hfOeLI75zLDUn9Vc3JJUtQwAtUkq3
Knu4quftdlYDqxyANSMwkWJ+nMXkdIxdmGF1sKg2nxUhD+gFvz+mUOKZ4f8JSW+s
oG1o7kLblq8bebV1GhIQedLP3HQ0hajz1KXAgNB0QbYqHXdVLVWnhgPmgF4+se4s
FtdKhsFUaD1PxCqSvAas5W3YmqzkIOxkcPonj38m8gZyPWji+ZxbrEQXiRmgpmyr
BVxnfjQ42OQR/vXrCM3+rydRxISaL7MVA0J3GaveDQ8Pbtn8uW1zetBfLvKo30mX
11b66cBKTZwaOy5xsKus6XtQ4QiI8goylAl3iSb9juwkA+iWh6wUYReRswrwZJV4
xt5WDDdzi9kPfBoOi9wyknPI1RhZ++gIr+l9Uz2KOjKGwJQwTgtZwOUlJOpMk9lH
WK3NWgD3jKuTFrO1BcHOVimzrlBLo1GmlYwuBOZsaIpIwXZrSIfSeDBjeNACGCJQ
u6KPUehZPFbJRr9vYNX15ysmNkMxm8zv6M0gy9DwiclZVNLoG8+MADmp5HZV8e45
xjUVfawINmDBpip6c6gh8ItpbtEoaVvr0ZOsLmqCQQOIevJDQPB1BgxClkL6Wh+w
HXCoQJblEAbCpR6VzVoAq3UN9em2lxPDvzeYX2fsjBFy6pS+gFjocM+9vCs0RzaU
QN/iKJkVVwVhqF0AL+Z4jK8ozbL2Zt3PuBM/tV8WAwJTvB8vvY9NvVPQLnmj/pRK
e6fDOO/dGnPhpjQm99YtcG9khF0MsBQcquSvW8OvoWYtlwOuxoGxAs/l6k1wJTmB
jUcKVYYC9CUZeQEi1m1A61DaMrcSFxulys31sgFC5VdZatVDcK0OUX9GJqNO8gTY
YDC2t8Bx4/gUbhPU4Ydt67o7PibB0h3oc4YtMzAgn7KyFZpIrq88KDomYg0+Od6m
4u9+8NYfEUvEiUEtriV+8KA7XaUlp5snl5zmJbV4uRnOMye7suU+6fUrvwMkEznw
YnBIaz04NSyk8fAg7G66PQG2STHix6empp30HUKtgttA9dkOQVckpJ8oIzo9OeEW
zfPXaYRwLisn7aDzvgDz57CckzyDVA/w8tFl7oe5y8ehGV2vL7RCEfepYeY3eEgH
J0ZCvsRrDbjg+ONw+7RngjN1OJBFVDRt6O3AiG9l5PZxme4LYCiTeYOojbel440q
NbzDqyBQQrdoKTp2wNq5AZt90xy7R3BrM5IXoAM4XXpn/CqX0n/WDc9uz/Y4BSLy
0oWQ579WMKQ3evQvtR05d6uw/93qmkzmh+yC24OS+mo9f+Ym8I9Nb6ck2+wdSwJr
Ix23VIOWbTO0HIs65rI+ErjxMeVGJJUgabiXhTl7M06ascijmZW5hZpFeSYVdCSq
phV9+18VNqeb0Bm1p9QJj7dC+pPTI6RTRC+02oQQ99jvVCGh/ct4kbKAYE8AqZp9
xce+/0OBdaDMHOCYMWuUXKpJGC4iBfTVX0va4VS4mIvEGOBsNnhKMMCpfFnWx1pq
oiHTnWM4C7Kc60IzFMv2gNd9wogpkLFnd1FaBk3k6MeW1sOiGveI7aTyw4Y10cut
yd1TYUM1g6CZhPmMCfya3DxTlOKvTFbVOA291HT1lWwqH8+tlGiWKcyt2xAh5Vxy
bq6u5Fk1sekJg/pfymQDwUSiItstwAJtV1j2jzrGH7UnTjVw5Tr57IUV8fzP47hc
sVNua24S8qkA77/vjLRwhgwYbrnwBz/nF4z9B87zr5ZUbIjOOFT5cILGe2P/U0/x
RoxKo/LVsifQU80sQZFcNoIWixFCp40eCHnD4XWoiGJwKXMSuaZNhiHPQxTW4C5E
N1F6pcoP6K1KCdqz9HQ8bzMyN8/zQhmq+nQBkEpn71AH3ZD7EK+TfQSajMbP3/8m
sBu3bg0VASzYJ+pgnk76xonrEouUYo6ChX0fwiOPPh9HEN4jGQwmzwdI2q6meDQ/
GaMKoGLcNbjwpV/VmtGgd7ZM8Wr3rYmYbjg+Xo8XuabnEFsAekdn6blgJoV9Fv85
GqqU8AXjYUzMhNRtZwtgzFDmCXSnSn9T5mcTz3FHW4TIs3uoA66ODeX7ZF/It8s7
Nmup1iTTroKDKzV3Szp3Jf7SsoVkP4bKEhHNlt0AdWGQc4QdGQZB5+6KJsitxhfv
Kq0abeSmHY1/loelqtHY1DnuAQ7GdYrn8KCoqtuw4RJFK23ydB/XnaUPqFMSOA8k
Fsa6fVxXk9vVnIdkoyxNuCXLk2CAsVNzBhhyZwIIYOvMCkjIWVS6Vn5hUbUd2BqU
8cIzarocCZwdIHJNI1dsYXekTXLuUZNBc4FIyUhEQNRET7H2/d/Gxdbl2XbKXEOA
AlFxQA5viwR8P3z/vP+dWd/Z97IuTWZ9XfDvtvXydDNLyZ1eHTVryuAtMlyvWPXw
Vbs8vW6LIAqpMHWsiDpAhreRyowizDbsYlPN3u2JpKOfnRmeTiMKf9F+vle9EeUK
b9ecXQi75nhkPa87USSn8KiQt5LBKIj/Z5J0vNuAKJXxWPZ/IDx6ON9RphLimPHy
hJKp8i4+vB+ER16cQh+ZLxYiouueh1xT6FnietVFDS3lH4LULs+V291L6zgU9MTx
2s9uZWk6G1lnayIY9D7MUuKZSw6I1rm8521OFh/6quzViHAOaTeZTi3paAHK+eyG
0z4nJXvXPNADFdPKZctWYdZx3HO0ph/9/MovAOgV14LK1i6J99SMwobEYMxRAt/W
UD2lfEMQEmp4OI/UqjTWC/DOoQvFoS1TeOk3ogGC2tVxYyQAkD5RmaK22IyU7l0J
JBE+StredOdhPs9Ola0t4ucVFIiakUZKW0sQneWbpi//Z05SYc1HUfpskdJaWV8y
MnaVorCFBiOcZ6tOPH8gz3ZVFwttAZUId4Wqr5UKwqs51GrN7O/j4nJvewHXqRx7
rw3x4nadrSUuRrauNZ2GwbywM02MrSHX7HwP4KzyEux6mQaG1MILDwvBf0zb+hzE
F+hYEf0rVzgY/BvcKnwMtcPnuurMF5YFgdlbDgAjSmoTWufPOKGZST4fSW1oSVRE
e73qL0TQbR1rA7HDE1BLhyBraWlOVjamJhuNOSmZw78Byv7T268uENCWsu5mGxhk
69GjI/INCDnKUSaEUfJ+c7YjL6I3JCv3dvjcFA234uRaEd1ZQVVWozWwrjalcK9M
2hK1Ch7oYHtrzPJTEtuXF9XAhOY/HOIiuwKunlAFkxkcPej32sCgvpYc72rCqXcc
EFskkYqhunz8Vd6aRvVIw8z6G1Lm68sHz4Qf7OcHGI6rqqKDhWhDRKfZDinKQrkW
7rEbc+9eKl1ulqqeVh9fGkELW4BNy1yq/k/JpHr5Fpzs1pYF7GWT8bxVg9SotuLm
RweG6tLzeO7r0dcT7NcSaIhHbhdGZJygv7ljYBYsODXkolzsCmgUIb5onTL0kKwm
BsOWYcnmGi2Jk3+cq2BacJk1Tn89Wain7dT1qu2R0A0TVju/TQPCm3lqQ3XPikKm
di2j6UFY5yS8DBhpGA5/pva3oKupdXz2PfdBqTZKOHQwBPPhO8e650DiL4o0IOn7
HwHcFREa5JnaeEuvdc+8gfm2JeY1IADzEStD+lh3uojKKKBpmTsBR0r+/0Fc1ke8
ktz+OegFWnMnMP5EZYmpJjTUmLSzd5fnbmD4nQrY0NZVHvL+DwjF1CHsEn2Txtqo
j0DjJGHMi8q4llVplZfxMG/LX3dnze7e4Vn3tRTKG9Mqg9BYf11AKDYMOAGmmSFc
H0TLEfx3BDPb9phBAi6y2aI0iLROn5Li+BKdwy3HBxF7XMZT0nALwc2OKqf3TQhE
54Ih2NUWQGRb8+Hn/XtJvoRaddtFufjwXfNUPMW65j0uTM6WAaVly2OAje5cpWWk
lKguaUCudxxZt+4XoKdxcwCrm6+Q1+SDVhl2Jb8VL59E3bFaE79Kk6tUT+kUJy/t
hlfoTXWitycChWttSDRainUgRG7b+SvjsjFEBNhgaaWGo7TZeZzRn8gVo6ZZU7jK
H8OskPNYFtAEWMnNHxEY1FF5OJZQJSSNU2gWwZ1Ify9SzGzG8unQcfWvMFqKnLWU
xwI0FU9XDA7HjpthLFDr/EFvE34B3gAI0O+WT1XMiysls9Vsnru779A2D/gCJgdO
/TvKxjYoFewnTdNeK4W9BKZvwNMKHfnIvftpdRgLFQ/35zPSAwjlg4Y1M99pC8zN
R2KLig1RXNGfQodFWpvunzhQEdBMH3V8kxpNj2c77ipUB7b1lhtLn/cAL9gu/qXO
46hGzaXNOzBuUZKBgqMEReyjprg8Xg1fWWToUv3k2E3Jtqxnu3T2x94gcr8O9sA+
EIWS6XkU5pDWOo+OTsgYM3LWcp9AqyHOcQ+KXJ+/7ypUa2XjLAAVQu44HNDxj4XM
Af1ankNnFcZY/231yJ5gSHjQG2eVYoheGZS6mCm/QoH07qem/DG7uzNMXp7CteMH
XKNftPwWu31FOthExT1X9v/TDjhH9x9w7knKyvF7vtg4TELX2NSPZ3SX3Qrthq6k
NhV6AyKjZ2uhDJ+f5j3WwlmjgmQ6X8Q5ee4pc4P0L7spRjWnFdCm4k930/86ATCM
Cp1qxYClx2kXObbuFu71xEZGH94701bsEzlnNnDDtkrSOgv02866HTzN/fWWMv3g
+kArgvBob7oMthw0kjEcfKe4DpWEEmMWTwS2IiI3SLnJ4mtFTAp94rVqJG7RFKGh
vm4fLyIBdSrBFW/YG1PvD0x4xv+ev3bJ0ANbZkiZymtikOQ+ps5/Qz0x48c7D25b
kXlP4ylmY+CD62Z3ygONZ1r2rHJL9Re/kORmZzcYsbqqGBfYZBdkbOKbGshtcuxE
S95UzroiVRzuYtHdr/UsCKldpdoLBR5QoppBCtHLBzKLQ22qm5zTtQDi8ctGtYsP
n3pFxWhi/v8MTgiO9R2JJ5huyY9ZjfxJERQFuhTcXEywTpjPkpqNS3/K7vNjQCnZ
pypIhMo0L0k/Ik+VCK6aysxJFfnrvFqkhFp2QCGyEdm1kYN0pmM0ckOfU29nQoRp
nrf9Cnvk8JXosZNgLxLyO06Ei02VLDIJcmWZomy+SIwHG2e5giFZL1BSe/dvtkO5
ENelSvPKfJu44b1K1yGBz3u6lwYUZvOp8LM9kdu6zgOjPonJ03INUjDpd/GAOtfc
We3qv6uQbgodnDFqU/FOTwqHoShCoafheDb2usF5ilOpkFEl1bkdx84faZODv/Ke
I6dFTcY1XK1cyzdJ08LMafpjUdi3FPRo+ePT+wosYOw+iJBDu2BXVrep0FvvaeWR
3byBJIm9rdUgi30R6FM7woky+gly3bmwPLnEbUHJWCc/erE1Bzuw5fyLsrkDocBq
SBRQYK2wIQU5tUN4+F/0CXkFyDPnWBINiMX5tLsnwBHmP1fF3XS/+BA7MJ46Ncs+
EA5NXsU87LhtYCC3vCzuqtPhe37uGcUZqFXF+weChlm1nb94IYDewFl0yrWBys2o
IldV1ldvCE49eUVvsmk0ug9fQKFwGnV9697qvQlviLIvMCHx/py+baFqeoxTx6JX
hHnk/CI7h5EEt5bSsB4M361Jf44ufb/X9D9Gb51yVadUCRUmsgd1pi8KqCOo8Uor
UYGwCRWgyGlM/JdxnVS8QRCL3bY+aNu09MU6lnlh4qfuZ+BUcH6ejsFBt8rDKCgz
qoaa+qftPz7GGutUtCL5bD+wDBhRe8GnxdydtIbgO9RgIaLzNOJr18MiK+GRAPfL
WFt4wd87VpJ1YGH6TKYxZbQKKw2pAkuDNZje2LZDcsRjGrUT+0iMS9j55VWxT3B0
KMOaq15dSGixh5U+lsbPHllBlUCtqShSzyllPN93NnXbs+kMcHnM+YwNY7V07pQe
XbfP+KVCpSdGt95UQ6mklj3+JYBz/n7S9FbVVMSEfzB4750wvRknrMQEskGE/0W0
7jgdt5DGS/6eOt74cMCaBwFgwAPPlQsv0gyOz+kjp0vnCz+2HKLMJJxCNMiKmlbz
rum2CUc50ik/pvWApHH0E9IlPGA8Qr1dVAGDy+TPZ5djTmIf+GQQ9HjW8DLCMHq7
9gW4yJRe9kXySPBeSH3Ist/NG+z0VIpI2zVF5egV4nGdTQNnoBAJu76XkwiYUN/h
hR9YlcaS5lIDksUrTZ0HkXBTZMw37S9TVko2r3QXQfNrIVYsGuopAsOfbqT9xuDp
yeVCBN6xLjfOaTLDNGaTmOfmTM3Hk2y6jbfN24h122ounL9TUuYZHfW3fYVcTGQ7
xFjTdTa1UVg7VxjupfZ3mB4yToltI4n82+/KvT79WSVBt6MtwbvQXKVHbim8FdHR
ke2W2zsHDbVr8V+F4tpkscWec20PNf+pOv9SCbxA/Pc8NhcNsGjtD4oCDOG5nZBo
pby9Kkh8FUA4zqHzsNSx5GqVE+hltEagOGHvtzuAlnpoZDBgXnJj1dL/uH6gEdz2
D2ypxaOawlemxCm45xC22Unt57Vo+U8u1J4ovrpxkbW7emO7KQoygNT9ntwBkn1i
wyQtw2Kc7I1QF1eaq2DhsY53La0lMEpSTH1jR2Izdq1uP6iEyWI7Fx26oKrZNNPS
0TmWyRpwk40e+C+b47yOzfFm3WxLD0nJIroNmwg8zaSG2hJ4u9vZHMfFKu4D4HmF
vByqrXLcycGYbrhANp+/CNG4pDjgKn7n4KfF28A/sQjbvM6XuHubejM3F+TINreQ
y8AJ7DXIMW9cjxh4ChZ/wNSUq0yrj07SPJBaMr5QrmMMVZYG002LzYuw0Pf9FGjV
b25yHQy+7G9IvVLO40n+4JFitYp0SM5UumzbB5y5vIuMj9v/fHHZzE8myZfduZPg
uzcFpMMYCOao7UDQa7ERYLUGTjf8uE9fnBrzcaX0ZnzfgaII4HdXou1g6iJuf6DD
d0YV4TRqMSvDiSQskFvx9pElDyqp5polhYtITDPQrKi64FKwwU7s2t2bGIg9xFSV
S5XEx6eZR4tB/CTUIvTJ8zzVutguQiDUQkPyGVcnFUSnLVeT7GuzKCRN0cYlInsL
jkdz+PwwOtDcktwX3j6682fKu7VQw7XzWlQJcLfVlcuCdisPgh3Ifyz880ShT5i3
j5XpyUjFgrNTCQscIXpZI/Tbvak7e581qKBuX6qZryKEHTnVkbI6Zt+NgviLi6kP
KSHF/ogqYg+h8NIVcO7LoXlsjzCpZ183NZbIU3231LnPYkqE1W9qD5s0RvtmTpKr
9SmPRd8UwqYBmF5hZu0PGRd16YpyQiJnjltjtMYkJXGOoXwPnKFXLFKatCqM0Q8D
IS9Aeah0yd1CaO4AWnXToGnlasbAqiDsyjiQVj9wjZHuwN8ic1PZqOCZiIi+QaJh
G53oMeFIAjnI2TWuCr6AujwsrJ9lgqY996r8/RLFmaZYrsXY5N2EJ+XUjL7Ghoyv
Z/AevIfFBQPp/OXnFdj7N/tef7/cmkFbNRPfvYS/QJZag1LMiyv89fZ4lBntKYpE
mKU6bTO3SS1/arb0yaBTZYAmA5/lQG8lRdJstQKJRaSRVpfwesv6VH5y1RmdSNdB
Lluoj8dhFjpDiq5WkTfSrqrwVgMNT0Eh9l2qDlcVGNE27dn8DGbcz7jCNIUJOvQ0
J3ZwillJR/BAG8lOHmej6puIvo1Jnn6aeDH41tEtBO0jGrlBRhUBOheqrSVFdyDS
pGbWy1D/QtYa7LRrnO+tDR1izsyOUP4D2i2Zvxkx22i0N1s6ff4Rs3O1rjW63PF6
DYves43E57iBXk8MK1jAKgLwOEeI5XC20wK2Z6T3gi3dW3TjQ4Fn/YaTLZ8PZmCR
W9OyKWm8gMQItkG+g8e5/BJTk0WzEI4Yu6ovQ9XHYVM0E0YBsSwk0h40//l/6uDV
VyJhlEVJNOtwFUP1AHFRD128CpJ08cModrhHer1jNVW5o4p/Ru7sJMuWl61Z9Wlo
Lzh3QTzCKOPEkCLbKVVbK/hHedbPhvPhOn6B3vBkw7KeomtADDxrh6nD2jjnSE1k
Z7/GiZo+JX/D0QRCgw7BwPdiBkKGp/Y2hIBHXYhPkLTeHvYZUo+mWDVOz2Upqn9G
myvukn0JxQu7Pj0GSy7PjI5Omub4u/aV6pGS2x6VXLaqSlqSylYWS3x2eIr95OH/
Lbtw2UKXgfjyIuUPjXgVkY9vQmu1BVjkxvfGZMxEPmjwfdnLZMzighPH3W+sX46/
0B+CBK5/RiqD+CMbjZYX4u4tljBkSHtCceYoxU2U4xSoej4pLaw7NJ/FVZC7izFK
l4z8auiRZjkX2yIh0wM8BYQe90Xtz7QzbmNmltt8n4fzQSYyCYbP7lsvSTt/FIuk
lce0tXTLehCAnjR3txXbH6UQ/GE1N29KSQvC+w5MNmNgX2IrByBkoKOTD0TsfTKu
6AeNws2jyLUHgucpvq6Lch3cI5yggEo3Mdesl2I1ZVJz18G+JDk4gRJeNbWHYuft
50CxErb2XfcfTxW7I/SJkIyj6YqVSyS1WYG+2N5bWozcRvIv+pui05GsnERNyKKy
6nlrzLn9bu+/ZB8yUk/sFSzK1A6lCrndoOR1KMkTMKGoN5OhQ5Cz8EpeIgWPEkSD
G9mhyUFMPSFyK7R4x+vEhQxoFdBtzlDvmyhytCzQvXJZgOJyDij0iZy9A3aCnDXE
ZZYyYwUH7dVZiOU0HhAvxtJem5xRWCJ2LqQ3IbmNXBp/ny9c4um1FzSTUU0Imbsp
sqZvtK8SymSe+2lZlTYGRb5aAyf4sa+cqbz5LT+jiV5NMhCr5bDW06Va2ZwcggkM
nL74VJrRpzw3RD1i4heBVfm/2rJimILI//IqstHi4RB2wF6n8P9KYvNVfjZWmAwO
miB27GDDD/djyITJtbgkc4hB5WdNhAT3IAR+ougCVnc4zL+3shOwOXaLj1sE1vbH
0WtcJ6/xDVVXtRVRUJA6Cb0PEyO/Cv1u2pxHXL1cz1w5N5Nlzaww1+IcmI6qSpnw
wan0hdzmKo2yUbinYWM0i9Rm/i/CtTBk4ViwBiX2U3DzXlBoofPNTZGf+msUODKj
g7VtP5a/C8dxDhthx/7Tx7fDIiyfYcNB42lq+e7Fsg1dk4y2/LC1R8IaPt9ZQsgk
SJQysSS1V1YiMAbEvDBKOn5wdJyDPxFsiPeE71jm944PquhAZ0atXwFaO9LLGn16
n5Prx7wh0yBXiRpkxpAcUoKbqcZ2V4WkiDqftZO0JjX4qcrBIOW+JgZ70wj1D57K
8NM0m9+01kvBfHqXNKO5A2zeqOfqDjqVicxwuWaIn2e2lvcdQLGGMdDhU+0KiCOm
YYg6jZZjSmyw+1QDN83XbybLDu3Ejdyjfg1Fgozy1fnhAJ9Id62u2rPPMrEWiQEN
Fs6PUiSclZ2UblHCIZOsuG+wV8FNZ69z2dFkFnDUGqSG0UZe8AQjyJhOvUgfVNoz
jkY/ZWTL40Mgkeq9aiskem6THU9xjHnZNF8lmKysXDtOC2LVOl9Yrx/to+asfFRU
UOV+Qx7QE3VTyJn0JT5yWt7kyLsi30lYAlWKwhmQNx5kDBzsWCxs5ulHdR351SnR
/8S1GAvKv1qLI5UpE0librAW1hZhlKlqA65Co1+EwK/SayRVRrkYjhYUfG72zv4M
KtPoI5y2KfCOdYIiodDS/zD8efuZ83TdSAVYJhPfbQ8S/fB++X/SwDTOz1tk/myH
Q0WZywQyatqglBcynCDYIK+rf/uRlyE0etho4nGyIU2oMhKzKnuIPQF4xWf7I0fq
Li3jfIRNp78md0WiJP+tOegzM4+ArjsPMhSIPvBBCTdvtefZme5Qe14IsFXfrLTM
6BytkA+FydolgWVyR/WQAADYJBDCZLj1HL0sht42sVdy8NFi4Qvvm5vGeh3tXo36
0xP2j9wgpNXbVovIfJpCPYdv1kp6Kvcs/z/kh/PCHJwH3XpCiLzvuBHRlBeZltED
XVM3vQG8AU91lZwpuse555YFfUlW/1wbOhoytgUwentfK7lh/XGMOGXo7kRl0/Zb
phX4hUFkgBF7D2gGFixbeT+uu315j6lgZH0yAjg7M5OMAnvH9K+Tpp1RClMdae2n
jbSjWIsh01GpQ8vYpIpAsDfAKkhTjgus+GYznHbE5A1pTUDv5MvkR6Lr30RtcmEa
XgP/8sKUJmQz0w+CCsu0tB4X5wblUtabkgVRuUmDKsSEWCbL48hARWc0XvCaqfyV
ux9I7wZFvXTT+yVNv9y6b0fB0HATjZad+mtgV2eTB6wxM1fTZSiuKPYX/vjMToSH
k28v3DDmbkt5bDT5iFk0ZXyXqHCzRzfUMar/8KHB2O8kahBilmDZJLtzQ5Cra6Ki
eRHFPI3hw3yUoILOK51XOWGMMIw2og7WW5WWJI0bFuFOg7fQCBfSPDkqV6J9yLb1
O5UYG9NTaLiw1f2YxezM+BxbxPc0vsd1r4GvT4SHcW/NINDov07+jHhBufW4mnqy
+aumuSW2Ya6k5dLEr/1q0ifUEa0WNEyPiDouFha7qrE3FkIqzAfuwSJHiUOTDH3p
DoNLOWgrsk9wciGA6rjbWpM7v7Fr2pAIlcfzKbc06xX42U2UeEkL5D36tDmRJY/d
gM8yrxfmlemRFk81dTigS0FxxkR66mTRXeJzNqgUk/xkZy79UGjBQv7908G323/h
CbyL1XMpYP1wjQu7B+HW3ycxRTI8qIBWx6bpXnGP23/Yw1GpyK7wLaihnacaU/F8
v6Rdru7Td60WH0UeHi4uI6Jss5gzUQbZjfm7WizpeZottc47KRLZRBp+Xm2+NCuU
XTOYGo3VHFrvGymvVE+ouM3ZRe9Few48N8tSWxNm3eL0Hms4iPaUmIRQy5NKxmVT
tU8ETZG5mD2RP+e/PYxTfKJFqjO12WsafFZZCQSMvNxbE+i1wjtO3sRK0BdHIIrr
ymC8bN5MB6Yq+6bVwO8tn0aEqJfG92e1zJmj0VpZjSx7ImikFqSrfrR6R9eUFUIC
19kLhqnPOBTtyE/FWCyHwMtMsHot9JGnSLLh+zRVA5SKesVLwR/zbP9qNIVnb7uJ
5M6ExEieVwdycuqRbIO+s1Y7qwoXlTJIQFGHcuif4WxLCEVvcPzfj6ZVNQMjzEMC
/K5ADNWSUs9BxqvFr8THkSJAGXS/3wnDwMJQocP/v66xEwKrYcqYnaVtq8CTizF+
2dsdKbp+TlgUlSVny2QTxPZIo41+iDgIgnXr2Ze+fKic9y8sQDjnqx1tyT4N4S3M
ApLTPY9tYrWo6OF+yJmEDZqZGUHG1FHaR64k723Pldn3KCxZXWIG4VzZYNg8OpX+
RqVuUyhCZZ67jiSVymajgGR6KdyFyyx6qGv6TaJyPqd0hQNW68h8MgXqE9p5QLAN
PA0EutmBVWQspY9D5d5Rbzxn/gWO5eRp39xZ3cbkL0smcy78iC96vzJtAuQnRy/a
VOTWYro9hhBT6fdzOGNRuw/3wmut35yTsdo38/T/4gq1rDiYckCGuezM9WAucsra
DhcityqlcQcXEQSZeqgaDM2LENWNzk3V7sm5MzhArJdHZ/2/o5NK1r+Xu1dED8xF
sDkoBUeRkGjevugj8ert8daTeGHyNWCJHZt0oFX9JTz8/vakuppb36fT747oSxaO
+zcAv2MDb48dHjnYzGzJBekIh9/0DFHn1+dPDLYBiTT91JqG6ldMskB5LsXbuqLW
o6ZOOqKerKdLcFrURu6mZfsdMSIaY3BX8/aOt1vsglszJbUvwknFC09VmWiub7sJ
blbvi0kqVZ6g4xIjGRppuj2yOKm3nqYwNWTT/TAGdUA7dgBqtnXAJSR9rLJtxmuk
lBF6Cnf/IsPvwWdBHPMtaEtEU96TzYMXQGFOZPGTc4MrN5673mng6NCPmvLgRoa1
957st4DjkXHFkK/NSYgQLOcg4Qev/mwgLswWYRlFJBK8jFzt2nNY/ECaq6z2yP71
vaDquqD3zqNs7sOeEnBgLTG+fp18i3aQaqOVXzTP8f4D7HFdJUF91x+12jzsfc7H
k4W/rdr99Ya16Sp7El4sg3bT0ou1mnJsHSOhZzbb6Xr7dNc0xMDXMEljNKtywlKi
Zowh6WOQvdbe9L8fr8Wf6k+RNE8XR6j+0b5VnSfgjHPD3UJ5kd/9I5qWrt3k6Fih
V1S2nHcxxVI6Bihlja54R+AvwxPng5dXZE4jdjtTzbSRhe7t4TYwJuZigayrGcb0
A0Y0a58BhEHlbBYn+2bne9WyHvov0Y6BcSOfhu8Y0oicyjbq7PGLZqigCMbZ7Q4L
iMAX7vpKJuT5Omy8ltsq3zKqICLABycIfCjoGyqfC3bAwhbS/27LacK44e78Qk4h
Ho4Lee8EWgvLR11xUvF4ytSH8ynqFDqLzpl+GEsR77L8Uzr6cUeuob3D+NwBOSlW
n8LWsWSartEZ6q9Yg48BsnoO7IYezQMxRWjWq2vDzIrqDF7ItpfClrYOHWs7L3wi
4KqMxi2UeF0O8b9GxuPyDacwyWc/Gi3Zjc4xPp5pslwcLk4029fDzeNbTMioI85q
FTInKr0qkCDxDeSJClzrQWs+PE+ISF632ziuD+yi+3Nt8Ncotv3HE07DxJXfyosi
b0HiNPzBsMN8CHiQ7mLHMqCkgYjPJvodNpaJkC10soUXn4Abcs0EwV4cECoO4QNQ
uURE7yRWjGbw+vl6Hoi0IVhdRcHr1BFgLbLxj8WinM8Ow1WpEW6ipy5872NopBmu
xdVbpsrZMLtJI5Hh14RRnjiO+n1rTSJuYnWZYOdgmKMZQxFMOguOgITak0ZoCebv
SWHsyiR0imrxeCWHu0wj7f3vFbma6Z6+9BX006DvmHCEFp6EnWEimxupT8gkFhoF
zE9O/RVa7x0dJJJEr158qO+TyiGHmmu7WQOOFcBTO0qxW0AjGR5Y1XDcttfbXRVg
dhRjqjnQZJoYkcK5uYYT7+NKe6UJbJrf8CkfGaFPHcdV3IAO5k7da6pPzuXj8OGN
djDRATFRwwwCZjEddTOk7HHqzeGQjk/9H00H/pE7S7bj3umL7+Oa79Zl7nrZfTH1
caXhKkAxzc/lTm+M/WlRaVxL6JZ15SBQ2pNmy6PcmIhGFnVzehhUhyAceEfw62Hl
aXkHSg9PnTWIhO/n3YsTSKCnJaB7T67mSGWtfJvRb8fjx8MT/1XCn4PW0NQXrC4W
R+/WjYlsbsPVQvm+Zuydz3C+vw4AQqo7OB6Xpv/Wx8psCjCLgXUQ/ib7sdawDwda
PH6B8PlbRXHG04s5+USNhBCQOyabqO9RGgpAvXFknOn757wEKYP45ZXaJSWh8WAn
mLkBST0KX2uz16WvEOANJ4kjooKmpLEJczpMaU/MxlJMYBO5/JUl86VNwJXzT7fd
XfFBSIaiYP3qQAGUh/Thjqu5fMCHHLQ53KaHaRW8lpDZfQ1Hs4IfNdY6br2buc7H
xdF0Qkwa1c8mHRAgCVmPYyMoJViH+/M5Ax+DbA/rQEx9rdCPx6ot0YRhYLDyEz/G
PHU6w7Y9gWtDyZYGZCP7KJDzwBxVmjb/j3GPh8wRJOMZ24NzpvlVBj7nOqn0jtf7
EwM2kLL5rgIuRIhbF1unOBJRetdBcgUMQeUS5OZ/Am88JEX7PflCRLUJaS0D+mgi
ljqN8P3WYflHoRYibE0G9ko3V1SKLGV2T4Hx1VHXWmuYr3AFZ4AtMtunx8L3H9hk
lXg6Nl5vni30fOJtRsRPyTCcMl4+fGU30ajXCuYZmX/65lzxaepCuhuRBFZe+yBT
FK7aKLQFRuxngBLnovawasqOXf106lWZjt4arJtm4RxJ8dDSk6hG2kSzHatAkinl
UjxTdDHK/1zbm7R3YFN4zNv1Nw+Zck5VBY4zD4kX3M+HVta40qan9x7UKxKRoTtv
tw2RC/7+u4WGxaxC2SqUNM/dsRSVed4TLRyc9pdFFrWe8SQfc4plaugUoomN+9y5
pCDXcfkYg2oCKQZXJH6wpUaoO9/bEKjvE4UNN5tipOdNGUnDYV1hKPxsy+eKl8uC
wWRdoSopZ+0N+QFtRkYHe2NFCPjHjPmRZ5hm31e118+vxojMzoFPuXmZfPNtc2X/
Ge5zk/hXHLSPsJAeBPeVFRsh5mHSpw2OtgjrNZbZYZJNpcPG9BZnbBOu1wT1bOIC
v9P0nXo5trm6rV0R14ECv7HZhMUy+0CTIicMn0P4eLcV/7mkMnfnNn+bsF5iWap5
BThh1AQJKPOa43w03dUx9Lpwj/5bA+Hp4dF0yprWcIxxkb7uO2PhPmR18oFqzH8y
KfExYKbZ+3WnDolptPWYXZVhWjeVHJzRRabhOYDL/jpashWuvy/J8aCZ7NczKd3y
DpPbj4zSGeuFKBoTuxEX5i0A2nU3DRxrLS8ITI0RNML9Uj4em5ubP5IokCgv1viX
N0gcRbAgoAJAHWxObPYp2lhea2/hK45NOiMfwLYJiA8453LEZBB6J9UQjZseIiyt
46bATSVp0tGxa2HcIRHfW5JdloYBcIFvpzVrnelqIZaq/hdi5VkuIPbJCYF/v9ZE
BSZnkH1iUHXj3/IyP4kMWwKD2HC1cib++HpZxGzOE4wLrNlgpW6mMvYA6LuATxSo
xmwTUZSWslIswpCmsLU4n8m48MI2aRdm4xf45e14JojtFK3lUvqMy+rRdVjgmWpe
OxDqc2bIaNcflcLzpXD512Btc+KfqnScVzbvptTDBf9tBjxTUmmGitFxR5bADROV
S7gG51aT+3NXDnv39tgWzKOBLbhf9DMuqzMhqpIF5UC+8cmT/xF4NkjpC3iEp/qQ
V4na/GEWbK3G/oLdVU7QelVvYjYm4yGK4h0IVhtTdAeY+RuCyGgykFptTRz1q0OL
+MWjWJirj5s6IYSmt0FsgiunfF1Ljw6YiImL7HuCW7GWnL2KF7rGtEciyfSxHrkc
vmbzMzHTZYtNePHDYxo6ClhjVdMbhaEFJfQDMWfggMiRFpc/zaQBs5rNz5AnjhD7
B6O7d9dE1hOfy9bjmmdBmcyaKwBOuh4MgJJyDmIanf8zJDG72RF0hRp9KXRtW5VO
63AZRT+QiofoWw8bI0ncmE1RyqPp0riKTmplmOx60c7RFCjMWbGyhjZzDd8Q3Eac
K3lUGD5qG/fKRgXWstQnXlA417Bvap2X/g0yrkUfagGVxxY2XGr9GUMEkGDvSxfJ
Z4oocqJlJzhsjC5yflUtAp30UZqUi0XbMq6+lt0VkebOR6PPJCx1FdXpxpfZbK2Y
9CH2OIpcSM8GOVqtKGY+IG+UsC02OOcQyevXFM3zKuJ6Y9ergY7L7sKIl/yf+Y/I
IoZ1d2V9b6pRFIVQdM2LRzNWPVxad5NqQMmDMrd5rLxxr4gELrrTOC9ruGVQD5eJ
Wu2wiCUrg2iOHfpwv0TogIc4RyqvYHjeFleXnos0C6TMW1vlMVLcYAmzukPY8WBQ
3kTt+t6yeLd9vNmCE7H1Bn0dGWCmwIHl8uprSPTC5W0+zHi9qB/VY1ug8VtRw8AJ
sMDTNKEEFXq1t5h7admVqU9X9TsmgEpmImfuNFh636dQKkBSOlWfc117VE/+o90h
w7ZzbSE1yhjG97cQBM0juQgAjMnbWPrRwXdVrrG6BMOSNE/PcPXAx4PuiZ0T5Q4L
5Yra9EUtEInRIMpq8bm/jgAw8c7XMFdEX73PPVyQTL+qcZuJ/y4GbEPeO91wb1s/
JzOjL3ojwleciwPrudM0ngeW+X13QjA1Tw5Jm7jSv01Rkz3qGnOtYcFFejvCKN7Q
DFDb1hI6L0Hd1EjnWCd8hWc3rJSUqPO5V9LkqvOTua0fffdRxguO3NAmoknIJaIm
5iUHp84Ihyfgzfs1vFLRNnWwzakGQG99StD5RSFGff2quvpWuSqNFst5HSe3L6Ke
vG9PGiQJb9ij9loIeoUlJCgIwTDJMexT65qhDDyP+Zbzwn3ATu6mx6hRh+P2Ngq5
WxXNrbbKBeaTMlfLTjCi5fXOToOJSWw3GiJuCATSo13uHw9019/5QkCmlgVNMdBE
W3zNaR7mK2AHI5aqblmQZlNYjv+OEzU0zQM/sSrrgWokGpVQw1IBXzZhqao8vTGK
KnbIICtWKKPVEpTOfqIo9gFhQFZ5IcCnRF80guowdJOdSxpZ7sShfybawb4haiEA
5nkPY9ZuGvLGD8CdXtfwpsava7dFS89wHw/EFMn2kPbSVrkLhB0iY0sT+v4JSpnq
sNyMcDc6x8bMZ2hSp+ft0iP0vEM5KWevfTNArOnnpZV/0wpzlswXSFyMJKCXajw4
lh6pL+xbwI9MLoBl5TyT8RCYJTOvfn7cV85bRHnX0XVjO1UTTHCl0e0Oy7Kn68X0
YDWAZytpEF9gz/x0xIP7NFV9GX4hPtF2dC3KhvNuU0tanL4Oi5vYkvuX27X22k+n
ei3XV24DMyHUdu4SCPsx//Qlqu/CEDwHNvgeyaPaZsisZgCqGZ7E7R0R/viV9wWY
6S/22nkYEKNka/URldJwJY6w5bE0Z/NZ9PLwvV8UngGoll+HG+FtfbXn3aesWxmD
l1t6CiKfUiM8FgeDfCbYMU/nXThNa6KR4VdqAms59ktgheNcPxkyUm2G8y2Z1pIx
YcE9VrsfGEwiYSqfmblQAmOfdOVBgHJzxS4UOrKc3PF17fq5XCJnp00Jy7Vgb2te
VxhAgRVOIj+9ZoTE/b5iJSb2/DT4cYhSJ1W61hrhYr+QJvRQolx/M6hbIuPKhLsy
k0uuxUrSZNg8B/pxx+F7jI5OrzDZHsFHE//qjV8Q5W3T1t0ExT/IUwTqKjNs67r0
2jRqDMAeq7kxS3hoBvwc01lLSmqi6AUZZ97UZOnEooFAi24BIhXEIGROBWBXxx5w
u2soEI/L9hsDOVxDs7SyBIgeW7p1AvtKejp6eB3zmEcyiQwhREVzh7HvVjC6biH/
kgD5bMq9f+hygz1fTQWk8QvSmrpBgbwFmxiPDiftRJV6M2enj/p3uPn3OEqZVJHn
d3+J8v4clhaVw9ltnHR2O412HALXOsB/Gg0v42mC74/r+FGwbZC2RIx0MI77JAdz
nQLDh9t2ZKOK1tPfeF/k/jsaJW8eW0ubbQQCVZfIjH0zKU9N4qlF4dB21XNNUu1J
Jbf8jY/1sYFwWsD4pZhons7p1neHy/tA4TQwo9IHhNKJzLQD7FPcInjtYkK94DdA
TzCSNKHHTCZ2WQy9Q3tk1MRSQZyEURoidFPczP/JmIXJdwYC9gIatmNhfJcIWclw
Xs3pIdHq+uZH+sA7BRvene6xgHj9nOloFerXXdspZK4aJCYrP+pN9dvF3MXVk9Ud
lCFHnP2IPmAVXILfVgoXk/SdUSMxoGqODJ9Bxo1CLQ5OX/Jq1YyBkIHeciCOwUYB
3oEpW8reRjo3TzT3DeqPVXw0AYv2YRVfjEa2BOxP6MYExnNWxsWSF/VJ7hTyvLsb
G/+XmyBCG5aL3qFpBWPz4tZ4OiH3Zj3LWMdwHUMRJr+4VHlwNJFi63E6Pxyuj+G5
buswyEWUo4VJp7Xs3I9Q5dIB3H8Vmcv6YGzhz4cjAukBNUQ8xpcdkv18YA9SMNld
UfGAcw/uNzzikcp77uzQLJM0MIHA3sQjBIoG7qBWVZ1YPxtGFbqz3Sf4vQD6KPk9
zruCuOXr5OEk6Wq6kAHstMH7mx2SyVGwgjWs7+c3KfCVUHDYKIGOu1wkhrgXIPY3
gB17v56yeuZ9Gf0wuH3fRHhT1nY6igez1cyyy3bMjS3jJAWqMGevt2CembjFsX2X
O7LrrYkC6JeUWghNEVjuxgzPL3PrzZ2TVFVy/R8tWrSqEjE4ogBYw2hnXi2V3wkY
CMDe+AGJ15axxFfK28OhRKLUY7G3InSHyNLxUMixmJ8jdTO4A57BBX/Y/cL0wvjn
B1pDVu9KxjtKAbN2ZXY8CUCC9o0CU94G6iVTG1muMILKLouGVSDYfR1t7h/LKQvw
4GDxBupI8IutOV+kZWGJBUPddiDtAvOcznZGY88spXQuvrKdaNiILhzm7dO3OnQU
t8LQXTrdHwYVYSOawPPA+wXDgIZgNdJYQRRSNRkBM+ogQGKLqjU0gRr9xghDTJdR
1ueBNiu4Lq8Mws0v4lQVUtacqO10iFv8jr1Z/rr+xFf++On6e3vANOP++dOnv0HQ
o+GyQ0u5hmfeoQOhFZ3m1NmOCKbu656z/myliJU8+dWoiddO6hj1VK3/sxZa7trS
fycglSguv06oLcjOE8knMwC4HIlMEP110FakuWIxjEm88IJlNXBgmfLtR0bkWsVS
/1lusy+DTK/+IjONbjkeu226nxwU2l8SlVYt9NMYeOkjFfqUV/Eh1AyS/TZbWb01
hAac8ncjjX1fRpDh4Pcc+LkNiZbVX8GnfMvGRnQlbNtrfFymAArOV4LUvll8wKz0
CMU3C+sZRUN4L/MNxnmbRi/a8EYDw+H+/+8MxSRMQEcr1CcBWcCllf2SQSGBvEfv
1KGD9vuGUbUQosE0IHuEeDQH2INvBGhHcyrHOzBnw/0G5mTaC0KrEe6ULCscIZFO
jbdV5l48/8zVINl9/bPk9wBe5Oh2SrblVxZ4HKlmYDwNEHkWCzK98iTe0vZelhx5
VsZPDW4vyhSGs3PLE8eih6ZrNnXtEWlrR5UjZ7yZtWFrNsnn9nSC3TrUGFEZllYF
vyzKUwuAolVnNztHg4dx1c6JeoiWBGaJNQCecRKsROcD8azQnzJkZ47HERU7WRMt
PvX7ennnY3ocnBnld/lsrB/DHq4CK4ie8YBe/xlbYbumuwolVDgQSDbv5rfokgMU
eohRBmYlHU/Wcr3cWmptXHoFcuyu5fGiloTA+kmp+bmB43QFo3hzcwQU4ZUV7KLM
NfcgRD0yZtYBmPAqeBpfUNvhbTl0h6D3U+qLSb+oElkzaWUvYewfCAtCTFjVOiD5
GfC0qL3HsCc3VTDTT6c1WWXxHhqf3vsRxUJCoR/j65mg4L34J8TUhCAb5hbRmxMS
mZ3vwhh6jkrtZr08MbJoM7GXCQJMW1RuSJDNQM/IyJNRF1vBu3wJWcoclm2r37Zk
2o/9SlkNBtrR89o5ujcLChbF3kmd0Xx084mSniEQLYDa81Oc+z/raZKiQrso5rE0
scLDRRqkZloktfSlpf6CKuaBkus67BTKykJ2GrwbVv1J48sJuqLPSGeHx9rSzbQD
RtT34hmp5xy0KgX2w/Iy2NMHiN0rRMVoB4Wegd3+12vQ7bE3nHX6wUTrk9RNakrw
A4Vwyljt38hx9cAusU2vgrwUeVTVI0nF+uDtUTHDZp0XElaW/8XPOcBKOqBWwYg9
CmlYxdK+/Io2JWv92DZnWCxtkZyzFXrT/FqhtDqR/IS2UHgo8rjcxH3HWr1xzWQC
0dvKE7RdHP1w5ff683QUAHtCM0ysdZimTfPHh92IBWhfLGXHCvooE3RlPSuFOvNR
DMawgFN9W2c8nDySiirTSnFk2x5VrK5Ws4mtVzaTOIwRAT1KWl9ogrlyZPZ92qkL
XX5x30DEqhqt6QZTt8T3bTpfvRsVs+5O/bZZtOmCrebscBVjVXmOTPBD0uw/TvvY
WqYbK3gjq/L4ec0bAw40HAO8bTZMOlva2huqKvpu3jt6PD2bs9Gf/aaqT8O+LBYm
DZwhbwduNkcfRu/PppyrGqoqcaBNeUhXGuDq3Htk3UFaNHmQSTcaG0XM6NQW35cP
pNSC2opRUkPBtiCCDqogjIkBk9VOrIZRBI0i8aWvNQjGn4qRJSwsMudPC6Rtcix3
I22lYxBNe/rQ9dEGsx4jjLUqHSsSsfgbjpre6nT+4GJYjjg8kfX7kp4uwpBfkEqY
CHgd9y70Y7pS//9xi7CDA9Xf8UdUCK4gPV7uwnCk7LQ+tf/eWkgy/9bjeXq2RWYt
ATTmgIB280UVEO79xZTJ8XGzbO/LQEQl6Mmp84GAxSMyvxCOR+LlfR3ooOcQwq5F
7GlZ0Wc9JZ7Wgs4gsYCIq8bXC5QpWzBTMvh+Wlw1XYDVpeiBZSrHdyKs+nNmMLp+
Ps01M0XSPINRNtR0ZeN85KdrV4WV+saLc+zMAnQ2NhfQxnU9DdQnqTqvHKKK7cT8
ofDOX3UnUlSzVlDFu0VA3YeIJk33d35L0lqon3MDKvdjsOYeFJ1qNQqzOYWFDsMn
ZZ52FTUmpBplJl8bxqKYjkLpHNdhtEB1A/XqTRlDbguq0K5f3yxwUEKkKHCksfD3
39JF2VK4cdiFr9xbQtyecdxIGIP2nIoJQTFuFin4BjAKqKye59nkuZSh9vsL0klW
EawpQu4zT14iOR5AMj6BdTrOIrbJeFzVsAK59/3FWNHYKBsNnu1uGg2ZpYY50WZT
/TOzj4nuXud9LIgMjISLl3lbhZp4saS4m87YTc3ZaTCfVg3HruzMXZopbujYCf3Q
Pc7JkhPijJj18rzUvZ7dhsO9StK1xYCLNHMdScH4Vu75llfvL8cXSJCCh8fyPhr4
XmQ4obfMKFXx2w4VuOAoNE6ietJbwggL2cjd5FVAqpWf6on+2NSdBR2gNdH764ZA
dmMKWAPeEwRsY5fiuY0/5WPuYUMMera7CK5jsnX3Ks9M3sJxyvLSgjOMw2nTzO9v
tWxM8U01jEWCVxj3cQzuN+pvaiLmYqyRU4qhmE7duFC2SQ1CLQvavQal/nHNaAa8
+6sUWL7L/SHWLCW4KLWr6brL4hfntCs2Jd6DI8ACJ38qOwmTzKYiWIPk88GKyuPm
5fjxbYEyAC5J0YGiAlUZYgK2c2ORVGe2AOUYExaj8xbgJJJDTkpyH3qHsEWXORMT
fXfWv4i/hMTUwH67lRqFVp7nzLiNz4V7/x0Z6jDNa9EG/kDdd0Fczq4EfgjluLsN
iphaDzI4VccPBGqL9mywWmlLD88eACaLo2jhj03EsY/bZaySz5hVx/4Q3egzjdh1
elwwUjmNFB9qV6xbsd8PZECsZO0/d8BYYtagdPgFSynNr0mRgWy1/VDEcubrzxYu
dyjzcIVWGlBt4JJPYREu7JLGolhEHDiJI/9nwU9B417l9hsl26QbDGE/Stz8lr4j
U7YmiouQEp7ph7STw9O3vHS2+oVPnvxOGigiLhJiClrg9QYkt4YYRpk5TcXeKOty
8jWeTx4jr/Lwdj4Gs7/+Hz/VAaFJkv8YjN3ldIeLAPMqz5SU9/DZagHMqLyCxpCG
R7F3KdLgS83tSHIGimjO8eM8mFg+Kiat89UY8yZyrCdIsMfS3FAVbUaGyEm3n+Je
p35cV7akbT0UyIpAKs7kX1y0OMIRg3iEgiZVzK7SvoXjlGwpVzfZjhL6HSUO3tEW
xiXf0yv1kTRo5ORvSFelTrBSjkNCjN9zq7w+aqUNrpBmxXqKCgce9Fcrpnhzwoz/
X4Wxocp08uss8HmeTxh2iuyDMxYa5dCpdv15NVAC49GDRbwO3RvShNgxhLCAYDUL
TfhBzIf1Wo7CM3bYMnkeItfVmlweIXPshsalrAd7QVGF9wVC85WVd+AqEJGxakJa
COIWqpfnuj5dIRkZzMqoYyRfpKI5yCUbX1ME6kgqz9mZZCLZ+kuGoJ6fMyu0gHkS
CEB6zPZeeXraR8Qn509RrGk/04mRhkUGLDgcpgq4jIDU80i2l5opvofA0/nKEd/M
9oSH45lCU9B1AEiYGFHIMEdSUkmwN/96e+rxxJh0ann8xdqKXy4k+p/dgle+/iHz
azKKNH5Epm0fCxPeb2j6kwoYQUVb3nZms4GizbMf8lDu+K6HpFgfEctGcJXuNRHd
u29gk4aT+Dp+iKCDgOzSXoRmr6eUJJtgs3awB48Nq+cTzurCTvFYYqscPh+Mq9S8
nxp7dOOKTtwmz900jB+qUxmRu9l5O6yr7MGv7LAaBIxTHzU9mCvzVYGPjNz5Bg5R
n5pBDgIKULJfrSIxCkpg3ecvmOO/9wNCckxFvrPNZ8iGxhlO1lVYv/D1gEJdHaE5
9oLzuOaK0SDJDMqXQdsZjvZXP/b6hqPghMgbDNoYtZEV85VWxsv9QCigabUaBDbb
Q0R8IRVjG4r9BtKATf9H/QL3uRYp0y+TS0wjfm62rtRwI87zJtyKT7GwomtNaKXJ
DnhtEl0PRZ8W7akydDLg+GuxHPfG5Gv4aGp4RmpkL+TKxAvuoMBKEBFos0P+QxRy
C3Xtow2cNcIYFrQTFesTSbwnIr3PlVy0Dkm/c0X0iBPpwGYYmq/lhyOkJXWkQ3sh
8s/FLq4ANaL+/CCLZ0fE4Jzk0DTvVjRJpm3NVN2C9rvvt/fN+k4t/86wCgQLfeYP
OWfyrON5OtsgNZu4/3i0FNFDHRaMqOrtdyI7U4x2GcbziwNBwUouYPVqjM+V66AR
poztd2cPcnD/K7pfvuhI6IjPEScefHbZs4m0CiTQ6Y8qhFTE9v3wI3+21I3wP/rQ
pU+4szsabFHsDvbwK1U6h/GTu3jgu5nWlINPFHuFO5atHbbBGeFcHypS/rfF4tE1
3jIk+W+iqx+nLNWMypxkcK5uGTN+4Kwt7X8xQS5PUxfEQMgz7eEobBlyKzlzDdJP
2RtdW4e84bZDfvMgMYh5WGJcTDT5EyQj6+quEYClIxb7E08VA/OA9O/r8wZ4eb/m
t4EkozbPJR6xBjOzv4mP5AN7mcc/L+c+U+85LRiAYmOCubP5bNA2F1TWXsxUobPC
lkzxwVgHdt4QsegO8YAK4rFt/mV5MuvdA5iDJSyQJjN4OG8aRnBUlv8HT7w/qvD7
0UPFJda2U/BjKixsXKYl9X/4+sz0cLSKMEk93XGpi4CPXTAKeZgLLJssAKuEgN67
3vjQASb8aMEiCGq2ffDc2jw6U7ArKD2v+WB+4mCNE3G24zoz4QvXfjVdSbEuFzey
xdT7DsBtqSSrmqQ4aA13HTZsl9B51K8gSM+GJV72rK9JS2PiMAuQ18DBYLw0MfTE
Dfx9a5EBfXB6gUhJ5AYdS1voSCOc/piFmu6YvNDOI9VQAKhC1WsqEmsMIdJwPQuk
H4Tb6O22VsOMDBv/bCZ+AjfGzFBSkuEQG7FbZ1LP/o3dhw7Qc1iKxvVi8TJgajB1
5pRFj6bGOsqkB5vJh1guzo35FqCo8yz3sSpo5qhDE5cZ018ovvyo5c2MbYtHDV0k
T8gSf/wwyk7jaem+fuIOdJdE9Wh6dUf2yTL4fpNcuqOaVRd7bl0AyCuz3Qq7Vmf4
xh+n6qNL78JXUBgk0rXY8zrwzwxMulexCozFfCvGDTwhKH2rnEGs2e+JII5/1V0y
Dw0b/iYPnUAoIfN/S4fE69cEPEu7sJe9GTZ0QWhzFVlcpq3S1t7OKEmsXmsmootJ
kvCDi5MgsiCLPSu/ozPbl2x6RNzxF6XnFOUXz3nudLXG6XhtJ7MLJ6WjcSM+qpWC
2Smtfh3fQuqWlrLKszQgsTh8iD2i3DAJ+w1A0yhtQeW0kE/ZWWBGMnA1UCQHPGr1
UsZFEvMKIbDgmDYvQurac82rfFM/I+Rkx2YTnVgc1aAII072BZyy1OhcHIc8UYF8
PIJMFrKWtgVV0qawmju5dXLXlm6SavuRHznhvivtlXAoHmaYb7/+djshooNV8KWg
5De0zJ6zxYBqmjz4qK3PpqBILLqMBoC6yv/3pbMQETVzcp2ifJEOXCXlcs/5DsSD
xYufeo21vb1Hi1qdrmdAPfWKZD3BGYV0KLEHw5kwI4FNBDDufdBH1Zxq9H8VTk65
LlXYD+hXQqwiVgd5tLDGeguVZ8UYqvi5toXJZfH8gjManYI+UYadwjJoQ7MT0yyY
X50ya1AxKlXiE5o3OiRNpT5aQlxNn719LdFoWCquyExqQP75zweTnLOmFsBWBxGn
yhjw2cJquZErP1nnA+RMnEJoNE0ztbmifrkNqPbvCjVi7ox1/ZEDFVwtpbh8tyD2
GmA5d/ZmlRYqhsBPnMkhDyGReA4TUWAaqepe3tVm/R5koP+uTwufLZ6+FoRo9DlA
bS3hyrzyy6jP5E3Z4vqpEBYO0qOk+Xed7O63AdBB+bFKMsK0I9Su/A3uUVEBRPbP
QT2JHK8Paj4G/W92uc8xhekyeBk0DHegHlVjsahcy2B2wsxbYP0hUJs3hg14rgkv
698irPlMFaRoDPyLc/mnvfNfWQ9Moh1A57BJ003RD4Aq3t8wfevnfVK1CFhJgGO1
hqhKsFg1dbB3HcGn4mAd/T+HLK9dqR+4pwtikeBlLcsJCkefGeODtwckOoVP5aFS
ouipJSdLcbkxetka3xUjnLY2a+OvBZUx4TU1pefIjukXWNV00q0FG5BBsRJk32jN
PncvCoIh/gGP9w6xGuX5/r5nvNZBrVkOW9z2qDa9url6zQDGIQ2ugNeGCTCyhD5c
eOp58nEE9ElSmF8SkkzQ2fiUhacPifiel4NjBch2Onteh5ty3WBR/9aBG46sbZtb
P0p+1PSvZ7FoZ+I5DakZtfUrveLXT821vnM1xSzZSw/Kh75rQeaZDdYWL4H8oAmW
rtlXkbKdNYL1NA0xWoeRafLE4SSgMnElx37Dz+Br02EQrd81XiB9N7YPPjSXU/cL
48YsCydcwodGD+11m38gmh1UtBbxrtNGkmig95HZK5PQULX+OvQRZ3q/xQmhhsx7
iuo+2Q/v9HaFwkgImtR9aMwWrfpbgi8EY7/4NG4wfSWfjiPHu8nU+Yqbph4C9hmL
qj5kUrYzLqmOANbIL1/y9MXrDa6ycVYl/WLFAL2deOZRBdgYFKKOEp7ZrKH7kD+R
GSxcfSkY5RMpxIMTQphSBx5kcHQ9ZTLPe/uGG0/dffi1yAtNsJr2LDArDaSaL7L2
j7K4Pn2TMYS5dkDs7kv6e7TCALbS/DCEP2SWLtlDyX0D+aIQAQolfD1ccVE/vRBW
WcnAg5J4Fp9vCbaOiYlSsteAIbPFnUKE3zSCqjXsX+zYSlg9J4+rg2cRIu7TSjzk
mB+PoUg4hb6s3sPsFszYVCXxv9thjbcirKCzJBaVPeOP+Bu3+sXXM/t2UDgpWAJJ
I+9++aC8BEb9l22Bg+87NJPmGcmyuCTUaHjeG7wPB5wfUKBC1blFRBPGNsj89QW7
0nzS0CAV0aUQAgTxNgljSRdsHcoGl/EPnxrHQDIZLV9LGlXIi/K4XniiHBZrU/Vg
SIyUhvqowd/T5OlWQrhGuEzDSJo8kmPF6umNSb8KbfafSi5xqb1BqJKZHBvEkrNY
VvUUAdoYXFq4eu5ciEHqqPW6dWFKEKYBDfIk0LTmXcAoB+tVwIN3OLyDVaX/+js/
mcSx1/l3fKkmZvcqL6sOF4QvzVJEGjmvB1tGbfD0i3KVh0vHtWG7OJdTVL1esw9X
8K5LMXuDZH1I+vEP/RUwhV4+BK+lzK5dCGiC/j9ltI6Ng9nHbQjF0pP+m/Svn+DQ
cWMGubk3iUSkA3VLwRlh1nH9w0/8Vv1+dfY2ZSBkslay9oWwe+HAiMlNFsmt2WsZ
6naamR4JbJZgs5b9yAbNYCJXCNaUu6k/a+qjeviQHTyesQPGL6XHcPKc1/hvyPuK
qkvu+ssCuNMp50G5r+yYxQvddp7eMk8bRlt8Na+OFMF/ZbHpOVuwGNMdcFmS09Oh
VnCE5/zV07GdHTnOwyrcBsltn4Yh4FkQRslduTPEVHS+wYIhGsGnKYOiC+tf0RhI
XsYxveWSyZYP1m46MBM2pcAAjE/E4WHsSG7ubhVCdbnVnTjoDTIXWzpJVekbmAVC
XIcwX6mgqXcdhpx+WAcaP/Ll8cQIeBKrzDLBIyQZrkTCEpHrrIErOfst6LxECAjr
/GTa++rXYL5GvtnBuG1OEg5GZ9VkWvVSyINIrv+gCzKPiTtN2ZJ9HAGUo2/usKwH
ZfwsU0eBhxuZ9BcupjuFluZuFbcweYjVZ1sE5zEAroPWjtQ3gSEqfz504h9cVozJ
u4CQpU4LZ/ygwp+VmM7wcf+/6HBiAQlTuHoJjDkfw02L/LeEQgtq9+lXDYDXRt/Q
CgjcS1KYFlUOYTyN8IgMyhbsF1/gnTA7+Ij6TEi0FOuLSD6/Vfhw6JUCP/v3gcf7
JBCtRgrohX196Kbuc5mtHSMux7lhDx4ZmYUo5ZIjsRcUfgT/0Lx96eJUnMZMAQPv
717QAXJ/USAclzgN6fI42yDswHRAfPqt5LqMhWtvUymnvJM281EFpxjeugU25CBN
Z1rVbyxrwfMXDf3px6FmdG5ZFu3HYc6oaXwt6T6zVI1UKo4Pe8YE1Ifb8O7lXFhr
HLiB5tZtvnSvHpnQfy+g199DMiBlFa2uyyRXcQAtL6ViVuPdfvsDenef4y/mkZ2O
+m/yWj3tigLpOlvB2qKFtEesHqByxR07abDF8gXQNyROZpiKKZXGlrOWd28t/Any
hhu+0EjXgw9b7HqnzCLleF+I3qpTdtJ747R3UtpcLZSIQH/eI4zRh+H76nqEsPzO
siBPjAlB4gvKqbzP23D5o+/ZZNDZNFRuUGPb+wQiJjtI5xIup1dj7tg31wQ7JgBY
y48Ty8YMPDaI6uUGsG2oDHUhqzMOVKHXAQy+R9PEMRfqFJASVDMgIpzpa+LnEfNc
GEY3+R7eSaN8++fTZpuHk65fqxpZtsPI4Llz1OB2kgvwozUDjvq24MG9lfaI6aRj
v/AEJezFIvfM66rmVzvTG2882/dXi5B3XM2virBnxxpjBD/XftJruhXAmfrxBjSk
Z8m5NXUYfLjcLaBK9g8Tjg8EsvU1/1SdR+KJVc5J9HFT+Oayh//xhNsKI320MO1j
HNgMBobKixC+BVr+bW8/mXu2yShIdQcyA2TT7NRc7NO5PUkLU74rgqCIyRsiZmG0
kAb60Dgnj16KrLYHn0Md4qGYl1KQJVZqP62WwJdBiXlIJNFeZXGOGRaA6xDgf9bY
y2N6dPAqnKr4dQNesxhIYrXC+qDhmm8IYhHgiopFJVKdSU0/obnHTWCV/TYHbM+j
poJHhBVPLpPKhnoRbEq4UXZp0LqUUGLYqBKr9QoHo1Y49U5Nrdl7cOI8Wf9xk5o6
ot8TypZHy50JtcHcdLrDIAaTt0CHyL2OMv+21V9tddeh7kYZXHTjsHVuhArssMQk
6YIycg5SUHwoLPKiTUVkfhXFnZOYmHiHNzc6oCNGvGXx7ZpMLkWblBVNAbhp89Kl
SvfocTuVx3La48Wvgk9abUzjjjib1uwbtRmb38J7W4M13nrFtXFNnT05G3KCvD7/
pKVjCD1bcu+UCGc9xmcfRhG7lXCIxJwtXI5ol8kfLB56agG89nsluqb4hTXrrtN3
ERO+EGTKYOQhVanwoP+otP931jw3D3bvnvKdL55LlsT73Pq9hPCEAtkxmCqFRiJA
l+IZZcPTh0Ixg57VbBMaKT1qyMo+uMHBeT+ItOJOXpL0vBlUfavocPrQHLzdNzkE
oDxP0At0DTsqD7Ij33eXJn31SYT4suolRaQYytw8Mj/DHRu3os8+jXU0ZXMKfsaW
v4hTsONtgKHb8TLLlrxlfV/cZ554HRqA9wMmBPPUVTEyhd1avD7Mgz7yV/Vz+bYF
YggnBjqXNSN8q7bf7OLjuofK8gcowLv2udvgBv707k1JGlFz7RJYyoyPxZDky4Je
xOAp1sBivBwC5isN0vB/bws36BUdWQKDPT1akksikylNKXyYS03KxvZu+UVtgJ8G
0TDkTDqgEF//L9/i8vivMlsSbFBDqxlg/c8QXQr+OhF2R4DePn+lqua5o9KXzHVz
jBYldnC/BuI8vAc91DIM17SjMgMibscxoHW0fYfAmeM3+yorZxppz+FQ5gM+S6v4
iOIFh8WrS9A4flYD6hv/3KHw2WFJTu6YD7PeMFnZZf4xDKXjY4OVpKo/BNDU2uJ/
UYVDcnHvUrVXQx5ycnR9Gwt+Tp5qij2GBnevg4gYObWlU+Oh2xN+nLOtHsYb0w29
HMTG4a9unvXkmAicXHVl/SeGQaV++8pijqn1u/0fYzgGDg/hQyfaMD7Y6BqlwR67
tRo53lTZbMw8EuyPRplMSPU+vwdfiJS82uaN6ftc5LYTXzPlrzCvHMGvq7hVsRiG
qawvodCr2xkBgp24OYay4uKcddsw/+/DKLodO0neDugcWR72CZHtrD+feXnVjNg5
RIBYdf9DnT0eTpeHee3zzEcFdTJBV3y1cZVdUZRTG9Qv7R7/13nxBhINMidTZLOY
xBetTLSsycEDqYVIz1uicoBSi4wq4t+EGoore9WtZa/RzW/GReyVzoJHUlDRqy/g
qoxh7yJmHxlNzztUvlw2oB0y9OgHzUsDdjYz9dS0tWjmlOSsH1zyBkRTFJx+AFh/
yCDTazu7Gubde34XxKdnqU8KOm/fyLIuJV+u14qE5HbsbkqoS8/1f6tf0mDTwAbZ
m3PCG7zdzG35APdGEZXhNnk+cSzB7+g4aWbzBU5quKjlW1QR5SEvhYkAwmk01cv8
YkRK/Y3xx1zAluJsk0gVG2VwGxbS2cRf50GAh3usZMC/4TTrruuZ8yy3Ud2KUho4
xYNMMmiSqhSqRTaA3OCKO118Tsk4Gw+HpCyPEF2m8RSaIbWaz+hO4K503zqPRL+1
6HrYRnoSiUS+QtGmslRumdKAJ8DwDYF+AP6xOmknjFbVoqI3Jwlr+yFBccsCge7Q
WqiqxMuZ752LAhwBOH2Z9sTBvFfWDaDJP4EAJEYKgdHaXk9lerteEfJ47sOZlO+f
T4/kDoIj5OueZUM3rol57pIz5r5ZmoeP+KE5YcitXEF+0V5AW4sJRQ1V2bOusPYv
OXu4KX1HtpD7fqH+/ogwhQXh/+qtij3lNjuVfxM2ic8RACE08aZQwsMMsiaIW++a
0SVArMk5JRDipOFptntrxVbnHC2gVQnIBGBBpDNRynQlwlFFpYADLzIHOg7NIgcI
LzvMyybSgQN4J9UE1+P6A2oApRSD5Vu6tVBLndNIlX0TPTOaw9rzNfGDapqEc3ut
Cg+s7Bn5aiCwQbg1C6fgv+GRAQNP/oRrUf5S5Om/z7yGfPrsckv3bc48tB7HhBwm
cvjzQE5rgISqa3RtE6sQl/B5Oi9v3IJSJBNNy/oRw/qPwkuipnxB+X9q78QAhov0
8Svg2zT9f+CPxWg/zKSAMAfPBhVdBdEkuRiHE6cBVek0xSBz9fAZgQF05A4nfB40
wdoPXKAq1CHiObsUjIRq+iFwu2UbgtZy+WSey+bf1HF9YQFTnNDjuem0uQUE9Oyq
ZPczfztwNKZH4cuYHpejLDdvPucZ+AOy4QjpMjLgzqU4NG6V5f/ByZQK/5/mtfqF
m8OdzmOScu5JY7ULOi5GPAjEkYQt2ndSbK6PIPzKPDh3xByA0e5gkLnQQX5f/sog
Ffq0Tw7hNOmjxgyuVkC1P+Ka+rHWBXWrxITFx5P48G33/75mWUqqRzXiYmAEWtjy
0q8izIU9p6l4nGnYvobF/RASWtpW4t9Xh4lu2rTXgR97c92wYRvUBZNxA0QpUt6H
FzNXI6L3whm48Aasg5bSt1d18E+1SHiM18G1LJHUEoJNcy2GZRED5FVs/oeUae5W
VXo/EwWqqwwH9IkuAlqO3NabZwno7vC8B48arMGBh853mtDDoNp2e8vPorf9Kab/
enenQZg40jkshF4crLsoWoK5CnKvEHENgoXoPkTNeBbXygd4Zf5LRK9kfShsFVAl
51e1DcTM0IJEKxjnjXG1RhWpewDDOHJGYEHzFsukMp+/UiXNuhCn0DNTy/woFp74
xt/S5QFkLfoqYND5l+cSBrxbiBTEjQNdIAhkd/x29v7imlzWJ7bUqs0gLPn8XQ6B
qPm7MzQtCO1afT7H+BJTTgmiISh0u9Ithtn1MjEWH/i8eOKBubRHUmp9GCBbUUgU
yYiSRRL04IpQp9vLfu09zEBNLicwFdO5sM397JEqZdybTCFaQI4wno5qAGrwHMF0
5PSS93lYaFS+bLkacJfjzqH7mdvt8IccF/t8lJ1uEm9N9Y2ZPAq3lfJWsvDNchIk
G4I7F3lVV3bSxct9kTLqU0NW3d+T/2sZMqVctHbJ13ruUfHxAvBRRiaqwcq+LxEd
STZQT5lWo+qZNkPh/hzbV2mvfO9kjTRlE2AYi2b6EtRMQlGKGHqPBJeYUikqblZF
6DSaLDbaFi3MfcZtxerKB0+dMg7p8ZqCD0IM3epuEfFZzSLnB0nhusbyz/dsTqsw
s2Z2Tc6dNTL5dk6UyihsKbXU571yFSTLa2EiSiWNIFBwbsjeWsfFPkT+BZ/53sYK
WEjx0albOH1EVxENN2Zb4wAOVm6r4ekG10ZcyXNXZAahiL8YTTEeSjWiE6av9gS1
FIJVeB+CsoXuR2NRgazkRA1TD56L6KwV6nCJYutMP6X9b4lyQUw5p4BRqN7QicNC
bCTTcTHiIFeoQXdpf8zjA5zMEofx89jZlWsEaxAN29ZQSrzVE8vebzeXiGGTb4QG
Q2QWbAfy5T4r4/PZ1bZOQ36y4e7DyFSjAJit2oopkDS3/ulv79mL4XqApAMF82AT
+/ZdGHfvQThksFMbQ7bAVqmDKp/oRVp078QfAMKh4nvTwQvDdke+9PXXkGhaRUCL
D+G92iiVlRgkTU5HrFIE6v4d1dST8yZK299r+0zVpwmQCPuahTa/93BmmE3lnIZX
sxdL4Sxk4sUtn9JXb8e07aD7c5QCGkZ5fdsK0XUgVGY8iKggWZj+zlA3Y3sRy+Do
BhgwTeJYupvaQAmBFoVesWusNkjFk1WEs1F+RjhKdt1JxFO+vPYpbIwD0Zj4t0IR
8+ygaOAeWXV4UWRB1LoONqtmuSLZ07bBMje4X43uC9jAEoY6znTqoFXDDqGaBXP+
vbcRwm/emf+3U604od7Srowt14sexZP2b3iT+F1tyVhJR6NTRV8Y9Ko/wFfDIDog
Qp85eMZXJg2W7WTOojTjTnW4jZqAoUhXmOrlmO1XkH9JjkwuCemh9ygOgDN2QqA3
JAPUR6XhGWGk8S9cv9PBWgJMkm/zvSExLALM+IpS/8zwWWRxKpxlgAiSCWkaSXZF
y9x+oefvAfAqiecDenW5qP903t8W8iqsFi1U5qjmwK8YdNx/3Q3H4C7KHnaG5Bg7
HXp3u5ARTRGFIrnEr1T/MDszmqs8kNnbFDWJN38twBRaKb6lsZq30I9B3hmNnNqD
DZFewGqNxev/ou7jeoFbdW7lkJT8ws9kbGgW9/YqYEW0NLq0lFx6bVAAMm93RRNx
plEThVZuWKjciKfAE/3DMVuVfsIVubWJQNuQTO8jhyCvRtS6Cqsh6JhsaaBmdfdT
LUc15kSJjsFyQKeQg1F/e68qD9K8YUwEJUM0q7EeFCJonXM4FisGX8hBquwm9M7u
IPWGpJIYNQEJc/WBS6vxpY5sEkvuVKarJZGqitIu2bcDM7yVSzEa5qM4FoA9v2IQ
Trc0kVqQH+s3z9QsV4S+V+eOkPGpUf7nu41vyUuiRsnryJBV5z+gxOIp/1E75VX+
LCCG15SpWPAGfX8qGACH8MSKBgr52rI8rtzlEvDWMicZfk8+y2KHJWEuQWMJ9k8e
eloO1pT0J8yBn6K1jBq4ivoyFHQqKMgrtzjPuLEDNVUJokmHHZJUA7wopWqOgLwS
i8qoWwpqZGavRF9KvXLwfZJjfua+aZlX7Dv+invocv+JkKWH8LeZFxeTwWfLAYDi
mCeVHpvxwe+XDt5S1bzRBWG2iAUGypXXfiJeWH+spBLGO8YVrHlDNMNj2cmez4Il
D3p6QrDBmChXewp/SjQRr+dGhyhRE7z4KjAIR6N+jLbtuKRasXAmzEI//3PhQQFU
32Re8JeoSn9kFLjBF/1P+54Cm7y7dNLYg4knGwauKMeAZSWQ26KyA8P5I+6MvG5n
MVMWCd8wJlDvbQ86khXQOiAQ867s5pg7SWj4qemSRq/rft6de5ANpzYber2nw5XJ
Yw3gGnF2AbmpyMQJ5Wt+NpLtUg5nXB2r3d3GeFhGBVKgqNXfm/htEy74g8X4Zhzd
ve6Jtqay8HpgNmj29JDZx5LGBe4iaF+GFEB9cPy/McI/sYMwFQw73IwVrtq5Cmnx
ePGKkugJWYTaHedYzFWoSYJRpyArfEinybGGTF3+YtNbMpq41zDL0KU/mbeK7Xnn
wMQ4opPZT4aDnxQ/8m6NxpxUABMO0WSXGpcJsulMaajPHGuAswN3EJxlDn3VClhL
iTth7ffqYaXs1As8lQdDGM1AlXnWO9nxqUxhR4b7asv2lIXWPQ1rInBeFEsAiJh7
+gDTxM4h8OVuNSv6vbM0HpWZAyjYy1BSpKy/OHh/yVMq3xJjxXL4Elsmw2u/vToB
FVf9jE6OFPjStPS9BCSHFxq+CrL++QoraY6yKlFoDjBf6F951P88U7izUWobIlKE
6FYeE6uSHfkiWEFGa5+QQTXgBQqHo3AF3an8aNvw34yoFvWooJvFshrUkqkk2Opg
PCf1kCGpra8n/CrlXXgg5EeTC85yJBRTEtvZTJ5zRBpBsbwji0NVbbpqWb9nvzSa
X1Km5pPYlTb6LJXQIkTHA+KN9/gyWyOwdoEeZPs9C4X0cXS9or/qM4tK+W764C9P
UHy9SyC29R7yLwSF2FuTt1wTbj1PM00qnryAMF0QbhQ/ZghYh2TpnMf0VHjw7sWH
Oro53Detw2bb0ft1YU6HHKDK1p7QDqNmy2Po9sKjJEgGmlq4eBKxTQQ61iwkDOXJ
jUOVbuEXyYI/QhKAWzU/1+WzuZoH5elykzdeS1+EZ+W+xwbB7zh642am9MHAxM+2
U8EiwwTk0mShK04cYW0emc6jUfh0oHF/i/bUdRiq4OwcvnaQe62upFSX8jHg8LrP
yyqNPTbaQWyuSoktPBCTDNyDvJa1ULyOS84qo5TizJgcXGShaDoqT9yxSDxIwOtz
FeMlV6+OQt62UOr1V2Ja0jEut/a3G5ul8tm0xGWugkiSIfUzWBMNep9ahJHYWIhz
ItLkm1awwi9AsumSF07o3hmuadDsofWHwZtpd32qm3c9FhGnECz/fctvRwGKi+BH
WgZL0jWL1B3lSAOYXJhf+VQ2yOrxbOjL+pJLZcDhHYBEbxB7Xv8eby/4goVr07dd
KxEon0YQDa539NSvLHqCXbmCOm5MrplhQR0b3etwyi1k1lGE+HC8moueucdWbTpv
EY5ovN04ub099XR6G4BjhR9vpcjMlEFKetvyClPrL+uP5wvGpjheaNlpNNNlGZX/
KiTd2Mr1vP0x/eTOmnGxdTWcHaNIro7axLSp57pT7iIQXKoFKWJFKiYp9MqQS2aC
HrmcR2kynm7x31/mOdqcL9q7vbkj5rJHhPlGgT9YVSje4shYp0/gUKLmiG0aA+Du
KND7ByV41xcHn3GhiydDIIHwD7NwicLPlTJDOBy6KP2wFBKFP4k+ksg5/9/ScTz9
dS18M1NHXi0R1OQMFyq/lCc5DkT1QCEjFKWNyYWMz2vAAkYp4Kop/VqfiSwFHi/n
ylN008duihm/nih41hALrgshf3xaXm0tZ4XrIw5L7L/1SqH65Rfw+6WrFgLe0XLp
J4yOlZm2b7HLl0J3l4azrSqQNGovT4Fp1b9vhhw3NLCom3q0VIXwunNTtR4LIa5s
d5zXKryzC+NKP1ubbkY1a2W6UBKUbKyBgKev3RKqF5jh4bxK/Y0OaY3PmHXDzlnq
YF5IaUOX3wwzB/HvJMPXNBJCmL498MFksHEhN3Npc5SGc0rWw8q09Ze2ekTI+ZTN
CffklnuD3MTsqtz73GcsrsJXD2Up+6jG7GHuSsXTA5kUQJ9Nl8ZW/9pG8wDHV3N0
zFGwru+E5lEvWkIMwhU9vdPmrzhBJI5SwrM1APIP5rLf4NTbWsTwtialb709+y+N
IOIeEF3KugFdkDc/xlOQ9tjsFy3Svb1zxzAwxYUPyYtQT8aPKlLvd5/oLF2yRbdq
dvPB8NcY0aInuAxRcq7bZjyy4JiCh/AnJQUF9QKP+YClf2htBTYAjR2iTN99Ff4x
tiKmLtpIrGKpEZ8FmSLoWWGDvhI+6IYSC6nJDy3sbVUidtWCQd6fzrK25qqJLiz6
GqvlRFoZys+QVFpamaHdQq/ZuamHz60hccqnMkvbJ1iBIXk61igBy+eUprY2v3sa
5M5A09ESC8v8zEJn0tfX4vqz58vYuOMUIvqfQDTnPCZgpEEJywoJEVeWtuJPIRSK
GjYKytSoVkXpZ3GCXaICA2mzWXrotH7YtOyvWpMwuo07YRrbd0AffR1Wof332+89
iCjjlPg08vQwQ/Og5TvcuThK94XPPR7ZSE+9R1Vo0Wf56FFmmxVcjMck236uUu8z
PvU4o6cvwL+IwaBRl2yuMUJZ1v3/vyS5vE/UOH7DMlbpJhyyzcumBEsaa9swKn7P
+pnhNqLSlVYfZEANrVAHHBDu70dcSDAzjxiAKz/eeeoheC1Y6+u+g2HveH/wqx8Z
W6+zFlJkG8qSNL/9XN6S2Smg/6cnHliUyub6mUl/1ubjNwVeHWSo5oJ9IVh01yBU
iDAuEUgqiyC+M/DXqkcD/n60offuG8jq4WZ9MAHEHqBLVnaop0AWry5tgdeqpQr7
Vc12s/vCGTPPcKa+PqlWYjA0ePfDAoxK9E/Ojadpx+2LJdnpT9DB6R+tHfqeF6py
KbJwqiVmMOhZBb8aGLOKPi3gBI9SKHwKOIGiUa8RJ0FX6Cut+F7+mmjNob4M6+PE
1PDJHhshxPuyIhe9xqapTnYggTW7dxt4YdmEAM8SCT+esAyDNqV93kf5aKXTS/tp
KOw+1nsQ6z+v7uIK/aioIxj9sj0f5GXzE9i8X0rt4olzyu6+s2kh12GvNCoxrZHK
se/MVQhCvMBnqIQTUoakv61Mrbh0u6mWmbM+l+/2xAHFEE1KetE7hQD8/F+XTh+P
/Mlo5XybwnPzSTcEnq+Hgs7CE8CElomK+AEO/EI/jOZGu6YTOKifrMlsA2u6nz/b
4MAQk0iL1ZSH5nXZreFMdhdqYVbGDSUJ1iMPF30dtJYm3Idn1LLrEKz7VW+mMrG6
iOSVNa6tk0SjxYDamMgpqBtrne/M0q1MCcICZD1Ke8gZr7YzgFzl8/oTeWPbpdTP
P6uzYRO/t2V1/rKtjjhXtmLfHQVIJACBUxhPATNxcqCBvKyp0cRX5SDUfHdbyaRn
NfldLgwya/bPd923MLXNBWMAKqRAeJyahPPaS0eRGfkfEK/zBmEZPwDgRx7hsTDt
sNGo9hhaO+tI8R8CgevjB1EIL65bipNVQ4Z3y+S7Gl18w1uGCEwhTZtj16DLPHFR
+0ECFaTIVHyknTS2bT9UjhgWMeYKHTBGhByA1Zlqk8w2nBCNuwFBHTZJbVnAETTm
loS15agpqI3nnahxbiEcbmXAC579rkKGwPXpbhN7i6uYLzrCe8cLr4XrnuLQz1PP
4vLT4Y64lLuIs+dnPaXyMOF+R1GFVW253bqcCOZZErXvqIqzAFRRHHJuCZlzscMc
Q3sMe3xnHBoyrdkElT0/+FmWKCwpTKKxyTFPZ+s5t23JunD8v8kAPiFVOT8xDg2s
/GL2RI6IIyf//dY/QYV+x/m+Ks9zLvTm2dqJKnXW66oApaMY/F5KWQBEosDXM2gX
Zyl2ciojkaK489V0lRCWqInzBHRauRNj5TyKzvob8K/8ZQNBl4XxrFaw38g3+5ij
pwovEhDkyUJccV7E9EhHOGbwNaLuINVsnrI+yd7ERLH2jbgOkHhdcXgpES1/C9ba
eUZGPBgr5M667E54rpAMQvyrEd3e/gckMee5kg1nGg/8w8qsCU4Jfsd4uLrlO0MZ
+1WsCfYs7K8RGUvPP+PL6zmzTOf9UpLiVgVLe6C4X8k0XAVZ6FevNn1Yg19LZzJx
NNLxQAOEp6WGPV1iTaOcyRk4rk8FQVTPRJ/+aL1I8n8lf5USHmMjB8BW8yUdVUOd
rtRBEjic4bhBn+mWUBCkYUqnaw9E7fie9jJQwp4f+pM54CzWKfOyV8hSK5jVwkjI
5oiZ/kHm7MyTpooHvrUkXD9icn/H7+82OsxWfUZUHMEPm1v/r25QXWEfT7zcQ+rN
9RZew/n5vb5IzhhwPlszn1xHdr1k6U3120faA8Ubqeib8TiA/PKSTgVyDAYomA9Q
zJ6blPWQuM3RI5BpW+tJMH9kH45N5647t1zAwOw5teSBWHl9ouYFT5/HzEAQ2Kv7
GMnmJjEY9ArnxgaGGGI8dap0E/qBxIFBTh3nURmGHCYnFTAlyYM1mr2OTSgSjzq+
9p+xJpxN3xadSjnZKD003g8Nh2wYByAtaVyR8zWyQPsjvDm9mZ3pqbwNi4RevK+R
s7+LBuAOm/VJEj7HcLJ9tki54JjRtVUKSDnMU/YRYxVbZoN9aUzBRnEMfQuSNssp
cz2sNRFrmTTOBpsB9lxe29/CAYEjsOQ5fyIDMnbTZhPPcahVyTDMsbk/G04+2/k6
CNQg5eZ9yMWpn0wd4PQ6Yu2BEo3bWmUAnuCdU/c5qTDZaQiv8HU9cURHwGOy3Mx8
hNYzji1aCTTX6c0ob/fVBjbKysQeoUoyj4So/31uTzw4ojx06FkNruplnk0MROHB
+BRPMV1dfQwT2+d+Ed1cMzRsw98un5cGSdC/UZ2ZygG+Qbm4zELfTEal+kCGsliA
JeJJmc8mBCxHALfYnBvg9jgKkBQAu4EAoBprVp2sfuzQ7KapClP9tLy1YxgkiuxX
+aMTNJd3iwoFF+9SKHUmhmPsv0oiMmnCc/7hRWPli4VEPLi0E/1wwyy4RFxj+KKT
kUvpzKk6nljshlmSpOnCdrmN7oUhFBJd7fXlw/5s5pfzMeZQ7FqqCjIU7GAlRhGn
yRc0tIpU8GTN+PJjADzboQcCrtoNLn6ci5eWEEwlxK+3RpnyKkjJFI9+bdhAuSNY
e1y7hpKya61MvqkBVBW2SBed44dztOaMeLHPFCVe6nwJ/v7Sj4dd7JjupT+c1d0M
IDcyI3y0WR2I3KCx7O85DDw3gIxEnw1Eafh8/0KPlOnDsvyanj+kAFLqFr3jS3ad
noiteinFfvor/1wA5TBL1iU3yyG4ywbWGAtEUM20+vQ5IoUnJmbkZqlkuOyEy6gY
h2r2VHDErYtK9yz6oguwhxgFFC2zfjCl1Pa+z/JBBqIBv/LuO+6uvVnBUYPfkljB
PW7Anvi1ln3gqHggw/KEsNkkdTCge74WnSzvu6SmPzp/Qid5qR3b2pg3/r3VC+o4
Z4+aMhCsW6jst5KPlB61Ku3SVyfUNI8DVGSedLNHkByyIcXiyP7DXyZF8GzWufqL
mkmh1COLG8lti2L0J0V/N8VuEDagsybVYdNh2ez3bg54DdgoBG2EApae6DG9rs6q
v1qkR8xSRHAsPGE2U/P6t3O83BQqwusw2hmOyiuVrBWdlpHLbMP4m6Q+LLi4eoHb
FGUsn6Mx881Ib0VNqVbravX8EYTpWuU1Q3szBu5DBecC6CYAkH67dkTLOty7nIY6
zW6DQR3b2y6ZVElsVbhJj4lkzNhtVbGVfrfQv58UvYYJo3nO/uuCyBG5Bw8f2eS2
XH8b53rO33T9y0MsymMRw68smHRs/jb5g0XYwB5b825JJ6wo8lXRwMZPdbbdxH09
azTxaZKasAteb/zLRvd1QNlwHtAFN5cdNSOBEEMF+x1uQRUpuPHy5zd6xYQ+3lrp
LZ2fUZy/Ov52if5wPc4vHrYlqPBbHpwtcLOFOeIXVgb65xcPBqwEeIBHmCSDHaKX
haXJxMKmp+v1T+vSp+cq78mxiUjUz7Db39npgz42jy1Cvw3rpKUt1As4H8gpp0l4
waZ3RrwhGIBkII9zfRhYsGwDIhk9WTfptM1M+mRXH2yN4ZLWHdqigzMaf4JoX57y
rsguSaZVZhajLEbfmCU6HTK7pLWIb+1yId/ySOhmq/BR1sIfr4TqEU+lHk5RcER/
MxjxrvfVCxgZLCpumMgNAd9UtbQtfGUD4l9XYlHOP60VmQw0gng/KFnr1UqKp5k7
/nrLuo76XgcxnXiuMPTTzXOO25LeP81sX51eKEbk9ODFrQEEd3KNpvEvsaCCd3uU
zxJfPRnX+8ZWbp8XzJt+6C+GdyqjJbYk7ogwLHdd77S/i/RC6A+XlmcksNA24WUq
k4TQynhRHmZjVPONI+CjesXkLu2aQojf8JG6aJjHhhz6lmBXlrW8w3UhNPtheddT
uK/5IxE8OJT7MTxqSFsbxq4Qh4kGHZI45JZTFOEHb4nKUEhGVvNnNq2owkUwuqUf
IHt6xNdc9W9Wl2qfy4cvbOhNgXqbE9pyKa8Jg4VXE/ZmArssx2jrpFTp5WhzdQJM
jGSDy5OBpI7kmVpYlna4RpRAGpLB1irx+ZJpegEBfOviVdCNE9IYUHVEiawFbOsC
emsRLo1u9hQA2u0TaABJ4Vj+JdE8dhVdLk738+74n+X++fjFeU9xB9bvvg0mBtEO
6ki0rWqtwLy4EzdmMQowNuWl10NM5tTMnxKpzEqDm0H6J+i8fJSHEZlEckcIb1q0
Y6vbJhSzi2CBIi4QuUQyjCS4BM3gYxRhlghCUCYOyY/ukkyehPihwKmt9mDFn7ev
33BSxo1mPMUMf5Oe8y9+I5s+AoxM3NHGCKOTyFeRdEDXqpTIOZR6F+rYWXH9JGdR
ZpmMI8w0/h3iOC2QZF1HIJdz8/sBi1mzYQdZMF6PvSSbCidSEShL2CLS53DhpV8L
aRLtEixo4QnAHwG6PT6/F0JTNBDgQZaNAZg9Dqt2icc0xGwRUgNcWdhNG2X+OPTG
tlqon9fcjhrHKHDoHltzbejmBwW39BP23nW7hStiZgTvbt3zYS3X1ScI5WSNG5cq
hEYFEZBfrvLLA7VMTtzT3xoxSdFLT2XHIBK5d9WTSh2wl5yvaukwIzHJMw0qZTN4
cUROfsJwE/4ckInrDgfrQnnBi1854+Lm2/G1bs0cp0uZSi9ihNcCdRRU8PsHIoL5
OS1/pr3bbHOsJK15Tru6NTNdiNga09Jt3QwWtdQtuWjfSur4/3iLqfcc0xrEUZ33
Tof6MfL1++tY/4zvxWbItQBM5XfEaqbqOdl4TX6hEFBikjKRAzIgYcF9SUNBK/K8
PxFyeHL5ZuP88BAZfst3nYMi0b0Furf4XPiJHS6bLQpfg7M2Dn73/ByQ2BGXAAiV
XplieCDYRxAYFKJY4Xeg4OdOutqXYfBqdLQIMfAQvhsauaPDfoPgqbcwb/NqZFwq
IuAaGM6j3zO/5K5Msq56hq53AwIjHEtR4LbI0Y9NKjhcnGcnXpm409eWvlow+Su1
q/oXG+QBcNPIcwMlQz9KJAcH0xpAKeZL8OWX8k0shqH7ZmDe2LnA6KmUr9AgosYm
6tq6AhZUTgcq0hMa0fViAifXjhDdsSfngrvxowOKrg/EdOsnm4jQ+dWyzxFNo8n4
SKBVzXwykqG7dazcmBe975oJij0HD0PWl4lEVQIRGHQHMHozySv7XWi5xus85tFp
VLcSpCX/nIdSzbgQbTWWKsRCIU9LQ5NYXccYKuLLbqYI/cm9Nv96E5StS7UaLkCd
T8kpIdLwxyVs3QD+uaXj/N+oKfQ9BZPyAKPvmYd9Qz2w3GyPG9b+9iKW8BAAFAg0
7wJPrGlwO4Pal04LQIpBX6WPwcTcPShU6wE9gbWPVL88ajmInLLWiVtMx6ntRUpu
2pxUSfGPRtmh4kj+9tbgtOW5QeKPL+7S4I3sc0txEdSy4gORxDOhBnQuVMWxYZbm
OOo9n5WbhonX1bTf68Eml/F4I+N65b2sBIipEjWR+SODb42KOL19BH5IgIxE6fNf
pSU8/Sz/DtE3fs4XMxrjLKUcdWFV+COOJXgJDbIGbybEjT0CTv5i7CNj4UdVyoLt
pmH0MHRpOqJ1ylDKgjdrlwqbpr7EOTqCdRAVpnNRDX3Sa76HX9TWuHzG10a1uYt8
LP83MucmXxK9ZtRpMA9pxSCXvOaRblOv4TvPVjqvuoXbgBusnFJR6zvEE9n6HHrk
Yd+1L/0khEt21WakoTEPwRXas+PTkQXZc1MyhASOggSE9xS+lXMZe3gYbrUcydWi
RreivxcbemgQ9c/GDRjm5ssUstLmV7lEeaOl6bKDWqHSOxQXwKVcrgNLAWhS2PyL
YXxfrQ8L8Wku1P3fXMgM01552Vz2u93Z7r+mI1QoxWSKDdtgC4uRpI2orHragt4D
MVI3737Oh5P97JHkZ94/DWIqCn/eGkse1eUoYu0Itw/xCc7P7NMEywky9Q1lmkx8
bW6npzABP7tRDM1AWQEuAKhJEQRRgx+kWWCYu6I2UGK7zwQvjS4KjoZezx9T6b1S
tIwYr8lUz2SdCzdzJkF/ORkM1JJyEBNgsBKizMW6OslWT1E9F3X2Jb/TTxP0T9eV
ZWEzFJyMVMRHUmhizx+fQf8BgfApdzJh2ZJApCGzKLdIysgP9jnvs+Fq18jamzCE
O1aXkvqdAf3IhT2x42cRFYPNpeMbNom557E+eZl5Z/EHrfCnKi5fsFjmG+h4YBcs
+z9a1f9hfLIQr8lLw0xWIPZXPzJHwe8QAootKsvl/SmIwI0VwbOC/Bo0oGUf4+Ti
RwzAnVN4Zk9q+T7lt7Y+Oz2kvRyv4yKDr/mFQ50Vwk7YY0NZUIypzcdOhBPKZQU9
0lomt/p0uEFZNBkn8+okT+ZuNLjIZ+CcVTmGbWIE7N5azfm2qQ3ZeKPNIxyK6VM7
Ib2D/4o9GXS8nzdgmV39h3J2vdVKpQHkuEAGba2RU4qNxW3IhviDv4kQAEaWm+85
uB2TrJsnmoxPvGIViXIyV7khyeJevisA60ql2WiTEeezTFDKfpHGODFU/f4Uyb9T
SCFgKU38Qpl3TilpjIMcbvo77Eqz8X+I3Rn36dcPDcEb/6QuimLg+9NYpc+pBRS2
dKGubJ5OkVjYBT6FwYiVq0xhbjUb7Edof63B4oFGV0Ha6WEnfy5BmPFDek4O6Z4c
vNmafno6vKB8JwG3GzmpZsFvrg2MuO6GX1Elfk7e7ovoRGOB7LtZadyYWiY7Alo8
Amtk8yH3zmKOEYPr4ipRtKx1R59UiH01G6VEle6kil0oINLIDkqGqUIvJz1WZa92
aqJKtu6ecyio6j5vqGSYDJpMJ43Ei1e34XKKHEp0lYmJEH0C7D0SZaBR0EYPsmBd
dFk/IC+upDQ1msKnnsL79E7mRrjRQhmdgdoWiou4IlbeRMYZBnFIQ0HEBTqfdqYz
oDCZ9tI24/o0a+UySOX6/Pr6phJB7ZRlrghGHjohJj7dxSB4Y2qNcs9JSfpdNcGz
lLJomqLSOuDQ+0TMlMBXavo5NYDk4b74iah0KJWGyyMgNamB/iCcieAhZpzylj7D
4Hz+f9+0m0h0atpwu0aElG/yBHHPdRVDyUmcM49ZWZbIAEux4SyUQuq3ZxRU+kxV
NCNYZsfKTGgypRiMx8RmUBl0cWl7cwE1E/mz9z/zf127hCX8ig7F4BID7ySuGF4k
5BANau91ej3ipOmctOtQDxh+7+aY6UmoMcB1D2pCXtCcSosC15At4/zfDtH12L+s
bzSTwXFjhISt4x+NHcuZaRhmK68hi3whfnlTpzoXTK0zXQlEdiBZObNwXxodWQow
+czAE3WRsIjmt1mlvnQrsTcbAv0E6b2avlqEGUHLqBrfjYyvQqvrHFJw/n4/W5BY
HB6cs0Q5hEgTimSAVX7o4g/t1acRAgo0PTrr3EJmoIndbBrPx5Id7cmtRn6WM8Bo
qaWh05kCZ5OA7mbnPcyMLRjGxry0vRLHMvBl8cqJ0qpoZ90pfOTIzkobeMvPdmKw
qk1ih7fL/NHThNyLMYUVP3I+o7G6ksZXaVJxCg20OC6yZOXAWK9LeVagd325mS1h
q7fbYYhEXkkIW30F5Jb2wy3Rme2C89VEa3OZ4iqsnanwuWTsd8g3nb3LFV7/q5sf
/5R4tpDnj0qGrlDB/OIp58f3YM3QGANZ5LbuJTeprmnquUjazH41ZcL6nqTxh8c4
DQJUElPojubJyi0N6cMDfUddmNLk1OYizNDNNdgaTuECjVh2BwYtquo0QhCu8mUY
gM5u8sOyDs6fHKmVy9k6h86njUQBXs3Q5EzSrsYsDC8l6N23/witEWNvJQpRUmRy
dYt+bNWVc4E6jM5ZhlsJGU99fH7icDen4aQnOAdUXGXtGuF1NS5DkoHV38QLYwrX
kK+wtnG3GTukwZmh/J34pCo72PcZ55ayd8LFUlmWQXvB1ouKN+3hg5GZn9XD3f8S
yUjTIzI3UDwzBJ+26tP8zVVtT+eBcF6aISaSo8+QC+L/b4pJcmxitQISZv6VoLgZ
ILda1SUW0hGAc1yhsZd8BViKrPFijjaEzryZJjH+ahH/fKYORRaWQSdFP4zhY+pi
AxUuMk80YmPApAAJqWH34ndqR8WcdueMlQdG7Fs8tkmaoLYDUDjzrkyHIkKGubqY
DCINnGBHuCEpCTKZnRzrZFL1OXlVVWHGBKYYskiARQ+JcT+i2NR3pS1WcInQ98oe
zKbtu0cL6nIwDF69XhvsMVwhP7+81YVUit0yGrpTwQtMaOJ98xRmn6159xymnzll
lsus+IrBNIEOACyYXD5dVdbJwi/sGMh494Phpf+bayyNj//Dqs522tt2kiM+49Hn
6N23ZyGQcsNUGAvWwVhi/ULc3wWJzv9i37ribI/pO2/hFcrlOWowsVKJigJDreAw
OnylbA3nSm2qGAkp9A2Nj52I0pMaFhjccpYRcdlnW4fnTIXlxNxLNsBgtkWOxF2F
W/VRIzjFskQnBl+09Y5NBoFxAHZd0Kb8sb3FVzzWs+pSy3pUBbIsGjFvDb2m5ayC
7pqQhqsCgUTHJQ8iHY8CwjodmVyoV85+SWJoGeCHXb/W5335vWVEnhmb5pQFJT71
AcU1nRnA1r2Sl83HgGO3o4i21WhxOD7XKDvjiNrz/0ZfklFAXkterCx4U/ziMgyG
7AS/AIv1o1ii1lrRqCO8rpvE0yq6YkzbbHPwZq9AB3HGgZfCMVFZ80JIaIc8oheR
lxLVm7BQ7MhJ9ZorhqxEBWf7GKFcyJB5g5xgGh9aEWQ824i/aYJiT9MUXB8xK+0l
Kt34MprQ2ffAyzu5hmPwV+XXW6euqVqPSzswKgmrLEhNf5fF4yrTfHaHTnWcBcKu
ftOzk6x0yRJDZpAT7jBSeyE40MX/BsfHV1rzGK2pMcte9+ikP3V65c8QUYj/PUt/
Ylwca/m0hyEcCwhFJGUk3M4BaoSQXbAaqUo0+osBah6yY8qBi5G2bLRSdeHWVjWg
9UmZd7/H1+yJbbBEZ/dt4GughDzjY6XBGtUi8gksQ2OmNy0D0kDZwgilVC7V/sO6
Wy+DCltc9Z0A6GTe1hUzSvBxuIQPfgS1p1wTl02chb/5OpTAdnVs/MW0qbS/fnrQ
3jpkF1MkPVABCV3YRpwEah/cOf7jikAiGCJw4Yh8NmMI8IYeJHFl6m3Cq/IyU2p7
z5Sx6xJHUaIZl1jbsvwTOtOnn05YIiDDaZ68QqQXhg+QFwaW2VQx4pR8p3ube3j1
W5QqXoqeQRd9yp34f5lSvxXhnFXegU0YECk11pz8ADJcbxXIB8lUroVNsOQWzhQV
6BFmV4CrbhBk+RJgQNXV9q2k7RzHDNpDXZbWQ248QOxJI/IWG8QKyFxHj2xvZnZv
hJSTlyRR3xAenda56LCotfCq/6Leh8hbe+eLDE/cra7vzjoUyAyPpi+PRqFzOB9V
lpzoQKiZjfue1Oj0LvKP4Cggb2xRQpA6ki8oF/ZF31ejHfA12hbd3mqDAmAYIHv+
VuHvvhuU6gB2sQMNx4x8RkTXxW1A4wFLlt3yqy69lcvdCIPArvq/LvZx/1YguV31
GPcwoKEsjCMcuIjFrZD6UjIUOA6RjUH2Rk3deR5UKLVSUdX4x4u0XFeoNov3D3hF
QTRtg438NO4WCTepOoQHCnt9YU2IgLFxcqFEzyxW/1i1tH94qNcWek3MVZzN1mn3
gDgz4/ajyYQweu/oEOJnRplic4u5C6ZrYe0gaasWvrkQC5jd6s+O/jrwqu40PxFu
EQTLgc2cEvUY8B+/W6GPzodEsEpXPKzsdZzRFye0ZByl7msNYZ6lbXpcRwoultsF
+CNVfBEb6ZpDfpvDKxx/O+EggrmBOIeiCFIP5FgeAE4dSbmnA4h0AnUgSsO+WEIz
Oei+dV9S87YE3alA+UZxPdlNQ3BUnrzDvqpjhTMX0a7ve6Sqd/QMyVsKnFVtAiCT
++oTHtdGJxB6kwlhvTfazd7RNaQYQC0SitMbmMsDcXAuhg8bpHsJO5uG7SYeRtO2
XvPfPsydzaIiJ3QJBZplk1f5uHP8XQhGAlfhBK1tunoLX3DNa9s7KTBD2es837V7
8qCXc+MBeKcpzoay9gS45xSLnANSN4k1/9geZ0zb1W4M8phiItqQ2fqboofjgxCV
3DDGQ49jsVfjd8lRFDbZOOqJTozlVHN6eYR/uSCts/WzqQw1YscYWpKa0QiXErYZ
6ygbhOk7gF6HkMpuxvRqwwU/+MMnSAr8U3NDMbTHZBXtRAoOHIQva73uGYeVZBCT
Ud5XYldkJy/K2PCm3julbLt8Mj4p6qrNOhpN0iQ5/Y2JjQGxOwSvUk+TDH7zrO3C
qTwsPGbE8vQfBBJB/iccyRhFFgaki1PwKcFxeIXp06m44oiQEUS5WP4sxKoX99Nw
X8+Tx+O4p5MGM/7r6iqrAFDOA4WVcWX/0cQNW4qu1Cd3DMjjglyja7EvQSH2OFny
EkhauADjHpSAbYrByvyNd22E9nWsCD+pWHnZ3hFr/AUbyCkGwc1nRvgPgD8E7oMq
5ZzA+ysa9gH1UJeUi0OpNexHhQjaSlfp354azB2wx8SeKyklvmFb+XileKiIcz6X
Fin2wBKmMhlcUYNCU0OtSgb6htCbZRnPsnNsxzE2Fcns8CTE+cWu0uri6bs9iB1V
6o4bWUa5XrxJlze4oXJ2PmAMdVlwffWUYxrAhRCL+Qnkbs0eRKES2qE1Q3cSiIm+
VqP0Is0tswRl/715zZhhA7YNE5PQYFBuMd6dn7IBHdnKrnkc4Nzz8StLONieYnX1
Tf5faXC8C8+8cUqmaUsVe380pisWP2A3nIT4oqPh/PbYNASFY/tpODpvh3xLuYsM
bB9GXKXEcqBd6dRNRDSbQLRQqo++nhgrZHXoLzCYBR5FSOin2CkHCBLvReoQit+3
a+pGwGC2cwNPr8vEi+RchpQ8IG+iKYjoeC20wEdKJMZxoxDW1BOtFXO/5BS80H72
+2b1EbZI8GUWMoSfXKVwTVON9uJUvm4rpjxBooq5VpUgtMhXXlDbzejoOfzV8ejm
PrEQDZwwtbcS4kk7W7lAnkoIOp4PnFqdlSyoafOF4z4KnegBVo6w4iCdBizWuyhA
/DV0SHGd4ZUFHdcvLWtSuS+GKQhiFbeRu9kUqp2ZuKZFVQxi+aJM1VWhJ9Bq83G9
ri8fUmkZ3ZjcAlzjJ9e7eoAF8YBySB3Vus1DQuRb8GZNdt5Ur20H0RBhIwjHKhRA
HMVFQ08LLeJLYqUXART5IgLBvTvH4xIh37URQLHNdFhxVwTMpzHKugbbNH8c1RZ5
1M73QdpIibQgOdAqiRlkb+/GLT21iPnYU8YhAhKg7am4r/odTw8Y+qi9IULNmXDd
4qxxGOAf9SFAV4Kihc0i5uQxQ4rrrtlTKdnrpuwBJLGg6B5E+FDsbTW+sZWXpk1m
lIC5tyfwJI7uOWcw8gurwB4Mgml/EyouJneNm0qhFHkAmmWJOqMuuwBG1ae+ijlv
Ihp4o0LC6K03f19BWy+AB3C3rl4HFzX0sLfSIzeL4t6GBjTKG4UyCDNELtq3rkSU
Mm6tn48ofOaq7iT/cdf+1qQ8VLdi1OMklW6d24TJbNUxDP6VpUvz3RFE5K+O7NyT
37VLi3aQRxVbsjt64wTOeC3xGiqIK5FBi7Bj5NGEpi69blM7hKZR0DWgiSUn1rdr
0UCVuoQBK1HTY+WcNGMdOdjgHYnh015LDZarsJbqykkbDWJ31APXJiybp0SF4qTX
IXaHH0IOa8FrI4D2EnCE3OkiJ+vsnYxws1t/RfKZ+QQO1l/j3/BtMGHKi1Ez40j/
aQ2GYN21wcDCPtIvm5jUvOVub/M3b1mJ2W6++QnUKJdl12g9Rbf6pGmy9MA2hl9v
3qXha5Y0VrPKAI4alWl19Kclf6haX+WqeYloQdBf3nNLtHTjM+GXrsLNHhZCfFEz
1or+q4RyrrNm+je0xJm98gZfYeHgGhPKeazTB3XUqvNtgN0BpEXK90RmCuMzLPrV
lXKV/KCkTR9I1TU9z+rvFYUsr4/KfOEWsmGLGbqoOzjadgWXv+b5umwYckizX7xQ
gpyCX3xNavo1dkY24EAXtam0ZDbhd7u+SlIIBlKL9HtgrrPPQQxL6IyKSXLq+F91
hOa1qgeRgQxZaoEjEpY+p7wHgnp8ZQI9HocA08xxqRosvS3taGfy7b0m1N1sujVX
DYTqrXItHHcf5VmLbD/UbEJ4bb0qLQA9TGuwX49a5OCKbwfo+sCJLEI0fMPoNOL6
/9zZ1TLQUzILQmp+P+3MXd13AUqU/DC+vApi0KAePd5SLRhbokM9wHgv6pw417Y/
LMAhL8VAY9GWDoFGJKCO9DV/9oBXWnRZu0dfihx0zC0tylcYeFCX7fXKRCSAxZuq
3Vbjg/9S9XRXkMQyvNCqIJ1QjyI4uTSowxZR3CuSVLplmilRmFd5ZL5XBAdzGv1J
ihr7FP67vQO1tTap9RYCtshZsHDDAbBOX9Z3gndC9ZfqKTIBj+1UWH0bv8pweiSr
6t+ayvwBaV8DuKwUGh4xmZZFSsdRGpfQMk5u/dCPgGXS2k4wxl72JajWKUeJMKed
KrmSvMhja4M0BzxD0h5zFmraG95qeIASiEG28YCqC6NFPQWfKSJRb68TD3ZWh7Wr
nGYY9UIZkg2ZrIkSGFznWUweNCBiTeVK3AuiVJ1NM/D1ziGBVrUwkRzWROeEU4mv
xB/6CWAdaMXUKRKLig/sztJeAJapM4eC8d9mFWNbgM7ksT6FMKLs15ersl7VCr5w
DutdSzUnN4zrHqbTUXWdsMErAFjZ0cERiD8vvjP62hvyyWsRguuyKap8f/Pbjmrs
00yg9ujNwZg+S9mk7x5AMy0BAZDrA/6QNVrQbekuA2Wg4zRfesBp19E+zQfg8ihC
7KhG6EeMI9FvCs0HUXgqH6k+97ysmhM0wC5abRRopPtbb1Dmg0is42o27l1+ZaGg
QEFWIitdI2PNmMlYbsCkgDW9Iz6abcZUm8GOp8/RlvK0Am+WgX+cm7GAxNvA8A87
ExPvWZ79cY03vdlQFT9lYmqhe4eSNyec545wHe0lQJJU/40YieNT98Xm6w4+sGG4
piD8imH7LjtbI8v+usMU//B12WCY/HoCo7BAYcdRckoCAazf3mJyETeb1ZG9EOYT
YzOAenWJsMzrdrjfMd4tOWOuqAmlveQi8u3daZ7ddqM4IDnZ/ofSQb8k1Izp3/O5
M3j0yvjPIgAwe3JNPhzjcmTaH5ghy4ZGtw6w+p9EgL6pz8L/JnCj5A8OQsbQDATK
2B0xJ77vN1r0mJg5yQaKXAVpOAy6c/6bRm0VI+mjdAAklgcTrNqCAK+4dkrJ/eWx
dDEAlyVbdeU1E5UdqT3ieCEe1wqKhCmki+N1mRpzqxCF+MXy1S1QQpJn2UtHKPzD
tmC9kKW+3rRKDq3gukpRqFuTrxNyWLH5b5AF+Glb8/+/eY1JeQiOguvPVzxn2vYV
5lvEs6grADUpen8p7eeg59UwoYHKG6/B11zo62eKuHuMuBScIZuzWDpJsYpmgmDg
WbaRcUHntCNfqOOUsyJ8WDC1kofQSk0I9dbU/bsELxDoVbeW2X7SqV7hOzni+/+R
2KmFlvh1AkdZmB6RksYDjDMp2/QQBnwBUN/mVsUfbfiFFfVj0BXDK0xwgXBndNDT
0B+Ln9Nn4OxmAbK/Y3B4QG0nvUWnLvMsLK5gb0iwmn8Hv2WLRha15d13Rd7hH5ba
BZN6rj3oapBN3J9h4TnzsT/7bbjXOPgUhXOV9BdKUzbmtBvO8acF3a+cytoGS3as
x0B0Vgml87JByZH9+90Kzvvrgp4PrGA/NupcoGzXHzT5FbjRLhO6NApoIkzzoDhw
Xe7u1cl6d/K2ps/gMvOs3csZEm7LFsbqina6CvYefvXm09yp9RJyIBk3WXwyb1hk
1vpn1NDvchO2HIJO7bPSYZD6D9MgPgjPqUuvmt1q5MjYgfyUERUUAC2VMDDVQHka
vNbPzf/ZDAeVDINn6TTnUnfKzmg4yvHaFnftbtWmFworFwX2Y7YqPu06qJEwdoot
/oDcHcPxwTjKHIbeYj46M4nIYVeXxotvKmznlv5MguhGA7jL70pIu6khBUgeHACi
18COJ/BUIGGxBamxCYjRb1UdXH042Ym1iD6TxEhJlDbiqyjsTo4SQX7pLhg4NlT2
1cMa+flOPJhK2+oYn4rIy9artGxOwY+QO/OHhQ0NIgHlznsnr58p0CaBSIz+FoTl
Hrc56yFkQZCxVVjqDn6YlccQ2VcfV6AyiCAz/y5m+YIUg1C3tyxMCGFE+Tzftycx
2PQEC0YUHEBbIB3+BzImO7nkXtJ+X9NHlYwmShyHoUDp0MEae3bs5k0Po9YNZh4m
HIYQO3eCEIim3O37J5kj2S6azUCtuyLtTVgsLVN3xGz4YIy4a30caHC10rlC1u7k
6AyQAU0zNuB0JGPQ85FXcLXpPFhxCa5CB1ibW9wkJ4jf/aL3XhSxIAszzWtsZM29
7y5pD1iHu+ja2w+9hQVgWJRd3MupTEqsiD97PVCNZUYcs2Ue6bXO5fMWBohczE+m
STwWCZ2/qPR2fmc0Zlc7oqImsqp2gtMxf4370td0BHugnacc7sw1q78S7mKYIwcQ
i/GRzsvfhhZrt318YpdLmQr01uQjxV+iyP9uLaGuc7SrCBmEuvf9PoGy3be7y6f9
XASo9B/9yJzmb10hC/eimJuyyJ8B3mHHzG3LAoW5bsnQA1JnskEgfzY4bRaKf+um
Y6Uq4rDby5psvYd26q8aS/hASxv5sXkr9rMBhPRoH2SrfhuPbbutU2jJED9SLpbv
2SGbwohZGdn2ZdXSuF/jA424V4B+3q6SfuEjz6litnLORAXxZTqfkSfqXWSkqJtq
l2SYqfNrn0uQ3vucohvYTpTiW1ia3jnDNJeql3cCwg9J7eJ6em/robtLHHo9fVis
OzHk8ov4JlUfqaYfd6WKpLggI/0Z4il8phLGDM9Gcxkw7xCo/pobyfeikIs80ruz
d9DgfsXvrluImVrjXrDgZu+/aTfb6sdh5HVtnxx3Q6SWi8XYaMNUGcf68Eg9ZtwN
l0ErI2KmQxSSYmy8lOkZhDVE7zUas3yAhTzhfTaJWH3GWbUdZoYhrhenWWnhaO6l
OuFyTPU9YD21Bh4Pf33RaljiC774OAbQjau35mItbLToK6cQl2XqYCd+Q61kONMV
qRR/9fZKQvFPaVAXSirNm5IqB4IhwCh/dLdvqPln1KK4FcX4RgbiK4BUFkKaTxjk
Tygrjdb2tqtmlZtDsLYsh2xxrg4cDBgBSs6wII51KlFYKND5yMO69X72yU1eZVKw
pX1pTIxH3xa9XxtAtswf5HyyGj/t+y8DaIsF+YnhC/SCkXjYtSvEd1cCDl2nqIUX
wM9uSna8d6E8uYcTHDWqDiBeWezqunK7efral1HgUXEgwZgrYi25UrN3a7y3f11l
qiJS5iFXzQag1L0i3+prvQT7YDZ4TkubTxAp0T+YLyc3vlh0wNRYxHRio2ZfBFW8
GBmKxOoMYo9/C5BDJ/xkCqyIpTWt9OOAxc4Nt4XOyuawuBxaAvLT5MzZN8iIa9nw
VUQrYAs7eV5AR6g0TgRykYFntIx+bUHh9fLeAnw0wDThVMN2oUcuzFEoi4j3TFIW
UarTjQgEB5V3wnWDwJI1KpBuTDpvHzKIKMgjrhhNHaYUYuoqps0BGWbiitBmly8u
TSfAK98uUsFeFymvLFQPtMG6huOkhScpmsAaTxaB/P9QFGGPB1/qDQ1xvCe94yOI
mlmc9exImQBQTjOyB/QLJEfsclAoXyx4npSHH3RUUmppQN11J7z1DOhXeu/FXBLT
5YjDSjUcYHxS0ZSbOBTNjX2dHbssadVEt5CkFl2PX8YGOf7YNDYebf3qiPvQMnsW
3lzLJliNVaXBFemJyFT1fdXwaJgaKalNj8IRLJjpOJX1wJmlbrGtKXPuNI8zWL2+
ChR1k/aZ1YVFDHu4dI6isuUFC0O4iRgs9P/meTfxKv4Y5YkByCRYe1H1AoQsETLY
aSyXXdLAP2P6g48jKc3lTgOyFOOy9x3dVM+N4DBnJOCRS9BePsrQKWAT0+yoyGKo
8M3jt5CaZKCYxzLTEX7dJ0cJuor5hTwIPcpU0b0x7Rwmj2E1OJ5X3+Zygir3K/op
TRECtZr6hnpEP4s3HZ0OAMjXWNjtiabqMbbWBR1EFrXeZB3BbrQHxHsv5qQGFUcg
Vqo5SsVoQdBnYT7FNE/63/G4xknOjGbLJzTDVXxV4qgEGn06jsl57EXZNgvwp8UN
UmeizXY5WrxlgsUBHByR1WQ1mAB8nmGOc09ZyB+zQXHE9EHA0U7KL94VbRpv8NoU
1jbkp+M56SBfDrxep2POk5X4BSJLKQaZ8A0BdVI6HumSunQUWP4QD4HqCpXY4zDu
z7U9lz+SBMJD4E48SKnSf0qUSEDYWfco8Edqisk2BXGWmJ0Aqkw8Mq6N3UWSbxhl
HvYZkQSk+TxjZDypuc6uBaSoI9p1gF5lyJiZYQJHWwZgR3QLkWaaGTuSZyzLxFMd
E/CDm0HGv3Gwhle3hZ+fRo0UBGsa/bL4v2wOEkbLYXe8jJpCIN+0tvpdKmI3bZra
NQv+pMXcnhSAVNLNb5nFI2h+zDhBH0kBROZBZDu5+A/QCzy98k6OGO5niKMGQZEx
Vv0d+w8+6zIGDgeZZVlKEvN8O0N9tEJTzbhoFNgTNLKNuIvvypJAEHYTbtXRMuMv
32aumlBy7yNEG5JVZ8dPM9Akzu4czmOuFvpX2jpuvPDxbNhAxMenFsiIVK9zYVns
4FV4irmDOKFCEm7eX3v6BW0/vz1OftT7TDeij+Lh68Y3Tr+5Lj5Q6NMLvkasa1FT
YAmOqZCHKrp/RHuhZ3mtz1OXTSISnlFvZGM5AT4k+McDDAWXLX2rzl+yaQ2j5XOK
qelO07t0i9QUgom5RDRw0Pt5NH3bD2IglYOWljmcxvhZjlfomixkmsznmfpOCW88
Q/x/T4UdBKJgdxV1E5yWEHfidSiM3sP6dKI289BA+JZ+HICkAyrElgfPrvciCBkx
HeypwTQkPss0pfVj/Fd1EmDvaug2ZmZkntppn6C603SqMcy6loQrcJqbJGRe5Pcx
HjVxf8bFXNzAS14Jah25mo9wSY0LmCStGt8a07d8g4SrtYxcKG8L56958Jd808Le
qseh49m6JeiCDl4zpKBClW72z8ilEO8cwSexz6fwYhgweb0Kv2JaGorio+oLZJ7L
e8fJSU+JXOXH3+f8mhI3DX1hFcN28Wgboh+6BCSLlWTw9tRVRGMBicCuw4ylSWlu
wLVdbDcUENep/i6+zy0Pwv37xpLNB3s5bKJTOPApY8FVbDNuNtxmlIiXm62TTbPK
0MoApGajF8NXuN+/XWpLM4sBo3NxWFbNLGW/9JHHZJR4TRlRoZMhZROJkcl8pHgq
8PcKe+ZkvY8xfxY/o7cp5NZ157RpSKIga4ZeDPcv9vzdReAo9MjAqKCs6OP23kuO
vepRAKxom6dTfzh8tBhYX3QvfGzaxEEzK176CgUuJ3o30mchPaF0wTsC/xspGWsB
szE2QbgLE9hKVvZSzTLE8yjZU1YuHdqIbZXmeUvq0TXqaLMvUj2rUfgJRKPv617y
apvHjSNGpT2KiV50Mn/xk6ACeZRpt4kql7z8I0IqnuhlrD6im7bshdbgzsteu1Uq
iGplLJB5NazdcdZU+NwVrGM1PuLSR4Gst3TlpkUXTWI97zjEa1O6Ochu6d4Y8VGb
LTDISpztmC3zq9+CMvXk5n3BnjnfEA0NGuevbfagceD67TT7bInFL7NR+QJEH3U5
g+ARJZ26xRKggZ9s4YjTzqQoWL/YSaa4On3rwpK0oQIOnjljglAITZE+6/9pAJnr
RGIe0Br7SkmSU7//fb20RnhPqde6B4q/43zJoPrGVP1zZRW56UPKSuA6Hyt73Px6
iEh7jclAXpY8JrH3PE1+e1rqPInorTCBGPlmGQ2UUCXXgdjTU9AGC1mDasktMD8/
Gb0gK7VJW+iDdel9of9RnKsjtCXaX1UERYzxujSKuv2ia8MBkNCmPWj7gAxYzyMQ
wCzzYwcypOaa6WvFhBXmO2GdGP0v3m3M/KZ6pkPgeY7UmkMshdenrn/yYAemfXTU
id1ZTyaQtxEZuQ0LzeOr1MrIeF23FgIODmlMYvSQ6fRBETUBHgtgfBl7vDv75I1F
gy2LXZOdk46wLJpr0FmliwaTu8S1w7VLlGzkI/fcTFy2iv051uMXiRJPgl9I3u+l
Vfxo3Ld/CCoGUJlfbA1HtzbU5kkbR0M3KRQ3UcIG79KubE+/iW7Va9/dXFKD94VD
6MGe/jxaszTeRZ/rhll7+OTQOh4ta2JUQG/e2FCxOnLDINVtABnETANOs+lWMWtV
xNXIBuJS9PDI5iSbQQAFdW4JVWPe1ClvStxPloOxl1ShQ8SGug6nTCsENzsGA4Bq
wjZROInx8b3NeatmggOfBTOVgLEE8hGcrDT+CFYNvcZUTHf79oz/qur62cCeDMkI
7p8cfisQqWsjsFFUL7/EpDEAUlGjAwHsn8XoErCKA/vLvgilwjW7XDnL6GkU9oX6
vJTE6SmpKzMznDFSByPdZ1oMdqIPdqp5+7vcHLf+wesiP6fntqmUvH+CX0iyHn6g
bKQCbpP5DTInw/1/gfQTU5L66c+IAXbOS+NJR8vlQ6og7BhWLuNhPd9K1oyHmcqM
/UoN2KdPB8KncxTuN7nTEJ9vGg3azaFHDZFYLVhK0uX2va1t71q5BMOEP6ogP6ig
57ICmGQdUBi/wRnqMur9zCW9dalrHMhn49KFYJSOqOuXpsa1SEf1OB/2jHgqdJLV
qxjix0gjRQs1Od7skzPiGJmjB5nDBtCVgksIh3tRjlbcesRP2+9zItQ1hiMiT+wI
+C6H/kVnK+PFCIvFCko1SIahodrAx40eGbzKwP5K5/AUvjdgMVGwu01qxYkucADI
P8DNgAZ/pHa3blz9hmeEoTBFWxUR8LBO0IY03jj4KeWkk3+G8/hF7w585NFHjd2m
rlRHwkcCEi/wPFK2vbMdisgorLiaFOVNdBJoPD2yiKlQbV59V4uBHHg+OcqOaLgc
p1rjHq16yq/2AWhrEz5sVkqlUluwARPyIlfRmlPbhjyVn9rNpI6caSNGpl4O7ZjW
XrKaxnOnD26lTo74L+M1Tu37enn5Ob8ewqiK2ZuTJPNCJrBo7jAfJhPhd3t3umlW
xkzjUvbF5Y3oY0C8Eg9ulAasMBpUf2oyY2poM6gaE8hhxg75Z01c6G3EGReIcZA3
fRcmzB+wBJ3L+oJRpvtUpLSjXOmWhcrVt4MbsZcyAya0kXj0GuEmEjCFH2g+Uw8B
CaNRKZo1yIgCjVrmwhFewv4Es0fAX1tChtJed5KZ0fwB1eyoPsr3JkJn0uqssubq
QTMej+2NP+FbBI2XYDXT8GwDdsGw6vQ7rhJSuRtJAowrQ3N/26JclSpr+Zh64vRS
90oIZNhAN3pDPDMi125A9EVpdBBSuhfAKEo4CBimgOXSyrq9CZa+QrInt5W9Qmpi
xZ86DWH1k3fhcfsElc3Z2t9RvBYoPOV4xgGHWQF4/oMLaWr2sxXh0X/37JfW69CY
ADFFPEZtgQposoJwDy07Zswg3Xl0fQkyvBbfH+EaKMq1siB+kqSuo54iaJPLinPa
+0FvzlgSM4up8qYETA3g9+eG3DdPSMru0AXldOUZ2mfloO/GOZ2jP5riEZHgy1wh
qW3EQs6j8tMeiVLxCE+B6ABdBBp+MEcY5SeYK/VYSDjfKZ4s9MqGzlKWrdS3jQ6b
ILEh6+qURcJ2JZ/lSDAuT3vLNbO5lQE/uTveEakeh34CLacsM6CmK14Ogd5L2FsZ
yY9TAoLlACyv2eacfMUtazRU5LOzADUPeeJfXJr0Lk8uo4LjwZgMkafCvt8qXbff
KeOZDF2LYEs9r8muTWuvLXdoj9D5Pplf56sX4vZXoIP2/5A+KcNp+Rdn7wySv3VA
RTvZWWJsvwfHdGLrAAygArLsdqKEVcq8oPb2jdrEDmVYLb3fOKnhGBUFkYSDXZFM
l4CvJXKfVAdD6wbNBVXxgXMc1lKPkYj2nRVCWX9k5ORkPziC/okphvJeewXILiy7
ZcLCmyYSuj3WWIkgiAsHxQuPhpoCctZMCXPaiNLjwMCVWEWlvqSglo1i9ZhAatCJ
nJj55DjcHtmdkVylqmSMdstwGIE43F/rwVx8MooMzy0Cgc8wwIX3//c2wr6QpQoy
aNqyZMPv4QUb7nmwIaEV9h9OGnZIUxhZxK0n2cR+QCJsTOFfAr4CzREs5yt1jCjz
ctCpfKxGJ4TenraTz4a9qSPKq6hq/933nM2i5yFOSRv3/tuXWXPfpuXVaZYO3NnG
My2bX6g/O+JEzPBpfZ5gX92Y3A+NxFK5KYjyuyLf0eUKNJEw0FPfajo+5SkC7E6x
SjrdUOf41dpSgI0lZ7nuxbTChrFA32z8adVlnV1RXELq6IvqaIyUJT0VfQBDIkvR
FoqdwX+Blc0j+ZiMcvfjm2KFtotwt3HR7OALWlw/yq+Dwl077heMO2EAZZktofyX
wjyb/y5FD/jUAhmmIWROWWDRJMZGbzOgmQ2dXBQnZpD4Lev06f4lWMEAIm3h6TMK
HdanHdddRKT+9O1AhqvjfoyRKEEb76Vafgg8kFcDFmzw8V48a94wYV0XI3SDLJEl
bOwuGCuuQgKkdW5jtwpUeWua1K94129bRYJuZXd8c3NC/TxNrvVtahRKbIe5oaoz
X/6L7Lqbp/G6Qs3ZeG8oloyYfvglTHtb3XcOGlmLNOhWw7aSKoJG1NnPZk4VnM02
GiQduW9on4QBD+6U2VBTaMibwz+LP9X7TYp+r3s7JdpA16zNtXAHJ7C1qwyYMBDJ
Cm+3GePcAbjBDKaf4DyLAm0hJX+RCGm5I9h+WJdGB4pifpS9ykeRxRszrXZ/UKQE
CfZ4gom1g1fUTdv1jhBmj3F1TJuxuSvRA2mi9v8kreycCbFUry0BRMY+YaUNA4ir
2Lfdm3R6lUJLxutwVh8jhwsgrH10se31og4xiIxxoiYlvIOrKwhFVOJLh4VEFI8P
VQ/5ePRQ7S8v+u6OANxf3WGpUzuyEn6YGZaEExO6sWRHyrm5Kgc94dc844zzwmlg
TyHd1GaTf3HiEsk9zvgmeH5TZGpFxzS1/g4nbgsKgp1+Fy++AR0Zrpsubv/ok7ZW
8xbdBbeexHgU29DHzjIEN+oB8V5G3omJVgh0rJx9eDmMiJJi4hqhji0lnbKR7kFc
Vjd1RmZuXWLBCxfsNuy9gX5+2R4APFr6KTUBYsWWOuiq8WEJgpDrc8yJuBGy3PqE
w8bWm/4TnxX7Eer/14qihUWVbrtrHFg1zAlxNJRiDKxu8xMKt+4flmbFkf3y0WYV
NFp2WwYimIbNnX933X4L+2Ypf/ZW5EqSPLFNXJIBNx1YE5uyLS7NVVsRrj506dx8
/64+1vukVBmKDtClYdewTopYKeiwu0idRGmHw6842hqGCN8rNoOvD/gE70G65quG
ZSD9l5Yst0MEVlFVyaZD6ioyGxb6ql5Ss0EVbHWDsUkHLYLhXfYh3Uv+lSZGfNM+
tb+lTXqU3kXybXkrpy1WqxfV3B/doqa7ickUQs2HvG9jJesFlr3dx0vfffjqlzav
W9pyiMw0eelDvE9JIwxlq/qINTQ9YWFO1jXi25PlfAFAQ/kZOZ41HbzJl4Yh7PTq
WPSaawyLt2e9ZmGC7mIkv0mK8JwU668PA2YCyi1X+CxMqwF5uoNZYR6V/6fczCTI
GRWjSzszLKpUXEPJZ4obGLC+RMQEipftipQxdZ9DF3WSMNFcWlOwmNtWRvkmsRne
HuYIrPtFSYCL0EpfXa3HWf3QKaQC6JT0x8JGNPfwnlTt15ldVmTpMsuWdzTFawHN
WGc4Lj2tNUiDUvUOLa1vp2c9RuTFTOgQ9G2fcV+1+GNfwh6KWtn5HKuhf8aAt0A5
h0dGgRMg3ua1DEpJ+XsRm7m2CyHJA3uACZIKBMVJWIy0DSC+FX1zNu0WidxSBfnI
Qvfqwc5LPuGMqyAfiwC6Kxq+VyfGYvf2kf3kKV2OG0k/EpFeMhuACZoxuLiJiGX1
75VZnlpNepUat/JS1guNPPkOVGItNZ+Edp9IdFLaRUaRpbT+dAViBw68jxzl4V7M
AoNKcN9Qg3YlgMWH70s2bN0FG5ut5LZWwfqGfijyUNhCgoIH+B4IpCU4DUwN4yVw
iRfCFL6j30plUTSgLs+mqFUqdfjpWexyjVUR3BRcqWUCRkVG+/6OJa6vcBHYrude
hyWIXRA1w7TAbrrb2eyD1FwTr2q1UCd91KivoBs3VqG7UE3SwlAT5Ik0kkIriojg
iq+/oyKLlQyFp1i0ODL1axgbAvF19BQ67V2rhkJ82gZ40/h1osoo7fnL2guxLNsT
3uOh9fRL1XV7IPMVa7dRobvMMrltDDd/6v1Dl4yxmOx231723x0koUJSTGMeHh4W
oT61HelS+adoUqSrdx1VeXcz3P2vhNsjX75Q/O20C9nKaXduMhY5rm4zfcFaFby2
FbMT7PhRpSM5F+FQhy8VS2W+9GYvgtSs3yd6K+xr5SiYAxdTXoUs5iu2QmuXEuoY
VVqrUymjnwIvlmaFHn2ttWbWdU2V18sM+EkxVM3FCuu/VaN4KDUyL9B2q/LybqEE
1qP9EtxOEU9BWEILfbUXoWPoZNFuidRlFJsYlk/cB2WtW0r0gAjQBSK6gcKH+KMf
EwVjh+vNFAS5uksKSGXiRz9+DTUmec6UsXa2+nmedNb58nkjxJGKzgSXlii8gGpm
FSDDeDPYaKEKbhEXMfzaCFgreKx2FWiZ9EFG1U5/8RjHPaInrFb9CE0YZXCrKWM9
Mrgyq6ZLeo8QkWLJzmyuGc4vR3SylYtghdBp6c2Q0TH7NWPb3eijecFRhtYbEqYI
EZzQx+MZPzSXpJkoGGun8/aksKpjdIunPVxNdWif+2W2R7uP5H5us39xHLeTZuq9
vNvI9Q0Tw9M2yU3hGe9M1SWAoBIU+e3aeOOMIOvTR6CSSrJ9VmIgXKNNKm5Wak0F
k/W5oD5VYl2R2ZR77tZ17qKNlfv1oCEh3h6d57WEag4PX3Ir6cb3/JekWzBuREmx
Mj9Gh3xpgmiGUhxmlbeDNg3P0ijPOAxzLbachCLTq6t/NDLl/abL/l+4KQ/Nl74f
joBacsOaMMY9zickkaamWyA+FEtbA/P5oBShN37hv0IILPIDycgcAxF7lu0KWfTW
ESiFqnLYgVhStt9W5rnkNLuud1yR2fgtSJFl+4pws1HzKTWH/KBcR0U1zsSwp8f1
xS+ift/k2PUCZ0n1TJRArJd7zw22+jiX9YPBFEF45rTH3hK2vHw5bcfYJw5YcLYH
xmc2oYnLWjN0darIvnib4roL5ifxbX6CjObeULHiG6URaRBqQS6gQCUS43lC2MYw
26r+G818gzafVCk+JGWMPopK3T/OJSCO5+kk8+uXwQhE0WBaJi93an8ePOxkX5m1
fo1LjwWBMUkWRi+44XaEtXtvvHv7lPBwkdkPrTN42/GP/itg35zhZXVXJRU78GGN
Z9qN7vRE/n758B22r6KPWY+01K4PdGDI1zUfx3g9dqonCE17loWzqmwibqOXuGCJ
w8mrNgZLzyp/4rWL9su/GNYcX0UU/FABHUR/1GNxDQi3ipwLkS1JnU3MQNfhbJ42
eHYjw6DPsZ8QqQxhv/AXG4cjogp3oGrgYOVoeCIUxy07yYRkVDXZVus8sWvsYtpf
3ZdwYpulBEU9v0uqEPyKU4LEcq+IYAPIFNpEHFfNiUi0ITtZb9JasMOx6YiN9zDp
zH/lM8MP3Pg3GRQ5CxSkT4Foi+/16UgwvfQ4gVTNX9JyccBNUh7LcfvbVbowaWeW
1BpJ12zCZNe9ZhVB2FjrahSRr5HMeF9m3H5CWKHzBIbTvTBCLp++IkrA4NOvqWBD
g28ZWSRBL/Iz0tFwi6UQSzkLRtlX03Qz8I6+Vo3MNYjqL0jG/agqW4GJfm1rPWKR
0iCYaV/J4rU5450R5Zhn5l42ryXzfXTeapRRqo/7QmHm3KWZWjVnPRuLMaeZzqW0
EM4MHGJgBralGO6p0PO0oRJOsSWTZwYL09HSn+HLoGRczknrX04tl3LEHby/Wd0O
A1cHGSAFi0G8P6QRjDu/gvpAdc1WPjloaZvmY9VOlIPfzrkcAU3GMgjtmsQNAkNY
og9i062rX6FvyMrK2RKz+JhiL2+FhHDw8F7A2eAeIrcObgelNaNmWl7BilTRJTbu
/HytAoDZRRfFqamOPIvTtHaU3nZ83zkvaLJAymLLGWjUmqaJwT9e1yO8kj1vFaiQ
l3UbxGVF5HU9xetbJoFhxE/N4clx/gOhgaJ/EZVocRWt1JWUR/TlsijLntWePHpY
CmPxWWn6cYp22BdhDQpjLeiUegnXRCJ7a8RFgce8GcVUTrWneFHgO889cLClokA6
Asa9YMh7ufJBU+fOL4vI/ehIDXh1VLCEw38rwop7D6rEDRItbGCcpGEjCygpO+2w
sU6b58ntQeOlm6g/8z41UnbzjKPib6WbPkAePfAgqm3UybCabFm+fkYEcsv4FdJM
gbYwOmir09LGy4aZzQY09M8dtPhvsETBc5YKm/ifrCpJ+pJI2ratcEKPk6P5XWuO
xx1LkVX8ZMxtABeA4xrXF9oJIqDsFguMg8Biaufv20KOlYSemwujBXFOAMHrbAyk
RNW4hllCWN0RBk021M/ji8aeahpx4+GujfglY7x5KVe/1aOJq9dDhZ4PL/B545l0
TNsOkNHJzSpaRA9Hls6HEsOGAV0bMxErIEjQqT/1oF9jAqDCuF8fbJMcw88L7RQZ
gpv3DmtecQzKPr17W3DQaIUb0xrnCGpFdiYqFmqF6Ti1TuxOgaYMRsuMAGgzM2Yg
jqIP18jVe8C6+2no73WxMrS9VsU4m7IvKTUBGj0RztPm8MyXE0SZDE5ZBHi3W5Hg
xAWu44kLxYgrLDZ71uW7t+Da9iAAW50t1RU0qGt2RE9JauhVN9nZdwrlnlCrVA1r
vt3g8cI6oh17hpvOYwVodJ8TceMHXVgviCECh9B1he9nZAPvf6uEVtKUQ12cHRSx
1b5t83ZHLptcLcN9XTEpQG836pysDfPb37B2M0bU4Ic6UD9mEcVysBhfszzOUcTy
zYTsGh8qPvqn0N9FTgx3rxGza8kIptNwr9APkmg34WlnbnLsJXQLa0BwvrvvYSIV
CPoks0HritmUjvxKb5wVz8lyDCy5XIIRXgTHAY04NYr3DSOJ247RoPCeztbgLE1D
R8n9GR+cmw49YO4pp5MyvomtWZlURWG6Q8byRGI41tXVngMuKR5ddvNWzO3IIUhF
+J9ufj1Xf4L3rHGRg29mot31WYEcsxnUc2g5KhOQCTGCgD0TamZRYdFDiifD8qT+
B2ayhftFryFo+bAhP4uDECSa4kRNgXuGHIgf2P1FxmbkqHKeJZKpbuX9zosx3XlT
NXjwLUrqyqROJsWCBDKkM+NT2hi4bHvDBDR0AHUPjsHWPcqu6EFvVqDSLKo0Dnfu
nF+VDAy9G3prxniOO5PfaHEFUheu9Q5kSxlGMhMv3K0/gYaqRV4oo03QQmtfzpvc
an03jHUrT5SzEGzhTc0piN2hysh+l3erND/WLlZ1pOHebEYsEih4gXk8g0WoKL1/
JRkdWG1JhSIq9ZdkNiyCAUAQ/xg7EQaDJHRsxekPYMTSomoNoTYFlpPKc7kwsXoR
DMHu0JxfZ+PlEMwabuoicCnP5n4eKIXWLtpzXLUlzu4qOa8Z2BZ0+E+hAE3kRqlx
52gxeV+1bC5H4zgkyf8Zz+AqhSswBYAsA/8jAbSmRHfrydTUFLNlujj1cta1kreg
vQu37ewdIPtdVMYG6V2nDHetAMBTDtr8/7iFzBceGs8UzMPu0pWIIgUKCS0osutP
w25snq1AqDQLNwVB0y91c9J6HFEXWZQCbzf7c14e+vExHh5Xz1vgOMGfI6MviKnZ
xgzBLCe55lLBv2LnY2/gSscCc2tJrugol2SAWumSr2EAx5/YLR+pUws4PwhX9AG+
uqVMIMJUmRzLBh0FfLj0wvck/njzp6uXIutjnXGLuBA2qAt8S6D5t6ha5AXD9biB
6Q2XznciBNR/YpVc5VlPVW7VNd3kMxP6hgb0lhdrxpSgBtdtkxDY70z4MR5I7DeV
iqXL207nQAP94ljtS0uAakcPi0axiTTgsPuQjx/32BOp4Ok4TLypv8V1mtA2C9Qu
FNkWHmBUda8bGrrRI7Ww41kMUdcGLRjGcXKEGpk+qgLDDFro6LedDnQkJCqcK1mK
tLhvolC048LH/3sPZzG9KeU9pZ4W1TdgUVrDom/peNK/ticSccU5RdXjaS/e+w4o
t3pSD3t4+qGlXgbCf5C7/O89JDB+mtv+r4filLzYugkRu368pQE5nlIYYS2DcnE9
yEET/+HgQe+MPkF0AYK59LYcOJMJCbQC24iCI1lfbA62PZdYP4zgacu4Oe2EsUoX
ke96kRXAq5I3rNc/Y3OpzbSDbEaqkGgpt5xVvMerhYnqUeFIJziGdar2us1cv0RE
mxL24+FsU0m2HOoX+lpWdXIadFUu11/RpZcj9zKvh+ko42WD8MPdGo2nJ8ounn1E
emWnKjx7/k52CYip60Dc3jiLBhW6lBv9aAGVjTxBtsmvaJZ4hYL8FjpMJrZ2ilZH
16y22KJp8PzAVNSBmgQui7AA+Z13KjZ6w0qUbOkxymUkMkRkKz+VppY9B9Fos4FK
Cn8dmUndRlXLqpMtWMhh/k5K7di1lexd+3raUSycJg7Q21N5hLx/EYhzkIwUaiPt
eIyl92SaTjV33VZFaXt1zcENFCIyiaWm7IUHBs+ZNz2ilUzXcvCccOxhsprop/C8
HrHTkjD79cWnglWz2xABRIDytGp2aeUn+X/Loq7XIZISVw4AD+y9CxYlAUZtXn5U
c4a1e+zbajYAM7dcv/dSgeDps1wkb/t74i2EQ+pfeEG/4bEd6FgG2EM73ZR9jWpj
W5YACl1ijUhPFOY7DSB3i3HaR+vuLTXdf+boStQId7odfDK5/ihjWTlpYP9WEq2y
AWG5UAKjqsBpRf9e7L8B2xhTS1HGiBw7m787lYdU52pQZYYxIx5LRWqjkhmct0my
SZmmtRpay6E15UuzGZTbGhjO91BttDu/jOWKIKcXvH729ZzLKcrH0wtx9zW7XqKc
ANrgW5FJOZrNkchDuhxtExq9qqA4VoD54iIywIGY1WiEhBhGsksJuhuA/PkD1784
cv5ENqeNcJjIA2pZ/OOmsenxI9xTRnEZvsjvPG3neJv8Jh41xWksANo+wg4qEJWO
aJxDOscObftw6vRc1sg4q/CpCT1koMZCaRdm3iehFMsqYLWPxXQyqkc2dBpwewmo
Zf8AuKirzEfHYhmOJ7jpouKM8vAK6g0RODMcqSLrbX/iggYHMkzPeMfzHuRnzc05
uzpyXk6BNoEAH0iCKYa0WFKmc2m36HQgzLfHaGRzAXV6D0q3F/a2tNLLhrHsOVGJ
qm3IEG8sRr0A+e7iphShkbLG2A+f3cSElUHfGYTXIta6KcIifGQHwKZixcF2gps2
DCPsVLQFc9fM/8jwo52X4gt++U016j5j+4zB6ey6DROsF7V36Z6dltYOsXTxn7sv
SGmDxiilmt7vpC78NU5BNxEmsAB5X3ZJamgQlAJ6BwBILx1psrQ4EhKL+mL69fkd
xZ8waSLdyQ5q3gCJ96FMRrhvONp6yCzbW/v6t16obSEuJ6qj42hxpDBeNu2+7Wyl
PiRN9ek9M0yi3FBfqmXkMEmaK8iMsNApkLy7HAf3TURwwej8iahX0FdsAx4hMLGg
h/cUQFwyC+syUUOJExL9o8t4ROW9EOyWnIQBId9/8Y5kEV4y2v+GQzzON1vRILcw
ziuRUClc3BqsAKkc5SCciLDlXHrNfm8unJq1dReKjLbHxok52/H2erNEWNsOARC8
zQ+4UnG8gvmEBVy3ydJr2co78ElOCAlIK6eapHLDfD7V7A1LMUz9hKGiY0kf5VzO
p9x5dn/4ud52fs0wKbpHmUDc41TMDBjRouybvhH1rBmR6dbKx3xpqlHq9wAgJr2+
2yTncZV2LPSHQRonCKKx6P2/zsd58660zGntRElDhLEtrBTaZGdiAjwRCHpsJmXp
PHRulrvsdquDTbPzTqhGRDQtpx10gdXfNo7+ucPWQcXV74ih10WiuTz8062KAhh1
N+1ZEAMi8p3B1nPrrxkLtMTv11GJnWHnLcjgnfUPkftioU4rbZBjPXtIlvV/i+Yo
YfA/mC4CNxFGMw0EH1F4jElqVhmtkPHy5WlRRvX6OGg2j+sAHqgiS55vxl2EgMLo
LfE5c3yjyWC01BkkkLhegAVceJARfQX+Qcpd7jwcLhe8MuqBq6mtevgC+6Xr9Moa
hGZT8QQdNCdVX0O8Gor4RoIb5+SgkdAzSklP5bY1l4+DYMbHEXZZjL1d8yoXm54O
5Gys7UatfIhIDuu1EwUeK77f1wizobqMMPwfTF/bsX3wC2zUig7oq4g1tb6blCvQ
y5dSI4Fm3GvKfl5cStnwJWqBDgg9hjI4qXgaOdbti50zdpLfT0I5mOEwGpM6pcmI
dRlOu68saO8bMzna4/cfaGzbhN28pSRkqvCe1W7IMKli8nZKMU/NaBKMjNw5bzok
M/gL/POwOox8f/XXVZE0SP+QzDfZetKyZByaUwkQ53G+vsyWczWDNI9YJ1D7sWim
96Pvc2X3AkVo88avQl/WE2EMTJ11UpZ/pdBEI28DZgoY6qbZSFQeSDZGh23vgQPA
2OMBXRqKzJXhQQ0Lcevjm7i15f7H7vepmiMvx90SEqe6suUaoAe8r4FnYpSDIZja
jQMo+AuI22MLJBqpUd1oDA1sRIMloGOFxup3pTg4rQ+lnG5GgGM2k9erKWY1FrZq
Z7F2gjmgY/dCqc3kQjD94xmsJ2kYZnHvGxpcj6RinD0PAHJBwrf0gL6ybpuH8/N5
B9dyyaSUjarYVJWIW/rxGdJVVniEbO03fmi08jOSCOp1SF23uKISgDJMoIboE3Ce
KAgQgV7JPTl4AAL/I6Uz7fua1GXylXr2CnikLpjtdNtlntv+DLN27Xnnj253oPKH
cgjpb24+3/nxfDVkdIHa5fAXraSr6rCfkddYbwFkQEVG8s+gNH61Gkx9hYJNkMrC
9dkL+iWvY8mIATHOSh+ENVi4WFTRYaoIV8fIVVaMA1JliC3CIbtstU9QDQUbwq8q
a4SW2GbUfgnNI5o24WCHPvqnHSKE+aIG4qWoq0b/8t/0kNceQKm0fpOESPMxUR12
su24h37lhbqr+J6M/zwEzhj13V+7uFgKKae4RQki4+rS8EP619WjsdHTIaJOMmbd
JIbtPgclYLk2LQtM9l5JWLJ1o38XD6YzQw9O0q3CCzhbJuTC0Y3JKiyy++ffkOaR
/UT02kLmUsa+Hg19DBrI0XxUR2lxh9Rno2Aa0eFsqzHa1zgfuz90VmmuWrnz00hn
pAQwOQ5596SXTXEgPlIjdnaf2bdy0JkWICnIAc1qEHE8qww1sB1j8BvszRVq2Kni
S1gLynHUmZOheM82KV6m5ng4KM0IDm3Q0IMrOo828b84IxG5p+plipPUkRca2hU1
//9Yl9yWmRLC2anh04ansBFM4Y13KuZanvuTCj27qkC5qXbSFwE4zV/sUP349XAO
HCkKRuEO9XsX0Xd0qryul9CequGVvLj/6bni8mGpv1w5IqPUsaHCflDgkhbsMR1p
VxsgI/+jLa3ooegXyfRe/+A/RkCSUY2BYG9b1Bm8UR1iZbS8mkW4RTa3PcEDixpj
GhyRx5txdJcovdAOqtnPy2t8B8osHbUnbIFnjAo7hQwtsgt12KxmMp4uyK/6r6ik
moF/j8N9KW6LGhXfsSa5EBP6yBbGRzeCi7hoHKAPRNWEkyZkQ0FCeWBczWBJLNRm
hh3uY+gx6DI4Th/cG0z67B3EpDpMu/xVM3XddhllTZ0iHfau4w539a7/wilTmEML
5UgMr0FSJeYYua/8VkHSV2wc5C7lGyEWb00UWFTuoy9FjmUB2N+L76rHGy07CytV
isvX+8g6vGQXQvM7YeFFwkcCFTvT0VN5cB8oxjqdDjKGcLSq5R+mtp6ZwJY2Y03+
aK7qS9ZjvYStcl5H8UFyyG1//r3oRqBocQGBZcsMtHgs+nyjC1g+nS6yPOiZGWjn
MBnymBZyQXnGl+vj0zyri7lPdl6vsO+vJpybHzQAnA66Znu7dHR3zt7ezljDk0M0
Qs9D/smwfMtN3NSWAHx5mw7DneDP02fZm5HrqW/AkKwamGh9/07HjRHNNriKshqo
+W1hD7zQR2mHSJIFlftFQiehr+jpM9KscadhWNkBtH1fDEIF6rWOxJlJeLlQC/h6
jRQahSvwKGZilkuA/OGLWkNhj/QPDU0ndpw77xDD+Yge7Woh9yy8uorsUrgaB6HW
BPyFDNatvadVBS51zuK2cYryFqQ5iPd2PplZxAYz0IW/GVAL+AQUi5d+fEcV37/v
QnikJynO2jGMCnB39thSimlfytB6ehXzE65upP9FC4efs10D0ZuRNbQvjQy9P8pg
73FFeTonzdVY/Ic8LSQnYdH94RXtylMT6QKW10CA36RRmvYyPL3nlpEBL5CbQZWo
XnqPOp3rdQP7ISM/Op7NyXTzMP5H3yfx/7UUOe/mOaIVjDPgb3wdFV4Pso4m5WYe
QbT+WFbMhACLelWd1Dnx16QZ+IKfFg8/oElHcmSfxSiLE67ll9NsmaZGFlFiBWvi
rVTPnTGfPg7laF8WK6on5HBcXl+2DioowHk9fKbNklLVpvsnuUDefArk69TiHcQU
CwIjLxNjBNBxdzAnVrFVlyfEsTNcp0HXU+eRlz7FQxFFvdBOAYLQeepnAECMk19Y
U0hEVUYcxp44PH196iWk7FUiAn3RokmTfa+cRei0Fn7QmA3io47UXF1tIFMA/qrx
tSEOlTGt1qWu2AaixC8OdiMxN9GL2Ph3bkOpVNQvUIAvEBd+6vR96isdTpbdf6qn
DZONeWnU7RWz7OSNUASVTriHqyJcRFapJj4WOW71nIljaNBerqXALrGiV1VfeIrj
w1ING73WRaQaJNm/sGRDfPQ/1JziFxEPf1Cm8ZYUjXCzxRBBDgVzJZN5d3SvSucQ
7P00+R8CwU7ukNBe9TdF7wnQq4R49RKNk4VysaDRciJeOAp6IAtNUHOdYX6Fei4r
j0dtt5qfVlbEcGN/M1Mee3iHP3CA3lbf7DCUEW7G23jP2BA6UPTfwv1QvFwC6/rY
H86MNfGjCl0mXs5OUPEbeSTQRYzDqCc0OcxCAUyDsPvr34HiTgJoa7wx0Gqk68n6
qvOvPJstNQtBnAUec1UkulIoJFiNyihMEF7ECPKmDKErraACTWxmfYcdMzflO6MM
qnHZ3/yy1kAE35VLJd7J0lmMN3HqaZ1hS9X8LQ2xDx57tsGlnlBi/HoL2Wx20b8/
yUd86XQwa/7N0epdicJX+ZNbLa77PBS1FFUA3q3r4nRqsqaJUJbX1NvSGz0wwhLU
gVdW50ob74ETMeENM9Y2BDOBnXGLsSxgtWxd7GgluclAKu6aL3iGd/w4aV7U7YA1
b12AN/vfam7WnyF4KHfh9mWO/oneaLrWq3518E7nUYs1WRaToOauR97RRyqurAnr
uXekFlNQPrXbOpDDo4lrUNArKkxednonDcY59P4RBTcrWV6XX6vZBRrTbx3lN21U
wVvxeLnhrF0bMDNkqgQU2M2dmBv3cM81hsah+UnQwNhaJ8sdPhmyLncfdGCBjro3
nXLdmD/TiZ4dEqIBGWnlbf/h1c6kiblxzmYpd/HZu29oo66vhlCINgfN+IsqW2bm
zzYm5lKZrkkCQzpLPx8gxHRiX9hW8OpdHCPmPXFrUeIsy0IEVgnTFsd/skqgjrvV
KC705cqapXfhqaXykBwJsebGlrMDlw3Y/fDx/MGKC8RB1JlZtaZ+Ld9GWrDb3+E7
1/FFhr+yi3f0xHw7u/rRUkJYI+Mcq9ZvQHW0snCUd5PCcyG8j5lXiDqlZnFckoZc
bgam0RhrwHYQTipnAgk2WIgcZLf/JrTG/fErkOS3la8NUWHKHTAkU5QpaE4i8MRN
y0ftjujWZFXhdxyyur1WfnWEv8flgqeP9D+aoBxkAKToiAGbbifm0JM9O53S2Yrw
9YNf2aqdckkjN543HdZggCoY5Czhfspv17miEvWFsmHiNshsVWIrdA1VPs4CsoLX
u6dQDsoh5wwvTV/KJ/+cEt/OChF32haUP4ivmStzuVeTpHJ8ODj69WLgrRZMOIGY
Qqf0Pa+84PJGAmHbyy8aaUltkPS5ttthgGa2UMWpagZ9YgjEjvdrqLiN2e8xYqwH
R1KxwmFuuZVKV3hRs49U58l2FOQ/RgnDliaojPwK6wbBpKiSfV7Uvr7rV1Mj4krL
r17dLfiMxWqTSjh/ty2GufLFH9AeC7kv2bAkkYt2VAAFijpyPVvoznCzHiEY9YRI
AzOlOdUxF/pOu7AjjX4WFQPvKnOMio8YIkXnIWJxID64Umks87o2PEzh2Z1Pqzaj
jUcuwqlFywV+rr/049cghdHa+l5irSl/sp/u62z5kYYGyhdXO0w1pYpjAiMc+ZW/
6yqenkvWmR9TJ2BnBpQE7cRPyNOooNcMtzUI10fVTeFVuSh3MhdPkMLDkKwVmkPk
hsyyK7GsuGOCgsFmnqSkVKWJDUtO8EsvyMVTm78GJbQPv5x8qdKIRWqhyDU4uRIz
Qjfaix66OXwzL+tdqfHZjjL8yGRf1qgBbcxXu92NZT8HkcvsGHAeifytwM2WVfbx
eS4ZRv1ZHk8PoNMe1VU0P6tQgLW2O10VU4dXCPsPQCLX7vzWuK0IPFs2YqWy/LP1
S1g86v0vV2eVHgjeIgtp/wfQ+roq/GRoVC5MqR6PUQ2OH5G4jUr+ca/ZU/puobT8
65I23HHhU7Zbqe17LfMXLB8XLP2MK7Q1AGDE8HRzkIk9ZB53vH+5LD1JWjwui0Tv
YowA65H3SzOen3HICAp3InWpiwxGFHZtZz4fsa20CS4IrHSMKZEFrt20yLZAT+/k
POBwfOSa9Vd0Tbv8OlYjGhuI2nzqGbFR2KSkEaxOg7oi1V2Gx4TIAbHQ2dwIJk+a
599R2UNew0CjLTuc7xy47qMveFo/ejRliWJj27IdLzsGMyG9FWOMiPjeSdsvEZ8X
eFmhzDCTdaJKMtrXjFGz+f9eiVRpOJGr2Kjhe/59uFDJPPK++7pP+61Z/ykdwslv
UnubIS6u/pAyFqdce1NKZ7/USZztMZ0Lv4yltA97IcRCcKu35vn0HpvqMpYnKlf+
15UxSpj0s+xTG6zcsW3JulOI8VO7c992iOIfWm7dtjlJNmmVIH4FXgohiBeLPcii
Q1q8slWBIqVlRb3zfX/CZi0nG/wMByN268KZ8y6m/B/K6PVBkOoPjS44EhIJMV/e
kveS/hYQtqCuFqRUEN/ZwTd+UCs/pi19UDDj74p4sliMND/+soicSZhitHjyJ3zX
28C7kFHkWXJQY3FMFwkIt3qTdZet5FmDG/oUGVQ4/Qpt0Wd8jBOAPcgjLO4cassZ
6X+b+mRVrbLe96vylrp5KZktTOfH+aHCl7Vl0K5KyNnqWx/0lL87aEfO7R38sJD0
vbHWT5NsyZoC32bzC4/fiI/tlKMjaNoQ8rN8wKhCDL7Mx2hNkbcJTZRHkxWmItcU
3l1+Xx5jyr9pDuh2ZKlK4SySKVuZiTZizGwqzkjYKUpSJ/HUp9ZuQYdsvWXjE87J
J7tOxC9ntfwcfG5nDGkWSJZKYTo79XyIHDBj4Id8s+83YPYGdXo5IbSlYns55Oxl
zaNImcnfHQsMMJJyh00hHzZ5G2S8sktIDkBKGNoUtPRJz+3YmCtxowz09FQ/pPQw
Cw51T01nt8yEZTD/RSky8WCLqAkpusvol8REHJzfSVWSH66Bxywfswm9alg23XF1
6DcT9WQpg2A9GHSrJNAEQq4WDZq1CrJ/pNgFx+J0P/r06uwJkXEnEtXYiPQde09v
NySsG8dg3HGda+xGUL6hI0rQ/P8Zf/iKfYNK5BzzfHZAPxnbZwHJs0xT28X/2c2k
kUScNr+UIAmz9tc3Alycle62tEN73OkwyM9/ESz1nMLPeBGCfsj3GBohnfE28LjM
nAC60RLSjq4U41u6gOFyDE1ZP4hUce+caJBsCjKteJbhIBGUCawzkLJ2L2fi/xDB
+N4P+QO2uVIdp7l0GHU8dJnveE/oHGP9KmmLivtGowrzLTs9jigOTlt9EddPgAFH
FgdvFiU0qVm2VkivlGLB9TKJr0aeUEWLwQNeFRT0HnhbwWXBlHU51rPV7tTriVs1
/KamVQc2cnRqxj6Km5b4Zm4v8m7R0TlxKE4gtBkE2/0gmi66JypQZs/RoL2ygwzW
145IVJgxfnVPSdqbovU0g38nIpJ9QBzga4MV22tIhKo/XpQc6V9A71VAyPMcBl0M
iVn1Tyb8omATtv6iejwwXJMeYHs0e9jJ1aFD2pa3pu4SUsBaqcy5cImsPjad0f8I
yLLszwDyZXasDOd9XnTJJ5WFSXe+pQkabbGH9eM/nZ22OHhFKcDecAGmjTG4ncfY
g/LQoMoayHZrsGfZK/TJ1nMdzuxxbVFml1n56ca0SITznoT3dVYPwWlfQBfhejLo
AmDYXrecCG66iedSkTESeyYeG82cKM7OB3a9GZ9g2KJZ42eDE+rjnRjUcf9NQG09
r5iSSQljEmHeGIl3vXc3l7C01HrMZe+r7NKKTkJa51u9i0gaGiKw9Mi+U/g3UCvI
Yduz271oCuo7ztdPy/NZGNM9v3YRd1zsNI6WgpeWJixbeBT0H8JWPQ/UXsDPBjKZ
NuYWZ1h6RyIxzdqy0CmajZBG9F+FNJIax0fgR4S1rjlJqeT5k9vXQBVfhnMSLNvh
X7dHECgc0LLjJ0cewnyIn17QvRXNRl0+yqppPZfEt+Ln8a9kmWZyv8iHWcmfSXP9
9RVVQ0gfAuJgjplPQEplukgxX0croxRJp0RJ5fQR8TyfrMX+K5QRI0uE4bFWXgR1
L5zYut5PTr5XkdGq5Q/ECz0085X8dOcd8lexngUxsNCPdSPfeS3Ax2nc1MPYmei6
AUM8Es8/Evi9eo/lt6toTVTNay82F1FivKfP5M+tvHNrzZqlGw2kiNeyBQX5pWI0
OZLRtafFctyxnRQV4OrzffPTg2K5HNxBA7OAzLqSiwbjxsfU5fEdsKvRrbRJVT9w
Qe3nqr4YLIsJka0Jw+f+FJ9cPDXEYmWMLJto0NPe7tOx0iTKt9lj6wM+zWd1o77S
l4pkdYZORS6AIFV7oyYdBBiVQISSBV893Yq+OcDWx5b0HZ0xfBm0HY5vhG5vV9le
wNoa2XNYR6+u5apD6it731sDg0rzqo7lUEPzglIYaQXfSc9X9hbFu5Az+X2xSgvM
D5mooOAZaJZI3cf09G/Ha+YpjzkvkUca/CtiwuMqgqwIm+gk5HtBFz7arefUbHRD
v9f8YneqChBaQyB+KiBxEA9zr1ns+9Gd043CdhDMlpOLGcap+J8/AWc827rCFIPn
9EqKfEZXnZv+lgmR3NisRj4P4cpTfNhJ0wEE/LwJHSjV3DuEHkYBunBDaXFMfrxQ
hAhZDQTs14F7ZqEpy/x5sX453VyRTM33pbO3C0jBzIA/M39h7VTd5cVYeHNUw8Hz
Aoa6A1qy8qpofYdFUJhs9YSDHWi29OwaJDboYYK1KDfLhdyHSUnxjjcl8SxeqMjn
zVH2HBfBNNB+usMIuMSXmIA6BopCEAzhOWzD7Is7FgBUTSsl7zqfPWgrmyR2GK1s
wENiuKOjvpdD1mGtxTfByztdBY6Fi/2WDBSLKAzCbzc9M1/t+S7B925mbVVtHZPl
KJm2iAk7zhBiZH9ZXnh60fMUeguSfhZXmVEXgfAKK6wN9BhKId4wA8tMwKUYtxAe
gdP9G7oVWO3ZRQM4V2Na8kmdzCTihOH8tT8l/r+6YYiOmQeobXmE1C7jfXxCR6wP
VyPxk/5guE219QO8j7MWvhp+Kn5aWPOAlqYNEU2grK8QgH3V+dsRk4Tb7B//MDmn
trn/S+jbp2s2e0pRyBWXwZKjOKRdywH+6t4tJWbS1FMlCVVpd+7KR3WRLIk5pH8K
p5FK7L8zSzgxwzpNJzupfPM2BDjy6RdcDCFDjcvGMckj13E1iYxDQxsmf2T4bhIe
mL/3aijKhNMCSquZxfwqQN9WGnJbYO0bBcvJcel/yz7FN9LYpg7gcoJv5c+VEQFQ
84TSutfthJSofH/r+w/Qqgeo4oXmkOpFRdruVbWvUObEbG7U5I6J4ejNDARXdNun
xJO++UU5HHVBgA74QxJp+Puzub/dZCJ8Yc5VQW2nwppJKN0epheimD27MXgHXnj+
aQC4U/Miu1C7KeIznPErUWcpxgYBxRS0f/Vvwzj6UQ4D+yN6PwLvp4Y4I9PxtmyH
5R2YYhkJfnsRU22fcPdwRByegx9sE0j7G3LO5ezIheqeeHAZ5v/Vg6JyGy/8v4sg
QqQcjey+pP6qAgap8GBN5GJOT3eF2wHkInytuQgCNSdH7MLZvI1rjWZ8oDr5MS+E
ZdjrDr0vybbd88s1jgub9a+nuXfRMg8ZtgvpwAdfwfQqQ0JxTd4tPu6xqBKlZOqJ
oN0s0FiQNC/aigBOKnfSMM+0/ssmPdJBnbssfoh7mdoRcCHeu97anpEQr5doklKZ
4QPU8mTulx3pkmQsvYwYZMLXpCNHRFTfuplKu7fG4oahIer5t+fI9iZ3djzf28s7
82k9klKMqDVrW2Siv7AncPHGcAsWXHbxJk9hInogLbDsB/jWk1GdLPGtQDJa+bYW
dB/XVUVAaHyOqMx+hi/UJOZzrSDqoIzl924qkwENnS6taaWWLzM/cFFyMXMvN8NN
wIIrKHyN3Zhpa3XJdNFS+0k2n+4+o31SKbHQ2Cb+prXKjFHj7FhCxxHlm1xFR+E5
79flD93mLKL6U7bw6C7iAgaWogTopRXbYmKFzFLXNMolp+kaAvupPVXfcB7lRe6M
WwfsPAoe1v+WJbYrpwHTD/Y1VoNPfXdT2DWfD5JeXcma0ymKQXp6ODU2Yb3rQ+kt
OvdkZH4BEMCcURBE+eBIXa4bSnFCiqLS0nJxMeiWibqQVgKtYkksoNZY0QjbWKtV
uRpG7TY2tgjnEWZHVkvks59yfgeqbZWjNwBM6NTRgXc9WvW5b1zq8yt4MwlUEdYL
ahwxnjzbnbEV3+yNXbLyQe/B4mo6l6ATuXyROlFTWiRC/ZyNO9RSpXzTfUr/HEwK
LqsGqj34hyWEUpobSDBo+k57xC+c1JACc8YYhmMmlBILZbzIFeSkddSJNu2vh4+a
2ReKbEWiLKJWxkIdSbvJlRK719MCDyLeXFyvU0ykocoM4er1+D80TpnlogFsQrJN
2FPSAV+DAxHde7b+cLzhfC2PigJ6BDPINxqXyO3M0j+69lOQpQOjR/KpB7pJxH4X
pF07gr27GzAO1RAatQzySDvev+dNuasFfx3Nc3ofh2z8ASXnnUGumu7oa/EHTGUc
qbdVqOec0fQcp3oAixOJneryj3vUNNvwvL9OH7yS1XWWJXehCg1z4IoDag0ZEipN
cNgM6b6VVR5Q82UdCHBqgAdx5lXp9yHbtCg/F7njlfZGmSFTGmeZZihcau1C/Ihf
b6J/OCvHEAzH3e1UUDx2aHs7MsozalEY0FCmA9rhDETI1DB7muK3iYKTlQZW3/kd
Zh7VHXnHQkfjhHYSiCclHTotdtD4lpUGeoIhy4P93sbknjXfydZGX+hiyiu8+4nO
VSXFUkag/h+gDp3chB/iBaDUIzNoKUy7rkkliEjpcPrHgVxSuqlPL/ko1K+H0z1z
/ySCz9qE/mGjU2BBhk2OqJxCVxBh0fRLLK4zKONSU+OPVpnwB9VjzshpUAhvDOo7
r9ifxIGaFiDxyqVCl/lk2akvWOaruaZ3gUX2GDOywruz5kM/JLgdttrWRTOq+gEB
2TAHQfPNpqYAfBELmAzzUmlzC6gpplEkhmx++DpZ8g5KCsqPnYu1Vjs3TAhXj04c
diB1/ADsCeQL6WFmh2NFv5wf1hcA0LgDiWyVVqQmTaV5Xcc7AeL+b016gGqOTval
z/a4vlJFX8NhWlM8k9H7wPg66MxeItNkXafIwIxT0xYiZ+TWbhsfWCOrXYDRb6PD
U/5yiXZ4Bt1pFAqY9fDbY3MIMd/bv7CdoL8KOGIA1Wd9doGmr9hkICHEBkddAXkA
ePbxa9Ri29HnRPyImMCZ4G/gZrEx+32tGXjpaInhUA/Vz/Gu0hsZqbE5MoiTckEn
K+5ZQTFm5PLFtM49vKCqVJYIIpy94fF40cN7G4FtzYmWmhNylvR12h6HrR/AwQ5n
PaM4pmXckSbBec9q5hBjdsveq0yhiYy2VL4Tx0yd1jQP60038BlnJbS6LKtx2Tqi
k2lDl19bylnFqzUXw4axeoWHiN3YdQfcuA9dkDDYFKs/Vise6+h7371nFOMsq0UE
RRuFRMbJNrRBlM64h7jfuEaWIE+CHVJL+DC1vx0+2SgJHWYion5USdRxmvVlbThh
8Zyv0Q0Pg/8eH30RBySJl4WCiwZr3vBzswFHk6IwaW2dU3CXR4EvQ0gScaeNgd2B
oYTkLM8CoGChqqp4AEfSFp61Zf9SxElqsHm/YN/j3RcWr7pbG3B6Ti9pjOgtdKgC
DqZ/rBFCIgjZotWJeJwYnuJ6DResHkAQIPSPcTVnL1M2xys7+u9j73t+aK7VuF+W
imZlYsbvKrIdzXttv8fc+3ieH8NaXFOzeq0bASt1Hfze8r6JJXktEQRdFgOacIo0
eGdFAR2iVc93EFFrT/UczsZZ1Z/z53P+0sFYVAN/y7OEPFLq/xHlbzs0ZDE/vm/e
ykTNoB1nAGZVY0CZvQ+3B/GfamJAUIEd083J05eRVHPgNp2A5mZxCuO645oXvopt
MitPRL8+7fAr0lSGdWW66nHk3ubtaUUjVAdroZYKEgNmuM3/3XVA9aP2INvyVtiP
cq8F4g5+mu7uxbjjB3Krh2gwE3UzYVsGPXThf5k6f1u4loV0XG6JxDZx4OAujfBd
VwI7aQBmDMvyeQREnUF7UOzr9oDxMfDzx4CckqenGRPv23vr4M7gh6lhWT2m82nQ
4ZHsOez9EqAb6vFppLLYN+oW2mY4oBjIIHIhiTP3T3PMTo+KROEhR/HjodH51Pyv
+DnjH6IAlNn6FxwHoqm66wMvV+RUVvCn76bWWvJslDfiT4WOkXfGL0yr/MLRQ41t
cOfLfwdNtFR7Sou09G+JOpxQFAYt3M836oAUWYHRpewwI55rT+m3Ru+gV9DddkEc
a2bdr2SuedH/XV3y6KZZ8X2+LMEPYr8/kfh/uSe7/dE7Nu57HQyzHKQMQj3xoKUB
ARKpwq80LzMBVKIIkUsO6whsFqVbSvEvjKJOYwg4Dp+ByQItHLSRMYig3Pv1Dici
CcWUk2GJpcivZfvpxc/T8mSiubrFtr3kqiVUF2vG4RferQeaJNnuUOEbgCwrpQPZ
ltKRVe2Ap3dhy5TM0w5l3NTPLtdLED/Nb9Ox733OMJJMbUmbKxLfAKU/ddC4JRpe
XaUGD1tz220C+v2OXJk1jccI1YStvv2wOfBuQr5AG+B6hWTiHPXl2HL3HTBMR4bg
lDDwhx4Rx74KaB7OCShDqhNhncWCGs6GtGKNUZtjr9b0xUNGp+1oDwcg7J8vV62K
29tKPQBJ94OleU7fxom0pCa7d+poKc7wNPADZMK79WLwloMRoV1d5ju3vdp725Tl
VWGrfBvRBEj4GU+u9MdHKHHatLHlsTh8V+lnoDK8fBSMummyCMglcdgo8aUCZBzs
dCaP+w2SJfGSbm2U14+LL3CMP0HNi5DWj86G/j6S+6I/46H3xTXzpQYA6dyXHErQ
Unqs4dJparxSGpVqWECo/i2iaBN8nj0zYFTWP0hGWhE7W5zYhfnXz6527XwS8/1y
kTVLU5M+ksyjI2nnTrhsOztV3mzcnaWxI7WbnlmcnNTkEDqWyREfRO3gvcSBp/Yb
xVrVT/bCft2gNVzzUpPMqgV4wyEUgJ7xdBDHQHmBgmlCyVXiLigGTY/KUelVDQ7i
chJeGDNglEASikEe3HjdgfCWfX5qpdcDRVUknM6uo6qZUu3xs3fkm04iky3H1UoG
cIbAxDvHSVwOt09im0iU3S00ItGXmeuOJ1YyvPtLtEpqk7HAnQaeafKrZqp4NwxA
k9/1qoNe4Kfv1LNngDRrlYM0JnS1+cQo2nUCehgphnjrRc9D1f0ZEoIArgoyND9N
nKbQFePAMBL1p+dx8vT5S4forwNcy/ELPH/Y0I0NiCIxH1nsKPNgvJsKacZQzNZH
tGRBg2NYv8Gu1duC1NOmms/s9YeGAyurEMoQAaqbde4Jd1sKdTWoDLAbHFNGdzxq
3z1JYWnUdo7kH4zm6rjb+1gfQ5sFZ437AxBmNrGfjaQMkFN4Bdtl2+zqYA09ySpr
0ut6e5WCsQtpYywTxTs7R+KWqBbc+/KqtmDq8nPGGsQwZ138zS2no1Q7/571IG6X
BR3XmqGZEZvKtrxXSAviEGCrLa8rocQb8Knp5rGK7zAHSQYAJGkpOOOLzKPJd+34
qaSA/dlYrH5WozNlMEy0050qvG6irEiyTJhf/72AJQ8RiBilnT8qmolmbShM32dq
zqN1mKXtu+IKcHmK/OkDJfGvXApXtAbCWnUl8qQe/Zmi+b8MPMPfT3nOLnfQmPiP
/lJDfn0LtTA2ReT/slWSkSlzHLJL4LuZoHYKSpisD6+XJ4j93youtMTJGafDLTDH
dbo9mLRV/A5BaRVjXTmRZ/Z+ZvaPTycymMa3wcHClINxoOhyMGo+4ska8GTRil7t
JEmKqu8u2MAJTdrsw67dKUcIM9b28pvLE69NyCR3nys2YW1f+rPeqaYvB9LflwZL
1naqt4mLVCwBHT5pygMCj4aIvGPpfH8rhhlhyX3l+m16debvLnuUYimbPM7MIvvz
DQzlIzQSz4Y6XY+R9pr6l/I5iaVOkwuxi0ZzWT7QVEhnyGwTFNWn1ogGT6GOxkRr
v4Jc7CnJxk4+w/qlc6s4K4wYAl9D3RhZDNzTJ8c/2nW8YgFVcZ/rOFsbBCi8JhnT
9FKvzhOiR3vD89kxBmJ6XmMBnoj9Ye3sGapnK5YATPb4unA2Ki+03AIo+nH+z+mz
dn4YzGWH7yfWBnjumtKYqv0d8asMDCwXN2CODq5fEO5CVi1mDkGtqwXuCXni+OrM
2IBlPeucBZBdtzFhg9hBEC79jwItCBjKwR3Znwq+53MVUpdPTdeVgSpc78jd+986
gPgeNEIAjgf5W2Tb40bkw5VTxP0MPOvR+9KqxSMAz0Dlg5V2DFmEyJOmtkCWea6P
yjCoKEGai1as1sWKfpSvFddcelPQos1GAguugkkM3opYdk36gSQS1l+AMyVNQIOq
BM2fKs7sKX8S1306p020e1c3KIEjUi8U3ih/9gpaKF1lqoo91BZgdd03H3F2/M5v
nCJsDyN3QD5t686CYFH3B4mebs+sZO1j8nAVxLkY92USWwlmvgQb23gliImg1kiR
fqzB+XC+/dJPa87l2jUtBJ1CRWErMlr6m/W3Mw5PpQkZyELX294pZq24W8AdAHGU
fYaR9o3kG4EYmb4Vw9fMrR9HZL1CumgbBdj/A1Rk4CFhRVj7wUWyFfEmPk2yUyFd
AKdqeOy4t6cFUc3D1TYryIQlCey8tWzDAC4mfUwpsnlUdaAaYl44tT3vYtDBaQu4
Ttb7LIx9sUGc7rmoJxeeWni2IjfynxmEyrFmP5/3iiKTn+jRwvFj3Zgq/AMikUYP
RXyAyfWMvo3lHpCa0GGI2975QzBtnQWMAoK821h850HKD7u/FLGcPads8cqRauYQ
q280ewMBAz4Fm5KWXCPJh78D8PcRpoepVIh+KYvBCQXzVF39i14yWk3uM5J4kTwo
cTDmgjGWZGrFIrnib8u36ZDHGMJssEOG1ZJy7zrC1Bg6CxXDmB1vXqljNbOJXnEN
tkDkcUWyiIb1cpnvQ2ADtV53SCo7AV0hQfzryaWw5K8KdxtisyU2Ov3VJGjTltly
hyqzsVMfSnXDIVvrL5B/28Q5PDhQzylMDU1Uyw5KnZN5A8gw7J0yGxiWgIoux0xI
kvx7g1z0LutAiBrDAloNjwqkgnGkpbYRd35BKBhL4AkRcTzLMRs9cSXQ44HzJK8+
7lLklUYF7xM/m5NjFJo1+XvWE2+w87lvhzGkKq0FX9XmGL16ld36cz4QgYbJgVP5
ryu8k5jM21CgR1pv9+mLQs2E1bYmJH32LVO6GnuGFT9uVuulPEnUJEJPuCE5I0E8
pmiUvXBbDJ8FplZuWvYnrVz7Sz0Mij1MP8gVzjjvsvvpfZgYruo7iNXX7wHkRFwU
4vywLNifmDxCJYfV5pDA/kiwjPSRhdzrrpYX5+0aNJKf/NvgB4J70OPWxWxTYgiq
zP/3y+mgeVm48h04DmRdauS71dxORtwmZQ/gwCiwogsLQlQiurYGcN59enb5FEer
KQjdpSzs4pxwZsCMEcl73t0tLm2AFLn3RirHQtrLiyZ8sFWThbi7PQT+rFTpwZ5R
UM4+AvW5UwZmpZ0nj2wczY3+3YpkIkhT4KvJ81VTeGyK/Nvp4BxKBBj0mac2CuNg
lmVbKgZ1V9xL7ahgwF0NEs/2sihF2IfT1KkAbq4bSG8yRn7YdVamnjuNDgVt2jc7
GBRS4it4c00icddCfT94cCfASBRb6ZZUqYtvZysAzCgiMOG3ewt2NAPz9k8+UHVi
geyxWqX/NHsHtWjntiIG/A+NGUTEaDo1J9Lno3jbgtt0qNwNH7dCHUtiEUoFNldI
yvoAzZS2uboj4/eK91DOfrQGVR7ZiQxnWVF6b6+lSBfa8BtPkdjQ6+szmjDBaUbC
SfP+TC+hLpmtmmtwskN/FxkOO7hZUK8QUYi+BUkLG439drEBY0tqb4hoPYkSBh3Y
lT081ZbxtjaM9e8+f+WLiz6YZ+eO1ER/gzqxIjbQNQTKTOdBln/jYFUtX2WblBMd
NGStTA4Ol7rQCALSQBO44ypkhYPYU/KMZFhobNZpCE+o3OIGANfMwooyV0hle7fE
Ueaj75oNGeaxoSmPxwIhyV+may7cSzNgFfCw+wiNcHXQ1Q2gVLLjWM3h/6obqETE
1KisZYFBy4jYEmKT41LOzuAIMHRMyvmJ8my2/pZRarfcEnH4rgMxe8YjCTsRR8cr
6M01PonDuJC7VcFkZhFIX+399DIK+nC4ocZLkPNbce0XwRY2POR4tn2NgbkT3S9L
D//XVwh59eu3CMo8KHsx2cqazVFlmWUxWULA4ddXHIJvdZGnRPnznE7wTT5G+DvT
mArsXBryCUok2LDUJXbPwR0Jhs8w3MjLxF0OYiIj3SeqnpPWectYfoMKvj6UXHQj
Y+NwI2B9Dtn3W+NgLGmHa8VsrlICHX8brhLJKG6TpV0gMHPLLUPsNU367kZqyfD9
5reI5pFzRkTcWIwew2UeO+/XJYtrfjxtzVfeykl6CRRwf3ifvuBVlOFFnLsD4tUt
c4hobzowX9MbIdBAKSWJBbASuQPvCF+JDaUIsof1MMM+/9fCJKT82mt8Yy6VAbCW
uhxDJzdQnvpVy3Dgwb68B94bxvDEoUuAkpEgOPq87Q8Bgx+yXZT0vnMwpR5gKQ0e
gov0uMZ1kqzYd2kfXSc7rFl5jNJ2FItZZYV1/b0eliMrOR8vFuOuFcBTLbRu7yyP
fD1mKTwunix/XEKGMR7HDCFmhWgJ9G1FHn8AwxSNRvnpRu80Z2+tjo6LywAbivSf
GZkcjjgtc4PoXyo3A5LCNEEt0rWO+DD4haAhYDU8S/BCLNub5PJplMoBxB+uLUnT
AbM0Ax9cY+n/tsRVdBpYsSzuKc/mg5UtJSBwymx4ol84FSi7bmW9GcDdDj+q9Zav
4yz4Jz/2Eethsy2S8EA6yucMDYxGpPp+JZmz8DL06+3PeIcWywxu+JfaVXbT8aS0
1y7v3yMzIO+ROSBIjUNwbV9kzt1bIRVBJB1kfQeCmpOthllthKydAIDtX9b+4hgQ
15+SmR8Uz+JJa/fHTVbMireUi5K3/BJ7UgFnT5YB6Lw49fhPJaLWwC9W7OYjsopg
E2D68aivtD4cfHOHSYMnQ0Cn154oOdgTw27f1iQ/GArZ68XJtcp72rGKee/KbOiX
TtmIWhjPNbn8fhs4zd/NEP7hm4CSVWnEw2hOrjpxMyJ41eaAvop713Fv757PrDPT
M2doAqLGw266BtFOSUBsrAOA5hp45ErcRN671FHKrkWHMr0zu/MCxAJ7L9mmhpia
NHqGb3S+A7n+YNhY1k2uXM+Nln/7yy+xBwQlI8dmKRjob1+1uyugUMTSn0VvwP/l
FBtOC1vLHIr+AbW0U04zGgNUAg5u6PuzcBbRGvLSkrh20oiECOrm3yCa6MONvS5c
jNyoml/5sf7cftbXMvz2EoBTPLqUrzT/AAuAz2F1G3isEnZzNeNtCBNnEaPOxFab
Z03yb+ZXXx7AO6AsaFUaK+fL7EjmiSevW7w6OfvRJ+x2NuO+N9X/twKOyVCOtweg
NAooPBxPpnvdYFveAsTfxC58aRGmvIjUw8SylFAnKeMplRGnHFxJr2JVJDGaQ9CP
HwHQWmiK6I2H7XS4QmWeQRWA/bANHLDts5AX1GBd5I7SBSUklgN+PdDbPGYBzoMf
12XNAYSv1rkdE4xa2VTegm91kDC1HiFZrqkDdreh9TE+cetGkr9zBgbOpOy4iI2H
eLyVE0i0cmhk5SKf6kCiPIZHry4n16KG75UUjorPhWcDhr3z1bBlSUP0sjbtCYO4
VZQ0t21bZogpZtJgUV3HnpgGiwZntZ0DSz5R3hAnri11m3klb2bbmAt5OCfF2brs
nCSfbF8jp9nV9zjvos0eAJ66ntHLoP7MWkEb/JqAxCOeQ0K2SLI39ch9ZiT+bSiB
ilkY/7EjApR0sjplKyiE1HN4Xo7qoTax8fPnuVX/bCr/+W5QohXmeeKRdhVPa+Rt
WZohWDmxMlDoAXFraX1KWMax/Izqv3y4bAtoiMoI9wCM0LPZ1TVtFUjHl4ePaXdt
JuAB9+Vl1HBrIvOgG7AcVovaFNJU9hjDr/W2NDmSMo1A+gqY2/THbMuYd+OsttS1
AUxVqEfyKMeTLxS0V4AsteVySCQMZ09Z4CfxdDjZR+BRzoAwFzXSqfnLDkNjC6rw
DcQmG/nNkt1cs+GeZKplC/Xd0DWxyXKPzpVh7xuTds3RDKxENnJC3iIbePVHLA83
Obx5a7ZXQNPm7EsC6VRg/7nGDPeTNUn9L0FVLwWxvFGbWgV9F8FvX1hRD+DOJCcJ
sOw964z6V5oGCW6PSBNViI2opBYsZqkDP4f1ssFnHtMjvt65vCP339G/iQe6YBqa
hxPXRodXB+tFd+DHRZG8kkGV9ZKswamXJR6XusI5OE2aZRxouUc/dZkqFP5mP+IE
VgPJoEoTNSWo5oTp+UxvUeqA0O8+U2IKVJRsbOkVhHGnPnetvX8C2jym1CG14G4G
9o3EwGbzQ/wKmYlaTx3oAewNmKGuSQMMyv9Y+xJQboQzfMfFly7HF+Zo7s7BehyY
T2ai1GZj0xxHTol1oojULtDByWECjPeWwLA1qUJRj/bU5urVHbe7BAYh2WyOdH82
KDwsYGyefWbRaOMqn4oaE4wPwL+DShOB2EIJ3HRPykzriC8IueXh5iD3hyBxWyGa
jCUZtoDQ9tvy8hpRXHSbJqPP+rE+j7sQK0ePF5Lms5gvqR2t3pJ+yWQS7AVrSyKA
CSNqUa1eHG/BhvP3F2B75e4LXwkBFwMqGyankl/Y7sTgU2/uLGTa7EER+AiIaOsC
x3IPfAjYNO8FByMiUi48jl+rFH3Oq261YZnO9j9L0UpG0TBXvCm5AqZaNSpygIWv
OGMeBzPmEPWuU0WGq4YQrcPNvTth+utERQbEXhy/HCgjkQyq3dV4HSj+6wqcVNZg
ivGHjmwJ/yjbzWjUsK32Mtn3l3obZ9G2AQ3C/+jMGEBYNFDNTbDvhSVNBK9zTsaQ
PgTAoixvKyMzJ4iTk1o592f3ErOwADytZCzKKv6kLTQTeA+JZ+MQdxZBIiJjHcGZ
Q+LyNuz+Zg2ThSqGBpPW+U6x/nG7iEBuY2cB3TcrDQzgEzIckgciJc5HkUX8m6Dy
dqq3mlW6OnuXHBo11CfV1UQeREBW0ZxWgvkq03oV4GPmnhqxHm7Ha8muiAEWzdqR
nQbegXvDGkpOOj3I/7P4OAbF8FhXz4M1BeSgH6zKw4r61zDfVi/3mKHaMbjjhQv/
0anIGMBKxntpOq15n0oaqpurYOd6pTBj92KUb0vSLwtn11qi0iAV+25agKJHIq60
slr54jqCdEZnc1QNdMrJ3sDn6maSNKaVPN+1agEWInP0OMJSjYwiw3zd16KE0tlQ
rjiVv1nRJZHZHgs2yZWxfobzOgZOFqmtluKUS4lx9fBS1YnFMn/rSSxwPxABKNOn
UEtsKO+f4UFy8XMgtUP/vn/m4gat0ThRWop5hyjoN0FBCKcDCFu1BHXtx0HPbeMB
RWlvR2Rd9E3BpG76lt4ROgcliqkK09Yd83yrrbcv/bXpE9cbiyftf3jeuc9mWwpZ
XwFdc5FTtpimUKtXJy3JS31dOa3VL2YZa/qFoQyemWFSF6hXxio8/IhEKvYU7AN0
2wP5Q6w8h8qKUz10nz0+0gfvTOy30qL+f3O6VzWP140kqXLFTD7AA+XNwYbhNZ3q
iXyYviqlJJoF0mOwuT7NzzedwEfo7y8KFOpwPZ3tPVfygrwNOLLAs39VDYTPF+XN
6ARNRmlRtDCk+mRA8goaxjb0KqG/QbbfnaX1rA6mQgGUk5YLqiUaEeCkeM+E7/kV
Baj0U7PyQMOVeEZRDCT79O4CPb6aaS1FCRuas4aH6ztN95SQFEd8iED5NidHjd59
DlbrgV60GUB+IyrPHhl6Q2vclSU9cTt7LA/GduKO3Orfvlt3Anx547eQ2p/JjIHA
JEIk563uXwP0ZzIE+1yCoc1BwPULwiX4vL0YoAnQQIlM/QmkO67LmN6s8+DVA8N7
1crBNRBMqVkWP8TYseMIfrWiqbm+34diyU77UolicuDV/AZt18G9onC/GP+6A8EZ
GG4Cu6oFD0gkehaYslG3/IXkrdd5eCzSscPHhm7He8KnvJxG905NmF3CrAARWA+/
41L3B+Aw58yPdk8qa+AV6JDrjgSP0yhlmPUUpoqD4Enervr2P2eCflkB9h6SMiZ3
j0U0llM6x38oP4WesmkOG6MFjP0Opj4p+8f1m5Tc2CxWs2tz3vdLJBhVWs/rRIQa
DiRq81DJIFVwWFNflzx8FkPbMHIb1QHkJTUyMarppgM9QZaguHxSrdPfF/5o6b3T
3T3yjYbtn26n4cN68kiL2FFJ4sqxOYyEoqZTu6dHXdig8nJvkMBuesTse2oNaEoT
ZFHAcOvStoSiOEZGMyckgjGEK5TBWJqkYbTdCEpmYJuZTZqyDwUQ501Zem5vtLZy
p28vdh1JaUgx21rau42c0zG6Ec5sdHhwlowPDi9aJCjjw6e/qO/hwH5OslRX8eCY
8Kl8IleYjiHmp2ZF08xf4MH/GNr1h6U2CBcfahniUlz/b9kKQKl1heMPYR4zZuO+
2OBmcV0sOoYdWX97O/y20wykK3i85/9C/9/T907bZsmzT/mSwybL+DBJJ07DBIt7
bqaBOsnj8YA/wI5wuM3+7ya4onL+8NOF56SWaVVZMmoix/3u9Qp/PO+1TFE5BhYX
SIH/q40744ml11fIN42ViJGccxCahiIyJ+5aMetAAFiCGhY87q3LadnXf/KpWu88
yBceM3wvhoKiUyfiV2RA+uyYs+DZ0Dn/pAlNl2lxc9bVson7MO9nL+AzbUqjnS3m
XHQBvhoDyh5OYtXoZp1dhhNnXdwoKl+n0ak/vBF/Pl72SMu9R5A6gTQWZaGTKnIE
C07cNGphqjMmCONoU3RRmtMillX18V+Qn6WLfPGvbdZO57KcZlxYM/0J7a5ky4FK
GHXnQA63EYZonPe4rOyHfL67hIhTecpqJVdu4xaSeiSiQy7a1dgyWLh3yXnM1sWx
477puXevwLzj3P+R+VVolVSLlZoyY7EARAoFD7UpKjbD+0jcjT52wenn7nQlP/f6
N8F9irmmUbmaIYpiyu53hAXjXxiAuECi8kP2MEnKXO3TY+UN52XK5irCDUUzk+P3
FoMuc7M/zxhki4qJxgj+Qd7oQ3kTJ20E8yYTLoWsu6v+wN/kKYOKTv5T2yke9T4w
VGXxVDwqiOBcSeYi9J60IZkOQS3yjL6V0pAHjIZxZpkX7nDtNQGHR9YzqHzLr3Ak
qZ0WAzNFdrllr7d1xkaiWCTHSwOlRAU2Y1kDn7itDpsbwQSn7nKA127kkAxe+PPG
HGvXCJKACjFsP7DHQNGakZW4I/7SOY7vHS4/5Yb6XbqPeHd7IzMc7cL0FSo08wf9
lvm58wbxqGGempTSVUm++R1v7SD5nytzzFdPyz+yOx9uoUehZKDBh5WN74A60Q2A
U5NuAi0bna1TAVn3uzWsuAiWc1CeymFKZDcwWgROhqozcH/Q4kdSGg/EVsTozGo4
7VYTiqHdYW5jl1wu96GnymBnL99PW2j0BsvwZFlQeoEzwFnn/dGNwb24TlMIMMUA
FIEh3oqlKdFFp648H8sXD0gj24kGTGZ/HlF/5DH8sK/vroX3UteI+1Rh4NoA4gTZ
PLTw/IVtLx2SuZ9K5+3X3uy3VO7oDicP0WcRYBoLnbDGBJbUQQRZ8gONiMy80DQd
AUQueZ06nEW1eU4bWYIfPfuWFM91NOU0kkoasoUJIsNsPxkopGxapZIAJYd9iC8K
KEVXE9Fz8Vu9jwMMwH09U/FEUfoPFSOZea4jx7e/cZk7QoZHBgaHcb5lFrrajS0L
OrEGpvVITLQN2vPGeQfFZWoXcIxDa3k9gioztfOOQdcKwMrX2d5EjV1HOGmyc7U8
cHKMx6AXbPsRbciIKKJ3+5tg76PKI7I2lktakOgxLcfQAF6hWIL1Q2mnxMudU6SZ
voFie5AqIoIgGkaGGO4H06bvTHDvkKVLJMc5cg/DOXU5Gce+BV1UON4RuglRqRQB
ewg4QY5lPV8+a9a0pXZwwtNhLLqUCyGQGydRUmyx+6V7gtj14l94PTnUZnbzeOB0
6E0Ug7AglvY9A/xSiZc715GzVwQIK+ermXpZaJczEuNPLbsMp3KUKLliVdzSgbvL
1969Aka4ehiV1g5PpVkpmLc23Fv13Iov9GN/pewWS3e57TOyCGJ501iuw/jt3hOq
Ap/6uf3jeG1dBRzGi/bQHj4QECKXLP3Q+TrNK9LU/jXR+ZECdWcShLnvwTRmmImc
SqFOyo5Es2qRAEeG7NuCTgaTLJAfjZD9TiJiGGMDHRMRI3MnGnSNT+PRZiKSZQoC
FLBL77SKXdRuQV3aJP4tHsLYQaL/uhoU1sz5tqmdirn8cvIHeM/IQNa4etPB13n8
FoVFxwM/YJaCB/we0v7iPtYYITTXBPLqxz4lzrnbcf9a142q1aU6z6e/YSyC5uy8
smtb/CJ8xFX4wSPqJ7X8A1hbQOC5AuQ7YD+zAF0k4ITaCqRqDtIcwJFrtBPfE3Mu
lblOs84dy8YP2k9XJNSfKI3/vKQNVvHNyUjoDQXdeLn7udt4aSVpy0UB/6lMRBBJ
iJyWInZRNS1djs5H1NxAvm5RAVnyUDSd9UPTtWnCmhv+/1xbriRxavu/1HAcE6xP
L2hqIwbH5Z0TJJKCHf6a2VjY514yS2izcvU/pzSowf4wUxOSneMblYf9aPpNezkS
PZOfIIa1tPdHowgwxWZbXsIh8/rdxuNkqz9xZb2nIhfAp3flKAcSdCCodRCKzihI
YwGDCk0fyVGNedy6mMDdNBZUncSnBuzmKhvZY0iSZKu0S35QPogZOsd2Y4pQNwMy
Nhp1gR+V7XgCaYAr7Pz3V+5DsKF7eUiPN/q4MDlA1Q3YSkM0eGKfHragBUxKBEle
sUxFVgADbjHZOhHBJRtDOQ8XEGEkr1iBRtYlKYvTzTv+TIZ/UZn0ATtlCcI5GsRJ
lv+7ng2yrhtkp/Ba5QYfmsL+h+C/3GhG/6kqVeoYsWuDpfQh0WvIfHFeyoSmQWx6
OZ+pUqkR24Z6nOtBcixQTf6v5kZc0wX+UhWEys5cShjS++0a/iVSBpq7HHlu76ul
20LTakYRmAEEVYYYRVlA4CNpe6qRL+wWOMNZbR0iZWnJzTuvGYpMgXuWp5qi+aEI
xb/9g4KeEzBnbm0cLcEV2C4MncXM9nTheOI+avZEcKNnEpUiRjMR5+03gICgaPFh
vgzFcr8P+asR3332rgrCWuOe0+Cn5/54GpTMzVymz253H+RZQa9zcDDq7zIDrWI4
SiRi/Qb9mQqmCqx2fxpSIMOi1M/glWsX8yhMVB5g/vb2vJLroSxzP4BbOlQDt7NC
hMHjoKxMdZOML6HdT31uv1MQyIBqfkzLO9MxN/7gt8AgI8a1VRt4Q14n14BGaQYr
QNN9z0OZnXK2BaA6YgNhuGqK8iClug5Zo75/XmfD5b3FjX5zvnB5qryXKI2ikPLG
4pytct+3hkQ3LV7keUoRzIhaGm3SxVtbFyafkZkbf17iBrwlme3JoEl4y2b+Nu1J
gcvnjG4KpVq6c9zBGi12Vzh033p6gQ42bXYpXhF6wIAvE0ERuJ+Tvl46r3lqLmKt
QqAcdmwy51TPSvg0udIxXuijuIqndzMm4aknp6O38veh/HY0kfYt+fFoClzxOux4
/CFd0JKTKC8pi8CWSsEqtkJVsxDKmBpsv+1kbR7UF0cs6guFUMpID0QTb7MKGXHK
OivXdwwsiIEldf9yh5g0fFk8XRLXi7KXClK91Q87t+V6FyN59A5AbzATY6N9r3EW
wp0QIk235NKlqwQIIuz+kC5tu32ZGkyFV5HudrxmUQCbWaDFRTWL+xR+G/1M7Pdy
SwRW4c8ceM1v7qQ2Ic21Fpo3rbbmQ2UvboULlKxfDB9RhoQ8LZPeQpvzMIevnhl8
pKN9ArCJ3fvx3cpBLlq9pLxzFx1JfZQ52P2a1UNfzi683xLEiZLgPg3fJid4pO2E
127hDpPIAId6p5WejIcPN1SxinF3Hn4Du/JK4UJ71LwJrf8NEncpvhTihi1f1Bb1
jLXYkF4vRSxuKCkU6faPcAmLHVuff6+MUHXyZNzSDMwunaskAYJP42UwlxhkhZp2
EzBfF9B37LVGlszANXLrrO4GxmFodFUhzI68MKD9zOGSTL9y56IXfgOdv7k++itk
Dkp63TDSn6rjhR01lC2MHf7sQJCJw+3vUZUl7p4DXvf4Id+FdCouCSQPHrZ6ZfmX
cFAvrTM7Hp16WYmkmMr29yMJ1T7djpthNSbDjLe9muC8vg5lCegzbt6YjTAZPLEs
MYSU6Gs4JF4ULDmco+9Z2FRT+Lbh0xHZ5M77IbZG799CFWxSWJcGuk5IhAbRcyVZ
7xbHKmnTi5t5D+/biKwAUk6h4r/GaAaLZlP1qWpNua+xoXXwIZQF5UOnTFJzPmCx
eu+jc7tlnSHLDXiQP2hIXLxrJMIXBrRElI/KKygWLfKGL4+fWvf39bISwhrL3/0u
pY6bVw8aF7pbsxNusbTVyKllV77OMpuCAtLXZyotov8ua5/31nD7iHuGPsOfWye5
OkZwNreosUKIi9MloAsE7IHB0MlVpeUhb1hy+XlsVatzvOOPhIA4ji34rUjIZDJa
rCD2iA8xGzp0j1wyiGW7+pF+vjPuuDQDt0fXMw7EQToRi6XchF5Wl3eqpN/5iinA
dK8HdNc9Haz1m1CqpApf8w4XPyIGUQFXZvECaFK9GOHnG4WHST3BjfYu3mWdT/86
u9XuvT6AWGA7hfXJYQLYSnmc5sPTQERMKK0LKP+BH7k3aqgb/belY6XcT4exRlJ9
KOhrO+flZsVdE2BJO47nNOJFL5mhcv7NJGHJJk3iN9zW+yK8dHdChb/DkjhCxPwH
jTCWKGDxxfrHktnKD+ktpn4DbTzUXaT8k7z/jtsaeUBHRD04t5am09YFyGe9fOSB
pOXmWpVIUJUZIkNLHBGp9x/WUmvORkrJmigx6i2OoIdKx75nrh508gQTsm3sqMjx
f8Lpip5PoVk1klH5fAfSmK0sFlxXTRXibE6UiURTVIKy81JcvQxQ+Q2YCPMphoa/
2Yb81AkEEoSGJjJsGBX1QkpanFJkcQLeS/GwHbKAjqvfiGZtmgcXZcxh6+BxhKCk
lLeipUyZGQLi/UYkRfuhB5Vbu2ChXG1jchXB/0Nun0w2Sal5zhglljd5Ov5WemkV
pZhv5+xvCoZP+SoOzVcrwkxYTBiVwJ3S59tlExif1BXB0EeUfhDv0aO+eMabwZq4
ZvUyVjPJyH8K7hsR+Uhw6ZMN64tIMZUROc7EcBAlM8hJqOIdEPvNi6demHSgeLLM
hX55EZBg/uLdQf380j9AO1s0aNKmBclQe11SIA6U3bwNL1o7vvk0HW18AUqd2QCS
Xw3pFKAVPPyIOTg07jAgTyPGkd6J9MoL9l82TkVpfpdFXAEoaH7oNhlKoMoturRo
ZolGJg1Wfr3PYoEa3G1BkEy9Kiwmtxn3IM0Csi3KzE4L3IJ/JSBpQcI4m3CvI6Sv
zvFmA4b23TFICdlWHjWta4gVUZsy0qYIahaQBQ655yt14a9yOMc2AXT05xeNvsQ8
7s8WtdyaNweMRtaM9Rd1Izs/9FHDyFRLXcG0C4Hp6TVrAdZz6xs0TUbtrj40xmwQ
7HSWZMGR2BF6BSTudq2zb49TTuz/0mQvOq7rd6cKySMrQzlnFdVWpnI5Of2IDV6j
BDXCszRbnjsWBSA/np1j7vj46qyiYFbEZRRQp/I2NlBJnpAJKHGwlb6fQsRyjZlH
ol+2cclym6v4qwOKDxecY7KHBkMq/913ZOXy3+pIUhTRP2lWFh9QCbZ3hYFjFMh6
52WvFn0M3O/8gtp/Qp/8BOgCzi/ABcZg51WzneV2ldHV8eSH1YZoGONEuQB1qKoD
HeLTubyBWOg9y/rQKsMie2FK9slJ4POjOSHbMOxjZy09I66mGZ15C/5AlfNT4X6G
iEV/f3dqp95NtMlSFslCqUauXZc8LDBaIex7/0r84ZGKurR+RW4fQVmjENg+kyx+
wAotZVkC8Xf4Katf6yigNg2lhr/AiXKcGyl65IOE5ZKMnGUNVXaNySbdM82wWoyW
bZGL/WPuq85pzwaa42SWPc4eV1P3EIYDHzQOW5n12XeNQ7zs4xRthNfv1kquQgrW
n5zDjq0g52inGnRCZ8fqOd+p4TUbvPWQtghk+9ElTaC/husP5XvNMFzrp5R73m4I
U7z+l4c7Blkwr1HIwpVaii/rgrqCmu3qNydfb5jl1f6ovz+cC12AA+WkqtofDm78
NKZWnJ0Q//Ji5hA5dnKmy+sNuqyeFv59b45zetNm7NidWZLd0/ItjI/hzHGfLw0i
S5qhxr5QQ6ugQWWb5QcjDPUHt1F+5NmszwQM2NXFDnEvU/9DgxO/O+bO+a7bNRAv
QcxSB4eQ1K/o01xovUqCNDFQnVLifgIvBZLr+X2z1NBHp2m0L2AwEkGUo77Gy3L3
b0G1MaTi5UbzvgrEPKeGYn7ftq9+L3leuiQlNGz03Ds7UkwV5W/5GCFNvhlA3m5P
RkjlhaF46cJ9xKOv3NzuipHthzUXaQTUq7CfWUhN8NP5Q9moEr7gVg1y/6N/0XCn
WqgFtzIQBA6zIz3+pR1bRCf8/5vpEzv89eJr1FoQWtnjCjLxvOr+PBze+U/3j85U
xjZaiShvhM5tC0qIzknnKnpUbf5EL2H4G9/RsOR/tWB2Gf/v/OWSP+eB4yM0IgYz
rzGzb/2/Vi/BGXJhTQruYa+cviIS0gtkb/TV3jwXfFSK7FuzEdTWRV6Wh19MkAps
aEayGLeAwbC5ZtV+IqRyJpOLIrzkhpEOhJMEeyOAuFTE1jALrOJZ1GzdliAJ++Pm
LvGKI90ZExxZdxE4zVjU4OoC1OtC1zLnASfEGleDIHGgS3NGQ8+6FDhcHirPX8a1
HFmHyUkTZ4epmxCNGwgYR7nLi3yt91oPGge+45lTsktV5F4eCX94+e9yBAL4O1Cz
Cv8LEe4lPZAtaJ6GjmHzHv7u6mSj35x/DqBz/06PvRqmMT2gZsskL3zSpEm+HB7L
MCmf8ae8+91qXt97j3bU/Bh7dw3U4/3Yq8XBMDU3NMX9DfS+YrOyQSfgpkElbri5
055LSRpehfDsgVExeFV3eXklSyFMOmcd/ycNN+g8ChYHAVEiQKEEX9bh3aNsbyxj
5z8kHtNX9png+xlU6bKzVKXZGAjLWVeClzWM4HBVc2hyqDqCFhSaCVbHOcI3osZJ
JXOyhhKkBWg2MumMSi8vaAsF3Aubw45dhifqSoiJEb2bJ1ov9gBoFHabf30lKVCg
iR2pPijf9duEuz6RFX5tABUcvZpio2mlYLbAzmMOJn8hBsrbYrT56UfHDikktefG
RxAKEG04IQwuu3NTmtHWLBJwp+8XkR/bUh9+/EaLKS9MIB4YpR88faMEkkkYuKlq
IOpAEm6gc3Pexbe50HEpITe6+apt8PboRdI8xbn7MzXToQq14H0/RShTvX7AlSI6
EtAIkS8nyY4DiFCK3Mc3zxlIEdiEA2qFZPuA6Z6Go3bOQcjnDVUdMbuy1wKKQBhu
W0FsgFmu1anzqneVOglj6GgVKmPXvxv6TzvMVmjKNCYoSIS5qbQxrEQoq8Wa3yma
UqYjhbN7+vvga3ZFy+dFOmHdPTkbAJieGvhxQkGRak8KGFlRs2DOZ0HTv9BpLU/0
xrlL+Bx7Z6r1RZYeDzeKGjsJYbeW2OZsbvTKzdiFoHGWEag5nwO3grw6HnAEodxJ
LpJD6kXDvE8ycsQxzqCdWaYSeRtyG7fcZHWDTUrJbD4BEcxPJqbNM6aSs3FAWCKg
JQDpxjyICUargfI7oPZfjuG8+StYXugaS+Ec0Y+OADDwjAo4BxXApreAYGp3wC5h
uGcNCS7XETWY6KqkMHLdEdVyFOOhZ9+zywkylnjjrV8H5pyyR9C5IDonx1ZrIxTm
JLbLHszTfG/v2Qw9W+TfZsp99Rb9zNjv46n7rQlovbpZX/mykjetSVrcml8OOnjx
w+1ln5JbvfgZVfGHxrq9lcz7F3EuUT+TCjrp6v14ya57/BxakMeye72H7LUNX8dl
fp7W72RGOtqYxUXlHSAv7iwtouDAIZ9F+5CAndSxHUNt7p8aOeGKDgedD8xazToX
ym108s5v9dd04V4Blx1NU1axLd4SDCr67z4tZsdN6SpSTT3O7TKC+Zb9CuAWE4hN
6Kh/K4mdz7DE+fQwnPSTBH6mIKyyK3cluNEz1iliAPtIoyUe9OPrst6U9kvVYqR/
i6+TZN2xzTNknLWKKVK4mV9d15PcbCZ3cYVanowqEEOUDTxbO/XLBEo3+h1hfKYt
nE7V24aW4Lz1BWKV9DbNC3tiCSnLnnaxTv/E6FWZnk+wssrcHOHfybYT/nJPHnc+
+J+N8X0XV2Rc4Q0Wgztp1zXDYuOx0f3K/B/5OwY6ktlbNBEKJpGljX0SCsIKoOPP
lBHx0wd8ybEp2+onOUAaE4PQGFuCCwLhl6cueo7zUt0hDZPkBLizqz5BiHWW0OnP
tGi8zuexlB867mlV5GV94/mlw/SOfD+FTgWg8TfUZ9mHtRHNBQDgKGdA3F9rlJAv
5jdCG8zV7OacCIn8elh2tV/n2SM7gt2a7GeD6gNra81h9cWQH0KFlOP1h161UZcE
TsWixy+BIgBjEtuZlkXTpgdVCbDLdgXK9Tp8AeXUDJkhHX9anGJdAFtHTXhuBbty
CP0Wv/8GMTheITW2w0AlMnzV50hHaJEXsbMT+ZqlzHcZIrqAxp4qQFWLeC9r9dHU
wxejhBZUk9FOSelIKW8aTsPncCdOKlNeIXLwAHy6w9DAiuzZUo3/3U3VDpNWtVUF
RhLB/mVCqjmVv9bbqULK4CNbFGXOyYhKUo26wwAMzZUu+sBiQWut89a4jPyPUA9z
nolPUD0ywXdrKk3d+Z51XQsGhGusfJ/P/N9R5ueyNuIiqm1i9kq5eR1o+WrF0gme
8CWMZ2+r8NOzqQ6BGXkfRv74d84Q2wNsF2T1cYwTX6Xc9JhkK2iJJe/+sjG43rA4
dKVC9fDs830rFg5ZMoCOBCsx2wvoTKnXcVlauTfcOZJiDdnwjkpDnhXEfl5f+lqx
1KraJ8rAA7fq24fSE6cZ/Yh1CFPt8G5zv5Gn7rpkih7I/nPY+WB0+HAy/NEV76c1
S/BuMH7rwW/D3DkLOfZ33Ao7SKzpc/Sg96+0zd0qrYWjzNDEiaSKzJ/ND/rSbFtN
CLG6YLGzQyCdwh81sHkEaTXmrFt2t4Su/XFpT4y8Mvq5O19hBc2rh9grmVkFIxbv
/DqaYqCSOF4EU7p/oBkL/PUAA0DVeikayCAx3DifKXsHzNl0ifsTz7QSRWE1xibM
Xq0qgF1JQpTcfKiK+tkdM4P/2Ql6G7hnH/TxK1kAKUoMTxN1ta9Cfsrh0q7c8uTC
LdLRVUTk+TbkNoJMWd2sTEicX9FOuRbmm+6cw0m1e2DerO/BewhMcFMygjVTIYyt
S0iLtuAktt1VhPgT0sAsC1BDUebiLs52kUmsst+kufGO7+fz5vE7T39kyLNd0XWr
bLQ2aGb0lYrD4aAePhSiPetMZWdKpD7qdRYik1QAGoJNG0aSwI5lbONN5QzcBq4s
cn7xPFVE3ZJbtVUDB8pegjiJbBp7ASSqSv+sRJiuTRg4bQA1GS1O72nQqYLhxKXg
566itgw5KB8WEXDx0TCnhNeL8zWrVu8oHmtfPsFNHDSt/IT6rCNVztTdVA4Q26x9
ji4DN27nXvftD3xMRhPNXURmHhFrGQYKj53faGXsW+UkIUwPthdODEGbFiHAArEc
Rn0iI5Vs0qUPmj++Rp0tJIvaF109O9M1M5b/+l0k8eX6c6Wpg5QrESxLTGj5D0D/
REF2PMl5Fx7Wdnky95HOkNRcXI5BzzPSFYUZpx/Ers/F6gs7700jmA402KptQyy0
527RsEYK0QM/rcOPBuE6F1avtJBIIE9t7+LWuzMKCZIol6NLWgp6LsV2bHJ/OGsL
ZjQSeIdzySJlttuJvBuc0/UtQ7zQPOG/bvBNrk7VGoylch+GpMLJqQMHkINKLOO/
v/rD6aiZEV7Gl+4khb8wWhaotuHvraUIEwsSei+CW6dlq4+BAESXpXRtN+3EY8wl
6T5e0bjiOyqTLawUpYywa28t81u829hakdmGhQQMXz2TMSPwz3sTscwta1YHRz9Q
knSxPBGoIXKTY1tPAHYWQCHDzKjGv6jV76R0iCMIFJ3I42chNRBaBwWy0AP/Z/cc
dtfsN7kVUWNAPkeq+R+zcQ88/wpcn7fbkL+vscimHS1AQfqD5kR9DIvoVYYtMIMN
zITPkFiQpcAKaV3wQASGjwS55rX8oNzlTYhI/VqCoZse8BGzdPrTUHwJrR0gsVUY
l2cgXEvkQ7K3Pnb+1YPFGFc7mhzTxPmgyqxT5xsWp3fjfG8QEU8TsYfmz+8CXYVM
12UzYCtEJmAzcfwztBgzcIlntgb/SUUbyD6uqkMisqhSSLMKtWOnAAk9K30fAu7H
O1LqnShwlyvGBzDBRYMc2GgzsGU83Oc5a/QE4zWNAUsDrQHUPeS5K59v35rWgBk0
+ismaZ2dEOZWgrAmKoYIULuK6evf+gdR4seSr9kOsW+ubU0op43P3wZi9humM+Wg
gMKXalu62TiPdHuVh8j8XCv+aCpxiY+1/Z3MStz/Kqr0bPSdQKdy0yh0QIbNZB0t
fF0OBA+tXqVYY5SHLOLRYxQ+2rGa8tuAcSjNzVR01ZOY5yX/U6k9jXhbqUxEoe2X
ge8GZLMlcSDQEkqLmVAqENzHAsndO9NtRxtU2mV4QpgLLoiX2UWQfxqZm/7vlQRn
Tr+M8/l9Y7DfeAVVZdr2O7uJ7SUM28Y2Bg1lVqbpcR7SD5BEH1AiaDoURsLjS3Y8
CPZfzrXAkG8j0aAuDgI/oBxId6/mNv/ks0QUTpOpAy4gC3gfucmsZ8eF0O2bpZCY
Z1iJUKWSY1aDVPpVx+bRSSkUcsQBcXCfB6vlkoL0n5QgK0QHH1Wg2G3uYanYuwMT
hpK+mZF+cQ7Y2jqxSvyLc0R0rvZDuy+iLKcAkyv9JO/RHLJ6zsBMUTnTHHXkHr2L
g84QhSNDuc1L+a9Lsu025j+ncPAPib1yhoYCpYbIJunXBvQTlxVzJ+RzT6BJE66M
+A+ktRss/553XG9iJNpLi1G5bw3aCz5nfJrjVrM5ilNrTRrc4t3s0QO9/Id7CJYe
Ml1F85oSRu2L/CYngbl7Wc1yqr3e+jauryHUwZN5Nn5qBCh/JhFGAFejKhPbejDR
ZR+qbfKohY61Msr3rq64ToQB8jIZJxRFPTc6UNUBSYFpbGx8vDaCb5yY21bruTi/
/HdIxD0IWyosQgBX9yjXHkBjj1Gns8hMxmPdjmC1kQZ+D7pPqREwkBc3EXe2YyBE
t9Obk5PS2UNapOmS2h25PNtTWtwMBxm45hud2sbmz8N17EeCQanlBbZPUMlA89Zl
bOnlqh5EBXOU/MFUrrB5c0w1M6h3qYEbNpnjJ6tXQmTLXKO7ZMAes4CODmGxHU/L
0oZ3WGYaEQINmJ5PNoG8shzZs9E2OPSGANbp9Z75J6EHx00ieQvSZLao7f1Vz6Na
H2nEwjIvkoKFkbr68zLbFHGn9eZnR2peSsxcxtBfpQWhwppXxvt7qE7I16ja4gfM
2dsmhEaYIz0wQOKuH9g+xepT3n8jLU3dxIudRa/mAiikAmDwRYSZjubxRogl9HEM
hX6FjCnAtgwTUEUQCeb/dcyTzEt/XI7kYNQZpYyVShTdUJuq8BQ+ocLzp7heexIL
KlSZtUVv+8PYQ8P5ryVdF1lqBLD4TjyMvs5KYAzwbds1cBnoBXfvseLG+X9VpwY+
AOGwZc9r4NRx3742ucHDCCTOkZAPD9+yl2oDh5ZGwPKZq2+126SD5WZy9PBcskR6
IMmKf8lChsQkuXi3D30r1QMc8uzQf4sIFoQUeFbHS/kC9Ncb4CSvWOwv45z5TeXt
RsDdN7OfrH7kdsO8vDHpns3bAVHBTzl3CM1r+lSWB6BuVrXkAiNZFUffy/F+qP5c
DVdQW5Yz+WJYp9jNVptetmvGwzTJ9yVpHhOaYD+vr1aRf2zsuHoDtKhqEkLDOBQj
E2gW+17EjikcxMBNNm93K32iQ3c0jUpClQcZ42habp6/Z6arja2ryp45qaGAjbc2
ju2iSzETzYOFLOFvstAfPhf96fnm2x0aVQxrA9SN4q98YwItJ90BubP9X27rFtfQ
ybZSAvVe+N6w/+nVluSt8A0VCEdZkUYLBIjkZkGToo16fSiwwnRWyV3g6Tlm36MQ
h4k4DgUD71ET0l9SBawPd8RzBy0M8e5b85br0f9FLx/grQYfiych+PmSmbk/IP0V
VsAeU1BVPWxCXbV0ZcygKqWkajNhst6FuNwnGZA+gFDMvauBGXrBzWqCKyMb+U/K
JL/GAzDIj9ggBGuwpkp+uabIjO4DxOmdaUFjRtL20Yz2smWLDvmVBZRXO8zK1qQT
pDy2duRrLSxxr0N0v7Hr94IKJ+aIxTevPH8H8R8quzXSLZ1lAMR0yyVQbOCKdXUR
4KgYYVpa+/JjRUK3YI4jsdzmyYeBeRWMpKkaebfFuKrEvj11F8yfY2FAaNP486Qe
OnSanr/xtHqfKxorTD2mkaPt0ohhjC0Le7n7s0++0kk2rErCMBHjlPhinHKZspy5
6CaH0N44O6aNrA7KDb8a8s9kRuragapDfvkRUwvrqz+aN+7iQ5nokWec60p2V9yb
nAvx459zDpAB02RICjx63+EZ3jvtScFN9AleZ1WbKHqPy2Y4RngdVzQPWlvHN6lx
F4rkLN9FpQm9bTd1iHaCy5efOZdFvdAcHz8MVeTbRbEkzonKTVTNp1AXwM2nTmHn
kkGaAeBRkUCupgKmeLcIO2guJN2kE4hw3JRHa2uy+RfDWrTxBL1Vw8ZJD53m33g5
frluUKC9YN/MP5IsNr3oWqViDPSRvEVk95H5JIrarJPuBQt3fDH74qEfGnSMjRlN
Q6kDjifeLW/MIWjaPFMPqfOa4qD5O/0Icnn1vAFVY0NkQBZ2nNzWal1p9T/E5tBZ
NILDZcSSDNwUpcIqTRMUoFOmM8xZpXMNgL4dw4RWKylpSQQvMq+rngLFfFaRaw6H
ltZRqZMM4okCzFaDeLYECEg2aTEAs5AGn3N24I4v4Zdv9s3rA8kVPN+hz+LU+sS+
fxg3XIcRR8DZpV5pzWEg+QkZrF5s4TvqP5xV7rYcHtWqLB9HstQ9oO8HPR8UyjPi
jUElqMU80oSmLfCA8ErGCx5VWr8X6LKx5r4HryNBqrDPvFkgeCSS0ZGOOqOxn7RU
sKUxHvmoD0bREUViz9wyl1DrOWFMprg8enohqyLrjSJ8VUXpfrR6be4kzDCw+7uU
JkOGb3zZ5uJjKayyXREhmAhjNEMjH9D9NUuupR0mXFdLQV7xACtWrCg9aCMOF96t
U+n7gTAc3WERXr/vKMF6Tq7d48qCBDxGUeEE8SpzhV1TIMh2NkTFvMTGz4Plmajh
1OjEhuLWz3LXmkM+scpCYnocNBZyddwCnkhfsEbGTDoAHg+L/7cUVNIdMNj60/hk
RxJerk1RSWCqVXvZMkrptJlMcoHuFHqZJyhPvY8Hrf8azf6Wwoo9oluHtwf3W8x0
ObYThMoIFn38A+82xA3b8K1xEXoWMz58RgXt5kQsf15aP8F3z26D3VKnhBes3U/w
JB0qS+mnai27sZNj8YKcxXsCgsd2q8FVI9GZ4eFo8krtcPD6xlmQecZGve5FHWwm
hXfgbCFMfzz/Px3mN19sc0RWWqbdNq8KF4u2CBO8qP/0S2thc2gwfHiTG7psWmZm
YXsX5z3OUFeUQlzWUP6lRXQmnseSuwHNzH8lJ4XHH/YPpkFErIjPdjfICpOsNEDM
KYek5PUZBXL1R3klxwknJWv+XxEJLG0LxlUH0SFpv0C+DfuPncHkqzBOP0DU0l8Q
0KdY6ZUkr9HTpm/Kz2EuEbcqIzWBcN2ZEqW/SthXUGmPiPOCfXvawUgJ5xb1pRh5
FSM3f+fHIsYFfvTeSniIDHwFjWNwKxuJqqWOvdoyJjG1hPWxsZ7rx5F3X7Dah4J7
Q8GKK6RYXs+L7OmcTr0jVv//a9uXtguVrLdz8ngjP6qDf1dk9Q9o2xzQRhAiFgiw
d29+PTj+BpHtpv9qgF9M53+bTJKMCXzEpVo5R8PjhW698s9fr1D23xLrPFzuA1Ed
jVfP2tpSdrHk8CJaGBCj9/Ro38nWEisJxJ8LwNsJYn6FnPNvAXg8XIslIL6jvd5v
tUGvSKzsfHknCYK82yjJOg81anecr0zmfo6pT4WUgUy9l7bMJps+BVsqNi32ubrI
GAbJn4IsYGiQleafLGM61WdsL9oc/q22gh6uKWaszl2oIU7UcrDDKnLo2iBuXY+P
FIm2htzTtnCJhaqgGr3QrRg/gs1HSqrNypgdBz7pueT+1kPxi7Sawd/F4kKn9bNw
tMcLJaTTtq7Hv9AkWH5NCLg1yAjhvJrlVUjH3AH3mGqiQxJLOQypcwfpxopCHOUK
zbOrmdZMqaeNqP4wV5OB8c2ZaHnv8VbJjjkQDGTQ2fbZofSi6XE4X6zyn97DIkSN
rF8s3RxMeGyzN8qcMsgk2W5WjkTjHuEkNMpK3SiS4b9LW5M8e2p0L47OGzyzg5GR
5+MTiDDyZqHvaFf/CVJkTEDq8/sHEQ+spccbnY22VBuN9zyu4WQDlzshsrV8MBMb
bx3emf0s+QVXMqGjFo1eneJCgGIEG2xK77E5Mus8zaDmJRLg3GAhiUS/d+AoorV2
6nG/pHk92x6Q3moEjmA0C9UmXmBsLjww8JUjaE7S+D4mO6bbrIM7J/zV5F+l4GPo
cZcZIG0TzKEzS9Gv/yrXttEySoY+yWzGyd0ZzDbfUmV0c2tyrEJZiXcAnywRTe2k
4QhzDktGNhesGFY+JUdPuKUXbc3aRwlusq4QnsHvoB4lDq4fdKcS9vbBTox6f+YF
LwGgqKwSP/cGvEZi9cdDT2k7rg6kxp2wSzRBB5of6LOVxM41YdPhwrGPw29dzzv/
k4bzlknXof/m4slJrWV1H0ozfSQr1F6d3Un85a4cQqUXVYlFC/RBBuFJ36tWFRvT
Dn4yEx/VJD1CjUTnNj2R+1E/CiGegfqxXe5rhq0PtR2vmp/JhW/fyMJDZRO+XOog
0qzmOX8PCIfwXWU/J3tuAW7OjXuaYv/DAa5Ab7vASyL/jAQfyojEaioDstOQFRdv
8uq/i0ca4hi8A+jQ8Lh0NFHrlZUBScagfrQ57HRWPLyBOvooMSLcBmfMCo1d2Ge+
EU2OZyxvV4L+jBAr9b9JdVLooL5vjhH3bPNttWNvBpzGktP8jkNAzpaxsWvHX8da
wTqtucA21oog/esxNLfh7xq1/enfkXm5nQxE/9OsyBH1NUYjx2Gyj7cLGvhX4kvV
fDSUA3BGDKBFieOI/cx2jttnW9DxD06c8wXV9rlbRoUllbLw0VnbSnxKsjRLx9CS
pW2zVDPPDFNBfKrTKjQsaBU7R/vENFuvcr4NFPSBIF1ctHThYk8YMSsgWNp727i/
vRuszTvFGXLTYJ03wnvV9pAkzaKiQIOg/ZQddHIUtqgKX7Eduuo36nwL9IBkdtmL
KRJ0SAB2ocUBm9icF8YoZGvgJo4vcNQ2Ufu2tLKrPzZhjoqtdIXZlyyD4nWEj2Vn
h+wvnORP87mKLXKehkmY+PezSlfbG7BlfYQU2Bid+CAdbXJvUC1vSD1Gn1gO2y+t
ZLm0uqkUh4gXWLHLM2EATbTJ3szdjlA4dBTIRbPNJbgok3IURrSQmdCTN8RjiOkl
0nLXTabEj69uNLpCJxUc9i76PEnoZv3/+yBXa7IHYuQT+uK5Alm/kedaePdUd6Z6
2lLoSPjrmOy65GyRHInwekf5Hc0m+8CeGnQfMl2ddPjBaqSlN2CSjjbOxAIf9Dif
ItP30awh1M7RgcYnfNW9VkE4SBUztNfHt99IOvicNId7k8vJVXSClp81OJofb3SA
zjR+E6Kjlks62O2f8GQ7Gn+bIS7aHygyFdxMIyZVpP8KT+AyUTlcZBhLb5VmLOLz
ZCn4AqHZWFEeSXo4ZNbwUdJQ8CreNUXXyyv7Q7hwquFehTWGSvOr5UyiawjxyX0x
OxtcN368ixt/xJgoiupIb2AuJma/ZeygaW3AVV3dHYlsrEbY1LHW7HzXb61Cm/YY
cqizDjfs28Fvol2Ez3Gk9BUqkX10ztV/VpFAkOqd4k1ZCckBmh+UAyW0ULILUUVc
rAgL7OuqXPDQDQwWOf0iv77giuTy+neFWIyq7B8usv6HbZGtpp1DwpxbrH7Bl3Bb
3yHpso5ziQNW+ER7ZplO5NtwefcFGgzeMUhoKOS8Ic925SKt2VnW6U+vYh1ikeV6
uKr4MdSZIU0M90Acc3wWgXezwp4/8ez3ZAEyRSFMRH8MwGfjr6xacWWFhnDeAKI+
Q/kfu7VuT1TaqR6VDQfiAiJeHTtbDVU2aKm1OILLj1SVlqeS2PErNtJIUJGxP2YG
Z5h6Q84aSS/bOxmDHktTnQ5lsJaDpB7njryqaQp49QbyJTCgXY6BFa1BHNZvcyaA
qTwTCYiwfqiNVP1Cw7PE3MbieT1fCiRlH6FNYjbTXlPc0EULILwj66vV7OlFG+cf
csPdEUh9ESjwkbXr0oOk5mrILhwWHw4FihW+pDkUjbq9Bj17RhO1UdSjKf2Zdv8r
vHvHTMuaXp9OHFVi6nlreUlliSeIvcFkOEC6rwnhQXUAOX5CttjQz80piZczc8zc
B9WZunPxkvnGbJge0cIcuUOtrmOt2E1sLAysdM0qPERI5F4Uaq2vYXMLxutSJVC+
N3EC1oRdyabI7Iu8+C643LgKRW6R3KL7JCLQq1GNCtjzd5F42DNOFC3Np3OOIydU
II/fw5HIf22Lc5qtS7hr5CDyfPiJ8nHl7yKRKApf9t+risiR0PT+q7mpekraVhgm
iwb0NlV47r0ElW1ikbxtxwGNnpmV5O93pmNCtEV4mCNGLMH/XRDRamOh34Zshr0F
q6n3M2Y/RRUys3YS05GAPcac+c2SnH2fRioTQzFjkAVlIoJdTBDwDXRFKo4WCKX3
8t6FdV8mtEFm9WEn8U+Jxjqs1CwAj9tT3Y1gqjo1X6C0qYjDYYkMu433cQTE9aMo
y8l6XwSPHYyr+qPibfaIv3Ew+7VEzFYoDmgkHzqfgoSw86BUGeLsqs21kgnMs7Wv
+kURtFdubbkMM4Zbgk1XQ9pWW8A/TUoNJE8T4MtXeIsVe0Slw2j3dlGXuSfBKArP
8bd6434YnOkmqVQP4/7xx6uoZ9E5VHQ2HEDaHGk5gRUNZ9yzdAGg5qJmYdH3U/gm
fZVGcGZdLx9rBGTj78Sxx0uv+4yK3eO60rYr/nQCXlzS9i/6lFyromtynSylgMP4
N7DCGtAkO0eEFNfJeIUSY6206LNrlwPVgsSc3v0jmJI/TLIj42mU4Nz/a2xEg7MG
8AG3Nlw+JnkX3p3VqNShjtjQFOVPRt20h9cs7FM09TqUH3W2BgzO8My7AKS+tA04
vyrcvr87vHHnjPW4LF34VRJW87S7N/YbbzMQe+Nmndi1QtOfB05s1Ux/v+itWXxZ
A7pw8RXMNmJhfmoaDmyVHmKWLZOF6PoHZ7vZ1mhh4Fp3Dfrl27FchiB9inkQ3v1E
tL9ITKdz6HaCXlJLO5b/dAWdTVgwK/NOc2U+rVjilXPGXtAYcqNH2bbs4gCu1/Ck
5FvpyBv+4GG1jySWflYB4bY7UmkiaWmB947FieU/NRbdoTSC4jxzGpwwAQSnbWih
O+8wAIZ6saZ7OSfl25Pw5MAGh0IIAdhBVdZpw8vhxxibfp1KsU7EuIJLMrp7SGCz
qA+ZfFBp9C1zE58Js4SGaKvmX3dn5ScKx9hnMWZpfuPY/MbHNMCzJNZiQxa2fU4A
wC4gDh7lH6udzaLs2+t6YWLHeiUJmAMXjoBatS6dNQ2OrbD0mX7NhD6Vr0sdhypk
L22xhozN290KBmrumH85F1CWHCeYgKkkKYzqsK0Hjbt1WtlnBnKyopmEVvayvvHw
7DMa/y5P947FxW2PhLpgxLtPQKqkz95xvA3NYpCyF/368F63JQbAVEsGgUrnn5aO
TMHCAEDN6ZoJsWASQO5AQv50IA1KTUvSiw2RZTKZXRVZx+MvPU+9ro+e8altN/s3
lVNQHdQrvfHEPkQSyBXEBQoicFPVgfllEOrygHOZgkAL/msvq/QoDFtFAXuLG9Xe
+psqSIbLhUvON8ovGcSI9ACS4aS5jSB2aoPJ/JDSFE1gqcwCL0uSigTCpjZ3mpIe
a7NoArlWwjsJSBvKSLre2CAysr8pYJrcvAoj5+ypJuvBbEG+Dmc9R89y26q1LQkL
LbRtYhOoyh8INMDuWRohyPzgPiAUOjxnQVdU+hZvG3pNKcgPwjS+vVWi34MssnBo
koEjbrXUyA3CW32UNDO3Zz7mQUz6Jvit1Z1snPG5wtwGeaq1t97hNLcHXDFH0w2P
kmVt/AFO82S0NJ+wY0iE9prjIddHL0yTBQkDbm8lggyMxqKsW3O4cWeIuPeox+8R
cioD3wHspNNWp2gPlK6HPTVkKSbJtrtW+q9KqihOIyfBQQEekgNwTfGK/SCSXiq7
5s78DzQiqbIjsECVmj/Q0R8lwXLQVHvr2yn2JNoZE3tZrvS9Hmv4+Pcw41SXT+dL
XXnlV+NmAqE8Q6DAJjBCYTr2G7vvrxrcWE574dZ6v0yljkuJLDUVIpyLj9cst5aS
Ua3AzcrhXYRy5Sahpv2/fRYI9c3Yc74QVu3kJwdtC1w+gQctYI+6PrAQYNSQG0Vx
3fWK0KiAM3Aw1aUk9+MokUxNr7nTKGUvlzcdR/MUFmCa46lP0eiSYOY1SIxb3aKu
AP124N9SECg7VNI7VMQXBYkfPzicroUoLPR3mOgHtLpcy08bREshpSXbIXOab0i2
6M2J0YqAfJNmQmSxiwRItkuECSmc/QT0L1OjhTVpsqapJ+l4bSQ+eCGg252yIlVu
IBltiNh5Dhd1qUTGYbLI7K+C8jiYqS3tPSY9MthllSgvnXB8yG8vRwhSmZCmbm3a
3E2W10bQbzjq/3FvgWOT+WnR+biEqP2J07Yq2Cw23KDp/g2jkv5FKfJyJ8Towpja
7KgXHQSaGr8Z8bExhlJEG/LRHIa6lq3LVwUIU51a0SyzSfWT7gDaOzDcpEc0WYP2
ewQOSrEjBkjXKsa3KCbdLxHVIa7xS3uAMrC+Z6nmnwmaXcuRWzg11Ywv9vdKOzmK
w7j5/Pq7igEzGa2zc4+4QGhofn2J6monctJW1o9rm62ac/RlT1IVToxyB+8UiLod
hcuuuDc2amZLiVcUtoCpACMC9uqlYBGO4Q+dsGS5oolKlv7TbO+THyi+iDAfFb18
+Z1QFoguOPQxIiixO8Ohy0jfVV0Df4E+paphZ+wOy7FTBTaGm+t2/u+a8IcVYDyt
H4ZsiZB+CZ8y5ENlA5B+O+iyvx/sbhu7y1kiap5u2fvmA4fiBwphO8AUHKxLDNa0
QHc54O+5wrQ9zoRhN2/LDIRbYYbjok7x2MX6RzL82pu8oJtHSuiRkF1S9Yespw4y
Q/YA3LHO0KmJuSxwcnkwl7YGqNoXKzpT5YxSp9MEH2KEC8IEvWKaGhF5q4FR4425
RicDT+n8wmPeBsnOLOozlgSgxqs+cQmrTySa2FrVahQvOM8Sk5SBCZ74xqqVYC8p
bfKeTBC3/TiVXgPOoTMn8PunUW+aCp4ek6Ver79dGl128y7gaY44IxYQZXp+hyPP
j2zpbrgbZBSERaDcZvWAAuBP+VmgW4XxQlSdI/40pSS8Uw2UdMIJZvPquXlTIh/Y
jhZ+cYbguQM2s4o36B1dSBKNifYi/chVXOXuNXB+L6X1PE4+blvW6GYMY/OXsQ8z
/Kq1EaLtXUTKxr2ShWcBMptAv/66Wjd6TGd+TW6gCqWF2eH22hHQ15ToQ60zNR8f
EAxQJxUxcI3yQXzeeJ0wTlM0+0tQf/MsmMpXhxBmvJoWhWDhd2Po7mroMwrlpLoE
XCADdkFIMk6U9krv2N82diU0JHXm5ig48Cii7/mfs2s16ldLmLOSfWKOS6yPH/uM
SEQOSvLE9pMx47uWb2qi/qkfFR345ILTHWyIz1HrZ6UC9TUbc+dEjnTRME4Gz2hc
n/A2IuWc9KWhdzvebxl53CmRGafRk6uuW8H8Jpkonz3QzqhoUtZbBmCVHrLoALbm
gpoI+suP968yl4tqpHnhuBMU+0NiBJJsJnYn76qY02nW89N6LTS8800YHdSJsPSt
flxkMMHo2vkuQdXfuZEnsAKO32wbVjj4Bmi3j/TkUvdF7WTJxHMOHobjGyyYMPYI
v0JfKHFW1tn3nw1TvdYDRzzw9tkre1ttQpTubiYePM1qUJ4oK9oprB38/jx+9PxD
JMD+BOD/k6BwNYLW0mDYRWmY+ERu+DDcTLM1wuIEeSVNMsO8SXsMAbuTxqrK8mfH
DxXyRsw/TFQOChbrRUilYM4jwcaVyWAEyqAhZ3QCgKkDnaNKdmmjGnc3TeM4Hkf8
qdSzJDuqRe3llG2hmJLeD6snTbIntFaqF3pkEf8hTn8NAlktDRwc3HQCy3bMaKiw
zbjEk4L/6XdCWUmKGoQdVg0MWywtzMBZt0+hTAfCtaDtnU9U5uxaemj+D85siYu2
91I9tlwoUp9hnR/3Ub0bShDer6qiCXvEVJhg7e+4dUuB83gqNO/Xk0C6IMt3OsE7
H+hP2Snv+Bj8mr2SHgroY49JLyO7c7NFgqfCa7jx/7ohAM8LTPqXzWm9X0AG6WbX
+bzmDfd/dDwTTzvjiP6JuVA97RwcZcEpF+tmEqZAD3K02WL/43ATwgMzzdy33fRT
bOPKmDj3O7ETSYcavlComvOQkiRvEj3JQ15Fzwp4d5VoZxRmtvp8o1FuKc5ruU2t
tmMvLNAvOvxExgW6p4UFE4Dp8grTjwdv98VfGMYBpA34qPkyb6vFO8KO7dG3HnM9
eI7Heg/kfMhkArynllX0KoaCKYk5GHJewGmRnzR3tG3wA93Rf2fg59GBOn+KuRnK
Q8iOujU3eBY0OF1/7DqUkVj5icNmHK/tvLsJY8uNHK30n7n4ifHcEaX6WOgmrjwi
HWQlg3j7LM3ucsroRtCJQBbBerXvoJzdSF8QOmXIF0Xj4irL76kc0NfOYnXNqYai
bkBfbaQlENcZ6QXmtlaG8IR/Waen7LiXHPnxyT3so/gsz7nqL0bv4dCSp2+4spoc
mFTnHEpMRGYOVOm62ZekDud2fs6P/nSxRoj4rydutI8DG7imo3brpjvU4ccaKNrw
KiKu4gTQSbuNaukAhfR4IUaq2ZvEBNJPS2u9KkSwCuDxCzYD3Q6whBnwDRCA2KoT
ZgBckduVFL9qPJXT2s9OIl7mwAQo5BsJbtsXK7zLqefWev60oea6n2NRYUMxTuPX
rQyyexAq0fjUggmz2vD31onx+7JHB17JBOZBo02cfXRqLCZS7vp9wN/+p6TY6r49
3UEFIAkmJ0ueCbqza169FKxmY0NFmsarIQib6NuGqQUDDCld6PfF4rs8O52dXEA6
hCGW8Uk3AH5JkRWJ0KsFkONEgVlwCcjBSbNWCuOOh/cxSYrZo6Njo6+ik6AVbvju
E5KK6yDmSVJIoPZXMf7PfNb1OQdZVCTHXMCs5WuL9ETfRGHahm6hLV8wnNMyzW3J
wDt/rnsU+45gNVZsw4QAt6VOMNophgWb/CTBv1BvrN1Ck9bEPVjUSyazZaAUWCWK
sLHqZeEo0avNb8agJ0++JWO7RuX1OmpRjjTYoaB5ZXehFIhK7Ld0lmzIGjxh7m8A
YhINZnb5jU4EFIG/rM1f7YU0BhXB6Y881wns0nsIWJAvH2/yxKuSjxujnd6BrN0M
i+WA4O1QafHhJ4lW/E9ic9pmp6CDAPp7FX2M5vV8Gn2RlOl8rAe37UO92Acw/Z3k
Jmnw2bRRDSIwD3GUDlAFBNRr1KtlTtSxS9uQI0IveTdT0FinzeRjKaqc/B8IkCg9
Sq4gDSLeAweFzWWevWVYPg7NK+Q+YDev5HaT7KsShm/FIkjL/aBqrMGinNh9Eqwt
A1f7fZGu+JpSQOPzpS1EXehrOmZhJkxqWY9nf5gwVhVQQaDs5A+i2EtEkAmGAiPe
xZVPe05kP+BfcF70i/abAfq92UaKmBFzIimAPmkUYm0HU1uUt0ERKFPu6pwG6RKU
VAtkrQYc2H1357Efu1G7s7qzwkPgDbxM3aE7VN8uVqMbE2C5yTutJhuXCRe+BZIC
nA59zyBd3Tz2p2eD/w4yL3DQc4S1c7EG3nR3XuP/fzo553DMIdc2tk3GuGsn0Aee
0T6xijshyx7DxvPrGTDPxktMkOys/+wSIqrcqJ9OGLgDXksGBMgH5eJxErHXPJHl
69Lb1XxZcdTHlzfYn8Y4MBdS2l9s6VbCt5obH0fkrvaNb8VdmRQj0JdsgEiAP8aX
k2LuRZYMYQSufC1XYwjCIVTjBC04gCO+FR5tpzN8zineYmERcxPaUB5r5pKu4AQN
t1KzjoiONIreasooHi1+yVSSX0RTrPpQXPJgXYkA7VUWMQQNSwgtse6m8Spel/nw
hQznG0eeS5BMYx7WnStHNdYypvTESyMoGACLH0bp7cAVIjIV+syPL7uDyCQp/E49
Vp96Z/tg/ZIVh2XQDow6XALrp7NrKV6G0q8xkTEvU0FkRv5BS7k1Hc2TL0Lo9vF4
I3Md4RKNI6G7zyXztRrom2toB7s6JPagvP2aK285UIxNzqHgEFSAYQVEAn61iFIN
TMf9NgNzzWUZV6x3Q0SOYFul5DhgcBUmZ83MTRxdu0fkuq/+Cca9CzJ5m7ruZ+iQ
L8tCW1bUNkKMAfeFQz8Xg8wJ+mr/dQ8nZhd6UCnZH/5u8aVVdJ352vzoaE2BxJLX
/MVFuuF7yP1j0uRgldUp0UmsdWi66GovjEx/eSizRQg+wD7kP6MYSBhjADfcWZaY
w63owAVaphNBv7HqSxTRXDG8RMYOuf1aYOC0r6DpVNEftNffGxQcBp24jfvT1a2J
dbpOf2XZUBqxeQJDk529nBg2k7HWzTRmH02PHZfI2Iot/CaSfUBcT/yAN8KF1K6C
B9D541/tFT0s9D7qCG96L33Yh1aVR0HoyjuraHQzvJhLQlPPgw83uM0/T3bNyZul
lergNqpk7tWZUyFXW2JFCBVcqw3RHsM3U4uB0CCNTX2WjQpRnrR+oVcV/wPQLAA4
by05LahVUGUcQrWUIpr42FNV6kFAJFfoveYSctovChc1LtPeEBBb/Bvh2QnXrMds
GkhX/9VnPpTPOKneOjTSALTp+adLaX/A0fZ4ROT2D97mS+8xAAza4hf3FsaZzSAH
RwhTRtezaNb2prhYTDnOqRxMQLtEXdDjJyLGvLj6SOvyDHNO0HYCzq6xCyDW+DtC
/3NeVJdhuaa28iKG/ZDvw+XhVHc/6j6QL6JkoZcvIosPxQwae3Pz4QuZ/dwMoJUU
evgolxPJFG7F36OHU6lsvV3lGDbE0p964xLh68ryuzUzOObA8pfR8616GKLrgSND
HxhcdXkQ+6tLwIBgY0zebdheWSEdmGNmMOLDwB+AHjrwj5u85rSli66gxHAtvncH
8Pj3d7NvTWjHO/I9soLXywk3jKGkyRyvEu7BAkSnPfhNF8G8Pf+Th2TDFQJnwHdD
VX2JWJogPbmqWjA0pcpNQ3HiDiRsYMJhqGdDXdP7kUH48dpHDYqw7hpeXhiUZ8ns
ggm7Acsty2uhncsmjyccHNOK0hkRJdifGDi0WPYgfVzSs2JA9ydWq4T3n8iKMln5
4Uyb0EyQsFlGXxMemYNxa9n96Ry0B1XSvR/zKV6jBjc0c3T994xhLz4gzJfZtymc
6S9EMJwQUlEvsCU6dy6ba2p3Y4IBEW2speRea4Xb4kJ/ph9swpvJ9DAuvJ/yOtNt
PlhSfCc7Lb50oWSCNKJjOefGHDaX/VPuxRQg8uyindHlf/4+o3HSqALuZp00aJb0
wlECIFicXRGcmWzEuNUL4ke1HB0pUpBMdAgNeR18fxwDezD0Ek5dzAP3TSQgq4ku
DaQqp1qAK1VRcu/aNdsI3+DbRCR/+MmJBm4Q5cWwcJ5eQX6ihbUJnWTq86oQiCTm
2PbHrUOVXadPQnSyLH91b9Klum7gHn37giXDp4hXDuNafeRC+fp1FvBd+tWI4qiH
Tg/Ky4W4HHpo0cCVIo1QVD5XQ6hHkNa1Lr6gDEZ1AwGssKZWw6P7evaFixgxwQKJ
AoIWfzVQ10BmDUuhawwW4WePjKeWhFFxP/60CNpd6do2liw6pB9CxZ+zaHLvVoL9
IDeskEe2pkgaBVZCpNvLUJsGD7Nctbb3pmtaVoWNWFwxbZfcZjZ0G/DSNAcnQhBF
5n4GqxTn2xWyAnUOOc/t0CLJWJt9ZjFpT/p/gcFcceu+fWYOoFhJ3+TgAWoPpNnQ
kjzRYJo7iVcfJ6e0GQEP2TyRHGRQe08uvDQEn5CwQLL1T/MZZ1uXo73rSFEwSSBd
KQV/U4Nbra8JaEgP5pMwjv64Ov2MusnFLVASCoeEzBkPXU1pj5uIQ4iGuyBDNg6e
QJqB9JRbYvaB2s+v789TZLxff7OHI/7W1uWZ+sjLle+UeL68zVKgSkgQU7WoKH2Y
72+2g8st6i8j9wSE3ieC4S/tTSk6lsOxiQSeY+QCDO4GUJoKcb2xbSaio4m0Mime
dI1f+ufctLqlFWIYdE9gKjJK9Fn8JUntflfD5VdCC4XG24kCf3aie0OwsiLgWWH0
PvwnYq2yIGZJZODJ7diLwzS7xcxP8u1wSqHu0YFf41NeIoeZXQPe135SHZ3vxG3w
L/v5kA8Pc6DlsktPlk0zPcwXKcJpcpVYyx7twB9lcvG8Aid2GF4dlCNz6qIjexCf
u6u3sebxmYSYhEuDS7oz9LUtf8ia7QzWKBSfCbMuhf+p0sVQaXoicb8kfEqX1Y8N
IV6CjbpcR1CF48icVDewR+uEUraFz5v1lNaELLBU3G822gJFkwgkVT0NM2OcBS5t
SKM/yB5p9bFghipEHY9xkpYK+AuLqH/kM764XOWoP8YKrYLa3g8ePIlE9jYLrbDV
SuSVPC8k4OoHnE/5mmZpp3AwLncPDVjGXBvnzac7Yy6WWBrKH6LMY52qLXKgBF/Y
hZvygWWJyONEyyLKm30Ncc7CVloUuVOrrdO+FiD6qHgS86laIO29LGtOu0ug8Q7J
SqVdwpXYzyHIR8vnjRFfCGbcZfFORYoMGSi+Cg6GqCXmPhl2X/a3LeD6Mz+tb4g0
V8sWwSO362kZFpD3ETwg4Dg4+SljGaTuqYaxA/oeHsB8gbN+hCS7CSOS/PZpil4K
Rc66hvOEuJjsizT4vVFL4FFHxjScyi4ymKz6fI1FAmAnahTqPc4hlMFIeodbDZZl
UBoN1d3wB0w9O8eqtrxrFN5a0DK2/aKbJnsnotZOT8QOhRep0NrxTyFypmZmH8Kt
Oernwv2oi+jVkJLZOoXGb6aSTMsEI41PrMxfy2x6gYyFXDJnnhZ3ljnBWLxSxKsZ
M/RlDksu53bqzr7ASmo9nyGJUIpJbvsfmJ0JK9u86PNzoPJpuecBlIijC5pXRUsM
NQYi5oen3XNCX+KNP4qeMvaAZqGZciTRQrk1GDKz0K2jp0pQm9enY+y1vx43fRDL
NNWqGmJGSh8AhcmvoyAR0h9YPEK3PPW7Ltb/6Mt7RlgxWRW19iEKB2fGtqZVbKBv
oRz9wlhzMD50jxMERKb9Qsjk8rDOF08MmyFLZPRfW/sdH5Jye5FoBgm33B7bqyQ9
W4inj9EVjpDXg3jhjst6iHOh3tYqe6vldWCFW+LFyhnKOFGryV9eK3hIFzSD8RDJ
LzgU0rFAvUmQZSNzWKglHvTbgPdOr2XeHK18MQpZglfVuUe//z7QfXolNfHJSDDj
iNlmUsBgFdgDKrRMP2QacO3aZ9qAjYhxGp4P99Sc60gHBsIWjCQIyLkRLsGmsjkf
Mk7is1Rz0wYWM5xYfNGefFMM3RJbAvfVmQcud6WMrftczAimKG+7qZ0aStV6lGyj
9oXVYD+BmD4fCj4Tz4/tn4xEyewV0QGvrGa7JgZDXq8Z+WQPaAlJcL2wvGhVjUsd
/Hn19sb+orCODjByCia/wP9HRdLzv6dkvEFzun7Y+04RDLXlgjK3EjR6klOLj56G
fcDPaWd9YH1bqFKo0SxyRkrgF4poFDfqFBAbB5NFx2DOZNuOkVTey1sMRHnv3zbK
t5zuKviNa2KLwne3YlJfFcHx4PoJxqlEAQyy8CRtmPLBHToBPsfKDqsKNQek37dH
0AssDfJkiZfpxQvt6Q+unHObvujmWin0NWlTbJKjUIkEde4C9oC7+J8x10N2B7Sm
F6GR+VsRD+31SgyYikvYYDyQs+tZuJNHiguFVpsyIIp7ch9bQuQ3ZXlbeiqUXWYn
P1EFeLSqXoSUFflC57IXVnd5LFNUwLugfGNulaJRW1MKrqVgNVP57Wj0C1jJRuwi
b44agx4WWw6jKzyNduLBZ+Hpfcinviqhhdmbu0akK2ZnyFHqNMGp1w190G/pWayq
jfGayUX6Z05+RODI9HFXGJg7fez4M64NZhnHXq0X0mdKpVjl941Y+q77Y+Bd/BnB
KrILSvs89ojJGcwo3JFwAPaIoOiRiSOvj2mxcjjujcIEl8Ch2IqdjA4OOQdzpaif
8nLoSjvnE6xdE3XZZ68qUa5xBBGAp20oD1n/BIVCGH3cCctWsr728csnFVF4+xD3
2bBxKjzQW4SUqy78dKsK1dYBygEnQC66yaVYeqfnHO8yraIz5vhAgr40+hr0plvF
WdMdnQEae6/3jSrF/XaRWD64BvfQek0n2Mn32WsBJs0YsIynGbmDBqmNOskhJyI+
TbmHkoBgr6SvK8v20ge+J1HEPreD5z0UTn2GKVoJiEngw+IjNfbeSa7V5d3wtD1u
vZRdfhT13APwAP5NTWwYrVkQG5F0UW0hY+herGKlzXYdXM/+Edm2ih3L8ZB+3SP+
8So8v9/mF3LQeE4voEQbhQcFmY9Jm0ZfCNUPQy4h3x09Cj/30nSKnN5zsl/J1u1T
wYuTktCNF/mtDP6XifX6/0YGhyh0DEbDEXGF4u4rS+TnSqDkB6P3Cc+1+PNRAE0p
6eU+wUlnGOAr/Is4HcIAjgIUOnLVQ38bxewdSGuY86kiWhWHVrTB9ONaHs+lCUe0
uxM1FD1IpmKFNi/I4wC/Jm63begrlRLKhv9yb/2N1GanFdsGo2uLN1IMHFhat8Jv
q8KFQ72sH9/JLF2dJZrEhYLVAHSeS8abVXw+PSjzsM0qYqLy9SGTQ29KGgY9MAM7
zPdDt+Of2buIv3IaHUvWU3HKbfO7GGPPb87WOSqSwiZrKxjrIS2m2Y982epjb3/5
E+OHRucPvdNRQyjF1/0pjUqHNEA7+ngsxIwjc2C12brOxyZ+0jeXGDq16s+kmEmt
vqaQjrBgGSPQ9+nC679ZkHbkHBYWd7Ih9VKQfRi5qwbPZaJDT4JjopzD7A5PI58M
dKpZIfiYofElJhZLc0jF2EaqPfFzkAZ4u1X3FfX8QzeT61y5QRx6a3HF4tc38WF3
J6u1Guu6iFFMhvudwQu4xhRF+27Qo3WpYr7YQYGnHYeHK84pNbNmY5QErvq4ynT2
mL0dFhiG2Rkww2flNuzvzXr07rSOMk4H7TRpPqdDSGIvr5WSjs9OYLwtVuazWKxQ
t3dnQLnqRpsd8pMYNu5q/j2lJu+mEcHWl49z+iz2rcfh73D5Md74ihiV4xioNKsR
cWRMB8A82idkn8a7BliRXAneeu8ZyhGRt0S/PlfNPifdhE6wgYiRImc/kWuPXXUe
fx7Sdab8yVbHeCPoIz06C/ehVVwn7CaGKrrlyKno73d1KD5TuGkYJugzoxSiG5Cy
7r+qJaeaxqLtDzjkQ4Nv6oV6d/SICvDPXlNU79i9lIwWQ8jkVwkNQKBDWeRuYHHu
WfkzoUjQsTGvmvO7dWId0UFqEzR2yKlnsPvjRIyAZURjOlBDlRC3QFx6Z4WJzpG8
tW75O2qhxdblqdr18EWcmRWbva0jGqAA0e5s6vhYyTmR6bbGTIBrVUFvXk1caQMV
CrUx0kvGu/Hjuym6e0JX1dmluQgJLjyk7EtyXHQdw6Q22zj6rjpdwc90FSP5EHae
FUVuwMjjmlwkZPvxZ8qmpmlzV96mbFwodgJXKyFgAjw9obIvXTyyTqCSSIwlgEeQ
5/vJHvayAvvlYZXHGHIM9FGxp9tK7JVv/N54UydJ9UZr+um+2peGAUQ7r36WddZq
teaIQZjrO9zM195/6kfkDCQC3BIYZg21cqNXywZP0K2W9qLpnmdTfMrYusvP0H3H
YSEp2KSojKY3WfQoqnzsoMknlfFdsYUIw1VOEaoe1mgrVlZPdRmG2WrDC7N90Dz5
4tQ0kaha382IDSobnTGX7RQMo3ekg9Y6ScW2JYeBOIBJjIjp5kcB0/7f9dRPNZ16
5OY/romW9caeOK18bPFAB9N7L4uC6i+ADgPPwOepnjUhnS14MsT7jhnjswHFFNpq
2Oq7brCuqdifpzSwHjmTihnrqRUFkzeCLKiClcQyIQoMjvi8O80/eSN/2aoNAAka
0tNp9tzvcUee6+Z1OC/0D997bMnH/iJPMSZsKzl3O7KTTNtoXYzyGxv/RT7GhhkJ
UgluCj7PUPiUXpzRbue7wCC5vEpQtc6DbGrRETk1LhcKC8YQRSsjMGrTbbR+SJI5
L17VeumSxJiJtAIQi7tphc99gKJnYAZmhgi128CPOfaxfjX4PpL2Xq2LZQL1i/5n
pjigLSb8F/xft1Y44tsvnXcHyhQhjqD8TL+VlzfkNeJ0bE8NDkmrdLvK+Kd6g3wS
bUueodoZDl6HLcRU2iL1AWA43ZD7vKI/H7YUziag42HTuv/71P6zMN29cHo34h0g
ektnGsmNeIOZDhii0dDLEfUDbXjWloarT8yrYEjWcPCTJIhehlBSzFgpV0rahDaS
S+LFL8rNH+2AW1w37NFugESASCgrQy9QzX1ed1qgOiPvpk3FeFW812Ycoxn35qdz
+AMNykT7ysOewPQQTh5mK/4DOmLBJ18rAs8/Iw5J9KWtTWbZOZf9bxw7a2OAXJCK
R3Es1nC6d/nTT/4J0g2GPuSCMYvK5ZhlNbGLyNhv0CH8nFojg+sudMzcRLJ2NtYY
vseiuaPOVjOHjdQ/y5a7+wRwEVMHkG4yJEwL/9YpeP7b8pgPKU5ycdJYotxW8G2l
gP17Cwra1B7SxQbH5Qe0Jg77np4mVlkRNnCwb8HevrglekX4C5URrqRbVxDiaoFT
isYeJdlZWZxKTt1qSLwLxLQC0ROt5Y7Be7FKal2KvIgxAMHk614jiRGSnoJTjD/3
Z+sUDNmAExVhUksRqP3MCmeyLZm4Jd+ic6YnkVwJH1YcOLnm3SzbS/NWUSo35kxU
aTOU1NmQy/+dFARFOdaY/HmodlBQj61mfuR0Vo7ZqNTqIpyoGK3er1Dp8pgdpriU
FaxM4/RCEsB87TJWbE7Fpz4rthN1ma0gMIv9dopOjJkv+V5oqLqzN849Ny+XDHZF
3yvOgIIDOOdo4P9xz+/PS3dywtI/EDymAQTOWwav0qcaMqQrhUsNEM9vKxkAUxfB
/vVIeKqsDohOGjhhdBAuMKx4jMDjQSVZM8aohVIOmaaPVsmGi/tzXpGEtEuM+6uD
66AUTww2r5LMUiFuyvZpzstRStcLNEbyrYSngT6AAX3XOiNd65d76Vg40xgAZqfw
cfm1H3wMBAV6025omKYndbnc/mgff8xPPHWWUQJPY1I5BxXIsKm351zIfbo3o8ky
wnv8OhNxEpiyEeL1205yQtKOLsnOo7GBIBb2OlDAvmZOzRJkGRebvrVhg3Mdp0lB
mqsMXQMTuDeIZmis2527he+GevVCOjNJLreUi1i9OfUXDk+Ugvs5qi/o1U/uVBLk
o1GbBe9KZSAhj8iKUerD6SlFLYA4hn57svQRSJnNRUcBdSXc5Nzb+Suk/Chyco0R
Q/1GglPI9EnCCBVqIYA4eiuaRkJpsMACdXjfD8QXS58VzwS1iWKpOdB2eJPkaUCt
+07iIRX5Y1d5y8T88TDORUhV53TTTFjCED9XtDGmWkPt0TCKyRXPWWnmSXBkYMon
DkVHtzp+i49WyPxWSWdP5gWreRTO7Hzhiq7VFC/k7H3oVt4/H4P0oK4rifu+XUG3
SubeOQT2fHv+C/xOtQJZmHWHGJoD8Dq6rHhZh6IPavIXvNKERifdml3HEqzs3Y7V
jNc3IG6gIQdeWLho5dnksUkThPX4SNQEDFKmN/gWQZDwl6pvSgjgLrdmsVFIZR5/
MBwcoRrGK4sJwVFjAC9KheGwUjMH4hB4qwFtipkIcJGPCjus3g8PWSGd8DaSPaV6
Hidm7zEjyDwH+BNq7mRdMxPgjmBZLMBEolo3ljTINk5FsN0WO32OkUghfzp0tCsK
zbdMCrY96Oh5y8sY3wVuKxHUZcWy/+0AW54udCOQBhJSnp6h6lcOgeB6LjufVnhn
sAhZadkfvpOn42nam75683HlW/YOb+a8/EnE8sIfdDEMOUF2TQX8RvXqvvvewEnV
CHzgbmh9WIa3dKJGj+HUdeZ/Lz7Q9rsgPxrtM/8gS/XTOWU7eYkFgyFJ2RewJ0Ey
oA/vXfJxSd0kUd4KX4d/RAzWfdf8A/Y2hMbIPhcpnMkrSfSnZZ6S615kT2gXNBBY
a7VWHANnuMMztBkzgYWHZTtjJmSKzeUq7H7wIONeHNMSHjPO8LHLxVwlB+BXo0jQ
sXq8rtpszGmhvXKGt3tX+7Bzfjn86VHHEKsKGX9Z5v48PfazyqnOtBB7ZIX1ecy8
bgQ2QY+ySkXpBdLcprPzFgAz1S8EBa2vXFPCwMzqk0gkonvYOWauIYmg2Nn7KGWj
C4zlv4k+LQKSeuUJ1yZQbC3T/A0OzGkKYOqXszgToPkt+9+opQH1ZEtZ64rdDP8g
PPgEySh3STDVQhK2GCYibFRhsS5cCujplsBUpb2DHqlUkgr3ZkyqB7kKUMh8k+TJ
+pyyFb7mzVsmTfKNYgZA6jOI6IORlADQjOXaJNrZUQoZnd+UV+yttThLxTEzHjz4
pXT8UXEPL5Osq8zA3ptxxHC7L4/mqPq/Dsj96SuKUbLGHECSUIlWgZGt9GHHTDJx
9fBcMhXNmsWy5+wK6gTLVcxWNW/fYhcvDWdFyOvoGJWmrqSWYIZL3RwqSsVnFvss
gVwReumCxNiS9xq7dpAHvn9VVsUfpz3ci3Y0g0s76c5Ta9hdpxarrurNwZyeg0t+
NdUHmE1LP1/C2ABI0RwJAYNNB564NYD6WuS+1UiShSPlhanJE3ns/g3oN3z5pKLf
vkz1D0Y+uiwvoIS8m1fLHuZ5lWDURg5zackLy3WcZqfhY+eAnBuY4BLW/nKBOPyX
W6Eu78UgBS0MGObm/9yj1d/AnRaNP32iwqkvNL2YJi1J+v48ye27JG+OR951qcy6
Se/ON30paK2Pl4+DnvEjooKdyFtgUoCDPEqySkhUFd6ALuPs9l+bWc+Y4tUH4n/T
I7dXVfPmbPhKNlhhKm4yPDqNnwCva5aVEzRv2odlkDbvd0ACcopXCJfyxtA1iHOh
bS8Jd1VegRDrwe18B/0iolYumUfXcurSBRYqLEq62kb7LSl3rJ9tkwG8Il2Q6Qm5
ZtBVTOC+ML8gOBwMmkKuU4eaOib2L0hMO+3fVsb1LLaGDJsVJBBeDcal9xAZiIrX
VCwu+Fek/kWvjW4v1z3vrDhY8jbO3kBLcZBPaUEAvc1vT/L1BSOcwI7YHkowt/jQ
8cXCEgPRgrs+i1yE+xtHIP3TwPjx4YP/xEnjLBEHSVeU9KbaeA8LO85LsWhpdtEc
GVVxM3NsSP5uHdoUAdZI34mTZqkV74LrYtg1lw3rOFRydOcjifTho08aNMr+xYyC
iYbvfQl/qc+6M/h0VflUAvYEj0mQPTUqfSVD3izDcgcFr9LM0/EPd/3iJIVHiDzA
uBiPwRPGV7ZKZqucI28+Y5vvhkqiHxP/qs/1Wo5kl4NWnp9Px3gI9U5SKEtZYiT7
onoJ1TFP+wRrs2NGJPv+b3HbZQqVuSgnWQk3o2au8W5axXJ9RyOVRacOQLgqg3N0
NWlh7vyf0j2PwaTrYX4I+M/fCZ54duyVRtOplV0Kl8Wl8FtNG+lFuJbtr3RGrtap
p99Io7T/Vw0S86+EmHDUi0rcProqY3mshOwRTQ4Zkma+L7kPEv418d6UHZdK0gWg
lb+7ria0IoBho0fhNTgtJVgGvyaw+2fXA5IY4ZkI+cHwUtAggltPML8pymkIhSVg
E6nK/1huK7K6otaUg8vZYbxZ8bhOgQ1bIsYetnc38M0IWs7rVLBNRJgkUFkIGw3R
5sIdEIlWtJAmtX6GyfQjZFVSoO5dzKJ3qw1eZ/YPRsgZD9wW8aKCkaMgYYTsJxb0
4sbK7TIrOMTNLP5+bP7Pd2QgcTGLXnKX7/680c7QdPWlOV6mtcd4leGKDiqasgOU
ry8K6WM1pA0+lNqj5e7kslXdqf3RCGizSsdg/yB9iOuASz5Z9PVQXqdra7AQXI/i
10nGz+aoqaWBBp4Kdvb4ORFOjeJuRIqezAa/uUl5hrYfrMiZE/UFiCIdaegcF1BF
6sW7ECIDrjWcu8RrMh+qFnL+Ap9TT4I3RXtpyEsHLpN7bCV9xhkDSzTMSIqZ+oyB
hKFOLrmhaj9H/VLpM3sOLnELK/jgSZLMXi1YTOSm8XHDhg4+9vwtrtC+eOInfnb4
WsIAGUmpqiD4H2q3dcILaNQ17qrgWhUtRdFfjdiEbPdkFWC/ASB4eRzM9eB+FNyz
tptiVgossC4B8cIiqOtW7eI82OTRMyedz0AQdZxGArQqtpGQzCvRAHFM8N9pvIvS
VSt27sQ/bEEwci9yAo6VNddUEr50TgZ/qPPs0B5wmWPsOC/taJLLLSGpYS4tmh+H
Bej/uvWs4EJ075c5CALO6xj77+T/635+bao0YtL0Di0MzwDyLyw/OZOskS+s/ZRH
IDA24ynrbBW+/gl7BKbK39KCKAzdPY5VlFGiDmJy2EyGUsphQRCq21GbAIxAiRKF
s3VBl4xns5QkKaORVR1JLnFa2OPDyuttlDLI5JyPOgzxGL2AlPEWPExqb+bXqp8d
2ava1v10aNeO5f5BpRTYtnx5FDK7GY1C8LbDie8wbOEYmluiylBNCyYEGlZWFYdU
skj7Z022iGvqkPYpHO9TuFxzaZlESdNi3YrNp+28v1wipRa6J7/JrPVWo9V4nElT
2wYEUbu6qtXxra946xYbE9eRCT4IePH45P2NjDTL0jkusa736MrtoqTbrSg3KkEU
TT//XmmvRTEdM+/mDRXC+hrwCThUnICansNy93Oex9mP6hIy63DhFgR2VQG8mhTi
I3mmNN+2t4u3DP0pVXlRLvGjKiRS7q1q8PxwoNisUvzAE8kgKf0XcvA7JxfAXTxw
+aCS7F3SXZde799dqK+sjDEDByDrwGgrSzqHmpI6O4fuvWOb/+epGZtZXyknuoaE
CT042hnZONWNr7wYYbqNUmo35WRwQWmEnoyQ1O9BlWBF9ATFOwprG7viBknbrVlo
x+y+c8+YxbeHPdvab6AQ/D60VgZkVjH6kC7VyJnjc43/PwIw8xVChMfaKY69T1+v
G3/90dmqw5FZT4lcBznt7SrlucTSrMnf1ttKqFOE5x8tyLMvSmN6eho5TbxCNx2L
PxFw5gE0PkOJOMzPOT8S9i/xWW0HSiucpDNtFtH0EhbCazUOW+UGRhfOfNaWuUvy
aw3VMbCKt3xqyQZ1BUexot+ISJTCrBqQcq8PkMlGgPwibWqfCcdA1dvp20rV2a8g
gpAEF8KQv6JH+VNatB72iBiZlfFDfLlABvUQOG6ELGrzKU8y/fA27m2tZe6/KD3x
nsiuUBTwEbSOPrBjHYzzkKw9rwa+rpzVDgcQS9Apv+xKYfMyI0T9TooKE8AgKXvD
Hx4u6gMHw/JGSrbOS9CNeinxxH74TfVnYRuqLDK7JV1Ej88EK35Kxvok0UWvWyVZ
6XRE9RZte06uj2wlM0Alo7Qchk0N6+fT28+bIgi1jyEvlBh3uOOWETNILybmt0UY
WsR1RrM7LW2zHrTIEdMvg4bZZf0OAhKZWU58P4QBKUoovxnLFILx6kcL2yX/YxZC
n9L5D3nGhYc0J2d7F37Zi1pc1s5/eXMpRloZ/hMufNeDPXz0Shs6fobEJVmWJFOI
QklY75jTIIDyIemjC/cVGQEFk0mMtwUzMDXJqU0zCnlPpEMpFWrO7lQBkqhpZXsj
p7XpSQ9LbrT4V8qYuppHt3D9Gas7RKgsscTlpohSV4Zi1mB1Z6AkTaLrSLVPcRdV
yYrE5tUrqyvOOQKdhGwy1W+G7jB4HfpJVHqOI0bVIpbimBzp0ZPM8wCAJaqe1PIY
9O1TcIhP6kTcsdzTouLikDeOFYMCH6L3hLr7gx7V/ALT65tA3ntobAG4OvYSaSQk
einFXkh8mogy2yAhhAPgAyhjVDlBDMqzeOYd2wpWO3TvY11sm6eZU3VFIS4nadav
HpR0jE1d5tYLuqhDGhADaKXKAyXREHgbipmED3Uolw+xrpdq7Hun1Z/IsLpXp5tX
3Z2MDpvLeuuwANCKBz1E4GJQ0eHPSnvaaB6IW6DNNOvH3Es+lrnqqYnh5eJiigWD
vEbGjdalgtnwZq+KliU2oKinlITmitK11sDsLn1cntHgjECiFHqNoaLcMHBHPoky
4G5MvexgwzvnZ4hFiDVUcjQVlw4+6ybFglDTNNE4B/rohdixPnkrnSipdyWXubLh
SJxi7i3hrEzKt2zDpXAzNZY22/VPkZ7c9mpAqeCmM9ILLgL+6id3GQg0XeLqW7DE
Laz6RgmhSh2CY6Lzc/NHhV9EqWZ/QoWyrkrs8OZgkhf9TvRum0dwmmEpbiDAMyU0
kYvqBSVFUCn0SMvZMCbhIxvQjguzXE1W+OwiUboB6fvznvJFnTVZui7yYFhM3rtM
W1BauoA6l6H11DVPhsP+k1PMSHmBvPSTPgjUrRnK8jBnkcq/Ni863gwwDXF8dk75
ODGsWANDfDdxplY2ilDrNgrwm6uocBEgPkyU3oBOc0TEIBfbSjrbVw/gcXb0sMSd
57llfckeDtFwafvgRPhowBCAxFBKfTq5wT3jdYG6I6pIgaduV+81SppG5wzhYGp5
REUViLUFUWOd9q8K5fqsi8C8zyv12+cHdK/LzlrtzSkv0twHOL6szAHigGf/PeIP
lj2JuxKsEhGIq5vjZ43I+Ikf49C3fvixsKlXGYWBbPc9+7wNHGEKxG8dEDSYihiG
KGxJJMdOEnUPX7GnKy1RDIbI15TfA/RP8RJaOXl5iCST30gtb1zWsASBLPVoP9R0
7XiErRntOhlD47vG4LCVvjS3lxd7GByd/p/xtVzS038ZlcNdjhbnxJzy+yhP6bZO
63CmEeKp0COZbr8VlN0/FmlUtGd2vjJtLfGXQX05K9qx5FbD0lt5NSrkPBbSppOK
JehekJhQp4CSGAYwKqKiiSphDit2ZEUJ9AcVOecgBW12v8RZzgMPtelZuHxGf59U
gHNaUXbdbFEeOMdZmXpssSd+ht6Cag1apJ/PZZitXI0BwJEYtvL8HDpH/zds4qxw
4q+XEpaQatiFzMQvxa0njOOMfmc6thZGaHpmJDAXsO5ahTz0GpRD7JPRd+BUJbG2
/NgFk2K7ls0Q4qq76gyANAlKVzgA3ADAh0cmMTPfALc5eDabhPSeSCShQpRlH9GT
cetf07raD+B9rU5fAPjyLblAV2dr0ts6z4hHWv5DX7UblAQH2CFnrysF+RHGLmmb
SR3H/fRDJmPMpC/Pdt1BjxPVfirIqcacEAjeoBB8pkwBYhzhmbvwjoKInmGQ177e
fMUE6oayNLiHH28nt8Fb4+VFy29teMXSgP2qHTMF6IfiU5eMP8HcnAT0hObjW/b/
36Y/m7R5agp4RAtV4uOKztqiNJRwk52CErVtflg23eAd+DF514seqpujRgA4VjnX
vkMK7NL6n9AS03MqUWF6jb2dwBBN/U7y9TprJ1iA8yO8MM8yKAWjF85q9c/2ZPDJ
MhSJPxv/Pnd1uLKHGKhI+FIuE8fBr/9j8CI8k0aatj5Tcc7XXQz1IyYMBU2pB9tB
VPmXGXYd+/VCQEtx8AGA8SUVj/2MBRd9FU0dtB/mwwnRxVk+BwrHJHpFH7aiTijX
ZfEGwbbB5SqfOaMHGQ6xPzbcgJXd1tgbZ+Mwt7R/qmQVvr/DuflfuWYBy3NCMpm5
hhngBYJXdTAanTyy+OaAb6Z/dIULODkT5b4fA3phocP8bUZHeROuBezz2+tekMz4
ysvvz0Ok4VZ11GqRbKaiUL4BaDt7x9PvHfnDZanLgfldTMcBt+gh0S/1exlDMuIR
qeRfOlwb6GfqLKzy/j8Q/VFm4OSgDJq+9KltreIqmb5WR9mpfbMFPC2Ii1j7UhRg
gvis9izGlinE1ojhJov1Sjso+N3HIRh/hjy+FzcD9pq6Q7yEu5xoNV12q2bFX6Gx
JTG1300blUf4rK545IdOlKqB/3zBzzYnmshVYbo6C5cHpKs7tHCf9/bw8msQbErN
b4ub2nRWP5Qz2WZ7hc8kgjdnnP88lZwcUAc/DRC0dNjE2qnj+nx/g1jA8LsZ2frZ
x324Y1D7r1wQSXiysy3L8wobNnQB95+tvb/1xFanA3Mp+ayJhGdrRMpINpBsSA9i
OrHNbv3fH7MVNE6WGrJPYXyvxNc2mPnO6bA5qQsJ6aMyD3I/uP5U9rSYo0iNX9VC
hmito8t3AUHSgLGnIx7EQqdVeGIbLyUb8693m55WFd0c8iE7aT82mb8slPtQ7TY2
fMpuO6jZFy6Vh0baxaymy5KYLchamZSYMNPtEQ7dqLIRUdGn5aB80XxPnuplublA
ZEPZXsxsLStjcz/5RluXP3fRWVkQY+8BCur8DNoKEQGeCSlJFtXa72i4NoBZzJEH
3dEvBqfaXeNj+mRqKlNjkN9NK9XxvXSonxzDQ1v3Qy7zzFLCTUFVOBqlA8w+v1/q
oVTqXbJ5nTPS64va5RWn35ysB5NFUvWzDY2NOpCMnEQRnCzIx3cVyf+n0iO8lld3
ULONVnMCyWI41Jm8R7vkC9xGPB4scXmVP3yp4Yw7paUTikG3hgWT8RsWWcZOlJyu
o2uGcsDE6l2ws1B6Ax74nX6rR9r/2RMpTp+DPCZ9e7Gt7MViBGsufhzfOPp2S4Fb
ndnU2NQP4vTkJk9t2ZHs6wBHV4pIkYjGpw17TtzRWx64UaUQHXY9roO+7cZu3HYS
VHMbIxnr4q5zVIB8wW5lwNLuoIGIqjT0FAIfhYPh9JPVuNTFb+ekjpRlPLr8ancT
QmqN4huFnliOhzw+D97Vm+4e06VMyMPXOhF+qz5yulxeV1D76SdCvDEBoWZuUsx+
QtejB/6r1YA6Xq8levlXIAmyRBu48F+WH6MbPyZObEuOg7Rg2MSsKKRJFdWgmHKJ
LSD+aoC96Smxr1zO+3Cs0unOyv1oOJNatAhVDy7EklNZEiJV5nt0pOR0bJ9SaiTu
y0pxm8FB+WsGSv5U+nVlYSKarbUAcBEUtMaGNgW9UoAXp0GsItijelJpTnyRo4kg
L447O1QwKp7WFqh73pLyZ3+FpOe5bIvzJFxQ1mcnrU0cpnnk8qF1IzC9/888JUbD
aEZOHUhEjHfJHNtxbR6Zw4gDfspe+CpdEg6BYLje8lBZgyqt2HB3tZrogjIidbxp
d/VFC+G+oNTtqBDpLGtOa7Z6YGYrVgohMCY7X1m3smaHInUIUrteggak660mh0E3
Fpwzv8QVKe0d+Ntg3GlhiTHK2pNhOqkceXWaIN50SD38L+KecHzFIeea4VRmGTuT
PmL7K2LN+Jm111IvNIxkKlX/XYYshZy3aZeOobJAb+gaEOOyC3T+lxRbViIURyoF
FKPwEzuIBAfY8aDbxSovgMLqdRyJrLdyYGOuz+vqhV6eLdU3Idx7cNHsUzmaMhd5
o+cgbYa1USNPWbcPmnfFfzW3hTgr5oq9OIU2gVvOdbyOuIubJmUndAAvuE58dFUc
Uqa5aOUBcr7dxL5bYenxW0O+KbdWP1x7zY+G9AD+tugIrzI9kgDipweKdwKLeeE6
rr5pw0jwYVR/I6k3WMG2A9GBdIv80QAqqEf9ar/bUcdlUeohqp2yor5haQpsU7Bp
NOLEJxnKyA2Rz4KcQL68Qjge8nm1PwN9pMIsV/ef85EDz+0I3gBME9xrGLGrQn5t
uAgEXpnO8at7XpJVaYDj/oROe8VUrsWMurJe/+CvrvuFZGiDTgOfO2/LoLRtPqPv
E7PEqmWvflRvJXJ94gbJb9dSgLDMQfOi7/a5TCLjizQ3rrG4vQiHKmNZe57eNjhf
IUJHyUR+G9eqQGZSUQyhtvrKRY8KBJuTPt+jRGicx2S8SLX26DRMH0TDEXMX3vli
z/OzA46wTmtTmoqTdlLv58mqyq1qzjIKFi7eJYDx9Vm0ebaaAZ2wVdIHbW1yYvGu
93LZjozN+CQNfbnEKQtB8wYN2aUPcblAgXH7lMcLyHKlJ3IKc9qhHTulcAONuPDF
936mGIBWGDDTZ0d+hl0dImKsNZdT8Vd1RxFXeuutRhP9B7wDe8Kj0E1waXQy0XFv
X6iBrWZ8tw4oP/im7inA0r8zGVmbt9ZlF5+qgpMfpV9etUwIgeVYzE5ERtkH/+52
yynqC2yda1/1zQQXznKfw8Oefn8rKEXbIx69Q7t9FsjHpUgGK/HSj3S/QvLPlyDi
sbPaohpHZJa91VkUO303DZpaNajD8KwYiw5uGqPvS2yBJSmXDYfkd0N0ah4PJQeK
H67wZZjzj+stYO2dXMiO9sfHFnob6RFmNFhue7S2Nq7eY2cyJkAuTzvJFuorWLG0
2fImuXrp+wXK2Pqfb2d43YJr3/h0Q5n6AwVGkHhlrjxMA0G+02biEnnypqupgqke
jsyOrRM39NXdTHgp4/ShuKJpStnEoMDbO9hs59HRXwFd/YDpIkMY/c+D35BYq3J2
mYfljQGcWCrFn806GlJnRJhSoxe94Ky/koZDoYvXEhiz/Q8KyzhArHIGnRfcUSAG
M7OWKbiA7JdyxDlAsw2n0HaWt/DcZynAxQdh6MB7zmr3PZY31DO70R0czMElMNua
Jeb6xLrMMHwLDGyq6t0bCAX2vkJWzudSWulSNCoMplenm/sgN5RFXU2i6bRVeBHk
VqW+jt4rrnDhFEQ8j1zYWQ4UszNHVMjHPllP7Sc5jWoWMsLyzQUptISx0vLxgblp
zz6iMcIVVftegllk8BdL8DJd1jUCgf7qWBQQzekL0h1qVBfqkRC92OZAHqKDXhll
UN4M8SWDSOvCpHymussxqobCsTgWQpnm8H0dXfPCYPqUwVIgVuwGdgSfj7JYNMPS
YTadvzITWExL646GvORxZGXxPCGt5leqPzyYpSOoUeRDDUeZbWqjffJ/YWNwqlh8
02JcIfcV2t3fTW1F+AHhFuqYkiW+cZhkpiX0V05+JPvNQcaEQkjeDHf89jea5Ubg
2MpR1lhLE5zTkU0ibqy0TU0bxdIuGzChf9veWEpCgf+DtTq701bxGfISvi2SlFvO
04IvUL5bF2p5gmy7a0fP9pCQHLWX6W52XuPJxmC+4hVjCazlQYrtENLVRgoNdske
ynokTs9lHPnhBvR5PPhRxRj5pXqTfvoIW6XtobviAxDJips0LWodZ00BsDVt34k2
FkSw4bah2XMABswbTUKgXuwkG8Q016Jpc9xVIQXxW2w8baamwWPSagnuQrBUw30P
pWsIPGjJbvYdG2azaAYW47cO9/4qN+f18NHmvU/mA33xStxhRlN+HeeP5/l2Y3IL
0hgyCiVl4knIo5BZtUDFJs0IIp478da1mMCyCdczJHiV8SXER5rYycqJy0Vh/WuX
vxNN1S8xFe2V8Ei6/jOhQ5rA7PeXum47jQOF8ubgzN+exCR7i6fCckn4v7rSILKp
akaVUyV5YBoqbY29RbIoKk2QfUWrXLZZV2lCNQauTHezPMQYVDFIx1lojUTfYhy7
oYjwQiDEOh6ubJpEu3kZ3HlVv8ZJCByug8BkA7VMxrzjCm/CyxT8SMfD6Uei53d7
Kt8kdPVKXoJvy0NRotSpnx0zmcd9SnBIY0t00Yl7Z0RsK5x+kwiPz4ROJFMHhywe
BCv86lsWKwJmCuWOQ1HgtDmQAhXTlLLfQ7cx3B70CBDfmmp3oLbTK4TmxLo+09Ra
NJ0GAi9LARlJ1A96C2jv/dzJrBtUJ8Y5XI3N4oYZZyQ9kVyEwiitdZGJKYfE+KF/
41PqlKaYQHZOL7Bs3ved00V/IqMJpgUIvFyjTwpmOiw7Myj6uycACRVwNP97bPpN
aBeGauX2VhsT351a6jO32eswLerO9BE/gZq4jqyCMRB1ielAC3g0j+aHjtiavcTi
7tZuCiIhgG/4DoQz5c5IEJS6TW6ZbwoBnb5Uy7lJ/h1zkjZVN9O8Nw8SHEFhWgoX
3PPPI+8prvPByOXle4OACCR2eEpEL2Nni3rapEupgMJi42BUT9G1F4CanY+Kr8II
GahSmiBiwOKJdvxOWo0glCUJO2O8FtGcx9Rc4AuAtoNX/0VNmiBZTTX4tE98piyv
F+8czQkFe/RiuN13zXnc/7bPSyVoZxU0XEbgqWkATVMgm76S1DYyzHfqz0ii+rFX
20xTaCQn2f2JQTfWuwQnBPB6z4YryHeZYMkgX22fNn4Sz6KpHFBK/DgcezI/36bA
k7Ju3Ft68BKNMVRu4YLBCsC+hgqQLbzfTF8+QhQIX0YJJjDC9vcYxtKcH/E7pURH
Pveaj8balXLney/sTTaWIra3ZI986QTyUaxoGBt31/6LMqnlBwFWjbu3phWGkaKy
8EmK3Qdb5zKBoL01E6kRX5Zf2Y6kWR2j/infYvCzQj8ENfeU2GeELtjL/xpEefF+
J5f1u+7PHpCV+ZgtFLNdCA7Hzw3wtNUqnQw9YVYQ1QDnDEqOB0KvvrG+5ZWWfoQv
1rgiuCMqdEIli/ojgTChbRl4sJYwoc4Qhb9ELw/TpCpgrhXE6NsOnFLnfy9tSUfR
RTM72Pwt9TzXppXGEYo56jAZD4aQTSnPXdnMuWm8i4UvRh/IzdKR3RsyACo1baAK
eMkqvQtHDNLgo4YrYKjZTJy+iheWWRC96iwIRWrEU3NhrgJsbAKj4unXX+CKAf1e
HtTQL4liq2hOAxOx2mPmTMzeNxBH465RwuW6EbbmIW3Men31flaKSmgKZHbY6mn8
OdolKkX2TsWDUpDz0pI4bqi+HyFjd48VfALthy7A/vDU3lmbzYfyCaTe8i7VpTy3
/PiU6W9jCOPE0t3lkTmamP9gSRvAaEMQ2AVAKrIGWvLMBtL7NcRV7OFU3GgjbZvJ
ocxmy8hrE44O0LrvS6mN+GL7KJm+erfiaHEbROKtCWMGL5hZjEwhBSOtgvleJ6L5
zIkKybxkxamtoj6TsC7MOp58C1m18v6kbbk985TT4iKxBRrFgWcpVzTJ6AyrAeL9
6Q99g5wXfEABaWAnNp6UeefQSGf3iS5BPFNmqVukmxy6NJdGnbNXd9ivBNRGGd9N
LAPxqDB4OPn27ComUydY9yKK0yVj+ZMsroBX9n6T2K84Uu1S6Jy4/ZpGIr+9Uljp
O1I26UYbWfuS8BRcX06s/3idY6FbCbADZs1o2ZyjmE8pPUtN01mwhmfRNuw/zTIf
IOwNxXj+GeRKWpLNBBVB0AZSNbfo6AThBwjAPWtcxWGOWIN7AuhFbNQq4vY/pu8E
K7Pphl7+b3rlzkQOeXFp9EWllMKJmc9ZViLQrfWooOElkPT3Zj44FjG92qYjEWVF
SIZOHXXJhIVAwXKoiySVuoeo/qO59GiW+AM6b52HpHggXVvrFm7FSpjMUaMcN9pY
3h5ylDCUim/kmGdzPljBfQfY8EECG/55GfwsaSV5j7NBjifSW1gsJgEhpdAkk5gx
8nGIoEi0i8jY83Y4paU3nhyX0dOMN+g3jLGgNZnpQ1n0wXKS8m6ZXSjKTMqdf5Ka
XYGGIBseNDIcBEoxymlhVOW3BHBfg+0PGgKE2maJIIcFyWlQmHF3K8N3mE0inpL2
VXCk66Sl55DbPLVgsPoCnZKYAfGFLOf+3W41/AjtUxHC/JMPjsQfy2HeOKF9xXGq
25+vqeu3FYfqEibyoV+9t5Uyg6DsmwVxTDPjdFjHGe8plR8k4hPulBtQn0vvdLmU
BU86C3OxbrrhwiitaArgopqoXP6TJu2MQalWSFcOC6vORawl19E35xzhNN0wFwYc
xQsCUiC4L51KyXAUhPIJMUaCy3XSXE8PWR+UMfQ4/cGoXqhjWq+5j0/mER1YHQXJ
hzdBIgcK3S3RD8nB3UHrdCHQwI/x96saICCYio2BJv/7ZL3eWME7nFeHbbQ6n02L
QDnU8jZ2XM0NNWtCUE8lHzm+bmDd0wvGesuPG2/XXHxlyQvtwwXvAHRXsNkHSgd+
yk3bfzgc48LHSmqZucHYsgMEQMSCBNSZMqSSait7ufAHsLiGkvdNF00tObhcrBer
jpPIHIu9EFyaJpTzzVvMXgf6/pOxLomIZRD4jOXleTrkDxWIGWH1KAcVdulxRzUi
df4NmH+LYvpuDEVDSZKoaRdwUeKKykjD4LhRAc0/y/XNV3DYRNGw5dqtKwHPbPjC
0YTSuvcjXJhJCj4cIJdmRbzdHHV/NdEMjjeeqDx8aVrR6ssK1FbcEQR+UjgcmEI6
uYzC1w++lmYOS4mfiRxse4SUkNF8Tg+ncVNBq1XnWdET4CF8in1hwTll3cEbV8dw
LbdbqbWB0L5S7NNgE4qBJzlCUyiye1SkJk12eVIoiUDq3VFVnMQM5pNNgHADRfrd
7+mG+zF9bBfrSBALWBdA9h2udZ6VYZYLIlPx37sArMdFsZUdAq42rRgsQHi1lS+y
RvOxcDpOQY70Zn2yHweyYPg8IuJ3j4tV0X6BefRRpOMhoaeehRLZwGYRxWz85rlX
EgMmMsjkFIGQ07zIGwKi7yZektjfXF0zRsozRxifT2fagF7Yn0CqYQf8KEGoq0Gu
GaWT2Mq1GQZSn/HpUtxjRSaD4yryNOcifO4oyoBSrdVmptOiDuJnFyKflECmPyri
Xs75VgzsKU+FEznugUFSnbn077RabBt7hf6bCriTHdQA20JC89ek+VKWEb0tW4zB
NlUfCdcPXXh23r+uWDD5OGym/BZXsjE6G/4OkC+frHtr5xflBLh3B1SsaHttnxbC
SlBlaAhzLzWZEr0IGGJKktf7KsCYTSyYIOMOddfktSUlpsuMl6c+k7s/tVsL2uIk
olAmkNpwxWsOrGwoHdS3w/kfh52VMHc5cBVU3Z9CGfeHwk53TkctCkxQ26WxFqnz
lfVVtr1EDfZzVHXt3futtfTP+rEz0QL35kEkp1nkH86lkicKocdpNXYvRUw2v8Yw
ojWMtVqV9Tm9qxc28rMegF/3ZClLluNIavkfHl3vHql1AJJd9yhF+LEeVj2IODw5
pgrvAsnFsLu2254MzkGv0WLpn6rq9dNP35Pm/lcF7GIPxq4XO+G9VbtzzVdrAp25
5i2tWz2knEFb4FRDpeT9tsGrA3qqqfX//yMRn6sPYCKcMnQPlEkMEqxkymuHDrWf
AP6a3JApZFJ7euGVzSLLjLQa9GmO1ckNFyoNnIXcKD4Ab4k7Olnj+qcnySFFXRYR
48ufL58HL1142/BPv9fGuGLmeqeHSOkrrwoWP0fM7uWrMTL6JUSXdRMFyE2Qv4KF
8XCksKpRDLyPB2w3hC8tpgiT+xN6nXsFyeBV21bqTHp7s1ZJ5nboVAD70zUbPGXF
KIOd0lwuk8Tqp7TPnIHZ6M/1Ur4iNMy+5plYd4i1FAR0yruBK6WRjsf80i5qq0GR
R4kYYy3XcChoaMSEbnx3YAGB2q2f4YzzWl4zkTpYK+XN09W+yL9izZxkQ/fNnMuN
UCo8I7nAbk0xFai5h1RxnWumT5bXDswJ9K16K73tPRDTCHqjFl65kllbVyiOV8IN
JJeblwzrsCwLwwymUuKVFPyDtAOMOpTfkOTMuvyr2WMNRlKRDmhXIagPe8E1dPES
aXEBJ8N7KII4LuzLKMCfZtMJVacVLGj40gxg8wvyF9gphWLq7OtZT1Gvs4sYUq7I
ZwMHU/HXRjgd9vmmrT1r6jFkpmFxc6cSzWK5DgU01y8yh7Yde3ifWzABmDTBqPFw
n1MbHRc2n1811myPwxOoZMy+Cbn9X4oPX63vPcoRHfgyUs43oqSgH+rszPC1lrco
8vJ/GnTvypXdacITFI3Vv6Rh9Gvb35E67vtVn6hojRkCnWvm6JmeFLlCZtGZkESC
qSy73fghJJmweYWheY7oeL4tklDcix16CTezV41ysafJnt4LMiG/Z1Xqwfrb5ame
gae+cbDiDpmgCD0/YMaS4B57fx7jwUUysgQxoIzxEox1xBF/VM6j1Sx25TDq3DiU
OqNUBvf/K9Zv/pKNgwWRoxU6lX+nhcW5Bf0fzrlndb4ivdHiTNE/38YPUgzfd9KP
12VzVk9vYbt9WOHY5srxB/joR5vWPu7gQ/J//FISiRwEBf5RZeb10+JjI9t53jb9
/LnwOE0xnZkgWWmx69/4hYpyBeTSkI0O6jqntQCBUpqSbbhqdYLMbbV02I0xR2vR
lUyyZqdWXtk5E66yMMS1YLYH1PYfm6iUzW2XZE43w5xKRYR10605YUGd/e7RVAzu
0MT9OZbewssganRYtaPJkB3bKxIjVqoQHXK0lFA9b54ZqSDcd/2tmFWW2GeZ24H/
Syt8fraCPY5gaWvJTpNx3h4iv7mVMAFH6DXoDsUbIKpQmbWwPwstAucUncb43TeY
Elm04c48XJf/HiQ8IbhLRw5ortgtLdNP0119wgCpiPuWMBi3oMlYna7+f+wrKHtn
S0eImlM3qLg3fQShV2wCC884844P2uDQYp1UIkr3H/E2r2rVvH1H/KmGGRSSBKBr
1cBkUVwsErmf4AokOaklfBY2lZRCdqyPKdncObTay4uZFpBCgcJ19rfDEAJaIGiK
g7Pjwmnnn6AFIhorjHH1X2/+7iDbd/k0EXAcTwCyWGT0iSBEsHjXsKkG8rD5YIEy
zTaOz1Om6d6ABn0ENYuMdfS8etasfj+VLiKSxb1QbttYB7M7R1uD129pM6WH2EOw
PrT8xhg4ymHLdPAt58ks2ohI1gX/o+bqvH9ARx6FmR4WYnXExTD5ecpSdO1ECmme
ER22KwEkjiSH0gPp4fUN/MZhSA5iGvjIyzDQRP/qpci7g42kZIi3diGJB3R1vavL
uEHyTdtQ+jl7q7X62ybIF9u6SzOSQXw+BHtp2mZAqxJpFna03Bk7R9Emm19eXDZ9
9qpXyCoPtJOY4ZZwhOCxBWF2LhHQDH5eOBwV8uR64fMkxUafs28YpUwFf9XNYmjH
UpP9XYR6GT1fR6CMh68Pi+fovhlHu/utaxdZ7DGEYunNBZNCkBHtfLp5KaK3G11Q
LuEAnfuDSyQIbn5Vr2uliklFOsNBfvYZ1s/UV6Kx4gnV5oBc7rNgp3vepxGyhP+m
1RnWpTDlzxuSQd7KgbwJAE4+Kn6LEBeE3xclVs3RH1fqL2ZmLJ2nSbxehBeNUb2O
nbmg9Qw3+/M+tjaHG+eZplguh9KDpAReNS61dBa8f9bH1w5wW7cYHU7H178CWv4M
U0NS8YZ0AW2dmbMo/fRcj10A5n8W8kNez3+vohAXu5vI45sUZcX4Fga0rLxFwuNX
PQoIRFRJJrDTPlK3kI8zW+TR1Z4UMEQ0RJxlxyFK59myZ1iEPr+lccBz/ZjWmTbp
MoyKIgKakpdM2aifgQIQNp0EJeXTwbxqfbvwELcDYptQqlo1bB6ksaUqDjwQgR+k
yoNzqXTUrY92Ef+XvIb7E6YHVCc+g39Nutqw1YoubTPfYfHmCiWsYAZQ6kgV96jZ
kukabILdG86+lns3GV5L87/ZkGOmVs3/LciPr5mWjsI6YVsI3MTLal12n7Rxa0sn
JeB//YqBzxGm4QkAX/AgFVWzLx2qeU8+vycyHcShJ3bN0vJCN+km+jfPe/Sm8Ico
XapLX/3z6bkhbZkR6l6eY/pL/pwsZAPmDUewJihvwNxRZrtcQzNO+l918PnwgH4X
DOCV8aABdW2jaDYwwa1bM0Co7NgjrwNLZicqcXRHIUpWc7owiIWB65OxaKIOjkJ5
enCBe9h4u48Bp/y7PHC+SZwyYGfpuA8O3W2Asole8O43EDs3KjJlj/15kErh2d/D
zf69Ii94fNpU8wamfGiF2oCKERoBcdYZ68jMu96DsrlDYchXmlEMAp7uw/A5tvJt
qA+1MLqCNToC5wC3h6OwtwCXs2n6QhGITevnQBjSEghjqXLwe00lKtYFjs6SKRJR
qkrxrU7S7oWTwxU3oQ0J6r1PMEOlj7pGIikC6+/WwABH/sKSM73BI4Y8Iayd4YsF
H4dTc63q9JR8a6FGhDwrCUUQrqzadWNL32nb8KtQRtREfSg1jQku8HVsCrjupGw8
1iZBf4llq3PchofXl9BqzDUE3+j/dO5PWRQV3ei5RdTHL6DBdvjywOypQJAjkAq6
NIVGfDw3Ux3OUsJo+nRkfvfJLf9xeTKlm3PaTC8Jx5tVagHq8O96TKDojLE+EKIe
zg6vG3kdrr4ZYVQZ8tPc4fDPWg3sBlcrE+yImF3yYnG1uvtvoAVSws2iPgQLWfG3
l8QoIPlkxRIJYEIFlT9cf/FJNvFU6U0ijtEMgDQI5mvxFFyySogrvzaJRcyWXwms
GIzOfPgTb9ehaJR7tKyvvs7ufNdP4fyU4xuVAtxGDt9FDSWcrBC5xI4QGmOmFXiY
bCHfxFqOHLjPCqJ/wXWBJJQ3Fy7GbRYglZwjN0bfgrCymXw36b6YKdJI0Bg4CkgU
EWDwQoKrAl6F6mtqxj1WkoBeFS5GXhD1Rn+FOqAmocLeFk7elBJYtcejh0+yxEgL
Sz/KsJQa8+rLTkDF7+qr/l8wHxn+Vm1AOpGcNH4CoqyiqaIJaRC53cQ0yqkkYZCM
xt5kzYy0q8fcbLedpByqt32WbtJrUQD4rUc1U8gwZe12rDzk0g+YQzIIoFTDD+Oq
Pld2/kqw6C98ba3gQdPk+Bc39zZIakEBNU6geVPvytkKXaBFsiNOum15mVFlC8N/
U0uQwqb+G1eGSAfW0je+Uzh+a7HNl/E9pjp1Cv158L4PLmKtyJRgOPal/gpKsIwx
m+0OgWzl2qvhLSIHua3AfNPj7uG5CDc8+fhHd7h5JGI6dqlu4GzobWapcOqMJGpa
1Ejbr0rDya/8tl3besc1ykwF8gWH3IiVrtUtqy3mwm2oz3qI+P7jNsfEt6Lr0JY7
0inS6mfZN83IOip1Epqatat0KDapVuyOk8KdmSA6oQhh8e1SPFF5elqWLuftbqUh
gXoT+LkFpjj8RSrxfMmQ+GJAS3OCSUeTzmgWiTTmSvRFrhhiUnG+aiefukIi8ZGj
CUtov20wQpQBmm1jn0v69XQdEN5SRkW6RNwCeb+Xi4m9E1QyqjgUL9GHXc10IdAD
4TC0Qev5j1E4xj7TjnALfu4S8uCmut+vRLjl5IdXAw0MwjwEtI+tvipIgvXT/agM
36dZcz0NriBEAJ7+QpXArhZ3J5p+GhkjH46mlVy5p6eZgnFumylE3xJj71DAL3gi
j4FuycagGfXwmkA2IADFE3yczDjbCCG6FqecPM8OJPntsDDhadUcj8AAlTDVXsJb
CcUGhAM1T5851k3FdQRyPofZkMnnknNxKDEGaX9weuiJoyw+iO5C9zR8sO6ZrCmv
VTWaaHc8GSjPPyZ3tj9rwO1yE5aDR5nh12oOU1z+S0j9sveLOC7LMxZ6Z95pyjQM
Dbv719fWC4wKpTiyHIRsg6TLak5KOJzVUSWDHiCvqJHx7diSqTfbLonJLhGrRztV
O4OORX++KLy5NHKTo6fJ8wTVsrEcqlSiCckLClpqU+hwpwq48/QN+5JjY9fu76e3
Hnz451QzYjXa9PbMqtKOy/C/Y6cKsYHbpb4WJCqDnQcHVRSBjhkza4j9h2bmFdYz
cE6k5+A7AQYm7tJurwFNhdbsev3VXdWdfYoHnoJpXoRd8e+yVzL3tcejNBc3HyZj
AsYWLt8BSOvhUQCSVMzzxzVMALKtj4vuSF+KenlRoel7cy+HavAuhc5A6uVD1VaR
9U6Bsh6S7yOGLf2h9SfHLMviOjDQ0mfE99qr2YfvcezymE38aBDEYADj+qgsTe2R
obvieyGWOKHB69Jg+fmoO8hBU3hLg6ixLHRNlevkZXZmLdr4a79xRCDGwnDR5ppl
un+Nz5SVF7rKCMVUXKZzxYTKAHvHTcGM3JY69/yZZb0D8dMvQuaKXyvXlRTdbRzx
lVYP3xdZizNarHWlSdqY/JS+UuwoClIJ4KSmjz2lz6GL9Rk5syTcUtF+LFRrjfUi
zSU1Srjla3zavWaqG6bO506YQHT4oVdxchIMHFPObm92MEGUjnXlEysijCMAtVBe
yLYjc2C6V/x2fjwsSjpfcfrZWQ2w8NkoYwt3uIZx8qUtp18kR2Q53awCyhuHEHkT
t6JRCEpOGHH53VKjslrm2FkN1FzsktbauqC9DttgqUTGM5akFoJ4AXH3GG8QPP/g
C+aNj/R7Q5ifUC+i97foVae5D4Rijqs0quyvcJegKpeIP2QitG/bewkoD5pZvX5F
zk9UkYPrVYguSjQrxcqsdxsgQhO3AUkGnhdSX7SkpT1vIBsGh6d46R4vYwz5vm3j
a8NO36kuTjX/xikgbCwPlzcKVTlyQvn5eHwUkfV9oCuLHorCfJOxeW7/5EjUThUk
I4Z4SGd8C0b6AKgwPP7PT4hro9+lhSeu6ueNw6GkH4AXII8QmWzx8BhcNX4yklNN
ZcCWej4Q4qed+2Db0DQj26a4uNK5cd5yk8OIvgJ6V3vz+uiiwz8xU86Nkws2I4Yx
ipvrn3kGaARXvy0fAHIXfrg60TWBcLaM8mMgGt/beFe/2AoHH4F5q/wjqwLsAl95
o2n+8gIWgFafsloJ/IVO5W+f2i4P0MbOxHZVkq3e/pkmrKyBMAYsZEnY3VCjjh9j
dUexTdDJ8Ilsy2WoOs2tnx1eao1ITy0YaWkAjUQjvjZV9wKjDkalRotFk956/+HI
Gc2tSSyEdwDmkUoHVomzE+ufS0KmgT7RHkIgeG4OBOiK+zAB6boEvZ+y6GPmp+f2
Di2iD0jdYf7EEr8OvEkQ2QY76BUhIKC3/AsIesa4x3eFjnZqziW7wdq5zIvUtIYB
WcQpfEHAexGZ/wV+/mgBfw+wxBZ8oEX2Km3tKFqKbrnq7lK4SkLmQOZs4qVjy8r0
K7lHu/lI9sKTGo8SVwWLYJIw6vzClFNQ+BNESSheB3RC8EVcMvwH9N2yDR19TvGf
JJxRnQCR/0CjDGCk9QZ6Io7ZtCa3OFqKkKLMWJk4k0tn8b7r8G/lxZLvR9D1PmnL
RFR317+mkQO8API72e4eJ5fndEJzW/+jYf7w9y3+UChqOWcSAqO8PymofZp86Nh0
xwwk51a5ueukDxfxLUjc9OLdGrSrbgB11m5JKWyUWNSKP/KgC1Bd6GvaWR8/7qWw
9UEUMaKv9p9yuyeK07Pf5nyNNwcNlVBnTw8RtBmXATM7YEzefjckRfregAFAOk5S
2UBD1kMvy8HgjqLURbiq3fmWJmG85n7YgR0CIbUOU1IckdlTvzDlmkoZddiYPdx6
VJpm4fYgYFduLf9UYNGFm2A1lACtWYA1BIGzP1hMiEu4OZoN76nEE2LGqp70EG3+
IPWnjb5yyKSArvcSPklOK2PTfTScywInKK4ACrb14zek/NdGdM2TDhc/eDNDlX2l
zDErwgQP2Q7LQfX0VRzApVt1ESmIEvL/xaXjZKjeNNQG9NcnYz2HWgBnbsKDOA09
7W0Ot72zJmk+We18N2lQBjJWba0+edbq/VI56FyT2ZeKbCDlHj4lzMIbJeahaEzb
bSTUYJn00AdcuWql8CigRawUPGwHtquiIEX6GXx0UCVsmPR4ft0wR3AL106MFSr4
YLKcD1GohHIl0RazgVBUecMfolAY9IrRYw86ExQwGmx793K4qW68DjpiMyLno4tA
Rb/lILK+EDViitwNa8mJP0iOC05O0LBYszVO8+Fq/LOUsBcgd22OVhiEvryVz0Hu
2mEJoQUsGZQlm/jOhy/hE13orugbQP8wH3XNZo10/Flz3tP2sXC8o/GKA6uErOgK
J2PYugzh5Mxjw9EE3EJKGEriUMcH3rXfSyL095qN6mSh/8aWDa4lRRPj+bGJA60S
KBPrBwuM88tIKt/YbmUv+X5ACZ6gmbrlKZblXuk+C6NmcPPSUyAc23Sq095SrYUR
Jf0+qwz2ISN/LKYaq6Hha49ZHhReWuFea9DY7JNvKVPx0uX+LxXLyLdyOwtaTUD8
cnovsRs8QI5V663IEOp5Rv/dZ+MPkaBBKsi5yQpCVDpmMpUwfoFYuCP+aTlWDevX
WeJDUtxTpOhM2V7kCLFnWocs/Y9Iz/U/g7VnPuESrdHpYYaCmxzeZvrr9jLWNv4i
PQItVZUSLyKFs0do4flpbM+o4aLqaz6SpnJo9ggGE+57RKCDdxmEnyv9KEaLBqvC
IuZfutp4XU3oq4H6UDajg1kmzertCHYXOgoPKD4JJQuZ9WuZOrm2glFf6LLaPFwp
wB8H7pqz1ALcj4xlUappWVqgpvQSeyN2POYQD5aXsY8IvpMb2kGXXJFRbIvWAKuy
+JJOtUOqyh9YpBTIbl/9rNd//vbwnBSBrAlsFl3zSxShJ4o64dzvpRzBDdpeNOA+
YIRziNTpVEUgW21QQunVA0etWbxInDsZOWRdx/FsGUhANMMvQTlpaov6kz/HkUhl
5/VCGV10BTRsanWLYHyOtDK4wJMV9+ha6EB/z0Wgm5/sga+FCvCanYb0+uBvhE7G
S9Bbr+hi9vIUDVNfulFeuWYnGLlo72L0sYUFWgLAlaVj4N94h100h2XUzDDIfiJi
ZKrx/W8YCk0XqZZHXgHrvqcn509kANpGJ/vhlu5w5Y5Xgw8a8LdmffF9CtVb+B/J
gQ5/Q/kSY44D93bcMEFTkbUeAt370dBXptWzjDUKKxyf57sdXbZYIFiKLJ62XZMu
s3W68vwLdnYb5PqpeYwXXqyfjuulXIr/c5+OM7Jt/6IVN0M7nLMQymAPJmOt8kkW
qrll/tm/HqGhMJmDE7Fn1L7bsR+Nb0YE7FdWPzUv+cVztXSo/7V71gKqntVNWuaL
Lt8lfIEQ9SkhbPwIhyFbtmHUKe+/L25EmsrL7tvMgWYces5r8SwYuVFl44A4m0bv
JXcuNZz4uCF5hnl95KpQ7pE3UhuC8LWRnYtJBzc9UxWF2hpaBpjwJsGT1nnKpJZD
uZ9ZX6DCaQVcNa79arBludBoBTRZyVgt+yg3MJkdHaz2f+yL//GPRitOG7CHfwnE
coM17nhyv2QMoroqSn6/ZtoKgTC8ONYnRtJTJF1PPHM//ZzAts2N9m3jt4o8voFW
tQbqms6EZghKrOLCvqM54GjtQmDJGh+YI5p1RTHxwJ0De0vtHS6s3f4x1aqzSTtc
bQeDbDRRB2XYPJtn77xvYI3B2YK+cFIhc7roBT9m9Sgs0+c4FOobKeQl+K4d2iCx
cL2yP6wXjkEX96/F7yIyeMq2AdKJdNPB1U1dho0w8Mwupr4WQ7cBTbwi0oKqXIEM
orEGIQVRP5mmdG80Oa02rD0qUrvLqZLVhUHVsanMQPSxKVAPPp6pidZNK64V3jF8
y4tj9efENr20KZ+gteBEcxM5TTWr0SBZDZtUy0pjp5ehVgdNtNcNiAVLZD98JVX6
WqAe0Tqdaf9J0KmO6ufGxM+uzYOkUBG25vI+kP/VzbvbV+uW5GkAEqxCsqTBzEGf
c1o17Y1VE3pS8gHqv4t6brLABkfbNOw6v40dBRhHlIrQ7Mp+1oCOyoSUBOfRc1HY
tG8v0Qjz5H5domKJz095zCT9C4y5PPfeli5ioSWtqvptqE1RBcm9F4W8E7NgQRPd
jxoJoGkqI0jQ9aB+K6EU7br+v+Kmx0jSdtkay3WpMQG3hh2evDsNXuoXFyZewsy5
RI4wyjg5yl79mxL3ZSioHbc5+UFnP1l+DxsILrKVn7xKBxIRHnac5sQz9IJTkYsq
YF57bbSRkiG5rKKvGMCKl6actLs0tmPthzbVNNpB8Q8G/o+C+rt0XiwvRfFjhihp
LuLtYO8Q7TpatbDsjHk9NiL/hFjn42kaRTFMZWg7VyQ6hZCTPQjWDt28R2qNG7/t
ejzaZ2LN87yCiVtzx5c0JFQRq4zhZdUd6b2BAwpUrUS1rWSH1UvTdhKzPO+7Fga0
hTl96JsOSdBpssssAaoummW4dkXGFY8bzNnOIrxkq5Zd4Sw7C0ZDDsgLAxQKGfVy
W9mjz+beKQsqZPzoR+cBFVxZSmqF+VB0C2QA0r1OSF6LBgqj8tnt8LmMF/F9oOH0
M75oSccld3zTq9c+caUKFcLdd6SV768x/ZPeUHeOyKVSoCj/U1tAPFLUPbbE/JEk
ZZcCgch61LdZ5gwvUnc2DLPgQVRT1BJJOsTz15Vd883h9fQZlf8/MTLInAuq6Eht
U7TupcOtPxZCZhsF2aAt63eNUsuC2moudMx5KbbpO2setSTvhcsFADlFnfXyPNrE
s1Fe8mOk6ppwHM9h1rQinJCK9keUgvgb8nBqoDYBLgig6IFNNARU4T5wVGxtCFFy
wF6QnaMNaSC25dqCv0o5FH6ijm4g53TjesFDWAekV+QrH/BtpkH05ZqSmL32nYz3
JTfaCMq07jjZrO0kcOrAnZM5DX+rac0wklBWYmXcyhiDC44kA1zm0I8HFKQsQIrH
AMvkkhUqNCVBL/UrWRgV3AMCK7xLk0wh6kszOhZXsO6vnC+p61ad+pUXPstk4LcY
xY6xhILcGc3F5GDtGnCvKqvp/fxkI7tX0oYoEmeDNm48UJdll67UJf6ZokffVa7H
05ieaNBg8LVpnSNsS1yauYdtBNJZFXZ59bs9RKabDbTkmfbqzj8Zr6guu62QjZfy
q8ETlomM5bIYjtBKDx4sPC4/ujAdyZ800WIlR/35gJqxwNejMG0JJ19aOFnhGlGK
k3VWBRPGVfMoSDp8vRn5sQZGxlbMUqbQnbllWmJu0IYwbQqNO0i4oeamEldMPN9Z
LEN4JlyLgMFsyQTd5fGxg8kWASYkNbwCIXEMEWcjD0Ul3nZJ5aU84WTzjC36LpnO
J0KAxQQOuMX/Y0/hamPTTvQqSrnM0n+Iexvo5a/u9TH2LwaSt203gLWGax+H1Y6c
cWsMAVGtoZmVIYEdyRzKcHYt3kK+LUV6SBiI16u8D9Rup3+hCq7Hlrn1cLGknLtL
Qh0gBUBs3tJeeWFMmn80uVzr8XfwGySRiqzBlKL34jgTe6m7rISaDdj6IbFWKxdC
8ZEHJirCNldxRm2J8Un7m8oeVZ3X1KmHS1NRm2wpewlYY8Z5lpOnOgS0f2UAJj+W
Mt9T+yR9dkgy5TOZrJWCTgi/dohpuQHe25ZxkGxPG050fYrMCZ86I+xysWQJjJwA
721dD7opkAgUq4DuhCGFBl2NzPBAnNdXab2VDM9yHZCE3+qoyv3NY/eeDSSIqwGt
/FgeejSVElt+hhHJj0vyQ17jL9OZxYMedhE2BxfSPlybshDegoHfujVvACKRpMGE
XpYVYhkoQB2KIghJJlokNLYXqwHqQbmFz9OUIqpo03Rofm57a5Oftrvv3TVnXRs5
C3VnORZWlaEzCR6GtS6OUQ7aQIJ97h0GcTBb+cBwc8M2LLDgy7t+5rukz9onUqKa
gCcXdKT2ehkeUvlzbAikQSkbQg0QcmMj0LyOpgQb3GL6TuB9awBVchr6xkvNztw4
5fkF5U66fOSbj8pZ6U8ch5+sdOOAVqA+Mq6B+7KgYMGXVy72ERZI3CqRa/4F7Q2L
3GnsvAsGqq0COxVLb8v5Zt3w24nitmle/ReiLIcxLIqL/83gIFVhQW2+umOrbzqf
NNIUk2MfSavbp1fNVzPd/Bf7AFIPPfKRvpa4Liv4fIAvV/1eoAqfvSkiG41XC8sx
SkrRmN9z1c0K9s6zZd6ZACNyCzaKMMjbd10cmKhZ6iBKfQ49KasbWE6hf4+yLuBe
0sH3APMYU3hQLfzB5D4ubHvd2LRlgIZHTw50MFVbAnHOrxt8ZfsIV1sfUnvEeivm
LbPHKtxGZk/p1tRQuIAAjwHQ3pXtsrthFmWJHkZtAEX5ihVXHB6eJRmhVfTiQRwE
QVzeud5Xg8iDPltA4Cu1dMkt9h5FZxqXYNVyFVqfT+77x2ikKi22mBkndEsJbEIz
N532E3CNkvIywr5BNCmkwnGQfd9sLeWLF1Kif3Q7d/h9phpai3XPMai9SpFele1S
+6dPxHj7AcZC4OaW9jRc0BVGhSwngeJK3p1CyeyNhmi29B7AOj00GIO9woC0biss
tw6y/5UTfmp8JlC/Nngk6PHzGEIHWjr/7EKcu8a4EMbzqA5rbu+nlN66ugXGudmH
a5YDsKuxcoiYvQza6L+y8aKLratsWRP521YJcV685U4S9CRekCHf42M9Am/X3nNY
tyQTVhrLCscU/u76b2aiPtIfJ42dtzUhMdj+DxgVo1G0YuQg1oMhI7ChrRSJjXd7
1S4N131DQOLihP76qfS/pJXc60wyDRviL0rh2AnoplpFZJMvH8fuwYGdrtdhQecp
W18dyDQSBww1JxxYSfvtSqHE8YSfK8mW4FKTNdNxu1oRAYguAW+Y95CROW6UYp48
JvaZqf3EVfCGElNg0c0PLQ2I1rEDzSizGfFo1Dgs7bFuW6wTyny1tpSXYrrZA70T
z88K5Xd1EUmx5ALjlxX+vSs1V6KM29QVwzx3jfmTBsA0YLzhcV+bGzV3w13zEcXS
uy1hcwft7znvzJZnHdrSinl4gSkED0jaiKn2MxfOUCuHpj6+ULKTB49iVr/ymRVZ
/g0QJ+hU5Z6k+pgfi1VazV/83SZfiY/a9M7//4ZJgPFwyKlEQSTRHWRLN2d/XOuY
4cdH3eVaCsuR6IYbJ7rGpP/OqDYuuxfw72bYWavf/+IQLQMUiDNjjrrNJWs2ZBS6
v0hytj4J6V2eNMXEV3nDgFpaPGJd9HSw8aF3I3wDQ3Kp+k489gUxTNyLratHOmF0
Ige/lb6Nuslix9E+DMqyOjB3ok6R8jdxNx/4o+Bi2bKKRhqFLJFyv5E+X9pAfJrN
7jVbq+I6EhysQ4rkHXSDSNAwL6mEUuLRowUobbTM6La0sJ85HND6eYyeINXI0cMH
1elPnM0S+2W5G2vig2h+rIjCI5fUnNECRyEM8J9LTVlJEVnw+Y4jhVr2vU7TS7NG
8irE+9u20GQ2Ad4B4VE8fo30IohEK51hePuv2d61rAwThiDvX8ShBJAWFjiHi45q
ICe/7dx1a6Yay+aS/julMkmG+oAXNjanKPalCn9sPnQ6JZKKBr+ttXf8kPPLOFsh
raBvtraOErAbJtlMoiAVuJvWjhbdl1sbFDXduV22aFn6H3oyV5su9IxHGd965g6i
11yElYM/mj46AvpYdNBaYrh6uTJUxCcLranbmhfCKV3xHmOqUKHPSce0n5ZEIhlF
Mo/foOTFqvg+wPeWXlfK9YnQT6IuIgWpn94q8eBHAf5jUNzE3YkV3AoaQAnh7zIz
YRMbi1rrWqLzS6YbojVtugq52QT8KaQq9oIT9U/HMo1CP+4e9X6VhqaNxd/Db8bG
5Kh7TejxhAT2xCHqsG324xrKZYPOOQv6Dvg2K2KeKHsP2kVxuZWYUdE/9TGFWKCZ
SZFmqsfTWQh2BL3t54V8+sKsC9Kj2liKJOCZlQnRP4BuawL7D6+lBFBz33rqilH7
axMb9BLtUU4NVCwnF8s9SQ9L0ifH2zv4WfnH9JFrgnZyZrdQ5QZT8SecphW8bqqn
pxkR42twJjCmp+iFcpN1qcLb/h14pfxtd3hk7c+z344lD6GnlIJUJh1YvwCjSyT5
lIE+0UwGdOArl8n+KMUBXP7srX1qRcirlGm+ndBfxzxbngtFQiOy5x/AO5/CsD8w
rz3CklWYBA7ehAskioUohJA5JRca5Fy9Ll+oks2MnOrdTvmOCdEnZtNehnRatlJ5
DsbS4+fH4CoD1eYok0US7jRVDnFBPRVovta60NLfBYi8KhXbID6uPQ3AqbzwCah1
iw+9CaBp0f7riRwvcZR5TfXfDHSvMdtG9zDLeLNvRxPz2oVbLFJER6Ho717F57dr
lxYMTdb/QZbVYelZ4IAsWA0H+hZqyvJjxfDZ9PnDIYkMtEUX83i2IbNnqBh0iYIz
823J7bKvx/+06OYU8jkEDY5psGG6dT+VBz1kuyU4X/lswlCKAllLUg9bMpdMxVq/
TvCN5cvXntcyu4znxGUc0Oq7f4Q7wqrY1qRq39Gcave8qLqT0BppgeDwN12NDGfr
cI0sWkXnNI9YOjK0o7X0ick/+vLB03y7oWrvuCkOLaTLcOm7quyYl0ehteNf9ctj
aXflfwuLoeJQSI/41LcdziIcktJeKnUgFXEYCefT/csqYtxYNSmvlr/Z9yzXa7Nh
BE0Q+9g1ICdgn0sa8cy9MiTLmUNRQN6y3uZWk3lwJXW5XTXXNeZlbUZz0WlHibmL
bEmL9P3cYePMyJe6/u0I636ByH/EBFhCmWjddcmcySWI7nzUaQ+fQfmOdavFRTNw
bXZ8LnJ688svv/HPCnsU1DU7zs5BVXVyhBOjRSRTi01tPO96AuT7WE3ufdtib9RC
OJWr4ChuyeGyfCkYLob/lGgb2gmPaIB5NWvWbk/xOoDpTUNksF2GXI1n9dhQWFnJ
TZup4L1l0Iyr4HP/GAYMXN8IBTqbTwNhn0zhk4nwDSWeuWhNkAHNUYV49jdw8a9h
qO7DXgn/IaUnC6Q9vHhbBz2UtmrnIobDIV3qWqjAeiNNtJHRatzu5O0Dhp3YO896
G2aeDJV0X3G9OwpGK5KaXw09kASOAn9f4hmY1NS/Hxi5OnYhaQfvtD30f+BeoqAH
Zr/ztZl4viuckKJ+ZBqsQTUiog3JPdlEeplyAhFxFgs3SszAiK8sDF98m+wAna/O
i3ON4MxppsJs/tv0DfxvBNro/b1wNsnD5gC8InWurKNTxHCeJ3agCYDja0WHKvRi
mHWn2NV7/h+uKN4F0gf/7hBN5DYBLUrVeD6ns8VMM7jaABsbM+GC8qgZCGMQm/rl
K5vvobQ+++otV37zy0xWs1QY1cdwn+qXjLuV7q8sarIxMPc49GxssKY/f+/XbwEA
5D+THrtNG4Aqho7GAKeQJEqYDv/RtFGuAFcLzvyiEvL11OhSsj/YEY+o7/jyOYbS
cmKWXtKsJK3PdaZ+ZSvvTmC7rI48sGB+kaLjo5vA7+TGI+KvBHdzqndL1tjPQFm/
IyZOesPzdUVNzU4BnXZAt/A7zwZ2mQUDNqKFVbg0OBd/7F5OgUY+kdShRoFKF8so
59uSfp7GA0hjaFkvyBVA17eDfSaTkLacj0ATFjf+n2ly/YicCAvlkRueawY2Av6i
lyMrQomF3nyJ76hZD+tB3wACkB7TvVpcyEVPq1waTX2gjBG9xqOo6ML5HLYLKbz3
VwyF0LY5jArl8KpgcwwPt8yd8TAj7T6POiFEf8F+78XOQ3kF0Y9gil/2M3inpsxx
dbt1DYRrQG4zz7nViaA37K+Vc/gFejegC6la8/1Nd8PnunkmIC6Fn2MlTQUSUzse
7zKvn96XTX9Ki6Z4uxGVS4ZRr8SoBD2dyfpF65lc0EiL13uHEDzVXngthby0Xcwk
Qp+D1TcgD/A0WF7UFwe2j3nKYqmtk6SKM2PeC32h+sUf2KBPo47bjhVCCcrWBt/4
gyOWPCeOdqDoOyLBbIDq5eZ9gIjROB3z1napkS7loQAo4TDPw+mdK8WP+ryHhvhd
FC88iQvpTZS6eXqbWUQVVEecmQopJ8Per0cM8iiiJM/2UsR7d+PwfOEhO9r5pXyY
Tk2dcgJ6zvOqBp6/f6DQwjtao3X8O6DHpwZxS7kQoDD7sKlhBOXgJiUApNQruLBi
4Lj/wdmP85plWCkzM1HnEz6Adoz16vQleOd4RsKOXysSySlkB4P/xtsQENMX+ZSa
qi24feTEhokq8PiWJoIpyuMhik/W3QyxtfpYJwYggQCdzv9xE14RZAKcQC4t7fP4
1t619H6xm8rm9fo4EWZrQWf0OLltlYGttWl1u3jepVtL/W2Macj7wMwdmesJTlpA
pecTgPIDM59amjc56urK046ZQ6YC3tvVvMInYkqUR7Ju/+BH1FDrtUz4aIlK3xTT
FwZA9KttBpmnFBrIF1PxgqWxNMYk/OBaMqNva2BXQd6RTcq39VIX8n7Syf9F6wCD
a7oHVPmK+rq4gOTnily2gQUE4j9CyNNxRsEAAWlND5htG0OVrR6YL0wwOPkWdTi6
03lv+UGc0M3IGL1B7of1VXU/CNdjpTqpnpO+Ct4T+kr8HUn1WawbqQjiZTLSGSIG
vKKd8dk+G+4P2nC5SFBGWaEutzqoIBRf8RS5lP3CsrDFZZjc0eAcPaJwozjG7gKN
37Q0eNGaswg860TUfD6QgMFPsQ8dtkO/Gu0TpONG2zE9R+46f3tfzXZrjjEQdlp4
acqQx5zoflb7ByGnhCnQ1kYVz6rN0WViHp+48Vtl5aiuy3P9Qffn79EQbYl08ZSh
G9/YlhdYLKrayp5JDXCA7fR0S7H+sU9onAbKrrz0AMhgVdwAIyre8/fUAaRlJDd3
pN4WseCCfSqVZlkpv9lwBvqJ/BQrEu0UJm6wxDsU6xYkkv6x8fbRlV9TJtKPeW+I
HEQEprbRxT6LsQ03ZcdBeOFzy7qb0N/nYxaudtlPp35A0PpNhbY0cw4iW3vVafua
WC003K0mdPaKri2dXtPi5Q1d8Zk5TKhACm3jLwqDmXJUI8Q4AR4s+r35PfZQ9PJq
YDelP0HdoSr/W8Yw2jNf2LPg1JlvFO41bxq0xskIKq45GRUzM5r9hZJKEBph/8p5
Y83BtiEb+FncWD10v8LIaBejhrKoF+Qyk5AQi2seJUEnYR/C75Cf4XiyBH5XoBpV
FSCghg9l4Lu7Qv8NCRhsKIO2/UbVUQUK7L9wndJ3ZdQww36ms335iIlQKLPm+YDs
zvPHBPAZMOPqH6KzzKFxNkS1lKlteezTH3rTvvrM6RkgNVv7xbfbVfbjaD2haapw
+H56B2tu9VnOBaOZ24tlq6WzGSEPlTiZL0QCTZ4kV/zmN4PGyfgkYZuSIBeRFjUF
l1qCl1oX4vGZg7VeAa7fIVSpeZuuIHD9KzfrIl4Az6yci90J5Df7Wu6yVxMFiP+V
YCw1WMZjSYVQY1fKShaSCg/hyTT4BsxMf0tSl929UxFziTPAdApnVFLTeiiNjViM
/AWGqfE+CYjadjuqhXu0eEMcmEP3hDU4ngPrQRYk+IM9KNs5St4oVIXbVIGkRPwQ
OeQI+QNMyHziUal8IUITtCLbj6inOTp548gn7HMIT10xTyg+BcctEM2ULz1PdIOk
a6QrLZTRRc6R9cj9DRAnEB0y++TNStPY4zxtq4u905EAFzUK6/Bp0lKUgyaAWNOH
d8OmQLSSdKtXss1n80wpPjH8JHWr8LaUZx4LAhlrUlCSVs2/52zik7zJMB8BFjX1
MQFpKOhpOVN3uoKOSh69NlARfCl00XwkYctAfCE8bgEJfbYttjzRMkm3OJfoxZYG
VAshALOUl/RsBZKJUhdlFAWgXx6Pdp/mYDpk4IUffzsALzs/HJ2zxznkrsCmIPDW
kNFdUNkvrI4xkA6bLx/AjhX46gPGqjGphN81i9zP5zlmMhNQxR916zWkNHTRUPFc
VBrLGlXfcSewloprTmie7rvV6d/nfyAOFb80Q5Hi6v09acGaJ/yBMCJ43SobN3ay
TlAJids/fDsq3KA4hXi3AfVPMU8FbsvJjF6Of0vTCM8HNIGM4Om0QvDb5Or+5Glv
B+RB96C6syUFanpM75uy1S9YS4nphl31/z355YFeIkiLFSDL2hEF3cFG/QHNz+uf
dEZUktJEKKvTvuk0kms1zCZmPkZlTJWvES5AYmcVuYspAi9Kv+XnBIIYqCboZasf
llNA+VzMlgIAJK9ucy5DfgE99vjV53+HbJVlZSs6aZy7+Y5q8AXhSeHDzMZCiqIK
e8eH8YvgWLmbSiJWae5qjuxg5niD38uFI1/qvrgJry5nTmfEBz/o5jzjuSJPdjFm
ttqHddFZGF7mayaRGl78h3CwbO3KZHUuo2RR97itptTBcj9kHJVsx6RQZCzoXkPI
85Z5Y7ukLz92/byZ3RhywhrA64qS0sphwXQJIO3z8gMBbh8XISgOeeTUy/Dl7IHC
H7n6GCDQ762NSRGow/3IfCwEiExTwukl/pg8mffQBDppHcMY/lJMeMMw7Pn/z3cn
W1j6sxoVKPnOwXDzOhQnrFB9o4HCYOvng1Fc40ICYfvYYJLJ3Ap1mV1p81YQsPcV
cJZwTXL/sqfdEQzjG+j3R5cGIYJMtL802k9DIMVOm2q7h1N7X/xhLxi2G0evnisi
4on765+yK1+gpgwUWF0KAchOWM8VLQ1Kbr1IgY+ivN9hcZKVYndFDZ9ntutQpJYR
XckzuqYDWDKFqqChHrLyCD1cW6YZ+W4FmZCzNIvt5CiuI+1i0S7v9Eaw8OhSLEwh
FVecI2E/om3/N4/p5oufX3jYwJonpB7ZGbEqsOMrEfOsRWVajCzlLgIg1NePbS4L
uDeOt5DxCrAjUVD5Xmm6zTIDxUWOkMyZUTYvCOgk78c5hLEqEbwstilc/TYmC2V1
s4A6iNNKhOeeC5xVrkqxrM1OBW7biVcR/Fb5wVJKMbTQLmi6MBV+bMeyIurGte90
J0nFR8sU6IKC+auG6B8BKNpTQdgUDXg2H9Xg4En3wYwdx7UuO4++lKeGFwvNN4r2
+lIhDYzbP17rspBhzV8TfVdTCKeLcJMxHr5YB7KyQAy/qrY+JXAYO0rGAbmZjHBE
O3A/myV+zlopbdexQoVKG7FFNbBNFcmCgKbzEJvGvyo7AQWTdIyOpTSGEtIImp1u
TFsMh491VxK/7AYOwAntoXWAKWRPhEnhqZmA0rTGbaWo3AgTg5iXHyrs4iQ+0FL0
c4QXHT/gjmeRXqSavryuu8dAc6ybWIEw3R1KA+hdu3+3HNEwUBzrq4vpwK0hPLeN
ksSDQQ8ompymxgiy83aay7ovUrqW1ZW+tS3lLc+HD5dss8VGblTcySX8gp5dTy3T
Y36aGhMKikE5Ce6RzPFob9U6K1eydT2SUcZCf6piLqVbxYZLdQOolNDw/WJYTcMP
fxa5YPYMXR5r2lFfOQi8+UJr+Z4ME4tytLLGYkS8uTlTr1Bu0C0+eFLlHqiTO9wM
hAow30BNZhiIEJ7vgJCwJrrzkA3amQILx2VVpm3q0fFglK4ifFS8cCiQDpyFuUYp
3r+MLkKUmRk1yKt/bZ/x937IDV5ld8YyEXGleyf8DXF2obI4xtpgQ3rGGlcQRVdB
5qJPlC9xXoS93kHMxZUgpeYbb+twEQNOvbuSEGmRSE9qHdoTWXt+sd4pmoEdd1Mx
NvF7kwV+WtSwbLV3dH6TaH7ogY1KzAe0oEnov345T+S7enxXvzCG2bo/PNyAq6Tl
8kg0xWCcIabFlmBKGWr4r7Agnvn2+tljmNsQKRTM+XamZ05fp3Opjy+MWlbLgxn0
fRAjvKYQWuiYAbZKby4rbltW2Uvxmx51NKQ1Vbs4HzuxT7j+5PuyJ1/NBvZgJMO+
X6mtwZ7A2kNpCL/foLFh/m/LNVdkK0QQ6K76yOINvhhmVF9gUKggb/nza//a0dvF
C0kg0BEzYlWu2LRpOZabdIZ2wis3WiGywdrJImq6LmtfJukclWTEk5thcWhFkJLp
f/SfKZf4Mkms4x/saNQLYUtR4FffVCQa0gusQZ0LT+NXlwkP888miAwOPcjALI8Q
H+TonLZlJkQ7ONN4IboSbcLt1m0u9uTVQ1d7N516Bb5PQj22Qxr/0vYBxI+R47S5
7lstT5Ct9lnPUB/1aNNKto5rLjlDTpiNsR0/5HKPibsHJ6EYgsMC60VBSCgxNDn6
QWqPCtZp4Sg7JGIwhdBWJCOkhu3RVqHyQEWCSPC6PFT2l34LdeJKHOntwI9vBVtD
nYvLeUYs7nRKnU8wrnTMAQ99ir/NduiKHMNGWIvSvBbI05xRqipzXSfhDaP6BkfR
+OPE25hTylknT3VOoucjUdo7CzTaD8S+//rcKKyAwhar7MC5+D8x/ke5HkJgDZ18
P0v+CVjyuUGZeDpZiPjCc5yquEaEMKFLZCV6EqR3cWcUHODXn5EZoLpAoet+FbfU
kBgQDXwTcyJVj8EW4jk1dZUjRUZt6TGb868yf7pAIBTnHk2jURKv1PeRwmVF7QRb
Eci/mGNMcc/7rGUzWR5e2VOL8X2mu7naXfUTmDlM3JBaCnPm9LgosWvf5p0En1+9
pOOSXolzAqKXairyeIjwpMVV9AtV+hD5apkuXcVhONLj+qzL+vr95Nq7gUjDar9+
QGOwg0UpyORr80q3diy+ID+v7XLRRg2ZddY6vXw3oAPWUpdF/s2k2z8dD0p37vU+
pQIpAZU4j0201X5/Lvy/utwww3OLyoE4Klp7uu/rblC0pbOVj75R+Ha7ggq5EbkO
k+EEmnz0zpZdJaAPuIQrOnlyxeCUzbz5nOJM5lbJgKHQNTL5zLThTh413/ngYmEP
Pxy2T6vA+dUQnAABJ2UzLq9KVIZGaxgWPg00cnl3/hjL6H+Hxi8/VHWGw0qQEiKD
tX5nfs37YFHdHsWXRMalPf37BXWRfq88bjjpE/BQ/i7aOccBo9FqnAeCb9KGk7EN
uVbHNPS3anwvm3y3U6Ff53GGMKR0GPrddyYDYkE4tRFIfERN8lngDlEEn1l97g5J
BAAhoUzyVaYwzuJkws5IXJHueXewONRpNTSexNRiq9fND5MucmsJgiDAnlHPnros
lLZe0pg+qAtFkc0fbcnkUL5NdSeZSsHdSfZ7RTxu5oDI9ZX7W4lxclVrwAPIupfS
INGuUilCfP9angQQ9yhboU8+jkwD0D4Iz4WNoBAFl/4vqxZezuVYRL6ZOGXCB3B/
qfwNvbFrcwXX9UEjBsqkF9KDcL7cQ2VtlIZjzibyDPy0F5ovVyDQDu1O8TS5iNiQ
c6edf0ISuf2e2vjK/VbDiWyoLYZ6cUFBg7dUIVXUqH1xunK6BVy3yIvgCoBhk+E8
vbWZZk3S5YgvFK5jbBpyNoO96XyVTPxteR+JCjmMV3PrSw6LNQhy0F4/mgI0JtnQ
KnENFP2GdBeig6fTq8OtE8D/i5NrD2tT+f2o6x+Q6/UsyZJuYq83yxLVAwt4Lr8l
d6XUTE3rowrYKbK1W1226m2IuY/GTtSagi8C+33RPxYk1sAVtErjN1XMuq23XIPH
/OwwFIGlNs42xgKtwBZ4GwRq8KMcV9FbDa3oSasHESNbI4/AAkBKpq64Eex+pxio
+j3YMLqwDNGSisoDJ8yBujOmIfhVk/cV9rixgf8XWu91PNtYh14AnMLWtZMpfSay
kn5TgBu6nvivf5UA5aWvfhvPePG7boM8ZnYsfF8kZtC0C2Pfa2KhskXl44jkQd9r
77m06Osydz2mfn+3wUbaq+9DaSbLfh2JmvMYyMQkimCeETmu+ab0ujPupEReekgB
Og4sLI5dIcaml0bsMP0GawbA5beciTkdL1X6uFUzHW4ZSYIvp/OU7mu0QczrmAHc
ROp5q+1MK4E2IPW/TH5W6JHX8oNtSREsgkGLFWfUCipDWs3ovFzZ2ZXP5Il9BKP1
40QCHS3gxQC0cXoMiXShH7XIshtM0lb4l+F/twJoAuSnBIOusa/E8HrMK9qNYlsG
cShJ8TTZrU8VIhNGUWqncE2exH9WEsQZPT39QWvN5ASqP0h/4MW5LrHq0X3G/har
oazuRwGqLphaSx9mkpiQmjnb7XgQD8Rhzmydi6ljqKAVeHgvvsk/3/3R8UhJuKsR
l18ZWT7uetSYtaiC1Jezq+8reIfpMmx3EO/7W3XT66TQ+/XJ2+6DFhQjuH0CbYFK
IP9XW9V764HART3eUgVgkgLeuUdcVDHJKGWA8v14v6o7oxY/BnSKr4voab3iuXyw
FqbzLcIM3eZ3cBZOTCwuu+nxKL/Tdnstnfw/lyvOz9Kmph22uFFYyNNyvGEse5fM
CI1rUSldGraiNeUe1GQoQ10gGxVIn3TLDeJLId7s1RXYTGMVlQpL/DuuP4Z/S7rv
qyDxsVyQ2pkZ6PmKkWtGfhk+RGSqrp0BMDYtXuGbVGtMSVJl20PndE3eaDTRunWp
t3dAvlzNQf1vxsUymGvQyOGLhnA8ZXqVJhKKsy/835MQoKLCXz6+39tVoaeeIW4a
aN3nURmPSvlAdzaLwlH/bEY3o118DaU0/geqoRdR8oB3G3uWI6l1y1BR99SsNsNT
OADE/7XpsPNphzKL99wc+RpVFVfub1wd4xUWTgVJMsighrQtmmzLInTP7QU3SQlr
9MQMTqW04iootf9XAKEOx/IJZ5ng9ydc2xUbyooYbMfTwKketHEna6ktlnXaqNo9
TnHDAkYPLOJbXRoIf9Lnn7BrIXQ38OAB0CJf630EW9eKpDlsMN8oV9pHrBK9JURO
7Ht+ZIjQ22bDOCgFNJRYWhO45BGSZ0nzfAYk+JT8cPrVuDzhpsOMjDvp8qiOJW+U
deWkoB0i5x/cLMs1nYv1/e8a+wjk1wOM6QBoQN5Y4ti7Qw+0mNXCv5jAkmwEelw8
Pn30ubWGqqLRR/LGzmmhIbzETO39RUpw1/WlNnW1HLjfmyrYmaIP0LwH65N9PCnO
OX8p2Oms2ZCdVx4Y2/+brugze9nEwP9XWyp0N/wB0875nX+mPptAitlpSaaxRYa2
Skmu0jOBl3gP/O0m3jCXvccXpb3mryeyBwqx3eDSHCE2QcEvwYpIcMT9UKp8gxaQ
jkd959BwDDt1o+iI5qGc6oNAwl+PuP6sdDops3Qx6TfzHuWxogyvqKDTVrqeAGDF
re60oKr0tzfjH/eLWrBhat0pmrg51CWMTACsXBldBDcG6aTuYJ9lmxiMd5kQjBEC
xqWCGThpxjHd7hqFT7SZuXHJMYOYqEdaiopelXprRfR8BLY2Myu688MdFZ/cPzxe
EnDTchOXi6W+3Kh6N1EIDhYywhIFflJyFPCK8LApiYUv2jRTSq+3oB+hdvnZyM2v
CGXFzP/uttDFjmPnI/kYqa13GNGZ+K5CN8f8BjORZ8/Dp8JTd7WQjwyuYvNbjiun
E7lumwxczvMOjQZUyon+EePYWnapsBbwkFCrPwbcVkuFvE1hBziZKdYAkPwN902i
ZJqrbG4XiRpRbTewoJ+VdoCKUd86ZATuSBGsJlbGu/GDrcUgTfUFzB4tVVgLdgTN
U4+BLpti8xFKy5hZ7L5/9ntHMVuF7Pde7lS6ivWUkFMi1i0DRBHsZiEoHNRvWxvV
ifVgf5AjYYq2wUV8oEF5zVqWMwdT5W5L3h5RlFBwi5eQvlRpjK8VLj9N2r86pDfr
LnxZKBugpZkeIid7t/CV+BE3tCkCFYOXYmDZ/IA1mDARn2kcIfHOTvsm2SoVN2X0
DUTCKxgAPTtYunCFyccZMRGQJfBOITWKqXR7D1J6DGnEbZ6lcELESdbK36VjJdmb
6w89IMW3jKqre3ERHAWlHafoNASAab7z3Bm5F/DCwb+r7NiGNpXniTZZffP0/z2j
rmpyINgQnwvuG7jj5SnuGBsfOZ6JvX+BTsctpXltRyc/fy6lDUp3mu5Jj8SK/dK9
sHp3kHwUYY+v7JIHixV6uSFgJNeU0z5+LE57BBH6E5h7ODThHw+7KLy1gPhY2b+u
1GkhUkfsAvzM/28p67qA1seJkon6ezUVLZeVTIbnljbknfe0wFxstjAeSRGnicyY
zPwva3sQzKUPmIluNA0IUkxH/UlGFqOiLBXmo0igJZQ4OTsCaK6TFWL8ULnWgZGn
0h9uPBMufJ2hTiNIkzoStblmECJNc69kUV8c+Ex4pYHVBfh0QR8hdur85+DGf6Ib
jIHYNbmh+hnmQ9a29cZgbbwlbhEn3e+BSVGli8YhwwmXj7ACmuuuFzMZZ6E6mJEy
26X7woVZ9Hnxi5rbCuBLI1+bcqhL2f5lujJt/F9vyRUaDFzRfmngIZDHOSBT7zEx
TDKa1WnyvtB22+6gM4g0r+f5YfNhShhRCemfFWcLU9ZutD927ylJO4z2Eav1znJG
pQBkab8hNVevPqa/YborvpyQ9M0L7Wk8NBOlAQa5KIBfl3V3SewhBxoXjsKrjkNE
rLZZbUZhf7BXOKXdDlZGYQb7VqOnHqdWACFwkjBkW44txe1fWWlgrwXRxSfqPT7c
MaTfjA0OwTYyRzZpdm58QkIVvYnntnouS8CWbI539qx0Cng2l44ZXCPFiAt1a8++
dJJIs4W4MNt2xks/lHm0LS2LCCLC1I2ha3FPvzERCQXB1flMIW6FvoY/tL1O66jZ
viaKfjK4GmFHMnZ5KtEqi3o7XRMGpmcIov1lQnJC1PsAAxc1hXC36f5t+JdOmOFm
KPe2dAzmXS47aVTsqc05Sb0ZwRXkdcL2/7ArsrhBeQgyEHN7mw4doksu/Sc74Uaw
4rTkhn4dIe2zMdro/U8TOUZ86AD/1Ne/MMghsBXoXJB3HFmlkIBuFzFSzK2CNHQK
aYQVqu1IgSRQ1fg3CxAxXTsaYJ5fWOTDAg+AyuksfHOpLjNJMpdeGT3hF9OAgxHI
bZSucGJ5+kv86rPx//A7wX2ULQ0dIZcs7VnnM0O/4k9rBFNUJad+Srny9Joio5Ar
jcRf7xFQ1EzztphWnSy1oMHuh91US3GbxnSoL9bAEkP3Gfym62GnRHvEfapg6qGE
qh7Dt/X3O7e+dvKgw3vdoC07GHshXtnVRHZSfC8UbuncMALia5aSdAOBmMo6Oae/
+1KG3tMyv+yPlroRpmEqhn7S9FAnbkIl6tSB8iRvXNCYoYNsvSabh3gB0yNoMVZO
fTmSPENFNLZkYSZuSCYhH1y0DbTxGiFvIPjJYQiQN7atcPP+sqVW1VPeSNyqVD4g
xQogC3PKnRyP3s17n3r8+fzQ0QaO/zNUKQvTm+msdECdTEMKTqxMzlUni7tOhCev
mzwT1+vSVq9iPIigM7Y0j6EKG5G8NHCKcPklh+1KQieQqsrJMPKM/0OeRVEFcvgq
ojs517IUVjn9CzDEYDNnxm01ZL/MgFjIAnDSNlEhXn0BMfYkXDOKP8wn3aDRZxcl
RdFVXXphwtqr6UA3z6neFZhDjU3THSvPAbNmXECwP+MSOMuRk6In5hqggyZGO9/i
UP0g7Bp4UnhDUPEiO/k2z5CmBccarpy6j5jCJ39G5tsFycl+xdIqcFSWyv7wokBf
J1myQfR4i21RRq1ZdtD7cZnZAn6JDYBXUSa1MxiHNQdLdpRjWMJTZZG21x/xVuJG
zon/nXZ2xSLb6vSaGenjPid2OJd6M8HT8ru/zbvx3M3wqHIgzBmwCzJAsffCnzis
PZcAVMn6BYdutM9GaPxUX8STFDUSe5CIieuCu+xn+K5jiwkjoehoMMRMFzfIE9EL
0hJS9SzVMy+QRop0YzVlxdxiv/8GtzCYRJS3v6/ZAUuDx7Zjeq7sZCuawpl1fEne
imvFA4EhOlXWjgcZEzOSorbBT8Ii1Ra2YupNafQYIpDPRoawJ4APgUMPClDV1/3j
6ZQnpCmqTbCYReO/0prMM9bE8mkRY4uos898WMsHBWr0C8isMrMBeheQeJTNpcJL
2fxHvlhltuyoUmRuiSR0oMN2q0GLbHXTaCpotxebtQndxRB3w/kDWw3JJXGwm+Cs
wTxfzwnXkybUDcUxi8oZi5USxNdoKgbH1chfxdzFoAgLwr/RbZj204lTqMYkRFv8
RfEMbNaANkhlz7eNBreP/ouf29ibN7ed9IOiLN2LVXU4UYqTd5c0pxVGM4plC1Dj
X0HeMNjXH4Vo2UG2tLsUt/vQj2Av6cuC5huaLca6ySfwKQnxKZaTPPu0BefzmLt0
4opywDMTl+w1GrvQ1yZ6qJ3ICoNw2J++fXVaqeIZJyaLLzaESv9IhHzMRcz/3xI/
We5A6oKfShX6sifyzfmscey/06OM3lbEck3tZbsTnd9+OSLYvAvb/mN8KDu6e6I1
4b3rCnDgD4v48++c4RjEGA1aYcK+IEU/HjLu52BJ6kItOOkFCmBF6V43l0pgZ7s2
cUK73sncjvpVS94MVoIinLlPSCjQsxPB0ptxvn5p/KfMjfdyIXr90cg7n2Nzlmy1
ZQTgwQZPgoUh44zyemJDgqF/dzQ3uR4wP8Czq75/rQZNsEEHxZjxNmmPCqYjjHMc
Ofur9glYGC+HZosGf0g57yiG7AN14jQ7GNi1ds7375093D4R+ssaAtjCe5E2OoFk
G6DoUIRCuH0XzMjckD8c95nZgDh+IAhdsUHzIrWEuJCB7EtD9MxcSrggEGfMlVL9
gthgnJkdPsf+VRRfaIRC5CuGKYMxxFfZdN8ORT4A4nMIATayeBcnwx7B0S18Pt4U
NoHhNro/wZgVz4Otb8xBC6ckapgj3WqTt2+XILePGHVHSSaLfj+XPJTkAuhOKLy0
EPh3S3R8rz9SJTUtnUTqLMQpRtZG/qfwN4KW5GFZacvuFcHF+l3M4bLVQ9FGLUFu
kUEEFS3mDARvIQM3p0QeSULyprKLP8FdD+1ljw1UeC79BNeE5KZvE2LCkj52YjXl
wBG9/GABkc/VmFzClp2Nayg47UovjNqeSEWiuBrQ3FGgLCCYmI1mmBsJozSUD7EN
JKmA6ydwlxQJgsO3GHNaPWlcm18Ra0N2SKvmKjjOtqWpKethq5UEcz4fyA8OyWIf
0F0nypuagLMtyCKYU6k9+a28J1GlEG8TKmbYUUClWbLPy6ci7egW/nAJBEZO+DjE
U6cu+AijLRt/wA1eQsJhQr93OfPEh6nkjAP/6InLlPkLTSr7YCHKUpQ7oXE/vsRG
y9AzXrD2nA0K1F3WTh4O9mPdrpZjVoRJszWw4EnBYXQNvYgddZHlzsdlSFH6HlDv
PdoM9xG8byn1syyQpTdgP8UUWZG3Ci1CoBv1pAx0gYnyNONw0IZgI8MjIEYiVhFI
rPbWsG/ZPuHUeb6NiIPCYUyeVmeSsBvshPNymcLFZCQS9O6egqIEoyo6+t/DTzjZ
o9IaiKnyYcmKWymrYuElOSdvExXycnAIjOAr699nwQF4ZWeCavwCB/+i8BewMAzn
1tj0mbnv4sMvXX0caVEq0JrLjlMV2DMbvdgJC2T6PdwDhUhtf1454mPysaDRpNly
p86TCXLiF8tB2oCLd9Hzdh4yFD+LXTso5hfqiDbQnKw7D2ct11JW1K9jA5P25syy
O6GHzOFbMrwAfrwE9nH70nmMy85JMKgPG1AK++uIgF0g1WRmyJqYEE4zv81PEFN+
WLHYZqCeGJFWa/bxto0iaSYz6zCxgSQpLZdw+endyAcZ3sASRTEHNW45YtSFpoAq
7DQ2vYb3unpsGYmPNb1Fmm/uTbQdyq5QkBR6KeYTMK0DDs81LmSCZrpvXbZkmkB8
KLdWpvQD7E3NrPJdaXfq8sSmmeODh/XLpd9ns4XnhX5kK3A4tr9bFi2OJ1drf+nD
RmhL8NBmuayYPDnKMx8jcxWSZm77fXLldyKvWM0vaLcCUv84ybCaBkBtAxbHjNDi
Q0hObrmzLPtUXyRBstUbMLXAb3gCVKF1H+Os4IqFN7SzaxB/O4cDdPOsgSsTpqIU
aQMxLLu3ErOuhaPC8SV5KcfGp/jxB8HyT41WKb/+7aItGSewH+eOE441ehHttUIQ
5lKlZ9Zo4dWsOyuywaEkl1mg3TNsu0RoVB7AO1LFekXlXKhVLTVPVYPgdAIuoU+8
C0xstmqgexY+tndPlC8kq6qbVTDPjCU8tfEaubgOAMsnI+m24oMeOYwwlJawSn04
4WJpepvUyS3th8960grJKQdj6qN9eP74mV6OSSxEdrE4sBrhW8UaiHzXMy2szf0n
txsatmUX9kwqMWkHNu1n3K+mbtOZ7Vev/r+iBZPaDxwPQGEDgF/c12df1KphuxZA
Z70840olP2UzN59qthjVfN+Q7z3f8hMfLx2Nm4Rj4+OuCPut/ly8xsTlYsGFZagc
cuGp7M4EKMYKyGpofBLeAV580Bep1PLQJbTYZRbiiqxO+SJuoe5OqkCeGWpAPfVZ
XlkdQQHNQWCQGGaXjg/J4BN66yKQrKze8qelDSNWb4vlu9j8OLaF0xJXvu2cSPMH
AAkrwKttMnu7w2ZuAK1uko3eqfp5aE+0EoSzjM0n8h/+SLgZVLETRNL2RXcGuT+q
qvBePrSn0IWr6O/th4Gros94SUbDmuFT6GaaR4Q9xBWL8ToZIqIU2HCn0l70wAN7
SJa1VZ+DXfWFBQwkEm7QqWdCRR9ct2SvggJgfgadABf+xHrFzpUYGEoRIm0r7N88
5YxEP/SyRUFnLLen39X047WTg5zU6ejJqRk6ql12/24P+bP6v5oY39f82WWgd6gv
LRHCkHt4I2k6tDx2ITe5gaUFMvRuAxGjjixDM7PzmXnvQRHLjVZgMEICx6BbAEkN
nScaIot9gD7XXbSzdAUh+2lUCG8WsE4jhZ05r9egtoBVoNur4PYZFtzHxQWRLK7f
8Y0zeTw40dPxeQvrxRcll80/v8h4oOGdPkbgVec752Jx+1Z12X0i4N74tWl4cSvn
5+4G9y/5Q15C8igtcxCKQmDUCv9jmNbRTaw9EfzYV0gU7vCM0T65/X8dbc7TDUji
eU8Wn2gpxDp+z17E3MoBWyNCZ+fLkn8GF4yylPi1I+WGVDe/SD5UmUt3XJdExl1z
M0zHt+5w9EHb81PGohwYFfqkcIGlg56rJ2gJs0sw1C1OxNW4zThylyqWuZKOP7d2
QFfhRF6FhzBldLxyTHqqqVwKk/oIMvNsCImxFx0Z41qAYHJUvz8co49nuUEv+hLe
WKs8NBtpmpHdOC432pRkSQ9dcs4gi3bhmTCD5lwAPEWr6tsuQ0JyKmPDAiy/CCga
ldMGlCjwxRyA4ifLP2PlMy0GCkvPIxrJ/nJx1ey7H+tmSHeKl9WuwBxv1fHhwEgt
v0bbbZn+wjSSkIrU/eBlEwuctpd4gCcFLvipbEwZ9S0cw1BotZXewRDOxQ6lNVj7
Pak/qgC0Akw8hlUaRSQG2P7b5aNy2WjRQ+75ARSWUvCnqRCnV5XXeL5Q7CpO2bu1
ZLmvwypDofqeBJwVyl9mCn+JME/ElaZ5tNZpYRkr/s/gX9rVnX9KNwVG9PtGAaRM
zGSwxaNEMMcKzy4eNSRF5A5glfQ19vYX3DKZDQx2xNpWetp3aocFd2EhSkxI4Kl6
AhFaImM6D9NbmCsk/Hb85lm6yc2fCihVOyjIJcEYJbcU1u6ZmdFBoPEVkTLg+EnA
Pj93rmHszXiisscSPYr4Nqz/mhnGFAwfxhLGx56zLoJOfcpjNMIEn/I5rkWd8gZB
cqe8qWbgf1FNg0ZbNlNkVGGllU0Npu6Hul2ditZ60RCcKI59iYnuPmeuA5ojxsyM
suPCF24pJdbBImeekLl8bJubOPBvvuUGbQ/IEslLLcTGKI9Zs7C+ZnvqdIB8zG7G
aweGuYOKL+rcfCVKn1YS7YkXghqr/F6pGGPj0af5BqE90MlNwe3CBWF6z1mQRNW+
/xsnxFrCONvxUJGDRt7m/R3uhkbGpEdb71WlwSeUOVydfvG07gp2LZXTQxYOxNxD
vJWUe/e22VN2LD3PC87109B7PRSZzjgFW1+wEv898bMWabjhLXWhpqCkrwIbi02d
3CFOrWGYvLvroJWXS3Kiy7ebWVHRimqdiqBuCsR4c3mDqYRA6VtoR0GJ0hT38cmZ
gSPgE5vvXPND4qXsnAAh+JVWSjNxTL/WcIS6Xw0EKnTf45mzw0kH7TqGxuEIQRvN
1rR1DZkHnJTeSVMJ4lCr+QT2PJFxC0W09mR4Xqy+jrvirZ0K68AZoKC9KilZsVyN
Jp+aLcfU4Kex9q/7grtg+9FvRoIIu6lihx3+hRDf5kB0txZYFOB9t0WS09B67yN0
E1IqQyezDKyb5ugwqjr8r+9t5u7cc93PrEy4ISkSIQIdH3Xn4OasVu6H8SHAM04e
+jWfgBQUgQ+AgX2P//8TBhWm/N0qHouOQBDFlxdfe9NNJS5peCOymnK8RUSBRX0+
ztZLPq9YHSRTUJh5a/Twmo9RDPuu5ROAAkDZkur08ANrKJTp/MYLBV7Gvgpr5fyH
NSsLOJ8DsXpy0uN1dwu14GIZhdGfAtDX9WQUH4XVOlTFSiBi6bGGf9OenO5O+xNS
xAcnhK80quA4QucRBgxb/zXPQ1tEo4RvTIzIv/Zr5l/Q5Gy+8wCf4pEe3JlNA2IG
Enem7CD76fANQETiExw42H9rtVOKHo9A45EJ4Yw0Ec7aJV6IhPRPzm5iMU5oA2Lh
N+VKIv0fevAtKDmvGBnmGxQ4B+J8fsHj3ZoJ2He96l5PLHSXykAiB+W8ZueYDf0Q
EgPC51xO1VmaTyArMCxucswDdeyrFtfOBTYESjcWZC5TWMPMzCyHHuKOavBhfKWl
35Oz8rwH8H7z5Nh/5nuWLnUDerQaEr12pDS7oz0t3gNdLJZURrtcWCmv8WbMrjSx
rW+Z8r/hysuZ6+IVkkFLxT7pVoQ9Hu9i/yrL118iqTnejWChVb3jj4iK0iXuJ2XO
Il46dlaDWzEQ67lU6yWgaQjjqdKkj7Dft5JF9LqMPAT42h+gH2BGUOs5d3fug5w8
jwI7Q/0TJ/a1KJxTcow47zHf5MuWHYzgUhzBwqjYoj/DZDhNCBk7Fu+QcA8+z2jz
wEI2YrUGVT6jrqLFWIzDsuAGynVY1q7qXFZRpPbrd5f6bhudXq7q/dcuBc5HFjLu
rFI7Ro3PnjvmGffwNkiLZ0r6ccv2qhjoFkbMcxa0QA6pXuXTJyGJ8hQf1t0/VreH
Qac71q6YVj2Wmo6QJutrXnzjrl5+UguO/H7cYeswcXxq1gUNoJ43lKk/ZsQGH0CP
PetQzlALHSyk0V5DHR3useJSNrws10s++/PeT0pgDUHUB1SnJl5eZfBc9y4f03wq
8MrJ2kHvJ1DpCiiM/5FFIY1aR7Zcy/mdDPwHAn97O5rCR/SqnZfDQFNylR4BhF8x
uGXVN9XVUJossI3j7Sz2eiWYb0EseC0En9SJVbp1QX9gxiH4MWm8sP9CIduoUbVu
isTYUgny7UANcDva+u46IeNJTNQ1SJ44nRLH6fbnuJ/RuDnZWaks8NVIjtZbYEsY
n0MMwPWix9M9j/0Qsxw4MU8u0uTGbxgyUgJIfhyZjjWFwIsuD4z+4mGl2OD1icJC
XaXFh+Opil3m3jAnbpUi5qeNaFgMUufc4z9s84fVLrAGfdI/9mYAK1Y+NTJ2f18Y
nL4p9Ly1nre6bwO/Qm1Y6rZy4j/56HvUP1vuQAeLMN2ZNymDQIequ+tbIGtvus43
4ZT/ukfkEjG6x5siRfevkVlgv4rBxzt4+WftNR6hB9tg4WgIaSqFg8OgRdZoDNXk
ABUbVljLfksdJiomB62mWOqsEFd8V1mes57NTyp7Zi5WacSGRXHsOMV/9XgA0rK2
WL+C6mALpUkkcK7lAynIBmDQlPdj0PfAAcL3x6WDBYCT5DgPRnd47Ouw51UKVGdl
Ojtq6exHqv/vkrRZuSsBJWZ4dKftBsQ0SFKZjmn7WlNc3U5MgFvsl8VyvVGDOzse
sQ2qtAs6w2ExREFSMrCQS1F7XDKdwuqYYE2visQSR751c1DpLXbGgKfS1UBnd9GK
UCnZop/wdEYaQZ3Dcr0cCLRIpQWijgdbbDwQ8mSdG5DjIfxo0KjIfgQ64OuWIxnW
crMrvNBKPRklbxULOanuIJKMHsfl1VpBNLVveUkXIdo0YuxQRQBKXNSXZMnErigd
k41OMBcvDMezNFZDr+otVPc0PGcADzD2x8EPuDx5GrP8rfX4dRdmRNStE0l46RaS
yzAKhrNVKQ9V1utn0TJ2EubVN85wsUXkbRpHRfIJ7DugsydH7vSxN5LQSryVee5E
5TDAco/Pm/NQHhi6nMLSFY4N+t0q6QMGiz7WbBmU4MTkIUOVbcRtVayiGd7LlnTl
0wFq5JJ2vjh6Bgmd8K+MOGRBqlQFeVhKVEbhmWOVXp6O2UDW9hAxs80T4ozTOkDV
4/wkORD5D1Uttrmh+iqr7tBNKDIZQhzogl5G6Y9iyPheikrfk/hzFhtQNzbS36Qc
mPhQ86xG/z5gOPDY+6qq8U7BOat7HUrFOsARTBH6Pv1FZGq1jD03qkIDSceZQRoH
VljbIOiMWRS1SptXzIKZE+GxenSU1NusqAg+GbqBLAyrNHw6RdUpvtaAgAjOIpAn
4h1flTegXqY+j1qPG70SyHRjA5g4o8BUxIruUZlkTVJ+wX+bIH3r+IGJt3xhK4pI
gLJdzOgnJUHUWNjXjgDSOl2+whYA6/yiDZjP1dfFUQLiExID8EAeiefVoO0akBg2
3yMJhxUPCN7srmWxLpVA4aHDxji0CnqAjDrnbh+CnimdCv701A01sVEP3tNAj4YY
v3mJNCYARXIsGvVDqaD44ZUqKnuAXPbiW7moqyaxwzKk0mbLTKuS5k7QMb2cd1Rh
yG+M4mlyJE3BoK70+Yjuqb7vlLrjQF9aF+oBp6LAhUAd8evDmL0DRilKsuaFIMUI
TQoBAzcjOhZT6Ym5Xq7vMkCXJ4OKvaiErvENDV3ttC4JlYyjQiSdvGwSUxZcqbUh
BAoDIntkWzFc1urmAVwK7r8wHazdBRdadjnheI3WJ7eebOSO/zpHYfC2QoZUZ6n7
EyQM/sWS/Sdacc+GT1z5Hi4kHirIRR67fNQdIEXc5K8CznTP/PgG+efVlJWox31I
yiOXMbnkqVBP45g6wBUHdAUU0J3L44p0S4tg0q8xANwhD/2K9Y96vhSZHXauqqco
csfJ7aWW2VIMULzUkXPIFWoYjLWTwgft3C0zkSirdMPj2Ehcd33kRnxErtuv3pp4
dnfLRuPwvRhc2JzidX/1AuAitCCuTUlVbYgCjoY6ISl8ZuyNsgLmKlIlwNdF1DWE
D4NTpDWg9kyEra4QwzxMa5narYjwd9UqiA41xPArdlaKxb8qCv9ajpnkOM2t2dfP
UuobdeMHdLzV7mIWBRKKaatIGY8vrcTUweqt+2Uzkqk9f+OVeZcRpwgydf1kBHLx
Fv/U3jv4COdRKeEFJEZ3z+CtAVBYERzJq22+seFWD6X22fC1VEYRpUFnU9T2dlLr
rSoSql8M4GRfwlnhBOiL92M/VOpdY0dLUhFK6d55yh3Sos8uphKUujuVC3sJsStk
mSqPzAj0htL2vhDTr1DnTztk1fbNKoIwRcNUhdk4+0x0F8GhV7jQ1txxSLeJaXSa
FjRf0HiWWneQ9hjkxKnbMbLYOQTVP/5QXQeHqlY1gOmmiagzRFDF/ToaVGMqiOX2
N+qxeiNalnzX5rljGuHWCitOEA8uuGxLeHTsiR0XHsNyXlZEq/4HaEps46C9QJRG
2XylUcTK1RkczQrjk6m6j/1q/c3SXDXByBRiHWeC1qyzZjgVZVS/qYU17FGEtJQI
SwMXsHLu1nMvp0Daol9theqB/9cNMq3MK6pDwHR4ZJ0Fqkx9XNg9FLU6WjERqT4L
nUV+uZ7Q6I45iOzwwM5Lk0tjb5RSVikpmoELswAmg25Qsw59kH7F5sQUTISTbp/d
a3aZHS3k70ykzdw/so0e5ehFlKMhp/4DDXZYKcAWzXb1GK0cWGAy4eL6XIOXMXtM
leLzCPO1ib7cObzDEWynMfYgDK5GgpNFBiCGt+L6y9flgsf7fznNrfguN/2vnWy7
5Iw7MQ39XH2OWE41xU9pPoQW8BwPzJSIYuAHoSeHF28lNLjJ8Nybqeo9byu3elcr
0APXmDOKYZMDIIPDG8mfi/MKDBskIha8nZKqVwFZ4u7U0TUv8AvM2ZeJX8Pe1rt/
sWzvJ1TohmzfnvJE4jEbS4YaBGsfhD76XnHz4Q4pXCTN8i7WqTZOrgXDthTbdKEM
1gNR7zh11JQo2uLfImByztAuHU7+WkCjB5hz2DXSQ1ebbOQeRjMb+XYDljOH9JKp
qMyNfyGXBRfKhaEme3ZV/DVE+9NC73nKag6AbHZZY6w0MtXOvknAuUy3ksHNq+fS
Ef0+OQbu7ognGm5ewIOvVlB+GTuO4/e6AZ3sciF/XMfYCOTP1U7MDb5gXei9apza
Lh/uZfiGpOT8mCXLnVyu9EeRmTuzJlK0d6bkaquUiesUCCqoNUJL8r5Z0t91IjTZ
Fghj1jRNTClfr0p17e7JTJ+j8V0NzOYv2PduJsuH7TqDfZKMoJTCPBTP+8V6kAOp
XAf2bDpTHbCLHJdLcGtiIeEHZeVOH44GrfwraPWd8qgXOg7OP6OmIQ8N3OEFcBOM
mQ05hWTo9Of/MIPpwGE2RK3KKjejvdLEYMMo0zerv+qxpW0+P4kd2koSE9xDDk1K
YliVVrtZULgszWxOhUFuv9yaBje2XVEUZ6iuO6kSuJiUBDmXoqvu+1rksWy/TkGt
+jdLDTjslraNzLrgxhEnPoiWBlksbJkq/3PPLF5A3bU/lJ3pQ5TOyu5z9lVVaG6Q
QKfvqci/qReDJ4Jl8bftnMzH/0sbE1RyRxqjPcBONJ6Jii+snpk+C5sy1nw32O5n
rLPcadktFXg70AbvwSqpJbsTxO4Zd2+USur1Mmr8bprIHhg6jhKM+rOLHC6TTjld
zroq0hrXkQ8NofwkFGQJc/IRgpKLcQHZ1Z4x/crCKXVSVuxk0Mb69RSbk+w2Y8j6
PGFQSOH1TiawPc/u55fWOWU2NYE6BxbbdhDfhowRitv2KLrpA40RNEcfLm/Rqqje
OiNsEVwBuWrslcXtLly1QHtND6etm3SPAKiF/8Qvu9UUT/N6FkeF98sNTFeNlM+A
Jp3jSuFhUqsDedRle8TVbHkqKdpenSGOchT3VSOYAGPa6jFLvHAB+vuYY5fuoNKP
t9+8c3igF8cliZYoOVp1n41u7/DxN15H3l9zRy6NpBqXdYop3RFuVTrRLKGi4BVO
2K8621AAN6g5C4lAq7egkpos06pja1+dyCDAvElW8suCFrwuB2ecu2Xty2+4EPXe
ZoCFXqbIGpqcyajh6MYgW4esjJH/7BPMz/3W26Zweg/L1AqFpEuaXmOrAuPBLv/t
R+yI5pnGbJzRQwHEiq11pWcZfhfK/yz7hRh9pCgicRudDRmBzbg077CriGxjNdhh
Bmym3lkd2iDmsiqe5mqYqihUQdFhkgppButo7dZ/lBjE1MyNs7I8PVTesltt25VC
e608+1MNmptV86covOiAwCm8c6psN8ACuYUg0de4qaTFvZWrirOnHHHSbB5opH68
t16/DjEl3xXfE7r+KjzYfsAN7nTB8k4UvFqQIErY7pB62YrnQiH1fb1lx4PcJzza
IYmWele+kf2hn+fLOmzFWALzQw+MfwN1TPnGpgmOoEAe6oxuuIGs9LcQ/hLbx7DB
/PeG1FXBP3SJoQNeWw56ggOONmn14cuN/Dv5AK1+JegmPdggFNBhefYDiTec55rJ
Vvsa/bRxOP9Aj07X+y2ccltzmCMtJvdXHWd8dpeJgHODLiyGoQKxN4BTMNmbvGMX
zzEeTn5n5oPzqnv/pBfTXOf0I/sbALtLFVsgAImXFOP+1CqsGC09W3eTdYpkDFTh
UBM1pQ/cltTR9AhOe1xUhbtUj3a8GeGUlp7DOZVsR4qqLPPhJUuAV5FYvcWvrusd
I/IqLujFiXJ535Azg/Ki5LflQoTlvfmPJ9is3UVpSdLH3XoM7/scLZe7d24uXgGw
x2LvvbkMHFpFrj9l+hIR4/k6VdyowddI7RzkhP1O1NKjn79agGWAIDtev1Q6FurK
8EHU8oaC7ljXiW94XzqF8ZtEnMlpfjAk++gl4llYNQ2Lsfp6FATPasizD5HEx24W
//fgfJcfDnzHrpKjq7lBeFsEd49Nl7tpOHWnXBRgRsaWYbCVpoTtylx6PKKKD5V/
ludI+UpjYOMIqJXiDxoXzaA7xmzVJVlyn+ijSJzc+c1hQwQtOQ0DKbL5FwML/q7c
dD9ewymb4B5Mj9chBuKexWjVVFguMiXqzZM212v3XEknGLzYIUmLYdtguOC1L6/b
/SX0cVqfzhyUkQGF9ATp10B9bcu3fh0LuoT1fECGPE7Sddt68kYDtmS5LwfN/U+n
Yin5xwZOgXY84DkIcaoJVE+zu35cEVuAE4IuiqmBaUF+/ApHeTeWuLHMyETM5/6N
GSSHgGvgT3EXHAaL8D9EexxYJCRfdHTh/ep0Bh4P6Xu8xXl7AMYYnSgDKkxHDtXv
C8pOqZA2h2nIO2CfBURdmt9+dW3Fp9HoM4GZZFdTje0PZqjfz2ZghJ0/VDnuYzK7
4lEWgoGgTY1EwbMXiEdHui8WJnfcqo5LQ/sxHh/9FLJ10Lay0SIIB4Iud3qrIv53
lJUBiyEU5KukDrjlG9srdNjIaLlzpBdmfUKK7HiQBSAyZXXVw/TGDavp/Q58m+Ar
ytxvVxyzIqEcbY62x14dSs/nTpgMwYAIgfAi5QKIM0C9yY2gMCoj7iIraviCEpmq
IW4sQjb5aM+XsBmBFeWy9nNV2JysKYJbx8paJQlroQSVi7NbvGfw40uX+hTb/ErK
3nwtVPqYnKL722iSjVeRC6mlPKd036MzEOppHgUNrvRNpE6WEY7xFVauIJrIcjJC
qmLpThiG1SLXjLK4aNqnnVYOuSDekr58r2OWyJIpM+eI50s4fcXoPj1nCp76E1jG
+xvo+pmU67jrhgRHKnMjgEub5+7vJtpp0om/QU+5DDE/NltmBozAVdTq6uWwTAKQ
qOrRRAS7iAzCDKk2TjnQbQF5XbmkBTjsRycs72XaY5CHBvebuvcaniPA5LsTb53y
usu/0UlfPQkc4AkEOq0vIXah9BczYutCLn4U5W3TtC34LZ8c6B/doe7LOLCyFVfF
2YQbdac8RkR1ua4c1vmmNL8nP4vLU6MLbmigHOhyb4q2nsiJEuo2bsG9dCwSusuE
LvS3JdSLtVRv3cDc19lEhyNFFGQrX7xlHrdRb6afxtwXvcEUYHIG5DznL8aoQqyA
K1cHZoETukYQgF8wdBSDc3mWTxDk9eZJAcAUMwhMhg0tICzR29f4hzJLH2NcJnAc
evFZUTseSxd59E6JI44lzRqIC/o42+zG5dMmrHc9rvAjXijZ2Q94jyGpwLntmXH8
DD+yvS7YVV4dxcBAY6wqUk+7grkTgOvpDesIPZsXMDgrsOs73JIV/ad3CCtlMNVE
MyRvfRvxzCjRlYyNCBdWx4Tdqsp/jhawHIhEHY7imqM0E2/9fcARVbJORFtcmoA4
ZNOhPx/iPG5J++CFU4keNoPLKsVsI+JnirJ7zwEIoilP6ZkCgQvnxw5YlUrzcdG7
X8X/hiLr3jWW6/VzMLf6R+d6DjpFAerFa1PUwv1LGf5l7dPDTxuA5WXYvTKI0J9k
tN4SYvvZpcfPdycNigpJurLiz4swiif4aNnQWOBhsdeTxTKEcPe5KFphH4gXxD++
E7Nio7aV0903Fl0NRZNWXgIkgW5FyyCH1iFUd9VUg3stWxH0TaxDIuRoHELspGd7
jNBj4+lcTC/32E8lKP5EzVokqABXrECCHygb9xGBX5bP2St3lZ0KKDJrK1BuL4Rq
B5Oq1xY+pP3iYlptM6RlOSMvhU5WIt/KkJ8pGVhWKm7wWJeQQ7kRDkRtiHbjkKbR
Br76Z7J+u191JacqiiVX5h3TmmPMAMLTv7xr38vmPt4Te/wmCia02VnZOL367Wvm
MCuo3Rsdpb8EbvD27BijdBBsJWXzSuCjIIJRHrvPYp1C/j6hOGEbUAZwfSLzTXLS
66b7n2j66O9cXA1tWKsf6XJgJEdhfG+ESPPe4TugNKwXxC2uVZhR5EpMJNrlqifT
6i4Jwm9c1N67LhzZUWavazHHHS84sqlzkiQQc2+vouRJ+/0Wb/57lA4F8A9JeQob
IaPQ8MiiHDf1NXgwspU83HUMzHqtlsjUlsYCMo8dFn5iQ/lwjuaY3ixQMXOkYbRz
AYg/yNWbV3HhrNsPCQV+dGhyLnp8jUtsRic5Sb+v9iaLnGubVFM8g/5vBGTC0BcS
LSqdwHkLFj4bO4XdZ9Kzf6uP1szalJfBGSr6DW/Hk9F83uSl1RgirZ4v+q10CEgB
DtFkhtMJYfLKfG9ztjlpcLjTjyfFI2ntEMflrQDL0mPLuRfQRKeNipqVTXYveSHY
lTsXLkY4fEo3acSeraiLtPAQgFponaWb8kxJayU/ylJg/mMrfheFb6HQ3hcRUC+g
rE8DzdQvcUuK2HIHKT1JmlDi4nX2ShQhSHkz3jMapYX96ZRLKZ8HoMd1ikz0YyA8
cwb6cN4zojsBrpOh2Jq0Lq+Fp68AOH+xXyGPyk0GZiKfmdr/2oWowxKRHgYSRkpw
msFB0JWQG/v0yh6iIe5pdXG9UnDisQ5m643jqeHlH3qE+oJI6elg1rZdnOIfXR+S
lmHG1N0UzWOS2vSowAWINHIyW0UP9Jw8xYIBP0rHQQM/E8OEiSTAIIJnL1cwJFFQ
KDfJzOLgCUH7PqhLKmO+JjvmncGT4rzpCvgTXVvDtcTbUUnYFJHleONihOFNVzBc
L6KLN/FK0cTFEFFZvRFCytQvpVKONpFhVJmhWQM4dIAnG0/7uNPcctWf4lpf2jWM
LJL4Ne0F7PZ22XGPimnu4D5ClKGOXwxZWxYbhJl8+Ju/h3GLo/GCX6cs6unNdWaL
OdYsL9MC+yhvSdlySbEnSLxhrScYzIdHG2nAWTBHvj3r6HkHdrWxU9MqDG6Lemz8
3XZzO60gFln9HJXbjKyUoibchP1DfhLXruROS1UIabW8A85OVgEb0a9af0PspUM5
ArvQf0r8YkV4IHgIwrpo02UgSSf3d/xHyyfhC4MQng7RD7gub/SepprZbhdygerg
eOp0sxl2uNIGZXchfvQCBCbSgzEBpSfupIoQV8k9Ii/wf2DD1veeMvCqjYnxqieU
SweKdjsmRES93/ObbrsuQCO71c24N05Ia8DPuyAo2vSl7znpsySTOm3J8w+eJlfE
RPRTSlf3s7fbq9n0IhO/WjVq5A7AvvgWrNR9SJ2FMlMqAaMaaXZW1Z6OkCN8TFUE
E+vFpIo7LFgsYZpMhwo2mos4k3fXbtzPSnfKHe51LGIANN/HTU8gtYJiQEa6ymNk
Ar80n3CHLUAsyicYEEvtXrSjtvliZdTNjxhRopSaqEqbt8fX0Nhfx7pasr5GxNUr
pLCFVDEKytspSjcYKHLjSJXrc8QjL/ZTFWXaLICbNQet0Kz94c6yPwMBWQkr8XwL
aygmjwbJt/rjT+1d2PkT9TSr1rFp4WZrpRxBMuKf5O4FsgMzdK84lJ0ioSSBhF3h
rvAJS3mmFUOwThsOBE0vcsdUg0fX7DJRfgc7DDwLCDZQm9vQE3C5YOk9ZR1FgsTq
Yu0GrrbCJx1w52744l0L8DkFSHbTtXsy5YmA+gsmH2yoDaGGzSTAjy1HrkjgyBc7
p9eg3zrn8w497ZTS9VdnwlPscbWtQHkVPY0LZnDhsv6bCVDsr9QIxhQBV/3U5eoW
D+SJ2FlrbaaU9SGC5LhnZtQTUFtMQjCWkT6IzusoR2AmaV4O4qMMQ8WxHQLVCF4/
36cN0ureXv0F4OX8irD9oDRDlQlywl1kYbtKUw+/xKp8CYEPftYU1SnnnaESwiBp
AgdqKaMddVZ+v4lkfoPAwzLs9X2ELfWIm9c8sbOBEw0eQD44BiaBH1rb1AsU1NzU
dzFKJIUt0XdkLguW3RLD7HwbDoOn3wdGEBSizjIX0SZX2SUson/tPLl2U5Npnlkh
4gO57z9C5P69eKKDArh8kyzwqzZLWd+Oh9f5LJG9Fr/B6153UcviYkNH3xQXR3Nk
TrFlS3E9D7qvYHZSt1QGbYV9XsD7T0TsXfSKBp7iIKx09ZgduxdMFhn31+iiSxTw
nmsJMFXq+CdBzyE8apWtQ2/Q7DY9G8dva0VA1hostxVvDREjYJaDdz74OvsA+h26
Ypu4rXGzxF/b2nTbJrX/EMoAVsVLJypnArSaV5zkLc+01wbP/YZ3Q0l9mkOHCthY
EbdNPineaMnlqgzHyw5lzmknG4PAlfz37bzPAMLMTz8cmZJrePQlLVrrFdcEzToB
NFoPN0OQ2RuHwqipa7BQJei1TEmbMgzSMcpOgaYxLuwlnBQ4Nl57gyeRJPt5TesC
GZQ+ekzdPTMI2oiLUBTFGzyW8Rs/A8L3jj1udMMr6nEKLoB8KARIr0rvMqYJHDsx
Hf/feCwLqYg6r4KvoSh0WCWTgOBfrFZfOvIMpdD0mlaY4upzLsWWUjmHEJ6KPOuR
V9yupsVkbdX8skUy2z1vIqvEy27TqdtywJLxjB4lL5yyWSCS1MRPdBADCOFxMgb+
6+7HRoYaezBfB/6oVsuIe0lsvGhc5Fo6em9wJ1O8aZdKzzze84L4gpWiq3LpYRku
jphh7yATdjhTrJdTgqPe7v2+Urhnhw3YtFWwyTRyFnU535nkSzB44/50S/TH3WQK
I1EI8O30iOMzEhmGVNu7S9b4yOgq8XWmFHKSXvIsl8ZtS5c9bKFpCaa5pvEtYzML
KYL7TRkqsAquOMB5gsP+z75MpD0nJWmGPhJYt8S+q/eGRCLZ4rMLycL595/53SQ3
pn2wEaBcK94Yq52pXIo1kMap/YOkH79YhKC7Hc8EhmWPqTq59B1hebxk26CwHRA0
gIwjdqvLiGLYDG2u45TalVK89kPmOXqC6EqyDYo7II+1rQvAyHVcBYs66o4mBr+W
5S7E5BB2jajtJ8e0gx/mOU3ZBqxjMvZpgfQOJ900+6TpK7cP82p5zr+RQutUKJmb
3R3XL2w8Y6UT4Uk+8hQiMj10asP8A5f7pq2MbbvuKGw/ext/7H+GMdGzoTbiU08B
mhgjVR3BBQ1KzgYCoTMHW3KWS5eH0AfpLiwC2g7+ZKgKXLLIS7jCjSCgj2tuVH6G
Bga6xE5F1PiK/DKyx6IFZhz9OatvXNSWDm6TqsZKtGF43KBUJuR6nV6oTfj0hIgh
UMqV9D9KULU2Ls++shRNr0V07eFZZBOVP+phB8UiVz7D2w7jVz9pLugxxr/Ywt9S
m1jwgZktN8udjpBHQGPCGkyirFMT+7VrD+fedElXGh+2atzFS/I4JSLCq1U0TF9a
QSBxlxpTsKCvYTSsSQAWVTASTLODCjP2hu5LkO3pzn5a7mQaKMFdclYYoaGfRem5
/Iu6ZSBPt+hlh4OIaB/M2SDAcXnXt6CU+IRPy9Rx1bAk7BwLfsnEknUbu2eKlazb
926I5dVJxOxzp7xGGHO9pSQ73bVLp/PM/RqlbnofzPwbUg6K2CHLojiLoWb+cmFk
mphq2HQE7tjaOwKy8m3XLK3yhuEugbmxywJBH9PjKwm9sfXn1N4cHjfx1dYJRahh
7d2s+aBKNkbRaaDHgodyTjcIZvaPrJLv1Ame+r6succ5lSCDl7m3DbKkXR0WcKN/
w3acV+OSDm7x1tEr3hts4x1CkFPTc7O38REQOojIIw/lBA+RXwI8cf89Fo2swHd7
wzlGE0PiQ22mvj0Rpwx+sHtGb4u4jYoqNjmuZ9awxm6mMZgo/A4FvHxiQPcg4Bwu
N4bUsaAVQxlDJtycHn+Lu8w7KI0YJI6NBdcB4DvpPKAnVvkz6JNylfjN/aiNbj/2
/5NwucCRJCTsToa2jAaG88+UfzmPSRo/mFAOMQr1QWuDCR6hmqk0p8mgE4MJkXFx
bV7WFXuBxdGj75pUPFsOw3L6V6Jk6JgISzPY+m++vPMk/T6ktOeaivXiAx9QC95G
AmUnqPNEzg8hP5cbx+N9tv0E8vH2DJZ8S4Ls6+R5ceo+nsmcxrJAfLNFw6OnNjEy
59UPURbYWkqNXCYAdE1fUIhrJR5tPR0GuYpoVq7Mb5+IkE/nxb07IxVkk3Ad8/sA
Mht6OvTeJYSJPnhJ93tPP23JBMuat1n4VPs7YNy8Fovdo4NmlXBef7PgKiGj62YG
C3njJwo6xWhBXHUlcn4DWOf/veJc2nVBM1+Apm/RsPbpqJM9facyYVrPz9nDNFY4
nqTmqyOo10OYuj/TPqkVhnbMdsIwRkDNJ0BJUDv0T3nwm/w7gIlI/o+shn+iw8n5
uEZTzz46DrLesUQNiSQIODSS93Fhh7Oloi+qofF9VeGMe+6JGjUB5MfIY/4uIS32
GdyXQOwYfSMFVGKPDSQ6WWwQIXQw0txkCQgnkVWgfQSY2jBGCkq6OV1+OSUQbiPk
KOLurPKufQ+wiSbZBc09YxolS+JcCkw6OYWfJ4H6HF6fJZ18qCY43+4Z1ov2fBZd
a5fo0pipMmhcagWeR3tHsEoEVvhyHJDoKqckKJK1qwMGr+tZWUx4U91SCuGIeqfO
TsVzSn0v9qvjMQFAP2BEEb9omlBMxcfJs64hSbbDdO4MuFQyBGB/q5sygx2kQ/Fs
o/daAVZM3k7z+I6pTEVWJljErO56VDpT0oRp8/hRZBGrneXd6wX7NvOj64t/j9bb
MuLQGT3QCN9ShP1+syM7aI1ovIYy4BV4tvkoIdcmOATrHCaTJXEP+fFfSa246AxI
HT/FNKbD72rORbmnDIaBVyzPCY/yKNOFMR/NpjLRubt6DcG6FZ/eqB74TQ7lVScm
9wBsiJaR7y9PaUK26IYZ0JU1l0gRODrgX+QcrqLUBYC0cCktJqIuKLlBcFgzvwKz
DZF8LcEtMahVtXThvPnaH+Jhi423tknjN8qEg4hnc2/FkCdMmV1Cwf6XX3nfQ786
ZuqDNeo0YjPuHnkDoejai4NSpQcC3tdng6EB6w9pecEgUDeqNGnnfPvtZhTFZzLV
ejMM/8xAsJWu2+bOxEq9O0+1fBvlSkzCWg01czXx5SL56Iga5Xxq+d8VmcOSuukZ
qi6vG6P+FJPs0rE6bk9RW7wKlwyn2Gwos9LGZxZGEUfjMLTh0QNexrIzWtcmeM3Y
1MvqmaDN/h6YRuFIIxTydEbIwrSmP6AIrFz/SfTGXH/AMZj1RL39T2UVkILQ2HQM
j0ZoDahZSB644aVhPXRN7zkRYKl9cog4hSVHWbF/2GqxOdjsLZEcqPJA7D6xoSUF
3tjjUR5n1uOMenIj9FnQHOoFbBwhbA9gDdrwbzXi8z4NlMQc80bktzx/Jz4e2aY+
JVJSnR2succ+6fLU/gkkQfdYgo+B7PZdI5hVWEQlvAwg5E7SYPzjnkPeByrp8d59
3pz/H/vXw96E7YkcQmJYixXiNkvbHbOzay0T1RgaXTkDNt9PH+pqm+/ZZC4y+5S0
G7Js/1agz1xL1hVvbtmvle2fO1KEaqC1VnjcQezeALSPozzPqSD6t3U/Ik5fYQmV
dodV9a1O+ETRkUIYnpsnXWyqyY8SbvXCNJI/8UwYm/6bTGhbCbhGS+GXDHkkV6YG
Y39+qGL7FtHNWbU//pAlboPHV7291UEn0EVDutJ9VRTLsrMRE596yEwRPiWvsXcx
kqoVjQhys1/sSpVWurdBv7sK8KkHrXD50OLL/nsBdraYFuQ2E9ysTrhQdyJm6PfI
bLpPmD1/A+NPYO6c7NJwwxPMmOlAcOvdcrsWWdvVWI8eRtBnbEpfNJFAjz706jLe
SkdGSF4Pf6NwMRQEZamRyw1puaADkVQmM0QZ5IqNiXt+FzX9X94GwDTnNonKOr0E
n9Uu0Y32UkWOl1qrGzZKj2agd7SyFAY2xrd0b6XtgfYr/eCFdMjOm8AGbPyU4+tg
jRK+VpBw8g+knL7XCMAdbUBPpvv4P4WvjGP+c7zWEcHUw/N4VXYwciUaNVX3aJH6
73oSoU7a7m1fz6l8p43l/s9lBwdemDNEH2HTKNQwtGzeAbcViU1gny+NLjEpXd47
F2EGg6RfY13lOU9Qdi1yc7EhkVYfNtRr6iBoaUlypTSV3hYtzSXC4LVC+KfkzexD
1LK2QPqCBaNdT2QmR0vWLrHoJ1k65AZYKRhBFaETUhaHpHDTQhZEsTv71EHEN0Dm
fJIC4Il6fzdfy9cClEQzbT498FDKB1oVDLD+JHzkMTiWXM8XYQ/ZmLHsnKtZAgBn
FlMleg5c0gEkT39LCxvuftZCmlRVk62HVqzzn2ek+ktkFHz1lEk93OJi65+7hMoM
0UJAdo2yojxi2uH8C+HyUKEOl3uBhZsGngsik/nr8ln8aQyJN3WNXEvU93OOzDBf
50nqQ6SD8VfZ7rGQEzgYzoEvESwgcPeKgGk7NAAnU1NvwAK1otUmBcofWHYtliKA
eU6Ztz9CkhA/NHcI/nDtM055B8FH4meo3VyPoTLwbREevL4ll1bVwn82aIENe7dR
Xuc9ehIFFJkMUAYMvsIQvihmz51WFXA7QUrJEp5aV3rllossfO8+GajqRONdwNm0
+ru2vQSF7rLSCVYfmqoRwfom9pXs8//5LPuGFDW4n9G/DsqQHsWiXO/bWGm5IwJ7
siVwcNtfCMAwioEF5o3dNKdyA1ql8+C/JvkfnSPTTbWeE1XAbTSy2OObMHyFkRa7
41e8gTnu4Fzn5NP8/L9y6VBYdC4zw/itoUEZb10NM0BU7b5UDrmpZjND/UgoZPZO
GvJ1nPAvvAjpWu/JVM7L069oGpyUC7zqAIosCfUhN2tPjNys8D/wj8H9S/dg+9kh
4H6GUoYAnALlqM7YW3SSxf+qX2b5kmXA32rY8sVeQTintcXrfbsL2RzoGmuLRlzw
1U5JG7HPiWezTvy4VvcJ1oOkAE0uWOW2LA9usuWTuN6BY74sl3BRtJTnDNQCJv1v
s6iPJ1NzsP2us+xuYz23nC3P9fTjS3VJAhtooEx4PeqnlxIwAIgZ51vtnZZv1KMk
kX1kB8z4icJnCA0SsITPGJgyyunLq4gmK9OHMh9EkhLH8WFJ8TbRAX5z+qDR72X0
iKYw4UaLmCsI0KzYWtW+WJdexxkoCiLfgKQ80ify/DRD6A41DnVuDbQkUcsdtMYU
IabJ7135MlwjAllktTRZHQ+gXuPrlQV/xdRVJ70hBGXYT4Z5bb9A3LG7y7nGIoZt
fYTWnaXgPQM0yD9w9mZU7QppiSpMgnHHTwfMI0GVk9p7ha4vHFdxLtaBpUYpnXhy
AaNHUrHQjwDGRsbQ4bRv/C1mMh2Z4h2hihKrV8dBpRXaPjStA9xM7PaHB1kPRN2d
CZpmybJyor2g5Vlx/wE2KBQZLbLgjH6lVNIquFYHd9JZQjNt8+iO52YjPCcvLYKN
QA7rnTJ3zgns5T8NShfICf2je4Q5Dr5kGFeMrhb82PJ5aqMVVBpYokZue+uZjtdC
8y1epyBT0PaXWqR+vHLEtln5fEYr0ACXtrcwuUJUlv6+PmGNgLz5C5CX4Kfx9N+H
feZ0wqb82vHwgX42fR3WEn4AR9+39G7Abpm2i+PSFZ0oHP9j+oeE2p1VNALZ3FrH
+39/9THnLPaVt/CIzeWsiRzR7d3Soa5rUxY4qOilyBmyPZR4lmf6KnmUIF+RvSD7
YPNTd4oHGQam57tGiXteIBFWlNadoe9Z8W5tTW9hzcIZ4vlhamYtYXk0aWo4HcNV
1boudTTWbxZ27IkFL9qFOPvFJfYaPnuRLWEQJfnXUyMaKONLhw7W4ehhm0V2xNi6
+AF107rbG4aS1VjoLiMYpsmq0gDZJeoYYejBi647FuIAHMO1rd7xaf78wqfH5ydh
Vis3xfVxy+Hdrihq8DH7Jbglw/PQ97L4LqLdxHRzCGtsq7Jy1yWpK/yRmgoXvA7s
fp44QQdhBGd0nQqzq0ZQGzqTHiSiVCzjkYdiWP6+cMJYzJqT48CK9ZTgCMT7Z8YD
jYkh0w5pdtmoPTMrS5rgyLhNAPPEfJVtnxts4zWl4eaT1mARpxh748BtcZ02Ah+h
6AB5VanYmEK+IITjuNFC3gUWv85JJA/nMQFWaDV18cbJjqdn98njCDskT8qDXif3
hKjDszwrH6JzKbDL1tBLpcCQJXdtYWw7X8hoDPyHDitxYztFrQhYRIZQhDBAp1wu
cLeHy8JLsFXBHLMJKX2nKwlCCgK4gt2kJeJSH2mubHn9t8SYtE0JN5/k9hSSSwqd
VH84s633gfCYpGEHLJ3cLUHGSCowkL50pbtQ499n5XqAmGOuQ6vkrQwhFGlC9OHR
Wdkts3zHbUxnZev+IE3ImvShpRaJPpC4uyaMhnc3T79Gl7YLwIbkX0RZdy62mY3+
OFWzVLlCyLkwaziKpO2DW41Q6lGts7WgYDisYW1YdD0eCPcgYbts1OLSDLR0idTt
SZEvH8rclzPTxsx3jdiwpEM32uRnZzLYB1FF/LVTLily+nr4GZCkRjLbRwiokEbH
31sZNCKQFSN5+ml/94RW4ZqbDMvHgHVU3flds4UsWAAijzLQMJEg+xb6TDBz3DcQ
ycg5UZ5vMF4FgCtiIEok+5dI68UgEDj1HNAAXH0TzPVO+wFc/Of6IOoje4gG0aMt
bXSnV5Q3/YMXOa68oHWsjjFF42jA+UlnerNHR4/0+Xu4lXyK4/AgrRc38xuTiYLa
xna+wC1vb/0Jz9QNp9Z70EtpAq+L7UAHD+7PfwLB7RCVVfrcVGQnl+rPmnbzqWWX
m7nbzd+8l6eoZjWtlpV/d78gSP7IQP9/qBcf7+3TLQTxm5vCSlQHUvpib0Gs5p/W
JaI2mkfilL0DXmXnPLnZAhFbX3KHqp3M4zjgMtJIsoTIE9MSedSPSnIeVPdLy93Y
opUC5DHxdCc/8/YOr2FQbcris569znDmEFd4tJC0q9m8NqcIdl44UsJzhVRpVibq
gSQ8wjK2UzgBkql/QeAeWMm4FNEhFT1HZ0sh88GDQZUXaLL+bj0aEaPyxvWaY1qn
1lD5Dq2UC63CJuEJ4skB1+kM1IE22WHsB84EuvfGX8qKVHA8acmCG2t3OrTJYNUL
Am+27I6rua6bSTSLr5XxriObFDSkVQQtHhffH9RibH7DklHrrDiZn1JjimlooUGU
v+d2O9CiSFkJDRm/zk5lkMJ7L/SjiI1gRTaKWqUVmO7dbMY5CV1bJLkR53CXj3Oy
sCTX+gDwCGqGwycgbdgPNpCWeLZ4k1aYPqp4sWhm2MPSr45lzChLZvGhULJYhd/s
h79ZP5LCr+fquN3HpWQAz+5BXtJt7Gjk7fOkiVlV6/mo9PdZoAeweeRE7/omYYDj
wRKDNG/su9iHrmnkquTq8Zpqepem9qr2uOS8oVZ3c8VNkkBXZCYcuIojWOcQaWeq
Gj4R0s97r9PiA8gdxtnDy/qAw8mZ8djhfNluq3YOTwuFFmtws0BtCmkDPVlkh5IW
kLmMS7FqX/KM1uH+oyuAePsaxD3GShXFswYu895z73XMb3P506z/mFeG059QBFWp
yA7DLWft6V60Ov13Z8iuyAjaAQbeuX0OGF2EAtgV0yxygMV3PvshRhLkPfQx8uDV
e8VaHZPgPDukMV8zYGTJOdp44vRDgzbTySCqmBiTOoIX/be8Mf017st0t84vVzc7
XTYp4A8g5OXsl2olNu9uiCKnPqIwx0u6LCS94erW1atREagoTAJbPkzn19n7ZR04
ba7/Yla4bKD0F0w3ynXV09n7/X3kCdSLhwDiqMwFePnISHgYtm5nu/4pD9zshqps
qdilspiHXkav+NmoXAG4/odp8EUw6k0wIoYA6VG05bE9KdwcRw2fJ2fSSt6a0mnt
GJiNpj/QNkESps+w7MHAcndjLXqj21gt2MrI59+ghGj51JrzFY5cmkt2+/tbyKuf
hnWOcCFAO4uHbbk5Jozm1hGrBIm3zER42yOC8I3n0grO09fGZJWuxM3nbhiMwyOR
3Uhf9b11mOfTujq50u5Tc7IOAp47n/jsbBRUgolVA/htb/2eXdLhLu3jlXIcAp4K
vwB/BNuNDN1UPCOUowHl+1ViSWiNmA53Yk9CT94Ix9shTT5w/9Yw+CCcnXz/5sHU
yPtPqbmhHoajaLw3FIAXfjZmi2DyodssGnIQfUCbdEv5bhz+wKbvJOfJxUhv8rYg
/d5WI35+Lh9S616n8EytmuLBhRAG9StOQlcXKFRb8bT9f5DiFtRsmNTygZVZzMQS
4WkU6dUJffRo85jGWjD7HOA5oMxSlkg+MwlfMnnFAj8BGH5Mw07hPb5Y3trU1iwO
hCgt36NWgVdxFBdMVPipdA+hZyi5wKS9uMdSsfoWe9IEqPMz5TN3xVmqZokJjl68
4vpNdLSvJgmhIEK8LoqH6jN7TfjuZBxhGZBfKjdE0kyTtTu3JCzB1pga4wrp+uOJ
3xZJp0GYAbD/yiy59tINlQ6aC57t3ImtoAbPjzLbNAsGWIIT+O3JqQD6WFgfBfvV
fAB7XrPGOn9TF+c1UJgSC+XTONfFKQanuDW9JcWJ76vOjs64nyCq3J238HUXpHJ1
IXuFDerAtlPla9FIJAsG7cwxic/oms+2BbCo9iS6wV3KPatsVEoZmdn58xzGbmfF
I0+A8W7SFFQyikD86eBZFTZcbuUz5QNIF2EhMyuwr+iiHJgB/MD/yFS7VfA14tB5
S+ZJwQ2xnNIEWbcwpxp1hhL/64VvjVCH69NuESACpYdqxnbk9WC5edwfxVqBnFoN
GU53yYKGaqkKhNMmLeKcyZLzoWkJFbDotFSzTX9x4/GDacEqjGhQKEms/8v4rw8Y
4rA6sYy8/m6wmfWltBZvI6UksSZefQT45bjwZ65jUzkxOgyaHjFmfl1JSOdxJj0w
zTcwfhqLhvDfmulUx6ihLCB88cH1NQjK2w77LqsN4fNAbdTUb8wqsey4zI1Dz14Y
Fxuptd0ar46TMScrxJhtg0XzrXyw1daRejS0Vuea+/IuoFGLKnxwVeVXO4ovxfeO
go3PBu7emagUCDMJ2i5B0z6Mq+qrTBek0bDmp7i8K4Gem2OQhPv15zqqfJaf65dq
ED3eKzP7bMVZb9bVbuLbbRla2qBS+TaVRl09Wy5wpjIhhRsI2ToBjQHt7WcLFaJz
TkSlKzBYQvPcrBy8DdHCROxYVbpEw14UrHrnU1eBXjJLgHR9v5Z2uQl40aM4VuLC
irIr1tkziMr1KE8CFuBADD8Vof6cfzfEZSSVSbZNFus5mWqORh49R2mTtYmBpHdV
/19e72IwP/tWOas2Mq9/R7kmUR0ZiqmB9s+lwAUu3V91O1DIHv204iKjW/lqj7Mn
zE2D2z6AZdwZXuPBSTlRR8+01+V1EvuT5L8sDCo3QAuLvmZUPQdXdVmEtUA0ngjd
IZIy3IomUuQxxl/XisK7nKiS1zWURmU+0d213H9vl9S74oZt1K1PVhv5ravewbPX
LdJShqnHzayeZRqbvuWfMpBhI3GwgFw5L/ineokPp8BWOX/6VfNzzx3kxN3L2mSz
De7C3eM9EQPG6XQ9lUaShYTf/nW/F9Nf20fmZKf749JqTsBP78b3+9qZX+RDmMsm
VRRtbHVlSD8ljGFjRpAYFqBEK6vjJPBfhEabntob5FRTZsPiFmfsRay1AoUUuR68
9pizhsSYj6IFZLLSy2Ev8wFsfGmJo8b6pppZWqV2VVqizvASufU0xJHvbjUM+a3n
3XYG234uV+FbsJ/cDf6eJ/Xvuuo8do4nA7N5XK9EpLYhAFFtPBfy8E3H4GK8LWzo
FLR/9mJDKa99IZpbn3ZJLp5pEn4GvYL7r8+NSuSxxUkGnPb9KV8EFRxfXBHI2t3q
rgeou1kDAKP39Sx5SGNURhg42hmgcMqwpAuifVAsRWmHiScvJXLriTw2G4wDcWJ/
OO07lDGgr5zMO3Zg15/+vtb+5VswFAV173IwEuwmEMSBgttxD0JkJU9alnasUHhP
b+ObVyMBNLredzUfiqHwZOVSAJn+yg6Oc1LrkVzx3pGbj6Z9ViqDhiOsPv9LThjC
/iS3JZ5PrOnRJfw/Kqh8AicQLdwbyhly4ZXjLjNoWxtzdCxhJyGLGBgdDt+/q6tJ
mVF/aNSJHmDMlzkwNFFormqaYvCSH69kEH+JSW6M5OTgjT0o0xZk8leEWSLeAs9O
n8P4fOxc6KTzFWtkNcamA6Z/X0BhGfGnpnwoNPgdY5NF97ZStJTqcloLlpnU+M/Z
HsRKUpI90GX1ynwoc8vLOKtWMCq28rKn/lqknqs83/jLPJimi/1+geHdNH2864Vt
L96W/HvqTGQ1jCmm6mCQDY5izsUpEZCCl6yljIMLF5jZ98w0+jPd6a94PPdCKxOP
y6EcinBO5PFgUazZFUV8A/bi/K+GXuakg+6IT4ALHJ9wUJhgE7rKixSCewoKga5f
EO0HgALa02slvuoun8IjfumXLePutM1qR5FSsyaqJmWkrWVmQ3Yw9YbMszIS3BsU
OSiDiDfskC8/nM+DFvaw7bCjVS4UBTUvqnYaku6LdkOrWghoiJKaHI8FgINo5FLJ
TJkWDk0GGlnDK5OXzD8x+9+io2yl3MIogJgpVHSvTHWaKtJS3SpL/blY8ABQKCBV
z47QstzDhldI1NbYb5O6GPjhregWr3wSno0DZ8BJGLVveuqy7yiUFgnfsHCGtYN5
oSgbIEmaZHrCCbuX/70e6HkvXehX0yuf4vEB9bMy/Xt/fLREZZWuyVwl2P+jU8ax
6b9jiV96SPGy1BamyPv2VCytG4jMFYeH48txH/rXG4S7UraEilW4LXP/OeE7o9sw
n7XEeGj69bbKO5O65KwGo5tQvhpNnimHOQfAs84OXe/WQUHRgz9sH7xKSV0UBu2m
y2EFaMnKD59M9qjM2Uo0gq6tKPhvyGyUHmMC+kKFZUi4VtTKMUnLxdnXGPFn/97B
MLEIFxBu9gKVypK/ZOEO+Q4QRvTfzOkw81fbR0+NzSej+DEgx5aITATfUdxbEyj/
UHzVfOAjwOelOBMjbjsTclBgo5F92jlfwQzX8qXe6mwBetBc3vdzm5EWnXkFvEjM
Pn5xcaainMTqv3Z/TQPvv1YDaEOI8E74gih950psMrA14fCkJAmky0Sw4/nWpuF6
BGc0koDefFGYuNlfyfX1lxSfeXdrocAy+ii7QBBqSn/nh5f72DzWyUnBG5pV1PMx
6zGel+7q6Q4AslEJzzaJlnPiVOZEjdmSMlgNNJ/W/DMy0fKW/W9BUMO5vu1qKkaw
FU9Gx/qMXDkPSzyiWabyBuDckRk6kTJSXP3mLoAN5pGF1X+B+3Dbv5wkzBMJPlU3
/hJX1D93e2djKiNdVViOyeGzJP6n1S7FjsTrLHCQ9+Y9gLLljvps5Oa5tF6EH57z
/nDshsSAS9Y9eB6WFZj1C6Zy9H2+BY/Wr0ZfZgQ3Z1ogEbyqNHt+WrMwEWlsBjcU
9XP43QifuF2mRVpE/IKB2zjfTiEehcccGySYKWxAjEQpjjlqFwnxAH0RBU+xOr8k
mo/EbAZeJAgdZpHUcRYued/EpQo8AI5axPjufLgC8Fx3zNzhNBwt16Y4EO8wXEeE
0ERyoaqqqROBbeI18UORzqk57y8WsR7e1GpRnqaSbXuQjOk/rcu4OPPXpVIRXuEr
9zr8QNYSt6nEOMjXrrZ6q1ZATi9S5soG9lqcBN5KhKXQ3ZHKSEe+bIvW5EjsabOL
OdD0DDv5mHPyBa7atgJhKT609rPH2txI0kAj5G6agItppF5OXK54XmeTODsKwLzm
JsRdAneiNSThxwj9rAZGWYQ3LSB+PHLSp4mPGh3r+fjS1AW22Uswqda1Yqw4zIq/
KQQCaBl5Qi/8yCJHCI8Of+zj0zz0AKMGfCVNdN4VtjLSMe1h/y8nOwXPQYmfRVq2
u/7dXXPuwSx33ms3057R/ZRDYB/TDcPtFsLcsIUZRWv9dsCvvky7iRKLLpT6tFnh
LShRKwoeOJobrLMYU3oEqEOszHR5PfO9vG26SbyqVeyHlbCXcNU9y+MV+LyGVajU
Rl3rMA5PShqi69a9jjyVqYSnOsFbLNEfpiEB+seel2AZnb/UmF2eGE7CyCTjwpGf
XDAgIIy+R7qOuppL9vS7qdsiC7VUtVD5YPpj0IzhQFhjJvwkUVUJAz8dVok04wYB
+crX/HQoEXohpWFwHOah03SpIOxW06RYeLKjx+owlxkrml+DHhwEOiD7vhfK6pmq
/w9TlpqjVCz0m/Go3j6h6KZak3arufasVVN4fD/SooFOm7RWbuLcdWijO8TL9MC/
TgqbgnifPhStO+w7L4KgQfCU+6NTdD0yC80Lhcv54QyPtjSobkKGD3pveMo5qROH
JrjckfTF02dvmOGOoD4YUlxAWrijiQx2+U6fSHEadfAaqHrGIWMtE+iaaYrkOiT0
2qMjkXX98GRAcy0CpbTy1s/hcvzFVZ40BlDVsEGMOM2ysexpJ6byw7K4WiM/3tiF
YDl9M8B1M3OmJsLPaN4nXog5KRjy+Cavry6WxUqeWrDYEjTPMroqbR8i5OzsLTMT
dLirQPNosk1tAa/boIzrkK9cVEBIwsLo2sKvn/NG/Grii39Gj7sfDJVG4HKPdgGm
zqGcLeiAGL5UIDAr2wazP4Nqm9iB49/+cw0GaoPJykmCCScpAHkfxlCFYBLDnH6l
3HZtAo0WQV+MSomxoCjIqxMyZtfRybGE/iGJcNARHvk5MEyIKuNar67gtYoptAnm
qaKH/9WLHNBSLW3gVc8MqngH5TsZYsSguGKOquZpYWXAhez/LtWfiz86mejiXaPz
p025Y6HkWqOJdqHMm9UzAuO3i4jyhG8I3vAJSptm1RruxdYmeGVzn2ekYRXknh2K
/TRp4Kz3JGl+XIxLEDIg4mRTO3loTDhihvV0karU2WCI0owM3+dcepdGVKCBCHQ+
0xRUqVkT4gdAkMbFHJomNKsvNojueNYXiOtDNQyiVnOT65CETKu+cx1C/LJVKeNJ
ZbKhHDoF4HWFd/SyEU7jiJzukPZbzTrPITkKaaovn2KrdnTcdt0YcMw9NoKuakmf
+Ef8sO6+VFdRoltoj5PmPZsyazdCVYCGssnODZhUSAXb9IYRjaK+pnhUlyy67xAa
874Xtvq1imhSLeQfxP1d6+N2SeI/n6WJskuSrwNCnlP7lUsjyfZ+to0yj0t0LLhY
AotbwNnfmXBXQHimcgepbk4vWJXgTLg4feGroZHEqpNk1AzHSzQoaZ9KFg/YbGYd
CBG1Tozx9/PKTwycgnvSNwowTvStCFehkOqvvF4GHCpgKAtdqtw6i5ef4NhXq23p
SmVg5ESt7jUy84+O6UCc/mz1IWo7CzbprB6syCJD7GuiXqukqTSjloWWgAZhlSpZ
z8qqdTPELuA/OVGBItW1zYMhZo9NKS2NTyvtEHtzwbPQcaTW0OMSO7mSmBy3TBBq
GwCZ93OtuepLejDk/a66JWDj2p1vlMQlplcW96wTniLW3oq/eyeSTcqrjhYu4hvG
06XZd8tBoG80gTwuCq7sPlMvHHKbOWXeo5Byaa//7ytLcs2iVaDLOSqAk6hSOvmH
tc8nzrZfMvKqXP61BgWX1nTDtpJLbE6Xj0XaBva7E+UVvOyoOl5+KdHXS/Xtgman
lzy3NqEDypzp5JDBav+ojRTg3d5tSRxDPbDJHgsa1zqleSOqpg9/XHZy99T7qhy5
jc9kBgQYRlb3UyniIh426mwgLgJQLrpD64IiDAQmPdGZOcWqj85VAfcoAtbC6U0C
yidfec3RRkSWzYg7LW+1oA/1Dwb3h3fU6ECOege2itRHE79BFuBROrjes+Rj2gng
9IOZnKzTQuZMMzLY+iw8oiJLANG1+h2yb/+XLSQAXdebNdk0wIGS69GeSmRy8Uzl
mrsFbvLQ9822zc2Tb5tYymgKExbb9aziKTYhmyN1xVv0O2ikfxzAyTlIMg0l0Bkm
UYKKP9BaZKzXrdoASkSpAPqs6Bhc7m0/GCiql5YnvWm9uKMyZZD4fceFux7pE7zu
o1LQCCJS5BUeTc0wG4sf4FD+CiRWslliFxEidnTLL7bEpGyxahT7cW/9HXvxjE59
2PFilGOD3nJfq+lOoftncQBTDQTinZV1FVKyJUx+wjHyhoE6yYv6iGM93/1IPYKs
FU1AS3KRvSwxLTTyug8ciUTa641co/UIEXMuaBMpnv1F8sQt8sHtp8KtkQM/Ofn2
UWZqEf7Ijl7GJ7RFzu2YDDHIof82XYMxUyOrrVxwmU3JwPhCMFlsjZwTft2GiscZ
J4PTc/hP6BCUK/osv8TYBIj/1sqoMTDuQtta98unjfkyizswU4GmjnkNH5lldb1l
LTKZODoQRlnkeAMnqggQTsivAitN2NQpGJDwe7DoFf7pQ3nmgkzBrJe0Vo7vLxV2
tBAP0Fqad7qPFwabgpFZFRdut4D/cfb2cGBJq69N2YP/GTmdf8XoI/KR3CoidjdS
LtlaCp6IpmUQKmvr7ActOo5CLoPrNQAnyQoFfKxboRGqnH//gu1moMOMTUEcUETS
lhqV0ffTyGA6HZirV1SxpjV8jgzAC6F89OmGirLETmSHb+vwkgh+3x0mw4FH2+wQ
9oX/LnEF+pNRd5QEsq5PYiZEdbV5/3DDFDn1ATsRHVbMqv2sdfDpX/Dd35Yh2Yia
vR0Hah8Rz45UTRaT2CCej7vEIvlBG8QGI/lnyRLX4BJNV0TIQmJoLQDTz5r2cxf0
H8sDPEGmXHdMXT3iSg0i9Id4Cohz3iIy+lxL58W/DnkJMtsSnZd0ISx5gjzIpt32
B2H8rwC/QzgaqwLe21UxQO5ERJOxcil6Xe+gWJiYcoc1aavW9n0f9ABQagY7zMWX
+oQ4WDRUm89lRAWfDp38PeEc0OaS2AZ9fAAq5mpLc6i/WxloDKx/ia45iV7vcvL4
9Tj4dOFOzayMKjtaUaJ0IzUW8u7LD3Jf8vcugQV/R5DTYvcIE9Emu1UilhZXRj2r
Votc8gNU/guG1ZGCIOeDyispl/JP6/KCMcbc9sv6CvsnuSGoBTJC/YmuON0UKulq
WDDmeBsc0SIYwExxXRyBKGD3ig0k2zW1GO6wXrLnWIHEyiTHAFFlVcFUrMjPYXLg
fhihdWmAV3b6gDkeTFNQ2nPmfnM7NyWNtgoy3hdiP31mdlsxl5dZynpmSa1WV5PO
tPMJrCE7TxcGqkuSKDroyjSKGxM+DseBJI0em4HR4Jg7ZiTXxTjhmFaJfFXH76Vh
/YIj3QYsSiThsBxY6dp2VFB6bs1b8waQ+NXyykrVULbdJn2UC/f9XkBs5UT6Vrx8
9BeumoTTF/zCmWTmw96BPaihbQhYyKJww2hsGgkbv5wMWtCMHmYhTm+MzzuUqNPi
v/j+D0ZpMwCKfyvdMZ1YUwK8quXVoKaqkg87dXghnhxOIOZJyivUOXaHQ1Xdv7mm
WZ0rTDYwE1XcQCeVXlflgMEbkKA0qBjo6S91K7y2mfRVe+GUCQQ4zaQiHsIvkObf
vMHB+p0QFG8Ah/m1bBTmXsFZBPQN4SL4Rlrxby4tlm6mQaSQshDnfwa8Yjoz+sdt
tcoC+Z/ozne6xFMFCDWU12W+ulrcvO1Zl/zh978O9ZHDhg+/HMEI0SUIv1iP8Mfq
dF2j2tqcGtNFapdjaTV5cLRYICQD4GFLFii1Cepm2iXSXB3TRz0W/WclP4QR8T9Y
KokQtSIsVLchXRhip95NDBRmMK87Hvs8sZuw+hj894ruhJ/8BmRK+jIQqEQEeR6p
zQ/BHw7md7VCEm3zI1kqjtTwHivhjVvnfNsgFbxNK6aOiCx82/BidnTC5iYIVo14
ZkvRsE3DrIJUXX6ZyhK1C1DEvBN2lU1803W/a7wEUovgxLgbYLYq1kTHPKDMbXF+
8Idug/UpG6Trmok4YSeKFwsVZsgh9x0CulbeRmZTAwNL0MXSRkaCwDVOw7kZA4xw
in+7t0++ArAvdgLdMhptUefdRvfpNLBg5x/5Jviz4N9afc5NrIXL/vZHcZk3RMYx
N/R9nHIBCVKPs+EhAIvrQ5iF73kOOt9tZD0IW27F07+3e7KFGm9fnvRUgKOwhM7G
lW9MuAc+fFlEq695J4y05dP4m8YHB/UUbUESTYwkllu2xAriOr878Apc9WANjJVr
tTeOoal7s7B3njFF8MzZ1u19OuwM49O3ZIvKQeB00aDzWJSAtd0DxrIjAkuRg8NS
Ud52Zauwl9F336n093GJQFS7EdnZFD+ErL4DwQkd9i6VTZbjQlLlIDi0mhjlUV//
ggMxM/MphqzuiVGebHCWuF6C733hLsdNPkmXhU9RmjnIOQx9x/VUYceuOWBGy3+T
RYpPBZCnBjnMAyaXhl7wEXb8ZpIEEbV3XIlWh6elI4NLF90grONadZCt4nevqTqX
5FFbFoGFAMiP5G8wE0qZ/vY0dMBeGTvsSRL0gDvthMl7AWaC+flHNe8AELu7rSOT
0gTW71hPh/I6pjJyoTWTXNktHJc9iwe+ERWZJdwV9EOa8A4HsULm+0rDS9y8Jb6f
M5yXTojSE1t03BQ5cS3U+6ue1hIC6zatjiJ/Ugp5yimlallYq6hckI7Yv/jR+WdM
Cd0kP1OgCVaBrYBYOSUMtZtz/aX/hN/ZTWppo6CDbEeV8mvropAqWFYpvqqftduE
dqunBOQMrG+3J/XlI8dvW9d6Tpq7avouOctl/aKzyKEuFzQnfgR8CeX0M5SEMaco
2n8HEvRe7C+NJE+dE1L3bwEnNIvD0z5yb61VxvXufw4J2G/RskDhrYfZM3soO7uC
hff+JTt5kEX3E3QNdQz0/3hvrj9G31NJFzgt8L3LrXKerGqAzmaWk5moM+1ZyuAC
aKdfSSM5shzBAZPqQM5swOyamKg3VK9tT/5MttJDyHQSE9FHnyKXMGpKUrLMfcs5
PjflE1SRxbV0mcNE3y2LAp/+qkVIRFAuEUua4ALKiApvh0gqEV6izuFy211xwJVK
txuq6lggKmOgiAK/f4adjL0Acx2bIS4CCfkJdgMnjHND0TQ+gcEQEMpTDK7Dz46i
MN0910V2AxwsVZHSAZZhOFZWeRdSITq/JLJlIodAiCyth0b7aTwjKMO89d9ad68Q
ZqLq5PHbrAwMi0rEnkfql0LwYPPMCJ8LHJBAHS7vv4SgXVC6RJDzGA/tw2c9cdtc
jtIR81UnI/TQX9mAfsfzdrZSgMOcZQa4mNR2AU/B/GL5r3dEXk13WBqJsGVjqluT
5lR5wTJ0pWA3vKPZa3VMvD+3kpFaagIIUsKBA+eGCFQXMjUO+VekJUtn72dGaCLA
wygn30jtyHeTBqHxJ51LJMiRlLnz2eH7iNVYwszn22y1GCOHGjJmOK8WQrCH1s3J
V79SqdIeINBg3GSln83qe1v4GcEf6MgipeTUMMK4DIMuMxrUZd2WC6IpVDhiFVpb
xndFcsycSbSWOMp4W4VuXdxMsjehFXhTKSQFmBHwvdz+yLSX0+Lx5YbdeX94Wmhq
Qp5yDL793BRrOwKTVE/55bVyEz9Dotj0cnR4/F8MJMhViz9FLcW71duYicRK2ET6
My+3vy+wMXimqjeJvYOzu3Po/C4s4pLVICziY/ENhLruZ7hKSnD2RpY/372k2onj
P5qlICKCPEWKB+JHIB0CXBeFp8u0lEHV2ZQV4RM1eDWO2LXg79vcJLaVekdllZXU
fyEpsJSVEdkyMLPzVh1AZr63Woz8cYSz0tVh/Uh/H67BLv+Qt0ZtJnlHeaugqu1n
l1nsrHajMVSfvUqUV9lOsKCl7UTLqRgllgrebu/EWlp3Tb5kzD7GGE2CBQxZ+maG
3AHSkrNI7eWKZTjfBKD3iKHH6RyxLGA3Od9/as6qCxM03sO41wZoS8lYbAPwgs0B
Z4lwLIs/ZnywybHhJta7A9r5LnTsxaydX7OZqH3Fec5Ky7fPm4/ev5gKT9qkrX3p
sZnav4B/ZWOo+XrIGWoTjizwWxjwHh42TdUHSvc2Wv2nduEGXTKUGRlWp7JsyVen
XSz+91mPMqPmQZHm4a5z9SfNXq2H/4xGGL+d/YuvM7FzbBAQadKlqwIXFZq4yVWz
6TVCOr94GEv3En4RxelZOfDQUp2aBsOCs8tUaN8bCAlEMLCC6ja5tmicnbEiKPIb
mLP5WrLhKVZ0kRg8rhijWqBHx+I64I4sN8xhP7tUNGLfJek1xuGVpnEbi17D7TlE
+UC8KGNvtEpEnbF/oDIXkytlMDBg/Dadf1TOfYJXhb5zddO2NQWVb42Y6N1OKGoa
EeU92tRBoMuqDGG5kVzNEo0IPQk8cz98ZvafoneN3n/SosiUQT9pklYHjFXVZNNI
2PNkscQLJlxTYRIbeclmqXreNnaYYo6MHkIStDZCppccHnUJM83njiFg4EPQZvWT
nLLzXt1Ryv8Vh6HUaJy5oApLMibQbbFy1MdyCzSh0bbl+kIo32NoHYmqF+IilYtb
FAH4c7yw6fmQjez4CSmZUl4E+CjkUw/SxQh+86wTqDiXAW9jKAg6Rl/ncfr8V6sR
prQ8SnGur68kRdzpPdoyNRkpm25JobDziLgLwbl0PgADyl6p41eo66lCEIOppjCR
2Fld8yEgDYEMgdL927TMKoGDxRfuwSEcMkL9TkJ1nw86nr2GiNX5pFUy7r/CfJQ7
bkWAp2SaVE4MRIdHgC6bNXGRJV4jHl/aX5I6HrzkoVShr5G5cbHG8eWX3laPBXIF
D2VH82ec94oTp4MJDHqCYFMTaJP+s8cTDes77icooQZagKbl7dR0c/F2fiRrgGxL
C1FB03onKl23aDZYP6qfM+CtPEdzrSBAph+w7tlsIpeWWBDMcBEqZyD9a4hBvsmD
YptL0jWc25HMF/3oLRwg7UHaBdE0EbSHY7lV3/FmraINV4/d+QRiECRTUPuRJG6A
CBXvyacy8bu5ECWG8+qwWf4fW3z4lbT+sBNhlDeEd7HLA0TDM7SAgEeNCURTtLuP
fuyIFrypeV+YMiTYEqs70HQBqJSR4K1EXj+ScCsozQ0N1eRHIMESk0jA801pIIE3
sdExvM2shrufy5L0M7ZA3ltljmXfI+AGPayGZMsy4nxXhRvejP04YMbS6CSq2VYr
R/ePclGGhJ4A3emUVZLX4EihBLIDhRnzq8qguydrL61eVY6AmKCdvziNGTrMzYCC
lExGjrH1eNslnaOc4hCqNAOD5mvHqi8AAQBlynxXfRDUjKugjJgkNH4rgwz3siJA
ZKrEuGgaNs0qy+ZQ+gZIXS1IbD90PvB3l18Kh9ZR2S0k4RQK2yZwlXOzoNO3zXGY
y8lLvO9uyyoPUFMyx634LU0e1AEx3V5Ca4k27Y96A1qD5Qd+NcE/vLs1GL2wayWF
2aAP4pe+CZbaixtJ5RMtDcqZ1SE67d6AbxhqSJfFBk4WkBeSEFnvpTMZ7/f+xaON
RngultnbaxUll9qFRhyXV1adburDbSelEBpfVuJlfoK6OoxQ3p2Mtrh4OHok1EeJ
ODQOW8x45KtUCmdAfa2RKJmeBQdprERY/LUjWXS57IsT5pCJlukHajK2qOLXzFfS
LEAeS2SqKfJqtBRK3yvuTsiCOlU67qtZKKFnQrLs6ayLCqThs3VKumFjiliIffPi
rClcjFc9d3NDXg0yrnNeVsIstMMiRa6sMR0uVoQMPNpJMHSqgTXNmfSqA2JvwxKb
eT96BndhDb1MZ1qdcFobGGSuYxDuy+xGyyq4HG8G2aM+eR7YVU0kB+ffon6+eNN6
Lnim9e304BIWU2L9pHkej0TEgXLzT4aH180ovYg90sI+66qEkkmebePrLA/6S9Is
UvTneIdT2byZXxiFpVn5boGxizqRcvhkrzIsPaMWShdiGWXZCC7hw6F16TNJAeoV
Q0wvLdndCoSasqZoBMBxF2J53kcA3OqTnrEDTRj36mwzfXk36qW2Trmjl+SpZMBj
ymDsKaqZRQWbVeor8ZKwPsMUtdu61GC4HHgVQ6JaoRkxuMvKyvKJvsEky8h9d8Sa
fd0FbyFHm51yKsmkZVZNh0NlUo9L4gLzYyEvdB3JvkniAjE747Fc4Y546hfSX9OF
NW+sbHQipypghKWxRr3OqU1d7ijhPL0aKN8sxG/WcXfX5Kzn9mN3S4b6Zo8z+zpc
QFZRick9p8/epCYpXetFzfn9wbhwS4J6BP8lDjzUvM2p0qJp8cv/Zatecg0hRy/3
dbnQZ2Xw/QCuzRH3tw8hjWsI85dqqPg3kmQtzCEn7snZnKAy29pkTQ6taNcUZj17
Ry7P04BNUCgHrChdcAemOg46HE1QXsxLoKfn0Q/l4kjTmbF4rxqpGP7cuWQly0U3
xKNwyG3ft80cKGIzKXXbCkIGYYxHvStB9c9IF5LbReBlE9NyjTA2bM3MiY3O4pBI
UAqjsKqAXhKwDLRsrUiPBiXZfD7xb2L10+8JcmdPy7v7D1DqKyiQgymfKjisx5GV
jFRRhg0aVz9vPDpSsHQZjQV0A8a9PuiQ2kINtSpdshr56a7Eqghm+DUbZJUuUj1d
nkMed6cmMV15x6d/Rw3ic600Z1Ty9QP/4D+xF1j9/ggwfJWU4T3lyR9b725AirGW
hMtWosaG0s9eb2D0j1zqYecbKK5ZRbCvwSo3a2tk14rQghuvbhpx6pK3PIztDdOu
MrKvkIsZ+J3Ro4BR+EfNnpEJj0SNsgi4Di07L8WZ5o97B/S5fg06nrdK5JKjOg7x
JAQKVJ30QVY9cbnMIsQtXY1+gnslsA/8j9tIxCPIp5M7Snm47NaPifqFeUadKv47
d5y53brVtSAWJtUyatnQWCr/BJJXOYRARs/vG2oXL11nwUzQTUimdnkC8T0kctNw
yXC128ghnwfE+eflnk1W+PGwQRTkijBD2s7dnxywDmC8SBqCSzybaGIdpFlj2Tov
oNGqCOZNN4tLm6o4zi86zuPr9o3z88oSBibG80qVooGgmsZLg91UJOKxSqC25Rep
mkQBGxvORR3mwQLF/QxpcnTFelzQCmh9/oDFxUVvW0MdYfRlggPPjcN30AQhoI4U
qa4JStz8PwyEArfJLyXLQrKPT8z5uBh+3KhyKZKFRATOhWjdHBnSSjO0y7Rlp4Px
DCJhR7z5KlJoqbrndskjI6FE3fVWtJk8JfUNepDC1CFs8s7e4aQzxfrvs4B5hbTp
2kPhGha7/1OIib/eJ4Q5Xg5tAtuVwZcHjhSCJvPoRRDUtIZtapvJW8vNMBtNnPjn
SPwICgtNjc+To06CVejAYrGv06bMBrlajQBNrnXswOhOzFqqOid2MBurLjrhhPOw
hdAK/UpFXzRC90HVme+teO8f5FfHU5vbN5XekCtPOVB5pt06i3vSo61grLExd8sw
CWYNnRXFDwXDYtZGb2TzbLL46CttHZLGbp+JViK+JTHhLXI1VHejA885c4Re21l+
NJfHkhFHGmqM0c995W2WOw1Fu9SXBuj3HPNxZh19oid/1nrS5hIi8MTQZnQIjBMv
L8WuTzs0ELSvODuQ6sMoV4ClM3NBNLvGmNgh+SoMp5gz5H2eoCTEJnQ4tc+d2k2N
aVWiWOw1hiEcNVSCahl1750AG52UJM/wqlqGgF2j4ZvIb5tYXAc/7/8AP4lAW3CU
FDb7wwpfXqF20QmeyHtWUZ0hLLaQL1GmUxe7/bdL6qY2SKqbOHRjasd4ndGD928y
RbiPOOVpnQ2bkwJJHyn4e3kVAPHCOGk547N1KXxfZR0PuKL2OCcLGTfrPhUzC70Q
mhjUQB8jVOMvlJpT8IZ/+CzSELalna8zau9+KvK1EW8kYvONOpXqmi6G421KsUKo
5Ua1UqhKGue0m6RxLNqlujMezkWFeuUgxSuqZdJihMGXQWXR4uEgZiRmNdq8AGo4
HlWgX9BHaqpWeSw8TyINRUtJ5rV6wRs5x5bGLRqnriGsxkYWBNbUAFjKqjlinuPd
iOcLc7kbsLviSkR9t3DVwS3F0s+slFH8WJhVWrXzvgR4gpbrmDyivIRXzJIEbcBR
hyFnqFj9bpN+fJiZdsbzIvWNEGRso+ucIvxQEYZoMuQFLMUNDNq6FtaZORtdEHjz
K77ZxuhcLN2E6oY+xJf/6Ch2+Wplv5kqZJYCZN5s2ph/Z7Y41g4K6MX0bX25c81s
pQVSvcx1ynETJek4udT+2T/f+bsUGrG4dGd1sTiTm//kUCy+25jqI6/IA6RelRqp
Nj+Fa2j+j/S7sgBwl5Ae3Uxn4WNJoqrApQcinZZdyxWgt4DNeiwnF7BuOG47zaBO
AaJaoHKtolptqD2Ayqkh2B0UosGOr4b1ff5IsQis/SnZYGZuVoSh1Wz55V7DHASn
TRNXUkiM2yRGfX2omW4HA4A1H7spOknH5lBjOeB82UIsE4PrRkrO3l5bKGVmsF1C
pkdAKQCQ6fR0ijnfX1Lx15nhiua0U/hxyUplxcMeye4JV5tWwzx2l9kiDQh3jLod
15M/aoMAylBQaH82TvID28dtBcYIZT3Xs8qN3TmgCVT86Wj+mtlrvzyuTcQ0JaMY
lld9VvoXF0Eba+hiaBHeeSSrdpyxf3fXHdF91rNJgwlbrNK3cXW+6uAdo6HerpYl
I3VXxXytC/NZe0ZPzaSw2k5AuUUyBK7GytQJLdYD+/6tA70gmDQuQmEjhSZeNX8+
x3r6c2n/wnhDmivYeOhjoFMjYcUmZb9KYrPDX0MivDaFOuycaNfw2tkA5GkccXNx
O6tPGPr+JlUzcsFuMMycS7/abLVZCKR7o73w9DQdWeWZEW4IeT0kVkEUKdv9Gldx
bM2YWijLzBA/KbSKNTFwjn543ttV7kChKODabgWeZDogZc08Zvf+CM7MnLHRmPVI
gI1J1iTXaVrMT/3lrUzM9RZW9PLvGFkM0U/Puv9QXEonV6KePi3W45mkdtQ4SWFt
F0hXZC73fRiBqxRtgnoWBRh3/le7Qvpu9aTwe+hKeYEgLZnqr7wxAcodDMxbksvD
nK1S96Ou8ReeVpRlLhI1ywu9Zw5KFR/USJiAUyBfbcVXT+zXhUj9cFVK8jSAuqEA
NrRFRda9gKcoqnFsimD0pxsJwy3Tj13FgRhtds4zNfHFYJOpkyrBZ9QP/8aZ0/4m
P+LtOfAImshU/yEasLdMUVOp6k7bmbkHJGWwZ9ZInUmQ7oiYo0P8+UxhsRe91Ltw
hn5RY7aUmBC+LLdMzIB2zv+iyeMxC4WWqGXZzCoGSrdPCzK/ZMpS8Z5uGQyZ2hy6
p7QdSIhijI3/6n1+Wm/yoTqzvRXl+9Pys18mUuARkfAOqMtrIDjueNOS8zQiUWnW
PPk+Y6wwSZdYirt5vH3rEajvVpDwXqnVaqQXfQxj9Ov8+kDmBpIB3D0etTn4g1Y8
XerGr31c33OcLZirM9LAfa73SrcMSpZY2KWS6Kd7jRpE/bIJ7tRBvRIwabWrWubD
3Gezg8ag1tVAif5jVkMhGgWh2EtMb0EeCK5NkRf2mAnwk6FZWvVTlSl3Y3UZ/Nwn
smGVNU+JjQSCXVi+NoZaVdCoJmzWjPqRcu9PSgClrFcjV/q4P+krHD7DIhNfpYGC
QDcucLtU2MYlLVKZbd2JehcooF82ptH0DtI+mpo0jCY3w8BoLDoDkd7XwR02UYt5
1TmZFy7T8WSx7RK7Wb33nqeYaMPtSGcnRFTa1j0dCclH5uvs++SmHRD1qTVmeLxh
Fc7RUCBG5wxmzCFaeuG9TjqDlJTT9LxNNRDYDKprU5E/dETPAuApeBoazS/Ftf7L
GKXaeMelFvfFRAUEAllz6iw7neX0QN8BULbZv3u6LXtRYA4Mec6NNa4sLEf+uOGu
xG57sv/t40UTjpAZFhUUt3U/Pl9LCMGh59SYPyHJGjyfgA+OEVkVq0Z/rTD9JDMY
qYAHTx0WpRqf8QBaO5f+a+nLf/IiFOoCjVjIgvedcOvcj6XuMfff1bMvVVfcE7vx
mdGye2AJ39FGaDLMTx0MVxGT55Gb7G7hnPQ06flLHQ3WBDdEeY/jvo8KKRKB33+i
b9sh6Ln7OXUhy/b6Cel4pBMloxRs5nptWJYqjrdxRpU9nBtvNY98xxXdw3NqHKi2
P95jv/7jc9Jie3CUv5C20YjJ+IbkUFhyWj2snZ1sca0X0aBmhdB8Keq3fdQABEK0
xO80UD4OSdi5WZOhmxMMxNax2UTroLlnDPw5CNoN6LSfdDtHk9tqfI6+XRh3h2cy
e8MC5PtGNv86Y0/chbvDDPqi6VqXKyjAPOB6ennvyk1/jPSaqE752+hjHvpQ1gp4
SrNulwnsOqtSneDI/xMByrRhyWqdhqMwaqgxqIrOdCKDHZ407tyw+9Fb8inioPjV
BK09IUtuZUp/NFCngODV2uEtYVny9FYaqfpm+QwceHp5RRYjOZmi+lPkbie9hu0W
8qKs7mSq6bwDY+biNbLH4yHNYRLV5meuNh+jT4DXY1riG6kCcJo5Y2MCabR70NS6
LdkcDNkNuDJOI7JmTtTwjC1Cao2JNucAhcp1eCdlaAVdbLmG/JCgretJ5dhHt/eg
jlKsjzmVZxIL4+m+5o3htzdNJQJPNnQEEJ5DPzqEmKliKjPMIZ3ZEaeulM3edH7/
g8AbMVni5G5gmwdl1qA/CUc+CNTpXl1ulkxxFN54TUi2gBSSYCSH+6ThkW6Kwxaj
F5iu5xtSm39faudUMUwSSEhtUPBnTiQ1Fc0IR90Sask+q/xWBWp/V1r6Tf02mMAo
EaLVdj61hTFEUi21k9RuWBBN318ko7eDNlq+MAjkJNP225q/xDS9/lJ42uZEYQZV
ReQ3trRhCMZZvXHFtXcr6pyVqSyWz3adJur3+kYbSmkj9kLgZ4k090gKKHSMDH1o
rRDPlILGXXD8zCGII+3cVtUkb4JVIwzVnUxSZtG+a8cgOfIjRKf6PtjUALQYK1j2
OIrs761gTWuAN89inI4O/+4XGV/7c21ubAHQIgiUzXpXXR2jx939iPIPuIH6mE7n
J5JkOWPb98v2zmWE23OJhsP7gl0Z7TcilfTHgxQ4/4pR4nUCfivPeqSxz8r1KPMO
usvKOLdZH5f71KsbO+fAmDsus/dlj33NlQv4S/kcWB2MV1Uua/hAj4eHU25mIA32
S7Azk30mK3cFlcDlCeu5Yu0hWA7x4HBwNylStopyy8Hp1zfLkfp13di1IyxJo0NY
Oki/Sq4+F6cXu2/O9ofMM3qLAZamQ3PpCmrbJY8FLLCffNJs1PKj5JbTNLlPhlYr
GEozOd6fVeVNfACm9aFCHeUfJ1o1a/cnev0C3j3To2ZilIwRZ02tntYXV5HnrhQf
8ltg09tatoOThaOuWZehgStddwvx01GlOsLewVfg+4XUPiSBk/s92e9WBsJazyLl
jQ/zhBMm0EF8iycIjA03ODba7GfKwCl+x7l+5ur9nydvSW81cX0kyuUbpkvaCXeR
yOjLwj2ewYHXsAaHRrT2kFaZ1qi1dnvRnonF7SpjpGAJf6aH8wNJmNYsl1sMb2FL
39Z1geHx2Z5ApGGzanwaA5hKROponSWCIH+0BATqXSVWcsEN2QWH9YCiEowj8nJH
h1R6CYJq3Kfkcr/bgA907okCqjLGShHq3wToZ3wO3FEOv36w+5s4r5pdPGlP9Jta
CtiKHZ5lTmwZBXqtq+G7Sc+hdcW3kXVSZIAR3MKYRurCgH/5GASfqXCoWSzRmGV+
rvbRIhurMj5AVocB13u2QneNM2Gejn7MkfABvZA9U9DfBPQ1E8OvNFabDWouU2l1
hm61pksxu3Vc4IoecAzSLMpHCn62JYcpjMEtssK8kjbxqg78prs/UoES7qdNCc0a
bAqzQFab9405EF2618BiS0tT7OKx4ribLdketO5qZ9gYOkBYzDXQdGA/xAsx1qG2
nBchDhLJlCA8twvH0kPSCJDByyFpQEb32SqqnvHabVpXJkVVariP7toUcCVthlO9
EWdXsO7YTYrNWR/zgtNmGm4tVLLW2dDcMFZZq74b+dYKmLhxWLkFB9WbsY7JTe/w
5bbjnkhXgXeJbHDqDV9WudTsH0oa89E8wWQvbDiwsFCvlrke80tm7rrkwOR6W+Ml
i9+v+RhS8LJh5rh+pdANtbXbv8xq2T90HIGgu6Bh2T3jcVW251K2jybDQ1sg83QX
JHKuEgCGpWXNYLjHBDrLod1+egWh/zyhBRVwIicttjBzzTVpynO0VJ5tIAj8Q6yq
m9uDPzgCxNU/M0CufD/pNrWPYnBqUF4ASGgFDbzlritk77xWJ3qoE0ClGXqK9qBV
p0YC2EBrBYYczQUGteSscSQrrrKJn+LO9bRhhTHRiO6gScoeAdODX41HqGs9UdB3
hodWer06l2Mr7FMQ+B1Hm3oX4w924WRSndjeBZnkjeebdREDPkXTz6ayGRUDnwnQ
lWfvAGFhGTkTeAXXfrO63CO3EvP4SXGfjOHGbFmzY+GPTYKGPtKy+R4Ly2B5hFMq
ls3JEzyq0+GJJAWnGz47RKceyc6/MnMJVY1zFVyYZ1Jy6pX7zCMb30Z0RnjsvaAK
Q8l0wdqHJxF9JzFwvWKPSNf2s6EwOhJd61xTgIb4ozMVae7gKM5209EDd8PzxLU3
+V8uYo+AXjkNmqsCziLHnde7HPpkpeBZIvIEzElpPBILZh4aEhnAubm26g3SfzMv
11pCE8R/cbMtjwKj/GFJKA/4FySNptBlWr3KZGwLPepzlUEa24Mm5iGylPSl27EA
sntv2eyZXuvmr+LwmUO8dxDFDcDrR58VlwC1d4/iAijmhKYVJvLrEEIIyMGQJ+2W
+eOqkZb9dyHZ7pe/eYHYU5K1FnIuXEB4EH4fHRqFnypUM+sDLcoTQ7WDZx02sazG
/vhD9SQRvOubKZns+j/CvLQJcH7HQm8KJLsbpgLVyYULOBYHDLCRh+fmQaFfYjVq
QH6PiBcaxmwpEJVB6Zq9njiHv4v6EMJWCcrV7WDq04p+486s0ZtSs4lpanjhtWi7
gIQBbgCM7Lk8FcwNlZVR1jxrsa1BzCFrtBQcRm9LJZbFK6PKK4GVzd9oB7ocAxRl
yQVyTXRJi6dwaiGpZJfZYEYEA7ULtsXmquoKKMC9vQ02YRJy/B0lncJ+57j8O6IQ
ZFe6XQ/wzsq6e7n4vOEHtdwjbF9f4013f2dE0w0/cg5FLyKiQdCZdDouYpcF1Fx4
RzWLvrUDrD4E8HYtbt3hk3epz3STy3b7WYQQI4ETw0oBe0eIfqWT8VAcr4s1Xjt9
Ype8c3GWkK6IVsGd3bCtcxRqHutQMAhAr2QJWOwW2DUBma/WxBhB7eEHjs9kX4Fu
WFtT00ndwQ/xSAASSa3jSnZU60VmdH0H6rThIR1XB165L5xoQE5LAN4r647q3Yys
yYxSHoed5rCPuCktvOl+hEckJmbNc8lg9X86ac5rVnvqFqch9YdgZcZQl6EKeb3A
E1iNwwtaO0G06glQFB8BpLIar5bQiE7df9kmoFzxvTRRt4Tf0mKTN15BlEPdV5xF
IPcD9sIHhPTgo15Th1LtiCVHLdiW5LVx9vAoad9tHPv64b0z+arpcQ8iH/KJS+3v
Q/YlQaDZwvoaRuGD/DqNf3wdOUruk5Hv8Lh1Y+75ksMLEckfJIEROqrHFoclPOAh
r1fnF5rZzlAE/vH5SW4drxhQZG/Wt72yfrqov59y8SQkFgLL+ACsWqBvjzBWvUJI
vF+yLRmd46alz/ECEl6RHLZCrMSSjL0YPp3b7wWRyIv9X20U3tzmICT2CYP6T5d+
2epxk9SFYFGtQXnBPkUqYPobg5qMrdIUav6HzsFFTR0tDTJYRCkBNKrNO96pYfs0
NSn6JQO1Gery521DN2zIFziZsYNTPlBXXu4kolmCQ9qU/6yiuAc7OL3LPECVMn79
KFwvf0eebUEDZhnMppdtyo4J9RRc0sYh5EJ7yxBV7fzzs52dmxghkDnKI6EQjkuj
lr6FEzCvhPHxazOydlOMCnQyzClOiPziGeMervKiBpdmGnZnacUQWrbGhzqJt4y1
uzU5/d8pQuG8bHNDtbfHD7fBulgN0lPGhS+krcTkDaBuXCeHyo+POoz7JaKaOTIQ
K1Z+1L5clYwZv51lrGlCOhlued7Hh+unvB8UUFdIMJvHdAdWp+lze2ipI5Q8/4F6
VhWa18JjfIUIvyYncTxojzETw2snVep56uDsap1udTCcd9uyraz1vkvjObd48JBE
TqgF3OSMqy8azbiFToIcjlktxRK5Xw66VN58A6OQO4ZQJMgu2agRdRNRMKkdaDoP
lzZyIcZoDdyP/GYSvmULukFmPL+Krx3rdLCzy9sEmESjs53O0QYQUijaf+clQrUD
jfI74H6AG3MfLawPXdK3gxntQsmQHFWWWAZ6I5/hSfVrBHehVd1LAUimzTb3N4yh
MDhzvCu3tStIdvtA+sPyuo/UttT+m0Axn2/hiP20gfEc+s2gjaMdgGSx+be3Q7vs
Yx5aKgLtJK39R3PCmpeLlpdD2BkUvA8vHnFUbEKPAOfi4x6ikI15tkSY6b6ESyO6
G2FmdGfXfZnFsxsnwfiZ+zXt/tJ0/wMzIOo4TGDu2c9H7gZ5pHmO0eGsppXQ59/I
Un1xUHcgPw+c1nJ3xHigHhiXC2V5MmR75FkHS89j8w++6mSZhAo7NYVAEQVv3Jp/
EFtc75miFHhUdM/HXflAIgIbrgB9+ByHcvB7nCsUZh1PKToB/CxtkBcvFu9AD/Gb
OmsFbfsWZadHHyU7R2S0gJEUyhXq97wcL/VkJ8a7iZib5DL0dev2QSVaRK/9GqIA
KuNjDvM03arSf6jrZLLeDlI0zOvmK5danoaQvP5Kf78rUNiEMDkYD+vs1/xtmTDv
bj9ODwKkd0Q/InoZWZ6CD2+h++XIdYeFogGJ+a4786OCNYMEAb73fV88qK/Jb88+
PDXh0BCOJTbc0FzWnIL27pN+VBSrlaOFqYrmbTeeA7vu0o5dkQGJfQJcJBesk+BX
x7Yg+TT4wWA5Zswz+dk0RSLyA2QSNrmhb5GH4W9qHtv7bzVqT8+1YvcPAwCmSQuo
WxcPy/OXb1P71ZwzFAXpuhOi0GkhI/xf9MF9utC+koqYOnHlyo0i+0+j9VAsNPyF
SOYspSjeeqvqUQx4pkbsNHfyzAnKbSgLDxkf1o0CVY56dpAgUlMiWjr6O1naAWef
OGEzMan3lalwMZpPo5cZuhuxZMb4wivqyPbZbMLNxSKoBJlwgVekEJinIWMpDcQz
kRpqSnf58QmK5qYL1H8HvWMUVtEkGN/WDW+zKqWjrvaYnrO32+LwJlw3Wq3ZVeQd
GZwAY4ANWHhlmZqgaJC/wwlCUZ98Kgm5kOxS+Yg+GKEpn5my6kLiB8GuBS536gM6
u/DG0m5XwttjgmBsUgQy/659rwr/TSwOq/rtU0RAPM2ytHt9gNMmpKmF8CUXUykx
4FWuRpzYQqLA+41oLGJEHMs+z/v48hCJ5zucFN+Yng8ikL3dXxCbsz2W94UEIHkT
5OySEvGZW7CMBWAlaYKpGX0a7sJE1EipODIaYDalEgFxZ9JB7mFTQfXf9bJsDZre
6SLHCllSJmHTZeJTigMcQDTCgKI2CLR9sIExu4xRwqPxzasm6EGUs3RQ2v4d/yzH
boePJTCMSHD+VuL17MNG4xxh81Y+aeZ9AySB9LSz2Rjkg2Lc192r5AZevUqwstWN
oYuXun/ImpFpCDMereV6UJx1rECpaqIQ3g+57/wlz9Lmwi9ueudCrbe11pCojHlE
Hq55eNhbeS75ocxoJzW26C0vZlTP4L4xIpPmQ/J4Zk0SdtSr7lpw3SEpkN736CIj
GryUoCXzTv/A/rsIZeasP4XNXqtCU6lKV1/n7eZzNSSJJ5z181o1sLqShieLi5d9
vW+Nljq5tCuM57+iQADQiqm4DXUQMV07Cz8RFh6korF2GV3nu/CU41xM1rJsEtBL
xQrgmlmnVn/fTf4pyZyUHpOG6N/1iVlJs8/QXTIYunha1DLnpNbo+KoQIpDZtXgT
YPzWaCuwpOOlt7KFLqyv7n3pJg6d6AEABqDYWDOEftt4k8aDZf7j3v5Z64SbW43J
OxJKQ4e73BtDz+KUU2oUxn15mLpIq/BVdkzQGqqcmSRSGigeMjFGENkiH+5m3jYW
YRC3+6hqdbxgI1xjYv0iSW5Zu3VXxKzSlQ029T7qXD9h7QrtsJMndSsHBwCqWWhw
txEt5lHurtUwZx0HDmq0fw+MXS8A5xJF50/RLAijCouWwvJ6viGEwBcvq92x2TDn
eo1rMwK0lv/SapXJH4yCKQDVwbqk+7VM8t5hNyLDAQgqL4eumf6blrwMkuMhZ7aM
znkgt93EdEUM7dX5vEs6C9u3K9GXxlUXuKE9cM9pxbEbsb2KKPg+f42VkrlpNKIT
qnPWJBSBxVbSprEQjbyjtQDXVJXnKrA2u6hkhYgFx5MqLeQRWwjGg8KLCg3/igvV
7AlJji9vJxFVVhrL2XeRNSg0e51oPZIyFAk6nqoUPLd9B462hez2aK+EwNSD2/z6
pJPsZ+/BhnbLzsDLHA/hV6rYmCzkffaBMH6TPX0tNkKAnk4V9fjzGrlv/oKBpH1g
gJgD7UmvE6KmRcz4+nkYao+iaWEGN3L/IYnPF/BwCObv2c+iUX7SwrXgyUeGVbIS
QjzJyHN88DHT+nrnKt90ZZxWblG/uXkAduSxMaKKXFj6F/SBnHQfm8YgdeevSaUU
lU4CowiPjxg+IeXj7K/EISxCRd7CmQv0+2VifATpK4TKcfHmOgIzSEWQ1lLOGVzZ
xS3CaFkzskS7mgOyGazOFLPTr2tuJvTFJIAO2uRolmxgR3q4ACQfeADPp9LZZyvL
vkysMZDcrinJlAPvj/oV36g7YmLMzMFBmzTkHiT6MCqKSEqI68hBGTjp3oqRUcwG
I64VYwhktrOnxvqpYhQui1UL9l/9q2We+0klYEmeZKo3ocWxw4yNRihyy/esIR+q
iRzmxMpKq9RvsoBDTgBqws6Bpkpr5kypwsd6e9xdchf8Y5ZNvb0FmJxx2owbSKiL
HlDrTq1kLNueL6ieUudhfXBDwVC8WQ4zs3vuUz2dPrfSXu1NH9oKz7IeAOMelgmm
oEfCBz1Nn/OKYWq1/euFR4YQ6UuI68NUpFpJtOunM/4BVgBNRx3xQi8rpznEeQh0
TTZKPKvW9Yd6Ws/GTYphwbLu27teFI8tP1+QW1lXTKUkEetiVi5h7IyaWI4U83pU
ZQCi+GfcsHOUriVwkJDDzPjrwOZRPc3EKHh8lX7E3ojdAMP9f4/epwy+mcUd9Eks
JUtPqP3XEaFfCf3Oz4mkhZvhIFMqI+B2Vgf2yAWuRtunlyGzsA7sb0rzNQq2GZqL
zYFe1CeKYWOQPo/+pPAcnDaoSYdaajEqGIW65sFyRCRE2YGCFdKdGfaOJQJBLcqn
VmabXB9L37bIClHtoJruxKnjRbFDzD4IiRsoCpKlkWzqNRit/IJpQbvzZK+l9Lww
kcCIVynZjwGN3naLvKQ6/ROQKCKcF31s+FiqbqBiHMaVpeejsaiTfOTlbU0DgXwH
zNdvcfmgs6MqyUnsW+hYnVi/pBCUHfcraxvd3ekX781duIY2/JHpHeaK/aw+rieC
3BNeYB+aKIbKssRQIJulJ59ivpwCzVqk28TfH0PJLKXUonnaLDwMhJ25VUlHol4O
gTgEzTYcvMeBbxEi9rXz54jUzGxjr3UVaHkxQtlhNstKGDb1+UM7FpKItvQDrv62
sZ00CTQvdtscvJBHZ1G5AfZmNggBiLVCrpKmZ3fWLEtNnnjMHmyaRZxeN4FCWo84
WDWFOF3vEsQ/FI8Gsmg/L+iBgKbO9ZTbANaoawitReS8DACIMZWZ+qDA+/CGZe7e
1e+obtxUrPrDTEQPBd53HE1Es7iXv/MgeYypzMnARVE/iD6WZoCz9qUYbi9t/kbU
Jro52oLEDkdlGO2Ac9s50TnWAfm0UxrG/HEACNn8+Oa3DE2zTtcLhCE/O4/lNthg
5SyBnL50BO2iapybHpU/gBZvDsQ2rI4n5jti6J0+4/8Au6WO1d6VyvR/E6lL5Gvy
Yj0kXKk7AXLxNuh/e7hnYRcwhHxYMzbZ9EpQ/HEx4qevsFPi92qdY46jRTQpDa9m
j3hpQ3jAd6jrbhpywQSN8G81L8Kq4UFGn6IyPIGRcGkzRg3/zraDQGoBhLevgpCF
1O1VB7Cv2L0wETVuwqADkrE7Li8hZNaa12pmza+34rI4vOLK1qftWWeHZf3Ui2fE
FoIXnLds6Hvjt/0oD3yeZipmBGb3MCWdD/fp5cnbQGNjqtcclAwTBdJBqP4mby2h
gZfnxffWHddfN4X4As50Nlr7vAvuPNERu+P1t/fsPNHt6WDt6p6DxfCwBePzOkna
YLGVdKtuz2fP1DWAcKDNMt4stACxxk3zCgh1RQN3q44bcQN/hG5+9/ojbyWpKe77
9SY/+8mE8iKVVejVBNjMoVwxMqLy0XinVGAmSlWTvH7BpmSPUj4A8FYsbFUP1puE
7148EtH7WcPF3Hw+E5Gh1lFRsATVwIvL/lF77XyEe6zJgoBRD7Ht52dlPLTKzout
VBDPyhg1Pf/EdMgavOhAuWJi2TIQtXvvZ6247oY5nZ3BFvXRQgwm2WzjxIyD8VgT
V36kORrcIg6o9SbLlpKKmCW8T9GzhkJRsQElbqWrTeEARF3367qBV9IqSkiiqhcO
QeSvKK2Mwa8TOhYQOXh/qfJg6T2PZYfT4DXdHHFxvqWfJqxVKUWV7YRsQWoK1XUW
3/aymdRCkqD4d/Q4wX+DUwP67gRIXIHfDpw1ktm5xBxKqe0QOMMQAJGeRRdlrXwy
pGAhWZ96TU5Gv3NN0G3sHnsiUKVNzeMui1QGlGbEvGriZe7YaU1W53xg7A5Qx/Sq
UVfltpwS848tTdWA11KWm94MvzuJ7iVwJYvI8tAPdor0qudSmtsWDXCRP22gwjEw
uFLg7pMjpBG/9GlGU9FUEmkeUdblxkEOkCT+uqDf68eJBDt+sjKbvN/sVDHk2389
9ULVhJaAZ4pGf4+R8AvMYy0YnTwwe/Ic7jctI8bdEmtngjxmNBzfVOVzhz9saGjz
43Y0Icd8B1KhxoecWHzqU5Q/+Q23vfBGtc19/xQ1RPSf7vcGRRsI7f9/io0fGSmA
D0fV/+gu0+QNUjW9WtyRO9AHhiJSUjjc3+HP24MPZSNmDOX/Ns4GtVpTjFejN4nI
N14CEzeC5u993DEkJ+ScMuxycAtb61eo+tJQIeXUPVXLgPI4KVStU0/4I2dRGbCe
+ifFImGL94+lgQhbQ7YWRybmiz+Dwjz3YwqQvjwzXFhOfpWxpsP5X59a4PKdxUmo
SHR7DJS7ISR7graiUY2azkYegwF/oJAP38J+B5stw59mB4RStW+le6+8+dPWoliC
Vp4BhVs8HyAIbia9nKVotasxAwUXGPdrrpWjkA6YmrbKb/XvhSBbP9ea2p/TW3JL
MZQ+bEyirbhXBZD25BKeA7lin1kGWehAtII/+autLb6HVFgNRFWCOkImvbfDEmyP
fvpeGxvYQ4VkdclKsOpZ8EiZxPRvVYybeQa+HfgKQ7/5YnLOJFV/YEU5ApQqGRD3
U/+XwqIk4yN9M9nVmojL91Tz2aNKKdpDdcG3V96Ys8+PX3CE7/dUvHr82uNku1Pr
AgAzyO89p9P3of1mDNRgeIeRp9sTXQlBkGem5KPjjMqQtz1yaTaXuLyQ+mKLX+D6
i5hz5/c8t62cSLGur10YKIfASpw5677GNLH//wDQfQm+y5cPjycQ0a+SPoef/++x
Bvf4JElP+976vpKCI1Tn2epD+GBdc/iKI58QqW25Ib0cvyiM2d37lOV9AhNesGI2
/qKuzeumu+F4szATUCITa7uJIbwXxsZPmhyNaNCDUCZB1Y63Xxc7jez1zOU+Gwe9
dn8Dc/t91C48HA0g6L7DuuFQJUeWc3v7pJBi3Uh/ZGhhkM40s94m5OnslEuaZS4r
2H2g0rWYlOPYwrItewN9X+HX0+HHOs3MWMLcJ7DErARaPnJ7FfVeKn523bSGQZ04
pluxg8RmOkAJWSYGQ4pF9+aqpc67djJmNtfWw4Iv3VyWE1k1QLoDt47ECSKY105n
RiVqqT8j1WtZFvrufOiyClHCclUCQtsZzbHfbMx0cN46ZZSms7DmBZx+EZcRVL1I
pyn3nuNd1xCoJ0OnRrFF/5ZtLZpIBc3XXZwdPYmu6M3+j1CFA/vSY0K6QZVLMKPJ
ANuaFXWN4K+e2qo//GgjTGhkTcqUVdqd5P/V4+79B9tlmlviiqCmBr/nMQYDnjpA
UGjuKGDNUGcDPFsj/Y3iI4rMwa1X9stkH0HoIhUsAebhq6TVp2KtU13cw0khcauX
3gWE/YE5mutoSfl67ApDpfQMwuxpXgRmdMPyasHMs2wowEBiWLd0PgSavhdf8sSX
PtJhoHwJtAb1IZN6xMKhjTHPJUb39jKKDZKv7aKy30XghDDqNsmTKRsb4TSp9pUo
A4iUVz9Lac+/4Ul6LY+V3gH3sJ8ZeMXX9/iYx5iBgnuQmEZjZWFMX0koDZcbKNMr
ki8trPOO8PJBFOe0bZwWGYm3YxulApmnGWjtgKCgcWZSXN7BPX5fM/sTSfKOCqWn
7xy1mFfkE+rcOB/lzEOjLlJWllc9pWNT8Cqg5lz/WQfMZgN3yOX0S40zj59V2Cuy
6lsamp4KAG26wiTSP8x1vjBj9Hp6nUg5T3r2ZjQuyG5LeDLOGdFzPxk4qyrQLv/P
l+/Q957cFGcTGUMe4VIaknMJp7xkqXDZzfa5gpsOHOAdD7JO8gBElVd8sHV+cQ9c
AEYje4lqMSAPr91iGSS+GWqpYhc+lZ2aVDCKqow4CUS10YZJcKELuwRaarONKuft
6+hSyUKaHKwoQwbkJ5pgcWMU3YYLtLrCfzvJeCGd24B27Qu2oYKcTxbPFVtD7Ktd
xBWs2m6BfLZXQPY21458EPrBf/dQOJt2kPvvXioeA6iNept5PyyhVm7jUJw0UPZe
tQFhUV0F7znJVsUA7CtMBOgIwwUf/gp6jrKM4akfzKB+UaTE/f/SCCgmKqYAWiKs
vK8R6q381KLr6HykwaFmMj0B9cdHuS4XyQ+4m0Yvy4fYFIwiqfHEcKVwTG5WEHsC
VqhIXU2mXnyFMlfCnTZoHA/VF3nMZcoRki4z2SfwV6SY3CQg+IkeluMO/3V2/OVa
euycAhZMCADp6BCWwph6oXmvcb7+wSv6QNFSANvV43hlH0QEfzNkrKewszdiCueq
6FdqlDTD7d0wGwKn4/SKuZkr2neKT8OTLbHOXDNXyLVzqHw3SB9KC1i8uXy7ObFm
8/v3Z1wCWDgEW1swGQN9q8J2arU3kVpLBGi4zJ4h1pb5eUVnc+NojzhYPEIM3BTf
zrHNMFjOKGEmVcQF9nvhLjnCbb0a3N1TRxhkktlAnNUdIVnD7078IDfiP29jV1zv
KC0sj/S++KfLKnNslh6xzCDWOgn2ANP06s9vxfVha2UKN9fvdzbBcR1mKRcv4vpJ
u9L5VUOBom2VkbRCQ649sLvH2hCjQSZePJ+THHqpr0JUt3PExjhug1bGrTXF/eJT
bneCyK1wgjZsZI/bZijyWk8g19ZHOnQ066vPeoOxSiXrFBPsZmKvlcL7E+jsOhVG
/k57JkbMifyY1iTrhuUqF+CdBlRLQiBtoivQmXX6yinc24ijM+/lV/qC6dgrhyPy
XKKOrZK0S1HmlejsVyFgToOVPzRwJ3NvjfPAAV7NcQggG2hdpjupMN0EhSNuNPBC
NuK7NEOcY1oQqf4rn/7PTYNMOTFiVI5u6NLHoWS37hUrZxoNnt9SwwCA1WBGtUm2
k9KisJmIJv6uzyiqiun1yuBrOGJe7s5BH/GJm3VKsuXVs+WaSNI9klnPiFSjpkqK
UAXZC+ipIhdx+ZcmHZFBtNR8IWDnsDq3X6ufPLvBi7RO1Vk2owRdmLQUHg5Pbn8e
iF/CHC+/H0eg2GqxGEcD3ieCOfix6eaKWEJUo6bjmnjpstQZYcj1FyKSRVMhIe4M
AqZv00HHHXUoYho3W65LoLPESXR7sn5qsF5j6wCDBLguZyPcdryN3ASR963rjoxZ
7+KgEtGp+v41oFWHvESLuByzvBCL54N2GMdztLQhEY+C62S9Cd+gR/YLD174GRnz
MUKdR773IN8TA/Vxcr+wVwPMS7iKRqY4tiUsPoUK5YFrG97YI+2NVyjUIt/hXD1t
AjgGSvg6WvuwMy/O8Z4hop0rR16Ih9AwrlOlNI31znur1deVqa4iCzELdrq4suFd
RxR8QEQS4H0fRZ09RtYMmChPSLGxch3ybLnWjgjdeRyLRBPSs2cQQPNZOU/BDxrX
yJKsQZSxISx8s9e9Wakq7t8T5SskZUPLHxIKCNcUVToQVCGivvgvlJKl+wiqSowi
Z0oPniKP97j368hgTBo3dj+ISps7Q4TXEISjpKVfnP9Vu+2OTWrwYVGpTGOT5eWw
KBuShlaRSUdZ1Ob8c1KsRGe9b21fUVzPoW1Ib6gepUKcN+Pvsm4f1m+i1rGfTxtD
jURbpkg/C6MhAkasZOMezFSSwk02TYUCUF4UvFhnJfr8cqIAT590gczJuicifi9q
FfAtqB+ItKeW7QdPH5W3XzYWH5y+mWYiJcdiEpGr6mV3/NsNrFUK4DIx3lCiPP9E
63NBhDRFQAZfCx+hTkt9F/qdAGoLxZrVI7VlkaOHfdXBg8hT0k3NuabxGQSJcC6/
0gatAWHzTrTPRnvQ/NiLBzcr30xWEMHnGhbTmXx9tJTbVc1qtBVc92Cxec40Bmhn
F/63v5YC6KKddYZUtLrqxuTRiUEh+BZ9HFcJ1RYxZJe06Xfub5cqtOkoqQccC367
aoS952xf5Rerte1gwvsyupLBJiC9ieDNLCkqG97hsHjdYFxIcDEYh25o12GMl9pY
2apgDSPBbcOzPgTvh9g+dm8MmFzUfDVBXFWTsrpZWIWRtepZU62t2Z9HVxEEeP8T
ZFnJ6rkuGSKWT/ForX9tIMiajEa4LPJ5v9lVcZRiWGsWZ+TmBvad/Zrcj1Qv6BSp
DQUnUlYkW/eS26TkLaH6JwYi4Sfwcd/8e/0igYCt8LgvXDbC8bB+nOgX6di9Q1ms
PQ3RTI+7a3fg6hSqWNnyuK5oRawR/APHM0rcfEyqlrZi7GSPGnyY5Kz/pTHUmbcY
g9akPyPALcVWAEQIrTgoIlrmx5XIHAjZdt4SiCmxHEJdlGjATqG2tZYlOOKut+Rg
YNr+915Bz1Ya7JBMEB5pf5uS4+bfxXk/iHhTYJi0cyMZht/xGG0s2I0GU9lWC5sm
3326HCNfNUyRBFxF1P7F9ftYmnfq2U9IQ5MCrTImvyFEHfGdpiq+1YUY8yy4AJmn
GKxEGlgPWgW0AJ1jm7QcMBPm+dcR591thuCqYufwnOYr/zFffySjEHJIguYo63bD
jHagdvGJMGZPEW1kcEQo2b9KnCzHtD/I5/g4shtCNcpwAy/6f8n5CvkL5W8992Gq
StH2Le1TGIKMaysxIHZd7wz2QHgo5jiyaKonX0rUG1IQL5lXy4NukiZXdcwd2IAw
45SELxC6qhiVIg+l9pM+ZuEyyE95rzuyahsTpvWtlzjwAK1kTGplrgiIc6TpKlCX
cd7BSYCU5prDGjEipGNn9sdlvl5AOy/V9pzth5eJsKkMREqvI4eBI5rBgrN99FAy
y5Hf+K4vhkPlwZi0InxTONiv7G1DFSb3WCPMgximX6Nl236scPSQmTb7pgT3xqdh
ONQu98dJFpp+gyWrJe35vKrsV4gsxgcduwRecPHW78nKxuRxBfGflBYp4OJnnWYX
YHEZggXXb1LZLq4JtpBVsXntJN73vnSWLoIffPl/3M9Nu+2TMOQX8SQYD1dC+LR5
OFqmcdoBjzqoVdGeDQGsjwfvoMjhe1jCdQ5qdrNeOFpTdLP0R4xeUG9CYvw3s87Z
7iiyVoOhQ7zOvy3XjHi8/0qrhtQu3X0jqiHfZLx5I3ujOjvdEOAg+fl7FjEhz4jr
j1nUrWnMqkplxURmaxGVv5JNdwD5bthGLwQqJ5JIkG+LkU/NwaMeK0qxMgriqB3H
MQb0IM/AyHNQ2QAd9U1WvzfUx9h4ovl7uF41LxH3kuKcrf3H0ecrdxWQOqnr7C1Q
LaBu2CbVKlDYmJbH5AQvz3yp/VgJDtb0o30Yyytl6KelybMqPvZgmeaWz57pU264
DVMtJMH8HyEpZoH7Oc9O2E/jJGu9yKInHGB9+qmN8hB+crcgq4K9CmqbnUj0dEaA
LriFH6BotMk8fmnVTTlAEwL8Sw2xiww+dsBM5IBWp6CNmX4zS4VQMesaIGSQcTpU
y5IVErNq3hyCd0Qxh6fQpKo3esstt1Ec1Qo+xIkUG/3QFt1JVczsPzCWVcFbS3Po
IJaGOGLOoSUUWK+VNAaMDjFMOzGtQChAyoMI211dZqd7q7VrtaXB7ntpytcYhSYb
frgGH+AkuVfIeFZ3uo4vt2T0didKg30Zhet22fPHelDogyER0Ad9dunRlSObCGMf
+gXMLLul6K+cUFrGBp0Bxpmz32Nh5vv0wdp3va7bSoTapq4wO5X/qeTUNacQX5qk
dHyMbrLR6ecGujEfZcjnGcb4+okFEO2cP3AGJE9OegdJ2lmttc+GdFle1ABsRCyG
D3DRJ4f6ovO0zd24x8in0rITgNHL3F3ULpceSy3Wl7we3y5qB9HAdlb+2FA/pCiG
o4p6smay50wL+XRhQc1guQHWnii7aWbQ+S9aQ390DGfAagnyJ9Bz1eWGOD+2bKQk
HiLa4mxNX5SItz4r14Pte0Jsq3XWyCyw5Iq8CVlXL2+wRyGBjUVippHqKUD4FElJ
OdrkOeH5LPzJwaG1Eso6Fci7SjAHMYcyfblZMTTdwLoH/J2uIFgiFIVOExw7CoSI
Vj9z5CMf06hMc+gE19fuOb3EOQVw9zjB8pYAFT5Z/5GkOQd1yqEngeJ2prXDWgB/
ufFYF63Q1uhiDFLRNu0DHoeqLO5kp05D6H37ZtdjANc8L5Oq9RhWUgE6s2UtKgrA
lBwS+yJ820b8TfFkd6CkQje3L1hnEk9z9WMZdY+GEJED/ko/1vZW/gT9bTAOCocB
y8pCLLH9S90QcDtKDkp20cQS9+THuRFvKlsHlS2M1loS/1uVAAwbS75RkVbZaiS/
ujO6xXMHXoSo/L2E2gK2uUOn240OFSENzbZVc+5131NtnNAKE1DWF9560fqDzia5
4IvXH2p+NoOmNLXQwf/mEJTmcPTFG6CNvta4bb02KC7RjpQqvkFPF9YbyAi67RlI
BL7LB5/0++rXF+0NdH8dXJcOHc41WDXidbWyocFpd+gs932LfpIO8X1FzYTAhEof
0rnGEfQdeQvHrkE8hZjF88ioJZQzRDvLuPHetAmbmF2hb85aIjaMCDx4tsCc8K1Q
y+TQrXr+ErWZH1MGkdGKzzFSVmQEyDuJZKQ71SN25R3+GTVnuMCqGF8inmnS+7h7
WH5gD32thS6dFJO0h1Gl8mCINtpUOOxlbwQpuorShTfl6BiyCXBN/Z1o/FDD3IR5
C7cC/uVqVk/vhwmspjSsLxTDknkk2ZcBefbVr1rknm1ijGt0nYVWTbJ3RdA/rp7v
ZQLrJ/7z18DEM9efsg3I9DtzezUovCG/T8cY29T+nEqXNk+7KMlbkvZC2eKtahx4
Dfv1p1XPjWLBMrVJsG2YNEaOcz3cFvO8ZKv8h33PdhLvevdUqcRFJtOdd1+UuD+8
uxIYwZJs/7vK+dkjTvjI7NfheO8jJlGvG5/FVJKD/tmhmrvxD6zub38sCjbsFQZu
XTHGZatfwjamzqq+ISERA7cR2BRrjB/5/6CwdbIcHskvzJjtGFpvrk5MecRkUwJD
cFgbXLl6p0kas07vimy7n3EizzJetnspWTD15PstVZBQ/w2gRdhUOUDLV51rJuzC
KslABkQGR0GsLFCHgA5glINnW8CSMe6UixZ9MMFSrdDCb3ywdUvqcqlU53sBPj9E
Niv35wP3a/KT7e34wLBWa8/NCPyuq3qqhbIqnnOnSTLWBjcK9uTbr5YTUJXqro/Z
NkOeoZvI/UjEir2gliTehPBuemuxq0KAMVj+MGlYjbXraZd+AS5CYoCaymxZKbwI
OmIhtbcwWGpUdLOatS/XLSX3S9iIsRcQ4inDls0bk4Gi4tpkgWz/XpGix1FO/Mal
dWJrDfYIze42di0tzxZtPi+o+PXzGN+s0bWMuFrnJtqlhliVZjUEGjCCWA/4gm1r
p2m83ITgrAx2CNkysOskd3s9HgKAbcZPFZsgjyAr5PtbjjXGkn89KFP/SGe13DGy
szXNg0KBZ7FPJ2vRX7gIshol0VR3ZR2lBs71RBaN2cdTscc7G2wsQ92cvzbF8spQ
DPsTCcTYrdZ00FoxPEjIdU5Cjk9p8eyCI2Ohqi5IYsw4ytqETKRaX3bmXV2magJb
yZmaB5JoZNah20vkzJKTmHkXBrmWsf3GkxPlzQnmx8gPIeKQ9g4FJC9b1PHjGHpf
lHX1M/hrALZtZmTYk4LstnAZidr+ADhkFictktYL2X3V+sPouHZnu2e2932Brt2E
cXD9zxpfqAYiufCQrN/6Rckb5591798NaYWTFs1expjArYv8DuJ7+LFjdD9xPYg2
DlmpLvsan5yjcORgDNYCHlkPAzOOHKkjcLY+9FO79NUjsau9YZH7c60dmyGsNIns
SQuNFpfUOevBufxNW9xlOT0aq4fxLoEu53E9v4HEQbpHNqS7nJ5WM7bfWN+0ghTS
etH75p7XKGqaM3X/jWULiQZrHJtqotMxr/g5CD4Hc9Nmmlk4U+tHhX3hCEQTwdNL
BjJhXkmpTjwr/XH8ywE2In+W7ZrIwUqPNDfbEyJME6tEV6LjvI7A7eaDRKPPcUr+
M24ZET/jbVebMetQbavZM8S0VOUe9FO7fJfHn5RAOLmS7xUny/AMmDzACGycTLhl
RwAwfimUsc93wSg4pOeB01jkC08lkPQrwZASiEQbD0Qsnvi7gh/D245gHzsv4a9d
Ne71suF+BRSfp/KFcM45YneFGh5c4XLz8cbbzJDFlx4TBWDw/r8N8UqvaTyboBV1
C4vh7Ma8Q6JrGqgPgtzQak7Bv2UQKnFcAMhQs7iUY29Po20b++o71diGW9k/lT1j
c14xtCQ+8jvNEunhxIx8RrA8v4Ng4rtypmIyPR2Snl8PCN4HjSc7EFAPHBaDc5x8
oWm1RR4ZlCKRG7zp0GANNzYn5pES7df1kZ3si2OHF7ylrbij49tmCbNlpig6t+XO
YJ8Yxpyo2K6JjDK6uzn9M9DBx8IOF15HKkvAmzbzpIbpC1Hm7ElTH7krwuYUYvqa
GrdEldQGC9/0AttBCnaOjv9MeOFSajcNnlqK0EGQajyzrxhMJkw1s+kkCxz6D9F2
KmMtULIAg3TJNdIeceQrAWJtf/UpgVVKKp2+88ZymIF/YQjR46ofXmS8xAuQXOeO
cDHxNXfedZwteTXiI6CFLLCnH/uTx4K9iWW5ea7V5zLCf/VvW5nCUxWJ+ZDokJXA
xk7HhyC0g9nJTLoW2cQkl8k8LWV30gbKyZUihqQ4lgvWBT2g8Sa0BAZ9PkKyKLts
9pzdcSyIw50YhtN2rAx2gl8cJX7OVzVs9uBi5RWmQi4uow65LNsDDRPL3vrR0BSq
k5pSwxVxk1ugekHS/P7/Z2LPvD3/NRbRdAC2eENxOukaM0Mta1ykz8z+5AtSREct
Rk3hTo1EmwWE88DaQo13ipjJHQJX4pK/GZB0tCsLS+/J6JoamYMnuLW1Pine0Z7x
ulmk8168fuQ6Xet59UezwgX3HmIhG3KAv88bHvt7Jrb84+184b2KOx1hwUWUnxTn
OvxP+Upo1GM5CDg25El5jtIfamAFfmpaFRAIpOJVcFL8DUdo8HmhApKYwsQ3jUVo
1VJr0N4GOpGtwcFJp09WDN+6nFunOBapRvQ+4R5uFG5rpF7QSNLrdK/vSDjbo1Vw
JCTF76A5y6SujcHhrWi6WpGykpVXclaFSShrmxjkS5fPHlVLHTbdATsASvHy+fAt
d+LQzZB+APfxyFxKvPxiv2ABqlxqIG0rpdJXu4G0uo791w30s3TvX5fCpl45ofW2
E+HXlOZ4i2Q7Sr7TywAU+SQlBnTWBJzTl8hEkyBORjmwxpna+7HtaYq5D23I2rkK
DPHYRHr8ZOBxnH211Odzu95spGp2EoQOrfWO/wp7IkKwrQaI9T8vnBklYY0cxF+l
ImBB3NiRhrPKf3sRn7K8GW0P+g4j1+Mn0O0cyrEK2YOwu2AD/TzPDSPFZd3hEEEE
AMB66c8gsLyiFYkXnA4bUjXTysyKNhyV2Z+4rGgFHKJqjSp2k42yCsSr3oNNR1j7
Xu/vitwl7CVLGRZiIypffOPA/1jvbFLVZbzrKn69JYK5U9Bs94eIaHuYo4hJX8jQ
geA9xiCggn6eJrY4hs9zjzZNPimLqjnvSR9vKrQi3CfJpliKIzAC6MKLumoVPPSB
/+SzWRo4ZZFCjodXYYVVZ2+AKLRMuvvtz58Dsb4iuiHqVxyXvPS1uURDTdId2J2P
cTGIV8I79JSa8R1V8Fno1FEvn9nZ7t3KhSr003NhZQqeyzfvdWxpYw1a/5qhliTj
hUnbbzsKqc2fOicyp5qpu+tByY0L8Ro4B0Auuz3eGqoCl4xNQurFfv9w8AmjzI4o
i3ubelw3EDrrL4PROCUZ4/bhQQbJVu0H4vwauJTQQb0UM5vHfzbrht2lciuwhaXf
mQBnt+coevYeFht9WkI3mebzthlG6pJjCJ5c6SAIiTBAbbwbeM3N/LOXeNwvsJL2
JSauoroox42bMoa4SBQg9oqzyRScplufnhQmDmb9Nma0nzllAK4bba1RbhOD/aTH
Es60ADzgFz/xYZ/F0fO3p8yUAHZCKVKz3+yjElLAPUz8XN8D/B6geVVFFKvWn2wJ
tI9uwK1XcuH7u5Wrvo6ZWBRozmFQKQj4JRP1fh4zIZ7nPo/GmbFJ3Zqs9VgFd3q1
Ks0PjdoIbXxdC9xhLkQhMB6WLWECXa2Xu4fvZN0MnzLMnTCzqYdNli6PlYLwzH8+
rqadLKl93cqYLDG7vF9YicNtxlK9QVetHdFBNbTQFrrNQOEjF+nLUdshQpvXUnLW
68zhQbGLUq+/rIhbqFpsvEQcYfyk42c69BpOHY2t1OleQ+fWBsHnk8rbNwEFw5gi
rg3chzVhu6vupn5CArh28oFxbpzlrXrWlQhAJPHlIVuxJwz3nHlEC3N0xYGSK1yo
e4zJ5uN9fXqh5ERSjy5lBqZZCvsTmSC38Rf9tftRvDfnLhFoocqHrkF2IDmGkdJI
ifUsuIPIq9JPypD8NAtiKPBjq3/o/Z8FD4WRrAJ88ixJfcn+3QP3o1rUKoBzMY+0
bjlI8C0cSWpSqvwqx5LcJbbqU6Ed8cloHwQUM/Ar4WcS1XTc5okdvjMydtbgzBNh
HEvjKCx+zMcwXC0lu8txb3jruPALD3Lr93ypFp54+XasT8Alln1/MLvXynwqDzrc
vNjubxLTJltWqGlRJwkGXJioWZzS0xjt1J5mPN3XMKFeVzNQ8yBrqsee4t5JFMGa
dEHjUSwsDX3bg3mGtNIlHXUoM0vGFVtEbmwPAUapeKpxguKty2BRtyJ/ELtNQPnC
h6I0WGqR7h5KfI4M2hrfW1PwM3HCwGjT5FwP5NiZJ8gCJenb2L3FLNxr7tP5Xbd8
7kFwA+t2xXGZzcfhDQjjQXrKHGpxHDftgUn/G2YCqdCVEuVKSKaDYUVnMuQxuxil
j+2pip/uf66cV7IP5VquYkSamOzjUPRVEAmE8ysFC5R3MVJ8OYsCDWFN58mboc1Z
Q9qLvQGIJYYJhUi0wL6AUB2GMNVkSqlQUFD7eHYIKqyqbL5scqFX2ikjx8MsjLZ8
yV93HCcnTpDLqfmWJK2etGg7XOG7Ap5vi6s14MrptFcnHQgRFYLZ9DSxR5/tWd2v
4xbYDTszD9pdgf71WMl/2WeqvAAXxRWu5I2CpPig9+fQDl/R6co49L+qR3cb9cmN
sWYvJepzrDpwM3m+aosV6S4C+qtCwQOn4/W0Jd9TRRyEkftCY7DuLMJ4gVdDO/cC
896Q9lpEvAAnepNOjQXCPImCKI2XHhiDlY5sJ4WPNPb9E3pnzGqaG9lc4y9mHYox
BW4383gAGqLe4F/0n7kXK26eFaq6ckm9ps/Jsts/DSiDhKUziZMlbMj4iYmg85Tr
qgXUGp/xE+rbhBW1EH332PIKHRbAEd+U5NuWB224dY3I+jmnsiwBm74SVWhDJ7s2
gE/4PMpqvrMTG+jg/EfoXUpAMqVsF6se7pMIekBe51jACU598gsz2Nem5kPoDKfG
1QiL2tgwhWcC+rqJs3risMis3qyW7/c1GCfm6HNMQ5OxsVB6tYiNszIfNrSSUrE2
QNJ7PYjLhBrcizjNSASFh1vog0qhR2yNyp+mKG0dNYNmBkTObtzRODV0OLjngpiK
fIs89uPwJJ1qzltrAej2H9W9HKd3TSeEibLwEYt+WvHYjTN3u+F0NgrTfah2GtBB
uxPWk/rRTHmDYmF9FASJe5U5xhd9TZso2P8hJwGH+4SX81J0sKKZX3rRNUKCxPE3
eQN11pa5qkDU5pmNfTrfe5Agagh9Nht/8tsiPF6ivYMi4Y6bAc5QYqHl5N5SzQ++
AxJzUXegLqodOTUDdDi4UzRo5K5ZfH6OfrVzoX3dD6Xxg3/3yTwzLWuzIuQL+noP
ehBtleYi8kzxnTmWupMOEF1+QT33LFHNX6PYtBV0ZCVP5imEvu4ZgBn4mP2JuoVc
VNNFGnFnankjFnUkBQVhFHoj6MXUdX4/Toa5AtS7aOuKwR45d53LpFaj6jANwcj1
IJI2BSZIKNeCojwYqwxGeNP2EnkP4XWEtmGhXohBDpiBH0AGsJn1t6CAlU4WmoMc
RJdHtiRiqENPkaKf2gaYFocDUd3v9wQFbKNx2i2Ob/PRjZ/17xip7kCqzccmCL5U
XzyMF0EBFrxisQ8M/+ETVonLRTtFENOIWPGbGKmSjih3CsqP3cRaLJzXabO0ZcJY
V7IzOy88MhnwZxIQwjlLuIeNYXRHXYNvFejCUbIWHdUxcbL23pQnccysa2kdYDQL
Y2rSYdftmHAPga49YCTMi5O5WxtgoS7w3pTaaGPmRSKcnYaZhissaaRcjJktn8uv
ZN5ePVi2CbWqkNj3ROLwpijOea3+7R2g97z1B68kg4bcCwWkASOwRB5vW83FoeBd
72zwUk6zY4k7/PS3i/H84O2hYVv+ifgeOJaod7UDVh0oQio9nut0q9CnR8VPBsKp
YDuMXckGs98X3vdsfYErscvl8MaVbFhFGr9pELSApuoToU4NE0XTzmSyd8qJ8ePK
kIOk5f7DuHcT4SMjbKUPn2uxeDp5/OCBDiiwB8n62HdFqQzJ1Vbtz0EQp4cQ11t1
kytCxQw3j9BqyJBDhJTmZYxC6eUr233XKvwVhyv6SfUkQo8Z23YW16Y8v+wA3EqB
JzQ/mNnrDkjdNOd8hOlKU/F+XCD+MsEae05lmhft3iH37YRo+KtKrRjhy9oLAQj3
6aV4a+Hi9HSdQ5cDqJhe1cnjyUevBEmQAeoUbZY1cop0LXGgXKvDB0QVSpbBRvLk
U/HGTXZmwHTPXPytTcgpG1eW32z3TSwTbab+OjhTh/EJmYtBYzzTpTJbfupoaNfn
/VVgjLGxQtl7DOY7TkKO9PxvDB6jTaTIGpNmeJirc3O+BB62+4L0iToCymQAzuWN
pw2PA5YRP+p/UkSUi/ArTYjkm2z8lRg1/4WHf+ljTu6ybSyJLP5wgo7OIa7MtlFz
Co1IbuFoSOQQa+JVTGIVg3aCcdY1ktR+vyMbkSEBdiCv8EpTCgman3hcvudX+dv2
Cj4V2OUL18vE0aW+R0MewTltOQhQQUrz8FuxyxLUavNAUfvw7tV5m1YoeJFO0pP4
fb1RBZC8tFGnfpG7JP8C94osUL9IXOGD9Y6+M9Ga4E3Hx3XVXQqrwScypDrsktD9
9AdeQ0K4g/MXiUHSuCj3/lRKYKjjmSCrK6kOlzI/4Xiyl/P6rhA5hpo9yE77lQ7O
ar0s0BwObn7eq856GRJFPGkSphRHtVtxEYri+FQr3eLB8NfOawbDc57ThI1VsiJB
9JQAl+n6xlKFaZtkcr5qyssRWMNbg6WpugUL8VCo5UBsd+KI2r/e+VK6Jwth0/b9
dpv6RQGCjA3ViFnmfgJs/nEi7K3a3+yLv9GpF0dCK7ftYuHqN6y3lLNFPgqKKQFp
M7V11tiXijOpo/WQQGtuAHEkEkBmzkjwd9B/FcBPmc30JmVeIf5gMY2CW8RY1eHB
dnbJApVikzaFO/BNaBm3962Ldhp7X1GGRO7qDqVZKvNPEOWENSVmDaEwWpjrVbyG
V1DSZ4iTZkq/oDzmD8QIHPNoz0XOGf7MPtPm7NShL08ju/r450MRs3gQxQX4p2lv
u9r5HvpPrGwvO/a989njJIQNKQC7AnF9cWr/ArtaP/bzuCdZ4C9xkLdkMZBD1Fdm
LFV4I3hYnjUmnjXuSGIpXBb3fpzY0N+vENfg98Achze8sfgDyD/3TeQ5lBI440sg
Z/XGS9w2uXg2i0ElJcTA0SCqzpVamtYHhC6EfpfaQjWo8YBWRMtZ6evrrr7FICox
et1/2w2U2Mcp/5oNLDIStZoNqD2sY+iTt4Z7QYqduksg3UaB6VQxl6/pP6JRwNCL
V74pJTuD95u98IPUiq0uYafapnLjn+l2OJK3qzgLft1d9Zzw4XKTkm36gXp8vnXF
oJm2cXXwGMW9PpOXzj4D+G+PpdQoKqK4iH0Sb2HXNKMdph0K3KGkQ2FKHh3MXAcQ
yOPM4+KFC3MZetunJUsnyuWOUPjWcT/W+EPAbBmM5NDzoaRoMU9iAACu8GjkHws0
HzjchE5bB3RSUNOJcl44ggIEpl6VAKnRx9S8hE7kwwRlvOByZ5DhNgGGHf3dT1hw
2b60OWi2Ot2dfbl3mkq8kL91ujsOVcEDJbvpg889VicQ/6ue9LxBzCDndOfQ0viB
YsZ9LS6ycxzeiDGK3NWlVo75tTwSBtIcVKAIa3N5W9WNb/hSqYuGi2P7XLDeIDei
Oza5jy01WIo401en1aOXg4z4Q2tfh0TA/UKfp1gmylEanzfawLAKbdVLA9NPYmnX
ya/AyYI6Xdj7288hrNRPP5ftZz6WrxyioBZVbn/gjSN9hiQ/jG1Nqbnnq3e+v+bR
mkg4DVJ8mi2kupg3/yYjyzQsFUGDab1V1tWtzAqWuJJlI01sf0ElnMVmAgDUPgSQ
e2hS4D2VI96ho08vS+IDcoGg4vjDNF8SmnRG+CzXEHDqKY+0x2HFCJhESUvyFS44
OWo1RC6k1mdgYnktUCt6X405qyj3AbeTAQqvEoiXhWHQZddk9ms9j7rxq4xFyH8O
XjD+ZMWENaH9VjtATqA3sijJFpacwrheEVpBGRu5CJ8cUrdeKDUnjbLdOs3cK0Gr
FIhDHKjtwcSy23FTSUD6mi582j6qSyaaZJNhlQHgH3LP2e+KpFCNvuq3cIOFugfW
qUZZJRDbSqpoER348LnqFMDm749aKEBABloiqPmLWr8ehqKLdMOAqjdZUSPAB9WI
pFf6/st+1zNPiU3gWduE7Bezs5wk62lcwE4JBObF3f3lO48OtaIMe31V3AA692Zq
f2njocmeCKdSaKpWo8fCBybdYnnYdYWvR8H6gSjGitnvLqj6lIC2TV4Ye6pQsgZM
IzDIWM+OgdlG0UOvr7LzORAYqG2nOCmxADLHo9+HTkKMfywoQsX0En0yvQLpcjCd
gAjLH+iskyF24gFEdNqyiueKWpmxSxDxVoiWDVPGwkH3Z71vKFmCloSCSEUk3aE1
8nNd4ADAxrTmsfXrZcdPTvigD3aiDGvtoUJ7h4U11BQKpwVTzuy1xUcoGlMXZTlJ
sD0D3guhH5xOgsCCkgfU0v4BP2t/+OuCG+5El1jP11cizM8BiC/PTbeRDiZVYYSe
ARPN8blYigLNHgdCLB/kRn03hspUXXToPj/uMR0o/zpqeRYKjY7KU4oiZ/2zwt9J
SoFvYwDNC5oyuKKPQxIZbQ/+Xki3FxU+mAD5Qt8tPs3y4Mh/iRubBvcaEp4EBn88
e/l4WPYamxtfA1YKNXytOlDTJVpZ9DaQa/n0s9PPEJMOZcpm7VJutyAkYXb/sbz7
zHFXKLduAqF1KHtiikBRZARUaFmO4m7POz3tc3U0mNlnjpzwJjFnQllFAR30FBOi
V668aGvodd4qJrtp47htx2Hp9IJ7vtYe1QZbtaXJVpQZNHfxH9VkH1LudDpnB2FB
fKt5Ml9s4t2bJTYQAZGOLLh95xIzhmdlfPyM9gI6AARvaX1Lss3H/fH1gKIuhHzf
rKA2sT1rGKRGxNm20ieO1eIW3a6jiQXazTquDOc2jbmDPmq9ZU8bbWRL6nHmZ8D7
aTEmf7iNZCrfSZFw0/hNQOMO1D+68yb3FTP0sSaKm5do0CCb5KtuFX2pl9y1si8i
nxA7zNQ6eyKmGtr2qmIG87UiM2vaA7+37bnWn878lJmJ+z9bOrfnaZLjBr42EV2x
NhvgqKViGxUWdqsgs9JrW5X2JyXMtnSeUqXzSsMvAQHmm/p3iLx1koz8fAYSa38y
/jpderRistsx/Cn7Oq2IZVskDm3cQe0CzCokX+j5fiIPnfwYlgbisB3G/1tlzZ7Q
tjb7aNxLYEZVkkNUO2SZyRN3rjdDa0dvUmpMAdJO2zCtVaD5aBCwQ2VV2RnwfgmX
AneojhGLkNwh7/0H/ifqS3XzCt+USdxxwwBYrzZF9pwhLNtidwcz/zygzNdsQFAo
mOoct89g2EPXEDCagYGa6Fs62BW0jUKbNY+NdKjToWrv6XHtfKhKf52m4/5UiAke
atcAkGUrxA2bhhv9tryev60NYWgE0gef60UOqbPvPTOZ4kNvTZrWTyNrppLIOzQ4
YfJORcHZ0Yp/1X6AaALNNCygcOojXNCU6NqP6Khy2cvX6Zppz6uO1uJ9A1Y+LaUH
aK9o/fUKtPWVvm4L/C7uSgxHvWnQXEaMijPlZnHx+L2b7Jn+pvqDBE85yTpo5HGA
HL4kWliAKpgp2oFqeMuQXwwufN1NfmPlofeU9WSLGfqPUfMSWYHmSvBcJcMMFkLJ
g183xbBT/ywbY1/fvknVLwFhgyC9vlDSZ4Q/GIUNrL8FXg+CQx9Fxuroulc8cLWr
iyjGi2os0vRHBJiGuFIh577T9mBEDUoPrcwZ1XRebu3BxO/+AW6BpYUtCnU7Dbnl
kt8qzJjJb2zPGIQGk54S/dmNdpGWlGGXNqubR9lDv6ns0EJSfTdA7czJi6eXpkdt
LTWs4ro6y4VW16aot3z9g1zdJcVL5xZpl1KPPA2kcLJ8KbuzZRIcy2kEDDtz0Xvn
s/u3awh3E7k7HjKSMYi2jtxoRxNLtfpDYwlnvluJAzpd4pRy7K4JgfuynL/JK1YS
MZfGOn7cuiI3P/VXbve1AYjP1//oyhkeL/bcUKGp1dNvCijxbl6ayQLBtySIaxlD
mxyuAKUM8oKLIuk/zMBxkhPDvHSORlhe5hXARTxK/pdJDpo8RTRdo+SLQEpSJ88p
gRUQgj1GkAC8NZct6+57Hj25zQBQ3Cuvc6SqxLJRt+uNURt3Gushp1ihKsKGe8BQ
Onxh+Ys+a4gVtT81IfSDeSHakF5/kRLSUYJyYjwunLREVYD4hqr7gQYkF5/FwB0o
s9wV4iDli0McZVmUB27nRjfPbWeJhaJgEKeMesP/HuVXqN9pWv2ipEfA9WoRiAy7
XBgyNeysOyyrKsjiQ8fMKwW+y5dAMpMlRD8PqQZGg5LVxam4pE3a7d25jCyIF3A0
QWp2tUTuLTDWyWmPRGv24/OMUGbiOVadUFAqROHpC557aRtBixJYkK7elx7SMZq9
G8V7GRzHsVCobOL64zuHV2VhyLMwYNJFlHncUlMMDNacquCcHK0I8B/T2FP9o4jN
X9B1YeCQSAqX0Q5D5ywc0DohY1ltln1u1N91LnhJKSleMVKJze1UqoRgdQPKwdFQ
UpNzw88DTwESrVgoFTDaKPFVYmN3p2PIOWFKtSUju5f3m2fohbRXFpyjUjU1VJZk
NENAcDbwtLqDPOpIIqv9aOQhYFSkff/50JSmLpzoLjGHjIqmFQ7IG7xqa+odPZnZ
loV6x/oJD1Pj97xW6npWwv9kMK70INqKD2nDG3/mvzSUBUzKNEad8S4Vxtr4ed7J
Kuq8Vl/+yKuulrlsuDzEy55Lk45fZ0BgR/Nq4rAeD/XCsYjqvt4jFw0CeX5WwrDj
kSskxSZD1Jel1Wxfnn38z/mmWBblH1nn0EnkaB81rHICMETdXFp0sFAdX7qTYfTa
JItjd7S/lqjTIHIILbaGIWL4To+xpjRCieoQh799hMiled/Vsz7JjMM4vK3bZFzn
DQM2GMUZILK4r2bLEyqQUi4aSaPe6Gpw3rqbVYxV65DWUqwbz4eZhgAbZ6Du/Ik/
H1pvEQ3FUelsrGbBLOVXnKEuxB36UxcvHxxFyqnOztygaTIPnWzVbg+k55lsOoYO
sff/DaI+zfgacSrY91s/SdxuYq1+dV2hO//Mn6C6akXS4CR74DDaU3peCaS6zdqr
JPfcj3vUPYpVJtnYhiYBxq8SidlqfWoHpdkRTEbch5PaJKqpeXfuA3Iq4roaAazt
7fDonioIVidFxWY99q8jNYIU81RY/vC+VyPwKYibchKJlClNHy3YS77U5DGira7a
zmXccwnMIueSI+h8g+sXLXauo+SGzLvMadAMK7t/z0+nswhLpbXSeY1WPLEDsXyM
Gexq0Yn//5lkUwNeorGFV/5JqxW1mGa74ulXIgdghxRnjFvUlOVDnxCN7MtfFgTe
eujD3t2d872yesykjZo9v1Zaz1xFPW6bvYar02Ka4TNQCX6DGaNYjjcWPYi14wtl
nPYMyHhN4gCmZhawRZOnNlE0B3QPr9pn/uSTGCFCHgZ/CT1bOkRoc1qezXqorDSi
eN3m92+8l7Em8XJ6PIWVc8g8EBV6lEgh+ZMSMLPRT9dpV7FT7XxWHm/iAwUbsN06
mu5WDK9yd8sheQIDmBOpns7VD4NB/CxXMf+ADrCIxm8o9ujwjKoj3ejXYI5OeaqM
XqJ96y69t8b9qWvvV+3ND+YssrJhHZF0GY3IpOM9yzw/+s3Hdj4jE743oTu8zYZq
pYF42eccdQpQWczkfttf/6Hd1WNTu8Wy+05KbE3UOfQxSBN0CofQF/TC0f8XuJRw
7dgG+yzwyXaAq0ZL/Mt3aspWaTDi+8tljoQCfQ2sf2SDsG67SmBEGc+ArxKbRTUC
0wnauXpM/85iU27eDyKY0zF+G+dF9K7c8ejOhbgTi+m0h4nb070d7tAj9CVkbolh
/jVNxRtBeWKbC2F1C5xiGq2d44MLFy5E/qRelQj41St8o6dz7IVwkvCJ2/rwz+E7
RxrIXOroi4L+N+90Hlu8TY2jx4dGqziLXxaP91EnUOhll0HElTWHyByPgKFcFbcl
LcFOJwp+QMiFLgRjdeR/dsKawINy+/7Bfi1MRZra885u+B7gQB8GK1n92TmS5PSG
gsF16cfLhwG9PKl69FfnJHIdlfuzFQChkXFOE3i/en9cr/ylet8FETsDztPt7YeP
L52EmLtq/SYLw6m+ti2c/a3ITcDjxcdR/ziRywUIN8mPCbBJ9s+8pfkGyxp1trrL
jMxEYRSbhrxxcs9e5pK8QwzJw7YGNxKfECyUJFdMGNScZyEVYNr85yQF6Gcqv5DX
cTlWGZhTB5j++iouSQeAhgFBlXO1B2BFUoADd7MZNfsi+gMQgyuOdyo0gX88aGZK
/AR+wzBiKYWZfVY1XTZ5Uffcpr7Nd2euvgWImPBntv27ucb8fyshGtdZDQlGlFtz
J5TKZG5RiMrEl8oh0DYcz8YHlhJ5NPN5InKvHDuPddU5KQ4a/1Z8UOZyY+iffenr
vZavL7diTFkV7GtZ2158ezL36ZO44SIXcco2doQNIS3IhgzYvVZ4LfPgrQHT0Gfa
GmYXOCmVfx2SmUEWzszeVxGpHt/opZSm/Ya3k2T7Jk2Mx+Oy0ywnwLFnsRk4KHck
22oDiHT2Evphtlgao0qnpO4Zjua/bZLDMkO+aXW3nfwOqWrNqxvK7tTH2PtVDvrh
r7paBOQFNU59n2EshbA5nlvL5pHxjqPPxjmhBO5Uh/F1r8asuAVRmtiZHdtAHNrD
hfsGnUyKKrhIAXRks28LqXUd/1RGJytPSKXmZtb0ycUTjbQH+7GPt7muJtuXhd/N
+quEzaPUBU/xhpw4K3X4TXgwg8SnI5FdbOTSCIGaFuwoDhM4aNZFl4eD+eieA8AA
dTuWHSibtkADvYw53ceJ/sb5pio/4mw6eKWUTqr3YtmV1KkAKqN16AbXm8qlYtMH
nnO0rVwqUo8c/G5QGK7CGrsXQQp8+uXZ2kYLFuqWzdr3w9iW9CA/0znjbc7jg3Ll
hrJFzaqeZf+r21ivp/MOl92v+0Qj6FPxRbYxTrUmNbykmz8HYLnNrghCXwonZTEi
2dqDBoq+zHwMhjTfqSXYBBOyGpl7B4c/EbzWlrtEzOiRHAvsWX1ILzfRNfON6ScA
ymm4xyDR9elsfPy9jZIMxr7szl3owKt7msWxluciubw7RTwUldtrJSN9Pkj4I2zq
MudN2fRPuoTyxca6jvrCA5K3Iw2qHsU2a9DqYen7zW3bOGhz/LHHd5GDeIsYf39i
1JbSAMAocdwbUzRMGSo+aFJUjbghOFy7TN4OQh9hlx5K7fZ5cuoX4nQ8d5KrHICc
YfBJhv8V+wM7Tk9FCZjhCQlXsUtg/gSqwnny5+kT7CV+Pe686OKo+rj4Tu+mPg7N
ydEerGMJfp9F0jf6XcGAWvsQF836EIEyzD3IW9NjErv6wLi2TAiipyakdKUKCqjB
WBy83KeI4hnq1Gq10xVzc1jvtDuyh9ZEBg33b4yTDgUYjrWYK7UyS+BdAcPF20Wi
iv21OXAveYhicUZ91TSf/Kz0LF8GudItGZAqPBwfAwT0oFxD65zgPWwjTBnmKsCO
aHIteAcwF3waPnqepGcjbVBpKjvG0p/IYaGk0jTNY46bKZOFw9SOx8JKrTIth1Ej
aj6oaTUGzHgEcxnkGoT//SnJxcBnsQayhIN0NaWHhnyyDZp1oOUR8DzF1WE3dzep
3eBiVG+Va0aPfUU6TeXUov+l8F0DuPKSNA4baqmmac56CqxU/76D4gfT4b44lo2I
XXliWnR2nVq/yh9xgjCO7+Mb3GVQNTKtQGLFjpXJUmfmyTH/j6BOoB9VU8RulkZc
MDXRKpFSX64lcbgax+yRnwjoIVpDtfSjoyNIjKfXFQkXmx8IioL/NmnMqHC22V+H
iH3Z+L2coKZ0j1I58LXC59LhOEz2RMH6fPBCQSxfdpDBDA5NtSPPV3kWnoo5m2kS
bVWLsjsDulK9FC01XHST3BeM8jxmvzOm6MlGKZVU/IG36Cba5a0AVEyDcnHWBQVN
TG0In8auw11pn2qgVLsGEdz+jIBlusSMthAO+O4ymF+Wxx2qh8SnMdhMfYZWGJqG
isFA0zWMsUz5ywJSJ4t6PoLCc3MfX0ZugftQB7Qr/KpMzydbAmZIA500az4QDv/K
e4AXphbMQj4JfIRnajIXUfFFodcXv/A/6AV9x7kvg1uw4NSWJ5ndKw0WRqedkSGt
plv+m3J6RPLajytlF1oO7/5Eb2f3cg0c+C2/mpT+bC4vTzB/V62LQ2DMNXB+7l6d
tG4mXNl4f0zTjFgre9IR4+Hm10Y9A3SbYoq6UQgJNWrkpgHnMyTe42oyiNLAcpiZ
8P9PTwyJucj9/KV46HmikhbOQ69q3NV5dcMf5d0RvuuIgFhPFJxBEUVd2neH6GmF
NfFYLZ54S2nfdmw4xRz/9YuVQPa2AEiI+QKL9i15LplBHr2OMSwCM3YaAsPfl6k2
UQJ5UVPmVsb4+j6AK0yx6nxFDSCtreG2qzBDPpXF8r+v1uIk4y0akLMkVp8Uzp6t
iphcNAdbZoRjOVpijVF2td21391/oJRfMk8PzcxTdknmGAcGO5P1GAPA0SlfQqoQ
jkAtSqOqBI8QRYWaLuVMy9GgGe6IaI6fgEe9PpelOw+YTzSj+smZ4xZ3tiVWltlF
xYQz3RyUxbDzFGGrIfIJ3pz9eA1irib/st+r07SBYkjicC+kwx3HXU7GLKIAMOtE
X0XYGKvd8RrMjBlBu0eH4e8MuOhJCJdPgc7aVjr5Kk19CfW+cFxjh88ovgMMA9c1
4TuH1lxFMwEx+XvgiGxa6JNJwNUc0wiVJbH5wV3nC/I3HbQw6dp2IGVc3bOMSpU5
SVQ8LMjyrlZT0d8qrubtss1NNLIvJtxlpYteHQTSniyJXi/99L3emRPMYTBG9Hjp
AtFkxjPQYKwAE0pSFLFIxnEzOjXTSy+/K9/sZY5C/BkfSbGwet98IWYwmj256Emo
q+qBmBD9X6PzEa1Oss3VvhlMDsYEipixiBZJKqsequ8hj5Td6eta6Y5xqwANp9RM
mG5HGc5u+wPBx37bRg2dRSa3Qz/JoaLhY3/s4nro6i5vLJtgkq/o4Mk5nveo38uo
FLJvWLVBMm/6CcQUyTKXqT6QAo7DYDFLqgtesyG7v8Km/NrdeoDBTqNXr3XCxPlx
9JnYWV6wG9EVmaU47CGjbzmdAOzBeCknoVUDsdzWOcsAefjCBB2drAk+cUJN9J/e
SE80eN31YKx83PSa/6McuQd/KWTzlzE3Swl3wSQ7G5Yki7zyws/X+dyQQqNtN7Wj
5AQxBmoEerRF+sf17qtN6IYE3rx3Fox5DNaTo3HyAF9yv2u5jGOxucfzWhCw4t6Q
jSPVO7WpfRWW/3fcuVjQAweMG7BIXGNtfvl2MP0tHcAZOiDa5kScISW2j4ctsW7f
0nFvEOavqpsSECOck0GArZYb7O82YhDGdvzNEznuBk/zFwCBOPMh9Ib/BLJKUnvv
CWaXO8zGeExJW7rK6hNkpRZYRwviszGw4jnNxmglq5f3jDJtAnW9fmZ8gzn6B/iZ
FOL0ErhQfm0Tb3Fe91aCbtLgiRlkVfzny8bShoSy4X9egzAZAUGB7cm/I0bAk0OA
qhTjllBVZJlYBFtE9t6UzS22pwprL5sJG0prhGoP4u3qkyA3F6rnSxqUN4ESu/pJ
E9R4bGE54QktVNHHXYCvfTYx9QkWW1ojL3PbgLUPgR8mkl+japBFfygrJo/lNc0Y
GVfVHc4PhnBYwJTVxIcTv92EWzMaM9Gi+hZakbHakzMarv1Ptn74BYIQe9WCtHc2
c7FisJvu/UP/OS3xUy7kNGBD6TDK+L82va/RcFT/Gn/6wgwMl0LLcDwaI3B0ifjG
XMWT/68PAVVfDuHhD8b6f3zrS/ZSIqw67BdiBTN0kpBZCOpgqvzH8z58lodMuksx
P8UU1taM64Jiw39PQwVIEFdfO1UOP//vAJ23DDRfXbRoldNhc8Gs/D598q2Ptrgt
NUETJtRtXE6de24IzZnWyHq8UvwGjfPBnbnPtI1HrpKHQVrmQL+wHFJwhB/TFkQY
ZEp72SCv9Zre5v38lEDWsESWLrdDzOL7r5eDZkH8ASw0B2i9pJgFI+MqCibxCSh3
ef8DgeWP9as3tH/8eb2aK8rgZ2KNIqqkccB1/lQI5pDOWO1SAVlB9mcp0u8dboG4
iavEKbz3GgVL2NDTVakdJLiLZyGhXE01NXko646x599KJ2ODuaUXSjYmrb1qNYco
/XkswqL1/4TkdlsN4mqczmKyOQDJZYoYI88Kd2wLcfdjJLvgD38oTdo/mR0qpa1A
v49Ia3feLrwkqULc2XMhyxsLvTXucD4uWuViP4ZYfEY3wFcwB8bfWMIEsJfzxdcF
p5WZseKRbmPhdW4nN02wwSTGVxqBkJLnoiE2l4/47BRzVruBUmoVpOMlH8LT3JXV
6hw/AlhzUJi6JGED0OH8vxnInowtWWndJdgVY2fIWTrLMPx13gKYIbsWAJICzsFk
NZL7GN3WTuk2q6vaEIag0vAsrzVIbmDCU3MnL7paipukUmPUMv7VzhM0Sw4VRZLY
iD7YsFbXt/fa53uLbat6JBkdPpVSlilVvZBcMF1Q3R/29UT6n9RqlVLpU6h6Fj2Y
H2YvbubszN1pvS7IOBi/EbaCSxKTgX/aSTtmwrh4tKnewjgmxWonrqoUKz6eFIT+
jmXhRtyqJA5uHYO1B9WRaSth2zShxpmkhfKzj8FP4zTmrJTVNgX0BDcaENNCW+Cd
5PYnzpfXA4wBxkpaj7l5bLIdCPNpiKWO+O9JNh+4uQHeka9W/4LLLVBV368RGQ2o
Zt+mAejAF12gxZ2MlVw3YtpAx6C7MbEMxqHD5KWci8Sona8KPzj6sdRG7Uv7gBdK
MsRyaOV/UElf2pzjcAhGzbMK25XqvHBJQ8WNpm/w5WAok/VIIH955OdoMlaBwU05
/cWAFDIzcQXIwnXt5n7HOSV7y5iybcROF2aMeh+X/Bjf/TdDdmWFJlfBAFCW5NOX
j8Hc+rAokDrLbwHK5HhouxikJirtgNzSO5jE7l5Abodslj4S0YOAhhHdWQ5u7WWI
Gdc5K3xNEPXI+korhefUUu/UdI4kkMs0VUkspOoJAXy1+26vKnj/Qkvo/aiPOxJ0
sbrq6MGl0guB5eH+874wmLAjG6isi+xDvkr9c/DXEQ5YhZbCpoC8BAMP7qq3Doeu
zzS7qVMBuf/jAyoeUAg37v1Rmt+/AmV7X3ohfftwOEMsINANgGGynU7hsFaXIOMQ
QyuupkF0rgNRpxed12eiI7krH+/HcyQ8p4RgG9GhVTH2s0l2w25ByDA38Kz1sEtw
UotLspRs3hwf+KEe2q5B3a1hz00Vd5vKvl/6dDSG9fBFkuZuHxrUcD3y0fpSPasf
E6PjcIWvmBbzuIUw4rU2aGDFmrlADAMIYCehQqjOPVzZx58a7dtGAceU8OhFvbk4
xQi1SNS/s/ceyB6lUzPd54SuBD72PKjxTtVWDUJYCZwBNjapmbzjF8lCr/W6btRG
zQpYKlBtLXO1kTkVXaHEQ5SapJK5Dp7aXN/oHYsA1VECy03wbYbJQNCAbfOsTW3X
bMa4vVwakWbnIUq/Oy9YQ4L8+F5AyJDUmXWPlaZ00qS4RiSdBjLwqvMHzuJsUMvZ
BoE9exqhaRO6rrUnzcvT5UfyiuJeK9AWkbqAZawMlwsMqcqeS7VZyXLNBIprhrYO
ukLemR4UMMWSYEVSV5+cvmNTZq1wsjj4deWxDhnA1/sMWzGbsPDpjwvDfBQ+2Kfj
lYzTMjSJbHqxKU+hG2cWph/YF3lyMBY4XXPFYHWtUlDGggW1ZA053B6qRBTrP92x
jaLeYeeJppasQdCxhrpz2T4MC4Ao8Ti+l6F51ixkKLJ531+YH4uFEVhMqRkhXKxb
NXOSY1yVpfZYlCf6xjJXpvK6Vnnd0lWUHUt9rhs3lM7MdYl582NnuGSV/9RLz12j
g7P8AChE1e/Hw3bd25uFOEtvVepM+LMJ4wehizHidTcnsg+3Dm74VamEBE4LOLa4
vVyBNzyz/ufuvaU8g/3gRaweRIU+WieQMixovUB321G6RRyJ+8v3VLMB976Jnpqb
HerHw7KTxlYS8CmhibnftUz70tkS467rwBZbMJrdljFM52O0T1v+YXcI4wTaaSO0
+djCYviVBr8Y8XJ9VqE5qzU7YMg+L5Xb++DVuCoJORigfRZaK9JkfXMCdYGLGK53
HoBDo+AlikGFNm43F8AfKlEU2bbsSJfNXu/1ar8ykZ1p4g8XFS62/r6jF0GKnqwW
7fh4Hrt7cJ+FZ3gwEwtcNq+GewzaaOQlfSd78z1UEMohMqkrxqRMUPwDhwJJVZzu
QZcYlT61RK7gw4Y/FgUIuusPaLZZBE/sabftREgmHS3qXGGgJvKVYESWZg3IOhVJ
4m4hPujtJw/nmlWV78yMH+t8bw/I9Q8tHBqQcu0PYGJ2jfnM/WbNcq1jKhpKXzmB
VLvhZKZQ65QJ9ANXSZw8lr1APfsMPG2yc8MIytjAqyWMWO7z3Sb2qB2wMXC1T9c6
sosb2KQh0PDNyD2UsHtodyQtQue2o0tMm+Wy7uCqGvNtBOLLsZBXK/e22jlsCYFk
J3vc5p7UzpsEHOfvr85FCeGPQTxpCKyOXTii0p9fwMdiNeIrsg7G9dOcyR3aXBDl
1L5o2Mnn6s6x9IJJTK1HAC1kTSgZF9AWHz09Lz1qtm7te+2BMLillBs5BSqAMD48
S9eMU2OqFv72DvV2Q0/j2B75MzdNCatfmmJnka13093cx0UTMhJNwRokSJSdIFna
sd9gb+XrxZfZR3NAV5N33nB8kvdGgS2aYPpkil26r3W7xTNSi5Us6GxV6WBT1IvC
sZaYnM13kBoC9NPXtLDaEt1Q+Lie+cnavXy8fcKSZ/yz7weLWOd+dKNXeSl65CRb
eIO3fH9+DTRMq5LyDBugUwiLBb+bYS88qHfwb7TagQBqWaUHrMCQlzesYLbld/5l
JLteFPkUk2zjctfq1dXdC4/bHIA5d+z2OeMvQrsqQTkLae+xl+QyII9vSeu3ax7N
P7t4+gQZ4qGvxbyZBbEGXh32SgK6Cb2/uFkT1fjw+TG8CRO/aFN51tJBi0k4mIMI
XIQ5eC4pt4q+qzRc3bnCGfd7dRPeFuOU37LwGofU3sU8pshLvUqZFFDVDdrOFkpL
b+dPpkOxRxrP1EdYo2B6zFhbFHj45mDmEomAj0/8X3j0F8pqTDPbIUHjrm4Q7vvE
E6QOfPT5JkyuVWWieB9dOj17Rc+ynWf6ZOoTIxgF3W0EuviAMPhZqOC0IEjT9N1e
FV2vGfbDFW19TFUaE2agJt2HHuBfmnzj8W16ARRKUY7r5xdqlra18NEzZYvxuTGD
lKQteeGVjicGh5FpHYuJCvuIkFZA6BEO/wIQ9mTjqkAOTH4El4Ivg53ClliOcNYh
vouWm393ufME01xOVuSIXvlxA/kWGprs7v7jFOodhddFfmS+Y2qqVIM8F/LiowOx
BUSc8gUlxAdXlY2G0BnMWs5a3STXeIASsMxyihViEXJvpXfjXwgYWW519MoO87KC
v5DqztU/opxt9yzW/aTnOdWZwNUpbkmMLH5PizXAGdrRaTPWh4g8lu6Yr9IiFHho
T08UvIUUExy7h1+ycKE9BYZ0Tg6tL8kwtRYak0ynFlhiGLDsbd1SpwaHlWcBMRQG
EGoqYMfrEAI1YTVJWtei1o8j4WcLnP+2wMHoFEicQficPOlKWq82yRQjQ44X5uja
4YnyBJ0Ajxgh2fh1l8iM8DzqNH6jbiHLolGD6FQ6e8lBETfo9hOssPZuE5xoGaUl
XQ0a+mOW7iKwBnCC5EqWtglKBHET7Gh7bK3p6xQxPHV7YmMoHZkp2IHu59jXQVvD
WFtksDIE4YFNe0A9iVvQisuY7VqJw+lSCp/gcbMatE8PXCcI0rbPmJ/5CMgq3L5s
858cWPVNMYK5r8Y+fJtzbqS65xdOZZ+fP7lV/rtAgUEhx6PByAvkm4bZ2FEPhXPE
K7ouhtQs7zUakZoQh70S1o4ZIxC/3fnUdT48QYvqQiFKRxXOAWsiArVaa5uIvk7f
1KW7JY28ltQUG/S1MVQ0+vTEYHH/KV2GjR0kqFCtSPUmY80wZ1dAfrV5ONzEjUHI
ld1KAF8uLwaJwDmshCMsthm1QvqUMo363tYy9yL98MhP0afO/SuoGt9/eNZVCJrP
06y5BXig7SxPVe0KQwSsqy6LC2Og6n4fkA2c7P/yPdhJPztisk4uilM32BhxBf1Z
vEg8TjJUdkWhYmhFLhMV7o2mLLTX4ZX747DgXFPuaUmJInp0vCUqjujbLPoc6mDY
5LP5jeJp7tt4e+0+KD6rptCw+pUHb5Eg3fJ4Qxz4y7Z1CUmfTC44c9DpgJfhVYxF
pN9SEvbgFV1svkDvF/R7BgpcGU0gBI/+R+2cQokztZTYvN582FYC+fZOkHGF9dA2
bxZUXgQBHdWD7R+J1miaY7sFGkjDA8nUMMPwXZ4fbHSEs4DvO6L8+N05jzc+O14t
sc+uDQapp2M4MjajQeqJlD0vwoB//zJsucOU+B35b4ILSs11pNSIdEW7ypZlTUM2
ixyLLh42yy8kq1sLAAYC7FA1oYdZw4Rz9uuzSd0iFXjHosQTjxxU2hmYcAZZgYg7
KrPIh4bUTWaIkNqvbKIjevr4sZc+vzgB0OA9XmUuhQ7CwOvMe5IKnhe4Fm3Dyg7k
g4d4vDpMVcPACH8kAm3S9E5znV9YFXpwEjtXEwred9mEgncAoMcTWOquG9khzocq
vPGi59/B64uxbcvAFsAFEwY4hgvj+e4pKJR+NFaF+ZwexSB3O8Yjxi8ccDVpmg95
ApfZY7cqzCEgHF2tRYt5/YHExMFnQJC0mLWim495pOcgekjtSMx+PLzsihZyWaDm
khkugTpWzo/bYNxpuAb5f6ZWEXAZ5I+calaMBVA1CKHGNRtgQGwbNuBKpPHex4hd
5DbHZj42GNUWsk/1fBajRuRJameR7s6tH/mMpmKptouURNEB/ltysSwbj7/TNcG4
0blQEUDq5YYBVkfu7CZt4zog2s9XdOwCic3EOWuLEMSRtgDXXVUgQWoRbKj7zzS9
KomPFh2VSM8IA/HejxSSWAJ8wGHIsxpavgV9tkLUJYhEgNwXzOWmbk5o6IZHcTpn
v7+iQKGWOFRrzMDB61AAAZlCDJwnSrvuChChdzPOB1MF/3e4meBYhQzwzCw6FiFH
abbfedaPAcus8UfcvoWwO9Wr+aZs5sOuXrYNv3FOMzcV8wDwwug1mKOJcnYrXavt
7N178qRRVHxtjR90vayo/Pp1PUPfROoqeB/LF2+r5WWMv3RARqgIF1/COh80yBi7
P6hIfYjNcLC3BcuMK3yQ+vgG7as05vBfUwvkX5SkfzCOq+zYqoUNmPO/fiN2x0S1
yJG5qblFkaXcueOsTeRFQR6AYvLzhd5zV00dC+P3Y58isztT/rJ4DjZX57HPcMoN
KtZhE0bopmuB8imgEiGjWvAp/HYhvpAXcskgmbLpXe03CToL1eM7ujS70oZYgEeX
OXJWS0nii5wNRurrQ5P2iSy3/CXdW7EeL5DKhEBSFld2Eu94btdbBTgwBJIy5f9j
qBm1r+xR95r2zr7+DsNkxta0bJq9lUgdAM5a8D67zI0t1qVWy87Z3ImSL5xS+55Q
+F9HyrPpnQmsIAN7CUQnC+F8orRi7zbnbPzaAKU73Df9lKRlAT3Jxojyom56QBH9
luKJmUbgQncPNS3z0C9chTfw73PgCuSxdXt6K8dwvQqEijqV6YSt/vG+up0cmISU
bnIZfa4Mshu9wB7s9bzfO3kOHITQfVcJqBurvSGsjwVDKY3rEO4gcpea84p5J8Ao
Yj4rwE8xDAPET6lIDhnHu5Sfwd3qH71aaFfX0DQBsALXeeYOZYLot7xCvLOsng+J
xkr+npz/Uqadm8XhW0aRerUFtEA65ykeXCSEZkBlL5FCVqiuPJ/LjnAF2TLWXQZv
npfi9ELbASCyRSeh+8KY+KjgOrE5gxcsQ+lmCuykdnPv0iOfhAKGWL/GXh7eqmA2
gvvI6CKlv9U2gDIzrrWle8jzgITn8pmBAhJz/dBz6elFIHXTWzbEX1D0aN8EmUq9
Gtskq5AKRUqC3CU+pxKmb3n9+vFvO7pfdZGe4YLyNQ8/5LSHKEZPti4u2Zw2m1K/
553PZski+t8sI4xzn1hF04gIfD5uRc2LsW904hHJ9UNVE0TUzQBWioeHRG2mXqG4
YNoduhdhK8BDZhQAOSz/HfemAv4/TmGnB+7LqqsKl52x8Jetq7f08il7WNe3bseK
Bl7jTnN1WsCcrw+v8mCwI7YYz2YkxAOlx6PtLLbblcoUPBXbo2gWN3TnzCd/2wNj
XqCZEkcWUNZtn2EiDZDKQgqQxNDjQHY1DnNv+uvqYU87FrRovWYcoBIpWQXqyNDx
YyyQzVAgBFk6r0UoKYLeyXtMdD7uVEaT9un6Q2E5YD4plfx395caZRT/2mjDnsbs
9iePy1OBjdWU77HHIapLgv7QCt5n0nXJSo9fnp5MnZue5x6x90ueeLo2sbWNTedu
t/vjqWHiKomW1HruFv1TSysjaeQKeWXcxyiNgpompN0dE0TSP3peLdNIxxsTqJu3
pzD25iR3klxWwi/8ts4ijvwXfUtdpGJO/frmM8hXx5ML1bY+QdXKZVTFZfGVY6CC
Jz9ZxZ7AylMcAgKr8X/KOZhZmtKcx0vUZtAg7sQqQNA58rtvmBGA5AbX7lwn/5yt
ZLZ5yvKzW0Ec6zDbjPUBIRbxJTyCXG+J6DL9Z8s9wxDyNzqc0mg7Ld1eVALFSr0u
l1kJcomXHoOwA7eOAH5JdMvFyERNtHsJMO5jBgqed20vXcJ1Uc8ZxzkGlIJzltUx
pTcSUpXB1fl0gfo38oO1743JwkLIPJL3Q6dBZly0rmdSZN09BiHj8/UOtja9tcCX
NzqwPUO92h4bwBUwdIfqx7SPmQV8lEPE3ACFPO5jT+jPdzRPtHVkdlfndYmvrZFq
qJSQlkXUhfKnqBV8CXqQ9U0d+4/QqCEof1xZOvDdyD28BFP08SIgs5XM+zY/OpeY
YhyT26qjl8WUdnz2/KGFmBAOcK3J9nAOpgr5hXXFq7/1dkf1wELVv5hR8TVl4hwI
q/4yyKpCkIxJ9PaPZQwhyjxYgXsBM2qR1cq6tC/4qHr90JDEgWmMPTea0ImgKL9r
JRqN2f5VDaC5XLJfr5vsn40KGMadsEkNjG1Lx9PKW5oKvmH9B7zOA/wgIESNHidk
KgKRO2jU6fR3+4htGrrCjycc+y8ErO4Bqh5xzy94lRy0w+K7fuzuJBhdAezZGm7O
eUwT1SiYITbelEO0c/k4PwtchK7ypMxRT12GVrln2ol40XiHgqpj62EQs5y77A90
xyNLeAsBXKpCjcVMFzDUhJj7O9TDxpHlyYU3BRZxDMn9H/p36rZWSg08kdowaxbz
LcJEmsRWCiBQ80svmA/4dksk06ynp7V+3dLudmtLnyLXqfdfMoWUKptwsYKV2Fc2
hEFFQ+3fF3gdvN+4P+5H9W0dEkLlLvLgHPa3x99r/XZs4TV9P4wdju1zbgNGvzSN
xii6ZGlAvJFmpu/wnwcRk8wCgR9vLFCKu/siyusQEIBQPh+ioJ5PS5WLbM45OsJD
dQ886o7cLfypgmbkSos6VU4vQnLiz5N6VlGam9TM4Fh691e7YGS507FIh//bcQHL
3PHFIytGfXSdVs+LS6yUlqniKn2FMvwTzcmpqf8iFwGrrTxKIt12xkO+iBYd3SXv
euXQ1Bp9AbjW6jkBEeM7VsC7YOYM1mYiVkQ9Cjdq5ZnH6Q33Eba7N/ByWAzYkMcP
o3OC1TqKnVMwtvM5dTwVPgqeaxitH+FpsPfGvpF8BXU45F2AANSqhOxp4o9BXnwr
iw8u/yhktBxNMN7Hztn3YwsAqycO1GctD5QCUPudQjNb+L4enV0NoBh9zj/OnpbV
PggYMovta6jdb3FI1RC+JcQSOHpPkPK5c1vbipmRy3vfFaBJw159W0lDFEZ3pj7G
jb/D9Z3d91RACsU90Wc2QoxhPcsvkv4rwo48FGnFlLT0oEadhnDL0Nb/gwrZunUv
f+aChlKS+2MmJqOR5dPJsNgG6lZWJ95Hegi8915YAkAbk7M8va5EY5Qv9zYWwsOz
WXa6NXMN/0espJsLJ+cDhE26bhMQXSqGt0hLPRex0XKFmWUE7Aknm1hH2T+Jzu06
K7oOO6Su6u9/O7R5AOrd9lRFuOhvPGSpgGTB/WsaqH1j0MWvw5XjjOx0gGN6Kzs2
MeW3EoQCVRFMBPNcfOrmZ8JLfRUEMc50fSri4FD3TIvEKDgBTijjQIBdR2+PPhkR
LuVHGHPlLaEpJUyW3RqKKcaE28IpLGZlJZ/kO0WGdSsuZXu0MucvtITUYheWTUAo
wZ3jC0FPE5htjIN38zsxegBj9TATrN0KQiY2T16IfSA3RllSYN26Vvsxybi+DVVG
jsXN3Cjy/PefMj2TQdVygZpmTAPG+JLdYLvEF1DW81rgnZE1dZx0eKSTtnh1EOBy
N0e4FGpIbA0Z79IYHDbJbPry0RadxLzZJN7YCt4TsvJn+/Hh8l5n6PgeA3f8Saer
mR9A7fVo62e2IVvg3ZnYv6v2mF8qGWH7kZz+nOQC1Ah1EwrzdoossgGc2T3WK2WA
y0Viu/ASwSFpf785HhQsOsYmtpT5Zw2nroXN0etJqvtltscPjC+U12hjV3qGAo1k
MHcaJG58Yeq1dB1jiqIZ5/vQAXO9plfMVf7QK0g1yHESqxVEZ9UA70Ugba+M4Wih
5KTuzyvBmejpvfGGe72j6j9oyRuujv5cf7+OPJenQlCn+tio2EL9IelWcV+0w7cE
A1NTHEaSl8qEdmwmX24UiQQKrh/q++Thoqxg6zP/Adtlr6Ywq/2+scQARflwNsRX
KdnZTRs6x+6fg+QAQ8SaTSA58FSLLWGYNnYDZTo2R39SliBvfiM879AJQFTW25kt
ZhaItZwRrtE9Zelx/ietb0PAmxoU5/2iP4q3SKvD48oWRGsEYwEqPCQKE/cA6Umh
Th5d16/iyiETkl6eoR41m8qwYYdcRa7/FDTnso+Ze4kNTWnlZkRd+5jmb9OQuQtI
koB1ZC0kJT8BB4Sum27/L5znX+nG9XuHourWCBNHHC9XVRRy1bWQnzklmA1Jnk9F
Y5WT3iwMo6A8ojApOxkFQOzSfLX6nDKAOm1VsyLbDJVNqcgYnUgAjvCrhjUF/CP+
2Yjkbg5718rswp07OEBDLGUsc9cu728JA9PxtaZmTF7s6P9Zm3n0Jc3oVsvJGNI1
8q0QrkbqpB28vz+znk3/Im+50Ghyl1XoN5+4eOIV3ZrCuWcwsCer9pA258Uvw7RM
WLx17ppjYm3RMgYD8v7JHdmhYAONq8iaMiUmWyMqqUjAD7l+ZmlMQw3kN5V3Igfm
+pxH7AQUwLUJvPbhRop8sz/wQdHsYYU9c13UQiR/wVfF6i4GIq/g5E1gl6zERzWL
FH+rzkHiAxOjye06UjoNXlQMwVpRyMlXDneBl8mdVfnGWLpSwi5BUgkmdiK3fNJf
AuYjsLjGfJrcK/TMNUIhZ/DKJckjeBzE0y3OjITj29Wiw+K4cImxg0dtGgIsa7+d
q3MbzpJ7OhmaQalTSoW+aPyRwVGbDE1GeM5JF0B31rATAClZExe0OwJf4WvSb4MC
WIDa+p6B/FlFopFUD6P9w7ZwR785dCa++FDPfafFkd5PZXkK05xuv6mndjE/nROx
kIZNY0bCa9HiMnAXg5E/Q7GUZVYxmX67LrGx78buVQV3Ne+hprISjrhQ4YAvGFNp
qSGdErL4tw4EPOsk25ZL+APIrJcO6Dl84OeXDZXRGqHEBPieeZ+WFrYc1BvRs6N8
OZl+ZSYweOOGEUY//f1+0c4aNZJgvgxISrfFLvcA2PD3QBkBoOPLWz6p6Hk1+eCa
cGiUynSOnrJCXXhq3sCKqcopL/0IC0VHAtW0RF1SY1jOjrFCLZf6H7lAsQf2VYSG
UYB1DXmYzqzuPaOwDC8fbeLPPN0m1hu2hWQjQCAVdXu5feQKqSAOZhx1/+IOyxN0
Q9PTNGyhhOXmX2O+Ww+deEZm1RxOpEggWi45ubH2MMX4pecx9ubWjWnlUHADABKS
mbt1XCkaWF7U6Zl6HNDjHJ/hCBsOMyLfydnFFifYBFIcnYplu6w/2fBNf9NggKY+
UU7JD8w0IKTb9DTEc9KLdq1toOkO/SDZ4fZ5KaXD/NSRMpbwv6rrq0jCXWJAH727
zoKnXo387olo2HylfTPVAFOlkmLXQ2TvconNT4wOkrq5tqxaClHulN3IgVMCaNQG
CVWt7tErWjYdstMwepQoKEyC3EZGU8n+1s7qYUnVTwCXKQumkvT6864C1Bo67DFo
yfif546vuFsRBX/3Vy9iAqz2EiuzSoRcQyQdk3Lo+oa3gQ3NPtIQ/4CXabjcPw83
AOOGN47nKLdi358eRi0tDsnqp+e4G26RPq9iyyLyZZ7liMqWRF8LRUSzMkBiqVmV
1qWbzmDmcJtrWLO5NA/CKxz3gC72E/pV2c5xlRSIVqd53uko3XX/heWtFOtfCOwa
ouxdlSbJYc+cwfg0SNKYwauBFTAhS7whHgiuyJfaTlZa0pr7m44Uw1P/xCzPN6Ra
pQrEV7ayG/U2uASoAFQGDT+7UrR/pd2wILz/Kb++dr6JfaLdGRCKNS+Xp5RC7i6B
TJyi46SJzeV7l8/iRksQueSqXODKs2QF/WbLR3OOU9KxENvVe+6CUh3BbnHvKqoR
qMJzw68pu65kqvhANsqwUnA5b1PIFpdoyAkXij6/Nhj76ymVCgee678HiMNmoast
3Nos0A0APM2wombCOUKkPsG3JKJYZ3M+WUNCRuOjkmzo588Bp7mLoMDT3AWsygCW
4wN5DfWeC3g+sLsoCOiMnyy5eSHN6TtocD5/k4p/6ijTjPXtK+QYPtWdxdIyU5iM
xcJXiJ5f6Uk3N0ighxZIwWng2TSaVvTDQArbdfXPXteYu2aHAyXT4Bn3uf8kqoaj
eE2WmpRxCrksXFo4BRlIyaNHHcgnJ/yV4XwcdYb2plIezN7od4UVGPLri41x+CSL
tSC/TokR0M1bh6ApnrqiExuCHE80Y3cQiDnX9PyJoyEfkQ9+XwuTu4J/p29sNAF8
air2BYRDrn+lh8kz2diegdt4T4cIZG0vZmVVfMJ1HGuSCVRe40NAGO1LAJZF3n/5
XT7USYucZ3w4yiNg+k1IZyFE3m7uih+Ct3KjedaSfMdF3CZl0en+TrooJW9UyjJl
GvT2WiL03JTcTrRINawvUgeuTO0n/fyv8rlTDK6e/Kytp2yno0wLBnap7vjcD/kN
ymsEgPYVQGfW2+uQx2wh0Y3rA4LI4UKxtquoZDXaUMVByAepS0+AJwId+J2SLoSz
WQ7BQg5WWHz6+vViPOYLZqfJd47qO7Bhw+4bfdVA+0v2M4/Nz4eU7hH6/LuW390o
qoHUHAhVHweffGLqzTnYz7zzXj0TJEgw0QDzKUefICwhrsTunlzrAetaGfKWYCh3
YdQzPWulnor3Y/jZFNQs0GFciAwXJalVWPCHL4pOoDLAJCHICoEFZfVmNKk7uAZj
C8OeOMX0PZbQypDE0ZdMeO3N/VEj7yXGW9uMnW3swjiQneOttdvIYBEVKlDagAH2
SZ17JqGUAvu/vC7hkODrNVs+5uhbIjBhY0QIMXHZsixPGRGV97KGPrvRocDz5Ptn
7ROEyfdoyUkZPI1MQYf0ovYwfMtMrjitrBJFHPNCzamLz+A8NpG/bxDe/39y1l+G
e8p8EuhgJazo0QMUC7NFoZ8mBlBtvm2iJ/xzQfualLvWs/mfCmUo/IRQ0Cv8gyeu
TkmTpY0lhqi2TDcNXilLI+/06craHuML+2uPjgd4uGZeEyaCGZ3AbS4VouyO/vuj
9fVPdn9u6Q73QWRZWsQbf2d9ufHhb8mIavSILZodEmAqe+GvMv8Pho8GJd3t+obE
C/yJ7Q2yRJ4/Pa0CIVQsjuPaHwnL55ojRLVt288n1qhDcS4un6+5lZ8604TduXc+
qjN2ltotkSO0Jn2TtPk191yLhUIBh6X1dNLSKoEZKsiwm+bIiMk8QQp86aK6vYoZ
RTtucPj3aRpyT3DKM6jfVv4DB+cicsW1JxA+NOxrJL2jWvKuz7CET64TDWsT5er7
OxRDMhw62ElNmHdkieYAta0DU+ie7+tURqv868P1TrwXhUJ5jQIlvbhkSWSpaGqn
Zs+GS+83AZsg2c8+BII1TS680mlk9LzuLytXJzWzpvSlLM84zwbMuAdDFHTq1VR4
XKmXpBw3BJ/voQCtyjQJXF//Wjdl8YUrNqen/JETzyJBcMCc5duPDMkNUjlR5DkW
Ln/BIr44RDi5ofmmD/5vBjfZKgdSOH2++ugaJjCmGg4QJ/OYqVEZtQP128GRsPJM
3SMpjxGTECPPaFLE0B4iPK5bSxMxaRr1sD0dhO8chKw7QUYKM3sKG1QTSqb0UPMG
59Z7AFJ0V4+oNV3xVcUyrcoQ3a3yKlIuyuKxpBfGEox/VlNOBzPqz9GPBQXl+5tf
l6HPrQtL4LQ5y4wXMjcVeQEK62smnafr6qWzh4qV4yZvZ02zVyYmeS0oKmbFJl7L
l6KcQMnalIfq5JvfBpVrqPozDvJ7FSJofNdoL6ojhjuIdcOOj8LFroRNJQmQe9OI
fbNf7WjYCsftPN+zHOU/4qO7ggsQ5p4/D1I9zvpRLA7vvztmaGrq4QUM55Ee7jCC
fuhxgPCrWXmjGJHY7oEr9HhGHIICb1cle0N3X6eUeIPB2fY9lbj+L1WFBmPhBqHt
n2iTLEocQt3dNM0jp3JyBisuLhcf/T52usSGebv5u5d4fAiQCyAlitMIDXwSddBH
kSoJzWUUOAGME75OTPtclE3YvW71WhDzt10c5M9hvNiim0A3kjRO375odaYpYge7
RbdcX0kOd4Kuf08IL+2irrMAJfb6ITcZ96+MGUzZiohTcHPmFilZOeguqP+11aRo
zTobFdH/5FbuFFDebH34oqmp/QecxqnAH3RoteJDN2t/IVenySY9hR++NwWn8qCj
GEi6zLkdzWPZVu/1fYJaNiD19M7f8+B1R0cYfm2yuxZ4uasEp1bv/scEEb8+SIPE
cocmxvNlj2EOFyZ9Q3H+SLP1GA8/+Ipp6QB9lWs3UhzKhBgHWQ/3f/p4CBzFn76T
+03L5Sg2ZCJ9qh0TisfDJSaxmdcs0XrD1iX/gNjuOg7v5VblblkrOFfYkri5mK37
ts8235CmEeveoyzButjT/zdMbVusNsNNEyzcvoY2xL5acIuNDG3Xl8nRCarVYe2D
uXH0rGARMiJzRlh586qCKAK9A7wPuhBj2TO1kI5OFN/lngbWmCf7E5PeQn0L3jVs
J3iGlwxO2xxFsptgTx92JzZ4R8e5dcUo7G+suQU4DXzG4NlxyKuJB0Zx+3VAvWLi
n6w+JcJHnsgjrJQJ566NdkqmU7Cczl8lamv5D28dBR2yk1Sn2uoyf5TiBAggXPd+
dyfH0jf6nFDwyt1O28NX24xZumWQFVsGBLxmKC3N5/2OB435OKFAty6/TsmOzD9k
ihCPvqA4fGNSo3mAzoV2ybCSFZjVicDcPOflNii8dnL9liBTWhNjREoR4Pxv5sEl
fQJ00+yneEzChHEWWhxpxcXI8s25D2jNSyr5NPS/3U5mVj/K4ne39SKux9l91Xwm
AMSXljHK9Rw0ONSklrEbK/LiUUwNT+Xhqt80bRs4pkZvMpgEaMM6MoOpumBUMNKr
O0B1yJ1SKz5GtEDOFuYrqWR191IvOXNCN5fFlVT7hLHfe1v4vUhHgEgqD2OKX2MI
i7ikNOPANaFZnKZ6wTiMYyhAgUa1kX2d0n8NqlOCDDg/OY1GeyJ7TvQ6wKKkZclI
F1l1ObJ07SKfRP4yhXucIJvuztsy3H99BQZUqtOKIUyRCOrTDO9glxl91q90qAkG
mAfuJzhUNWEgTS6VeLqQY6yL/E/fjKzfrgp5jyK72c4pBLthOGYzFmZH3Ff8B4qg
eYm0QQf+9sznWB8j4/VXlMUy8rsdb/DQGPgdWANrHGAMNAzmqWfXnOoz/Bfsduzx
HusuGBR+Zzf7wvB03jvJaiRrlgxvAn3CzCeNopUltKsyNn52toZbdGSp0tpzJlrQ
hKpGAGlBWA1sCiP2X7xkU0WJcy2fTDIavQpq64ZmaI6Q+HX0nroaQBiiAVy2dd0x
nNiiuyP6rdc1z4kyWrIjF3J2lfto2wiEpzG80ttrBl6X0sv60ZhCtd5IhkyWf6GN
zWGAcAGyiN47WxeH6t+0O2x+x6NYOISzuD85ZDmu36Kb6VlKEK4PRZN0h86Wl0kl
x6st3Ij1mZ8J+0Middjr/KHPh3MGg72YIfUaE+Hf9AZQCnoVjit+f+z3HokwXrVk
kyCXErhWjq7J2OdxHnFUnbENlbKsKU/iXjRPOnA4o/C1oihnIqNTWNOk6ARJOlW6
Hdv7Dp/XxmGXpj0fowRIpj3r+ZCADiAlb5qX08J+CvHj3K4ex521KB0ozoBnILbE
JH7Syuc1VxySl3zmBuhuMdyc88WfSjbbR97PgCsfiFq6y9i0iO7iSU6huzSc6L2g
AWn/L6Pepnfk8riX/xP7QWsD5IevXmIu967Jrn4XwC5N0rt3uTKYaHRTDzaI0KFQ
yqfhmh/xx761TkeZIBK1GhmptA7pgR9VQBVUOJBaH/TA6RXcpj/BNY6MdLUvpyiB
gvN7eO6gvn1P3yYza4i6TBn8uxWMKHcQ/9IzTigtzwezMOP3UkbX4PMqwvsie5Pi
nOXc5eXuzV8oazI6/3d7NI5Nf7IJh1ycYR0snftZmE8VHo1ewGlCZiYLiVQGq7WJ
RIs0lsoULIhzLwJUBqi6QHB9hVKQ/L8Zx9zMGyN2QwFXZzeRoAC4ec5MTLvBmVFR
iorwKi3Dc6yljuxSre3pT1I8Sh2sLiq8pFNUeA0nHlV0z5ZSaB7So/ho0ginpED1
B4AXlO9BuldrX1t4AwWKAz7gzIdtNJcOEEjzgJ79Ur/BkCGqJ9p0ez3RH6nH7b0q
drrlOq18vNNH5gS/oovd/3ZpO7H1txxv2sccF7g/Ef4f1lIWHMS1ABN5DSgqtb45
uUyfm0ctWYawqAnQT6JQGOTmtu7llLneesZUzN8Sj5RHP0LoH6dJLtqCFOrmtKBu
94h4BOjPI7mSSh/7YsIoMS/AdsqvJWAz2wi6tlPXYmMgl7LBGtHMiKRvQjPBSV8N
Cd8EVmz+dTZjztvYYljS5drvcRAd/UwPRcEBZm9c+0RCxerXQblauPmZxJ7tk7SX
EHyHSRII/X9ze7ee6H4iJum7ZDXX3mOw/dGiQsdLB+YFhtNPzkbgVv2CMp4rXBxn
V30g/cDJiSLF+VY5rsntUsRq9uSjkCOBKPdEJQrXystGgHOFP3PyEVIoQDUI5qNQ
E33QZHNQeH1b3qbuUdI4lFtbjxcBXhGl7lLd0toE4LzEj9AGc6p3Yz+hR/G0sN3H
o8FCbakwPbNo3nid+/PrssVQzfhbjHrZ4canwEFwQtGWQAkCr+T6bGAPyPjszrf+
Fc3tgobz6nU5IHj66oAnXC4kugDdSSnaWkPSS4FFUC2BZWz2G7RCehbNDAw0S1I5
L0jNRLgkH2WmilAjKZ9KEG3Ku8aukr6RApn5SBrExQ6KDSUcamd1dU5khnm4tNd/
1KHfTW5/idp/8WOsoZl2ivwZzN/tvMeXqwOk8EbWspJmO09FenDYFCsiYfLEmwK0
qitLocg5w7D1YBBL6M2HeFvyNMyo+VEN1WakIZamcvf2roAB+saQm1JBUwHRw3bd
9s5IR3ESQh9/rctrgTA16T3mB1zScjyflw3u71JiX69txFhsXt2QSp2eLhpeFG2T
HkjKfAXot4fVGdPF6P43eCe5aaeaymBkAwWOv+/iHFjO3amDCHTxp0eDHzoT6vFt
FWCHcSnMnrKjJJ5a0tmqQbvvVhsNTGLjgz+XyiuuJAYvnEVle2GhXXTp5mgIY/9f
nT+Y5UhsLV9umJb5nbKtqgtK0qMkRK6tDks7MEnB4kJviHBgFF+AxtGRoIr4AQJY
NaHBAGTw9BBObjb5dr2u7yhYGZybQ+irqkZ5DvN6yHuX3nVE/ES6Y/ITzZOHusBv
/Q2Q4IGp7OJ7apSUHz1h/3s2o4HYajsNjk6oKCvy/o0YarBkbU9mIuLDzwIBO6OS
Ig3HVqzkqL6Q7hs5f58sWoI2DE9t2JWeIA2dY5DbhC7mMPsmMawIptHK4gQ1lXQs
EG4U0fmV6xjTjilXAI+B9evh7dC6GPSv3oeWVNR9Lr82+XorclpXJ9FZSGci1mjB
3ZkzPbP7UWcJlRLgNWIt+owdsbieE2HWi0q0xzutzL/zcGPhVBLHzOLCYOI98vKv
tsw6dF+x1UcSQ+DQNJecJHn6wzPJgqWIvrbBVyODCI4Ee8jgVdobcyqs7Wm7Wfot
DlCH4GiGyU+p4nVka1znn45EOXvfe2HTDcQtHLqP+F4Qicj01oeoGvB+6olvg7j+
9MV9v3Mv7rinXDOc/eEInMsfoEdxkMZQGzXls+CHggmUrkczCQNa1isYnquQm/LY
qjmTRB9XkQAlKsXXH2x/Z+QK4YSOpgwcBz4ZJZhT7ACoKIMvrORKBUZhsBm2EI5H
ohNDfIxOJvTp4lu1B6u+R7xv1bJOztzajAts1TQqKV/1r089g8pPPpBBOjj9c9ZR
IRgu/pJciax/0NIKFHTFVhMO9LR9Hvl+3TgjPAonxUJvKb+8fbw/fBciGR6v2Fa9
N2EYBnQNwuRH4Hi3r87sHWHyMKS0+qonuJiLAk6oUza1fFso6WEYlINlfAWyWS8W
IclsNKpsym0xp7pTOCy+Cr8LZ9Y+PGSONPjdjjNd9uskQi/omz86UpCDTnz199yz
p7ENoDhZd8WebX6TNFP3jAu6lDnRNFe443FIsuxAqaaU/WtnaKliqzazBMDuPD2w
ghUSrZAthhKovl3KZPPn2KaehF03QRbAjhx0Di3P6A/jQUH2rHTw0HqEpPaWqnlP
usq5hBAbGX5xHjHvJf9oyy85bFxLuwNfPLO5GVnG68oxHWKBdX3QhkjZtKmSlM5I
jYjeVZLOuIq/CVa2NVlbT7c/V439BkEBUIgOwEuWmJtM7hk9IdnZEoS4jhTItIPZ
KylHhBTc4L0EslFEpJdSgezchwAL2zWpUGSiRUZCBqQxkZStPbEiqc/Ldy0viwXl
rF9mqHLQs+OZm+Eu746/YY89k4zhqv0ytiZT5CQG1e4nWtt1C5AiobuU+b/MDzfD
hKbpdwXC5P3EV6EjyiALl6dW08IImHR8ViXp1uJMMZkslgjjzRCPE6RSuLtu+Rag
2nvW6Tc/qDpeGiEZua3IYw28QML2T2aDG3roIlLxdR/QsuB0FNBIl94chRN8vw+A
MaogIQ9txSTWzFgtcYUUXkwWTr43ysT6BasvCLAejtOqQDsxnYlQA2x3LM1JxqTg
v0ELp9wdQjsmzUnu313HU8MjptFbF9BrX9jo369krvBJAqpCtzR8hV9GlHJIkS/s
PvoSI62/2xaCR3Y9okWH050GYTeyPuSlkMkhMul0OjOZP19bm78JJ18PDyyynZJa
4alQTqsY2Vj54ZermsHkfzzp8KueDZBnM/IUW0JUp4O9ZsJV5A2754UMtlkHzxQu
EL0LJ3lSiouTumOg/dpp11n/vVm0xd63m36uiyDvn4oKynk+D7zxMmRkEJLOALXp
l9jrtTQD6WmKxdfvyZnQyrM5eC22BZM8yCF0LbxMytHphd/U5E89QcNi4tQFneYV
1OS54iyCU6DNvz/llS4uTuyxgld4QzvYVCYh+KDTMdB4VZuD8c0Z79+mndm771EH
RUZt0y8WjxSNrjeMwBk0U3AeMoAIjcpMNRzF7Fj0OmXdzkvLPUKdb8WTIaQiEfSa
tHmbKAj9Ro3u0cDrUlMV99oECoYHornZt3b2EwClLleLzbApdVSRg/e86oXWqwgE
jguTtTZORpGlkBUoJ1ehYGzRt78jL8u4GJ3BHLpHbhYkEWU+O0NwbKQw7xo24w91
szDWLwVMYIN0hyfH8wmMAMCPa+0ekN6D8P4OqDJX2pwSagT2tER4G2Z5X2k59ySV
9caTehysYLLk4A29Ltbg4c7rIbOixQgzXC0dydOtVkiQibNd7hIyBoPMAgKqrW0w
U3XYmzf0i3ouvaRtSX5UFWB8YqYsYfXxBsoUaw4cGVx3R9XbiLiV+OnfroxM3JAI
tWg7I4IAlCYw7jNqeMnsjNgvZ9mkCqdPIRV6zhc+Xxq17A7wlt4z4qqAmRe8Of/b
QdxS22rmLsR/wNA/DtmHahDw4vNG6wHVC7+Prw4h7GJNZa1JN7L+mq0A7Gf+1XKT
trbIny7An934I0Fsf0pZuYkTx/8Odky/XUIYSPnv8GLxjSp43/R8dzIKQnezM0vb
aq2V2uuUgzPtQoqOk5RKqaM+gXgWCPqesMhLHKiskXFwjT8Xhmp66GihIK+WBMu0
sSGjR8kEktIkPbqD6ZP8QbaauF5y+lXrYCzk4g2/Vbg28zbRVvfeCZKAVBv6aCNN
i/CcNrjqUrGcxValvarmdu+J2Qgxss1Zj09XAPvQfkLTeRuhJb6UZEwdPDML2Yg+
WQ+4SfDB6Z0zdVhtZmWk0d03ykV5Mqy0qCg8q5kUOstPKo3sxKCJD/6Pd2G3oLJ/
k0GReESfEtXOIb23hf+XiYyS5J/j6JpcVRZBaYRPGaG23xZFnw8R61RU8YLEUWpY
AzGgdnXBf37hC6E9s3uHg/ZdH4lE5njG1DyUA+a7E1YtdwjlEiq/ObgCv8aapxmJ
c5cr2ItaEz/ABoDxqeKXHIXP3gi6DWGGOKOxFJL3vaw2xfZdPKa8WnlUs9vQHHYj
EmzOq6LwAqLbw49fn86A/IzOK6oiExrp3bVoNlTnFI7PM1Q6atCBRsBYNCaBl3JU
ldCcsht/6stmdf8uZSIyyKyaoUrI8IGKC+2fRw6qz0xWf64+J+FZi7Wiw/5yrcYk
TbX5la0+AGqx7HSjFgUr4FBnpkqwu0MsW2Y7CuetRxipw4tVgY/ge6Zbjs3OWWUp
1HqXl5VjLs9xJGdPsHSjUjZUPoJ1vpJON7UapuhL9cIWGAtSNBKrS7TCrLfHw6MZ
SlDqXm/bRQ/RgfL8GXQW7s0s051ADIohngkeJuRm/FNdhRkkYyHUGIhT2sY0fx2r
G8eeEoEb+pBt4/txXlwldhOX9OcCgAvKyfIVMToR2aBZUdOF6ICTfPayYT4Ox9KZ
3T8GMkywRzxIYnq7/eIWTHfgL4mZuS6RYUomMg87UHL5pSpsGY+aDtWCkE1zwKNC
f01gYte9wlSi1IOXqXsOGZRKGmm8zHjvRsKHksT0RdTPLO31yMPyCPe5LY1cDbKT
R+tunjA1FEWAsAbOik3LZ+vze7RaD8zSjURnqAf/bkKF8SUIS+dDwAmqAB56Dj1R
0qba5Kj4spF7Mj0Ga6DcBWhVGQMTigOoKfEG/1CqARO1sMUj4/tz3O4exO6aRrxs
TL4lEvX4zr1hudCsyzQ/r3yCBjX4JOs5OulxsFryQn3bdQCm3Yj4IyXCSQusoXeq
enYSRsTx/WcKv9Cr1Ri8u6fTFflzi4UBrWs7wwn8QYwX4u2pjV8e9wQR46H2Rcp0
posASfIfaUFdvL+0V+pUSaPGBcEDEw7/HgqPX4W6qkeMnPTQ4U6ZthxWPMMxXGV4
a+PopVbq92ZOoGkr+uchgNC8dlmeTjl46NaXYBYRymrVfZ5o6TmZxiuP3F7kAc52
Vdr1g51xtyriOY0I9V5wFjyw3TcqFGDbzTP8hG1VSDOBXqqGFcmuW9MAUUlY1cwK
+0gGr3ZHCqkpcXdp2C+IkjH3XmZBiBXQVwLL19sLE2cP62WdL/TKOJmfyOokYQS/
hNzUZ4ztQzS2qvRoDfohLEFtSyngFMS+/BCsOR+bU755HFt2mf1be6QXhYIJRMH7
lverVp1WoccxclCDtCFmQHHjMx5BU+9BIrpr9bqXTT2wUqXgmHBC9HKc58bHeFr/
w1w68OSPyX8fttiMsVeY2Ug0rrtkkcsYggrC1Ptkzhjx0KcXDgqpkouXcZvCS5CG
X4bULgOB2KpeouIF+ybMaNzGDbnZ1pwWAe72B/oQxQJMheK1KWJfjiRLkZ4LOW2x
vahBIls5zbMuI3sjBgEUoxmNJXkXftmg/x0GMzXPkilvfcAjVnn+7CcO+CO4QKJY
DfTD18DAGviMwHw5mJQy+yR1u4hVDsPzCf72fGhIS8yerVqhkmR2fZI9A91q0YhK
4WqhXALXF+LefuhJVCCVnx4ZumqOwU1oW6heeFeyslIK5ajVc9somYnW6Gn0UUbI
YvR9qi0oKJw1V2Dgkkh8aWe+McDXraEIBArfm8xQF+hyTFYEsm+2MbmFtj5RcGxL
wtGiQUmm+YqskmCvzsFNM3XAkOrx0eWR4QDXsYi8KWYOrQ4JpBe2AitfiRtqeosV
2G++smTcd6nBBQlye6+S38VDKM2SyWas2omhyO55kvFSYZXgLnxS+/gWGdQ7ONIn
1XZchZffui3GPhSCEz+/lHfCOhx0bbd47LKBSU7BhadnHnALAdToEIUqGX9u2bRl
2OGhZHBRbAiajnl18H9DtbBC6ZMKQHT1d1bGLJNQIFgTJbv8qdPjipLiIlHE+VLU
neEI/MgOGVYK9ynp4z34AF4ofwR7Z4ATm+dUVUClrVUuWMVUZrsR4USgGRBP+GIU
8jkdy90Darpe8HjPU5yxngK4NxHGKRCceGZ8Dror/ptGsKPb6T8wxCZFoCeLLiAM
SWYjdFkZ/+jW4muWNZ2kN9SbEWVU8hTRrPDG7y0W0iAiLWNJdR6p9JtpAfeB+Kmg
bsjs3/V2Ecpxiglw9izFKZb0FOPqvmxCXHPalIYmJgVSd/gHkQcEQjlQampxWCe+
Ju3SfYajDhyNMsF+yct7xUTs1CbQ23S9Yzgx3Ol4v4nMwgZ2QDZXF/HJTmNpmX6N
GLzuaeCzoskRNYql+dB2W+AoRYaw7z/a20A2g5mcZZH0olMknOp1pIGt5SSRo7lN
vfCY5pDqzaqkEUlR2oby9zWRzk8gt2k2HZnIs1hCl8zn18NZbGtlrMNsnE5tyKYw
jkaJVnsBE/ughRDLwfSX1y0ee8B4v2AVVZRr92/yUXzBQ6xz1OC10ungl2Fm1s2Q
tOIB8TB71yh9VV9Ue66wSGVQ4V5fb6evI3H00wX+NfRbodP2Jfrk12s3eIUG2nnH
hNoFCebgUCMcr9yu3tR1pEZ/EOh8BVzEaz/cDc+ARJpcqaY0uSgam3El4JSz69vA
6zAZP65n/Kk50Xsro1mR5fAQsr52+2V2y2+AZ9cXaPSVyrPhb4H/Hvr6CpztvDEI
bKvP5w2GKy1f7n/Q78CcpVy8KDH+Ox4/S9Hjcyky0oR/u8TvBKIFuQaGTd9BnE1M
29D6LR7BIVnjwFe0Q9AS7/QHGcM/zeIVnHj7LAnLzywhT9lo32KJXTwNrcha7u7n
GTQp1Y3lPOClqwvBkVbxK0cpcqSu0lB7Z6Tr4R0c3tGhrPAFfF6lJxGps1ivCirq
PCkZ/DNMPpBZbD7MZO5HyxIUYQ8ilS1hO0suRNmoN9+bKiivsHRnnUN5q0wWBSej
QDu/RxxP8sLoA0NnwaBUwpzX5PLxOSkrRB40I+7e6mtuWRk0bknkNx849lwGPC1A
MV9dX8v3q7DVcvuEgNTg9Ya9NBX+B4GEW7ygMPGOonQIwYlCZ0FejTakyHWfw/gi
fgC9V6paM9JHd+cytl/tOqbL9pX3SpBSqXjZNubbT6qRXAnWTiTxaoe+AMk4BmBl
ARzNqp15NHjx89M3ZNeGzvSChLRLIM+pctvc7FQrQ8YbZ2z7EwcJbn4STtowult+
QwQJtFlF2SvDaa1W1Yt7eO55XICV+OsHMgdnomdNUKFgFanLPYw9hwBjFTvbibER
D+dJRSTycfTkc1NAmacwcDhu+f1LuAMaCPXQ3s+C6qrkGVslzQibStO2v4Redhd+
tNFyldz3vmwXSw6FYXYVPRwGzHQHzKHjCKjCVCnrxYiOjop32ZLWem7pp4hyrJ3X
OWpIooP45NALOFkpTcAsYERi0giQgDY2FRqmY0UGoqJ0s2JieT6Mq9mafcEJe5Lt
5k24g9MRv+pWr9XCWgt3qm6GocwZZUjGsbvx1P+YCC2pcdwQwswOr5o0zbpndDLS
OnfuFj5YWiVG3WhvTlZljt3qCitytpqvGvbpbbpQPfv5I8HNoL92ICX7nKwECi3w
4evtH/gKjqHQLmVzM6CCBZcOfxK6nFueKqsZgNiOcNyo92ozdKIePlVrvCqeg5qk
HZ2KAD31WJ1Zg7UaZC6CKSv5lLEla4afWRveM/KcQuqxFPCY8TC9YST8Jo2YGCD2
7h/xG0QX0WD/aSTQn9xkkigvY+oJP72DxDxOBT6TlwDGFvHQHYl+3PsXOb2UrCAD
rv3mZp7mPCTwYkx6xXHJ3WWbkPkuemFzG7gfsuveaKh5TziuXYtTBSdP6vmsDc+j
AERNenwQvf1HLP/e+axgTsND9/kkjVvNBl9/dSLOSUEQ1HIHq6sz5pfCtR7jl449
DPDYo058QdBSMe4uKVwAlGLkXAUkI15Hdt+lq6HrhzBTuVrNLli2ajyXG8jAKem3
pKCzMlCpU5GSgF2z8KKtQY/TwWOSasojG49yHo0l6+hfSQ8MYNxDfMPPIXPb4D2H
QP/UsWMcwbsYrgfUweUsMbgjRsGEpSlqKl5DVi9KvJEaI968tMszlkNC1lPaHJGg
yVL9Aka4PaCj2qFbrt4XkeE9SFTLRbTtcq/6thgyAl7HQZ3EzIuw7CVgHlMzJnZ6
NCStnNMCrJvLPV1XXKu7g8RdEONyPTbRWoA3nsYrSuXBafglsBGFRLaDQS1I0c12
ETJTd+qKeJBtTJL7Vn/fZnNh9xERoAt6UOK8LQjesJb3ZZr+gw49LKewcwYQ2iSE
FOehf4xLgTTchvzKn1/SBZlytw6tHmsdvUFPVLu32lYAcWoIHLSM1jbWmJzxX5hO
OLYEGXxor2MkaDcuQCXp25q/xl8Ldg1qkIzauniwzCxpW3SMn8Yo9Dk6fpGTtck5
jRueXg1nZnmoy9ui2PFKlHo9sx3pal3Ew6hWB3ArcY7LB7OsGdODcevAu/0IwBfa
DmP9h6oidqjPyuw+JDsozvRaLQNxCcBPLJSVGc8IvFP2ZsrvZUm/PS2dgPhWQ2lJ
klXhxFtg5sgfMNg5dhajl04XqcwT43Z0vvUtdqmk5Jw8e0FaTo7ryZI/754R3U1P
CwdZXTvOqb2LPy8jYARDY/uRoKARQAx8Azzc4psnZWo1Hz1WM98QkeFPEcoKAag0
a5Ex7YTuGekDcpTVezHs8zaXlU4tn5ZnnTtd+c0RlwsS+dl0I8irSvKWQLViJZd3
X/gxZATUHzQlzFvfCRV1dgtwDx8AZHa4z3Nqr7RWEtupLK1CPyz9Q7sHQMPU/JGq
ggnuaXG4yZfgr9FkOCPbye7TcqhTzXCkfT4XTGw3cfvWpJU5L1EPQ9iMEnSGUZoI
eVVZox/m2ajQFMqj/E5yV1m5FXeZn+x/FuBINVDv8jnWPQe42qLpIFO2MXrTn/ia
FCuWga1lMJ2Hw8jCVYdKDUrm7THHqf3NxG9jslZ1x/vqsfKATs5JN36QD8D+CZH/
Q7kU/O45hw7kxxNyMmEj433AaqproOHyEg8Jn7GHq2Kja0Tjm6z6TxDwYoG/tyO6
BfW7Ev0e24jshT+UN/yPAfGg+jAcYU3oaLHkVo1tZf9Q4oqB4GoMTISIRxKTlfpB
fY4PUmF2kKnSVCTUF+lcuSy0v5s9gSCBjWUdPCKqX4L971wfF84Rv3CLpeLbsp0p
IIMkH9pkxzlQOQWfSbliDZIkZuGu5iquqBdrInupZiHfu91VviUsKcNRE7TuT7Ij
szQonG+2ommw6Jq/EiTaeAL0rdF9RuXE9rXyEdF6Tj+AAxH6KSHDBCkzupJWbpBR
G5JOaNwy9hY6aR7+5+BeMdgzi99kvmc6X5hpZ00E8O4MDfNsfghT9iub0k7eoG5i
cCASWV2bCNeyszS7pHUpyLHi3SdAAtqOJVkcpPPyeEJayW1sdQ8isfMYnG3n9I7V
w0lUTaY0uNVuE5oXI41tm1T2Yd5vZpap51puY5qTce9FR4trRIQ8qWp1b4JD7Vhh
sSaJbjEMQ69Olw5XpzRYizcdm3nscBU9Rn/n7QbNM9AHg/Vpd+ZBr5u+VbnI7AH4
grGXJjrBGUb88n3gbGjgjF2GLJ2+kfVARzMmABbgLMXs7zvFA/F2swYvgzOIDxJO
kqhkjzSSB7XD6GSlSXUvqVpF9Mosiig9VURavCY3JmNh73infTKfiaGZkzgAgwhV
e5GLqc7if0SvzkqDNC9gMH+0UMNdygFzjJUbPYR00Gz7wYlpGxqO3SyPcmavSZXQ
WBK65WVDCd25qVFgojYXoqeQMGgwq9puRHHIjjBRlpmxKpC3d5sUzr6Wr0jnbAtc
LEHwPQx1mlPJYjClMQK5Z/fPrrosuUPIMrvTp4CpGktcmmaunRzn1RDNeSRy5vpN
ti9R9x/8NWtZD4GfpIGVT0cstPgw7xklKhlmkoEtzOGP4QfaUrpHz1X5TkcRgRxu
SknwinYX7eePSiqRedF8PgoJo+OYf3Oc7y2S2MVLRu9wkNW/aBrsGW92pkxLyAwm
8ouC3Zdj5SW7uvIlwsi05Z0Nc+DMGj5Gtsr4PQY4MlfG5boJHaG4fUqoRN3eYElt
oZAABirR1qoRd/hAUIpq8mHi2vF3Cy4hnze2+RMU7SyRjdgor4J2zRAHDfLeaAF3
JIbuYsy8WxFWjxcQzCERq+TEzNNkCljK/hi+ObfHznVYMwZOEhvLwGrLNod0RSFj
68K33DZiHicdrAK7xIpiHQuKqNUkOzLwtAIMbpncFk+3uMNDv984hP5NtkuE2mAR
8WDXMZixQWgwCSzSoz9Mdp+JdLeA9s6rpXLIiy/ovyx04jTfWYGVAFgh/zW2zjH3
4TjwKKvPXtDEbsFbTJdJWXWQAxktnPg77ISMwYRKYeEcRGGs225/04yPSyQvlopu
oHm9aQ/hvCxPPM3KVQCYIHoCkzbQWIT9YUIfz+QfaOuRNjobJvxwhJtCTE64G4Wk
iJWqjGUizzejzOdb9kFvx/nTjgN2M3zuesKXS59jjNTDz+JykmRRW0ITz7sfpbkN
w8RpxBICmQHXWXIZ33Gh1PuCCw5cTEUBqoFZ8UKEupA+S3SlYY+KU7jz+Ejm+VuV
9fLlfMVMvFZ2GIbt3ztdIXYgj8nlzvWGRgvLdKmrj5QDhUKz7eFUeuuXRD6Lndyg
6ag4sv6hVSAstkJFWrh11qZ9ZUQKlDQh+FEJDXJTugHL3BlTXU59XOfwgaxPK8dy
eKl7Fr86l7Uzhc7yvvwZiT6/BiWaKCcPVIHCNFfrITrixMdxoDMc6VpX3tI9qVX0
i0wa41d2Mr0bDPD5HZ+ZaEJ1r7c1hz7i61Gsl2o9NR0P14Lzx44nRVgbURJZDDQT
6AP2pQZA1UFPqzgOImeRpLOp95KHbVmZF3NWpN++mtseyjh6VtRai5xYzmtGmey/
58L+IdTopwYR0ME2mfcQV4JlsLGNi1KqbFvA/wbbgWsCH4bdk/urufWStJAJI/Ny
ZMi7a9BVPNdCWHGo9mdtvWtJXQ20/3xy8wtnZt3wAYJqCow/HDzo8RviYht2AwnI
Kt3gqmmLAAPSXfdfRv9IDT3SF1r7N/TQ/ExTS/T2RIwz1ExhfqdCqFVe4XzqHesH
BkJaK4wShHBgZT9NJ7toobSHvgdnJk+E9mq6vy+KWrZdzk1BZybGHUX4L8naFDX2
gV6HiII92tOQKgvBPjDqUGhX/M1d/cDpgafSc+x/WRMklagbClLPC7Wzsj3jtdcy
yhAU1WK4Mml6kWgJ8rFq0wQblDSnVko7VyyIF7QkISR3UYGzewUOjRcYPtRMEgWy
iIsimprEiOrwnwzRpAXbCJ9TqL5zi/zMa7DFem6QSvvdeMxqMuqngaUIH6TW07dV
e4CyPkQJl8Ovp7+4XS16+mo11j+QuCoayG+06gxjEX3U+2lCWvpAWicuOYNNT+k5
ALvfBhPE9yyZ3bEj3ElaUzfR1zsd8ccqAAqAI/Hh5BzqZRnkcOQ4lqXz2zOv0HTd
Q7wWZfQZBDoYRCje9mQlDqdWgjtqMk34sXBVEj4fqYJ1Y7WZ+ETJKhEO3QJOuuYR
+LiVG+BskLE+E+WCW9gpepUKCj1g3zHelDfOz+1AnplD0F0CrQG8rzU7S8PmEF3v
eo01wMZ8HMpBHfYujv+xRTDJ8DXCVpaxa2Nd0IR2gYfSlE1OiedtN0AH4E7Kdkfy
uchUF3Zr9u6vg5fof6I0kqTz6AjTNKIgYFQj2dW/pHzznjJ9/pPf6zLCfctKRgf9
bBSRF5kCXTAZZA+ZB/JniS8g71yALnyx8+cFt+Rse9VBORJqAboOzKTr9dQMYj8L
AxYzkafWArETjslPoawFc0FxT1Xiw+aunt2sFrspA0ysyJFTL68LYJ0/gXNUrf5r
3ttIspJRJknTrYaNumfpwYRS906UuPRIZQQMIUBLYX7M7ZscoI8XN3D31wf10UFU
3bD7RStQMqxSQtEvmSveuiLEukKZx6LMHcGuJ5R6W+rUFxmGqUtYx4irTZaOvbh8
86W6qgrlFhohtocYdBLQ5L+YnMAq87vHJJmSnS6AAStTpTaF1yBjPFLohGM7H/Rs
5NQMUTxx2MBO0fSnAjGxjS9mAZtZD8CQPRBCwLZFTIfn/zwYECO32aTxuY1LALnE
SiwmZITf0vfQMR7T7HfCg6YW/h63IkyDWazxq/l+9Tcvy2UBik5WMIRy7ZkG0KL+
SyDDVxIu/bxvpgitXftMC0MerIbs6pY4EfXcymb6I96rRdiiaHcE0rR1Ys3VF1zo
R3wQKOrgVeBk31g5o3LgEKRJO9Vo1gYnlbh5MO9nKP572gej6Nk0gvAWYftyldty
MYOoILIguSG1SsY8MmctJx6cT8+/z9jl6zzQmVld44z6QkM7hErg+oSXURRtCTpG
2Ys5Zx6xhxMLWAIyiRZwDNOIm7yf7r3zRzn2uM20fTa4vej9kWFNGGrPhgCEOwX3
WGc9paTSeuu4DnnsYCsjEYHdhGjyea02QRQv0r+KVwf1eaLx0uxlx+Yi2RR4l6ww
OH3yQFBswnkyagtII1ccuUqBAOWVaN7ctcpitRWCz3ymVk5jnWe4H9Y3K7oHehGZ
kBYk9U8DVBTKqyryRQyGyG4DwTsPM2MRofpUVnexnkBAC9BcUskRCYWUM7wYOF/W
H9W1au+uuSJPN8wPro7cBk6AqvnaRa9YDXcFmJG/xpwfmLhLYYpmeYD8iPpUTJ4C
kLrMIyA4CiJ+SAqUezRHC6Bl9GEh3Tdc10TmCHsy0zrVfZmF6eTU+JUyWsXlGNUv
84YkDbzi2h3wBD8yCBhvSFWiBRq0+e9nlwBG6HJgJ+6px9VJ2FxOncYkLtupLl+B
ikSNWLBEohnt8pCBxOzXcz0OQeKJo9zulX0AqYWchbh0dhB7zJ8dlG8iMnsfeLdH
df6NNIyq0/rbEW7M5P2kQHhunmB7Gq7qri/etxDSDmfmawR7spIBgJxoJsldQr8K
ZxHg9hHWJJW3UnMPFoDDYFqzjGjgB43YTRswvv39TzurDMFWkcVVxpAoffdzBnDr
QpCw3qozkIKKmfptYOVupRYF9gEb8hLXnstNE2DV55DOaSxrBcC3qCUs8ZHsA1Lc
6D2k0pcB+Gqiv9zRFQ9UzVltBbR2elnVM17a6NkaKZgJtOJWEBAEKrZMQgNSxnDd
NflYnDiklREKwpMj2AhZL47PqI22Dzegy9KWjbOCs+JcM6ba+5mJNpaTGY4NN3aP
zGinDae/osonZWW0Raf9ZCijdcuSWs4n0PLitaruRm/oTGe6Fk76OrSfNQxwlVrn
3K4LYYuTlQlY0yDNNcleygaNNmwR+9r9oZXvz71RRGjIv+5dPClnUzOYCsHrAL/D
QkqwcmT/mC4iNTaZn/udXhqoZXWK0uYXV1e4EwtYBS1SONt7I0p/IJ6z7ZR8wGu0
UWE3WaBAFHp7Bqp/yBLvDkfqezjMKZrmU3U2JOxsjSmvNjpkJxyHXxfA1zAPDUoA
AQikRF7ONRmGuSUtEsPu46A/B1Gbycnwg4XJKd3w6pkljWjfQgS0aCgFToKzncBX
Ru74N7ltphH/G9xdKWhpsfLpWg2gs75GkxlPN8zvhiKS3kwlGLSE3L60g86MWKw3
tcykQa3X7KsFC5T2cHJGIgyasY1MTBIZWvREcn7TjixscU3VeE+bbtCyANX1GlEg
SN65yzBeyxSnwik+gsJYzFy6kKwiobzi2HbpyWr4/6i9FyEB4V0PtQejOowOWu71
Q9oa10dDsmZvtDg4j/u+Qa6Z/7g1qYHEr6JL9TnuLfLwzni2lHF74p9vYrclZnXd
XelLB2WWgE5ng5xc8dxCJmqILddReb8EBdkqb46ya5oGFl0uOq1MZpHWZE/QpnJR
uLYmfPnMLURREq6l2zYdHm/DnZ4VgtlUgaXeExKTfCeDth2XmQy7JJrSu2raEzxc
mWoSqGqu8KUtgQf+s3JXtPpv2/UyR5KS1TqrBGHINVxjS+OFJD9WgOML1ZYFD28q
xKTYPTuJikGyeLNsr62x75LdFph0/sEThpAv5E/K8+0JxlLh9Agltvm+RHzX51V0
6ExR3ODJ1XsDTF0XExI3PvswuQ4E9vaYwxpPOl7qpX5AQSpl+Po8R861eAJYO2G5
Mw/6b27noiwjlhA0vwTMkpHuansNawSmwl3DWzNcvHr+R1Z3j3ohSeOG0EIdTo/i
Yl2n49mmnDmJ01DDPkW9jTAUmfYAb4VWGLot682SLo6FexsHG8/U8S34I5aSknep
wBuogZh+26UQekk2WWAcy1hafvG5Pw8Y6AB2pXXB4BonfOKQ6yFyMQj+K17ir2Q4
5vCpTbuu5SvbQEDYIJ48C/ZRNiQyYNny8nRiKwR+4QWlhJ3vwFCk3LmRB8trI2jz
7cMN/ul+FB9a3HAlEfJk2qDgFpCILSurztLIA7FP9cJEW1xrNOriYjrYC1AuAA5m
Xo10/gmju+KLlgj4pMMxp+Vcmd1kKRDhItpgd0aiHu9uU7/6SosjJO7h6v2SztCb
2cnKmbLHtgdVW+TsbYhg+d6DzFkxLiqVLhUmUGJjoRWWecFZDxMCNRCrY/62D8Em
5T0dQEuMQ142QKRANVDY3Zd3VODgJH6FMEUuSfhlomW/QA75g9aDT1k7m82m4lJs
/BdI5cp1G9slqoltURG/K/5N3TpVKJS1il879CITsCgZtyEQGK6hpO1B3WykQp1L
rLYyYoYyzJLFP2os3vRFXpCD6VRNBwDY/9YaV3jDxhbkiXI3exsdJr8xy3oQlRkC
j7wdIL7gc8tPUEvG8Jtmrn3zOGMjY/ADPaTKT+H8EYlkymMMAQkHD74aFSGoY29/
8MDBUXe23LpHh+d0iaG09wLDEArMflQVtFFCH+2Ed3P21oiLA8x8KP2VzUPbAWlJ
qr+nFUua9bBw+nLWVipkQZ0dyVD2YKlXPsO9dCIsv5XvMmKrpN8a6Cy+kP50DysA
l09wiOpl5tE8pfZDrE0Zi1TdM8jRQnKAf1WxkkU1CsZLcDG6ATITBLrDCeQ3yo2t
GguOq1WHJoZkZw+o8zG6Vw0w4tDcL4Rw4vcqDNx/lYyH/bLlY0tfZUjbT97k0SCB
mFsy9qOA/CmQpNxOWD5AtLsHyBHwRn+JKqx/NJWR0saCa2h0eTIBkh3KF+axFHB9
tKcP/iffBihNFFBoIv/VlQmX+tZifrWuuDysew/v7xn9IZW3YSSVsrXNH4pR/SxC
0li7Pt9vs4XjksOEEIzXNq203GpPWgeoVkjJWbLLZKWGZFKQDAWIH08AzujXJu3I
jQ+bEBrhsFScqyryeWBg0fhuzU+Icmjm3/aaMMgHWYkD/8bqLNhLJuldZMudapVf
A1MWssARqPexLbMITiZCQk0qxZd+HfeeDYcqn0f7xVvJCck2eF9PpzKf8yrBfjt0
SD+I0Y+Gsdm/Fy3BldmtOS29VqF5lFA5CAUyYJkacE9hBF4a+Lh4S078dL9vGNwW
dzEswRhzWtKRCUKw2xk2w7krcx/aCy8dMWQja2o+U1P/Xzt1LPF37E5eJuzy9JBt
a0b5OpN39xgVUWQ3ZoaGISpqo4YPp6loJI61cEQZWcPw9FkXpgdAe4mwOXSpnKWw
bszv3PFZvsNmnh79OLZF7JDPOmDBCf4+7UODJgTOWiZj1BehofkpzhPlE9CcLoaE
X1xVVxNukBfewNp3SYIH0ekcdRyXrO6dPZJkPYNUF0BIg5dSx+kPQL7b5c+UG2Pt
nyzNmsYiu0mj8dLahwcJR/weg1tsNouxkzFUQ7hCD9lWkCRTmLFRf/AHVIXj/U65
mrtke6UvTEv1URN939tckP+8LEg1rNhPDN+JmIEZXMsLo9QE1lzwh1GE9L/MYHTY
tpRcHk6egWgC2EfunZOcFB6HWENSQsWP6Elwd/OOu7sS53c89QZnrUjuH4Ivhf48
abUJyEsvlaELBX+OeKrMSkc55RdhI45US8f0YYXk9NrxSq3ZgvHMBpMHyVMX2tGn
2YZIxtkp9qsY4hwe41dXtW/03dyn2lvZrRRPOItAFMasjW/Xi/xiwErhUBfb0bYZ
1IjCdvtbqQO8rr7bylxcA9780WRBT5clycafbSXvKVTWadUGI56i+Tr/CcXLXtxa
pwyIuJL8fEIVOg+rD1b6usN3RnsBtipobE/1L3UGo2+eJtrp0JEvZG8mZTwE0t8/
MuJdey0KoEq5R8NEzelo7AL8qTTtMo30dJAwIEDgvpy0t3LAJPUoPMWFCat2/Rzj
RMt9NGJ2c+vWhrIUoZkReL1YyiVeU7w/dPmO/dRi0fzsTi23ecMfPibwGLza7IMz
jBBYSxNa7iq5C6sL6jcVw8TJXCed4YDog926oH5Wa/+BVCk+lhoyvRhJXnbU0O2D
ntC9E5/FAk8xyIlBKuzTh+NQuhDAQh+SAz27ip/JtCLO5EvaejIY1ciMGKzvb/qt
6EUiHokKBqM7GNBTrUc4RKEnar5BtZJsmTgcjDMHeULaU99uCDYpJKkbwUUW09xk
Z/V2tpYn1s6aWy9I47Gx3WXlOp949qynFPKbBr40nI4e7DityBzkB7ETHX4H1a8d
HnaOMjHX7lVqpVxQGLQd7gQvn02EISfK21ymwFluU5pzAKxKwoh3AZC2kUkYF2pH
1wrzElqGPoy1uR8wDDVOuWdR/sDJ53bF0ZyfKPGGBSvdYXZG2+BFw20kZVcs5sWY
Yt7YdUu5GFdd2rjrQpGIOwwOBx42jqMKiOZ7KO2t4V3j0zEkm18Tf71ox+1RB3Sd
NfQjxnjYO4nNxmhGxUyuveinn06hJh35+3Ux7aTqTBImgOKS8J1s90BzpbOW2Lbi
K3lYFAgb1lvaCms2CwZnNLwEVUoNmM8g4Et8EbhkzVitQ5cIzayg1JumHDK/7s/A
oVK6NcFphQPDttnO+8snuJay6iOMQp94GoiwtJLgTjaHEz2vCat4i8ZgZWG3g8sd
JhcwwJrYipHpjkWjIiSxgy4LLiIfZjiU9DXRxcUenIBuVI4LaAaDNE9CgIjTskEY
0dNw4hUkDuM5fqJrg2Jil3/9kyx+1W/tliB5BA5O5ZsqbAVeo5yDvvUhsD18ChX6
XJGVoqQ0+se0+mKrpH1JgNzlT/UJZ3X99qvp59Idg/W5XlZuc99hG0sTRiKWgAGH
jtGOhXUl/NrZkx3bRmiseAaezgjEoVwiua0scV9QeGnTv4IlNGoRfODf8APAqcAS
6Vh1h/wAqGL9CrHrAYb2XC3HRA8huJAMXpd1RBqbT3nHRdw0KFftlREt9Uy0Ig1q
Y8PAbyDYO0yFBIeiHxEA3FpCv3qCSyO/abaZ2SVbn45TWoyocBjkNVk9hstLQ2Qm
yWjMFz5knFIsAeWCi7winga9Y2fyJRl85itS89VFC6Ue9qyC3aMguB5JJWAXUjV4
s9ZSoy8SDKF7/z5gnL3QA0zE3xDEQLibp4e8ejd7/XUIw3aGXhjDrr14UOFliHgC
FpdrMZxyRSW3j1SbNefPDqY9d6pjxO1UV209yyroIFG2bZ9inmtchqKHjTFbyFUe
L4vGo2GM0SBv2s3jg6NyjgLRm8CpeKOJsSvq+lSe9no05L2MM1NYV9oTZvyEQdwb
tNHD+OkPeyH2oEkk2nXuSLN5yK18/BoB63J5FbiceXTXABZ2COHdBE5b3Ys8rssa
APxtpOeQBZr91Acg7mqTCTXSLcwRTLNmw3rHW0YsJ+0BLG+k1TAK5ISa9waz6st6
Hdu67qBy1DAWeR3H56dx5oLl7L0/Ew5fNfn6/e/nvRWu306/CLswhKJhytfzMuLy
7COn5r2ftcr1mNC6CAyMiGKembtNJtM1bYSjbTQAzHx5hVP+jxG2EbjoDHhrkGVd
UfIKZLq3CByrjVQQW1T3WwNyc2HYdAD0WGtus/K5MkVeazL/uD/bM79sD1wnaoyV
NODnIsmLzmgoJjjnYOXFg3r835iCxCwe+sF8qE29UUAdMnUm84gX2Uuyp2txg9p8
Xe5ENnZ31MDn3njUgmCKdplung3uIQjiba2pHs6c6Xd2zqMBTpkJk7jzDJDTkusC
8ehvbDwP6MRO9r+XimEE+VAnCZE2082s0Nzt4r1GbbDexP8dU/HuIcy45ah55V69
KG3nQzml+H9S5nAeX1HD+iG1q84wiN9FmtlObeH2ZzBNgpZICEtstcyumdGYzr1+
m0dQSkRLNF3xzKcmAQQeU8Tvb8jLI+1RG7ezyCiNgNEGzjc+INUwGxv0bQRsV8sm
Y81kNxnCvAWF7j+19V/n6jaAbGs0tMjj8Ruc2Ay2XXWw73twZLzIBukcu7H9M2pc
617PeqZJ3R0PTBkj85Q+Ws0mKGz41tFOmwhgilrZSOElr+4XGDp+YX+z7yBltX9+
tLw2LTBPvCmTo1f6RMHWvZswA7QsWb0vQvI5vIUfup2zl+ybAjXuWKYBAHLNVTK7
NFBKbgQQ4X18JTSS6Jew/qrga3pMdYG+VC095LhsyO6tB4hvhjqNDkLvaZkysgMq
6C0sBFgtUnCzUk7a0wgdxHA3mrSUcWdqIfVDXUghGovszFd6eLDFqDkllbY+uc1f
PqtSpyp+hlXSQm3zYg+OO6gi5OSbxU/9wbusJB3rkOC2JdglDONPKXRocBAoQRu3
97fzfhcJpIAQEupAUgPr1q7nWH6ef+EZ/fOSiuJMDZm/rnoihSergg7L+qblv++M
LLEfewu+/SFyRVgqHnVAj4nc4D+reJ0MsWmunNP8RdxRLNQNbrYBQWVmCTfBpF94
ExsxdrOs7V1ztLTWQjDMfcGO/52ZtvxwpkDlfzU7/iSLNROUv5OSkctZl1RM2Yhe
f6hB+oAW7Yh18LPWdtDLNv6yjhnVAVO9WNI99ZAKJ1IZU9mHhacImPmqRGSd0Yoz
0035X+sDd4eIwrhYAobb8ACIY59lJ3kMOsBR2esmSJ7tEoYtf6wYvti5ph6xGsZ3
uNmD1dTYKTWjuCjyhWdoDa4qhZxXG5z48LyKZX32CjbiJcLrw063ONFA9kaMBGq2
yqTQFQNdEaUKgQYIANNaUVXIO9PTR6UZ5Pi0aUJ6NLHgNCrJcizzU6UO8XZa+CdJ
NEoS8pUJ9ebaQUinmI+8ND53aMo+vYE7KuTp7WZ59G3vvrmpGq0fkXIJS92aYzp7
LN7TPMyPPh6dxfZ+Mu53OfhzQy04a3c+nHChpHIbM1+OzlGvFUkAIUU03gQcGb5g
UKkYvfdcnDpl8iNQ9SYMNLLcDSd4ENwZOQpRkGMWPC/K6vHHZ118HpWvzeHonwn0
QyE11K/BEvCb/JjunyLY9f3UiY4Lqsr7XldWo+NCtQC4M+G6qzuG1a2f3kzxOg0j
7s7qeyECfWiFCr46mr0T21KBnOU3Csvt49a/JK9GLK4FXohW6if2vqFBeVFEMVk/
f8WyIrn1G9NW0bsB/oLBQMR7eTOvyCc8+EmoUXPMlglMdUK6WeCZd+KoLxfIRFPF
wo0IE6LNOhLYt1TSp4Lsg4RloBten38Tf/d1yHfTroyQGg33X9MxGfARvGXxVZ1U
eO7gzlF1Dx3DdZRW68EX4Qk/4z4HdxmJDgNMgG7IYsewnPsFSiqNkwFyuNXbM3pE
I5d+n9gWKiCC8p2zQ3y5czXtlroo6gX3g3eegVUAQMwgUUj7IRuLVCkGvo4sviDO
9RNruwg4u1yOwQ8pcZBJYww1FedoDNmsD6AFa1alxg0WIgI0qIkpRwf6b+YfD0Wg
jWrRy5Bqarkwd8p/p5S2i0TRMLO/DqOXQSrpEFUFBp2hcXfQcg38BXtTXEeMqJkM
6vte6ChaOcKkVwi/YRiPGjsRcYSsKkCQhcKh6cfl3gFBMLtfLNrG5iRZNMBtVYZU
i2EWdAm6tsaThdQMs5YQQS/ieUBMheA1nVsAN9CYu2V8O+YPNc+ELXmKSUljN9a6
2W6yoZVDqnfUt0g8aKv5doj9PBh25lkghD5AdC2OXiOIR+Xl+Ndh71L1KpmcjW90
w5CsvujpuaPXPb7uORzgPIL+8zz3s17kKe+zEr2CabTy1v4SDf3tvVjG3mNcQqE+
gFdBxBkbc9CcPbsGI79H+lmYnrOFfhVJQ3HUzxKRH1eeOjHxqDTQBAa2WbiXibRd
8HwSYNqZ8iuuG6y3qKxaAppN7wzd3ZEbccHSf6VGvCMP/5uswSvdG6yiY8gfvqLu
yycrgicDCL93vMZvjPkxiea8/CuCCQ2iTqg7rNvWvZVzB20iAxGhkJQMExh3Heta
JMN1ZvhVFcEw9PvIVHnRHF0CP6S1v3S9aHIr+/fGDGeKY4uyO6SlUyxSMwIU5qpQ
aLMGyiyhLAEF0kJMpHSKGByI8NV09y/EOzi7xj/C1o7S6poK7ufk/0vLihfm2leO
7b7IGuzpgIKjZgf2SJ2X0hshIQNyu3PQeMwsmor7OnfClT//bfa02Z9pf+LvrkPf
V2KRB+d9l8je27y+Mg4tvqHX1ipBpbPgV0OCsNe7l4dpW4kxr1gc5WW05Ag22Mbx
0Ldr5iH1yp+x1t3C964NPJIQk5O89fNMUHg05WDW//WyOv+RUfqgjrnvV1ph9ihG
VPH8F7vX/3iZ1PPxI/wzx38DIQryIO+qUqVz/en4BNh6XZkyLqWmVnPT/67ZfJoh
NsNjk9lnf00wYhdYZYEu8vtmgZa1Tf3n3A7/gdZdAIVtsFFZMX8a/tZ3xV6psnnI
nD821ZOBg5JZSxkDna2WeCxFW0zS4rgTP61ZVanTvHenuDLFzeAdkjQpr3ueBiEp
Puuz2djZQjvicZ2bodyh4ciMLSwcSk3/AtGWeVccWmud7y/hvqDyg5pP9NZxDqv9
UEVo3vUAAZa8hC0R2ZCch6zFvfTTlaiXCnArY51ekJ+EODbwGggf74Wl7D2dViQZ
2HVV5L04D640VxRdOmInKIg8mDz9bHBVEoAzgQkRqtR7YeXx4mmI4xslFjOY1D8T
WzsBiJxquX/stEGIP3Fk60skiUFPkXoX0t5EVwPSWtf4UM47OcGzZJu9kW324LE2
CKwitiw7UjEmau84nMw6RieBmf6WEpqz85COPpAkKOIrrXCU0ii5L1QfQxHgrqVC
zixBPp5rjHT2GymUTTNN0wPf+hZt1e9iTfAqrVx6kkCQ3d6GAITp6kfIEjUFtjTW
WhZ/PGO3tRkYs8d2wxmGhV8WPYbseKe3DL2Lr5Cn3XqfFs7InNkn8ESnAP2I1m2f
Ebm1h7CCL4O8bezWUE+2iSTz6nG3tKHaf+2TSKMMTz6z0PbtRhDz1PSiymFaJZT3
Ym1yGZmBrKcRWf7sD8qFYYgH1+4FDIl4W+O1ULfubVi4Eezz4vpQffZDoEYPKqlD
emrhdQeJIw12O7+nkKhUvr2p8OWYcJMG4yKbn+/jnJpjFL2caU98GB9V6RSUYCQb
qDQhB9KZvrFTe4dlDsQNUdYKXIv1k9hqu20agAVk5lYkryG4D8qeMhRZIXjBRPNF
/Sxb6z7JTQvNjrdJVUJlZOA+NuegTTYSAuEFCbMNTuepowd69cD1889ZC4seNXrb
OU9lUw1ZsCJBRPqcQx9YJ2gpieFDq+h1NLnucEFlsx/k7ZbRl/UV8rgtZWb76Ubw
1FZFapHE9tJmoP7+dRTRRSt0blJyZM02PFbCtE+HZg7eZVnFHlGk2siGdQlI3zXs
qBSxRWpTLsyDkP1w8Vq3m28zj7w8hoZ+R3Oupk3svQebRYqJYcJSarO3MzGgx6ME
086E6fS2xiPFMS7nKOZSceWEvyYMOJmzs61k9sYHupOMsxA9sIJ9bPuchoyp60nq
x4FM8Mi283oDnrUGs/xfOvC8LfGHjLywlP+5ZWwPl1+ouWZ/+5ef/PWSU/MUrRmH
/dghXwjPSbnNAHu8h0YpWq7y78IdxQUYC/jtmdzOgH6ma9430gjPV2qRdulDdyHe
Z36Tl9wItlN/3ftq53p7p8U6LTNDHxYjT4Vm+3I7mq3KDWy8a2qMbnZoy1FTBQcL
zRYcoQT00XVAoBPQKep3rB6g/bHDL/YiC4AlhrRHOYe3dvDFPG6wbsDdPL6nvU/w
TQHAC09dBNPW1yDf08zSxd3mUaZgnO42s+voC7y8uWGwYVHT+eddHwbPvUveWCtl
F1MRCa/O0RZrFocTOmrlU7bw0oAKtafZUdXK/cw7WzohAZKE3PQV3OlOgTDhuRqj
V2kwentCId4gX1GgQw5dMDq75aj+Y9wxS0/YgQ1rS+b4KeyPdPtGyAGjGOHUsDl9
En+PxfJEu0I+8TOUn5HGcgn/5PqH3eqgErQaCbkxM89JAB/jS2Tmp21vzY+3E5RZ
z1zYh8lZNPXCWdzK8tzL1ido75pVZgZ/BSPmQuWT2J0xC5bX5zAUJedaXdK4zU3P
Y9OzF3MatJgVs2ghtHH2XQ5OXxjP5A+yJla9uODc8oUdRkdoXGVnKMlxysFjXWlZ
7qxzkjO+3Mvbiw1hnx5yp0vVqAs4OX1F6kdrlp5SQQyLwSStSlDkyB6NnPb9dKjF
KBety1qNJlGiB4ez4cdIatgtINYy74wbjsQ+WhtoTRUtiMS9HVxXQxQ8EIAXZH1V
7IUugFjoyBbg62Qw6rfC2PMpsRT7NJvMXfDp1C8/ubJHginzm7blyxWwTWW8/stm
RG9rEqljpncjC3zxNroNbMpQFJDUPjAkdfasL7ZSh2DI0179xEL4anofyUwTD3ga
tt2sv9C0OCHJSb/+sClwm7qXXL8cslYqTmE1VV0vW9WQOcaWIcSC1V3wk8eKm9lX
JGRJRYzlywX2jfyTKoj5cacAidPkJcJBi3KxmvZdvh93bt9VK2rdcHfLdEX+JPR8
pLRDSkaaRVvf6gTMxPelUBM6W4Dp6ebdJLWbxmtT0oZrQ3xkPbURP9e/g6mBuTq3
jggtsC1OR61Fy+bHuIMecHX4+DJ8y7EzvlFEWknmMj12V+H7mmqZdka/b+wTJhiA
9uAburlnrvMa1hSGNy9WnQlolaLTcZVnbPaVMNAOR5fmyRgdIDb4QiVx42Sls+jz
7zvrswKQify7AEuNzbD/kIJFtV5+X1WooKynjc94jMR4/tskeBchg4R+XFunnmAK
qY0pYza76d0pOqmqmXVQmMJ76YElzjCTzNTFpwVJpSf2rVt8AifN1KRhxZwBkw+4
D3Xx7AD/bDvrYYxQB5gHO2sYjgWx2BQOQBw+GXDOJqH+b0fc4klg/WVj+ba0rmHi
zBu9M7xNFo7yeKh1ntUUqXXhu64KC/jCeIOZ8lP2KSqei0LABzBZCYko2vDaLVTO
b50O9rcu7bBlqXzDCg58WUFYrEIdBTTr+qc7hdVzvix26cTWxVlo28YclVa6C8b3
FazQuu0tk6w06gBd8FLVM03G5NENZ7n+KCJmFXuPjfzhOiqLntl+nQ77s69gxw3U
R89UCD7s49wBKCHeLgzM5r2fmQerzZz4/3t7B16iCG2G3YTXCbM1+YLlAZ7BXUSs
q6mucyboKDNHmIQENk1oZWvzACT+j2rAdc8gGqNr5jWAnOHVbWkQ8XEYoa4WDAiw
lAhyE9130ZtaDMJAncki0uEPgU/1KEoWwLhwPhs6epyfl0Uk9wyZZSUBG6smYWrS
KiZrIek5eFF9XGFXskYHjBpVeT010OjGss8IPMi8cnrWjpxWlykkV9OP56y7InuT
jwHv/H4mMaKD4V2L18kXp+cSKG/+Foeyf27gdXk9uObviVJkLytrDQk3ICB++5jd
QnuuXj20iIvXq4CZpS1chBfml9G7qmFt6bP47W4Wcbr0+nMOdORM7VKe1utDAmJI
ctCuJMvCLjixPyxiRHlOzGy1yf3w/6kcYxpQiTxcfOIOy9wwXVjmKa9rxnkAfBYe
sH7PZVZ/4STIe+ruFS1PRL4ygnH6wJoIrMjvx1f1q2KDP85MAy/9kmOf1LRIaGVO
5lhpVFPi0Su+8YPFtIJUPCbOa9wRkSg3K+uAzk1qQ/c4ksZt4XY9yFWkF61PJ8kx
2mMBiKlVKRo+V1tkd+IsQjI8ECHUaYVxnMA7r614Ef8NqBxOkT/dh+YAI6ne3n2v
O9yZNXbNLY8BTkD5ydlPwX+osThg6ulMwVsUFuvSu5nG8v6JxBKVf9WDJGhlz2/T
w6EbRiRvc3MSyYUaUjV6wJff/h5ujRmG1EzSLHsHx/wQlG53LsYXZhYkihNNSa/8
bipYw7iIBRWQmyAvXbWmEhWqP7AA1WertG7dEr1iCisfKdQh5efs/MUj6JO6i2hP
EfLkuyVbaGAz1/ZoFJC+BRR0bGkP2K1z8KRmU/A7qO0Z7ki/vJxbYiPx6GHJztlL
3KskmtddBVIq33A2O2MW//QnA0D7xWjtSxMLRLi5zyOegNNI1Qm1g3A9XA5VPq0j
1IXcJk2pSDy5hpfS2EcAXx6N+HCTekeRQbHF1qmIml9D4vJMhFdPBJ6xB46cAnKi
57cItlgF8xK09RRE/p9FlYkjdwTKhr8RW5ZGiw0WrwBCD+cQG3/1SCLRK8jbLSIy
AomrGO2azycQqHi9yG8yl23WGA0im+nci/hJrjpiNEtbZHW8hq74pzziHco5Ifm3
KxNXUam8yEuQs+YuOh+1owcmK+N0odGZGNzR0yHZd19NjlGnxL3M/ficOITX5T7N
P9FuvPBVbi1BOApQw9Wdii1k/QJKvYGBAysvcyBKH9ylEw4x+heiryI0lncZZyJx
vqNgSevX0Ei6XBv93JihdSELS5SNDz0n9T64E/3C0MiIVDTJ7DvoH4v+lkCdhJMR
8LIYAPB0yN9RmqHIchBLwnQJs2GCurNxCPf6umQLOU+3Vpyfcs/7+elee4Zr7B6s
R/Rx3DZLRf1Yp8A+SoGPRCdn7dq9pYJY6tyV88Cz3I6KtKx2h/xJVjD9KCaESdy/
m94Sj1TDE39xecEp65BNFPUvhciF6DtHDUqorPnxTvxG86vlNtYCEoqqA+shME3z
6POhEq0XxoO88pM5APPyOEbtJRB2YEVCczYhqV+mJXT8NAltobyyWnS1WkzwjPG5
z/o8cW2AY5QBTE3hD4l40M0UDB0delge5AI5e9pSuCBrp6yAeEnHqPti97x8j29v
FGZTl4BoMjOxBjMf52iYfXoredYPSpCQIBwLj5UEutfQneDFYC7HrLCGe8FfMhWh
s0FKEAE9p5adecEyzR7IhVyXSRVSUjlzpnsGixLkGHnYbK/Ze8le95XFjbKe4s3A
rsX9L9EydkT3vyGJrzR0O+IW8uqY6ex7LQeLjzvbkERZhxhN7s5HX4KLHlnPNhiX
oZlbVWcBZ2Gy3mqCXcgIZ3QP0Dw5vhbuaouwVoMDx5z5fY52b3kY21XfpjPlTpYX
nUjuLJyA+Y+IFMT7UmlOmVw362xK0OTfHDCFeNHbb0r+XALSH4TgT9THbEP6lkrc
5bFcXBjU9njsmALa4yORFFBAdrB+Wkqe+9+PagpRPO2fKXrcF+7c7hWq1wUEXxbq
htAinhA+cMxMWXsfajLHXY8fWpGSppXsu/MrfIU4EraK3UT73Y9HbHvpSNNxRBUB
yAYrnp0aVAk032GkDAygzMocXyySiWGfXg59gZ7Tkoa67VTiwLSjpdiRp0kffLbO
FErXsmqiKD6/a6Hkyu+ITXc93SridxiA4+U4jW22Y7wRIUp7+teXO20bGVJNyoQO
nvOI2nxGabhrwjBbAFm2Uhf/tf8v3ZWummF71P9OgGNFkN0OnlqN7fBOtk2V268f
O814cf4geOxM6RJwT/2pwuHlVjKxCmVUAzRH26b5yB4q/1ivFBPoyfWuTCguKhlc
Vi5+SlrNap+5lSrHGPslt2pL7yXE3sxyGx341vbPv2n1mlTwz78LuI9QAFcMB1l7
A2qswcWOrYXbfb/fqGi8hVUknknx1Vr0rH9sm1ssv9NE4fxyaxrLD13aBxZRvBr8
ji2xT6qXS75DIa6XMa+YFsusMk4BrhE+fMIqDO0fRDNWjGHDikWgidBeN9o05JOq
ZDhIbSgmdKD28TWKZ25nq+YBsNhaAcxQIvp0B+9/Pl7PNX9rhAxyq2Hk/HM4eVmc
Z6zZGWHQN+tsyexAlIv2yTmSoO5tRIETFhzWB2kHHZuXN3X+2YaVshFcj00NA0fO
VeIJx5o//SX5pwsA9uJ5uUItqDymd5re2ZkRClBCIupfh8VdKm1cehHboNaxlfca
px4rqQUZj7wW1COqYDfBU+cg/L3fLTMHmXxolpqlD+Ah6daeEftcp0vfTeOO54b0
+WA9mKV/Wh7rx0mtL9LW5Fr6V6E9ynvPuuC+pCeNV2gma/vyDDV6trRRKt7Z63mi
lzI7VyZyC7yymqyvaOWLoZ59LdUlO4qXHOEIrx6SP3oL1Pvdmr2LvfGjw5F/Syso
LjiA1KTrHbFt4LbZKWRvKzg1lWz0Lh5UWIzZGtRoBdV4/RLxxkKh3+amS+T44UKB
ubM6y4YGJGQ+SgdHRQ1gapJFpO2TvWuk2nExGhQgFrwHkYtyLjf4pz+wSlFaMeTr
MYzT7WpLTWgEslnPY/+lb5uCFnh5jDbzG+9m2H7jma8ePpZY2IUWR87nOnA6G98s
7KapSRetNvX00LM9uihWg7l4WSSuLXDxYUik456Scv28vzhVWbqi8670zpCpq1po
JujePOCAkYizWA/AX5TH+iBUzcpRJufzbL3rLdUS4OPRL2ERsY3HFEniiBWvlMb5
TiAMYXAp2w3lkKlVfpXQn9jR/a6DfEbZUeXROcpGkD2NxCxckydeThE0M9ZnSqo+
3B36jo7UO8k1ExvvtxfV4ffgnj3+IhseR3r6jiu3WxploeVpJff8B82vOdgTYd3P
L/eTms7R11VpyYjLSQdcbEgynWG9B8btl9dyo7e9PyAmtu24qsAjQZAKIwDHAKAr
ffmPmbQYwUn1hLErndSnU+KweSKM4EbxYe7mP2LzItv9AVVQKA824/dV0MK1Lsah
i7siLJ7ObaIwVuknr3EMsERk4KSGBNRaljGk3A2VBf0PFxEmp7I1sH06HcA3IV/7
epEi0jW84HpL83S7CV2lxCh304r8SMsv241Wb+4Wyg8m3yNgU0HRdZJh8k2sHqkO
nTGNrSJEDH9Upp4HhfyfZdSPVOlB4XCPOM+oop9a5CMfCAEf2IOW7sTP5KLmDZKu
LpqnikMxvmETZlZ6BwCuQVXGbPjvFbwt28oRZmZWiqqwC8jxbZ+yozTGum0iDi3I
/ECBXWx+bL46s7jx2N2fVb4NbFWVMVH5mC8aqnTfwZWV9NwTM5zVL2dSzxcxtRbv
MDzt02lDpF/eon3cWnKs+vq15CCW+ZcJdPjr6hPmwpdd+6Xso/PYd6EsIzc4m7ol
V+U4BEy3N0gasRsp1DA7Nu7Q7+aU08Gl854FZAZ32YNC9BHpgtB7IwN9642mk2GY
fQvrNA9G3ollEIQ4CG/le3xBLWVOlihHyQ9HMyQMaq3mvfgGRaQ7N0ZggwJChzM9
jT949ECoKy/Jb5Q19tGBQwGcSBBhCjgeVPUKux6A8XxOEpsiSomHGGaiCwce7/Rn
PGy8jBrm8rcGUbSt9MliR3/jnUg01mBiNY0lh++wPaWtm5kodjF29VDd43q1jJs2
DGWoqqNgXMSE5qjTWUUsjtiroQh97dHnxqtRqI+mXA5XasZmxcVMJd8JwVbdAlY5
xa/tzc1TM9UeekNM6MhO9es8gm8M6SEgEKw7WLmX5aQQ2V8ZMMRw8RYFxio4x663
DJRxCN4TFHdmRzGIXYMqX8T6Pa/FoKb70EykeHNeexnHBNQI+nmyFBGoThV51haB
uQuyM14n1wRnrGqrhSj82mGtmT0S1Mu7Y0j2P99/QXuc7NkHCW1TUWjkWNplglFx
7Wwt5k7sUPV3tD++xn5TK7bwrE+vvjwvcWR+hAgczNkffgNDA8iXU/lXxD6rrKg4
thiKQyrftUmFjYo8YuOA+AG9pgjBNq02kHOLbN7t/+HvEHMZA01yd46/JtxQtFNh
RWADFcn2EA0Z0tIeu9A3rquzR/ylTHTWGJylV/ZCg26dGORhlVqVk/k5e9CDkHsr
/ktK2jDaxj1Cxz668sUVokkBdRv2XYsXvGpHV4gChWBnjnJcux2erttqadvXwnXa
Nhsez3g2m1ZU1GxBymFvL2+GHSo5K8IH/CZIuxacFA7JyoIao+TwLEZbmivEjwH8
m8Q96FGlthXfhwuweJkpfJ9dCqCLBi5Dj4GLsZgXNnzTCR6gl8VYFrPv7XbQGiVp
HH7/kTkW8e2cHgh3L4RblX0+vUCdsXuJp+u0aJ62M5Ne7oLzuCN/hOGooIL2qXgd
A3BCr28CYetgGLjJXjZ0YaAHYbLDLXA6obZwciBpFH2ran1EljiSPcBdGGJ7r6Tx
KSidiR8mgjpQbO6nMsBAe7eC1aPnWorXwKUvKuPYDpTeAKQJvXSZ5uM7Fdbrun29
6pUiMO78V1hRsjxtNvPU+OxH7AG8OLRXQNPQYkk+t5udjiR7RqxhazrgIXBk3KnG
SQMyGwCYHFfLkFL6CX2tjkg10T0HXJPUFCh1k4UUFw5iutSQ/eq4K0K0LhhMYozb
LtMAMsFEi2fJkbRYqTUAKl+muFsEKiPS7HIOtn0SRd9wmZujuwW2zglZmHXEEFcq
W5alw+DNb6w2TnrsbRhOxOolzGQldBeMSvbPVzOlgknBjdjxMapfh9GV/fGaX78I
f8Pw0U7RIif1tAitGWM5iVZ/REX6C+UZ1Y9TzU6gzpmVAsxiQjDVruFkMb+Nou1p
3XzVqx/wPtsESZ5jrA6hYS4ndW/I3JdGUCNtuyqCR3u08DnlkORKrmMp4CoVSRzz
cPrgKr2/WY73Zep9GVr9EHw1IQMahi4Mhcq6f7fkpfuaGsaD0Eh96n4g6mEo9k2/
fAa2vEs7FVo0Smh/qVl5zKPEKJO55NaHPxsu1vzQojgZNGnxxexS3c7XtZSt+6hD
VP5FuuTfN00h1dqi6IPbqzM80KMoa1uUFB3oiupvmz2wER8GyNMBPSxnrNJ/JBi3
vc8u32/byGDtV+bQUTvABXpVBWwJLZ3EpKFOg3Qkn51gyiVqhzlkS4sgowhzXXGS
oIyZ2cHuB7VYYPxmBOJz/HOPyK8rrJU/g7SQR+QUxGtcxv7mShgfaqUlv+4hQxvU
O1VY0FLoWDRpI9RkvFnvGDqC4eIbAPxISRqkX9KrG4nsclxq6azGx2xjpPIdaPt3
22c9qw/x1j3+FkFtfBE3OI6I27iALvkTpUTaPCIWyu5g7ttR6oCINKwBKkLOq7/T
cbOCjvwMyLPa4vSA2NEMzzZMnhF6NI63pYU5GDB6kluZvmi1Y5fCkIHjAxX/+Oyw
PC1QC/4gyEGTy2QbdKcyutEHvJR3S6dsXWlK6Jfrpjj8pkz0Ksx4MxspAAYDc9qQ
m33k91avno3WZMzuT4B7Yvw3VR4++7MC3TulADcnGEIoWDzTaBrcH7ZaiCoPafCb
GXDsqnDT6yM6kJA1UyNpP02d/DtLq+824KFSuTNlx0j3gCuWkpdHtAXhqfnfI0tB
YbT1s9LR1AqeWk8QdBvImenWVJmPzAU0Lh5bq8bKKoRHQdwBBKsXFcVKtrocjLOi
HWUQ8pyr6D4n91wqNiMabEOG7l/wKqCA+D20toHTCDF4nhBTD6vNmweE1YhJl98z
u2Y44c1CtaiXZB2IiK0Fjl+fw3kKipjKz3JZ6YVgEwL/I0ymb7faf2UKd5hJM4IG
8AnztNgIHtMOIBdUNRmMB0k8h2C4i+G1Hg4Eo5YL9Pqc7MzJfipf7VZybpgRBiln
pdcHbJ7WajgZdqmBXFqI1RyaAzi213fpEpeMssnUpRY8JYaEy/jqtW551AkI5fS8
MCjraiWa9ej3bzqpjFnRRPeWQWoYc9zHXTjlf23mZhz+2JOG+KyVYXFVB0eNSs/0
Bs+Ffdlwpb7GMLQSNIaekk5lU6f3lDuX3X498fwj5kYmX+N7zbDeAuDDY6taARv2
u67o4kkPJ8vejXzvtY1vQFgrEgomimuonamFkUFConndUFU/JU+cTo8TUbkNKzMo
/Aw8bg80gqr2AbRXr6UNPghxIMhAEiS3geMDqXyamKTW9pmR2u6KGnKWitAW1bwt
d4Q30D+YSo0zQWgqC2rwq5n8roAjC/hWrnaiVEDSQ05WHadCyxyk/3QeuI07Yrgb
sOXjAv9hsqg3QqtYCz3fekofDLhRin32ROmvPZu+AI6VefKldfh/k6zvDvKuzYNP
Q1iT3Aoa1wnW2mkP/9zZLXR9Lyx/F77BOfMzC7oFz/+UNuF46c1ZdPMAGkaVbvzS
+VIM5xozTDMqR/N/JwY3E7LKXOpaLF9NlxFdzCJh/dsjTtm95Xt5+8/gnoilAV9R
oIPcQMdkSIoyNSl/v3iC4Zfhr4UY7qCyRVqwnqm+oJQFUdPUjpTPWoFNz8H8PafU
z0h4vRfo4v8vYjJyENLXBeW/d2nlg4ISD6h/pPAVS209IqgvyVSUmUU6k0FddReN
766yY4yfB7UkQ6jyMiiOAs5xbhTZMrMX68rLFM10lakUPZRo0/UTon7lwYGHPdUX
AzHRqBNLDD5822xU165RbJmKu0kOlZd7aHxPD2aWIpGChgwwvkMetuL8+sFMt68b
Q0RWqV/Gzn8htk5fwyXe/NS66zwq8S0ElEe8petoKh4JCdtmcoBMr48BYr1Tqh9u
yLoc7kVB/1Z+PEmz0vcKS6DCHCxkp46wGEu+2dJfSiYGc6Ogge0C5KPsPkvYOj9L
RRXPOSjrDOopFRpM3pdEG+owTXKgBxc5bxfloH1nP/uxik2+SaJgVX/Z+X7alN/B
EJn7mN+7+knlU7vNj09JptyYwYcLMtRLmLWs/JDcYlSyLX+iL8WZDsSW74EzRObX
dH2YveRk4308Bt22bEWN4w/G7w8uwwaS6YN7It4o/Yvu8vnY4iqiYhsg+bsOrQ+k
qEAPAP+9ryJMqgqz+Iqb/Uc3uaUgLdsdJj0Jt7sUR/+MensxEQqCQ9jgwsoelDyJ
7cKeb45qMTzx5jhiwUBJysFa0Ucvpgi1fyz753EHnCKqDKT6FJsDl7zDNFiwfOle
ayuUmTGHmTdoc65gfFvKE/svQQV2JhF7qV1D58LkO+9KAjyTYMaULSbGT/zAjPNP
YBBE9u/UdIc+ImJEyFfXJ6Qt+j5fq/GIJEpUT8D4XwJn5Yrgnq+Im7C3goslVYnq
3d04g4Dgz3MjFEiL6fnMEpBOHJipE01zHkA0+iSY9kbLkOV3A4SenWQmdakUFZSZ
DOsJK8Bt704LhPL0fFNaSWOUnWLtgCbu32AzlMUJV4puz67t0bF/BAbQpHCPp2o5
NpSgOFs/LRm3X8ZI4FPrN19kgfSpHvAbFIE5X03MDG4/F9CokepBAdJlpF8Irlu4
5xFeL0dcgl0Kzx8whikTgswX+nB2dXmj8VKJWefZi/MnCdB3Ui9HuQW+Y44x9m7M
+3eGZCmJ2vVcTIhCilUL1JUSkEMcPyxYnCDW1ihNqfFLBpP9/cjXBW1B1oiqnVms
GD2VNJPoGVGV0NzU/Xu5LFhbPaRXUSyk1u5D3ykpKqa39/fpZejMXEqLCQbWP3R3
KtqVuXTE1hxc/CnmKQ0t6jzhwSLVx5xg0A8ZEG7OeMBDGZRCsiZpzImzxJ2GGIOH
Ag2evvDdgKxb5+9ZAR384UE+0A9bB3yMqMF/8WQbgBC7+MHYg7eu1U4AkuK8vdmg
ljBjugqcuzayg/Bu9eDm9mae98hJlGBvCEL3zxCHKIVh7NJyikd3VJKDuGF9WS4w
cAhFDsIY0jp0eHfzLjj5WhWHhtc/S/OIAS+PqNht9fL6FmureLezE4VBPjn5sHY3
KS+C3SYZU2N25mHVWTE/qcH/WAmJIQ4RHOJjoRLVdnS0l9hUy1UJusuZDRJ2+mGu
q1Hv9Dcrv7+9/ULOuBCT9OUkXVCAGXiOtaLlp18LmNdWmmRNmXvh22laGwUdJsQw
H3Zg7BwB47fPp2YyPJ4Oxk89BPSD42INcSM2qRFcklk4KPUrEt1UbJQPQ5/xTRYL
zLKrqX70UVYbHvppiLknY9NGjTHsUU7NqHziqJSeOnyjuZd8SUj3xk1130096abX
pw+x7mi9kSznloM3L60x0qBxY03Y6YhBMsHVJzgb5h+paxloqmsKqqzU83V/rjxJ
paxTr6oJCHosJCxorUqJ0xP00tQl/E1oNO+plvGovSTaJoRSGPzgfkjuR2kjfWyk
P4S38JGBw6eOkPImrP3+2s7CSRVhnB7GNCoDaxPMOvQmeD4odLPZaBFrie90szwJ
+PKGSYy58RGa+yA/KiUJtAyyzhXfwmb215KYxVxi7WWEK4fu6r1gjA7z1vOxKpdh
DEQNQCBMDCm3lRY/PppQAw7DYL3n8ChxyVcCW+52WoG+OZTQu6FFk4Ctbr6IzR98
rHgawjPFOAAu1AoPxnG6JTIdz/LioGyxA6Oz+PCOB7yGSOcNYdd04+ZzbLu13SII
dSHtf9reAqhg9rjqfKSRH6f3IEP1y/BECYxNnRCInr9/Y5g01Cmxs7slROcNIrqi
WlDRIFan5hJr5/VmN+jp6sH8CMG9NqWkRUF3SXsB1t2S/2SCwpyfM9+dpmmv4OIV
XXivF/iGbkoxe4RQD+sZg+98XjcRUzo3TZstkbvHx4g0Nuhuk+ZzJDz5H8YT6kkH
aWu8pNEAXfqknmF+32iAQEu4dHzBpyNNZRs7d2SWefd0i3Gyg4cIepMqmrF3EQLK
1c83c8RTHcMRiAi5JpVKV0p1QtwBxEQiF1VVV6dR822s3ZEcnZahHISVPK9xrlsz
hoSl/K0d4nh9//s8iLeVEVR88amcgzrDbm8hEPSsXoY70YBgjzmUgKC4IzAFH0iw
6Q23i0ivoaxFVryl95Xt5KLKqJvIFjxCUWYrtNAwvS4S72zJ4ZtEGczgXow53mDf
BkVdjQ5EIfdMjE8Fe9Y6nc5hgsdsvm/UXRac7nnMbyNifjKjLZuIsLyFvvL3QIuU
hB6xaBljmCrgaQAiQVcu+wjFRH1OZOy5BGreVky9tEK07UWoxfcTD+AGuzmV6Eon
ZT1yd8DXP4pR48H427bP5cHTEX3ZFw3kUYWCzw5K+xgathnTH4imepToAbg0UixT
m7DLNr4FpH7PJQaWVpUWQ05Y4FGu13hOO7bcIYCX7bj6x8OdD4umZ0mfyVRPeu7B
4KV87KOnoEzU1tIgjpzJJ4GYaEqaj+OpzYj4NCzC+txhY1pBONrKcRt+ASeqC9og
dKw567QxIfIiZ4lySxzP06Xdr7GncBsN6VlFfH23K8Wkx+whsfTSlOH8k7vt33zm
/iGAQBzbrhr0dvpuuLaSN5EDzr4whj2SjjJdv0EhmaYz17xabKFUdp+Mu/Ze1cO1
2xju39tLvTOTbiTsK+FhstJvdrUYuCB9ipB00CdQSyhead0Hssd1NvXyBQ7AILui
4IwLBAAGMZ7R8W2m2JZBL8k+5xQAQu9pmW9/mHfXDpqRLvgMjlW2WbqnCs2tiI3d
njWzXTkDIo5A3RL7zqGFBDD+P80e3S64XPdzzBZ7Rh4/1/uL9GyMe4qY0XoGLocF
WcZ61+iGXUxk4IQjkTJP4C4wXCZxhFh8IQh8m6hOoXQ96mVV6UxeuDhbBNFbTFeH
JYMnpYzftPjoPxH4T6y89eK42xkb9a9JO7gip4HBEN/X0cArYRUVSK0LlF1oAfEQ
CHfmE4nGvrC3UCN8qhkWsCx7An79n1QVLyqy9XUOYm/AvXN3tVDVnO3YilurgEvk
ZV1MwGOumU0CGDdZxiJJOhLLaezNbam/G0x0355rVjTvb5p2eDMWcMXoYl/wqTA6
pA0AKwRTmbNIWQtoWVJA6yF5YgIXMouanP/1jKdsgARRHJirpuYWjhblCYW+cdQl
GmsQ7U1FTjm26WrfMVqqOaz4zl1RolB0o7779gBnX7aTzBk3R+CrjtTkRyFYyTrL
y7Ak7qOpDYRUE3h/xuwPxZN3etMdYxPj7xLXVHohFl+luADPmxVnxT+M6N0YSsDA
KBoIFchW3et8hvYApZhvkzlsc0Nd6x60Y7ACEKEA/KkoORA9TVsypbtgILJaG0d3
EQoUqiJ8NLdae1Iv/JYWci9p5yhPIKjVUpWN1r+TXHyiUDHEAa8YOEw69crWnNr1
r0DK0kID7xMPhnTldz6rU+95ujhRnAv30KXwl4nynzhrDYf1qyhEXMTPeGsRZnXJ
IlFQXjRkMstjlmOwnC2W9UInCdMsGIpxSIEMygShrxEaZkFWG79ncvnGztRqIWew
Ra/rqaHnIPOj3tK45r56eBf7yfy0MJodWP0Jg1qJ0Ib26fqOO/DmMm7uyg0zseKB
bPtj1iCLS8/Zh23lBZBKKIpElXPFxSRHK4n5l//nRLfWrMLmTWfzDWFCUIoKIO2F
UYZ+25Qm0P6aNKut8kQfR147ZeW6S29lBsFze6kA5qCFRQZrzvfVAiaT2MWHgyR7
ShFVoVsDo0U9jxkrf5ns5u3zMG3ntycWDk1YqnlomcbJRrXkoOl0AWulNPJwnbOm
+njrHJV5NCQqiOn1qR66mFZcsoufq91UVsKw99lLB9csJm7WQyV1SHrX1UiyZeNf
Z18Wg0xt7DnijJuXXd8TQiebXfqgn4J9QCrPIuqNA/iasBSAjOVMmUXZ0IZQlraa
QB8QDZlH1Cbhk15feSMe0XeiFlq3nHSMGeCunL6H+/eOW2Cw/NWtdaHyOnfX3Bw8
wKWtZCbb26P3NYsXxSYna7DEUU/ohQ7ig3PupdN7xAVKB9zKDH+jxAeGVngG8pf+
jXQDaiKuoN74fPqjLYIIs09oQIBDJf7QOXlfYb4aKXiWP8E6mQM0BRGZp+xLTZKi
/LzKd4sfFheh0j1CHTYhHDa+VPAInI2Uy1iB7prOyLazQHy6lZEY1Wq/GW8JlVgZ
RVPGyOCzg6cbvn4S8EpuVnznWMATIOE4cW29ikWvdIEwl4AhROjzoNJBpS39IxWk
v0/BqXPfixU9h5kPort7kZAXfa+Jmehtv67pEbseSSlf0Ci+Tr2Wx1iO3QaK6+QD
TsWki8Ur3jfAyxnz0QplNXbmrP53nrsjyfV8detlUfORr4q5T1oGy1Tjq0PBkdH+
KvqT/cuma9UawPHEFWcBC54LdNUFi6WwIuK05a5KSimV0SHRbq5Nvpgecgwkhy0+
AgFnz4C0tcOVobJftuoiBqrn/y2Yn61p3LgWbD0AqH1IRVmxj5upR0HlXd8PA88a
/YY46TP0yISu4n8acPw7hmtVGz3lRSO+tqr15KXRrp/mrbGAA7xVjBHR2L6S/PBk
VjWgwlQVFcdyNXEszOcRpYqsxnPcOYN1303kzmLC02HhD8pWXWVeOBHi9BnBQkLt
Yvt1wnbbv6EZDvDBJKXAj6gRySopynA2yN3GqYJzCrCD/iYMx3/zJknliL2dJXVw
gu9lVtdtxhRG6Q3d4K+p8XWnQPSTYegYo5IfX7uSBwX1fuRjLm9aA64IHJO81Bys
UnT4HOh9x5damZetgQY1GSQGSjNarA2LwEPirJU8BubKbjWS3lBQbr6bCebuSQXv
P9s7d/nh4iBmillD2q2SkVXgM4WOEEbXe3NHkHQmiU+wgu90O9jTiooYynM/TQRa
pF14wc/QO09MWuPswDWq8YKEwHpejJ8InnuRWV832mgTAOVtlXvD6sdl7oEgJk4V
kHSChWPRWO+gbLHkqIYH8cwb8uCvk0NEVSfbnqGDw6B6p29ecCYnGdE6+RmntB11
h5zvpoRQab7C4Q5asfiqF0ALYxeKW+H+GIkItJAyGlulXSRBQZxUpPwhXLLtgSi1
l1JqE3fWAyiSeHBBsiiJqN1u+D9d8Z3doc41rYZi0tnCxgbAx2KU9cmFr053M2SE
FSetRC4dXVFaa3Urn5x5hMG+/JncX8JAkem4D5rlQ7JoECsuYQgwd2HtvnWoL7hK
QRE/BGYvKXUC8B36qA3BdOnt5o/gv3dyWsFQQHzvWy1XIVpdfrURFr8Eo3g7D8XO
myqGQw7lpw2I+c0IEbLEsKuYYPPixhPS+2qlpvPqF1lMbG5HdnjjCyZ5lRuEflax
e8Jqk4qZv8p6fZt7V5QumcddRrOX+VHDUfztAtYO48zEDimA4Gn0MD8UMNTaKWuL
I5aZtFHnKpHhFwYTuV6zC7nI9IZtn0/lBbrrx7xd5Uc/bQJgH2JCdhswViNW2zLm
j566UHtmsM4//oht3YzI7G7W17e0fuURnNmrPz6GpGAY0i/5JytxNKkw9roouFlX
GfSzErMEguDf7gCXjfPrJPH+CiDIcBZe68s/2T+wvelyh6hfuUjWmzBfbHW9HvHT
3i9xKvmUoMj2fZgqxDmWADq0p/Kiza55s1veJUfDe3b8a+cYzFoFt7SXM676t2U3
95xAQi5rSfuyZkPE+EPlwTNvVO7t2t2DIh9EPfM/is5N/vHt2ntaFnEPrpMkDNbf
/O7LsYXenfvwo33lMW5Sww2DqfHfc1OCcnYlLVFqu41/aXzGenDaRyPLrKtuc1sx
IbFM4uG7hi/630cHFq4iu4sNaRXxYurMnNudv4h/pQBP9ifGoaKvP7wHJws2TQCZ
/KGrfIC0cXxG9rykv90kW2gmJJRr+esCe74/2ynS5yiIkg7jlFRopgB/DXrCyF+D
0Cbg/1hei7oGT5vjNsNEayy9AVFR8BHlnps2NS7x7lqaAYSL4QvhwDSzbjto7XOa
HR05eAbucYy7l+4Fbt1uV5r33mp4q9Ptf2RFVGsOX3AlsNaObCdgs9iH4kc01e48
fudI6kNQGg4XyHfR1OBX1qn+kTnO0j4veYlnr6KOwR2Q5ECH6u8YBBy533ndL3IG
WbECghrdlc6fCW2xl1ct4vp0/UKuMRrh29tY430aEKn02jfQiaMogg8dvHtJV16X
J6+8T8zIDGUoGUC0k//AeIgdHw1wrJw0V5mKxqH5YW0EJ6cKcSm863Cq97mVQ6I2
6kzG8PRzm7PX9mLpsV8JqXs6EhSF45L0GZY69h9dLXmMYWRtq8ovuP8Q4n1v/lKz
zeY3sNb3AG8f3Z4r4o+wwzpLYZfNadjdWYmowULQ86di3euHZsaIDXnsUAivWpak
n2gHXxqx51AMeBQsyGxlfTfAxx/TpPmCD791sz8ERBPlUeriMaVCzeuyLixISzmC
8nhQz0oJlSXAmzKN7Y9nRY8lasGO7udPAOYOLn5SYQP3eYHiJklJxAUAMxFtq6kq
m3eAwQGeb6ZeYE3mWyQldvWJVfMnb3Ujob30VxdqTKbnRB4CVygK4Ma0O1UC1gS5
/TbUzT3GQ3uwsunyX+txufdILceWcdsrMWzF17HA88SegJizfzI7NVsWiYGI/qwf
qrcUJqZ762PHDLkU9cUx/Bk2DWZTfgOM3seIdhRcftlJkGvFNyunI4FJMZxvzPci
Qbod4QAzePya5H/DO72KfkjiUuk4OS8IqKifdh5UXiZFmDSrMtkS/mzc0v2gjCq9
NWQJORIPa93itZoaUIxSqHiQpYV8Agy/BMfgDSOHioiSRH4XPQdDR7evlbqqflM3
RoihbuCfKEqm8QNx1/7mkMn/lEhXV/8mHzYafHmGPwCEyIBk/bgNiWhG3+/egJHS
4sm0pxe5guwqvuaKVuBANXWdN1ZMDJtFY9xyOqK8ifwhadfbvmriFtrgNHj9QF1Q
Tc9Ykf538OlRHCNaDU1ym1YD50UA1Xt3UeIKN+3l4qLSM4480PPi+ein0sSeixB5
B2U4MFpUzsdlLhHvu2QYCm7KtzWgeiDNiWoSp/caNz1ZDWHLV/5f83Rahb+h1+O5
8Z5p4+APZgQfTuKg8Rhz+kjMSik02b7WhtjNCo8FVY0DHnop6YLciTnjEyHv7oyR
x3Xz1OmOJr9N0Ot4j3Znc3GeNdlK+mGbwmJkz9SxXB9E4fhMvL72ypTvljBvwG1f
DgVQ5rs5r8OoMZTx0+c788zVdWIcXFSHUJRiA4DUYcA6O8n4zGf95nYqxK83MlHL
92C2sEdmhslBQrqX3+3P189j7kxbjZQbtuhaYnBiInbWd8WIhqN15gZEh7AK8kUB
dcDejsLv3peM20fAOvtA7tPHU8Dlq7WnwFqRg+EIR2CiUnbS6+m91Cz5OECsz1jt
ITW1M9PCzEBOi/fOPB/GOnqYIl3SQXITRP5UkWUqPiptBJYcpcOqosBuhUt7dL88
SJWGL7gygmLaLnMKUQz+Xq6AtJ26O2zAWPU24GKoaPSvhG9SSmEfFWO18NGKyERa
VwaFBTZqKMN5kB+gFocK4W5NOXCYbCE3hbXt7pND4xTl/Bq+es3Q+836V8+Jqmf4
TVr7WaTqU9leqirYgtpDfpas/V6VHSiRiUXdmRxCRWpXkGkYPr/xF+1PILrtZTHH
RBnOfcWJkdM9YwTqOZDlCtZS+F9mb9B50y+WJpaPMKoMJ4DUMUEFWicCCePgvEg2
q+X+HU+Jgn2BUku5/dIdeLq+mOUuxlh2H+Rki95ElEz8OUOk6OPSnmWNXj8l8IYu
w0qyIEJegb0eHIDE7kEZXNx5xLar/BXyekP5HKI7lxAUwi3f/xyenk2sVO0+1nwV
1Q4zAsLO0GlC8tJjZN4lyeUxGE04qW3HgVRSLZ/LNwwUQ3nqdGtXWl8P0Z9RCDax
7WWNbXq8rHgecoyfEzYnXaPwGwx4LDpRBp2O02zbL/+HD7n7dP1CTb8M2MgJs0Is
4AZ9G3ISYjq/xWGMjmU0YpRFJxpCITsLuL8Oi+XDv7llAu8nOwRDCZude6JQ4Yt5
Jv5XhNA9VoW3t8FN9aJgrE1kSCcgxRRAUVLx7/vXKLUQQ1iER92TrIw8LBnndPl3
l69xRZjdece4Wqha4fGth07lJhGitQg8x0tBYFO3OoCHX1BBonz6reOgYv2bm+xb
4Uj4vg4O2L796CdM7yyOj1BS8haoAsrqeIBeBLDeMOolP18BsJ6Sktgm/DuNBiZH
ov9X3b5cbaOY868ZDEtYhh7iJUEyIhosrzw+blq1GEex2hSEMRyvvw2ShIDRsyN/
tp0DYcft1zNfc0Mzqq2T0vykjUdPcErVqqB8JYlEeWsmuSLJhEOywqC3X9gfDg45
gmnJ2qk47w1RqC155RtT1pGhc++SvU2ota9HHUUGg4GPbX5Y4C+ODxtXuzheq/y6
oGnT8duvVQW7q1qPY9BYxX3iDtImOdANDcvYh1xFzO+pmkMU4YVvBHJBDqeieV0S
Mxvd0nLbStAuZx5OrLjutiZLvC19LhPU2BbvFBbxISZzwawhd5EusjI//+qZA4K/
cYeUzWOCpJSPzWKDrjzt39hoxzl5GIxeZxim7G8LkXY+eVPX0J8tYwpt4GfZzoRu
mX3d/KrZWZ/OCBv/NYWrtl8mi6Qm4v5+5nXCmviWsnRhPKa1+/zpnVzht8tjik0s
7bt/41CS/frEhANjWx9ZSk9/gf6iCjwgOCa6JihfHiaAxY6WWhDx0R/kOHdxFpcI
PMdApuYY9YkzjaqxBpZIxPFrpCRwtFynsoE2MLRJtWVSAej3wFxD9aVovtNg9bpy
qOFS/BiOzS2YtO4dgtEdqTSfT4gSBppFgVE1kX1362PdjB+Sgf0bI6hPgGnOrei7
nKgm+5NG8txU5fp/1dQKAgylSM46/H7INQT3+lPyW7kdYD0WJbXDY2o3MM1iuffF
HeYmusKH/KEd19Hqvz+e7l3AElBtM1H7xuoVWGRfSvqYPEpiVCztiB2U8bqm7PVx
Fqdb406LgYpM04gmOEkC4M/l4ywFCG8phYLAA0MoDBSeBhS5mvSUZVavz361CWnM
3mxwQUVgApD/d3Y2fsb/86kEl6goqFMmLXxzTqsCwWExKef9fU7Pa0VaSKIMVDqW
Qcw6g1cucf0g6A3vt6PLbPDaEy9Wc3Jl0Dr6IZbVBISHNef+sd7JIDDmdw5jiP7h
QZd5bP4Pv1+DL9+sUfSEJ6+L1WLjZ4+2SY+KakxuyKdl+7G+8YMhwiiFx0IwvqoT
q9oN9MQgTY4wIP/rM+Gg4Ycmxkt7TjNDRsYgDQr/CZ7cCof5OIN38ZGYBaMczKJe
Z6yot3VJ8xnbZkc9vEz/QByc2O8O5c+HRRXASVlQ9+BtV5rbBBFLyzCisKiR7N75
7yC7I1ntNcaF+oH5s/xphu6Hc+zQdA/QkOBfsF98Zv8sBC+A8uNBH197YA4Clgi3
2AD88iRunEmWC6Voe04K65dif+uSnFaSLKDqoZ/4naRR4qguZtCawuNmYUos8e8x
nCAswxe0g59cklO5kP5LlkT5+Ta4SjEwboESfkNgiGl1pFHnrw7uj/6HXz8V2b2o
pPq38yxaMSXykcBqFLYnup0lgNrMPcIuZPNLAgh67/Os/+t8bxFDiH0m6ZzZ61R/
45w/Un9k4F4SZ4C/bRSLqBWiQKlMdTOB7bXfSAE6JejaWup0TDaGK3EycFvqsOnM
PPQgdxpn4rDfxsPNsgN68n1DbyqGZScuu3qPd2HwcGxS5IbXFDUdTcbAkWiCXK40
H54kEUfZdOc0Sw7F8eLcScTSPaqzy3OxcS31PjWJjO+jtGO+kECBVPxiQwLia8Pd
SOkSsldOYsBeUSqJDCaE7zWg0CxFxVTVV3/NAWL2mQV2SW/QQaE04DlrFzPDkKP4
zGh6WYlRrocQJ4JEcmEYOeRU/53By/hshTF4VvGN9PwED8wrQY/Sg3HmqLm/YvTk
zR8OqzHec5Og8UB37jO8oW83EGzC1NOINSQx7wpfa9HgO0um2Ama8j05MNRqw5H1
6CTafUjDX7VBLkhsyoQ80+nXWlehDf/JBTcrlu8g4InjgaOg2g2WulJhuW0nmxc0
YBNAB//cF3FGca6o3IQh1C9Kai5GO32ql5tIZTzLEzU04VelM4sAmCfQI08Y8WJL
2plKKQPmHxmRsIooYiWCDcwDesJI4FojYSY9kdIIV8PDVTh9tN3qzmUQkKC1mTc5
wdBB8Vk9WuskPvvZgIFjX0LXoEzS7LBw5O/9sSX6jKhOFx35eOv3U3zICoccNOP1
y3AYFZQZ/p8NJtTmRNTkf0Stt5uMFhTqCGIlLWAGMCSxH3ywQDK0BukjUMKgpggt
irBA6pDjBHhRFf1l8Sv0ypn1W+bXDqR91TvHk8klfI0b47zl5Jyprtq6Tpm3AHr8
ugdLZP5eMH1IIHMFjRq+3ZjXwePipMbOZjeIzpkWZgBl4YpZ+zrlG4+d/kui0fgF
sR0xYlu6Q6u1koY4eeuZea/7aO2jFJrmplCZS8/bL/E0631D9nkfQnvTr5j0LQtT
+1QVv7xme/yQWiNoCfKlDnWsuunI6IhuHit4IInwIs+B1sOs0s4qVn0FbQSBn9vY
wu8xO7kwVUn9s2SSsIcM7bnE+O8BUy7dDeyr7P9IkQWqqp3Jmqqby8S2xsSE2sU0
uRPRM7cq0tLrsXS3ZZvOSuE20AAA/Z31EBucjEiCgDhYj9XHAb2tnloUzmygTQNC
VNIh6/C701P56HLVBIWKz1l+vvEcqJo4LZCJ2ix89ifvl8dsxouktv5vm3v+mwzT
OHa+9Q4tVla+gTkximgao5/UYCJ7YTVh0wRQsQxAZcpGY163zZ62qPQgg5yMkgWD
9zYw3YFHVwxVJLNcdnZqdOCcMa0vzf4FUj+ThiB2aVwdMKIobgyd2jOTbKTT3Lap
ciLnSFmpFC3mxmwigSQl7dFd9gnQ2NmZFUez8PdBlMeFucprE9hqObcrkNeQ4xpz
j8csD8T2WhQGfdzk04IHBFTeXoBMRLzn9dsgwFk+pLWlU4+rwtaeBSWNvjxYXb+l
OcXzsIOQ9u37Cp6i7LenwXw5CBoQzfkUitkiq2dZGiLV+MvC/+0tOwi/7CU0aq52
sK9HSD9I5Y5yJSn7RsU9jEJW3gJVCDsxqnPDvIzqU4TwR1wbhNp4o3LLuU7pBB6N
1EjRuiclw3ouJSb7Nm7LVUCIm5sBbRKt5uCkwdXZkfQFXJLHKPC0gf5EhAJqqwBn
2vqeSVLw3p+lmCmHbac/P9fc8DzHoRzmxoENvAbG8FnKCtlSlMBrGkM3e0nkvRW6
5Q0sJ6Zcs1p2nttg3tpCy/qdxyrIfJus//t8h3VunJI7iWzkcUkeGUhhuD5WejlZ
61gv6etraxYH24F/5MlSQDrTy1Lqhv1Y4Uh7JcFp2p8VN/TtnIN49M48K+ms4cgN
LGGy+8Sz3hLgbGgXbuXDTBZ8MwhvLamMgQtueOL/layMKWHOrru5hp3H+Jiud0RC
lvCnm2u1uOK9EchZyOtbGe9m1MO9gUxLLhvxsLTQawGkAq95gn7BC3FJkPwwR7zZ
ygF87/aRA0YU2Nh6X/YFzvLFwPSzZ51dbIqtPQJtIyvn2aTKIv7KSbiTTLEUqhPy
e92QvIW/mlgGWbUbNf5Lp4jrngwqJypMVp5jvAQ9vi5u0RCLy2swcAhlwJpVRJHH
R+/2zKS0fcSKygxxNNR7sTzoZkBI79KunL/XjgZUeLIl3b6LhIWJokUDQr8CHK/e
R5+2XKTR64BYMuVObSYlrqgW2gUfB9yElLSiLGC0n86fYO9R1Jsn86BbTzL54s3g
EbPycqItsbaxctIvRlfNtPDu7bSfIrhADd1+fayEHq+bj7jUKVeIlIxWIs1C1Vru
FrqjHSospjQI8LLFZAvThUrGEj8S9DM1UHfdiUX0dJgRv6ANn77nXGDWU/79j/1q
t8pGJGSmgKYhbCaEJjPVoOkGLO/0ign1MAQXkn3bhVTH4qSiSUsbGgucuGcfPVcy
Y6DZXjsC78empYWL6eF1oGf+Qop/GjabxuJBNTJpzSrt/DW1QwkIbcjW/6vh59NS
x3PYRngUxveNTFg3eAmd8b5vg4uaIp0Q5xT31N5wXw2+MuJQqZcht829sMIN1n8j
Dga78Fn531yW5WzEIpXHH9GA79l1FY9Y4LynyupdA+aDoRw/xtvbwm730zPYs9W4
8XlJ+/Ano1aCg/u/C2OhRRjsXWiLeofQczsarnU+Pi+61gwoVbyZh6Ayr/Kd4HwZ
uGONlAK1Zmt8PhUxL52J3TdWr8F3LiX5fJTwpLOd4vIyymrui7Jci9gFipnOc8v8
IjCvwYXI6kMLs97OEeHsGvwifZwx1ztbnWHFzrLMMA56hg6Cz6XzcFEXH6YS9lTs
CM0AD+EVpcIGx80tG89xqnu3IS1mP9MOr0H0RDJsd4bqfiDYUmjuNEZ52S40H6z3
by2z4+aT+j8jhDBdONvbDGcHhki3smY5Fn0tgSVylPIEiKJzsD18njKPckcp4lok
u3MFyBbkQ2XzXtwOSw/uGHKDGhDK2b+ntHcsZzmrtrSYcoDMMQ5S+fkc5qQBF40t
4dQButPC8+dKfU9X25bJDD0tnr5xZvx9YKgM6nSlPjY2lOOGFe0NSJPbLFtyoqY6
+fg0TW+Z4jR5rEJCJ85IAR+JT5VsguYcJS2KldH6LkIy8b+Bc9aeNrfUqfUsNmBr
7QFPyJWC2WW02asE/Fc9fk9PxWkwnXvvQrD2T0qDCw2o25nDm3JNu/FFynla5QYi
tfLKLzQazy9tG5Df3JG7SBnOFiE27wfSaWyXcV0nsLFsNGESl2Veyeg3ErMtoVOe
Bc4WGtU0i5jKNg6HrnF5cJjpPAbLa26Y67YFG8yWCQH+w7WDQ/6ix2sjYhlT+3CY
JhJAgqv/EwbDs2l+yiYrVHHfKfE2+fjYVnjQ1/etUUw0FMaXymVxr+JjO9cAHbaT
Pcsuf3gqGOVf5hqFfgEyYV13hKclXGlmIiTr2nDSsrNfPWapL3eN8MESC1kyYpHn
wDkb85fY3oey9ioAjA5XlbORb/Pm+4FE4dF9ew5OwpGPMOGCVZqG5pB8uShGsMUz
BrG9Udqb+aMg/IedyEkxaXDEjnXrr8HPv5yJox9+CD3OBFIZFSWp+5TxL40oIOGH
PDHIfRQQG41QorjH2SFpOcFzCGHdeFgxJpvmNfC/HLmOm1GwhtDsR5X1ZXYE1XQQ
cyQBNQpCn+K320HO9w6bWW6XlxtbQhIY8BoRbKJEHn/hS1cnpuow9zdr2SL0Ymiw
4LodssK6r/Se781lqQWIg4lOErBybCE1i9hiOnAOmZPZesum3O2BHeNHehtO9Q6a
hMKOkijPUK2Ay0f0ygcFC5wrG9TtNjfmgW4G0wX+33rfnwgyVmUiLWhmO1eHc8eC
r28zutedSSyRvdigdUmJmXhmZO/LtHZ/wylHBEV8Rh47nkw7PAL0Fb8Rse9yi8ng
o7qo/ZPIIIAC48l25JQXF6kesQXHLuI/uhhlxtUdp7LrFYqOXSzNPdaqGI26h1qA
CadkNYveyYSfPh4KdA3HEk6tCi68rObQwMDPlGMlWogVAlIntOKSIgu+zOC6bP99
CE9kKTFtJPirTdUNbsy00Y06fT2oU9RKHfI3eBN5/g9GzsMmMWYI49fnjQNUuC7W
/DFTobL9T8OfbhUqOAv2tfDhntL1V3PS4+Xzs+KAFP98ouP5yhlsxpaJAoToh8rw
WGpCqHQWUnBzCkIPzYuVfiC0iV3Dlp9/Wve4pZ7UImGMrBJDjl6r+jjfBqCUJKZZ
+JXkvn/caEYFAXHvhbJsuEKiHD9ah4PJREfrS5NvMZkPig7DEX7CqYCfhuPs6asq
C5y+xUz8+PONoST3X+k/8HgNIgusq/vtoMLTY4Y7oqQkz/PNb2fXCIFiRdXnUwR7
XqQtzrUlq6g6Hh02/8YmnOOeUWXRGYPGi/8ySEasp8raMSionn9ztTVd16IlGuVZ
27+uo/zCYdI1jAgA6au2dZLC2lTX4W4VcwwxjaAYGnF92Q0T8Xr/CBEIY3WsPLlh
qd/LJcYrdlPlkcKsoQ782E6C+j80uAMbfv60QZ/c7wsAiDixLSbQOaQYP2a+kAXS
F6AFp+KlQjpmxWV8QxgBYR5s0akzqGVB/wBcJ9Ew30IdMQXapqAr0G813/eCP5xv
IGdrKq0H5WrWmooL6wEAiaOd9mhMSw8znh5zwZmyfDoKRMDrqbw/QgJF4IHcR277
39b7pgirHHtGNwWc342OAH+nXczt3GIR1UPJ5F1nSEDau/d0iHm5O83tQOUKgxoR
N6sfavomgM7dmTC/ScKm2g+0YLAq/rw4wgoCxyojA8PHvxzESc+rY4dkEQcpaMCn
S6sVLjOMS6uNrciF9kiz9diZ6t1v1FQoo/aujh/n4cfNSTf+AIKTnm95KuRcePVB
PCLtW4ROFKzUoRB+dfrhaIjcBEhkB3w0QFmnvdXp+9pQ3qTLuzZjw3b/2v8Ezbni
FfYvxc8psmUCb4E/22ln8iXXDBkzIyn3+d5AkL4amIEL0A7jj/KMhopAxnjqnl3u
Y7gC+ExP4uflqz9Zdmy1o8p5y8FPl5sWhXxQ+bP55MjORq/kHpNgIGWT6cCpK2NE
OIFG8Hhpv4CEwVvcvtAq1UEO1+aVMtMvlBYgpQjHt421xHSpdJhrvPPSICMeUg5b
FFMg715W4l7GpCp265eenOQZgXqobnIFgRcXMa6NdIY0d6u6+hkHn0I7Ty53s7/a
Hz5/eoG5Juaa5w+2BKpgkM9en0e+jX4uPp27R7a1M1YHQfwReR5KE2Bt7CBfj8WB
9zSgGaT0BQIS8mNsBtdO+1f0OdPjf/vjyDt+jW8pU5LcreJZDa8mHZAm6fsgCFt+
XAOHZ/EXW775Ut2GQO83XYx6o+6BGt9tTNKG0UrO195drYrgJp993LvOiN3sXgZa
J66RTNLwRXib/RC2Bi61vtmB4f0m273u3TpndaGo7xtQ6ibFu+cHzkBAWQuKuH88
Kg3D4HilyoMl71HSD+LjyKjAP3MMMhf/qyA3svt6HLtWlYXT9ZI85/Aw3xX09Lvp
Ftvxi39IVLnSmPyg/py3mcnevamKM95wcU9rJIGuWFETaoVakolyy8ci1D5vGdxy
AzMTtUN3sNsQRdzBvMt5441nkelFv9I7LHJAYuBIUFqBAmaT32wCxctOqIh8uH79
nQ8LrY6GCxDHvfRy/a+1ezHOT5x395CxTFdZ6zdwiMxRr/c2Gqn6D9Bjzf2ku3Aq
rUUTq5tLOtn0U9afJAw/EXiwoI2HRBmXFoXTDRX3fb3mjGz5QDJEKlHvpnRv8why
n5FG0HLCUxqE92Wzp4FiaiqeLMkqzilUQlWmuktrwIlM+iwLZnHzn21yDyCgue8F
kw7VwMpREBXG1dZBkp3z0Tnm4KxLKakrB23TrhmZisBznEzdBapwgSPVy7C5sw0d
MrughQHFc4Bbs4HjaJ6uA3FtrgtBgIiM7daDpVF3aG5TC+4qKZgJTmzTBMiA8GWH
jSsn5LLNPac3MQ4NNQTVYHQtWU0kQL9bFdu8TQ1SltGFvEvF91tT0eKra5B54L1m
dJdE4HUJAytnxcqf09qrjVC3TWWMURgRnwosV4UGYmrLieXiiXu4D6o4NRDUeL00
oGo6qSP+Wc0HTfn+7kuQh85ptCwVqF2PIjqccTPAt8dBtE9877tH6daecZ8raqjQ
N2sWCCgCXxBsk8PlYmbT/dnXf1P8B5lQLv2PwTNihGLAc+yEgR3ESBpANgC50kvd
qg8GGMyIrAi8n3drgVdPlHB59gjwJ0+NGX75FHZYarb9J3wjQsztd2YKshVuVuA1
9TpN6dgxuuT5wv+h+g7JXV+xHNw3opOQZc4cpM79i0//0yMn+++6O9bu7MjMmhY9
PchjO4lWZ/0b27bWsK5W3iUL4JE19QEe+Utq3uiKMNh/zPt7n/up9A6b2hLiBEZe
ob5xOOqPSdrZgpPlkSRQsc5l/VaSKBSB8VJQ9msvlDRMCWLNwL5dNzKaesNQ3bvm
TaLSj1D0nh41TIuHf0NaCyHuMdNoJD7v3lu/lOgdOdADj1fj/2l6MbS5xcWJXBwU
u+CgZINpYYdFE7PJ65Ruu9kcO7lnxh7byOLZPDEeFH2GMZ38poa39tJOF3LOZr2z
qDQ8V8OJ1k8Y38lSgevGlfO4TvQbCLqIh9T0YqkYT9P9xKnxZbNm9JnBZ0aGWuAn
1jM2MpCCATKQnl+2T6IJ1ev5488JThvax6mKlGlIn+WJlUHUbB/dRKsVaIYo4Um0
bFWre/LN3ecshRU3eHL6asbsbPP1OOQo8k7F8oOI0sQdx9VS7LLr9ltr4YBcfvvJ
LXadHL+uAc626uG0tKfE1xD5ln4wK3DsiksMzYYTab3VtUlwaufaMSkXG6l47mHk
2BPSzhMfZr+mEqjQNF/sMg8SpzhGSH7itfdhotKCler9wU6d3tC/cE4T6G0Vp1WI
pjqrXLlNO0VLUs0tcKttttME28bRESPPan35iehqap+lhgnqY6aAA+DM5gA1Vg1x
9BDVBCsCf4czkYJoEpA4VCdrz0mDDo3z/Eo6YBcQ/Tt8stZvPlapCkIzTe9Gfxju
lCaM1HjSSE0xIRAk+Mrm3I2Ukb+79oBa84lqdWvFc/LXXswuq2C/3u4XCV6wGDFS
zHbypgbxU3g7US5ePwU+9aes+c+J2GQKQNboQ71dDloWRDIFCkYAvGae5iSQUxXO
S7qDuoeivDqFUFnUdSQUMr4OKDc7GBQ5D/wt2TX9FXs30BJ2jjMzsA5mxcf0XbWz
oTGtN02XataiTFdttlVi1iJ9WZKpck32P3BNzb3gk30f9VvqNS6LKVkM9KqHy73V
eTg2MN75LRqOhr7jQiigU4rmVMoxD3B+ktbdY85Bd/nNsm5Eae0eV5BY2CiyvAjV
Sl+6pS42G7Rr7FUsgxrCC3OufC5Y3I2uhKU28Td9tpp66XNXIzeKK81BwXMwmpqc
qsp+6hDQpX8o3MTdR311ZBBeyHtshq94thbe7ETZ2kQFz6ifVhpg/g3aVJRQm7zB
pIgbkieVBgFtosOdRheF55SQdPcuKc292lT3m6JP0YOAILQPdXT6CBcU5M4Dceez
1SfYTvz/2VKdYnjLh/224sKPMLCH5j0AUNSYoycMhOjA3IHTh2OQYirMTK+UpaAj
uY1d4bpJPv+Bms7FXpFWeOwWZLz1rl/P2eBmy3iOS/Kuth7TO7Ct4Z3NNj7hat4E
pcVCDuSe9RTxSiUVvSv0bSINHgsnNi7KaE/FyptY6nfwrIrStssSYtrc63GKnfYO
yO/Rd38B7sv+S4p1bdjnjKJT36Y02XgK44h9/kx55nlVAmLZzEKe6hCvGXJo/w3f
jgn+8IQAb9UFaozVu8n+0xy6OixNevI2uRlPRSOoF0FVOi4J2Rwmc5b/nO0Gnqte
FDBZAntyBVt29vy26nKczZQ2EeWat2i8HYtxYBcdELZRjdRVMsBKgM45Mm3EmY9e
55EZU9jqiWoh+qe1DxWzLYW6EsoseNoweG4NYVnA3oKZS8L4giYkCjse8gi6QoqZ
+mqmUqbUnZXk5+Twx8Tk/uB0IELfY8v2bI2N4X7njxuwRKIs4BcZD1z/dwdpC18j
9L84UqXONmV2dMijNraYx866BXcuQZVRKl+ngxJ/rNLBCEAl4M5O5nZohHZgvgr4
3Y7EyS/QkRIBsi8eQCLaoXAOxBNN5f4mqbyGARwYS6NiUpmliaeMUAYM00CVvbnx
Z3bFNTXGcwOoLjRb93rRHSlVhx74ovyHVmxwMmShQybejebR0lfHyQQ3o51CZ7y7
/wblv4xyL6fAXd0m3fGD4wzu++Sope26DESAZCcafd838Fatw04TdTUFtpZwPwki
8NEzCIk2nSKWigwvNi+Tr5vI2CH0mCpKnnhG/qRdADeMrb4vC2hyTEd8gLdiGVWh
1i2GLk+YRANizxLbzOHXYQyUjHTUZsb9jppXm2FaWrx4V97KCHx0AoBQBph8C9iA
NzfzRsTAs9oeSBQn2B8t8a+KCJBvvyGty3gnPmujvv19GzJE+8NVJsTo3gscJbqd
wZ1F/ywwwRHOEmcxe+9DOHsam+USk7IPyi8xmMn+udPAUhycfND7CtsF6jMcPCZN
5/owoAqafti/539qZ/WpRteqLHNXT6BwTVG0kQoJqBPUUtgEgq1QRRorm7+AaKlO
BEC5MBuc34KYz02I4T/csoinPI2Za4/gIYqPmIp+yxioh9e5l/zJH9rVKnnWRiSS
EWC1NZ4AJHqNeB1VKtmZnm2DMv3lJctLojD8U1W8NXO1NijLLbgtCUMy7I6KV7Zk
BxrV9i73P9HhwXp7Xz1NQRqZgZATUD2lts1R683pP2MaSNUdWmXp5tLN0mcKoHpL
Bl8poCqCTC77T9bVhHGOH/iV/yguHVD5AedIyHE874HjPUQfJSPGJall4RJe/a5k
z3yWEIAEhrhdV1wEmy3IyK6BGid+B2cVLvXwm+BFDVlJoZvGUc5X7wIOuFJKhuEb
1ptXDL1UMPnf+nS5yanPUz5TK4Ok6uOcvvrwf/LeWhZ9sloGl8Gitt65cDAugibC
jpRDXIpnAncSHYSTGG1f9Go+z3zWnt9z3QfTQp0qaTiivLWASctvPFBiP5PXibP5
CF6IpIO7TpAFXmItrbDfUcHyqudTik3QuPqcbSC2SQyhX7yKn/2rxCPfWrDTyPyN
LsQu5fBNg/i4g0suheie/WKEhUWP3Ym7F74kw2elNwfaQPHCgZIRaXIpw2hpSTOz
zf/OnTUb96/XVp2LMuPe2LuRXi1UkBzY1Fl2o62uAw6UDWwmACQfUarTmMoVxZcX
qV5sxjFnzOkX99meG0Kykth8+vURs2UxLkmKm0/MUWN1FaN47p/q3JKn9CmaL5vj
0IXpSncqDV/lQ9k6zohuujmNRz0Ps5DH+ph7jT5pc9sFedTuNJqvRhEAA1TTVF0n
KIT9mJR/vPlb5oLhlASqlyhg0k2Ph9Cij2+pTgdlissq74sR74wWMnV9UHK5cxEi
m3xmw/ayO4+iZwYH96v0qlU3L9QZd7RWZRhQPjBxmm+unSsYTh6b4wA5RBlXORWV
/cSd6agZcdpNQmgeqf4RS/+mKNL0GsS+s32aXGUzL46IeQR5aOm776lx4sLBRe1T
I3rp72h/354UImp7h6QrkMsqyxiD2G8e8iELMSc/3umPB6BWBYaFL3KUJXBPMLlZ
qLR3L15m9XWo0efsBuG908sJKoTKcna9tcLX1f28viAtApAeJ78obcJTw19Wh6kW
+OCocfTCSAuLQZuiu+w/3DNVLZZOVmfaj3GkUwruU18IOpcTs+X85YZQASPGRgsr
4Sps+xxto24yPCJXRvXtoTpl2jBLN273Yc5yqHAT6O+aDVgpVBWtgrRBUbE3A1a5
Lr86BkHyrEIi72PNCQpIFQ+LeWzGnqoBeasL3Xvhw6oF78ZcSy2s78uiEq6opslx
hDXIBZxBCmnotGhTozzMGgGOeJgP39WKnxRKMKoDvXy1CsOByrceQ37dWj31DEnD
0P29+djBAkur4haHeNpbWBIqpnnQmsEelndLKdTZFBCtyWyZUvxu2dgX1BV5dyYc
mb288LXevfagCM3MSgp6hwvKYjG6Tsb4teJLf1avT7yhmWeBdM4LPvkvLLtPUjGa
7jTW+V4dZkzhsNDW4HcsWmIDq2Iwqwi0WOPfKf7xOPoM9CYKVNbxDGvlknPBpc5N
7RdwHG2NeFBk0Q2ptkYPWvVPfhjBEaZqHumavfiOt9zKERlxfTD/G34X6OuzOI/+
FA9wojfEVz30eQt2bPn6dRSZPk2BywsUHpRftq8LllzeKV1qOye33Fgy0Z+4Uuiy
6PCWzrRKfJ+fhc/EpOmaL90QPYern2VX4uU1PcgVvDBFi7tJcLmLVfQorWEkTf20
1zxhbCo07aQXNBDjWCwruYBfATpsCb4vhWGVTMhw3WwPGxmuBaZbTQ/em+Y+E+8M
TSwtLoGTfpBiSPNfMDeQWnC0HQr2bgab96vhPxPKjEL1wyYRy54CTPbJ4VeC7U2g
2H7oHBDtNU99E8KihkiQwssEiMWUEhsKMcdSamGGjA3WMBCwH1yb2FmJN5ZJRJu5
KUjLzZRvgD3Q1L5PW0HRYwNbXLU9c4QeqvSP9MzbO+r3dAHAokNnOaFrPANytzws
ghM9OIjWNWW05KQ4LZUglDsbUmobFVDlnJhvZxz/Pxie+c5OiPpBvzpiFgzccIEA
eLCJbBFfeb3rSr3hES8eZYNKa7F0bHFkAVajx8djwNKqwrmiNYk4VT3t9PuGKoql
manZ4sd5ocsuu2MtuDuTYlTIHZPEWnEBvUp+HegVS/Q3dhpZ2W8yynnjEzzm+Wpr
uU12Q6NHiho1MrLBjpLIXtV1wpNu90xn2fI233QTiDH/Vh6PK8ATijtgSlpEBw58
3iT0GeUWKwffeDRecVpjqtNnJha2cuvxArsJxti5OE3kQRO/OA5hImnJ4SOEdonr
YF0kuNh9IuaVB1anhjlgE1PF89qqaS6HBemm05zzTHq0GRqKZ+RCCdVOE7z5jneT
+UkRbCec3HEUAshZHSruHRctnaiuYpI1vIACz+DVa1mWcLNRaYurpG7kn8fxnRG+
2Z3KLd1q57uvXZBEGJxkuJVHPywKwXv/jVOejoCAI0azu9iM4RHfyBH0/KMKfF2U
QG9hWP8sgLpr5ZEL6g+o4QMuq0wKc/QsurRVVnnzaQyZo9qnQrXdchGg2ng1eeYW
nkouyK1fTa5luAuRrrRxctLO6TTwTEBBVB3Pbf5r/Lekf9E/dJ6qfKG8gRMrEczn
UImG4EOYiWQ5lw++naV0EuoGzWTvrV3iNzvy+Oj3+Ql5VMjprGYGglAQX9bRdTC7
BSd6u2zQCoMDuFoA/ocraTAwkvMRvAuBaR6rS9k3w6h7pFzWU6uMt0X0JbDhXDx+
ueq1Zz54CKqXvFHKAmq8b6is6XVCRoTXKdotoumNlYn1Y47GBK8pSaOy5+LJANET
wme92FJlVNt9onBXWCrBRTQKO6om1xaPNErm7479Bd7grmkhSbYqGu4YUpIEsI48
uyUL9D6JAsWr4pZOlNot8SDQYqrdduok/5SjR65CwgPhtW35XCev3x/1EGQNlL5e
2xxPc2hAFmv1tobG27WHQGSrjWSYNlsOWpwqTGmJcNLbngr8Hl0PBfYaqZm0opnx
JGVPfSB9ewloBzeD15RThGR1yFq2vNqKL7TgRY3GbFJalS3dBywvLCoOM98BErTl
9121Rc2tEjbXmRs+eGoo06aTa88xhnCVftx1bloNBoJAQHMizOHIuv8P/Adx9Dlf
QSRENzAeMW4yEv6eH2Fhxz/i+zVA8GpMqKhVIKgYbdZ4ch5+9kxdOlZy0VabhVrq
G0DK0IUp0frCZ7uB032kkqnwvAP/vtOLVi8mNcUKbGzHMaSnq/XoekfZMxmdpqx1
/j/DQle6P87yxgBohf/6IVGvdEwhN6973hPb+oOiPtZmFRN4UePPiwkOY/enPyN8
YzmuoA7p/MlGviG4gSsbj78TS5UbTK+Anhf8GSrU7IYsYEM6LH0oAdUrRG4X8qUe
PnxbRtppR9DMtL1QFzgwimDeR19bc0o9k7hEU1bCyj/8mc0vSljAScuWpBDciLZv
+cPfqeIzsCetA8WinJM4gRKS4C5WMzBQCZh9ncmyXQvb7bwWCfw2zvUsCwAjHC8P
A5PSq8cKvrH4UnqY4b0Eo7JW+jt5H5Rmx/XsoM2IeBWASAKzV3BzDh9r+LYBWaLi
8wUlJ1BL9XCBxx7J0aWNhQ2OYq8Fmgy7R8q5yHYCIuU1oMYJQEEX73SBw3O19Mdk
kQs/cIesD7lKXXzvEbGK8Kkw4zXbEtNV+AnQTxbnwhvITVagdeUWJw1Vf1psWSVc
102pzzpIZZwTVrOWTQxhF7yD2vI9DocbwSRLtz8ZDxJaKA2I2/IwAbVbx5JRZq2Y
opceaBRd6sPA/1MywEJhyp0t5qbpQEXm/mRywodfa69HBLqDOVlyA7bxggRE85/j
nizONtCIYCCWBWZZsgx1ySjiQmZnvDWooFp44IUctvzLfpyZ8Jfl4qxwjv4t+nHq
i+jK7B9R7xZ2zYLpMUCmUvvyGU+tU0z0yYC2EppbWe/+mi3//JEGy+rQ/39i6kXv
K2MjiMeayUgShFDK2fcHJovO+eKTfeHoB4esNnc9BzjWeCQI7lcDTQaIQAii1x5R
mBHNOe36SzcQTuhJntg9H5Xt9M7CYOSVrlaiB9bzCGNA/y1O25ROCVi+VGL37d+2
D0+7PF6k80iRExjf5pAz4lPzKuyfVWJ3D2tcmfQ56yhtYcFBBopW165l7Pu11BUU
VGEGHbyeB2l+1fQqVmHC3NDDiTqVvNDhEFagktdMeaegqXg0HI0c3kYklHyib0tD
cJoTJlSasjxW0vAIuK87Pq4hY87D4NXQoSp1V2Yw6m2Faxkdq7wk7eHDHVfYwK0C
i07DfKetfCn1/ev9Tyt3xqEAnLDNcoFeoOvTGHmh5vY8fiSWr2LbzOy0fAbo/eTf
BRzl/RsEJaZj3Zywj4aYqp6ky3qDW8PCd8vYg1K8R7ZL/dkOl4dtkuy/wBNKCn8S
vm/KqdZ7VbI40X49KrDBoKSYnswmnWY+to33QK4h2cb0fCap2zyBNBBqOxCNq7Fm
jCqq0YfrmMtAYyk5PNbHr0LWQzF72DCNQdB8CqNFIAEbrkbdNLEduw0uKsGQ/WwK
IvKv7NcMc1CZ26JEiHX3xHyP2V5G1ONITeUVQlmyRWuMUMC1EbFIEsAd1ejQ0tZn
2Vzwmlox34WpSH/tiNWo8j62n/nx3bOaSITk/gyf9wV+281L623mMsNVrBZDph+V
/TKYOcXk4D2dvlekDxl3G15N4uVfHCm4wE614gyrN6nK1n5kpZC6pv6jbAC2WZz3
F+9lsNArPKrGGWYba5xsj5rF3LOqaghaOo3v8+VsUScXJUK6bNY29DV4dw2+QcNZ
8vXRKEOdiTU26e3cZOkAGsewOQMJuO67OlFjPNa/dwMBtE5Bv9ybnttUKMxV3h4D
44hWcnxKG6lO6a+BLUzhfozw5/29MUnFI8FIDHFoz08dl+Oyv9vL8czOUjt3S312
KjOC4S+Ow8Ue63SQPphfDLa5gbRJddPtWQn3KhRzVh591BjxYJqHlOgDf/dXZp4u
Eljp2CMvCg8XHrD1aaLR4LXwZ8k51qp4HMFFBY7/FejIEb8F7AwcS72b2F22dWiI
I5/TyjKJuIvNSKss/ud3N+kGgKIKcSd7VQUZQ4v+frSnPCE0zHaavyeNt021YkA1
X+qW6pfyOX1zBAa1z8ylLwzUmmZ4J2t2r/hfgitT8yUeGHppuiMq/0MgWDms9e4X
uQ5dl9KwoJUmrl2AUA8q+h9fhq8zzoRCmPkxGxkkqaLqCNkUkq94f2rK56jjz3d2
RcYpl/IiEZXGLwDEVhl0axIiWSb+fSpukQElAGOsYk4nyNI89DiwI9XNXAqX/J5x
4hmScQVyx4wPEFBSVKisgVD0ZmuIPUV786UJTqtfgk9rDs3RN9jNfVAiSbNL5bVo
s9oefhEiSRNqtjNlNbOay+yRx+flcSKcQULysJygtVVlaJXN9deyy0ivT8TXPkR7
Zxo9mkau4Ny8ZOIBzK514M73TcyrZwnQ3LO3PCX4514nq7KwcnPtOWHWw2q6yyn+
qSo8e2YgsymgymIMRM+C2DRBkvhuea/qAc+mGT3a//GgfrZsE0tYHvBeh94LxOca
ONkkCaDGEam9GWtsd9o5HSIA25yuE+C+/P0lN8X4sjA510F/XiiBsu6ZYTt3UolJ
ids4CDPl4QvkUhU3zOqOmO9GIn0pYlj+Z3nssjUU6MZskXujOkUHJODldvPnhsEU
wTHRO4uCDtZ94e7W1PNC8OyVL2h7BhtaayzcTOcp6j8rgl+ZK5o/3qZrPR6q5uPm
eRi1ADmiqkRAzfhjbq+C27UhZiH3nxMZPQbpJiwnBGP1L27Pl5SBHZIwZq+l7z5E
l9ZRWS4oFGwwrS1SvV6c+Muu+dVPpyeY8v0MyMMj2rdhoO7NP4M+yvWWzPCPx9Cg
3Tawe/mxNakylBG5LkSi5vK8irqlMU0IEpTfwTQTZFn170A1dKymRG1lh8DQJol3
ULf/GImD83Klye5kUBulgMQycTZhIhomLtQjEh0sp8tma6RvDVN3fznWJDxqPtmF
wLtloFI98opJ2/Mwn0NbecUzvIAn8WAGzbfY1Cb1wr5Qdc+G39z78Iu18Jn16KIb
wWTK2nn0NFZS9r/qkMIH5+XMvHvSaP+Juo9nFd5/0Tr1+uX4fWJMVO2rJyLXbhXA
tglN1Wan/NruSuXYaNAxU/MyVLdENZg3eH79CRlej5hkPaQeFD5r++RdqPDWKcp3
edcQPfiEGmeO0eqfaN8n+0ay3bUsRTb7z3jqpRe17ctjZUl1OFtpXyL7PUGgSbeW
rIIaiKofPI4UKhL+Gdj2U8CXGoZ7iigP+uPjuctDcN/qIg0Cbd56U9UZdZcSVN4Z
BkqD8ptCNVcvzCErjDNr8gAe7JAoy5vx3NDsvUbyMhRdpXNCZO+WLu0MqJfbUZkh
sphk7EjW5XpdQwGvcDx1lB+gUerov1q3ZRDeQnJtDsel4VpzPZ2B+h7mBwvbiqH6
N12n/grUrWqowR6zK9OgpPfwEOS3XlfjZlQTS4Zhyyuv8nzvwbr3w8nJ7MSnwl9i
hytKcU0wcZe2fW+1YqEd+Vsj2XVS53j7VBw+PwJ3/Jp9SsNPfPVJf2DGoBnEbbrI
S5fmw8WsUz18r+mbnPRVrudgPoqvMMhQ2o5zui8mkww7RorBVSVscPH0VXI5pO2R
ILXkyo2hbIZ0f5JCsY7yEjVH/kzm2aZKm4OPI5LZjTPB0sVlmu2mjNdIB9Qt4nr+
aJAMwShq12StmXJJKLolcWxuMud0ZdV4A0s+I149Owf8EED2K+Q7SYAhEhT0YsQ+
RT1HgqIFydOh11IfJ62P6WOyGN6h2qUrzbWMrA9Gg6IOPPSjZoQ6m5DEVTmhsc7E
WHx2VvAIx/vWJMRHGyeOhEd8SzKqRifUaWmh0WtaQC3nq739TPasrYk1IRCl7/V/
UuKrxuhSPndhRxO+tg64+xkoFSr7/lmXZA2J6TjDJI0vNFOtEJyRYmqkwdCD8S1E
R0F3itHnIBcontDNF50k2cqbYWYjeGS2HkfKdm0gOudQpwD0iGRhdbNdIIdQq7hK
oZNQjk1KzW4yaC3XKCwbkiVmbXfZaqYd/uPFGqgvUS2HlzILMy4hB1WXRj4vEww8
aNT53irkHOsFiA8zBhCpt85xq1qvpLBnhO60hfo1zE2fEhRpn7vGMmEyvvftjbfQ
KE7piSyoipajQFpclis6r37pbtCRI89IE5O45d7IKo/BNtxDNHiSirHzbyt8eAXU
8F8v6IzbnTH0pFgRd6T6Ng/rs3CYrB60vSCVPofNx+Yplpw+iWz3tD1559zm7Bty
JrNPJAFeUrUbnhYVXN/CjNhDRqPx0nA9tjH2Va+2l01kVzvhQDOA078Kp5WSJHYW
uHHXaQD5WR8W4q+QnDBfa3DXr8ObsIf2bvwhTwHmZea4RgoCCFb5dfNEinQMMLvw
gM7xDBVRSafuTXpHByQwXzjKkdpp2WZu6wK3mD/fZMtgpyHbxyEtjaJCvGr7BvYz
fs5G5mqNual1eoGstwTKe5rmS3W+RTXrbmb3qEvI/8UoYv8v5T2yd441+kjz8jVm
XmzoVMhGeR23gHzU6dnzEUCs1VMgQgpi1YCswysyTk55eMCg2iyfDZjIEOuZ5Adn
J67AnxazNGePHuC1aMTLVgJR+S5fMEoe82JXZ1Y2+xCZbmIrwbHL/3wof9aFaegb
L4JqG3tcMrsi71xXhO5M4Eo9V7eiTCvVe7OPDgdOwmneApjVuO4fxohwJluTt4xl
QT8c863+/ldCxAlRioTNfQjY3FpHPGkns5nsSmdcmWsTm1lcPaaGwaqMXPKBTsW1
xG7te/IwMxeyHKWKP7TTvx7Ff4woF5a6P/yXDe4n4qFaHyDnjfKfQstQ+LFF5kXC
0DP9SBK6Oe+Zw1hutEvvUEoLlPB/qFhRiaoybFsQYyQVqNgeVh2do45YFoJXBIfj
LRvseIX8cKpZdt9jA2E3up8A86eCsVrjkbMgkxcJmf1XM6G7XUsmDKo3a4Gyw08/
6vMADl8lH3tJ7GeHK5rR0RfoOdGadRiPSzMABu87RMK7lHRmxX6+z1oLg3iQaEb9
SFpSNTFxjivOcdceys5kAfOUFnAQTw3fDrWwzrdlRGXDvgM5c12BxGMqRPhpNcyE
pvsofhPdpQ03Rgvh48E+jlrd3a0cw9gHmPNk6BfI5w3QgO6BCxZmBKTYjt+XzK9f
vV+0UFA+uhFoboO1V0P3f/7Pn3EE9gregaMqHThn4STq7E2OCJJ/8wuWrJLJIlMu
PbuihGMgiEd5RUKJuAFnK6xRSHzHWtgw2o+kX2Cuan8TDUAqB98clU6mbuBWBr0U
RrDg3ZyRQWmxwxTj30g2PKp5xT8xwb80f4FkOJNZ9e4OjfzGQitAPARvtNSIVPEt
fP57wpPqZ5kKW2E/4hTJo0J4ZYH5AyS4VHh12ACW3jSLUFDWPnOM7+vCmtJg+T5O
0O37tD45GIXJVno7VYidiIqzpoKwJ84ccXe+7NPuB/DaU6NlvYme+IDBe3uJA86V
S6IjB0IOUov7bE2QN/b4+LCRKG9h4JM1YwwFUn91a6CzNPC9jKDroeBun0NtP9Zm
JRZ+HAcj/ZZbi5v1G0TpWe5B3hLKQD4UQl7Dkmtu//3QTIfOfNw9m+BxZ6WVSYSV
d6r6KGl2KEd0YZCUBUa09qmAOaGYYlAMO3GNs0fQuFjV6WH5L5Orsj/ldkPZD2UI
0+zFr9af7X5qgduWQbqTYiFmRLmJfJhuipun4mXy61S482uPIydysNR1M5skBOLt
nMc9UYU8W03xMLKhc04Dj85C69lplDoAzAipLd8Qeq+Nb3NUQolZ5kU6pg9eKpvN
QVxLoP7cA5WIJMUK6iM82Tf/v3x5RMmP96fRvUnqJDQTHkug9oWQ+c+LrvE5CNqh
8fI0Vye7CdGSYmP6fCQRleEY35AEIm3x0waTBw+t9MMzpIfIWldXOiawZU+DZJ60
lhl6MjZAVkNBFiJNIo5gYhluD/RhV0MfeAuW4SR6R0uRu9CaZJLxoLDMdlu4Qqf3
79er4T4L7NXPGsHigDKGH0lYdmbxjGkEV0Rthlz6/qdibkCsb+8t+gKyvDrHRlQM
jtDtKDR2bX9zl7XY7GXNSudf2kda8v//GLIS4ep+ZS/PrR2JZVHo+3UqZfJHqC9l
ga2JHOgTDAYk8ZhWseBrZeu8wW0vR1hcttL0w28eOUwMGBHbCtijbQf8oukt8Vob
5FV0MCWnF+k4d2l4vRD9vGC6dPKwthcQHnZnzdO9fiEwwHLYTN4Jkm5SFoxI+pMW
tQ14M5m8QAKYbQb9ekUIGUnhqnJ/+MZ6LNp/c8LPPcNObMKXakZZ1NQgvn1P/INf
16LotfbncSYGlXH55XGLTIUDmjIsHJfHwKIpiecfQm9MJW3LOKdxlfsKdD8DkNWC
I8/b7PVFNuMT1AKhIEYPeJZksjspquTjkmQgFo1EDDHx/JJM6S3wk7F9u0Cs5Ok+
XSgIO/c/ykA+y8Yhgw1TVpcxzMvncGyrGh1uY3SRUtaYPN5Z/Pp/DJkRQ12uiW+t
ARMumXst4wLCtT8tRGglV/a3LY1QWPSVqNKPesQMXdiNsjqGWfY723QymxKh173x
2pTb1kXiblIJFiekl38+RWwNUSBR+kH+yPaiotSLHYqHknNHtXERHqWLngNAmptE
SoC76Lr6Kyw2Y6izZwGrv/0wC8y2DT42RLNkUmjmUxG+ymKO5YUStUPJPOS7sSS9
8PSmTuOn1FrqriczYM1AiC44loK+jJUwt64XjnPxuMiGYxAnEB+sYOKkyz71dXmS
6lK7Ek8Wl3f47pdKQfsTpHFURYwVy+PqRI+MBudmTXOUy+IZji0PxT2s2VsQm6pc
UwE9auuR7lPoFSlNvlUt6RcNR7xyN+EytuBbHqHIiRyHyS+Gu2IxuFcV44rxQ8Uy
9Yl2RgYQVk90VcdNjOb/z5SqzXoPiDKV2lCyF/eBbBggRby/9huIywixBfQM49Bu
sVpZlxmb2UcJ8xSSQmTFzJYeHUge4yEExS/RN4VP8dsYDTBQb2whXyxvQMbmLX4W
02Ltj0zWBOExZLqXdtRHC9+7LrtySj99ytQiqhZvSaHS4gIWkTp5IefDhSBOp0E4
VUCw4sBSda+1lQAEXMLxZOPWEdjVAc6ffe+DTMPkaJOPcAHNjwSFupK2XYUJm5Jp
JvTcFK/TvlZL5wGHy2EstoCxayS05tbwKNbfdmxmtuPHzyyfapRJF2ofZXepmV3c
jVvduXRhV+pmj6tY7Y2lC5w69P5G8AWOaETp2M5LgmysCuhKy1/suCy2rdvZeopB
EUSHvZpy16CpdxMsSq56TSEi9X2VedVl7TCj2CNNT5PIi3iP5ecY/gRaEJ/v02ps
5NvO64/17e4qY7D0ZT7x1SVC4TeUGs8ptC0JSwXvhfShxEiysThUzke4UAXmtqRe
Md2cfFVHXsMY1zyV6URJ+/zdIy/tTVo0uFk7whJDW7nJAFT/HbmXT7h48dxq7Pem
TTxZSvoDNCyz3YUQZpN6yHZ5JT7xznGGYs1oWl9y7RIAqFmwq0HBUi7dwGT+3J37
/7U31UwWcLmHQosfaXwi180fDA7vGZzSNJdJlAhWL6vHdZTyqn4t8HTiPGLj9vAQ
K07kWrxQxxdMDyOJHPO3yViweGrYgAjbuCJUDFVX2Rj+o9HGML/V6XqsS5awlB95
t4J+zzO0eaDoV+tLyp6HbEWyeaB12S1OV3gVYZZCsSEAGy2QPr53XuMzTKFzSlY+
+i7hEQeKqPQfcwdtw06e553IbzY8ZcKOs5r1dPD3YyGbHW/Cmnr0PMDSm7ta2h+F
loKyLfvO3paSYxUi0EPaAdXmDxekwo4gEAy723nb40FElLUSaTgwumr7nJeS/fk4
emlcUP69kcp5sFwaiPfzTLozhEoEe4kCYIc7gUAuIlb1cckf6hRclXPiEL2C+20K
Lcj3VOunCV5HkSXYTsJKwKTGgus89yFPZxuwSTm/6hc5b9joYaTE3ggT10Ox1wPG
2hbkeReFbJ3chGFu+jdzOettabJKrxA1Br53aenJaqV88h5lSn+gUKakdZjNvjjB
mO2RZyMseSDNCp/KrmhMSHailLAGzixQbxP6j5sY7Mn4UxWQvcLjC1PXR2323IpS
enOXWatUBTM07pGRNIloKNBx4IxQEZud/GDMV25w0rioeZkUL1C9ZzY8NLaClvOg
PdHKot/rEoNZPyvKXkW4kJhP07psbBEzzbjwEJPWzSa46tCmk7XS9k4iKp3yr65X
lZ17/mX5zI52RlOiQUz1u5gBjMjBHEdNhJgn6DbIQfxI/QfXTICKWK/lezEOyWBH
gB4df5UtIN56YmBHUrAqfizyjlR8HbbWxtkcciSIZ5cnUjYf0k80teXvdxkPkvzE
zmdjjXyJS1OolXfi+qRUiikagsNLd0x+CZNUMEan0gIZ2W3xHB15bm1vji0FbtdF
ZDGdhA8Laxy1NNavejBHpOn+msqDbqGIwmDP4yZAZOhjB7TXan01qdXykYVU+J+Z
nsOLIkRbSwgpsYW5Q3ZPP/asEW+wjbg742yXeRGzsNPPStF/+aKz24WG7tIRWjN1
vaNqQq3juNTOOBNJV+uID7VC4dp4x6s9aTMxxVP+v/aYjiUs0XFR0PSOm4ASBLVg
50IYeaIT2XK4aHw6hWIh/SIHmJympW0eMFluxLkuE4Aoy2QdlikpUQ4fcSF21VFb
cElcNaNzRhurU2zXzsS86DTCqMnU6MphZVpQDhJ1FqoHc8ipliOUSlYbXmvmwbF3
h5/pWUTsfS3h9uoXncryGoutN+fVIk/L+BmSAbpxyd1rXdf8EBhEpS6iLzd6mrRO
qQXjmiyHZgi+aKp+oUMFqSQcujxCtS/PlR+Ewk32cMxYalMzS/EVP0TACTYFFfhp
YlwjIUq1vOOb0sOc2WIAYa9yBNlYd1hE57FScJ37pVpQ06noMckfJfQ9fX5w1yGo
9FRQgXqDIZ5I+vnx2CNcF+vUMflDWOnYOK7wg18oGsNGK430pq2UFdnHavaSDwaR
hs0/0IawPoepwBOZtXluR/8hxa3lhEgWV1PkSvB85NuCkC14ha2yTIYxgmIUVjmQ
VcGyu7CNg62F8Os7m1ya0cszy6qv2WwkqlEi5KQO3xsKClHAcl5wZq8iiX2G4bc8
fe8WBFkKloorMtohPnu/lM7Z5TxnHIZqgZoI1PnLXfENkEWGt9H2U7tQnOjx2xoA
tY4HL17L3up/+4NPzhtoc4RAEkzwKgzxQ/qB2rh6rPkXaY6rzQBnCcIiCAAs420k
rgU8cYSFp+U0ZT6rA2OUpV6su652L/P49mzH9kBJT3jXzlWNPbqQj20Th2/acEgw
XfQ0mqybcLK60lNkIn+tnFN+yw+o6LYoWDuz1LoEFJVsaiihWWGGVhtPWtk0EHlj
6xKWSXn9fdzh2PIGSj0KyolDEa+Fsv1kg86lcgq6uxjRdevQSXkzy+GIKS4cdUrv
93FQTBR7OIjOeMfZH1UzPVLXU1tc+XjntY232L8klp1Di7iLevqI5zI28/opMSM2
7iYkytecLzgtCXYn4TCCP8d3HYcf+ZdS2mXoPmtDKPVT6vhndNNJMgtji/1Wb2Sg
EBjlLnxsDcmpIBshcdcBJ/y+m+3yN48PVwEglT0GQC901c7BMfilwzXlvYsvULDe
R8nN1a43hfMiqyc9sLRd2vvsQPlhK3axUyNXGhyjX6Pd66ISPevMKEPVkbk9ybSL
ydte6XW6JMnn1jDzHO/MR/LzbMNoWS9jBScUnHowwn4jNAayhpM5TBNLGUJAtJzb
mkUjdfZ+n/MMv+mQqppRbgzDI39YN04Ax75RVwJs/xT4zKgUhIlhiAOiQ9xJPmFa
Zoy8+yUfUKH3kMI/RlaqPikbb+BK9Ol1vLdE4eMv1UrY/hwdnQftTLm+0GNw9m0d
zU0O8ibYe84GUYG1gjvTGT7GroVMzMMR7S0xuiA5g3EBLArQn4RdpqPCBWWBpbCD
gI9j6q1FPBdiUq7Xaxl4fQ3gUNqFogALtuwheea/Z7nGgcz+MzfEj1gj6OoLH36G
3OtX1ObZD7NmIDznbujQumiLZQfqM3P1/QaIiFs9+vtjz3ezxIQ0POrSDB+s3cPZ
N5akOx9Pf42/3MDTtYvltBtCUICzcK+igvxZ2r+bxMpfCVyt6+l0wN0vWSL7XXeq
E/2HNyOG9aHh3gW/HVWy/4LhMSteb68ypBiyWU3U1TQdTFXWLExMgzaGuWffdD2A
HemLPh0TkwmwDz9R2mNe184SoTwrDj+QGaahCigWKEernxKV8eRawJq8DVqz5CTh
+pPR962jAIAnB32EF5uxD2iQ6DVwhHRo2KGzrSD5ReKksvGoyYiIcWEgnDWYsQFT
X1HDeZ0oZeEgWEBkOvqvFWU94vd7/pHeJUA2juSNhSWYafvqD5+1M7JcaOd3j3Jy
eRx/WhbFICBDlmzjzYHVMj5JBlmhQ9e8oPh4wcagWS3ER8LtLl7ay+ASGqL5eWJr
UJ/mHDlYGzr0JdhiwRW+yI992dqES28gYrdt8uGbWFPtWAQr4KdLqKPS0hoDRQoE
TfuNZPHsejPtICKOAz3QyHGE4Y/I7pFx5VIzLK5oYX7AMKzqFkOtzxGmO3tvkxkP
V0ROt3rTJxUcGuXhRS/QqxfmzqVnVpwmUA1OHM9V4Nd1xGwyAB2f7x20dbdOtIBs
m7thrPkQ9NL7+mFb7FJtejSUZZhx3eos5veifaUqa1j58QwE3sTIpc4okoAfElvJ
CrKgn3Km+fNoDSpF394h3/VFQjkigDXkhKxYTFgVXovHZSCxQy/SvIsleXu8MG+H
zliHIPUUYTlVSxJFiJZQRevq7dC5hVKTGUEvzLnJQCPW//x+RfvjsyZz9ib6oGea
ptJT78SJeyWQ0+L7i+1iR1z8ZrKO7btNRInU4qjNt3j82ZJRX43ttwGazeBUyIi5
87FZDKPhV2punzZCO+vfve69SOrKWuL9NGGncvH6/NZe30u+FoxxDfqbjnWEZPqK
OocrY3hzBMUgHuf1P3DE77D7KRLbgbohQFEWPKq0rWRycjbmGOJlFc4MrgLBxaOb
DAAKDetIDWVfuuDB1u0mFgL+U6ti+OJLoYEnJA5SFPSZowQz5+h3eUZkiIrpcV59
hb1iR1Tgs4tHaZjrL3GZuiNzw2zwzfmXzW9G5uMRrO9pbH8BE7qldcDa6OXSZdp8
qIk02n+JjPWezsoMAjFPyN86qZyMHUmD7sft7Agkb3YbByanutOIQUmG7gKqkRZm
l8lDj7c2jq1ZPEzLkJz8PSF6VpG2XmBY19ytOlbzj/BQysofWyVdhKzmePcpfNZZ
5vX/llfX1Y9FM4f9avqR5oClKg5oL1XekZMktmH2r/P/BkJ64nrtOuI332ijA1YA
vw6LMdQSDzfms1iPZk4z1AwQ9NtuHEOUMfGbFKz47DhBzW730IKQvAZSnTi3kF+I
By+QMRBbVu5cxUVr+BFkGiORsCc8OYo4+iGvCPWFJOJ8OieiwRyoV6Ri4S6nZmGF
1u3uyOBq2XpnFpOecPg7W1nshWRm47c9nN0aeKilx4n766+2ov/GxOcx7vSD6y6h
hM71s3aCp/GGvnlQ66fDPryDI4nHY8EzlV1Mh87Sb1SECbQMmja9JdcFEDg/uDee
vd9OPuQfSTnvQ68dxKqHurSTM0IL8ooBR8TR1jUg6gHRDOIh1rfywFNMsrSy2Z5/
0WnYIgTQwGnajDRo8yUV0HqooWB9csuqY1jnb+WfGFVI3AN/wIy2GweRUsAIqqoT
vfcz8deSlhCLGTlC04k6qSUxlwqJfWr61O/O3PO8tpSTdWzN0RdcIS4y/MWKimQw
z1WE6uf6ZKRwsRGlbMcsCnEALPfaHSyVZZXWEV91LlqERasVK76werX2xd7i/1BK
Kw3lP0ibTkbxyY9G0Q7daTo/B0r3EYXmp6JbRzpdfWC0GSuCTIGVC1ypYpPrYriJ
GJSdIyVVoGcCJqOaeAJ3fAtxrLYplHwwyZ3XVvoOUXu2VUGoHth0YLOGQTWr+ANk
PZjovo0uy/6b0dPyVRL1ldBpQhC66OEudSzFDg/dowUCFMae34h64BOGnNbSAbfM
9JDNGlUkD37peqDHHLdzWOeGimwxA18HYsKBkYbKMESG/bzl3TrzK4K5NKgDsKZr
W9TSJSFwW+PslibtiJiGg80OsZUbrvfda1gVLZotJbstJV2Ha4TY1rUQixg8Ykps
/++CTSPLs9if/QuanbHCdOxOcTa7QvQGoZCls0Z39clAOzDPcKXc1DnJXocYyMcp
1afNcb3OpKL+1Yqx9GQpR6ZTjj23/kPHyVCvo6ajFZenFsK9aSIgF9Gq4XxzaSgg
acIzCptoIoiUcl+ytcI3qerCHQtaFdB/M2lQ+kzHPmSkQE1SaRaUDGimQq2wMYHl
GZNqhrWHGO+32taDK3scgUyR2TylyJpz/g4h6YsgFLePxK25DbB9h2/1/uSKhQXj
EI2TV5G9NBQQaFhyH/IkGEReGTs3HmhA2PLtCwBKnUZeP7fVHXtoW92uP3UHIxyu
BR5ooMxS7AXn4ywKXoE6wbDYb2ipQax1IZJGGkoaEQ8R1gRH57yyUqihlovBEY0E
7qPbfLDPIixc4UGbuAnmaSp4DD6fimtTn8Ki3A4wTHL5oL49+NiMDkIfogOEmAl4
+as5NBLce8DFv31MrXzbGOtTidCboXrrvPKYd9NzYay9vtvEGRJd8QPb/I4KYVS5
23w7Od/XLCulsbEGdDn4R6Urf46JtxqlZl/8FU90JqsKfWK0cEu4JO3w7CP2oxbH
BXfvSc2VzrVqkcx8YUczvIOkh0R3enR/QMKwhoYyv6CVOhulwUd6pahyr08kJtrW
OWZjvkLerEjCEwttoMNVCEGGEojFYTrowVBYFRhRENzj3Gj9pK5zBvDipnukqbx2
z5Kvejfvi7Ea9wq1d672qlbzOKDvxX1h3Lmv3WX7MIsWnAFdWuxj+ebAxdoWSgOF
fbzqhNeUxVYSuMtwzmr42lqSO63VToOCQfWLzzTbms7FU9Col3zjU2M4IT7Xn+PA
euFR+B3U2Gkgr2APkLzTg+bRxPhW7w4wnN6dpCYpxgVX7kWIOhnJhUA1MzFvcVrj
SpoXGwcbMR5jkxoPRdPtjrSVZTPpPSvaHtO4JWTWLnNlILHoWKfXDQz/JBQ9+uur
RDv6dBnhqm9g/lrNfp46YZj98UtbDC+qV/hzNcn1kYyRS1OCnYpg0zX91o82WGj0
uVxiYFpFJIaIizMCVPFmVWw1FtTyY8H1ZD2UAM0zSYNvN7JpN5HqakCoG3jFxP1N
R3c0RXdrJi76hc5+ysjBkMrPNX6rjdQs/MSYafQHLz76bear3DIJb6Ivikylt31k
PaaSCHm2I6WPO038cQu46giaQR95Y6VxaMgCdTVWPDVlRvpnLrTqKe6pIZjiTg2f
v/kSMhfcf7RdnkS28M8ugwiwP8lDPIpsO1auQIVdjCRuT2nIIUl4c+FcMImXJr/P
3fIIdjC7pNhJubOmvha+CJ9L0pmgvRRFf6o0WBHToQNtt7e/jzluPnuID9ditQMD
IPP/N7Xj+cWHGlUSFcB1zlm33KgNGKIe7MX11wWK6EG2epgRR1B1YHiaTCEOOX2B
MiThgjHEB0EsJu5sJzB5nEHYjHRIRTx1f8FyMQg/+clmGgA9Ejt0m/rNiVUQ8q3W
+qlMktOzwE3LB/wQH1EUwTmSGTfVhQqpw5+mkZKG2TAz4nNj2bUDL+0FeFHvbHf1
+eU5uNoPpybb7cbr2yA/yk4p5Q1D/rn/frDJhQPZck4RGTBdBYSVIHFLjG3J0mXU
/pJDhw+Kd7ywSnH9ScmAiwgbgSjp5E8Q/iVIZvWWyfPpYhuN1tD51rF1CjzUrmaE
0IfvPPYT71zlB6nbBvJDFi8yewZwBeCPxDt7OiTI/Sffj6qNa6bTipwF4l4pdgGR
awrsZK9d4V4C5C7kVLmWSybTDCPJj3E57Fb7l9ZIbv1klTJg9SKtdnsdTitbKFyR
uiPEiFCeQLKgotkZi9ccmGrLWV5dGsn2Z/XX7FyYIeq5x/VWUJsIYf65iCIv1leC
AajMiJKs/8bQuOZGHix3ii4VbrBbw14sZ8TwxZD1bMKb0YJbqssG+xiAs5oj1UwB
tlJKkv+DjdJO5ZvVVLHc5U9KekwBFvUcQ14yadx7JmOAO9sLSOLOTMtc6+v85GOM
R5Xby/tZYo8BpQbBReVdfiRKc+zH3Q31R6vWplaH8MtPFxxgppwlfh48HmKznzIW
2beVW8NfZ+FxsykJlB12nO5gW0nB6dTMVyBL0cxz1bDAkQ0YldpWTpNV1T2XNhHF
ia09Mxtm1clpAlNbK+Laiv3ddTSFDpcnrKSeurmmeFtjN3wJtsMmZUVVEahfus6O
+7QrlAO9aBAZCF8o8IqovnVU4uTmXJIJX7Bp2giF9XLJgPwEukoRJrKEwtpn1Iw8
Hjtfw2N/ZyvTR3kpba+ud7qnyIq+UkkJReobcgq/RH5bQuEPHEh2X428ebT6NVIn
CyImaRDyXdIDxkKDZOR/53CfP8Nth/k0zyyrMRG0Ec7ZJMxZ4XFdH9tjePcAXPtB
27XgtOJ/EoDn3kXugZbnWBOkc7u2uhOPbBTnqRtub6SXvg9uMpLzjpi4jF3yXYrC
UAa8jbwQpgolS14yrWoIbekVBFmkUUERvvFikAXWd7PcLFIk6b2SpAA953Jtwxn0
P0Y4hTuw4JPmpabdSYUApU0T7QBiLIt4QOvTcA3+3AsO12SevHaPjvQNEbOR+75B
cJ04FWz1J8aVGktO9ZHxwOXEC01x+TBBsQ7hWZoceLR+J0lmnCZHalLi13cYjAM1
SBKBDM3atTdAN1sZ1y6KqHFcx1YjKyTpAjccGwnY8zxIqV65nxDdnX4WZm9JA8Gm
JHGKrPxKTUeXFIg9FYMy255xpkUm4cfEHxwc+uQ6B1fjV6sZS6KxHAclmj/Z6+7w
0zlvSzmhQLY8n/8IhatddFlX1YSCqPyFJWyMxKz0VB+BnMw3qNJ/rBaB6FhRtF2r
YMcNhNys+syoIVoQeU9o3aD69ZC8wSkLQs4VdGsbZ6WJPpdqS9yvilsr2GwTBBb8
7UkzghQeIod24dHLbCTlqWGq/qyfv+Btp9u449+9TAWI9jDfRl0M57nWwnMG/Jyq
cSi0nbTFQeX3X95egHa+I9G19MLsyjCAHbtLgXMkO2GxU1jwPc09imFj4WvzlsC5
DalqYpuI/Lx5kHuk0StTPMTwU2WxLoSetkqsshBD1m5gc/EPI4W7paraF5GwTqK6
SI1Uz/LC9Zv5H6Z0T8DNtQkd4nd83TtLyd2UDTb0OFp8ukaHiryDT/GE2S8+Ko0S
sgqlkHv7ltuSTYsYIM+9Bmy0ST2x3MlRXNG5WP+oT3Myqbc3gSVmrWaHGm30Iq9J
JnVUoHJYJYpzClaAJNvDDO+DkPz4pEJZXZLEvSq4zlhgnx3B5/lgN4OhH2KYeZmL
HDbOG9MVkqDCAw8qpQi1tKAgdqUNZyq54+hR9k+u6NL4jrDMXW4c3540gJY+y8Dd
ZbrtOEbwQfr+aKrakc5OZflWgE2hHnth43KManXBzjQn7JlR9u1e7EQ6ovjLTDeo
Ukpd1kQ93VnFslPuuBqXFgVSH+0PNPZQ5onQCJjDACLpVdfh6v4u3fAh2Ow0vkML
K4aCMslFI9jBZTmJLiqSMdd/ZkKt7Kt3XNGUC6lnK4OdlQMceNMIDPQCzecAgUx1
mlxFTlVPxFHemGvypEdlOnu9tA7emrRegOTF9ElQWsYSPreOy5c8t7KWYqAJdVfh
Xgvnfytnporv81Sins/TSv+7wVcSx3d5rL1Jpc7dETi6ACuhv9VjXcyFjYx4RxqN
zGZ1CvV3+OPc6E++pGTFSY5pfWbnMUxO1lxx6ct/ub+dwcKf+ACjxz6kkTn7Ke8B
d98H8yqkfDVmDyi04zvALtnSa0ISA1EiKu33y4mlKRDIC8oR6NA3LnzxaZioQCZY
nZFOmX4+mEhdxJOAYbgzBKHEZpOQvQrC+/sKtTikMPH+RH1PouhC0xH3eFQzf0jT
w2j6ofGw4jglhmx7HVc98HqfcWMdvuxmSXW0qX6BE4JSXZnMMcvWhBXSFkipDkhf
Uykfjz5yVeWUUICbxzmMfvDmhC2QbVB7cs8lFVLJD7wSOu/kc6LSep8glLVzCKsG
euyT5P0BFO5lG5Pa/thZEP24LEd1cTn3Ojaz8B6Q5oloWWTm1wGYrwjBZlB07twM
Vm61oQMkvR3GhjRE+7GUF+4Rr94XuEgPxWMBanalWa5My8TuN9KIiXHkPzb54wAz
+jheKSiXqs9XPnpgiRdxAV/fM5G2ywSvrmpPZXXAVz+Rdz1sGpWocXEH13JFMLT6
eNWUCgINCqnO85oE9OBc8rsv2PhDxA1xNj8tm1VWrUdeE8CCQZ9tus9lwR/4MGcC
jn4xa+m0uo5iv8WpM0XCDG0FhVaM8whrh8p38ax8eVuCvFT6OrYjAxHubQx1WsIH
p/6dV80e46tLDXU2pPq4p1wPZ57bcpzfc/Xbo8qGGbhixb/JlfyrmoKDpWQkIYaC
hZQ1KzF2BpQM1BTP2R/EvzS/MRgdnv2ezDZBl/HvQUuzlunIqW84j1mTBlvxO/e2
tJvuXQkgD6eqFW2JvBbKeW84BBCDWJctolwnDRfcBKfbwCROkuDJ1lMa16SiGzw9
8s7xmjHPZgTs8G3CA7eGC3O4SUbl7GFBMEtxmfpUWosSQ2Xh0ZSlypDaRrql/ijB
2LA+mskS8XI84RAIF7C8Y3olI+3pQJuhxaLDjGQAxIUOxZWxHE+eHYd2Rugwavgy
jTQRQJ5oERdTq8xvo/Fkjo6TNk4QFc+yaaaJZFjJ01Fe11Ljv8M/gfhTdlGsMKWA
dspbwbCTo2E/SA14A6uWYzPmJKrnuZYAkN2jLDaL/Eb5xpY8A+r4xLIdKY2RacKL
y+UGBLkcaBm6T/ocAjsPpeB3opExiFwZqCAMqB/Nb5DUuT94DEnP1eAUZpK3v3/Y
wPgGssMNpf7jjk57PEWDZgFYhVVaEJYu6u3e6BPqdRGgil5wyFZg7HkhHJ7tqV48
2Lu/GAQfJAL59q0/BYauQGg0g4yU1JblFDSf1rjbh2sFQvsCvyTsniyaNqauDT4r
jjioCbPIN6bm8GN8AcVVuBgfb8Y2mrEC+8y9RgXxjbp6E0NbaxKkERivvJDNuA/X
ZzK/aTZhSi/VMO4eFVvaTj5adLBzt47oiuI/eV6sFjHTeBxdbWSUsyGfE0V9CMxQ
QUD5apTM3Oo9DcgzPe/bSjtgCX/Ry2znKLOzTbUFaagNcfoikiyNFUELwqu0GvxN
XLGz3cfQqcci3gFc4p+RCcJ124k7r31tTjfcw8nU7CNOeaDEXoWF7iJIJSIrJnEz
AkwPtI9wZ0TUa2c1Ivl39JZJmZ3Q7Bgd//zbUoMMnbUMjO8EJ6wY6X2mQ9AnParR
MMs2+GMz2wpygngCLkz2U21TjIzeQRWdUYSJCsWuSC77YN2+JBPD76FQs0dK8eZ6
NX3PJSK1wefLO3oCe1Ptt4gHg3fM7I/bBMrQhue9lQaaXbjYBC+GybxE/7UDPntk
CpW8YiaV0kk+f1Lhc1LbZ1vuYN5T3ns9nfeS1IL3hbsEKAPF4jsruCgkIcpSnItc
TLTPwW/T1eKoEtmAXlpgtdqbXQ/97yKmpMq5El3AL4ZmB4hlBAUGYXD+MxItZDoL
OLp5SeHHClXaDjDE/lVHluRATq8oG1Aon/Uta0bfFP7Jr0Ns5s5WkHehMEXSG0Sr
9eK5MiMvjuk+WzbxpHtbLQyeOgvVUF015Cqi8B2NwiK2PHI2xvSFGBUGKupIj2Fk
FQ942sEWOEHB7TZ7CdTuojZ1an40jOvVwVHdoMNLDhXWfeoySqarBkT8lcwgLZG4
XOynNwlW3dC7B7aCt+fcPrHg1KOiGKIdT4RcqBCcnhhlPNdDroSZfurAkJNPrUpO
cI4hB36OehJ8bWtxX1afJYQWR5ZZVhvhmAh2hn1m2HIjsd5RcPwC0PqPQ02q4Yq1
iRhQXz4DkS6AQhWxBWtQXEJBfHVmowT1LJrEfKgYPlgjCQDJc8fgoHGUVVgHys3o
i0Cp1LLtq8eCWe/GtXLAMZw2S1pIFmsKUFYaAt+e68CpOmSjBYWmmhyLgGAh3EJY
b6F4xDWoo8cqXg8lDqbHQUd3+5DWjBeYLlmgay9cSQFcNAegnsgcGpDrDU2nMXLw
kxEqQLGMlu0Lc7L6Wr+SlizZ7psxA7KyDMP1bFyhb3xoeL6AvBe7xe9B7CF+xHq1
iSYkRh+UPa+mWtTKlms1UZb5Lt67K/x3pOsnpJEyFQh+b/ciASKPcznn74Zj00IZ
mmSZx709wydt/dLS7Lk5rF3EQJcKGHdqrdBw7lRYZtClm85ee72D/7jKWk0ksRpU
0jczZH+TYzG1oE0MFkpFsR1oyddVjmYEVMmbj+yep5fuwbREwkHYfiOD5om76QDQ
eBPKURXv2By15sR5Y6rg2l8TXjWk+kmYZb9DUV8mCLMVc42mlk0XzMXhjzjBCu4S
ifNlMLEid+CuVE3i8e5tQoJDenPIMKuXEAenZzf3UUZtw65igSlXkUE8SdQeTxzJ
3aCC6TWBr2vhGj1PmuydWC4rVg89ZbkZtoMYfaIxDizXCX/i0STUo2fmkbIhfM5w
AM1tlrS30Sa2d/ZuMqYw59L4XGjTJaI1jWr5THk00dbauqV6a//NRUGbIxpS4pXg
7WdWPrI8LvBo7Wl/LsHCAcglIpPUIR4wzL26VSa4anSVaEeO8hHxZDK1gBlNrUyw
vr5IrQmYWJRclhuKbZS8t1v2IviA862sbD8hdi5iF9nkQ0XQt2zxpISL3G/ZePHa
YOfWaT9keTcc2SKNcJDolDI912FL/utSE9S9CpNhbsj6WueAMv1ZNzhiYjFlf57C
q4YP/fdShPteJDh7o9w71sUtU7IbqUg/3bZWa4LX/ezcXRCcr8SbqC+bQYJR7oXW
L/IfqMK4niAbB5Zsv4rbVdi5kDkWfUN8lpMUrl1GPUFVtsImvpggTprvPh+KM9G0
o4o5IJMeFk717ImWyORjDNr8MWGTTAl6JwMg1883dda9la0dsHgJSSTVk82uv5C2
+NAioxGPgiLn8qZHh48Mne60H+h/cui2d5WV80djogHwzxhcrl0HLeFaoKJ222nS
Zzj5Kl10iw2u7tAJfEEfz7t2BY7KUzj53sPi3iAyJeFe52CBE+0E/PXw6P46ZGf9
M9SHAbmpLOmFUYrN+7jqqFTQG0w/hShDN+scMSpe2NFX3lrIvxnk4AcZnbLWbwM9
4MJmNF+DfxVB9+E93ef/BiZ5EubS2LQvn6JdsSSCdfRY4T9Iv/qcJjWherllyyj9
08c+lalbNZ5NGI8/tKstSxyO1HMgQ+m6XgVaVwDmo4vef28h+uElGTnDXqd2tx3W
qNofF18b8k9KJ13W/T0n4Uf7b3D9Z5eOb0s0uiKTKL0bLs9dcHg8abtQI2Fx4gBl
jagr5afVsR+MgUJqx8sqqlysUQ/a07nrmB0mmXKqLU3VPtVC+TzOPdBhEYWcc35H
Hr46ok13VWVdMthpv8Ob+2FOeDYRmFFXmoEAxPo13g885nnUNGuG76XT8lkBXjIU
zOtGTBgIqyDdBEtqSEBp0M4vGx10edT8bDvpUvI9Li53bAKGp8AokmMh9nyK3eRz
udBanJydUxLpCEtJi80zAOu0ZZiptRnhJorXFLRxZQBlVwMfUV7LnUzGJQZQubvv
7KFl4EUAjGK0gkFQqbt5Lai30vHNu8QzfiSqTVfnRVYb3r0FLp+Lt9nvo6TJWCRQ
dxFKDFXozPy9gh4vvouDTS8VFmaCFIKyudJsMFvctyWR7rehv6GnkW6rxVfnTh4j
jhQsiNfqSWMP1IBXmJxwnBhpD99HYcuiLUeU//ASMx2Ii21xVRG5Nr8oCPr9juOp
EZVVJ7evwBT9wK8sbW1RZvd7IfK/XP62ADLiC9Eu1CUBgpRD8gyPBtf2xP4tU4uz
Zsv8N8LABz+wefVtV490YwGEpmooDw/19eAYr4YzGr8bJY1R59OKopTxM9hWsnWW
LGdZBKT02R7iYCnRc3TgC6topRsgRwYJ9EzUzVgNgY+AOYH9J9iZoEdizCZrYBqS
zro2nvX9DiQ8HplzMwKY476U7wBuHgU6CDFMvfIVTElowyBKSOvnowkF2KxVHDcu
Pl2rVVmb17j6ARdCwP07gOprstj0zhD07NInoEDAfe5M460RNDD+XXgqDPv4uB2E
ZoOqZrxzzEpsr4WSXi2IAekws229FKRlI30rE/GfgwQF5hj+EDCdqLTg7TfRVxfr
u6BR6uhkWNfmYwr1gtultH1U8DoiXEY3IrEbmG1JrSV9QG1lV6OnNk41eLbyS/6Q
xfrfpN8/3hxVh22Mj6yjdC7cCDuX5tsXAqKcj9K3NqOhFVycut7B80jH54jMkxPJ
lhvO+TUP/JbMOMDqv2lhywZHFSuoHKeAhVF6SWuSVhQCwnGWAkgM7stxIKbFvPJO
GLvYNncx9ZH2ENXLow4OFwa8np/G5ltSdRllH50/2ot5segcdlE/Y0uiGXGzug9I
iGahYqsPnczGfgB/XZ/3k2kRUXi3BIH3j9ztEk3fwzBIQoD9mKsHgxj5WxExYpwu
AgjS4OgVCjjB/gaD2WyZrfR+C/1w4i4DE5zZ8Q6H1/62xlTcH/CApP3Wao+MA62T
B9NLAVJOCoQ1Ps2ZzDEBFBdQyOoolWu6F/pQFhrVr9jyL8FfVQzaeNuKzZeb3pne
ZoQVf0eTkuWjr6C93SuGOBUN1nO4+433I/fbsxgdl0WV7GReTPQxurv/L/z1d5OA
0CJP3hvkcjB5GRNO8aKlC63KaOzSCTr0IGOK3CmOtZG/4SXMwOI3i5WFzAraA7v7
tiGC8nVYbPAuxufFKjybZP/+Qdj+ckSnEWPXGUGn7MCnPrby0bBBjNDnibS1sY0k
a+YJWOtHZrNx3mT27v/qpymOHPv+BdhYpFOzbiQGlWkPSL1SZSx74B3zJH+/Ypvn
mpSd/a+oJy05lRvUYpajXewhKlQ0MOhMlU8776BSGbASSNu0NFnzjjWfLF+Rclh/
4V19ikfeUDD2e69MBotBdUw2QWs5RDorXGFI9vwVJFjFlKzSda1I+OeSBacfChyT
Ar+GTwqwHI1Fr4P3DY5RQtrHQ0nKHmqEJLMsXrIL+NYJ6SMEk0Wes8/uYIAdRhvw
grA1YM7ewAoF4oAFy9NHwK+cNm3HWjwTJk3QZ+C+72lXE6Q5zjoQ8VFduHOKtDpY
8RvZu5xhxbFaKCBrztBP4PHq2eBK7AogMJTMry5GIMC8zPoKIWhJ7tCDjNuetGeh
tDT2tbG7KDaeL4z0p7E6P++as0FhwcVf/0T7+AXVx69XA4OYoMFmpIKkMWQtfsM0
lKvskpLV7wJtdeSjKqKLQVUifeU1+UdkWdSTe0m75TyERgOQsn0GCj/AsXOf/QvD
LphZ0CXxR19JOjz4YF4sIOSLFHloQzZc8Pa5d4W1FW5fGl7UxtFirksa0tUOCLdz
uQ8Wwpxw7x55G7XLjHdA+YLGifAi682x2DNmfvnoEejf6rDA1VHZyB0qDgQH3BcL
ydRLvVmNrahvw1ftYsy+Ay/yNUMI6gKSOq1W3ZvGAE5fgXfLdQTf04L9jcuPOuAL
8qmIJdRA11AfybIIMFijwS1cZY3Wndr4Vge7jHexjuUxz764f7f9CzoO18Cdo3SK
makadi6T9RwAiojFUCvKk5vZ1bIM9vZFDa6/SQIhbXKF3OhzEHDvdSjrSvgu9wjN
0Ge5PirqLeqRm6vxZeU7Byi7u8Q3x9EneszC+JGmmfeUdfVDNWcYhAW8ze33AjGF
qaw3fxQZIiXNxFNMmhFIOA+0FUmXwsXg9KbJxDQb67ini0+UNkNMNn9LRzEQAyct
pK6JByuFGTvIYjtdDauTKDfv+lLixjmMtXLd6YyxxnAQ0kOs0K5ZJOH6LodFxEPn
IGey0ulnctF1PCLex6G+Z97wjoaWw0AbRREdAzxZj4S0/hHlO0KbRClBmyyvgLqG
F6CMkVRdfUmVSk9/uZQe1IXfuNJkS8ShpgVCuLn39SVu9NTSj/ayhpO/4rqPjBHA
2pWYzpQuUReEsAmWfo58WunPfBu+PrJD+IDTtdYWYozc6nHkP7bm6z4Iob9ENtQv
XYpwiOec7Sl10jqQaUXCaur0cGi864SXxF6hZHYgOXZVbawb6fb3Db44XtlYpYGm
bwQj5I5hLZJw+nphqz0TY80fEi6keFqVEnjs0pDD/8AXzjKtvrxSNE6FyPJy4jEj
aohSnz9Z7JEGhB+Z9AmmBPVGeaHOPxKvB8gCjMjP+W8JT6J2vYfh5T3yq6K27SvI
ocx+pZayxEsVBWrsHX1N/daWbD+eCi6sSoxPft0dtwqwSpc3+Xj5oeqd7XXUzETs
fpl7UqdWkGYO6VPAvZKYbYznDty1BuQL1RhvvekoK/oVaTITTwFfp79MVGnXf7zn
ujjMsUw5hAGcwzm7I2xhX7ZBtL/mA0fXe04dFDhmwLhX7TMqDxlfhP8p6ktBJcnx
zm2sS1G9uBu1l4TseKo6/SG6qCRZt7YbP2eCJxijaRpcJ1s7WNeYVVyb8Ov6NUbH
j15Mr/eCFQ/NUwzXTlsg7Ez8iD5NkMzU0VXcY7+p8gpQd0z7Sj/2DK/yB7B3bKe/
soOWFG15Fi6DNrhIbBfGIiyW2mw11aWTMFIuFz+zSQ5rl5m4q9yUftj1gHnE03YH
nqZpeE9OcdnG0E3J8iXJDu+qygo5k26QfVQo4I37NLCyFG2FqbEZ5cxZ9OSoN5oA
I5AQgpfu/1F4s97xvBW8H/7H3xFc6+Np9h09+wzHGnx8osvzm5eKz+tT854Az8EH
2L2bdRnkaj3slhwpkp0Gg45dmLZIs7XEdWJLZqB8JuuooFURPFrQkevr9Yacpm7n
KQKjt10glBOBfobEbAgevboI6dOaTXbEl8Ni4XsR5hPOPS0GM5YLqoUDVD7Ed/72
IvfkxtM6+jLRYCafLGQmTW8jbPEpTiLYnfnkAVzZmCDX8vRzBhl/b3QMm3QBbLjp
fljdZc2h/5nKQtb3JT2hWJCyTaPo6Notu8bcrnQDm+epJ/aA6jnKCNCuc9hIY2w/
1Ps86P9RPDxiF3xLTnCaycEEE//zHCHKa/O8bD7Bqc7lvb24BCx1bSm7EnBH74Q/
tL5MOV/iQ7qo9h/Ohr4NAu/Cf4jmsyBa32Ue5VpOVih6I7+9uhNcIrXgCvK+Aqqu
+rkLArGrmLas7O6Ep1DeVzrU6gdv2FKz0iVnhMQ622gpnl2glq/Blm4xLIHtYdeS
ooxFDefjgzhtPgjucFJVsmNsgMV7vZGAka6fBKxxxRGMgCqR7LHOlTcqr9atHmbX
H26MhYBbMkV1+PYl/n7k/JViZNOgWeZ9MBxc8Dapn3gfa7mj/DQInAxj1dcPpeq/
705YbvRAVEC4R2MO71BJ7iwZMOwwMwI0w99W/VV4AXr89L9vO1gxFhLCzVx8nDtX
ZU3y2/9sqBpWqbBmssrflUJvOFRjQsXYSWQ6h1QKSWKd3LgMy8bi9CnQ4JneycwC
SmBVjuvN0mBdVbbeesbr8UIYa3DTE6dDuBouuLo79X860rlNTn/xNFNVX5hLiq0t
wIwRK74BDBfotAuLT0iydbEa7YYu7AvFa+uEYvFJZvh2n1HY23on5fuaSfOD7UBq
yNcTfTlr81FQg1QRm3qY9vGTNJjRybZ6KN96YJZKip2lfTK3aydKNOCR6Fco9/tm
AJAdLx7XxJAuVcVBw7TVha/GGSIETTZF/jaj/1tgHASKg/+8+IZ1RLHmUWavUOfI
J+ihQwas9Ozi6h0hJKE5YQEyodsY9o5fIBRwbTjldGpdadux2tLpWrmJw1XrcZHD
dOaiW42hduQt7G1o1++xDG0pA1EgLuoRS5qpNyRA2G29AWjHna0g2ScgfNQKxcwd
Kir6mq3fkaq8FK62s18oQrRbmRp4dkSV02fysETEs3BtjVEN3WTCfSfaYqg2P+33
VcI0hhBdZbxIC86ovhtcqf8MNWmfHOobok+6dZ2VPXVWL8iCFmJCsSwT5bkY1fnW
smH7VxnPcIizFtS7wNTyNGN5h5TbJRRsnDkIqA9hmh/J3ts3ESwwWwcuNXj5VGje
n7W55TGZ2Ma8o4WHzvBoVBOvZn0ZMKaCSQU7wsQ8T5E//jP771s55W0LSlVfqqJb
x0Y4/jo2JRCAm+TT6zP5STLJSsPLKmAymO1fBobNzvjwx5RpHqVkXiUcBXmjSO/d
yzNoi7av95Xp0/GyssoRG/SXpn4oOxWUO2uRA5dvnoVv90lcsrjiwFU8dfk+p25B
qW6msDG7p7BtgwKfqwFZ44gSW8f1OquVQv5hrWu4cmsDgV7A0dKDinBSgqjCbG7+
zuP8H4QCRm1JrLwWqQJvLEE7FUKvZwK/f/AABopV2QEUpi6LD5zbK759qcslEgHl
cOphVzVXV3xK6cilAnoaaIAdEdgmhnuQnuVRMoHI0Py1+NZK7hMcPpPP7zM0+M3B
xt4fzuQ4MxS03lJBxd7uJUD9WOaiqCnS607pDxWSsxU8Fdg5kwh1T0aZ2mphTzWQ
3C/equG5YjVVEPTxDsKoSHL/GygtZrcPdEg8v2GosnSRFx3yGkny228UTkMC1DCR
NZ3PaCwLv2d5+/4v59ZxLbtUYuQj38CSpn8XImyuiNW0o4i/KP0qTBZuAR4hXGKR
m3mJoc6hAFP6DIqpUpkFsQicnMAuyRCNmnJq8nDhhKMmKwN0ByyH8Ks2L+leUZ5U
R+NtLY+uLMp247BHoPvT8STskyrga8a/FrbAmPcM84jsn0jpoIyNmqag9jk5B0QE
BxomFCO8Wzw+Ku1vJA19QBiIYK80KNs9Ski66RdxyhiXLqRS9uesq8Ytkw8qYJYS
dhnRhKia3IEPBPPSB1IcArrKBucQjeu4VdjRxRNBKhzf8B73me+EH3ld80TVnxvD
HfjjUMkhKfAr2iS6l3YOUb3aff6bybNlxHFFREPXRck9r+UC/TM7+gYbYoHcFPEy
JUUMQ8P0aPQBTjNRYVWjIlB2qXenyaChZUyRv2MW7/g0g+tq7feeAr0JyfVYExr8
MPey/dI+fsbgaqf8c7kHLdT97CpmGfSbUiu7WYn6qf6qkzEvD7LkcrpyH0spW94s
/onMjIYStidGNfBT9wwrKQoTh86bui/9RkjgUc7r2wH4SEBB8WuY5nz/xWfyVtLY
UV8GM4C0fMv6klO3nKPCZK6D9igQjF7ilgQD1pUZlp2ong2+UBM9FnO5+3gS0XMW
WmWlcRADE7MyWk4HpeYkhKHRUwha98YV5FO0LDsc+6spGfu+8w4yQhmS2zrpfxkA
uvv5ui25W+TJZFU/SnPM7m1EzU37weRgkfRatMzEPUBZaDH0Md7/ZsID3m8tU2W1
rbVqJ91+iw+9CV1e6EFZVBqQVZE6WzMIyIrhrmWM4x9rAXDQoCHeIwW3ajpLx4fG
Kv3+OercrLWcC/dkSRo0HQ6z/da+O4skGqMTzBCBU8iGbCpL8SMm2x8De8tGY6qy
S6+jTmn7inlVcNo5BuQI09MQVVRSgo6bNvlnfqqTUMslGGian5UXoEoYFrkOh9ow
lcn1y1INEbrzF0RgxnkZ8pIlPRVyI1ln+/TmMobwUk4WlH2eWcrEssi7EUE5EnsY
Ueub78dqtf0XKjyEf+CcahyELPwh7dsYpr4tcDed39XMxvSCL8WDubGecfEt/bbp
oIECRATv+QetoXMyZENL+a8ZZcUR+mxAgTx0x6S1Yi1KjxCcCADv6fVMfls9duyQ
KCmMi6F0A37i+HYgBol04mmYjz7VcIvzlwjLOjcWG144SYGpR2pTnTN8i71tb7b0
Ay/4vyAyAdfzDUxvJRpBbaEyh2rmSRVOPhuUtm/MTB/aXrzPXyb/k22W1ndvd99J
wqKt/KfohvIP1vOyYqRLK6OyGKBd9YRwJ37hz9qUgRtp32ep/9xPh/gSihywQDq9
UFAUG0PA0XtEOcJu5++AGpSp+79kyC78Z1SiNDoGSo7hYJl0fwBol6G7x/tMWEOP
tGeJUcjR5sfvXevJXkFzb+7Kqpcmd1Q4NcCuqqCE5B5pdhmU3RDOM8uGFK+jnV1c
g5C8whpTupvS1dg6l6C5FyArUnynKgSyEZuXKCFIwaQxfnffOAGMhAeQqO5oVnO/
jrVqvVsKXzZQGjfmfy3O1n9ZqYSIp6Xyl6/Dag8SloBJcQ3wTkKxMc9fPrFUfMBp
naT75FOTVGjKi/h0KhVlw0xaaTXt9CWW7g7TBbvwGkKEb5y4uo+Sj+VBZB0pHXz9
cy4tk7KXnAQ7pS/rdx+3rO1rhuu7IJhfBm8Op7bML1xX3P4wsYvcZSMVJ4Domras
0F/vZp4Yg6r0flaITPI4b1Fo5ddGQdZKbopH+uz8Bm6tUxZuUEvuKHHx+SQkeSAr
zl9gBuO6ydkwsWko7SIiIJCBHiokGNlvt9m0cZdtEigiXBpmH6xHhTdZaOgDT66M
WksexOWLj0olCcgiEgXS3mh7CjiKsRs+PZJzhnHe55CV4Jk/JBx8ei06NvWkfJ34
blP/uD4mbl8t/dsmq/ocK+ReXENl4/oYoMQxh6tMKaV3Ab3eslfFrH5SMI8lKGqu
SaTZGzPipCmsluCTcEziHR0cAJ0TSRamgk8KYEgL/r78LO8vyOW4b0nMEanLlLuK
C6CmhF3W2SVQykKr1ugmsIUb2SOu8P+6nOyH49kQSe58CGx3c1yOQUhIXC7Gpi05
GNhaw9LZmxcZMr5baLSMtcv5+wNiWy6z3EKedpYaCLkGWzKDzABgwgwwmM5eXSSF
C9X+zS2VUjI2Gjzv9xxoaSZyGKGmn/wxgTzxiVms+LkAJC8zD3VAzaHVAzkWyWnY
UHL/Hl1acmArpY9MXsa7kMgBSgHT6ukx6lQYBTJyUBR+gF9AMVndFFSKSkBdh9MU
AwcxUJ8YiZDjm22xN4rrQ1whlxnxR6s4Z/yqlobI05N4aumgc6nGSgxIApsDk7Bu
5T39YmluJHHcfpeyfckyzuxCL49Xqdk0zmp8/Vj552QDvPrjpU3W32BZ9ouzqFep
ZUqDrznuagiOs9FJVW1mIBtIUeuyKoUJpmEULgLwVD8ij3s7WKNMiw0wAO9d5f8D
TYWJcHAOILm5/SucyreQTCu0lFiZYwiS5LXql2dlFHMPtFK11tgRowR7FDUhSNQL
2jxzxraX0H3oXuGcaffOtHCIdNd8CHXdV5YiZXQe+NqWLsAHxiMxxQMgk0XRjrQF
HNSqG545+40TtQ7oqRuwrSOmYz2SorkxwB3E5J87wxfMV4GG2h92HSIO4FBvPq6l
YYXMfQWOHPpvLfzhW0NRkRoee0hDk5jFkj6qCYtlXmiwkylrLIy3lXsXOLAfbW6W
65vCeWi9Eu7JQsmOkMkPgjEBu13ScoGahbiqKrCPXlswS+dFGu4IbWgBREdvb/OY
WQNcI8qA/9xL3avh0acPRZnnOwnhIxuYLm14kriHamowTuoqPnwa8DfGlBWzfaAv
taSWvorM1t9hSda6HCOvHeUP2NnMxouyGh8NLOdljQBghP39OePw+Ck13t8mlgIx
MG7oBlwjK+f+PElw3Eh3aQMsjpCHNvW64RHlasozKqOt+St3pP0SRPZTA+Q5NTYM
tKQVz85ZF6bUosvMf7R6EB0MwaycAfVrQNH+QrhFX++vj/+MgSjM/OPiDppSnY0Z
QWIcLbM7tfulJ/0gJgYfUvd6q03ATjnA7lrUaNMJeh4M5kQdFWuL81ac9SReD6no
VYZRJhqpQDYIT4q+JbcPXfl0A8STtEGxDPUzIGYg6MRKgcsFxC1bkCf1w3yl9A3b
a7n6gumCc8fXYOWKiAvGWg7rLmRLqhSEG16hp/J5YKjxh2xJLszVmFKyGVc7xJbV
EaT/rsgtbzmnmw3XxfzJBY6nljVJLDLh0gYuW11jhhabg9tL/5KTzL/vUm4pULZa
+PvE9FxYvA+ZdBDBCKyICZX147l+ixXpWKgnTUh5O2WUsBFVZ8GhS/tyHhzQotrk
zjGipbNk6YQxLM2UrJJDg5uCZPxW3zzKsXydloscAuDBUAXTa78rw57lPXhkDrlX
hZqqbefKiJ2v4qsQBcdNCkU117zUodcSWSGd8CTw6mmMs0nAw4cKyuU9JYuEINSZ
l6MaCcozpACQHvvBUOWe2qNwaFOhBpk29pTETRkCVhdd/oMIUynG+OCNU58uA73n
JNemPjDtnRnETFCWzlCOsptJc571IRGWBvbiUQfuND59FvV2aB7/bUis0k25xnZ/
IHwxH84nufT4+Nm1ISA1n0VA9pNSrHXGfKQf+liKVVQmkp454O0mK5/g+zRbqgy0
qiqMkN1pOAznvgUyDlZRL9bjxehHDqlNh2NMbSBdlXIbjocHTM2YemFZTKmnb1OH
zr5fJnu1EiNK0UA6oycdXjxRL1lxqX2WGxCOznBJamNuXJELhN5r4Xz9AzSrZIBV
hyCMEP5EH9mUfeqzuRfRrwLlli596KLVszYj4ODK3Q8CHAH9dj8B9t2DF3nlP8Em
7Vy7WaaL9Dh/29TlYBPfqkrLc9wmFT8jEtK3bjoHiCyXF/ITHLZ/C5roBERzXEv9
NZW7HHAcVdvjCIRoFlYPP3+5pfWvQ6ycDIU8n8fXecE7VIL2T0RaCwsSsvWJrrtr
q0FQSoxE4j7Xg176ljl0JQcP6t78XS9zaGoI9tbC3Pl3w1NouMu20eD0CYd/w7iK
8JilFFq310yYv5Phx4kOYHf2L1lK/cbboS+jwY3BjBfbrm6BeG04Bg/4fiHTR8tV
9svtu573iucXFcNqTnGdg988QvPGbqdg/j98seTHazRzzYOxYv2R12G3Z2gehiRz
0Ai5DeJUT+HgbTX4DeLXyaF2wT/qFljTG15UC+FvcGpOBvqPXxsGYwbnWNqilGbB
+VOYlISib3a2/HFOEpIdJTVn0vjvnkW5+ZVNKKnUgT27bGL3XqIis5c4K8CCk3aM
t9/WVTuF+ZDB3YhLOYY8sG2QGCSrI5cc0VTEGdvHWP3XpUil21KRSSdbqLh5M2su
f2wUVhw6OAk3q3gbEw/B8h/X6BdXrgt3hWLA+NFtlh/jrK5zXtrt25Et/d3rO3t0
EKNGFV3me/1ybSBP0FKPx9WhvVDAhFhEspJejvhtXSBkpvp+XM3+Uf4Mto/tMuxf
BNckoQG2r093cel7bUu2c/mJfXitY1kQWAQ72aFn3ixOfzdJqcymRETWN0eJDami
lb1XAHFX1HcNa3OTgIdXIxa4dtzrUWN0Hy7q5KX2B9qqM8ESd6AFNLdPwkoPdmXI
shFZXrJhoaRBvIj7M4yY2MCLX3K9eKWgKSq4WPwNYTiC1nf5ANptBnMWFQOrmunm
9XXZ6PW9GluHrgx9++Rww4K25nZ7U6F6LvDWs720DeMc2mJAu3pMbSjexB6bExAF
nhjZnSe07u9rQuk7OUHwocOt7ZtYRtbfMgrPs7eorsxNX0dB6yAIdkpjW5cwJf1x
cXBRrHqQ38kzFATgjrcmNSvA4jQNJKLrg4g4VBmpUhZhakl0ErX1eK4rybwbL2fL
GqxKUjRh7DDBh9Qzbbt0YWtFU26d+O0GPoOV+SgKIPGeY7gQG5IITOW2kOMaTGia
YchBlv9Gcfi31tBqO193oANcr6lslXDQRFlxeeCbiW9h0RRkubBtomamrfX5+XWm
XviFseckXNy/p4AWIewCHMxTlJnYfelj350cZcN4h9TA6AQh392f8XSrfnDLaLH7
I2cbX4O19P0D178QpBO4oca2u+TbqnTWMnC9yjqO/+2z2eW2f8QIupTYdolgAfR4
2XSwMaU0z6HX3qC8ds/z5b7I0Yn8eh/O8D4s5GTA2wVEttB6pvxGjIM5oAAvJZnP
2xN8RELPv8OHHofIeF3p0EBdINyK88vHxVn5+al/muLzDP0GDmmLb5ZRMLhF91HY
jTbmEgrwnEDjaK9QjpoO7WsY1kX2eyuPwkav3YrdW6meqReXpP1UPURSJ63tks4v
HsCRX6XzT1O4goVYd8hv9q9ThZoORe8WCU2+J1UBh4oOvkQowXUr9N7THdAI7Dbr
KomDaBsFl7iNV3rN2JbU3vyvkEXDEXxnyLGI1ySOXW0v1F4tgxGrMWnv6apac6Kc
BR3Ea1JQUOmQYn5P9n5NqqGnFX4E8SKP7Dr0I8BPAys/LEvqgykAXsKNAKrTfmqx
XTMam14g9+hend5XLJ3IWpPag0SyD6l0geAwbre1VcVizyq0s4RlUgmhp7byRRPg
v0pqKc4sjW2Oh/malyJJpynaM431+qQh9IHhZ+qlQKEpwGjJy/xwkqDVAkcdPfyu
SGtcJ/6eyf3+ESr8Jda3G1ETOiwkJDOkYgSZINt5PvIcwLVkCevljhgFZZNneLkg
AvMdbo+qqh7ZJnhrW1afJzCURonhKANPrb8Ek2YS7tL2gsk/kDaSurwDQv0z+bmC
MCVsrYQr4SgVuo+MPU5xCV32UhlhIbiw5o6VjWa+M4yqtSbz3YQVmJDF8nWldu5i
8KxRdEcSL794KPl9VJ4b8yFKrgDmRJqsXKwQ3uYdZIvhql7R1B2GCvMogdFDn1Ze
azvcrren0G6yI2pKjqh6TqkwjTXl2PrxYRdj6TFX1JKHoQCq/Ty4HLKtMmUG7LYx
Q84mj++jODFRUX+rtaND05TWieQKM/IF0pIOX1kYe0axHKQTyrRBmv3DTpnw+pgA
KTbDv8UAmTra4FeFckJfDHYMm3Zdftbc8LHdXHNbLinKLPrkoQghhm2x6daOfheb
5f1nNAsu30VzwIS4sEoNXk2Aon887E12JBzIYyeEK3bk7UWU+zMN+J9QQmAX+ana
wEpxMNyBeYtWTcxeC2b06bxDizbPMmtebaY3hhaOMG9RC5wBU5uKmSTWSjulsIru
6h394Pzy2ILSI7cA1jNfF0zIa1kx/0Rs0S0hcS27Yd5Jtxian/nvjWaK1ByRykrq
ErrbMo4yqgDl25qKeVhSl8bjgl6SWzWuCB8oMwkC7yqPx0cRZ6P4Ge9VVLOQUFK5
qMWMSD13ceXm0VoQPu86+rEQzYBOaBzMGwy5xdIS7TwDdiye+N6O8TYaUPq7y0P0
eEOikLEspq9zsvEBc/+OXWXUbmv0jfkeyuYMqiaN2xCp0yJb5LoUbRyHHiZ4Luqn
Qm+7nJpDfPO1CWsiQPn4UKBie8LAdCby2r6pgx/6z+xMUx5DTp0Yqkaw+NUMbGnz
j7mdoaYhMxKxrrUKeu2erNOXr1wQ6PHH3/Oh+sSGdrP30YrH96vD1v3nvM0YojHy
IrwHnPJ0uLJB08/3lN2J/+pGD88PwCdbQTpbu2++/YkzDaSE4ajZKOwkNQNlA/MX
xsgUuHtV1NxtIbR2K12CVzbt2B9+UQpHi7TrwPvanGeWddu4egYkE3CL/l7f408A
J4n/uz2l6+5s0M+VV8UtPL5DDgoH3Cib3K0IbQqO3XTN9Crvu1vSXZQQJw9Q8Bad
PMSbih4iQQcQUQCMG4UuK1ktL8whM5P3LSLTaguD4Vd8LJ50LkVZKwn0vgb+ds3E
6uWpZS+gLGLDevkIxjzkoi0Mm1aXIDVlxqqBc42+RbK2wdo7KqqRdQkaOcRqcsRV
yCIS50w2/T5Rqih0G2yppW6YkprTWKALADPlZBijawFoobCdAbEZE3ii9OHHRJox
/NwkpuIsBeUBDYGXDYRnv+b/+ZPDC0QrYy3+Eh7jVPMJB3c5vcUT7evt+QKBtxGP
0s9PVsGovuZd+IFAdq06d/OGUwDkd2S11LjhY0qbOhySA3cpni+hB7x78JilG+l3
CEBpDUuE44PHHB+mGVHdfHoMtfiZyjYWbJukuuVG8gDob5rFw+glIZHf0acN1AhB
t6huhVGHAsbwtpAyJCyv1kTdoxsqwYqtOwZ8oRuZ6sDzYrbI2uLVjYIg32l0h7jR
uf6k6/crQnX7toA4ZU8bykHGrjD1CV1d0ZBCeD3H+MPY6HrkNrGKu8fvMNS0bxFB
s52aAwOvhgPEZJp1yVk11SOcKl0PinE+ujeTi84HgKtR1Jv735mjCYwVCC2zk6Fw
GwU/k/zzJKdHGHO18zwCc1KJjlqQahbmNjFT8WtfHv99jnkRq6QOCoKMageBHlCx
OmdIhKYoa20GhMWUbzZqFEdYAvjfYMcIK1I0RvZKAgppx0AG1QA/mhfyt0/0UQk/
yS8u6x09WRCGDBD1axCPqB5B2NhCK4SL9/xmZZN61ROpwOoEc6EARQsyojaDgJkd
UrJv7rCR0bU0JhpSR1RkD30f+0J107UDtr1bTAQlue0yq+HP+vHYPIuFhOmZfliV
eTSEk2KDic8g9/9Imxp6em+J7rQyTTdyGEXt368QhxWb/i80o7AI+JiUBQXV3l/U
73/8CNZ5yEX4ibCdh/fs3Wsb78Mf3bcLSL2zQzdRzQO4g1MyL5IcxA3zeaiyuKvb
vKUK+kYWSiIxEgHynLFGIq9/esd5FBewV2RqH40RAZbB5uMZSyzjH5O5bUjPyyar
AbuwO//iuvptgqPwADyLDS4ITx2xuUFyqINQ+LeGZjw099mxKgJd7RNVY9+YQ5av
HT4pBT2TwVfi0Pm6eHPzsU5K13aklhGwlC2iygwtX633xJNfHfEriv7ZcwNGzrz0
QNwAOuN8ESMlKzF63ag5CokN/2y301WNBX0w0TxjRKlTt+ririg6k3D2AnX3NikI
Q3gRbO3kMtoRpvgq5ELqxs3Uy7keDvsux+FsTnjiUPZXEpxe4ga6jMcRBuBRppC3
GtWKOR8KXawJe5NkuIEozs8ljX11lnH+PJa14gSJzpT6LIGAP8zPsDsgGN9XpSPb
wxI8Wmp9L3u0Fnu1zCk1Qbf+bSCIfEEWnrE09LGzdoehLJZ0jIBw8IoIampXZzKv
YYftlc3AxmUVPEGE8cdxEzNyvVWFklzp5WyGD1jPDdNeWKjrpYoouXysouJvB+Ok
uLThlXbO7HeJceRjb1n3NC4eEXFTpmuy51B5rCjyAwu0wDp5q2hSJQ/VUG9u3NkW
sPC2qm9CmNAL22e1cXMu2Sohr5sHMgyforOQ/JoVywUyeUzkHTfR71DnFN2HBIpN
93xL6dDci4NtbwhlvB0iPESs7fGzPAwMTUxrPUuqN7A2jiUlur+8C19ngQ5xhLJl
l2oSz9uJKMlBWt9DftkX0g2LvvFH8HXXMaJhGdeeSNYXjAnLLKJVauzdKKk336Wc
guKqZg1t0aXVNEHZfMnPtUfHsSDDakfG8Km9en0+VfPstJ9/n9yX3J5N5jRI59Ma
jO4CAHlA69Qhaa/k5oRH7DLSaMOv6esxFXb8f8WegJaYoOxlTqA5GEfNPVZMJg4F
k7Zs4mRiz0artKlhZfZ3FROdUvh+GJmb6EpWEqiiGlB7/8hzIb9IRUHMEidu65U+
XZh6+f5qcoNZ+bNe0W2dI9I8j165z+CO4HTqVPg0l/tZ6CW3POSY2t/OFIMHVI+Q
adnsykASRGhcoU4ayYzTTRM0IrwHJxp01aWy5qF9J4FFVyGdfd7gaY8xHBz3ZHjR
K1aJvNIfFZb4sSwUOAbrwVujSW9k0LotZz/pK+XzfZ8ORWhy1jQ1+rG8yGBj8Rxt
dB/xbrT/i3J8BneQdPbWhERchl9tvEnwHp3K69qICCDEG8WSv49psRCNgTcR9gQZ
Oq8sGeW2f4j12IrX5gj+AXPeC2BGKBUqYfiNapsAnpEPiylGmoNoAvrP1ewmqoj3
HKTeqwvScb6vqCKdsTKtd3eSpOhyvHgMC49wvLzv1XbXmgcWYEFOVKwhUqMHLYcv
KmMAqeYMus3XIP+SphKeQendR1JjULo+HW+Ko4s2Y7Nx6D6W+pOj2Js2nRf9WRtC
G450YTpGIG06eecTm+bAnn2CkoKVB0fXjVIxBHgqyOsmPsTm9RZxAIKKFuy7c+ni
YkcQA6UsMp8YtzGiYgcyUDaumSJB9N/CBTbrpZsy6UP8WZP5R0vV9q1fcAym8aKH
3UZZcFN5v606rUK0Bd8WRv3oqJ7TKX4dywGj9N8Hw11qVl+0Fkij/rvNUJoaM2lR
c848wO9ur3o7n9jGssnPZUws1/xJqOKt19moVLlGu6BhfShc3BPpcrKln9DyRE5A
Sl0v3j6xiQzFeBTOU+LdA93EAx4S2lTDChSSbeApbC47E3TUbRdgvRsL8l8RK2ll
neoRfoxpDEcUZwUNqym1jmqC7/Yczw4vX2cknm/IyWZOejsM/UQqQC63ShyPdVYV
NtBIETG0phj3nXvb7tcn/y55kkNjqfEujUAzmGYbpKlmtgJZ8KhtSH/7mmE0xZ/g
CxzCkZaG319mC+bK11DmmBqEcNaKPjf6NA9H6Qifoe86vdkUijbHxuOUu6TiYI0g
pvVCiGy3MAt2/dwLCfBaBVZWP6yDJdPyEyRe4FIL3ufBBOQuXvTnYJe3dEQoji5z
iLtLUWatZUYK7EbF78BmxZ9YIjGP7RnkvQwwxSUcfHryQ+QERVF5IjLAIjRKUUpT
G9pMCw2m5k3tNTs/ORxsSLGD0Ib/tE8njt/glUNcwUdZuohskWV4KRBv2C6qMmMG
T7fj62f5eyB8RO6IRMf+T2xDEt0XnhRoHhNuiULty/oin+T2VHl3AI6c7CCZm4Sc
45ZiHxdTGvB4ngBgH6JaBqZCzbYghPlBtWnhsJiu5oMafnQkhYnPC0/pm3SG1JLF
3Gk/q3Q1nnrATXVIFFbxSP58QAhZfKVzKRtXDFNduYmw11pDgQk7rZlUbhE+dODH
WiIaI4hXhyKB1ye0CA0tbNip61VYu5g/MMhs5mNudsroRDT/OzGFu0T1grGhfqQA
j3R6jWNiHLmrGDhkrQ6nUYWCAenUpIS0qHc8WJs1aeFmwxfxIWxoVvXdUcDPPW26
RY/j3JQlqrl4ao7ls2118yZ4Jzl4m3bUudfqkzcJGl0ByCrr4KN8m3hCj5DWBrXD
TL3tCWvPRWviTAsFy+XKsDj8LQrs9RnIrOGKaC26pu71HpQJi7yB7yTQtvZnTNGH
8WtIeaO4mCNr5IBc2z4T+ij9Mj5C6A73YCrmYGWD6DAL02pcQAH3sFLX/NzsMn7Z
VF7fM2tCaZ5PcUPh64aNpoV1P23eSS9hPg8nkEkQTiEGqHLHjNKjlCrJUVVE9478
V6PFJgjXRb5zdp/I6epZ3cSzBhQS5MgP8t/sLvewuYKvAliWhcAf15lSHgaa+XSp
RFitAcv0BtMpicL2HDnL3/XC6Ietz7WWKfWvULUDwhZK2W7LeyYUg+dC4oqfcnvo
Gbl47zcm1ZcPl/0lSYXZJpKLbuhXlka71cdu8I0BqkTLfKlEhvv6UKt/TbvhrFde
jlc+jqpotYoorQue1Aa6qFxbaoBgiNUWkk8yPckwgZMYHch1bi7mK/Puj+Jo8z3P
RTXh08uzkq9e+hffjZbF8vOa8mKvJ53rC9rY+IhRgzJcMelRu/lKLdElTQvehdPI
6YoSMUP9eQod1ILf6Un4F/qX6BnwV41a3d8MggFT3gVjBroctD2ePYzJygbIpZ+u
NTchuNVKO4wWF0q7H/Xx2z/u75vsI6OoXGXPEkmiGOo9Kwb4LhPB33COToOR91y3
1H0jQmWdPFDMeSwAIJyxBdjEGALkLqZdVFQL8bM/S/WB5Z6FAirTgCwdX6PhEzAH
Nc5OCZmQG57S+Yo0uxa90mk0z3M1g+zlaWofJ0H905szBV0nj1BmJHmretpQt8tU
sVdzeuCQijeADbLQKGpubelkVis/LZYfmUULpaeupZPp0PeV6kCuAIFP5FqwblkD
eQJ5gGGcuvb0MblOoQQd4QseySvyVcG8R9lfzfwkOxLpLO/TdZh4/atMEdqOpRX4
R4w+XLvkXE0xvNI0UbeZ6QXDEiEBR+yIDtH2oPdt+ZZFCJ2B5ofzArFQ9Ed00W68
T1CXqWV5gSNWLuVb2imqk/M6T2zgR1ZZIqbRu2Gq2IHpBb+mhNOFrq9Omuv7U5e6
A4nmAJIdDQ0FaR6iBz8Cs2bhI1nmTns2VBm8qdM8eZLF0tktiQJsguGbACPgQxeO
7trasQzB0qxNkEB47kECm0r3mmjvDf6l9BWt/ZEDrIbjKZM+kRsilgxGy4ySvzW6
HN/L2DVMpih8RU6ZR1y2wv1KCvktPHOegWLvhEEwH5QP8ckkAiSrveGu5xAFzpAW
w9RcJZas8uzN3J8k+hdBIzA9PwyJfLBs23jgll4Th5LEW+9/jZ5iz0ZcUBuXhakm
EoUx+/9Ewf4tESRkf88rH/bD5w6Gjwhw7bgRaFwOtxHI0p3tmq7Q1bBP167o7hHr
UOfHtJ/SHrQeYXLsDYfvO1S2sro2NdvQFZMy47ehK6f0glHzfY6/5iJUsF++SeOM
p4jtRICt7BVpe4ivSHvli6GJlKp382vCVTql0j9t8WB7ew7jJ+AdAfgSSkXEdD+5
OMECyOFnxYZtYNLXIGPvjvCohZn4vtZDP4UQ2OvBNxfOOnMNMWoc5dHCHmrTHRE3
GSHrR39mrZiq8MPrWh6nj4GNL/XOivRJl3A5miSlZayo55rSKr0w7D1yhy9U4zsG
s04eLIR0yLt1SsXF7KfMTmgHsmMbkaj+rd1vxFZ39fHRJtcIltxtMCdPBE56iqmx
ldC1TF48i4v3xSJ3bKTlYer1h5GgY2MYCzHG8YCrdvT9p8o6CesLB41a9G4pbn1F
55pOFgE4CODGkRODbQAon0kZWAb0XLWu/eai7lbIfI09UPGf52iywzh78247GToY
xe+pIGwxa7CpLyC8d5W7GubzOAp4TAVntiAWqe1xHtXLBvvCJvk2UdiMXEtxzzf7
tbV86ceNrogGcs/7jP7vcQJd9jJQWAi83/hEwGk9RWwyZ0tQDjAy54tu9eNKJy3i
R9VUrqI4dpH0XqZD+k8dnhj5CMdMYQz7Kw1Pa4FhJ/UujQ0F3854YVuVBdRasXWE
g8DiOHkkqs8mT0QyBHZ3n9eKqV9020bTPsyfoe1eBbBzA5xf2EmFQhGNxkMecopC
5G+60w+xTJ84keEwQF3WKLtQXAAFRiISvhCl3i1ra4TGGF6GKUVzzynIp1PwWZZ2
laKu4QV6Y7tB0lvTF54KNdBIlMfB7ZorYPeC7iic+UrbJMH2tkM70WIdxWxRwIBT
tFlZk16PP46m6N0BYHb4qcyJnFvJHLzZmWQDscHX6Z+ssjqjARbbmNZ5PvtyJDrB
4iravp0JGeuK2YF+s/FIRb+QSkeqMWJFy2rTIv3nSAAQeBNgmusgH8IVEgpds4a5
wkBaurg8ANGuNtUG4zOl3WDu1DwIRgnVya0mIhCK4P0txcJ+VSeBneBhpIEWCfEF
VSgjInjs5HNEqhcpzzpWfY9s2QILTc8dnHwAZI/l4HO9RhVczaAmAkYt2GZWhlpk
kTLRSauIlp7nPjklnHTXePSIILCSGGQgvDWPQWnvXNQPBJsJVWSy+ZHipne+5aig
OKQdI3ZF7E84bc1tcwSJZ5iwi4dw++O8OR3Kh4SujPHWMy0Qefu9WJhdirP0M6By
ICOqUNVnqzg/AMyKw9jmnlEsuZmR8q5iXD36TZQh23qAFp11RO90rzNLxXS3mhTj
B3YySSaHjU8AXrFaNaVpf98GqUL8/6+Xiuq9DysanBTy2w1foZipzswh10wk4sSt
PKl+RBqvcop7bz3UYIH6j4HRPebS2uyvb00W0gxlMdvkCRqRhJu5Ou5cIm7kVRyH
VmuTs2xNv3qqi2hybamBAcQWH+HJQVYdL218O2u1MFCnhlSip85Lz3//CUx2zumV
zqDBZUCondUy5xacE18uRBqmMQLZ4vrgNUt1JhTAfUs3+ioG34MHsQTY5bC/D7a+
Y1nTrWx5Gkj327zJqtebcIP/lbxEJTsRYZTeA3jqAo2LgtSv+qbEmrO5w5KULU9o
vvyqX1OEfgrj9h9W6+pp44VINahZ+O+WZruWcEIdB+qc1JIrlZMp5gt19t6WUnNi
r889UI38sk50XX7ySqYGzFKy4IzyNLn9Kk/hrZ/F96pEn2+VMOS9FFOGgaq376k0
GahjhOHhQOAJUHjGj81y7jIKVPsxJEjIrL1Re7EGkbmoQKfv2fb6tE66pX3FafQm
JlJEe5N0Mu2HBnF47RZnIuMaBAXhI/UDw9NftLw8PQ2SokOV7HDJVaTYSyXcBPCA
yYhpql7zzplvtaGRzdPPmCtWebh7U8EOE1ywOcwPNkPw38AA4hrTsY0tyECVdSBF
suupK4WgvOkkK7bP6CG8wBWiJQtZG8OHR0HgxOQXnTeuIWDsqDQ5l4YfQ/d9GKpp
pcoxb4v+noG5EGYLjD1CsyrJLZ1ufJJro4WwraAjIWS1Ij5ExyPpqFWbLhYCqAKL
gznJfqBFyogaGNkDSVvHz5msy6iLKCg3MN5CvQoBpPxP5wa8wKsJtJaBlxlkufcH
kD5z5F2FmjEOG8KnzzGJGL6A9vDm1ogWz6S70KyIImV8G83dMiK7HZ4hH9c8TDm4
38qZGhJDWPmcIlUyubPdxv8/9/XLA5GY8RNp/Jz2hz+hCvl5Di+Mw4p/BJjN4k0L
YbhEdVSoiEy6BmTzhX6wA6Kc0Zc3sh2JYgjnHusjkieiK+t5OhUb5NOxTf0gFtCI
7U0VQBdx8ebMsUuEjqHhc0q23wNMZ7JVpoOqNAznkv3fCMZ5sREFYz8LZPIsOn/Y
KQO/s3sHxD/SD2/RmDigLTS2XiFBKZxoMResJLG+8mKOeYAhbFbwQXAvpmwbefDy
AAj0nEdKG6pURxsApOWE//0Bb3yD6mx4/umv9Pp768zeQsj+6UxjUbn+oWoG6zm0
vIUg+ujdHJ1/XHHyD9EoonTrV0PXRER5zudTmxgU2h92QTMlrX03V8EqsfDxN+x/
S3N6y1SH2m6PX5dc1rDZic0vaZfKsPUy3GkY1NpfiKkjbyGwZmiUI6FE+X00JTWr
fDmNg43CGedIbnJ2AJ9fyQrUVXE1w3SB07hdDvnBc+vvXho+TupkAipK5ht6aLJ9
OKYu8ay48vHGyK0t8pmrX4z5OSvVQaHSJSa08qkglaPI3LhN7bAzWzTfdHQMO0PV
MwtSXluHRqEoh/MaIcvuf/sgNkJp+B0tOAmoaLe29NMzSEM0JjIqHm3y7xafEbeY
CyEWEAe+BzMbG5+1iLoDbdgxk+mbmrXJ4Rspz+zB5PovLnSZRqxft8FVvHFbHb1W
3qOUc1IPoTl0JYjXmwJ5Yv3oFB09Ttvf9qcDOV/8n6g11nDF96FjJ/j0SbzFTMSy
tDeTM407Gm5lCogwqIm6bucgXXkSi12zRWog3/oaAvv1dzuLng7+/oTD2YtVoZaz
XJpRud6t60zftn8f11q9Jvwwh2Zrt1j5Q6gq7xf9FK08T3J8FV/5sqgMHnQA4YbQ
nf45X73sUiRmTDiOIDqPnqkLz846an8ePKFi7Fw8LtMSffVZG2HsFmNxiVznhApU
jDBlpIsVV61PVvVZDCZR0p9FTiDKXKcFJrcydMUNP2/0C+iUaJ3kGzp1u7VCRpOX
3LKKbRXp5FTAPH89iJO81e9LWYi7u9K9CfrJSk5i5f9e4f04cwPs2d9Wp8P8BpL1
yHCEuKaS6WSCLgQRzKVNxRGmbIEQvwlvEzUsIKZbJ1WR+nnWTOpKvv916mcYVEk6
N6KwQLI1OqGPfQYlVfbHfX/w2zVa5UFKUkMvQ+WuQlzvR95SqWMwlvLSEBhI+Shu
QEtBX526Y3anFGQcNng82jd9gh8/N0mOlnOVuFEG5A7IW19/uLjADE6+d9yIy46N
BCy0f0V6V2Iqek2JmLLCmF6jL/2y1LnBZZBl4CCwn8V8CCf/OxDYv8axVnh5EiPB
b/XsrVKI4azweIZv841ie668I7JzwtxtQg6fhsO613R0LjaJqRpENGxKTMHI69BL
jnteRjtPg4IzqcE7jI3RukJSmpnV3lUIih7jbPEpvnB9Yvp9dXGY8+Jmjp5brCl/
tSqoldknpIz/bFrxHWrcxktpYbMm/sDYqzAhI7fkgcWsTzX85DTMHr7JW3jl/L7W
0KKvvU1NOX7Z9/pJ0ANfFK2/sCjsKy/5NSEJ+D21oIQNlLxlGdgBkr0f58RpoZb6
ynj4TSXUYZIcbdzvdKmIeOWG6LzJmykq6U1dQJ8+NvOdEuVLgvm38iRgRvHQ7JJ9
77dd8GVuKhC7IckitBniBQOpv1myEIn8LpuYSvnrGns2ZNDAwbJcj7iIAAdc5Ttn
3fgpfIu0fzEawgpdFeuDeaD2Z/mBeScLhfiNA6KhVYWhRPWlR0j0ua6vub1QjVD7
4JjiDzMnfvUKeOsH0MqheaR+yR7zudshGZ1WHxJhEMValcC+vqiB8yy7c+9djfNO
3mp1XYx5xmFcMw+IPD6VyRy//GR8pYNTOg0yRVrMf4FJWS3L4z6f/K6R0Usufr3O
w9F4l4wgQR9xKPYl6/XgbZyD1JZugeCjQ5ocQjNu38IWx3TqxfQsa1J9TgkWaPv2
5OfIMjX9fIs0FUTr2s58SBCfT/NXyJePTyfLnWRrVDs59G/PkNEdE15czVI8QT+G
OmfWa2Y0JZcN6pN+qEG67qel2xoc97mnuswk58I1bkUS/b3pW7+OX6Z5nRTsALst
X0NjRVbwTuj8D0P4h+1ZXjrw7ZoB2frf9iBUDvImVpa/WOT+rxJsiHkn//8IOq0D
IsP6wKwiBFXxirY/zjkiGuK3PLvZITM1zgJJVKCbuddtJW8K0Yb93PwSe4XW30Ld
ZduHz/VNeVcYElmdeFV1Dwi4aR7tcWMoRCaRHFLP5sk9VzMmBKYXKVIMmoI254Oh
v9kbebnND1NNDk5PvzPe4KziG1JeI2Bjiad4sUCKN6YiLo53Jx3ONXTMoCX1LjWq
zpOJU66TuYOL20EDq8gntFcNOW4at9iX9ancYaag/J9cJdoDZ7AWU0bj1PFWJQWe
WalpWyp4pS3b7MWVApKeLiTLq+iF7OolQfGJ4W7R2JGExWy7luZhnLJ+ZMptSbDh
o485eZ9q/xZzD7TAV5h/FraONG2AUUcYXl6ShEWTP56o6J/egai8ExgDpUgL/05b
0repyUgDHJ62L2ZLL29ZTMz/Bn/q3+r/rEyCyR08tWCDGZSnRMWlab6mSSTV7aRZ
r4u21P2o17G5YdrCh9T4kGjKbtv4cy2KWa4x0I9DIFB3LLa0Ma/xqwSwAO18PUVz
SmBWHSGjmcWfjXhjlcCRZ50Jd9+mkmVCvylw5RpBgkduSDTR0MffuByL/BDO1SYo
ahxo7rW1Icxioj1IkvuSNaXgtz3eVss9H4LvbeAuK9ESQBAoCZgk5oTYxTeiG/gF
QK+U+73+x1QZQCOgzTdUm7JJDRVLGtbVj3WvyN8XRR7z1IdfnDwLDRHn5PkLvDrA
wv9QLLlUJCzBkqPdtioeJANYjGAWZTw9EHmpvhSlpvSvw8jB5OkHcnCw5yxM/7SW
Fv1j0hfKTUzBwM/O6IzXCuEz0iCGCzjcqPP2NOB6/KJlKkUPkpGceQ6m01IL9Oh2
xU6qEc6sSRGYjL/QnbkE/CS3iM+yPzCZAfNsxn0w/WXRAQXI4BzNh0CAM9NfN+im
6QkHPoHtLnCS4+qHQdMQQ76u8oF5wP7utRM5kFKFlXkeSsep7JFPkXduQUg9n5g4
umePd6RPqKMJ23t3yLufXwmK4EAFAoql9mZtDz7nIC/253Aq64v5LVnBRShIIIGj
rVh0LAgq3+37e4EEdRDI/hRXnGsCMpTf7xgNKv20bXTKYz4pEkZvp7JaFtpJlZ3X
zwbxMxBmj38NIObRXvkKrkYFaf8bA7CkZKMRU0HOwwRJxlYJvcmYjYhv4XG3mIYJ
EE42EdYbyIXbAJbNC3mTVeYTIYaXEAc+M/u+BPdfbyJhLdyTV1sZ6b13Aat5/I4m
4bBYwdEjpgPVudP9CS2zye8PPkT5pKeoVogsPYK6IBYKqlONtbcEfZlc07D0rd+m
I+0ILl0ODiobr/rOn6I/juK7tmwc0IlTnixvoLlvqpYYARJVqP75eJUNwkUu7OVh
HsCyNCtuZVV556UpYIA99fjJWpVIunBhVeIrzkRY8pZm8H6kU+2RGlbr5RHh5fGD
jU23FHdqqRGQnDZ8vmbmC5QAECI0yCG0vWzo5mL+hBYePD5Fa/ToXfT/Jl3MsVI2
5js3sKkuZw5cKB5Wt/zHJfU4FPlyvwVgjK0itAVu+zyQtAVV9Y77Iv4kNWSz9M6R
/f+Xhmvgwxf5ymv1nejSiJn5PjyOFFXWoA3kBAuJNPkLViefzD8R0nK3K0yidKlS
6L9BrX7t6JKniUAJfExlVNCqtIv9obhBBzaJFnKTOzlhqfhBYC4viD0n12d2Kcey
qV4dHCptitzcolY//SRrKbklGrA97+1sBaH9pHQYhY9rejWS7AjrC6p3HvVp6wFX
Yyek9CvMAnjIO5LmMka2u2kgJ5WsJmYQyazJ5NS8ESs7antVCSF+pwJPhCAbYhwK
rsh/F8o+i6gaXtq7Mxcab97fJlCQrO1tazx4QwmiPLjbmZ6HmxWTvivbrQ6RAdPP
oNJp304h0c0G9cC5xsz+mIngbyha2ixB2Yrp4vqEkdjwF6IdrneLqRB5iVCXuD2X
bv7SniNX6yzAhyJQny7yKQmE27HMyOAzimt/ZBhuYsJbcznHieuB9YQ2tEsHShaA
w2Y60LlMYZ9LDsn/UBMSrPdMV4a3pWzg+7FEq16+JLuPBe++ZMFWBxPJvUn5RH2F
HlofRzeGIKJmYowgKVbL3fL6zin4UZxd5OrysnOd/Pyl0KhkCdPd/4y/d20PrD+G
ASJ0NOV62ZZLkSBnppMdJ4mZhjqQ7Ir1mAYpHWHzrTHThzbZ7H3DZ4FvAxjdxfRK
rGBK+hm5wRNU3rvGGSUZk7Gd790tH+cV52d5TNaLWJaDFM8lBB7aEEihOEo8X3d1
1MMPHTdKNTXtQO+8IL8iiMBVzzDQmlpZpNh6QkokCC74N1xs1Q8UlfOO3qFcRkU5
6qRHf+E/GjXVom0JkzRiULSqsoYAQ8HQxO0bTDvtOSdlnvVQlBRmH+60jLZcNaFh
ye8aNC495/s0C5EtgnZDsXZ1YasLZjR5bLa4T0k+tJMLCzaF5E5C+DF3jOSWauQO
uJADns4goGSxU18sNTBpve3zDKw633HwhAVQzov3Prx9pVO6nmwWUTA2EVCBtcOd
6fwBT3ePj0HgDTUryNGS5PwSTUjNPBex3q0TiYcqr5KqkfHuQHEEtkasPnfyUQDW
lj5p0jcE7l5CW7Yzcuxt/SD0UuWOwPTLCk9KJrsimQirm5YgZeBWkvUnrQpTm/6X
i6Zy+y3sj8M/iau81G236kQrUc+oWoreiJSSzujU/zw6wNE24zupXeXkxGypjHqq
yRTkftN+lb1dOOonbOZsp5K4Z5b+Ui9vxR1VIi57lPb02sfFfpLi0HgqelKX6Z+l
eyaU6O4P4/0FN7+EkXxbUUO92PqwGxzTLV5PQ0Q1LKzfrIed8/u8g4f7rCBB0MYS
RXiSEd+V0pLS3nq9zqcRaYVSl/e4q7dhcbwqxyopYx5KCMytQ9fKsopvNeorLntP
hfVMgOsYhxLuTNGyrBP4Ce+EOUAyZYzoN88m43fLoZYdJkOEiWQjgXLUGkEdsr09
U9FXflRfjqoTkgw6U9IjcVEnoPn7exzeQdwcfdDsthdfMnVaVMJ5FLkHi+DJ7m/7
UxvGe7h6eWFES3iwOX3m/7fBufYVUOtjEk18e8jmcNieUBsPBgdMbLe0+9UpEDVn
1avmU2wTgGid7IAXkzQI+e4vNJCJ89eeFmao9twTWbOBUshJnRxdGNvMELj740ar
SuK/ORdndqVVzkCXwNWrURB8RqgCkCT1mQZnFfVCYMaVqSqGeApIyp2PoQIOgb7M
U2RqYM+wKQsi5vJl69wyaUZCWhZBRXPVoR+dtzmnXREHMf/EpinasFLREYTb0pi5
YXJ0dATxQleq/LP5vGOrN3flUmun8a1z5NzP3sR0zM4/IqF6loPz7XrZ7BoZiv3/
Mu3n5fnPtF+mt33wc/zQ7TJqAXzLO7FDt3Rtx/BuYjjr4WC+a2H6Rs3vj6N7k2ue
geZZHWH024XOT8w/jSFRbRx7+8ZiFjUl1ZEpIKh9aDJjqCG4bV87m6YnSb4uxNCm
V0PJ3SDcdx2gQSO2XulYI+mRtL21mUlkQ0AylNUaxVIW2j/qwdLdglbdwDwYeHr6
cEmII+PHxPSMtHPF6uYouo6cmkYzyIkBvsaGgEKOkG7LwBmSgCqETzxK+ClmybNb
QwvkVI0HwpUdL/cYDfXTapMk/N371p4TfIJAAjFD4jXKlx4rIlVeEVzhfn6q4HA4
ASIZ0YR6ET89uL3vIwLxl0pZ0FMCvxaAgVPWTu01kbQsSyWK9xYgIIWbXpU63Aaw
l3hIoUs3XOgXbaA44b16eCfza2IrBiNLBI74DSAqRHs1+e1jO0cyB1/OaRGWvvB9
iO0wbXZJgYlxn9RuhGgVyAhz20Gn6HOfcBqM0dYJn6BptbTaneek0ODHDRv5JJW8
5IRbtzHs38yrs7D/WZXhxFcEULDx0neQM5iyHsw9vST9+yVwEF5YR55kEroLmjzl
FZalzLhniIfp9WtDxt0EZYc5yq5Sjo1Eg2JL9vBSlxDMwxKXJOWAlrthUp6JPj/P
rJz2JaXvS3qfWGDEFaZOv5CURj1OlU65CW/+IjLbIDI4gEwdLUBzPXpQFXYOM9L3
dVVhdjQK5z3BRGrTQ5qjezSnjxZHdeMXK95o1nXTYVt/ua76wT2SabJ/Pt4Y6wzV
axy1n2dMrbuuAeZt2h3xxHvxQIrSEa3MembrfBTXDgcIdYGy9edwo1urOK261R6l
61r73p99jPrLwplLNtEro43pZhVizD5G0jXUHN3nXy5o3u5h8gssbAPYdRprP9Uu
jrGCpOpfVAuRYHxrWZtk8uDdzF/1yn0lqvceluoF/2jqannIdIb4+Dz7C0zSqAtu
FZqhp83wr+Tkii3kB8u+pWV0G75cEY+JmuhgG2Geb6i/AqPmQPEe5/3ZnUrztQgS
HgSqz8Y5nIk+gBnSJJfAfxHXFMMLp0b50wVP5x3byUjbPa8ZNMkd1nVGhmTDLsLI
rEWjy0shJ8ZlaBSkqzWrevU7rjqxiuoUwz4MKCx4+Q7nO+uo3sjblW2LRLnCBJJJ
tDpDTB2N5a4BbDGdItaDuhMieZ5cqYMIkdXZTUwccSrYZGmo/SzvrudRG7Je8yA1
FN733MDM8XftnfczY1jk0hSI5gNZcqm8Tq/DR5vi51hQGJ1pcrDRluQ1d1G5mAVd
UaEiauU2/1m7yJB6ZSHOuCXgDozSUDRiAI0ooSwGU9f4fvrW0bw5m0OQ7PUfGXVI
s68Thws57+7M889EKYqNmlGjY/77kvIikWvSJ0WkDG7HXIBdFBD/Xtr/O/SN8z/6
SMuJJvflNFllsoA/S1A/t8Rb5V97v71mT6MI7gsqA/1Yddf7PtVdVF/CvXG+xdXv
KeCi1Sjrc09erhmESF9Gu2KydZ0HWcoM9Ekjqv72VWAaxx2yFrUrYS737dS6aGHS
m1AxYygb23bZIjzkHMJDEj6vFrEsq9UScqK4ZTQ6No6P/SjO8iRLDggCgm6zwi2V
Yu76/3Zs3htA1hzYYh0WHJKH7ndCZiNc53GovoGqcB1E7Mg90BEoziwRhS6bRhi5
dsUf4WvWcK2uoT/8joDSufWr1I8J3eSZBE9bP7i6tJS2rD3abdl+Nq4wJTc4JH0r
LAevaSGThthfpapyYRdkR7ismGM/KR2VE/yT3FZGSLg762T8d/0E3PwBNFF+PPaa
aZIKxfnxtsAEyH1qolmbzeWP4TodQvG6paFk3EwId+gTdrreYdRkDcwMeY5ax1j2
mtBMsWv48+EjcKpFcYAis+q1RtJyxV7PWW7NNZL7J1231+nwV+40pzgeZMFw4oIQ
OiNzC5pL2ahMmoK9zAT6y/S/cSDuGZUOpB/urRpOMz18DX2fg39sxY9DEBs0XRYM
jmLV4OtBpWp+8HtT9GuXhIR/Rq4UJBaybsd4URbJDGd9iHCLTw6vIrZ0Fpt5Eohc
QVrfrNUngPm8g+SJoQjk/pymh8scrxc/LEsAenql2TwVVUjwAYLGMajyHlICkfL+
VTFI47ZTuRuQ4syX8I7pIHieeApCwvNkOFZ7i400ly/JMleCp2rhZgNTmMxbg3LG
z4ZKOPIu1s43ESLJ0i50h/f8/dua6TH/4FK6wlLVdBBJxHNvX6FEiEPe8QrrR2T/
ChnIj7H/ZcTQU0G7gVpRjvTuSNpbNz55J0ooH3L8tdbn0w+xuDGTh4PNKRoc63T1
olsmdiB5MoO7Rd9o2PBI/VYO4iFbZO1BBKJQjmvnyYNCSLWFZyKj0AT7F4qTILWp
ibCQ8kyduoyWRXJnxUhm6WIOfBkWVMp7qYyk4454gPxWu+J3UAIkLUaHCBuS1WjT
BYWpuiiBFItbwTDAXhLLYVSjuR8jxLc0ii7qDIYIJ9C+S4p6rC1NuceD9HQIRKu9
Ez7TOedJqBY2BWshiHhwQaFwu8scdMtyLs+1NJgYhgdzIVhNx+0fggdf/VuFkSCn
U6g/KVqa7tufM7BmxRiryl4Go4PVW2Cdqprdcx7b9cuhP0EQajK0qqr0ljhb5bvq
Okrx0wW/5SIfiqCRBqTo7YnunwJhYFMUeflbg9BBTH76Xk2ioAyxp7Xj+JQ6+3CX
YwaUz2sQ2nYKbGs2wBTrFslMVLDpvbfDscS77eHebi4Vt6G3rd+Z7vY2T+dIv0Vr
S5k+qOhu3Yo7LWXUZVUfZqMZcZlJX3Dm43LfkLJMFAOn3m2T8vAttapIttAMNifZ
IEIcj/q1Zu8kHGngRb1rW+2w9QefR0Wt3FHO7v4rYRuzKSVlhZyhmDfRDIBCTVP+
80sirVzsZdMl3/FysAN/oPRuvi2vibz8Vwr1TyJCceZVllCjr5vPyGqx3kXAbkVt
CvmnM5NP7jLQxyvQP60reGw0fYWrDVgOxuwXvcaT8UppkqVrROTR/iv8JklLzT+9
RKB6K6nDYiC8qMbAfN4Z2jCOKiFwzVZfv5YKuDMwuBjQtOOS8VyhQEXe9eUVEFx8
jGd62f5z0kXbdMUPwZXVQKS7RBiXabx7wrMKHLAQBoY6mJ885aBHwsxNkxdulC3e
q0A/7GCa2mMBs7QVslkH/HEqKUPek9izQjRRDvOOfwEoD9Ak0wcFHDOy0CscmXaP
caG66ue3nmdY8VM/hOXI0XGlNrOwScjYfNP+QvzsstfVIp47mN9noJxxcx8sDE2y
CI1LqlnLUz7ik6fnakg+rOqoR+6exvOw3j/R7Wn57Pf+RrRyKPVVxj7usOUnNZE7
U/y0+BKDv2S4J2/aGD+Dax/NeZfXER71dT4tnFCXIMo+Bbx9qyRx3oqYMSwqhlt4
Jzll0T36xMbtCHenl2HlMaNmo+QL6pKI7QyARJK6wpA/hTERJz4q3RjTi8aFszdu
yvDwe5n+VeEyjgYrGOzjKoZorzGc+4xyxktlM6nEu0VnPeilSv0yS/hFDQFoUDeB
Dx6GBKKziN7KqeCXOmmcUs+OqA7ZEjRlX+G6K5EGtTPcXp8DzudiAcY7hZ23gqXc
N8TuEcFaDQmD3Qe9m91MOwBpLwW4hHI4T1xbzqrxYPh1ugr29NeJ7qUQzBcU3SkI
kQBeL55vfhMoXPrO2EwK9ETGkAsoeieOjAXybKPMPzY3oxLhlmu3QmNQcVrOFKUA
iyJ1S12pd0SrM5zBfRH337nTIxYEki57gO44u+RO49H06KfMC1An7q1v/rduiGJi
gF6zpjfMPkgbrsUGzhpk8GwI1Ot+6TwvLymMGl5grtZvwW0muhvxEBVBm2ucQYp/
BQjA+7gzSPCd1fAWvEj3aTJYeylaUbtQXPd5CV/3j1yodXcWqyMqVqYYsPf030hN
F09HxlFStshFWYAEVqBP4aP0jR4A25/7ePaOnLOsnrSRm52zgjTuJJ/kbYhZ2U4e
y+hRhUThTii/vvGwJ9HC6z5uGb1b+PICmfqWsf0tNdIoOe7Ms3Z1X08iVnEj65+f
bcDopW2SgI9xm0K2Whog6CZXpAtnBa2F3etaVHYhxGm1D6U/AFEXsDYdAikq+sUo
iHdKy2ln8t5V6Iyg62aAtQc3/hH9entZitqTR6gGyn/k8T9tyj5YKixRHxlzdoRT
pcMLC+U/rE5R6TdLOTDWhTgm8YgDzj9MHLMV6Eo0ndIgJjjCuddERYBXFwucp66g
nCFGI7Ykl4KoEOh9op+Vol6cXI1J0coRhgmPFsdKb2ZJmsAe1I9Znp4Dj6znU+Ao
KbEa4CQt+4rivVKcKq+YdBXgIhgQqP/lKALOx1hLgi1+EnQK5MHeyRELrOp18Uyd
Yc6KPjLgVOMRkCJeg8GRAerKrGr+dIjjBwPfCKrsbBcNadO9zMb1gUQS9j3Ac0gB
Nj72GjgnXElsKuyfKbmPNodAB8E9G3evoinCl+CC9frI5tawIVg3HEHQXTAQ1uHm
RaAFws2MPNrdqUcZKODYxSauD4j8FqMihi8B1DIcSlqrzJejYmY/bOo5bK0sf3ZZ
5upKSOOfv3pVEOFFfsSoSegEhXW2g/vePqRJVEoB5lYi1LMsfQQnvE3loxF6bDtX
x8xC67m01WRO7j13Kl9tOSjnb7365pnQCWG25Q+30ziV+gfna3/I/CLxQB7/MuF0
8hRIVtXSfWTYMZpGXp9YwXyoBFyR0ewyXfrqffmu8wsxjHMseZiD8X8BcEABk6Mn
KGds0rOSOPGuRKi9x39vc0G5/3tjo+gc/OO8E1x01X96/yxbRFHQ8+1iUnHpjyOg
5+XAr/LyUcfM5joYacLGTtx7ORarce0w2f8crNy4jYjkgRhAy0wP3yaNPA6bEwAg
AlEcp4lzPxInJZXbTUWPaUU0Op7FrHXZpG5OCDF34u3WWst+gS0E8qtVJvSSaxdR
9Tr4jbl4YRG1E2z/Spv0vmhbWLeIds8d9fCKark4wVDfXGFL31gqCUMOz2NYNSXf
3qzfFDvf67Mg8bJlVsLTvNvJFTOvJ0nhNqvsHZ1M2eg5fA6WCS6J+pcMxu5Z9Rjo
rW09DWg7bFWTIWTPni7GtCVGQd3oP8NohgbKedFpLWfYAokbEGEEiwq+5rnOUMnO
yU5+QQHPNC7rTT94qBQB3Igq5f50/GOHbF1IMEpOubTw32/hHF8DpqYdRsPZtdL4
7akCpXxRAkVXTKbZrh4l+/vZ05L/sNOhr5L0VsG0JcuhN6MsjA08rBAIh4nXJY5o
hENgMUo7FalBQJC1Re+dV8YkcOe8rjgL/SvZCMzBQxHsah4ZFbfjWgWM9pgdpJIw
dOQTKw/6Rf58Cqs2ULLm0ymn5sYpK/ivAcUb5lxLyCVuOUNFrDZYOL7XNF6yOSjl
c/djTJFinAKEkAw4yBvBIWbzkyZUmgfW/HUKJm7gYo4NZ+VsshRNtLEUfSgjk9eJ
ZGc7VdmX9aKn1rwuDAhrNdV2jcoEUQw+AbmNI3ohl0zslhwrpZvngFIEMIZqvtvp
Cz9wP+ipSD0HlWEAdznZqkIPXMOwJbWBHgPxBLVg8W+N+arVMCGciLVfc7u7Mw4G
NiRSCTPFWlV/SaNqCgUfAR/NjYhBx4Vi8k3GCZYxLAsyCVVtXaIYU8THg2Z8UDEc
TEP7l7lO33RlVQEU+k3sKPuY4/4o51Cm+ObDXeeOKPY11kW51eL1RP7Qtl/+VNua
QcKZa1ZU71FKbVkDeYdjcAC1gWiof+bwXOxTolenIRnaN3UOmZEAyYDMqqBE1nAF
de13hDFYWfqNzoxbqPcfE1T0SH+yxsRsb7wk3esVyBBqVtQK+NKUdKdTUkCa+eqW
x41V+CoczqATAtXgTCCo8k7/Oxr0sKYQRUbNWS65Lqx8WcS6nd77A0rZYGKvSJ0k
aTfle8GMwn2syUMzWj/LqysWx53DLKju5McVUO2q3GAshmvrKPw4mbPiv6tr6V6m
cipWPPlpeAxN3FcJCA9t+NhoDacLKd+Zvav7Owg2cDp/Orc1cmfhVK3VcV1b38fI
G/WfHT2uaFFjOUEeLsVetkGuIzaFXUAE8AXbVZhmoSX1017ISknUVIuCn+cKJkRA
8rhryzYMGLi5ezGN1dN9LJuVGWo+c+IuJUsiD9xKUgsfFZWCwle8bYyH6atniZgH
GC6XzU7+ecK5LqMK1n5TWuY37etmiX+VrxAWBSZS/78oL8wfhkdF6ScURNwoC7Y5
htgPZGYESXc06kFeBfDbJPiMFniu9aW2y2Dp9ob3oFm430f8cAJlCI85viczB7Yg
u10mPTxkGmV2RgMrvQ6xknRk9oCo1KFT24/A6W6U2+7jyKXnXhLARdm91OAWMUdv
4hhu2IzBMogN1C9hKcoEmeKP+bh71jvsOH2Pgm7oPH9KzHoWw43v/2nyvsKiagLC
fDqFPQRJ2p3tKdmj5+Kbk/oQ3mM/MuUc1Y0R76s+YI7oSDiS17yUrfDk3glPq7HR
/9i4zlblepCT577YgCYTRRKmYp/Ny6Thyapzb3yv6oiWbu2Wovh8jyulHGPnBUb+
dHyRWn8Mi4iypM4qnZhVv8+nNFdHSvVBTgH7xoLluor7RH54UqkurNBdzGs1VY0Q
9NBJkivd8YDGDGJLrw91o8YCi4+O1tZdSyoKDkjD99lyz5k0V9bEEe8UQTeNTaeb
V0Y2oI1HTmbLezxqDzLKUm0ZuRqWkoW4EgPe56HAUNy2Gtq/PVFyLou8cA9Z/5uC
67WuQpM9mBZR5FLdYXUbST6a/zkk4NgYqWJSNVsuijMfFGxOu19LY5TfxM2u6EFo
zxYBmSDDRDHxLWzxzISzff/ZPAr3A4lSFatiL55D8dU4mXuUTS3tdVfLd5vAFdLp
QyTW0RoF3afMUdkAclffaBJ4dAz4gJs2WS09J84hX576IuUPkfrLJm6YY17zxmbs
uoVqWpRdDaabXZ+zqhCf5oMjJFylTpot433k8f9JHgIP0lPVDulSflp70Zt3Wayi
Iqo5GnsgBeDEJdB6YnY58kA0hDi4DQzM6iRwK/6JcdFCkdO8r57swze4XBRTtG9R
OHU9DBvaDdZjYZ0Lzrqy9Xtng4YhPovjMiT2nmxhKkItdiBr7yowKVZtim9T0LSt
3LiC5c+CAqI4uoAS7CkGdiZpjSmgj7d6Lyh7smcqPh+MXQfbAYoe/BLZyA6ObKt1
4JeyrkY+XGul7AVkyzJqJ/3dPPuFcAVNd5/peC4NFW9/1kXeKKn+rwR1Rztv0Yal
gUxn+q0m5MKU8XkNsDoCyXnCtZuio6U9xOAmkcjeQUV4HJa4dtQqILHbUmADZ4rL
kuQe7wD/s+oOfnVaEwtWj47E5wniZnXp1oSepRucQs0JV6eJDIE3uG1/Gi+aZiCa
Lrqos8r5OfQqIBo4Wd3TIp0TnH6MujU1Ft+7zqI9h70GkAh7zQGLNXVccTc5o5jE
HeKm+mUi9V9JVQYdYwDT3W5BRClTmkZUKaz+ZHaH3oGtTPzC9NjsHuCaV0SqgwoI
DP1kkTYkmecUQAmoDJdhIJAeU03MDSQLEKxOEJgxBanbmzZmQp5xoK7I2nr35LkQ
x50NPHQoGAVTDOPbQGCilDWOofShvKuUw8BKjq7e+OyRY+XXqzM+GM11RjDUO1qC
0/jsCEy/M4QzdWLOJe2gBSmhfrsFQGwyW3JkqIImNexwQTn7HMCn1PSB615knxQH
fGztTIHbUQAm9NACwMxkE+2iq3oIGuUqtZNBiWZaWFy5JyizBulnkoYtrEBD7WbF
qHMogWJW5rmHTHetIixW53DD59qOVoCbQ7XnycTf0EhURKycUUCscuwfX3wBfizr
CO28hU14ex0m/WecX2tp6ORWIt2GhrLwsQEzFiUaAhfuA8RL578hzF3IPyg5VmMH
7/zn5OOVMIch3zptbRy7mxlweVrr5flfOtA4AZbYBav3ZKKf15dM7juz4YlGxzOM
wrjM9EFyrMbC2alI4psuQBEGefK8nFG0EYeJnAiCLRRYJcaXY2Lm3cT+Xaes0BUY
UiUoU7B96uK/YJ1Jt9f07sXUSrgM9cvc53tI+8NfsA7oIqNJOxMlayHp1sSwUdXu
ARdXphehccBMQNHkoxADpb57Hdo4FY1XG+COgx1YVILlEcBZUa9LLWr3DnKX7swq
b+mHoFkwFAT9uZrj7KWYHkcpYR2/9Oi+7EMSY8Uo5TAMavCyLy3OtedmFVLPryVY
VDH91y6FGnTjiHOLXnezuYV7z1CCxKBkP+AtEz1J5ciSQ51VQa7Ljw0TCRHJSkDw
G4quPc6+7hrmM+fDNNkTBDUSv4NKlCtDjeKkezWUHjIQVPjKSAQHF7Olqh1ddexg
H8ZmJznE6n4e20AS0AfXDDJ9sdTuHzzRpWjey5udsipki0Hikef9eTm06XtNM/z+
rtCOSpA/mr2AcsD9h5NJW8xzsSbo5iI8VLCSEnJ9ch5j/OoYdTgCVhvkbxJeo8p7
aZJxrNVdTBzJozfVXSOkBOapSR1g3T0xhxP8iDN8dB8bDXWOIQ3RPLmXRMBs+0er
8ThhwFp2rCI1lN8yHXD3Qu8x+ohs4INa0Mj3u0+6ErF32txBfnYd6sdsMxD6GS5w
f5R3MYW/KunccNMU0kNJUglHFP8C0RPvZdiuxfVX2xoy8DDwYeqAaMvtPXOrDYWU
rF75PSY/CwtIvLeEcEr79+zVZVcpKfVOqQBxL63eyOEBJfh6hGWjM/xv3LmoefSs
jJWmzHq7aSo5onF95LWZ/u3FOjoi+J49ZQXvrZRpdtIHMMrOz4uZMS9XfqehHtd3
wRtX1HWRTJPz5n3HTNAcQcIsXdz55eMDZGgq6lLf48z5ZzJJxUMPwO//kmXtFCK4
J0AmqnalFwjDYuwo/un9IQSQHTmOhB74FFFQGGUxLR5b+zS3KovXiW0SI0grO9Up
RYBn0nqg4RSAEsZ/As8cfYwuFf7r57GBS6VaBaWEsaP6uHHdFR975QDWKG52TRLb
8jZM050a1u0cAnrNvMDrqkCeiweaFL3ZuAP3YOpe7YzatOmDp3qjBqzZ/9SRLc1t
PB8VURPOTKKPnv/EVkV++oaEFOlQUmBnPI7UrbA2WS3CTRs3WEBw3e7tmfGhjh4e
Fs5WDVUviNMRGOaPYr+m9It8PNo3AJvDnJwRjXaFzoXMpax7aqEKwR+ZepxUkhjD
tTWHY0lyMBlM13UOp1QoQ7JIKbUpxcW3sCgoctwS9XL6j2mjnmG9cMyHIp9ZjnLg
K+hTTcTnLPGqpUTUCKiP/RDfXkKmK74YFynQECkR1XNcuvrPRrJ/7YT5icae5SJf
cKAXNYzFRahlGFNe/2PaGNmUm+73kM8vYqxatb8bdk0vl6vBNROXPF7MaEtQOlwl
hbf/HOCyqHiMw05QRN9WlVFAIk5IboZtj905l2aC1IVlDCKrf0kcZOmXrOt4FhKn
npGvA9dDVExb3Tb7eEXBV8GeexEJtCRjpDLdP+G8cAsrRVPezBJhIbCpm5WY4BVO
/UyJcPvYIDfzShvQGks5tlKvG7VcaZ47gNog+KByGj/cLhaWe0Dr0rFn8BMahnVJ
eiGYJPrD0zgM6udWuQMifR8sYz1SMWTfuuqefJhzAWiUX+6eblnI0q0nzpUaf2Id
n9CajUwA7KuibHSXCS66mw6s0m3ah6dIE5g9JscUTCOnb0B8WaSROhrpMlUHmVPu
5MDfb5sKzU9PT5VwrdTSx+3N+CBHNvL03fgrrdxlikhgtBFd36GWJbCaE60CmgL2
/WAcGUnkp4HKRE9gn8b925KpsXYHjC6oxGNcAKRkUmAtORy1Z7Hm/8r+BjHQnRoR
R+Fhn58YCwlaj8NKZPsXqsEyMtFW9SkyID4YgcUxFlBKEIbfWnOdc1wM03paP4L6
JacmISqNS9VNtFAFbeznC2pgfQEd4e+ojZGhyhRVNSejloeG0qnj+hsZ3+syXdOD
1TUFsZ31rZd1Kc78x6t247CvxRnDrCseTvaKYitSpclx//VeNbyXTbqPFKfhspWg
J3rbyJLo0e4ABRvHpmQ+k2p5pDtoweHl4qur0M4RCkReAZ59r8pSU2DxDRupauXG
QI8NYpSpJKOJurICjhE5B/mxzIiM2eHrpVG/bNjngB9lTazRe2/DG51bSfhKp1Bf
PHbwplG/rzQqT7Z3ED8PTP7mTNQ3gwOE2zioOkiTXN2KiufKFX74qA90udaYX9xZ
pSkCGsmDn2ZbelfiEJlJYOetxLVtMxc4dCR4983fvGk1Vv23g9aBIrdl9NXmBO47
cL5PMjRHhydzBXHSTViBbjs8pd4Xoo+GI4E8auRq/ghecJlKAP63WtY8tUoHWwDQ
RL61eU3ksWf9DI9PjjM7Zdr4YFc7IwwR76fNi1kKhDof/3+WN5uSGaOOWblJ+f5+
dt991PH7q1EsCzJtIG27YUwrAkmocP/sRTa7tVB32FlFwLEOKX2Vo0PA/wf6zgab
kdOhfgqMheSGCeYVt6ov49l79s1NLdUnnMlZa4NT4kKgwk7gB9UWuGaWd4yuYFkT
EsJGRGYxWXLRMnuCLY9tt6qlI8KkRt6N2H3xDd52/n240YUfnPJmo5DxV3cJLtv9
pY9pQjmoD2sGsEpijgXAywPgxMK5+zVWo8sGMr0+81IYozF2XwrgSg/i6/YBvgFc
2yqTJgU5WR2uUezPfSNk6AZ2DcEO5tzCnf6XOQ3J77ZRjFoCnauCawMJkdDBjGN5
o9/VGNiV1GttdALBHBSygb44DZiPGQCllnxX0rPnO9yTzK7NXWFfjK7gLq1PE/vc
PVVeABYs97IsHgy2F0cglkkkVRnFEDE03kWV8qUBf9AFDAb3HKXDEMx+Ie29K8Dj
9Oq1Ctz/GGItxGg5FR7HkqoTzs58VKYEqtUO6BKvrNGyOU4k11R9jtEedZYczPbl
1ZnvtvnV9Nwagx1fzGowtXwlt2uwl8BdrTe1FRTFv/OcJ8AikroDl1SxEBiIHTgb
PvVvCg9Xoq+j/+4OQUAitLWp5KEcG5JL/dEv1OEMNoAVGmmtQL6BfG9Zwsp752ZP
nRucogRAetnIG6TGBbiE4pQEnCGcOch8Gk3Y0Ya+rUi1ne1a3uQNsFv+llMjYI+c
/p/hKpiFFGtkShp2Atb+X3uOC3XAMqZMVDVXc0AC92BlfRovYg4f99QR+C+Embm0
p1MWM+v3Tj90zWh8lpASNMuEvkRVvb1XyxF+beSp+Voy7RQCZrBObKv7gukV+txc
7eu2DWY7+Y9aY/g+q3s0OOujMrFhPWDofpIYksnbjNjg5glA8G9DdCQpS9o6dpU6
MGQuYtbIrDC5BYg3mowNfZnxH4HAfJIkwZqp1XMYYV121CwDV6C5rE0gSZ+DyXST
1KxbrP9q7bf8TcRLSg0Lw7BSTHqh1ydvjkSPrZa1bnN1gZg8+J/Qxw0ONN5RwFfj
yrq0uuUmc3plPfTfehnSg8YbonWKU6k3t2kzV9G/FAS+Cu894/fNzqIIV7vZY3Og
WtICuDwX3YaPgd5KeqxRh4PjTu3EsetpsZIx/1CdmWxl0RdkU+RPOgbsSzdPzvAK
hIsVZU9Z6k7J9hj1aLTOpQnRxF56SlbSQRysqbnj9eLcxc/JuVWwnLjIdD5Pq54q
spde0aYHz7OOkzPMIQN193fh66W0oLvrTv4TLTS68B7yIVtD1RrRWFs5s2UhLyxV
ohi5wxea9o3eypTxTw2n4YDgt/iMjMDMiKAypWrEafGDTIxgblf24AvBQjHXiIxL
QtfcHsPOZCqnAgHHex8rZlJ/95pwImGN0MkpnjNoM2RMp9y63WqOk3Of5smOqegB
FqfuBejyWwxblBKI293r4ZSE065NSnzYetJDWMkpDjDaKbU04Cmh477iT4muyz1m
8c/Ri4hTeJ0QR2yWv8RvevYH72CtCeoZV1pdHxmmTErDzr1wF0PVOVbvDWdsqf/V
iY1iIYpaioHMxGDvZBoPcmH7Jid+hlB/VHGvjW8LlV9H3CdD4lQ1R2BNUO/x2o10
cR/WFIkxjZe9+q5CC4jGnZLo2+QmGplsQfSMjZ8bOkr9OQbJbk4bQllriueZfWgi
TXWjUMcESmwY5LpZ0JZZuKfXUyuf/nvLaI4csl37Mpck2uHyPDcziBMxai9qiHng
pK/G4mcThszSuvgaraN3es9ih7XTJfjQ4mWYUaaKzgQYpFVRQl4i68LjnzQv9hEA
zOtGe25V7FjbcoHcyRZZS6BVk8906FPjAWMKs3o2IokeRw8yn11odEUCHp/p5IRc
4HuCrpaFcq7TWdzFZ8ZSvqNDicTKV1kVHCcqfazEXrK72JKCW0j0IjEdfqdIhNTj
8jW8+YacP89EgQ5z5qiV4jprg5u/k2zkqA81Aw9uw0+XXqfP7KajtU4JV+gw7tzk
LZE3dvsuNQ7C3pl4pbez3SLGXztv9X1Ce7qvxZwncLtd85tf6ID1v1G6nDtkFqcc
0xhgxQllrp6BxCotVc8/McKP/YqAgLLCROtZPBTwvxcKjjqVj1xRWEUy/46AbUnM
55lyHTk014UTU11HqOcMlSQBC8TZpaAa1s5AJw2qLkCFpQxhNw0Avq630P0xweVq
5R4oLRa6laxKYs7DYLn3bOoBfRf/tVLkQkZQ/a13jSqto40DaUMAkXkFy794OAQc
SuPnphUI/4hXlGD4pX5eI2OwgNG9gxm/DjKH7zJ6a7jWT+z853fulnZ5ogi4kn78
JprqaMl0qVTjBjrA2Bzld7w5hkVMVijwv02vCm1ZXBaS8Zf3b7IkILWkeWRmonqF
/Lw389U5a82r2TT83w/M7h6mlv9SVgzTfFMCFuO3YQA0kYfSOx4PlW7+qrVxnMPe
/yo76fkIfUpEnYsaRVAmzlpvcI6jRwL1vUKZ92EOPjpFEezJDNhipyD7DVW5iVuz
I68H7EbrxtZ8vPzZbsAicFPYBBA4O0bJLlzT9uEmh4LcMp2vCoYS2XReiciahET9
n5dplRPTKx7Qcx3itG3H4qGH+Z+O+cHbzh8yP8kKPDlW76iSS6CEhgAohUHOX7C4
YBUADmF31CXirh9YGFZ0K1/OSf+20DAaJfRGS80ZCbdxjUGvu0+wXymhSsrJpWXB
oHToxWMvGnmIgsBusPhxpmugyuMpB1GqrOLNqF6Mk/oGAkvwWIClClROwhsM0esW
UQTTPuwZf18woFqK2m5/lmd+gEZ1a4l7w/Il32VX4go6mqv+XOPqVu+iInlBd6+I
6WRWW5jtu4pBKHEZk1sDo8S9BqLZLAlKJ6JxzA3iF9/f+u/PCie+Gh5qeScBj18i
pnpy9pV85ut6RQ7OzijKgdDMSbNAOz3rRmrh2y+igNH42x5TGp2aCqcH0wG/b0WN
03EhBb3wpB4iA92ghhw+FReUgxBjhtT5Rmol+DLjmEZmU3pe7V6jBEn1iLQAEl+m
ZIjvpFa0TkPv87OM6fN8gZlIATJqYIFprRO2RlI26+UppjqlWwJpDCT2Rc07warh
v9FAltcT+oVNvctqTbRfqnfhYC/HvI5p5zXEyoGJE109/bh4AjzGmy8IDjzEe2DL
ysDnUZUUqfPHm5S9ks49ECB20Dxg/XPgyjI2QZRMBwYVWoM2N7OrcqTf8D9ZYYBX
fjAgcaZGB8ZUwGvtVzlxTpXlFfDYma3stDpzRp1mx4elKdSTas3YEb1pjsSl3xrD
An1Pdi+VYrZ/P0us6n0I22jpB/cqZe6HPnTDvagLll3OvbeItclwTcL8gkv7DoGb
eLf9DklmSaxo8aA7OCVgheoFAHi3DUWpg0n9t7ArURi0qvDVVTZU9uToVpsyxm2y
tKI94mtn4GFy+niViVeVjUj6hepraFBGLNGX8u2Zkcbay2JN79MIQs87BSuRavd+
gj1YkZGSueMvz9gefIC08fyDbA/atQDkCM8HGuYh+T7RqKEu3sKpiJ3d8OLHEFZc
BQ2ai2aNE8lkMrXYwsTTO+2woRfghd1gOcBY/jJbvE/f1ApskcZzwgFE9GvH90qd
p05aXzLtJlLR1WiY/HFXY6IzmHq5eCx+xIWAzNVxEl4uqK75XbRm8xNvRN46aKbm
XpcWTYZG2DvDTW1nhAUiWhWlsDP/Hnu22BlNeU4abooYOAZYXhknHufbqY6o66qP
jOyHnOwede08LK0av/Jmvz+Y4ovA4e/pfeJll59eIhbagNLzkGP6e8n52FVacP0L
8QceVmUMhdDdj+8z99ybo/1q5iJsnAqk0en+XgVO1WxLmD0RAiHXqTxv4Pd+5a/s
dKSVW/psl+0qmaakf5nzKA9L0ffEOjnRs71ced3RsV7HBdajMjMxPGt/fUovansN
0kC+B7ArMZBWGYA9bx0RvVe8+YNo1lBb15PPIkKMCvkQxVvtt6AkQDMiroFvdZZH
A32nH6fOdrk8b4SuH2xyNWLBtbJX9dLR5WIBqvBrCPUn78HXMa3Q3GcI5iiU3dS6
siu23pYdt2MDdRjq/SdhKgJPXKd4fWPR7gQVCzTeFsZYFR4dGVo6hkELAXoxPEr+
4H5LGmxkl3z179eWgp3v4/3MXymzvu0SwAjlgFCBMhQt6DgQIYoM0Js4thubrY8N
LXuGOplA3HH6nnYwHzEs+dg1m7OqSIn2GVEmdr9iFapLxNGfOPiuhio9hvqV14+S
qachEQHG01kIek6tIrc+VWyWSjBKTQSTdJY/88ucQxUgQBNHAo+s58YR73tGxR8t
AUBKVGy4FMv6+yytsEBJiHRu1+C1sh7OP7CNqk0FT/rm/+TQuNdxnTiwkUBRyLUL
+MOJo9eHCL1eIEN5mPkJxV7b8qAiCdgTeSNsYLtkGzEC7VZ+y7X6PQeHp8X19eZs
lW9OqIxN+9286lgbqX1PBgD+uQwCA2PtMj2ANQJqv22/5jyUUlBDjiHyzVDl4HaM
Ptj1Q+Wk79XnJP1WOv0RhuqOFNBWVkQyLMwYfwB42PmJrpVxLGMdUJfZInnl1MTE
ddajGSZsQwRtfG99UIGwBfYcTOpOU9S/vhHXWuwisWBNdvowdOBAs7Rku6bC5LCf
0WAAuWhlkeviP5LbAjQiGRcekAjnCpIM1O10fGAeYhWiCQ9AvGL9PRZcievWpzMP
sHffBX4sbTniZOrzdsvZ3kAVPOdocZ1b6b+iotCiSR9a6BxdIj3hoZpBp+eXSc3g
4oHNh8wMyxwF9Gs/vqXUv5viJQQFVHg+jU/7tjbqwcUFM0ttR0ZG2YnLBolC0xKg
KlLQJNlEwUt8AORPOAbh3umNRX1POA95HaMFQQS25Kpe1JJFzZaJN9TbwJT1y8Dm
OI1F6NXju/3Mg2RCJCFd+ibcJ0/BcTlYWa1HVPpvw5Xas9VnZ/HEJNhjC3JNabCo
MHU69HZhYH+8jQSPG/DEinv3FZWXin9V17Eb6JmGgLXEvvNM3S+nZ6zANrx5Sct1
/uwMmY9CPhPk/ZKYro6w7a/NlHlFHbg4+i9faCPqPCzkAMtRLCljtlG3cIviql/4
cak8kx73dIv2bJ/VOJXeIYQ1LYoD0EtQ8EoA1QCS9NeCiWTt5qrbDbyXs+S+Kfqs
N9huJlO17pzT3HjdsAPd7K2llLbpm8C5uB6subrCLc6idG+wIYkY/40KptHEHr9B
1N5kYKvUQwdhT+A2lIj/jyG4d4QDm/55+Nsel0LLJuz+ibTqaPB4ajVsoGUnw4gh
stNfrA7kmsgGgefLONMCteB4NbGArADM3wHUiUKOYFi3Ow5n2awlaxjDTD98Uz9d
T8R2eY9Zh3edKzy3+JT7gbHOsxdKrjwljL9qIwEMvO86p4KD0WWA0PxdBzwKt1UC
vSevpJkxXU4Wbwkio32FJV1e4d0QI8b6z2JyUCWHNM+u9wAlyDJMFW2EhPyIcsu2
0JzL0ZVSLdieGsUAJ4s6KL2hdLqnpC4hLlMlcVBJDDPliD4RZ8bg9UXQqIKQvmuG
zjfDTBHv0eMd/Rs1zIe1/O4IShCojTHS7nHrCQ6VwqL4c/e6TrW6wMDmjWQi541G
TRkqZP4luQk4bqAY4gAeMZLsNqJy0segpfiL0HZoXm2aEdrNhjt+p/Lbr+s5yuJP
nx9j0mgBWtcMfxqhQzuuUDI+yzZP8RgD75x7sYPeRPyDLIM108wpYi2jgafXGTp6
ITnJ15kzxJWQt1xSGaX+A4KggMu5vCAzJhttdiS0IAgwW17+qvlMIiOtPXmPY/Gf
KeJjEONkGAIPb1HbTXkMtt4bReww2jE9Kahqq3dDHP+zgnATczMBTrciW9TctoHe
A267kM7EUF+d1KXuUBwAEYcBWYtxgux57iRRuWFBcxbzEqlW+27UDz0Q2jJ2me+o
mjk+q/JAy5t5n8D6JKbq1VXur+flOlqZESSXNKOucyBd2+1iD/Gkt4sDlkWmJyVu
u9SvbnXB+sAPddzaFG3PkfqNUs3ppFTQR0RDeBHncolcxsSRdEtlUNSDjHL/Xcuf
7isKMR15QGbccarz8YpCDg4eM9cO76FXxJIAZ9sGkDdR46GChIbgZhUhOMH4eniz
ym7a3mIelRX0o2aK4/krxgw7LGDmeOAA240PjKG8qyTvPN9OVKjZLtoHwqUL29P1
5Tx3jydG+YWU/bdv5J3OpgBj5lJK97fniIqDO0K69yHJqJWOkrnhG3aZ1K/F3j+c
SHuQ/wRmz3aY1rbvKAw8NbrXyusUNoPi+DEbnmaAhy48Aij0oeEDnssgMz5vbFO7
5uYOE07AbWyl+Zk/9vms5uVmH+xgaeLWazNyXwKKi0J73t4KrB1GoZWepXU/e5HE
6PHqbUnG7aGSS1UayybMt4oBVUDK1Aj+4x0A73W7AD47tF9SCFejpfQ4SLynV2Ky
2mta+JVFBsRVLlrMsi3mZioetaqXw0o7CBH2w1d7vPnvYlOXNYQgQAnZHyeykLJb
MqoEMAiyIAGNQTpx97KAZ7xcsJuTbnhLyhjsosAV5EdG7h/+UDAbqUMfvaKnyPZD
rpW95PeqLAaxUEQgugPPKyGWEFf67G3M9gmJLgBLOXn28whkKqSi4bDL2UTHbbwj
Vj5MsgktiWFwdR1jTG61kEiL3eYxcxsO3JG6Qzm385IE9EdtLBlFLXhwIXrxcopy
dZynsGPX9LyvPgIHaQYYJpzgF9QlVuSRhAJWklmvEOd78g2q3kdpM3T3/DyCE4Sd
ouQcEZmFurIE+IxtCbpP+lKeYnWPk8i7uouRKa85nEcPJtMVi0o6/CmxAmxtysii
hk6RFXxhru4AHspWbXJmXOroQ2XRuTQwiZ9D7vsv6Pq/uQodowhMBSLypu9cJom+
4gp0AHw/hCB3Tlo5jukx98/V+19rmhPRlVBSTq80Mf4TySQrp/WFAhyalMhn8CPT
c5VvD2NVY5NHIpFbx5AkprzoqcQa4LieVWhTjClmIUu8Bl+wNZC5yqJNqIjCFA36
SNjY1hAofZTKoNcyWgQCo5PfkewGtWZXX+exLfP2SiXeagayuLvBZKsoBCB39rrG
etFXsJd24CoRqDDclKsD9zKSErtCTFsnhEfiZB+EXz5drxrQkYoOXpCfV1Tzj+4a
W/g8CPF266uSavVhMqjwS3zA5D+ky6+LQW7zHSw9kHLcs/i5R/7wyYLr3Jr8VT92
0tAsK+RcP8Qxi9tHw8XadAGo0qBwPeUKPWboNGXMnwOvuJnM0KoBLWdnNnz4lHoi
OE4HrwH0VB0YArq+JQhAzmrM7euEvm7Zi/pjzGaS+Ggt1/KqdXmLTbixXby5epnj
eUwe2f1fk3D695i+rERLAi78lRpKSt9WrRg0oWjBdl8VCfaw8ydXjgrGhuiIFwWR
TIv/fMpZqQBCsK+P3ZPaBsxO8SiHp9FOWaOxJNxo3r8g0O91P9vJ8CI9jTFdc304
qM9vPQzSHnWY37na7XiKhRwLWM5X9siqeyrQ2ARXBa0hq2Ldz4XbqYtMzTHKYlPE
sJjvRzS1M7Kb/GRzbm879L6nVuq9ULHDeBvQV0r6aIgy6OnRKYroKhsFRxoZmQZA
QUNECyo6WVsx0lN0vfL/KoOabk2iXKw9NzKCoNIn3vkSeBe0X0P7+L2q1KM+GDw1
YQdkkHPRSEmdzCJfyB7fiMxnF6+2Z+VEx0seUy4Q1HqZvGpg+1zkXuCjqxQUE75f
eDMol100Ic8foSpnUI5m/EapiFojNR28Q6dGNqYiW05uHpWV4SRQUck7zn5mFyEV
NO1OS1QSw/YeeicAPRjtpoprMDDeeRlZGtDNDKMKr6OxPX0OoUwjoxbmdlwzX5UJ
Y3IdnTnT40HlqjBfc6TBTa/iOKtyFcGFluR6dz0c1AE0ytbmG2/96355NEe8CdB5
d9iphALtddjRizsmgO7zwjZmAi752kjE8wyhFJ4AGQ5pWlAGu2TuX6LEM/6vH6Ya
wJFwH7w8hG4m4LvCdo7OM6OnrADNh/vyXfxBFVLOj67MvpPdczfooE5aw9eEONhz
QNMh0xOXRCBAU9UdhwGGdD+nZeN9fJo6ed9yphnb/SIKPyWciwYvRtCN0YvnUn4A
AEvVY37fOxa24SfAhAkmeWInQJqqLsddcXXUXQGOQt4nQ4nkNNaN+ph2c15Wrtu+
S6UazE5ERtooJEhUV019K2kj7EBbUpIgmHeT2p4odaPP/Q5M4JQ11s3V7bgybgvk
eFy9+3A7qnLM5BRCbbt0CPW3CM1GfbzdOmgSgE1gjeD209KpO+YroWcQ4bLS2Pkk
OuAN+wM4hU670smR0QdMMa7efzyf39EFY8Y2KtaT4O33uEkDqKrHlZe7V+L4d0TZ
57kHkmA6PuXetBQpHcI6AoqPEt1pygZ6uAX2XnxGS8YY2s1UQfEen8XQ2vHDmstQ
RxDLcfzHZ3Y02BuJHjn9iXDspTR3uNwbxaf3PpAQx91Y9fUmQ13l12XLP/aAaiYF
770ISgZZP6ZbAdOv8r4lqWEPgNUDI7vdmXHoCxfEkW9AHwmevW2mYgEiUmY6vMUA
RKEJ9FLiZQ1vl6E/9Be8QsYro5VEJnhncDNhSaJ7fvg9yek3yjZTV8T3Pm79aMD+
X6C+W9ubxOAfBotzBoWkegk8j64qtmWAkYv9H8Rz5/CViNSvLVmSCCD1Qmttl2/O
JonV/pDFC6AoGAx8TryYUQ9ntfsgftFvgdYN8FMLEpjGjO29AxzojkRi7X5GqDvW
OclKEfzcBUT+AEUgh0AIamP6ElMJZ60J86Qc3lLK+zioq+gO/AsGtVSbZkNmw5eF
WzxPh2oVmZJCIhKTFuGnBrP0osWLh7396zKPwkXt+9cb/CvXwdDeVbuHQhFYB0YS
DHIKsIjVTOpOknwFitxnxwZOwdgw3MPpidJpBumTVO4fBtwx/BvWDGCfybEoSlYc
+V/1EySJC52f6KoXmxdk7hgeKOSCyA3iIQrVz9SJjXUdiW9I+o7p4KfClRMuM9mc
ITInc3zjD/z+FYK+vxbA4qrxMcwpDHswiJbmD/Qdc8qA9dks7sI7By+OF1GTQUBF
6uzyPzTrno59Jd+tUYW5taGE14D96uAh6sHaYLvhTYvEh2WrujOlqDwokFBTHTKe
YBdPq7UUf75jVKgsRLDSPcHIxQnn60pE+e+VBFX5jOVnSlwGcNVmqklR8DQxgVvB
63Je9j6xAxktDsd9TI4O0AjP5+N8n/fc6YAEKsBsKjvkHwr/k2Cst6KYePR2DJXh
bwQNtW8K5U/+GJ1VS8MYXo/qorxAU6CuWI1vNVbCc/0gtB0F/C5NZXWokzFjhYHm
Mn7FvDSJVt4B4ZewlGSKZxmiBM9l8PeDFbMmbTokooiYV281k28vxwC8eK5ibKdf
km3qPk0fZeclFLvoXH3ZFZzJk1jmda+4VZff2V/XmgxhO7yiYl+f0ZDvIpImNV3R
GL1piJOk9BVreZ8UXuJuFxrvfbziIe9akslE0baDC5IKvfN6Mo3NtGR/cPfQVnUo
M5RuY2s22Vp/iEWOHfR+1EPk1eEgeqk8szXXG7PAuU1KATU/Kvh+Cu3oTS1tFeje
ug73QOZJfyoeOvjrkabu4f/HHH4/AJ1np5VHD3cW0VgxCoA1qTscNRO467Jgl7+i
cZHBwFqddsc+sZsiKLom1JPAitcixJLPFxAJXbLjhCG4WeweFzu1RMhv/ok7o+XV
J15NMRZzztWZVsJYe+4UIyHVHesBV1SjyiUXbCXmm9u/DLutFUkrdag8NRcs+48c
la9ApdNI5TBfgkmXl8aQUAvZ7DMKj6/JbE/bM/6O7bTpvGCoz9ZU34fQTcOt5X3M
qZXFGJPsJ/6nh5lJ3e6SAD9fY9Bc55KQwDCT7PMpf9TvuqXE59aceRqn3K5EYP4J
WQb7XmKnXGQTe0I1Ylsu5rFdCz71HxuS3PEbB5icwdBThRa9q2asvkg+uzsmTo5T
b53cvHqHwshaVko26xJMjlc5cv/iVQi0aVEV/eI6g9dsSHKbnvcgxlm5RtchW48M
hek/4rE6h49k82ml6hk5y1gP9eua2NEgiImQ36rXbe/Xgble0isXeIIJkZAlS2p7
GxWsn3bKGQP1Gko1Rpe97BCt5rdUPr6y1qXywRznTWR69GwaNHeXNCWyNwGG/4HQ
HkIWYgApDHrTudw9IvQQaDfaRRiLfnpB8cL92eqt+SMoNyijjFiIjr8F0fv/s2Wf
beyeTlixQO5aVhv4lFlYMv8NbOQ1vTTxKw8liGD8w0G+tT3p/0sJd0UqV8aNRMy2
TLpPJZXUoJfMVCmRigjYN4KQ/t3/7TdcvpIdU0TcRV8AB7VOD1nr0/STWaVAgGQg
HOtroifiP+oPZVZN/KmeFZoRK9EnmqiPvrD/N8ilKqlAUeTGkR4jUiCb57uSrVHD
a56SYTVD3pqZR91J5JMPbJfXjj+NGX2XmqNOApDivqnuW835H3IOQs07OyDYAAR9
Lz11gozI9UkMOGPKCl4oFEIIwYTDktuZKfo3Tfq9cdCFRmfTb4icgUvPTYrP0E98
oK6QAcS+UIXny3N3yVtWqC6qSXbKDYXKoETQeAZXBNyTPIlAsDj+3FX4ZxOOBQJ9
uic2DzkrUqRVmkp5fitMI8zIUc7CqJ6LGLX+nLGjEQ8xKdATKW3CHwxuaKlc2fqP
ikQEvHvZ2s8XrZYlBSIptsS6aoUG/i0fjgWbDRzqd9k3vpC+0+dB/wQWHAf2hlFN
jhul41rtRah9v+KdW6TqZ0LmV44gAyUGQZnXMeC1WQlXYJw3fQ9+PMld6kQ07sr3
NuEsMo3MIeHmp0Ms55+lKA/0vXhNudSqBmPCdRM3mR+8xAG1isiQNF+W6BI8q6QQ
v5P+TbkLzx7TDnNb/rCV6k05KtH/tcWMuxCMUgPrU1QTm133fszgcUVYJyiFjJiB
4T9GJLD0X43i3YqGhqg1mdLPhdQTOraN2dHNvET8o6kJ6hSv/QorR42Bwp4HkWmd
OMszklhItWYzPx3lh0FprjXJxkQ2TEKTPEhkvy9X3zGzdGCN732cLhw0ZoSvEknV
BNFoVliJZEUevDiCgjeLIYjzV7ZtV65GzJN6U+AuM8iYXXskR8Ls8CG11qGpCMrc
5cbd6ukup3TECVJB06t1xGGMyX/LeK+yiT03CFVorrDbSen+GKZ1dpiMpP+WGZUQ
I/OL2WFzqj4U8TKqf2M3l+EAZE4RJ6apxNbQiiuxbVwR8kosTn9oLO1oJKELs1J9
oixPzEjM9FbU8RRrvEqAIBoWpyAlc5r4rHZw0NT4Q0o9wGdPKxMQCPFglgoLe3et
qkavOb4tjD+0/JAwBbCDFiH/Y5pY6eHW08RmZR4YqzBrKUT7sOTIRwuzazjWlaq3
SnTq7LptvKM1aOs4MGuW63oMeQD6q2LeX6Ww9H/meBh8Ncn3hnLlFmWbY1Oxuezb
40wzutRRLNaYRxIJqfagwi3mZ+9Ztx7afrkBqv7u6G14D4I1s/UM9G49ij1UApRB
uQxdwqZCBB4wz6xLho7+PWxKsdtmDZcQct4a22iZK2V5uqD/jCHNeQNDRXWw2bmX
4Uugu2SbsUczTxbm7zocPM4weXJn6pER99EIg7ISyMT9ja2U5iXgQ3e2cQMr5X03
B+qVsU/rZzmEIMCsRLIur5nNpfUviLE8yI2zK9apfAhhxVVTozt9sdoBOsw/uYAW
7qaF2YMFptwFWEz/Q9pCmTgxvZc8OmgpE75Jrev7cD+pzLFUD1W7c4j5jyWawyrB
6hozIwHF+8qrZ1O425N2gCD7o6fj711Fx1+e/KNFd6WBp4S0BvA5JBvxEu0d+zhB
wQDkS2h47hywW/W22pd03RSAe61Yp5R2fAcc+CSvjTB/Gg1HTVZHBNTdQKyXM6gg
i8rhT4x0e34zk1hjW0m/+AXen6vCfq7aTh4lVouvnbE1V5Uq759wS5H79HdgG8T3
BJJ9eHeOIpgfOW3IKltHt9Qed27AMwe+0UtfXr/Sh78LfKZNmCSqYRif+zZX3j2n
G5t7l2AI1a3eGJjyNxnkjrCjOkFoaLowa49iOTcLmuVTBubjtT9B84UdXlfaPW20
BQbIVGav+pWouu0bivmhFn6QmL+YqulQBtS9BRanfsPkYdu63jzfeq9mAQjgXE1A
thr7jzbKVTwHzbXFZg+jU/+N5D8WUfd52jQ2Dasi99U1RIKwAt/RClObbYwyYDUS
c334qXscX5YuhIA1Qvp1/ZspMrCuRJcMLjx97Ef9WsWLTTvZxaDKmM+8m+jU3GPQ
bMHq0/CjLjhciZbRXZVUO20Ysc+NYqo5jC48V2OXeHha6Zudq9+DNVcW5orqoppJ
6vV/ctuwqIFSXlrlYg56rQM9j6/YSvqa/WUfm/5hmDtYf4GqyMh9nv/tf2vpSuBI
+Cu9a7kQeU1zRzJx93sZhq99zxH4rVI3ECQF82fYMtsAXQuJ0bbP4ZuZjeTa4MCX
va1EDqyGij0/V/W3wwnK0T3+awZXNhvhztHn5M1vfC0E0gw0pA1Mfb2DGn8FppOz
IrUu/ql1j/FAnJI5zzzHBpvgYL6HrzJcWLTNDfmuWOJ8RSy9x3DS8906cfCmnKTL
cwgDfnVDZvhJCTWY7F57M/ofqKs/t15bs8g+JPDAmbagum911PF2xhEOkgX7miKw
XPpzvKOoZvwNlxxXtw1IWwgfgYqBsl1sNz/bRgLAc59ZOkLYXSsPwqQnxaoJTiLk
xhiI2TT9jMLJt7YzLE1QBjvXe4GIHwbZJcO6u+RfIyximrhgf2WOu7R5Cja4kINy
Ef5iMAKjMlMdksH7NItSqt9ff6od7ZNEwMvY+GvT5fxIcyWdmsWXOM+gJcchhfSp
M/vq75TX696KqsH5qJFOJYFTDe1U8Gg7KHfxSiiMB3VOOD+DTJdNNzh8zVN3w7LB
kIVu+cte8bVCAbWttjibGujTvj/nL8QPPQAGxrtPmz4qXD8uxSvtiyqxT4E38+Xo
CAQvXM5M/M0R84i08tjgRNfNUyqrG+MU7pjvWoqTiwLfr23Op6thr3s2uLYGGCui
WoSVTnFqPEvNJmhhtdN0Q0EF5lbIQtwnC2p0Fbn/BxQqAnM1/1gtMkxsO979oJG+
NtMcbEa9kq3lvKBZUs0BFe4wNAdcrPHjMtt035UM0/d79EXWVUSIO/53WXk/rBqm
xiB+6YG0LFxb/bupBFHNshhWvMUT+k1edwpuzANKJ2k60f29+y1Sc0OUMyaViQVA
T2Jg4rzGaNEXX7qZ+e6bjemTiGyFrte6Q/XQdKO7Fneo+LbpI8MgfLAXmtzlIgx0
LFaANUOUzE3v3Odpj64x38qfQgJKG835ClyH0d45avfBP9lXjZ3ezBisdoRYK1wI
GBSLFttUGjSELvahbpqoHRy5s0Z0Bxax2BOxO11MDYGOyyJTzyjFQwgk4RAfNYc5
aYzbtE0ElcoZ0sPDP8iCL7SFBn0UPADiov4UbpCjauqPnJ3P0SiQzww+fg5b0JsQ
HsGfHv/KgxHvLUlIEsiWBNxPRki4OJCHQKp3+Y/4qPrYJGmVcpNH4G9t80rQNkiV
qA2yXIiQAWo3b25JSv2Lz9bVVu+AxD3nUJht7+2sVD6G8Bp8QTzrQLMmjDNhEgTr
l0a8L3HmsiBPXeAZRYBA8LjQVwvE5iQ4HGkpMz0lm8ZX6lSRtWgtc7B/W56tgxhI
ZlAe9NdFmt20UOLjtu/apSbVs2d/plKoOiKKh55obaojLWFvQ7SGfnslVgnstNwm
G2aO2kmRMFnS1I+uYxcsgaHAU8wDmVECJ2mgxLtZTfDrVaso3PK5DOvsCLDwbqCA
/TrqzcY4qO9AbToMlNP+P5/IH5RIlK3oG43sumUM6dwnj7IGwGzFavS03tZLPBrp
dSyaEcW9MzhiwGGt+sSLk9qLe2EBd1c7m7LA9pKrHZp8phJI5/uCYH0syBYqSgaR
bhlJnN/C9n+gG2f4yZK/lZPF21/yZSb8jLv/90j+baKtc/3smSVcaxl1s6koasMu
y22ztI5YLLpUkP0C0MEW2USrFlcnpH5kzmDMZlxT1A88LQdUqNa034WKoRI1X0ak
KCLe3qZtW0VbfZaVxdEcOBzKEXsrbHRMFp9R7hBfphG/Dw+Xh+vWG663I4Pphvi3
ivnSMwuT6lzjT5t8kmrFPLzJsy3FFFvOOP8kg+r8fNYdUzwQXPw2FRTypMlVuFuI
TLnWlgODrQytrW18tUIrbc4uxMx9/iQd89M4Zf+bmOo+Kspz0w4z4CgvR69zzqWp
QHWo0x88SJBIY+NBq2xqWwoN9lyg+oLdKlkGy621RrU165fVHsGmiQlswya300xK
ebubmJGwRqEHMcflBGYhVTJoBay3dwPOcQ4+QyRWfMtz1TFZtIwm7e3YvKkO4FF6
NY3Tt4MQp0M51+5s0BhaOea+eU66RERHRA/jimHo7T3+8m2l2QxjaA6tCvQ853nQ
iYl1gmeXKECDeCuaLwfx2LbMR3NgLbm1z1ZhawRCu8ej1Cw8mhoff4dAvIGAuHEu
zJK06AodSWf9k8ZoNBxI2PYRqsweLr0fpP/uBmafiW55piMVEvWBtjDMCq1ESECE
JEjXzc9mJ8Sf7oUNGQ7McLiMLuDePSo0io+63N9jJkK4R4sDACPAHQR4FmMvZsPh
UtE8HD+4BxuGG0J64CkrE+35Laz026DMG2dwSUkKcUQqAqWY27h2dIcZ/onqAZ3K
WQngYVX0as1jBdy9o/CjbEXL9YW/iRUzLGhv2XgugML8GD0PYvHec8vDYGHzPG1r
XkleHW2RxEZps/jodEVjlObD3fRTvam0gKHZ2x9/yaS2Y0hLv0roVrksZjfISiRo
1rvgNBhF72uhpY//VcQf4i/PsvWcigLD4cEZRv+rePXh4GNFMt3aPAv8c5kDH1sM
V8HyWjXClcGUHN75tB7TXqeUYfjcXL5Fjv5AOX86YvXcETmXAt/j3E0GsNdXOrzw
P/Jju1NoJdYnch8z4FYen7Wj+0y9HZVgNMeAfUqNJXHRAOjkS4uZX1NjD/gB5rmn
Sq2YqwROAjBC5B0mub7e5A26VurE+zwzqCA6eFeRoqvBYs+S6LhNssAZ2I3vt+6p
indVObWof7CQWJU6dFE+/YHBNbW3WqXzgSOsQVIF7Kg6i/8Dga372toiu87NlHbT
biFGU1rhZC81vFUVWKUXzQwDryPRvG28SwS0MFVYGfKOi7uYZTLsWzeaUnzdhGNA
KfbbJAsCnJ4SLF2xrOoHwZjfJUw33iI39YfiFJvx54PJX4x8Fvg4BKNEBPxbUEFA
U8NfqOANruAyXG1jAHgV/lg2FsewSj6q1Uce7xIeOYHZydO/X96973QZykqYEYEK
VD8ZS6hjci/7SkZi6rRxwBQayxRpdwkYuLdX2NVaWGuwxbCXDDFKNxuoKdh+qXaV
R6brtiUy7SsEJtfopaoKDJHBzZCWf6F5eCykW7iYvWMUIVLLY/UHTbyGYElzcLbv
KmgMamDUo5Dgi0CHUb3KHRtGox2RJyryE1UHQjPUJC3uE+kvafFWdMYO5t+YqYSP
V0Ej04eGohLXUHstVsHpvIcq4+Jp7I0u/QfJSDq2N/qloHIbheYhj+FHbUVGXUh/
QMOjugcx7r2jj/C8Gv73wg5N46bgcnWvEZZzxSdgc8TJhkBP4poaoXDVoVXXz2Kd
VrleCxamikGN9JmJTOnr2z2yw3GjsoT1pkexnq7l7DkiGAC5np0Ymak5VF+Red9U
otrSzbdbwuESxGoCZqOETnv243buVHhziToyFZBue8/jJZRk6g2D9W5sN5xUKRN8
QA98g+dR7tfK4MfSVggbZwf6NfJsnjMfkL8INTfFwZ889Vrwa1J9iB6BXpD0cm9/
yW2uigO385pe5U6n8Z+2UrfEmVeT90kzPiXlNd+kw+p2kWp/xoKP7E6Z/eUEPkWB
L4Shh1GMh4cOFOciNxBQ/VoVDJ6IjKgFvdjauHMIiQCUybTTReHOSydvwGiiCI5D
aBvVkIFVZJP9gVFRp46w60tJ9Ham0kjFMBuao0aZEpbWxb33kvZ1ql0PzpjZo5mc
nEkFkUs3/DC+mykOB9RGCtOkSVUp96rkWg0m82DVjB0e0stn9WNPEvX+44YUBHJV
rNQ4A8RcEMl4ElymM1XUcggfFdv89OL+rOLATEqDZZVNhz5D6Mbwt8gXbF/55Wga
dL2J56Jc62J6bHFVOC5kCGW6fnMHLdJXHHg/NyuY80SnztHaH0MpvkrSldrEuFJy
Uvo7mR2tV8xZK8clCzHUIH2pX1hBrkUe69fla+06MjHIiloixrgDoDkSF+aqurep
TPUV2CNHOVOCRlLDqBKYaKQuJMD0OfbzkEltS3v6/2sV1TcyDUTEI1l0LM/Jzc5H
3Uhs2eSQExdId8UTewedBOBclvZqoEAkJZVgPgPiWUqxePtfjMshm15LZzpPorYU
DR2WNGbp0A1vhmbdhQQH4xdmRo3sehPaj7jYw+Vnl9p2wb1H75h9hEpbm8JXFYRy
VM4S6aL0b8Tu0wpAMzMvdrsOdO1iZHvag8gqMS8RC8d86Izu/NaVPLjeRQnG4IAV
24l9tFGIhUCSxuZtQtTCe17Mo2uiODeLcEuO6YHpHWKW7pfBVbEMsK4SrmEAWsD4
WQv3VqSiIFAsQd8jtWmS6sDviBOAEM+Dc8NlukRiko16bs3HqhXBiOoDrJubyN1e
pfNJFDHJbOX+wKdSOpbnpbrrKUt9uex0PZ/QTtgm1rs0glKQ/HWrHSUjoz8wdDwR
1QnI72CUeSxibkw6qY5emo3Z75GTr4P/tj9z9FWloMm++4j6FYC/MmqgJboIQiso
18ugV4lo+/84e2opFscZ1FmfJthxCxIDgbMuSOD2kDkuC6ccqA+cEWYS7eG5gsSe
IMldFxTHuKxZFZNrQBTuGWvHutI1h1MOIBjJutJmSnpr/eUJCih/e/l1pJ8AXCCH
lOBOob5HbxxqIbA3tsebli04v2ojq7aIJqIbCcOVQoY7nkS3I2wbXZ7cPAYVaXQW
vMXKpUsWMdLA271Pdj/jsIQgWId+GWxHOXZeT2CZI38IRkpAm4rrzITu0KsFdDUX
FtdASsZvTJKrOZoQPUswduhyTJPYf/rWcPIN/QrxFqkdZpeqje0IBhc0rWiK4efL
WHUTodyOy/7YhQTHyKdVP191RDD2gb9XyWfxAbAD+2+M9GNF1j3lF++00ucEQroe
W37cUb6MQgouZbR8BmyxqQl+QXp5LFe19SLAtR4OraOsuf5Tuc2lTa7PcPnGcmLm
eI5QKdeZ1N1aYvovtoucsN61FORiteQoZiEUgQMK4OJYKEcoWPtB+svkV8o+S5AR
4iUWWF/nYIsxJ3DY7SYAk0Uo+6+ngiKFJqbMvXgzhiRbKcfZz2lr5bfdAYTz+o3j
baToY1CGjwevPeiHIALyaEh70qAT8plxMTJ4Crcvhv9w6YLQ/qLkpEuaYVDIf/6s
rSGChBn8IooRgZpOyqHM8oLaaTy/+B2KVDqU/shoYDJqyDgwk2z2jUrfEhR8RSW4
jFpX3eGuKNHLhQ2b5ufLuHe/VL8zO5+/RkAuE/9ChRdpzRKcdh9NuQ8ERHI431B+
juhq609UIgOoPVOuE0vWeWvZjvKN+2NgHHjos3ZEgjZ2xOsI39oxwXXm6NNbrpBO
gk9UmVG+fQ4fyi9y0uED21mKJSQiksuvoI7KQjk0sviSF5YaVRrAbti8PFX7/iDF
YgK/ketMz0HwL6PauKu/pPYSHQnD43+R2CWVlEeDagF/et8+1DQDjrmLrWLLUkbc
JgU9ateIYXjEJXgfKCX6UJlsMmmeTZmaRer+sMbVlViLCYjqIC+wNZIORuWaI/ma
ZwV1XBlyq6wJlrC4respwn4KHr0VpvGQtrvVD3gYc3Fu1DR/1Ure1Sw7prLyFR3w
6oL1GvofXxp8tvqQIc6awuxzocnHWtgHltihhG+K1SwXugV9DipHVolmi3BkEv8F
yxEVVuMLF2GQEL//2ifeWVezTsKYpym075ng4DYmDxeud/0ROciU0dlu0Svj7L+N
uLBwH5zKXXUnuDL/BVrZYz0Xrel/uNuZTLu+to97/bfGF4yHUQs5aqTRjBYwP+wu
FI/nhZClpQWPCl3QRPpHa4iWiKRHS2WzdwKs6bRrr2U78izk76njcuIWI5JiEE2D
CbK87doLiaPL584KQXNJcE2tvb0UtJwUYixyPlkMELMtG58A6cbSQJx23D1bNWwK
q44JIi9axDyHieoFNd7SyVDWYT1dgwJ4Mm7u1Uaj2vQpGc6DKBDmV4dGDrQ4wony
GRCjc+xAhdfNKPsKEEr/kpYVrklWl9tYY1AeAlfTn3Y37QvLgI9wPS4ECrBKzjEv
ZojRQKdbkswqKuesHY96fs+iwvwqGFYlWht9nUab8egZGRh/khRs9xcjLmAs+LmB
AfUXTmpuCHOm4iOdzKB1THl/Rg0iJJmfEEL5UkSAbfMiszWWcehfs3u/NxWQuj47
/fzyupDGcw+JM42SMVFaid/fFjIiIIZyf8ceIh+t+pkzHJhG47UwPEVwqM5on7Tx
8IBEx0kWjbWXRAoGoeR1o1NZ94yBkqxLVeqiLa3TqztE5bwPZ/hmfRCFeDlunHZX
QuyfHk38o0jK/0uPboGvKQSKmBl0H72onojGO9B8I5as4JYQuWT14nBQj3HXiJ14
4KZb5iYUwJxdPyglEufAdjnAfB/gO202mEFMplxqiHKtEN+dLdggcXFeZycvdHhW
icEnRWLpm4WVPW2zuawXUU4cCBdyKa82+2jFMOBRd9za6mAjsxV/2Cnq3M/Tl1fv
TZtAoXTpXOWfYdBY5E2u9oNmIXFLMDsKbczwF3OTXnJDlP59ySkaInu7M2UBlHcq
csgd3dIcN9KWxKtzcl8u/jWBxKHrqSBLoePyltOr2Fo7EfTQw/bN2OW412dUFKUS
rcrXuHX/k17TJRm6A6smMPZzoqrePwU5xbdfp7Y+9nQ5S8d/JT58ZXrWsiW5jSkR
zC/dyhfmd+0PTy5xagX8mreDirkScKh/alf1qhX/sLaVZlRbxZIPjwGCum+IVKPA
IwnGZSzuTfY09Li7GU1guC3V+abSBYAAlGJH2gaeqs6piqptsk9JulkZAy3LFUY4
TX82VzcmSe64eD5miMiRSq69KwZWypwR9dA5y5na39c0JaEP5EyYtPSvFejBQE5u
MJr4XkN10EqIJjaVDEYPKYCk6t9JFnb+Ewm6xIu5eREMJKiTOwVfdpebNT3kA1n8
AbbEoJ+Ag6BzUxcqhJQ7S930M/jfWYgXLYK9rb/R/FJanOKpCKMAoRYJe2sEWntk
X/tKxT14MP50OTTx7foJbgkSuz/+mXztdW8LlR/8T/1Wu8wFiBhwYuwy8FhRz0pe
+mIl+bZySzaasj1rRQe8WDljuIOWxAA0WLVMZbFy9/56MSEdPCfeRTXc/1XjHprD
SFL+Xh3kjp/NEpEdRAyWqnrgmNAxqhXM39CPS8bGW/urU3oP/IvbiDkiAWoPIZ1y
CgPpiNifRpC0ATQAAwFoLLp3th4aiD4BEUBdEgOWcHaNbp0pfTztd2UupwCeynH4
jnb5882IwH9vA8N4bZXVYCiDGIialWptqKXuAzg3jZ8rSYAnCKn99vnDSClx0+2F
Igcl9xLHZJpMOrujcrQ0rMvRzkoI90RrALLGqtWdHDARGrf1aiJkxpxy4eNti5fQ
0bFKfi5/LQls/xJ17B3fjcoIuyJkNVdf5RGUrmjX1SpyEFzwSkyQppAQ0M4urMHP
O+5+M6ZDC7FEYipuKbk7xSWrBu0cXIpVlRJnWv8UBHKW6iR9Uclt1uwBgbY2YEyB
iw5/Ff6wAV9gCZgYawyvjUxh1eTPzjrNC0Koi2Bn5jhOgap5V6KXJYR1gLosdJKE
jA+MLfg+U8M7n9xBE3dAI/4adMSsNVyae2ac61bA16WPhU/BYW+0V5ZXT50ws9bq
swB/dmaFWkXCbzrPWG/O3u5X2au1W8a1JvYFL0lBqnxnP52edDPCmvWku+lcywf8
I7R80payjfoPcPuRM/M9rR/MO6S5she9RsGt34XjoSQKqTELUDeZ4Dzc5E+XHthC
XqWKXR5qKmqFE1MLX1AOm2bqZqKr6DoqKilwXY3Wz0TagmciawemP26ZZjZS7s9v
aR+77265Qo8fBO8jL/KT2dH+mbScs3t3ngFm9A+QzQU4krAQkIhAIgPQrRbHAYG2
wvY+jkm988MIUGw2EnVkLu0QcBX6XvZ2OzkY2ZiQDr3Xacl85FXimpgbBpO1L2I2
VdQubENZgriqQUwsCps0AwQ7hHPbzQGjzsu3sotBdg3ggLMpUyubYkGeWFPpHJ3v
3CC43bSp7FwnRfTmIyJD7BIU48Pqtnqhnqw5IvUtekyQ/WyGJr4Fs4kaqYQAEK1q
B+uiY/PSz20nKeJ14xySOAJkKfxvKXqNxDEA+194l7VNCKOwddKMdzQ5Gu6ot/Ul
4QczvT4AJijh6qQrxfilLypxnWEu5c9l7dLUA6VpMXL4tzbRYFsSycqdHBYP+JCt
lnEiAMxRyTpI/ABtvT/TMAEpZVJLP+CFuWXBC67PXyrMwY5qDNF0z9vkrzggoFI8
sjWbVxmEng9LjVBV7a62OjU94YuNMwFJGznWDcs0Ucw3WXA2bKXL33Uh4PyTkErg
Lj74UlrQsUwSprd778tTxlOtQV1bZwss6MVzKmfnyu5sxGR38irJKk2i4sd1tjlz
ArpVwN+W7IabQOdsutNqXt87nHbc0whVxsHTmok2HQVV9p34yjiwenuX4HWYnmlB
AOMi9s3ELy3uzXSj38yJ1uHDZR9Km8K9KGWSXOET1rQcG3ht1VfAb8MxBYS5F5jq
ZzYQmM7WuV0a91RK8Gdr9HFa6PqHb4wnyqPJ06lF7Pc8ZoeXh91I8Gf9Etzhq81J
laENlGX2mpCZH23uQxBqzDacLJDkSP+dykvza/ByL4p0qKLKQ8QILff8ID2l3XDN
t2l9WMXU09YQQjjTTyuQIwbiodqmpxtmS65IgO0wH6h+Vq+irhz9r6VZFOl319zp
hLVbnawabgibjNugpBuTQpt4qMSmUyJUjvv09EJEhvUYiDrlxzFx2SLimhEx78eh
FtGS64LkFQ4BcALsBFRT21Pq0Zt+DkrBvXEJrycxuO0kjlLBaxLmq3ek+SLEyltv
B5zjJ9nTvNx2ERxm/i8M6GRanUWEcxcgLsAFE6487S35TlShu5FUrQDcWmtJCNnJ
z2naTZliWtGk1P5BXN4dMo78vW2q8Q3N7EctuvAi/jW75RrJZjiMrW3ZkJ5PhJHt
HfSzyiFaWfrXHOemJE3azAhos8QGUyO7iZ3A7mbp9oOK1w+62sewSRQ0BHpD7I4z
QE/EA34GqmWPLU2llze86ESgolAQNK+13AwxbLjcdMbTD+lfnG466nU13/zTFSEL
pwZKpgJ/jYwzM+2dnOZTVgPTKR0IJlKs5j8w+PuCbtqs3lAOjnPQRHsxoGETE1Zs
VIIVETb9j49Hj33DgnBSGoxs9Kdc0fxPIzW627qEZhxZMOfSWd0axms5GQ9BkKso
Ty0cBBO2tV86LBZqbbglX7gBjVtPrluBnULGaixq2/OLxL6pSuQQwreFo9G58EwR
SOrinV+K/zANwG/gQzc0TU3DPiAt6tq8KIg/DsNf1h+u7mStCGzd9Hgt7hmVujDc
MlXtgNj0GAk9IAEn/iDdZQO/DugjZJV6vliHqvuatSqUnhxDHAsgciauwLtznbyr
SS4h3DPWtoLtOFPAl7fc7oYdkM6cjjARm+QtLym2U8fK/u9cfkgWBZkMiQt75V9F
DvzdKX1Jq0SmWMZ5TKWNLEOf6+BdssGn4gXOSg8t9Jkbq2IaiFF5H08kkQU2eH23
3Kq1Tn+yULrrcwc1bf46H+QwaWnWh/1mvPtIr18PTMOBuqmdGmMEFAZKoivg8e94
pfwltCxExLYF7+O7MSDCPrRLNceWpEuVtI/uvSvEoWgSb/SuIjrfu4q+ZOFD2YZa
KjMb4j55uOXC6+xEMTp7FQy7JbC2PzT3y/oPLS6/KE0XW7jvJONKsfHc8Blqfi/Z
/L9EcOKMak7jxUiQPZOrUsOChhgpSlZHVVDrzrQEhc12fUm+1/LVQPFicEfZ8jVt
rXIrBaI/8jkPJL160DmTZxpQUotLwdMLBkjiAtQsIyK762S+24HiErrwXzXN5guG
A99RCSB+MN2ZhURtaFOL1LrJfOo6qHWTpfgHJCv/Wp039WYL0nY0QfzY9vtN2swy
UMKws7hbjNwgd/vfZkR3gKzWy8Gvg6GmWAGq83vJ7lsfRcsaVPyCEVmPDQypsBkz
rLSIjU5nEL1rmx/388XutRJAWKoU8NyMvapAOzdOs2/TOCCNNpNAJ5qnyx6J50AA
co18IxQRfy5VLXUa7pTlYwOPM6/kFpGK84GO2Z7pJP0U0eXfipVE1QhHRFm9lEQg
7V1bH7YzNxpuVi+NxDGokgobA4UlJY0aM8il/0Q1tMCfhyPrwNwKJO9LC4VXmFGq
JSdKfTo5zTT+I5Vmwcw8iVeBdV2p/QSTwRBE+oDihzHlLnAz7V0Mq3xC77yKERSW
4CrBxX4dH2hHeE58Hcd53aJzV3A2PAPyQIvXrCTXjtDCvn7cwc5VHiNppz98atA1
yV4BQdH0M4RyFSx9HYPuP00sYLJInbFXdaFIb5GMAGclO3GZ+21EZmtNLohcejUQ
jxI4OhwdEAuTo3LSjoAMmF5qVSqQ4CwZm9nEbyzb2n4cFgVrAwBfCCojGwQWJSZ2
Y8ds7AHWe1CWAXArAEOF6jYBznFY99Mi/9sMCmp7PNUaZE3YNB/7WT8P+Vdi/UkX
0udM00KYkp8IZ1wRCzzXOihJnmtpSLMxeyqAyLwKzZP9Ymbn/1R8gAugBjL4sOmP
ulngKvr4VP/C7EHktx7pmK3uP3XIXXq94tWekjGFLqkp5WiCRWYGhObaDtW0mZFr
DI72DRDgr/ZAey3P8GJ5W260M9mHSI+Aal994lnkxvCpx+yidZdmT7VW8DyDx1WU
dnna99ajXxgisdI+qTZArHPwB+3KDJcVzfJYi/cyIr7CX0IxdxGJ/EyB3koHxnFH
G0lIBz9mDH6NY1VSw/Wchn6Kd9cfcgenwCJdu/pCKGI5gShNCDShc8N6ziHRBPpo
73zyP8ahDQWSyrKv1i1gNmBDLjNFqZzj/vtW/DXSg1Vx3qGoKi0O4nzZWcMDVLED
qONa60EWZ4PtAjT6FXtDkkFd8Bg3XbBF8SNJkaZTgOdHgGyECVIsteH6WXELhT7b
/CGWZA5ReZXjAExefuUf3MZ+cX853WedoNHpNBi9eH+T0beGISxzwC/Es5XhwZlM
NCCiJ/Vsv8PmFtj9hpb0TQdzCRLDOGv2NldeH6ftIIarP7+4sK6PyFNriXUxUK6Y
nfbTp0Vd2Z0YzntndpNRxL4pxeJC8WEiilTdAPNflzAVIZzWxehOZ+7c5dARyFwb
RFHLvpDupEhHTqP5IhGiByNm1GyOXiJ+2Qy8WBQiVomjHf/J2DqgEB69zNB7RfTs
4g+Av7QJpCLqiNE113sa2Utfn2CC/TZ0DZ3f0mRzCi7mHf5gnzuyHh2dXhVeFln+
C6WILtgmw0/3k8kyiewTj6kbtCGnkaJnXuxCDT4j+G/CtfKSjkefBTta/NrinHxl
x6vKu+D3vdmFmX7X/l2YhL3u4FdooS0mzpRer1d/9a9pCqB3iFj5PiZmGBd6L6r0
GCttzl7R3dDP1n7XeDV6TAdu18m7taS8hCbHDbYFsulEils98INRlo50BWbfJdoH
GBAWP7NuvUhHKr0Wgw7yZc+AG69cJK1xiY8wY4eqAFf+yso5TV7nFRjM2+3BG92F
qF46xm4yhbp8hL2lYHZl9tP6bjdOob9eeMvKwIhEU1kXg843762XjhHg6gx2iUqr
5o9ctn5Qkrm3maGgcZ2llEFPubBAl+i3xh/LrYKQkqoDOU7Eox8aC5Cr01AryDdf
qBjBrv79eHB2DRs0crfjK0QYZ+mAugX6bCw4JDM4zJmLij2OHqjggcBsVR8FuucL
m6aQ8RfK8t5X/WaCVhDMTy8/rf1fQUnVXNqgqNykKUj5LvOM9vMwgtYCwqm6AYMS
3gShkcNwgF6b+rkUIzjWZ/efsaKcLe61NvpR35uXIZ796SpQcmPsvQvxE/0057hB
g611tXNYB1b3JztgilYnGFJdOO+W8q2ra3a5F5Fg6Fq4WfpaUBQWgKJ4RCzggSOW
fj+mI2KrdWe/6++pt/0Qz3yVpafzvPkxcZEAOvXzc3INwph3XteH0bs7voujDsmT
0KDsL09DQjpJ2BiTJjMRl26gNNJI+sCKjsY87BC7A26lynzNd0q2ZI2kFqs20GL/
C4xTgF4zOdNsiAJDHWLlLKWdt1He2OLiuhYNDpOPULvgpRRPH+rNUVUqmHbDa6c1
hdGgbB4nyFBWN3dSCUdeJg4Zno5Pwb1KJTWOt2rSY9dP3PHS4WYggasZ8qJm0GDs
QnDZv+qx8ERCP7LF0UqcCbvW8kHYo80KGeoRrEFqHsSW1JxEmAqP3RSNenqg7Ihb
vSoO6NLFKMc7qJ8yWvcCUiNskilDtCwWE4snCp0P+3sGMupnts8z2JryQ0/oNq7y
ThdEwfV65lb2TA+5nQb48TeOwYLVK+u2uFVkB0ENQJwbSe0j/Tye2+7Cnq9b1XGy
wKz1AiG+F1Msv6Wsxrf4YaWdJxVeEaB0lmPo9a9XfkYNNGwtONPngt7R+Vttpszn
+0tw063pY4m9RedBvF6BuhHXgWGuEByYKICuSId3lHrRTqjeb67L9KPKT21/I8ei
1KMXoSNGZmBQQyfJ3ejLBzL3c6NrbeijSbZgNpcEPGEL6CiCuRHRyYvqRvB6vkO/
8d0aHV42+Xm+DB/zlGe/0rlHen0RblE2rRvFg5+pU4mETwK3mtotwvE4k8VAksQv
NC1NgF8nXl99JxEjre1er+oTV0x5uI3dsUHEbC0EKVf9olcH+KTbOhZSdxZ4zq/o
8jJbQYuDdo1NoRaJigYU8/0hQAo6Zoi7icPn+MMZLXalZPs4Vcu74KIlXkDxbW1H
+kjwUWkAJS14jsDAcr40FZi6Vu6HhjqCWqUDE8nKehsYCPoIlKA/HGxtxAxGRs0a
sxOjGUa3Aep0Uk929IN49SpWLrm73K1ih+WfdCuz9ohxb9+LOE8hGtgq6JWXNOa6
ttALh7YQu73EaebCrBoaeXZKw9N8FVGUaKHeIDxYgAeGQBzdhppU3henEYKgLEtY
rnbhnolKU5suKqf7Sq792CsxtfWHyoy7gwlbyKezAZbuH/069oDBDybJCAq7KL4L
W7fTRzbra4ey14cpSh0bkBllSGMK08rD5ES+lVGANri8wfNSvJ0MBLVvmJTc+VQ1
FvpKqnAt1qCEeVm7DvA6pmKC7t9KvmrToDxeCt2zL0HLc6hH+lCKS0iGC9+Klrkv
AvdZ73MBVP9WAl6kKZQ5VjSRei5/Tdiszg2ANr8CoCEYwOklAR+7Z/P70JTN6Snr
csjhgwt4EgFfGamp0lEY2NesO/cII2WecvXhqgxRi5zIEoGIojj9eTuKsGcxypxt
im2/jtzkIl6dlQUVXWTubOHh8xB3aa1LiAjRLan0sb/07JKlMPMzjVTw5swNpe4/
7wUm6RxoyInfas8vT0vg7HnLRLQvtR0L14mvTAv4m7heGfeGjhfmR4N5aj1FbvpR
CFuO+Uextx4kwpyB9btw+G8SGj8WmeMNsCtbOSCw9YfrFl6QCs9BfeyGQdRKDBps
SBGN0B4Vyj2WZbPDiqei1f31jH51IK03PdZzXcUsji5cg3Cba+qmu5TOA6arQEvm
FFfR9X2Sy8+0Sam5+Irlqo+9rwyBrvazYWZVOz1UrSMt9wotRLDFwv81LKeBH1YX
qWzHqbUNO+oP+wmp2Qg+eJH/MRxuwB52oRbfTjJmbfNObj9A68BFHW8Npay0fz4j
qZfP7hC6oSCtr1TrEkfl42dgZQ06HiWSHaorjTioRTLlINaCP2ywRBK5FR/GxQIS
7/4sYPK3JL5tZkRmlLQw84XBPXqqt4KI+4kbNkc93g7yS6SBnsz1PXDTcPAB9u3D
vsZbI0MZpeKcC75JwYhGU0Y16ebmtYLqBxou7HsSolgvhrPXFE0imnO3JKo6lPKS
vNFV2j4xBkf2YDtaFmPuHLJ3xydVrhScfgpGjee9pFX3sTs+ZVM4KJbZufq+aiP1
ZXX9fSwH/7p1zOC9EDpvYz6PjO+q5NY2BlIQ/ESF/66BZR9A4suo7SAEybUMNWJy
Ave++wzI32xqCR35ejNqjkg4rWl2qs6lYz9eAzFSr2VgqrPs39//avfk8ZcikX8p
1auBDC5v+RypLydmYFbjvhp+4pTGsYKqOHr8GQuqXbFvIdoIp7lKJN35lt6QSOk+
YNxP2PxNkgeB8XLeJddn5nqOupPEx0Kln2RlqsLSY2FeqjvP945vaBnHfZz9DtUv
M1f5zayduHTHj0ojWtlHe502h+R89EYPFubHPGLtLuPmu3vltgp2MJfgofURdZlq
gmSdYgo8maURBUP1mdAK3G674lOwfDFmSJDHE9MM7lKNTi9g4KGq6/KIZtcGHAxk
Jp7kfuv1Avnj/3mPyUSwDIKxK3CszlZQ6XXXjHK04maqyTfItQwi6PPdRKWT+B+9
4+9gb9al49FZKKXoz+Xcw3hEsnV4ZLPwOzreUEzcBK5ghy0x1Zc7aInvSsU9wZM4
X/dpD6lvI/wFR1HX83N0QFtwqrzphGB3gZtoPtp9EROUUvHsfADKrUgykeKvNf79
V35l4pDXfjCGoHeiSdmxn98ZpsLWQeracZUHSP66PnDGd4+Q6sMJECU5epG/eOp9
FZ/3dqtEazW79ZTsdJ32jiTaf2CE+E5fV1o8B/6RXRG+1tynfPQSlpaAa8AcAFk6
PEpLeX6GP6xfCahZ+qpPugsOizK+Fu5ltYN1zw5T97iOe//DBg/pjgC4TmJ8XGoo
lfiAbIYWL08LOdP6MI6Od9/LLnKXvJ/wb+HUeNal/W+6rAs13jx6LtJmnUE648L5
Lmn4SU48cyF02s+sgi4SfFyIayQtJBwck4YyM5slToC2iY9s0hIwSktWBIHy0E58
Fl2LjXuZYCppnDNZ/g86YJJ+adxMDfWLPeEQYNlIHUCIxZxQgc5PPAOUGQDfVJSy
i7IsYXje9lS/sdri3tZ4qhMcJj+8rUdlMhptYk7ff7bz+vL6Awb7hWTDiXuynmy7
qs4Ca4+m0yDqPfTSQrWsfpIwM802coqQL8AEM8mCIk6NQDtDvRYe04R85IJXnWMb
PgZOJ4o+WlDA2zKh6Ij2lo2oDd5fZv3ZQ5RGSzSFUHVvBEUUnm7LASuTgKC3DvFR
Nd27ZT0wuuX1XF5BCBIskRpMUeNqzC3Mbs63aw/rF38WfWE/DsD5gBatllgqZPYl
a3Fd8A3fTxgVIuBfwDM4EtNRCR4hZe3WTFeJO1/TWM0GtRlb5znenMpXUx1L0bmQ
6OIu7xC8x72eQAMUL5gIxvHmU1qTLy+7rUAGwlUb4TBuW1UhmDsyRi2K9et96HDM
SzJtNd+4S5cWQK15bv7/qx/sLAgtvD82/IGCuKg5Ashnvts4ot5y+fjMDXy0Y/mC
fulk9ah6ssLCHNe7FjVRk7lLkeokD+aSuitJCQzpS+o33+fumqpxSabOUKAhvZdY
ImXQFC2G1/ent2e/0nEyylwXF9yXugfx1tzLtTQ0DzkGGIzIhmviacYQpq/CEM0s
2cN5YWeA7NdhawISj9BK+7v52rhZpJiYJea6YLQQ8SJ5tQfiz+rM7RJZ2pgXByeP
e132wlTk0QRTJkKv9GbsuvNlURlVnnm+Q61EHm8q423Ek9TJKIpiTuR/1x/iCcu4
a8zR18K7P48j1j5lnAzZOQASlOcjIa0jJo0v/D2t55pyACxtNyLOsasuPds2g6Mg
3d6ZCZ30vQEqbEQV2ejqeVkUEVydPbeezkAgB3z2nMEbH0rSjneH99nuTgphLhWJ
iG4w5b7CBJp7+pDcu2C63T/erDFdIupuWUiQVOB0IUhStbSkzVnMHqmDKQZLiuBS
Rnf2X22w2PJ2Rrh8NxAAxa9QzpKtlNnb00scyF6rgDZelsQBRTXH/Ki8L0yPgQMK
enYsV6sAuGW3A+i3+ovAlOlO7y6UmoeyRGd6qAxsDXBmNcUa3WIpYNkMGIUi2ud3
xRxFoAgFBkSPObchhJ3hdGjR6jNIYhMWmErSDbeGKe/bUrxFM/PQh46C/qKvIH1a
Hj4AYEKJznE8VqzZELoTasVDsz6fZDPxuXijiBxfa4TRMla9vqvx12rJ0UEyy9qp
fbj3m+huftarXkt/MJh09W/n3hCiVBupPwHepiYKcbLSYVl7EIhHbfU3yhfTnjza
TLimbTHtPaUhXMIKnWMcCfDbNHsMsDHS/HCYrSqRgtWX1XQ6eMQ27JazSw18Vf4g
m/6VnS0JeoWevSFq/yX1THomKQe+IiigxQGQ3DWkMnTKwSnKLJUJa1U+K+wyUa8M
WTgUX8gzrCxouJctAu1jhXJD7ItCTbUoNKllxiH3nBqbIz+KXt25zucpDfHzUg1L
Y2p58A/DrJvyZNw5R4q3B9H41FwzFmMlrRuo2yHKA/WLUx/omaB26fK3XbFrbxcI
wRBRhYOYRikVMFpBnF1IEJ+q+Fa/Ge4TxuGuaPDdNRModT5M5tzyh0lNFRQuaCnl
CijzjkvuIC3oiQHQ2DfnUAvR8Q58coqi7VJoHf9GGtIUyrvZ5X7D1gDih6PLpZI6
w128WzXuIIzHObVh7sSnUWlrB6moSpnBLmEGdGZArqCUp+lebsIBAqZpoafaGXIg
yQ7r8FEjJDlGUEvI/rttL1owYBHR6LMNZM1YN6J8i1gUujUjcKsfI/xRnW9i/ZpW
JQzJlvbvYNG/v4vYToxh1lFNj8GC9o3vdshHgU8n3rmU2oXBzGhA3EfTqvK9z33X
FFR+ZxChJ+PyrZc8C8SqXjwQa+mFNsoUrNe2PSgPdP23L8hVitzDnqJ+rR+r8UNc
9+fvGQtYWUb56dxufYCPMwAVeSZh/T9INFB8ZUydfx+pJJBZTrVCL3G1ZGnnBhsR
cV6PJ1YS8TiiZ1yyY2l5+myHZPKk5LZr8xBBj0BgjtpkMIA/pVjS/hNxI2icBNiO
Aa5VtqadIFGWJY7/JpYkg8TbBy3WR5IkO/00JfS/PipbQc14t/UH9uJzaesjwNM0
yUd3ZnCb+kiq+KOvZIucLSxEuNtAi7ahZKHQBzitNz1Ufo7G5GzaOIwYFGAxD6aC
boRWfRKJYwm9cfgA2HSaP5C7QYR7u+Odum54FPdcZ3XaLkjILkUd5Ju0XHa+OnrS
FyKV2aCYrq3wwZUKs6OQFIS2hZgNyi8nv9CEO5+6ZOSefLkE0577t0bboZq92jtk
y72zij2cFgUCjA8Bo3lfkf5EM3MSjJ0RLGIbqRSDlFNroU16cL/lj5IolioJtzXu
Zl5wEy0EN1SWz78iR4A4cxUjvnVsQ8gdtpAfm276l8l06dNNl4YiLw3wmoQvdh9H
EnndABzCAWVh4L5j0VpIZpuGxl+9CPgedCrC+YWhQ8C3sWAlt0o3HoLoDWWPgYQ2
LEsc/CklZy4359km48xT4t+Tk+L1FeL4uZOopC41s+/fPkBYtkl6FDHfui2Qf/4Q
7TKDE9MYOGb3rVY+kT+NeyzDp3VRaS73oXhRGjq5v9D5UrXY2qKf64JhMyMs6ksO
4JJ4icgBvi8OZeqFTHs56fIgU1665p7Vy0LfwrOzOos0S44RACz7euO6o9/ilVUQ
t62t8PkQpEUPCGMcUMM06P1pIirc+iiI77fCkXY7ra4XeRUYZr0oNqSP6SjD3Lpj
hnvJqHHVPOA8XCUVaVsjrak1PfbelBKopAkxIxanuaHhP59nDt5Q0mK04jJpigG3
LygwKXGoMQdL8ukwNqtLW7PQOiKOmpfDblXG5xxbqCET3hy9h3MFppa3Sx4WJath
riV+m7CK7OfTYSgEvMSTYlKqxVzqgps1fBC7/ZQtDspFKVpt/CBsTqYlv5tBqC1f
ZDkbBFHfxsRB8DnAwdIy6ErfU80AZl3iWwmtHRW66F6SmiTefLCs/7ua4n9nwreJ
LPuNAGJ3AGXOiacd2+B7sj6+CwCRpH1UCZsVSsXhi9zKbfRHVdfhb+eCOMsLtlbl
iiSPrACScyLKNjcIkITEGHXawnIsCFpa5xNn8h9idJ8vbJyNAArp2FhNEb2jzqxu
7qyrJpmsuwyflRcZsotqcvev1vIH0essZjKS46Q2KH3ijm3lEe7L9Aus6kuygrdQ
YXw8hp3bCYL/Iu0/icw0XuK2JTyHCpJrWRlH2uItQjEB4qCdjr634qMqGeMNVqRC
K0Uzo7b90ylQ7Sj21YhTWAsUX9C5MnzPBMC8kxPRk9EHDBcFSgBgKwOskx+ZZiOZ
btwVSpbvvetrQrD747mqEPtOS/cwF0dKguevIuS0TtgNHbdftTOlsZEyZPCeWKIb
i6OrjAikcj7ojyYjtcwHemmUICk6InizcJCFom6BaTcH5pi9X7EDmcJR/Bw6/CgT
gnQBikJiSpJ1w6AYgYqEW8D2ZX6J7f9f6S+Wjf+R8rparei2zLfMYAZ35iI2EqUg
FIpd9kBOWA0wVOwIfVNVy2T3+06OsF6W3eS/E1E256/5+F0lBfmmA7saZHsicG+b
DfFWaY3yZxj7H1sPF/d8KxFSUYo7mdMRX5JewN9mRejdqZR/TSwUyzv4njYE4aCR
oTo/JKCASG22VuasRImbTDg8KdtIyaeFyEyYr41nWIATF9zdGSeSqyJ/Uw+o4XMY
Xqa4GI5PFH5Fa0gkHuhPKYZuEUijX71jXe6BGYWgQyfFxuImZgEp4e19mVyOzwKs
vJ8tg71o0ET4gzQn739C0tcc99kIRLdgipbZVBiX6sIBnLBpXmOQi5zoZ6rhHbFk
Yo8af3O4nYO5wZHfPQKq/pYfSSug6CktXLHM/x7AC0GHeR1YLri7YuO/x7W/pj9B
w+0x3RPo1dA1H9Opwc4I732Nyzy9pP5U9SNwV7eSK/VPMD6sFSgA/lfoeGumhNYa
iASUvQ2SkoqZ7gLygvIBG6PJVrUeN2vPBV7Xl9ksQyrs3hfrqQuINNioAh67GTYf
lfiIgvYN+pryINyXkUaTYIH8hRVyB5zl87AS4EdLYNeX/Nl36pHoY3mGP/6Yz9dh
vauZ96P1UsSNLYxYEZQwqHh+tfdRExrYekZDxd/Ng0LhRCjL7wASNUMQf1lxt4AZ
/HfECXNIM6mkCr7Sl9Ye++jXhAtQ5iKRH7P1SaKUqYSltFPD7glrC+WrZqP2caeg
XYdeureLzJHANgi7epDHjOeQOEUMr6E2wOOeZcIRiNLOfJ7oTUHmjXJGUdUYeE5x
nbyb4E/mhQP0IKA5ZdZVSikPoSqet5ugPCzPCObhdIE1SNSwGWpHFZunSylzIb3M
OjXFcShtqJr7tdrtyBo+90aTZjpCG9nhzqYcGVeqHGOEEZmo83DZmNXY+5xpqWps
xflM91b6bZjbX07ir4G8nU7tIGWhkhY2Miekr8gEasJcFWpGVyF4gFYlakzPFkbQ
BGqd3Y80fAqdq98g68sluagaP4bMr22nEgQcG1BbmlizkPD1XqLK7BLXTjVUTN9f
pjCjw34nuOjCefFMPWeecklykKr72SxsB9tQAWAcRkc8QnENTjXwjE8nxijQD5nr
W6YywklJtoOCAvFkc9kwBKzNOEsnS8OtwlNn0aMllz5Ai85C3mPR94BPg4iwAs3E
S2yCGxHKBQ23h3LUiewYRyc/XqlUQSVzfn2EqevnY/uKFgE5l7xO+Ad1OyWNqZHM
F23G+5qFwyhiCvwbyYsWMuuRRmP4ABeYoBUHsv+JokfbrFXFHRsP29QQVEDA4oDh
cWMPKHenxizCRpgDkii6IXBMuhVG7ev7l027aWyO1sSAdXf9dDJndTHR9n/eYER2
/yFbSVQRLE2GDZUdLvqhJlV10JXXbcm7XfI56Y5oiCAjxRWoHvgO5o6UoodM65F2
e+WqW81cKYI9Z7JMHjlDrGi4sW/QZJe8EXDXT512NyzzHJ9CI7JAivEPHJd7rwM/
rz0vz15+xwk07NUVfTeW99AGwun+ero9/rH08JCHG/nLU0/bIBHpOKg1JQF310At
ztQD8YVf78+rTzSv39+iu6w1gnExMtUHG4qs213KEBgU3V2b7yQXRHMYX61VxJZz
zjSa2fbKd/hIzO+8H6VCzMF0ss5oWDqXtfZXIsYcZej9T1/3NAGQz7eE58es3xMU
Rho2a/hrvh9beskXtGWMRgpB4b2Z/TipAUv1wTqUVRpCQzdn/SATxp0YadnEvnZM
jVOznstVW85il8XCKfllMEKb/f5W5Ucv48gEldO03q1NariFWLs2rGVWck00nTZT
ZgrLkifjnPriqCd9t2UzdTf+yPtFhXHHN2LtctJmRKyXt6o0V91bpBc/TVU//mRe
NjfGCAVK08u1E6Gvwfag4Tv2akyyz1YlhG+8fFZ3rJ70Lv/Rc/HIFE07hQm224gA
PpF4RoWT6eFP/kzCgMyFIJNCQMd/UqE14Ae15QDQgLh++FNDZTTBZD1KdTpdYehs
WPPQsaveaAVRfZN6biGOS+l+843MEkmPJWIqjuY1tayFtxy3ui8s2hCR+MpB8JOW
cxYrV1yz0h+CgKan8uKCKwnq13VbwgizCR3y+jsv1/eZt3q2lyxc3DrJwsGUmymD
W8VTdKHKDEcpe2KDm3wQhB6BD0uSUCa2chvNbgnlg4c5ZXUPhCOtV42ElfOYG9QX
sxaMASu0MK2jzEp7ol2RkNDxnH28K9exx6lifobidKJiH2aJ8eYe15NpECWAr2RK
pLYq9GC2i6+JOq8gXxA+tBFlAM9YxUZHABDxGWSI0QNXjLGKoSgsaAxvxavnhVpU
JJoeXPkAkBW8yIp7+yAnEcAcvMVrariIFz619iHfLeFnUCuCz3fpAzng8IwbjdMR
x2RAcZoUI9Z12ZQwimq2K73ZczNe8eOTcm2wgyzVulqxa39SyRUW/MwZyAz1i/+9
WmiG8aTALDYSvR6VkbUR6e5dxNsex6knVvl3kkk5QOAGZFRQuZsfzk/Mj+fi1C9V
U3SO45voEsrZMg92fq0eiLKwlMy7eK+2G2fGkUgil4nfesrpO0Jdyh+OiTLIYqUt
VSwuWF95U8RXXgMQqELpF8QyqBXz46ERBZBgQ0g7jKJ37B07CGq0OjIKXplpVKkK
2/k/FKsHLyGB+ceHhCq1IsWkpoAt22imp31Uzz0DK7hS1AWY8RebQFByDIBLQyEs
31gIySDQ8OLWR043AcP7zHSC4ilT0vjQRj56hQKnK6Pp+cjdVsUD/6goDHDTlmQJ
CAPq4KUJXyJ93FPBA1w5wEvKpF7rxo4cxXIcxAkoC8m9M6sJKkrGDOHBzeK4QR89
XtlKNcJn+KY93AQUSe4x3LxVBIRqbW2vvNIOcDXPNbXFBE+BQxLbP8vCdGkL4Kpy
GRl3zOW6OAzOkgZLJe1Y3+cy7fKJRSxZaE/Y0ocf27tv5vq3ExN120RzY0tHaWQY
OSu/LWmR4Y6dY71jAlMJKXwe/hweJIqNjrY2CPqd3Dqq4jLptacQ1j1KM60l3K4h
2uMzQM1pkGTU3kAhzRlo3z6dwjBZ81s3lAryOi4FquKB04/qqwPMa68dzim5frZz
UTF3HTUhs5r0C4jrab8XJ5T1KDILtm0+FzymBczvwaYbiZxSFf6D2Ffl6j/WCsR4
id1X0AqXhICWsUqxgnLbqKufxliBQlDCbqFfgRn7laeGaJ/O74Vo/GXb9d6gdGId
hQwuO887dljtduzspqxs/WkMfex48Kq5YJlsuijc4MX9zEnKyEljjIolnUknvfwT
kjyzwuwQiUlliXgrtT751qiKNVWIj5ESTl/wbr0bF9O+y47G5n6ea87z4f4atX1+
SJQRZNKaaagjkV2XmM4Il3vmcowIyAVng4Ti6A6S3COg0/GpFtq6jB9HrDVuJkA8
REs7DI1+DZP52hqXEzLFJjfNxZp2gWt5YrLReKIQ4qpe2JQDis67/HALCnNzJOfW
W2gMTDBXI2bH7PKNS4lYS25V0E570T0VGkX4C+3iw4rqYoHoBjyKcU/X9+bnXzjv
rMN82C9lyB1BfqEWP/CqVPvFt8GD3poV6NSgsh0FQgxLwl8rJ8GOxDNj8mU/HIBz
zXJ2tq+T61PUSwC2gu4z6DpVEXDVh+pwgPtKA5HR9X5OaWYkB+vvc4XC9BWV2OW0
pvMW/PoK4MJvQc9enlho8TwCYcfNfbY22wfGWyiDuCt+hesdcV8B0S+mcz1eOqRo
cyNl6Kww/GRFsF9FXRfFnF+FodjS4XnwU10TIIYZawY7d9aZmN/dm41zbpQaJN/3
vjmsWitDXNKWopXoI7+VKBSV42Fcc7DidYthYVl8MDKSvC+O/E26kcHIY8X/sBUn
+pIPOsCrNA8oRgccNt9vfmm9lTowXGc2ADafs2eVc8kOTFoWmEnlb0U0HFZ9RzSj
N7xwYInNKr6SKeo0r48KFM66SPvBZ1UquTCwMTFfu+I/xqvM1xIi8zUHtzEu68zF
TItEEI4ndV+6U1Tn5gXmWABAjrQlbB1KAWsGYEMJK8PSrVhy6tXjMxtLwYZozyTg
ATAdai6yIe4A+p5MDO3eg9JGLiIrRQHqAGHZKzS9QhJVpiIYvIjowfDxp0IOKSYl
W2f6/QpuXSVj8vD5FU1VwmZtauvvfQXjrTy+FoX/feT7uj8jS41yWLY04YSWD2Oe
sI/ZXNCFDIML445qQYsRN7lRwMYvGqo5ZR8Vndra2vcYsJbwShs33sPE45Srf6WN
xtG0hVVijvt3UKVXuJbOq6Bq5zid686dHEG+MhL2vj8/8foLoMeNJpHqwl3wbyn9
XWtylN1Tr9N2ZrGNkouqnNIgQx001w+DP5fCYQvukiiw2RwcGzLHqtTPns/Tr4SM
U1iSJCMOmkWr0KlN0H+y7JATInG2BvaHR1UX8f/BPQ9bRbih5PnU9TkeexItknbk
AqTTl2xNYf14vhRtXCF0UQkUTkHQ4i+TKrRjCYX9KdjnrQvBY5eG6+QwqNFId0HR
F0GzNLzp7/1/lEOf8vQ/ynYR4YJL8IZwHRzL4PIx2lmm+q8GmJQlY2Eq/H3GEOLN
lTa35w0ATsExYTCWFQ6N8WekZFWJgJRhpzR3KlTlATeT2AroOu8Q0D9MdJ8uzRqh
qftlRZ9RKhFwjdeqsxd/9iBDZot2CYxlYggeM89G1wuGQw/1Ali4mNeHuXbrykVS
XGCONSzkMQhNSam0HWlNT1nfH1a0VWRIfYyk0TowTJq8kvNy7RwPR9r+sya+QLBV
s3pYTiRITOMri9/5phE9JIMGiA9raVGrT6xx+FQx+1X5KqGv7Rtg1y1fJT+Mqj45
hpsdlC5KkizP6iqp4AJfmVmdycnN9MF4jszOiJ4a3cmJcx/o7lTlexTXeC3xqiqf
kNzR66pvLwc0WDdj+MY1peyXTvDcGR0ciYmIhFM/lopDjvMKCy7dY2a+xzineMis
Bl2bhw1NNCGPNlNW5kGvz9t4Ft9c8Xg2GDuQzDoXAxi5VBAH6iD2H1CG/+bvROg6
H15wQgzgUFXx+YvmgGPapfnYzNlIH777ionKmogTk1BecEWo2EWtXoNkgu47OkeD
SEz9/0enh3RR2bslHnM4aT5a+32tOdBhnQkBM6Z0aQTwgHtY8Dzi52bmmFThK1yz
bSivyCSlYDVSxwKHB9/1ogwgciZcc6j2ZhyuVuPpAV75zsj46iI+fNADdboy5cMW
ww+bf0tGdiNSlm0cSzlRwCR7SSIBBVSwVFWYXSCIaXTW7i6zhJeRaFYYzEjWuV9m
o8KlokcZkwoSdVxheqriW2+Ylu7HeFrQiPQ6tH+EPplyoIsOs2eNe66DWddEG1BW
by7iiNBkK0mNqdh0DIj9bb75rSjqkWVCQCYkSKTtdAFagxUKq5byvbIgIPLR+I1M
OOYrMaVxabLP2fr92Jf/8tDgsua/tD+zmSU831Pbu3v18F3qbjBGb/IHWY/Apaee
Ze4ZIPz0WquguP+eOOkrkCNL9gfJC0m6DzCr/PUZFRIt1wJa0rv6pjxaBqFk4NWF
U7JEkmlt/8RVrWmDqJCCrjBGoxFuQGKiYkDmQHM66IfMfHtwL2KJj/RECW7MuYVX
9xJi0d4EMsSQyVxV/TuNKx+sQv8HfkarsGppCQzLlyFOLsL9vXXwY6mP3ZuNi8Qb
etjNt5dez2kE1bHL+lXTakcDqfWix8VNJ5Okyolf+i/NnIb0CDjWF1B1WY2FRJwY
oqyn+fdBuwIyMHaYlQP+ARyDNyZLK+36QSdaN1JOoOlMdcWKtICPBX73Std6xuMv
JJCJ3UlOA6zc4bjc07PGPbIqQHLJEbwrzPE84JdG3iAVX/BmWj+12dGaNLcQnzPA
jcuFPWI/bB35gXwcQckc+N5KSdQTfUIiAYMO3FaqSHBTlZgYDE0NNA7BXW/U3Zte
zzJqJCTlMLq/O7PiiO4DwLw3trBPke5my7sCNMYNa3VrcP2Hi9ZlNoR6ez7pQOVq
CeWN5xIA3hsXF0sxdCc+6Irh5ITHqShUf0SO44qgKX6KjtxkJyWz9JJXVRDVslYg
bbj8vMaTl4aT2v4gtV+ltwh1NFKt0pMPDzjwMPW27kUXupA6hN320G9kGNeGAsiW
nk1nYcStyB1aIkRgX/MNwmhrjqobyhkLORECy83Gr+noQeAfaNDKsiIFuJFsN+gd
39JCkKft1oYzC+ddixkYtiQpSwrkeDxyueccJ3dVpZt7ihO/ZF4Nx8qxQtM0h5m7
cb7PVCqlWIT7fQiVOGcDQgmApbdmNRM0yLZctmevjjPNMscsy+nRt8ylmGhAN6Vu
sVt7qwdH+3Oq45nHOa9K5mQFg9m217le9AqAssChlTmLf8rq86LHpEXU/yEbQbvh
wtXQX3PcSbG1x5LZ0Xu0rN4Ri6diCES3Acp0SR/l7xoxeJVYFuE9o2qH7WE3yjWR
i40qcye6xHPe2cZDHjPUQNhRJHZtx0DY4UJVUU/js0/swVsuUDiE1OcynGaBr2HO
Jhw8YwS886JGFF7Wdf/pyFY/FVMfOiYEQoBOwvnMyxIDNPLdrSYGldZuM5WvGAH0
L30VU35RCcjTFJpSzZWNCU428gNQ1aONMcOpFylXGB/CCp46mW8/6Y1JeTMdv6m0
v9t1ZDlcwgW1v1LhdUlLwhsGfoWznIgtmbJ0o4gdkr7BfNXvsW0xDVwZbiUQVO/y
ZXtd/+s9zSOnb3929zQ65yFILU0zdvLAbtGmgBm+GlF9Ki3RxAeGm/eJDNvvvXZm
hlwrjzm/v3fL6NHnPkn7tV6vrEuEf1o/0A2asmsvkCIq86LYPoyFsBLnQDRUjru8
Hg5aunPu9c5xt7eOAaNBs8EcJVwJo0Az1/K6uH3rHWzlWohs/f9MfU+cGjWaAA3X
5AV8m0+zodviU5jnw6qziGLCXoJIkpQ1EoaXBmYnSua4+nId3DqbcmzCPH7Os8jw
Cfg3FU6JXUL/KhlxD8wqWWZLD6dHdWBSure5bdp6QXhw09vk9Q2GIfAePX6pwfnA
mVCmemCs87XQz3vzXLB0ZU2BPoH5S4idif4Qi4BbX+a4VGrBn405o+D/SZpCCWEi
yTFOhc5v38bL204tdELpriA69cTbIMPNU3WBhNHflwcqgMKAbm9gJF8KKS+aJeME
4Flv8WocUwCFtvd8S3P5NmN+QM5Sq1a+Y5VSeUPdxoJhE7O/duApJcfX1G7ynTVG
7GmMGg4/fp/ZpLz45Vzwss4g3tC8LKJVpxoTakcCGOwICcn4zp3tOfc15WlKpwBA
LsDhnR3Fa7gtM+xiRh9VkJ751HYqpyZniGfmOM/n0Ym7hWETSF44V9qv/GNgSSHa
kvqLCR8UmQ9ZB++cRGEVHEXBWl8YjgFiRd6oqafG9jlxfweE3uAgaoKkKSVoAeta
EWzg3Jx6aPw1zurQCMjV+iMvCIKR1B5YEV1EeWngzMbf3Zm0MP7WG7O4hvRh5mqP
uumEyBYF0xw9qaahF2au75upIk+Vtcz14qEDYQPN00wyF0g71QFw2pQVDZaH1xt4
18/4WLN9usPu+Tww7JIXlEaQsaMQ1hce/bWevaukX2REb0GDUip1oNh15xxpqQCJ
6+GMwM21WA/+zEPQ6r8FmoySHPq74yrcL9VByBn7WdWQZad1cGD69nxb7vX67hCS
9oohAzyiMR6SvP2RM7w8sBIfLyZaWg5fE5J+cOPXgoZmQn1teqQyWYOzhd58CKxc
a4pG10xL+TAoZIqv9TNsuDKmczZlfXbQ0j6wxemkggU2uU8aejth+NgT/LjAG1GP
cO+tNIFgSmtpRxw4/DK0BO10/utZH2yw73uWntI5/BFUtXG8XIKQVbCkHGQ3P9XR
DcZKMP307FYLRVyQl3hbf6tpyT6R+7z8lfAz7Tx/nz+ehEBf4goytNeYGsw7mU+N
XFilrGH7TwD6okSYvveRcjNQGabbLkPt3Z+64m2h+9/J6wDR2mD2eUKruQR3Zllw
Re5YsOzaNbmBIKfaLXKsrabta7xaB01przWsbZPOaQ6Vy6yFC1lY5kO7afT/N0xN
Z3j+CmN3O4fOEJVLq5eASUxX0CBm9TvpnbE1bAIOtihX8+H1qFK9BJ9YnYtPqbsN
Sp0CKm25Su+J2iX8Jwj0z7ffLOnR8SEt5AoOG7x06EBxeLT0gC+ICnUSRgqDwo/H
50MoKdCTnYiYIadKPANaYININf9MPc4zNktyFAkZ5vEJgLF8Dfdos6r64i5vBdr6
+C2/sXRb6i7rcQknGDPRvNfaweln4yKrGlGwCrN6F6AkuW3aVU930eynCN0gKd2c
CJmm6XWrt4m2uCKAKiT4rfgMunKirF/lbcH34WJgPkAg/mp69vLZseEVLaIrJDs1
uQK7/vQ684asc3se3tarpTWQhrZEtTBbdG88O1mAu5nW/b9+vnQ+NG4LTrJs2FY/
h4LYLKquIMgfOmqnR4u0My5f7tbW0sQq+ukakJn2jNb4scL4e23Y+C96/TxGloOa
FZMTkFkP/stMgKXkmMun2HhyzXa5eyDwmon+q6NOiEzHVuoskOWJGgF49O3mZk+Y
Y/zqwvNX7lvoTdAbJz7eUMF8xIjDfxgmEJTQ57SuV88c2f3UyLIlegjc2Yvr5UmV
UuRomHyh28DSn7ZXKYqt+VSpIIH7wGPnAvHoYtsp4nGW8/NwR8dEDboL9vBNFPsR
3TFtmAy7/85jLtdC2G25WZkyETTYLfYQaQ4nwtNKYqTvQw0T2BO4+jaFaSHPTgqz
5hWwfFQ6lj4tHjo/5a+EV5yo9UK5MTG6q/n229DckcAWtmayCGBGXBROm3zbPkC0
+t1ixBZn/+nImO/q4u9gQG+vfcdeebekAfyum1AD6mw6D3D5yJ1eMcjPbzr1GLzq
1Q8DsclWnTu4mZDoLGYM4x7R0Q/ROFQ/egBRFeO2w9pYAnI3zVWimToCKaqKSntT
ahF9jCpKr/h3AUrRDERqWuNdBjRb/HFfvlPJqzDBU8jHhA+j3oZqG5Gfrr+TCIRp
dr5ZgF2iODaA+uywuRdtna8ibRusIsIr0jCe/V2NU2TrPRd3DwONRaerJxkPvG2g
KlnohP8L3NGfm6GbUNYzW+rE2VohBolGBROwphlqB6NszrT0OhrDBGUmkV6qE/8/
1+trXiujTPQIvq50H+4xmciBZFitR0KukVx2WEIH3p7Io0jYaCcURPBEoEBj7BQH
UhN7Hya0cBhxz0xsYtTdQMDKSctaP3F2J2DV3dZaXgnMBGaO9rn2nFzP0deNoF+P
YzXvbk3PU5LaWMRptt0hK/wB4m2p9kKmUV/IxnEyV++qCVdDEIg1ube5ZCeUQRLV
O86UXyfxj/b0Y1JbUwRpegQWCBEA6mW4qiBOsd3NdYsvnB6vk7lUbdFvCFTi/ysp
a5C2m4VHZ143XrQXB+xup5/8xMNDHBidS8RuYYQSO5GzOEG8weusi5kBJObuz1A4
+IxYMfkSOrs8HI40qrB1YFScvne54E/oHNujR/69t8K/GZlHyl2AVWuL+FKpWrBP
m21xpatglObueyrm1w55KkpwYXMoX6IVtBE3iEgv4OPLsMQvXZB92Ow+poSIuRyv
d9Ex0t8QeidmTl+pA8xZb1aTtZTV/wxeuPoDA2wSJWBkduS4om1s+9VV1kNE/Lmr
r5nkjTFLmyq6DEhu3EXHAwpzy/5Y45J04L4fWk+pwenoh0cx76IvzMu+GYxW64bO
NDllQa9I0QnA/HpwfDNaWiT1cX31WaVuZhpfeDmHyrCOvbaOC+UTw5Ck0t8Kc1+q
qni9pxexTiLnhPYZJQBj5y81wJ2S1qL4c8kjXdkMVnOM7sRYaxANgR0g0MiHeull
DqH+MiYmYgtSOH92HZ+oThqcfUnCBBr40ZYyTWUBaW0LS0u5bxJOg2R8GTbJTaew
5/a+eHD+zjS72bZyropTNL46EVFDSzTfV94PUpOYdWt8yKlOJ5YUcDSyv8k7JnY8
FedrsSnxy5Ehe2km1atDaKAZYUsp2LCjBse7mZw8tZaCeA2eBaaSOAZpP9v8zUEH
zIwghoXEDxvzeLR26UWexaUtEQp3xM/kkWEXtiX3kGDfTnBMkQrFH7hOaaKnAwvC
sqYfxnPZJxBLKUeRkgxMphuxxrDmK05IENxfBtgoFaHjZwbYXPF5FNx01XDCDfJ8
E8D5urD4Bzank8+mwCE/7dT3HrC6SOhypvHp4DWeVPM/14DQsK4d3Crl/vGj9DII
q8YiXJ9qoKpIu1XocjMdz0v6QjWRtbXcZB5rBGn+Hbk3itLiieqeV2Jy6NbW21Tk
gidGxMPAcwU1E2NQVhDJOv+00G0yCSGfy3JYm2uP2Nlk6jNN0i0wRX2IU9oPGbDI
Xc4/OQuuz52pa/4sabsxLyTShb6YRpXOoq1U7Y15PS2uc8v5Hgv/fVRayt1Xd/tw
jLvwuKwXMGojwWBhWEdOMgdfJLvgoW/8i8tXilnq5NIYpizduoekuaqpZGa1Jqtr
G0pqd/P6a+E9aYGUyYj4ZyzY2W+icQuhC+J7pOdxS4regmwm407m7c9YoVPCamWz
lbrNPHM7TE0lN6BbL5Tm9t2HUu9P60e54qIwWnBMR0FmRVy5WPIcDY9VRxDdLDC4
XR4WFuAkHGMNOwrVGiF7gN3dek0BaBSsmepnN9Q/ipZudIawqVa1dzf769rPTzV3
vHZIaTPYUk2SVTtZjSOf0dC6nWG8qx3x6HmkEJZw/yBs57BZTtYjbH/3efVOswBL
K8muiWfnWikbWhgX95yujTaQu8H+BltCY03aFqLxQs0UZjpf0z+XwhwJEbb0+mgk
3HspyoDPobz5k6q5y0HZ/gzxiLANggUa5A5MrB1RP7ukcwmpwHIldD5K7BSaVQse
QOf5iI55dVTbnpZYnl2AuWmDDOZf0nlPFMVoEMSip4VXWT9HvKFkB3Hnk5H/Ona8
nWS1f2tHPP4CkswMQiOXBP9pNNuPWhOLXVLsgW5Dj18/QEBxnJUJZ3auQLcaBmf8
/t50LAPQ9X9D+rs27z2ivDUjtUPuDoJ/Vefs/K1jZxO3a2g7WvG0sI8qxqFPZw2x
A6LUROHIt6aOn2DiccwbnLd71ba6kIlIGl66A3eRxTGqNjfhRnUeXSzjIIy/L1kQ
5OA0OlgjEwN+pp+9C1YNlXw+Cwx5wepwv2TDNObzOB2xD4O7dbFgXU5KfKNuFLBB
z+rDJiH7Wsb6wRtDYRa82UV9Sn8l2HDEN722AQHyuSBElTZwGFbwnQQP0FIUuhsX
OFmV7Vcs2Gaqmcjs736VO6oDW0oCSk5a3Zjwid1MxqZtc6RQpLJsm/+wD10j38dy
1w+e5Oi1am3rolp1SlliPivWzjbVXyOZf/Bysjhh3tPqk0uNh5uW/2RdNYonAUZv
TLHlaVB3BaJjkVnBNuxbZQCKoR+2igho8m4TOuIHWs1i1IDFgnRAUw/ahpyzV5lo
WiYmV/gyn+/mdvS688l9BcBJwQ+b//tqos+c/ZxCZ1Upz9n4m6+sHa/AGl9YKMow
QePorzGAG3HInYw1biPB0mIv1VeFQwWQBtGt0Jf6uoREveN/1cn5fz7wbJt+DcxU
JP03NWfLQGVWWGh1Rxqh9PU9D9tpGCX/VW+KGvpxC+gKPBlgp/GjMIEMQJbvxo2h
BmZ/sQ1LGhUWsU2huDyvrSQy1Zo33gj0WaLqnCmVlKkrB6rcuCsUXNhDHAGxmF8b
BZnEAiX03awJR9bPBLBVSuucoinjiuJbmU0dCr8uw9Y7LrvPaSUqSH4SRX+ySuai
3ejYtMTxHIiuU7L6haEiJkZcs1oK35J2eG0u2M1PotwwSmKRkzOshg1XwvLq0QkU
TrqyuXE6LC36909J1nwUHaUEAYdFtKYa0qLGfAu2tCo7V54lMEicrDokurXGavXW
d1CQBqeHuRn9iYTWjo6Bov+K2XkvRXALD308w6btbDEBgNwWCM+kOIGUUTTS86wi
N8BaR+rIi9PCn9fBVUbdBw5HwZtxgrEpnHcffxiNYdILcRrMQV3VQN9R9vgoatTr
+jSBTd4xSua/MLcHdJ3mIDC87FXKZBzoPnpq6/wrI4/N3BrVPTYg1HBdTe3f66Xw
XILFtmOu5jkqbM7NXxMB9wsOeW3JGd7jkIUFEiRKtRcheWNd9d2AazYwjWFZS1os
ziIcMSHuFgQQpwolAYL4u2bK/t4aXVRNViCEILShn6mhOsjue7vbPZlS5ALpZ/MW
Y/AfczuvYv0uOvkwZ5eWr9n2G22J78ZP06trSdGk9uo73/Hs6+RBWMNWnQ56avAY
Y8pNmvpCPYw4IXkdGCunk7Uj359dK34PSJ0mimSCe0iNwnEs5OIAhELksqVBO7sZ
rFeRgs3JNIw+MraDCj7DH9V4QkY+JAZg1Lbt8Ios9UB5Kxjpppd2iKg4C1l1uRqr
xwz5+UrDyJ0pQMNVWgOIh40q+eoMDgSpHaFixUyzriHjTifvdvrfkiAUB31y6B7t
aPvQGMJqUgxvWI4b1Co7TGmGXpw44+3m34zv4wKAXeH2r9WmK8XHLMNn8jAB/Fl4
CyrKLUrCEDyReeRK8WoYjvX7Qc3vodx8DkvMHQQfxmRXHK4P6+X1aaaG3r35iXmV
5ou0oct5PrSM/4zNH9NVSipG7lQCcivL/atL+qB2ZBy9cgemsBZIC7xwXTaXKyqH
oaPE1DM9lL4oIjE9nlsjaxM4KIYXkwHB783PDAM94ACqOChefkk85fslbAFJ2yCd
s5vgewTZ/0MVy6VAYhzjpVb32D/eFXuCs5IKtMYXYvxlaoMGBuLLU/Ws7fExcZLh
858c7we6UWD6zQXLffT17qYPffwK6CAFRvqlNOquYnBZpcCSQX/yLp9JEcKiwq5/
Re0Kjfz3hyuUiY1A/mN7EgyBkrLTTw6OH8kDdSXpJOPsbKxn5o30eeUGp6zxr34m
+J7uBcYjBKPzlkM57wcwfV8r0LH4kJwpcMdEJJaPaalQ7coiCbf6LV9blQCQEAvv
yKWFkO+Hcr64RJEcMFZusqAy6VtMbL3wdk3NQS71QbTd2c0bqhtOoCybIfjO3gAN
FLOfhrIvzktauzvyCgSUwZgXBSrp2FT1SOT5n9eQ4W9Gwa16FO/dAaTz7hBtA496
2qiNMVCMUi5EdFWhM/WPPPXUAUA505zIJVAHr19BlhOf/1X27D+o9gVLXNRm6xxy
RaCtu+g8eYcQcMbR1bMz552VXVW5u1T71+2OGzYPb/rj5IYt6NbX1YZixsV0fjB4
BvD/c/hsfpF+m2FxbZ3Knic3OhoANvIGO129J24JEyS4bZklmTO/GluX0Z/aXQjA
n5kq78uL8VSXDgVx069zvjijyUEbdVBLHGGRCK7hYEHghYHglPNTWGiokENz4VYu
4jJ8ZGb0SuI86QpifRuDzag451ll0dC4R7R75FLMMn9iWXgV9jYquWNJcudVALFP
ntB/nBP+fOxfIHuCqw/+m3KSOhAgx0sQVRwoZ8pDD04Xf8ADQtsChjf9y+ZHo+Hd
r96maXdeQUDhhqQjTg6Sd4Kh5zkyo9Vm70z4SYuYUXDvGIbE7Q82m9ahVW0F8W77
n8bGip+rVYMQtEt26AuATu81JE89C5/wSms5QA/VIyjQp3VnhJWsN2+Mu/IIN9Bk
a1pLjwmARTrHR2+8NJu7jLui9MrSoCGgoYIi13gL9IaIce1VtSt+dGbZEOmyBh1v
17XgN7ltb9Be7KfNogeYkhbFE0XhKmNYaGPUHc5mF3Exzf8fjBF7XeSxhbZOsZf3
aNzLtNsTwP5zotZ3MtbA+Y1UC+SP7Ttg/PWzsQqmwBIFeuLjhtZfqgTR5SCDEpYk
UqSeCSH8C38bkhTuxB8NH040nowR8GtxFGaXeGN59dK9ApNpMPlyIhfJzzkycOOy
QV3fm/xUlU9YkMAhVBWB0mESeH7BaJpRt8VSVxPpeg5uyOMTbKMwytAVpfdXFnvZ
2kwWObpVlF6b/5MERDPho9A20w5aEJAhTlHX5VhGOBznoYJzNEvnB+TOlDFEWFrq
wBkKAQoRkBzRmXWyxbXjWtdgpjQXBObHd9BnK81WtY5buZlgCgPD4e9hlFrDxd62
bLVU3vRYMu2YEVrh0TzVC0UuRRycozYY1txvaKNVdsjN6pLK4lSSQRkk4Eb+nagM
AwN7h8WlSkDlZmIvrhsg+9FdJhktNHpInND6yTysDU7Hzehx4Qi0YU4653PJECFh
ra+gCtVEqMmJg2weMq4iMSzWHQ/DFic/5J1/mXHmEKZOr3tnf+R+ojGDktjpUfF4
OnjAxX7ZQmkGDYAoqV3qCHuXISwxkiC1R07tQ8AxRxIWTJJVMG/fPoPidLrUntkX
WtoagY0EMcAfoxqHnOVa3TdRS8ILMwq2fiXc6ReA320dxMR9mVLVrsQ0DvXOJDmX
JZ8GLJx/i/kULHyK5qLYK6Rlh/Eb5I1dnvffyuZPYZ44SlaY/bVnAIOeD6F1JzWb
EDfIOlzSCBYZtv+IcsLsPd6IJigY7jbiFY4Nlk1jBDP5Sxude6PV+3wQbQTrrAOt
PaSC1gDE+7ZXUhkJaBeXjqo0Pj6g5thMF0ds/FE/YE/mRRzu7eIbmE+saE0IuHqx
Frje7jzI6QH4K/st6gzuXiHFuG0T/BvaVMddwnmAMbEj+agpHXpG/UbJdqsDBljz
e3ea/i3bkxVovid4Q2pKdFF5Zt02TlioNVcjFRK4PWpS40aDGNK3vOC+sZVtZlcD
4YRBwdnqaRi+inO+IAPx+4akb6xmrF6qrnmw5dg829zSKlbi/+zpUVg4CtbX5/30
3ZOsNNWnbjFEDo8hGUfX5G1eRhppWNfbGU54YgSm5hKaSzg/GxPFGBLt7eEsL1gO
YrRDX0GqE4Y7nk0mH57/yQImfR7kpHmtuy/u7k8jB49T7zd+IHMeAyZnN8Zqpp4D
4V6mRDs7cCJZL3Hg93LK95IF8qspVnnxDzggSXV/4MK+uaaDaqcfRY8yk545X1X0
SO9vcQXu5w0WkHfwdeRizflzgheFLM6gXW6wcl4botA4/8MdsSor5X3W8tJ3RvsV
jNZQjm/Hh2e6/dDgm2o4Zno7NZwJBidghEA0hGgsmbsS3ViPfS11MIcCB94RS445
GuLekyEyj2Rb5YJTzlasT+oxXx8xoJau/gxouU+IKQwjZKFLYIaKPLtWXwuMIN0P
Ebu4mSVFjZFE8EnvNqxazJR1NDxegdo37yDxYJ12S/BrjjM3Nyi6cm/2DAYa9Ueq
XtS9tvYNqZcFJvwjLpdkI8deAIR1yTfR7xsB/WdtCJZc+kQ6n3JCFRfEcVPK5ur6
pQvst6uCgQ6bT13XqXVpLhbte58egaxJS4AIAJ9I6O7/c5tOMkjoqZoH8AmZKsUE
JmoowId/iWyeIlOpLwdAcMOygTvN077mZicrXmO1dIY3L7uSGN1+ND10w3RoiTUf
mN4GWBYsdYnUsA8zIc4SNaXnYXF/jwDEahdbKM9R0Yxsi/g8ndc9eEnPTlSKqp4+
LylZVDBjr4vcBJw5dGAdpLpzmwOjwrdJM5wnJgGGNx1jEhBMvjRDlYHS9JHbl/su
nQWy6tpjeRCw6k7qHgshCNWsxVgbJlA3dqVgdU+6w86FplHtXccvq8sq/uKfjLnl
MzkuoyWywahUqDEuotsw7uLbUSClnkUAoWvtPaxqxRJIdku8/eQDw/AUzSn+r1In
Jzq+UZPz6QIH8dNrHlexIsSPtVj0TpRY/88NlqGL4GDo8O6DdEZVghSDalEE7ZS2
wigtzDRoHVNDPpxBm+qTg7vrFKP7cAK57f605HPMt0ihzx02bn1lFPPFF5fmSXpK
w+ejeS4hZ8YpnYX/4q01l6FKWvNz8V84seQKmSm29ldIq8ygr3/zikErQCFbCb3B
RiUs87PAz+2iut87ArsbiAyXvElzxiiQm/rx6XYT++9i7RsuHsXGCKNh3YITdtnv
4gqndPkSozUlfqsCJFzUBGn9bZr+ksCxcbEdjzYyYub/2OdwnJGm5hr95r7cIBPo
nvxD2grzfuRPNd92qDm5lYAByLMGYKaxz98ECCIOvmmSjHIwuz4Ha5U+BmE88oL/
70o6tnFHGa/cXghbqzLh2YUTHrJOJ3HkJ6ax6j2QX9+lAGmUbH6YVlw6sBj0Tvzm
N2PWjt833EqFXl92RTbpP29Ns9ru9ate+U1iJTMezg+YbDilSmbfrBAev4znqVhn
3pZILEvy/mg0VXsP5Wiz9nfff4v+iKK7QtlYxFPfWCU13WG6NjZeL6LWuA1wHlvE
yIMACk8B4RocDVzuadDIaSCT2ChWo3DOciy5xMRug6k4aWzU01lLfAj9y7l5Iee9
56Wh9FWl9plGQ/zYAWgOjabPNOhbkXmVIrnrovTgry2NqyXlN93WV7HFdX2SKNin
R2rzHnTiJCT6cdVpgda7J8Lf5voNy5HlCWtmDu0Yh0fWpcczd4/S0wl+zPhbkQ+I
rflXEpz1LsXAu1znRW8Rzo3gRWxMLxtZW471BP2wn12xLb7xw+NvsoqXfd7T99m0
Wczoq+EyEC6tJFOl3POQ2fbLVe1wrnMfTGhudlaR3Ctf8RyvTA9fnTx9/+fnKEYj
KkzIhFkjUdd4qTZn+9tgEsuJ01gnD4C/Mjeft8QA4bD6VkXF7IxIjm2FzRpnuwhw
Mr7cEOnuJlY8c8NzdflYf73TtT+4zkrmCwJFH5ionKXvhE03wY/Gtga2wN1A/7Zm
4QDm3TJEioHXY882ldTyZp8yRmQ34RwN87jP4hQrFy37Zw/nbuWPdUuxvJE9S+Rq
HsMn+sC+PkJan4IEvCOeVZ0gci5w6nV4wc5FF0re0sQbgq3+NAGmc50pkrX7mFhc
/7TvsQucTe2J5DkdNwOKgaDwtcugr6OOEAXKK+rZEMSUhKKOwWdN2M95xRQZhtSN
epAa27A/TrQZyMUyjZUAJHWblMSWQyfwgXmh62lU77f2UvU0HDZO/Uh9mAcrMqie
nTOK58SpDHwgPzH8co7Zj567cdoK1BH8A+Q9btv+WGwSh/YexOFnDxIUQ0lvTbj7
5HfOUMJCtVE05W56K/4PtXqIEDk8WbNTqXlzDepXcIOnzEmI3wxUWUh9rQ2gs4qm
RdHiBQrBmKi6im8ITYitxR/3OU0wIv2SZIZrZStVHfS7UQr4EwOoHj3uki7y3MXY
pFNuelAA3ZJUMRY83Ojq9CxloMxSGuhCyuydP21xXGB28FgOlHtt5vSyk8DW5a7q
VJAOvAa6JkWxReIf9d85X0TTRcBvunKxSPZ+lyv7EgVTIQYWGC2/I5kVjyxjX+BN
tPyVcZKCZHVmscDCXcmfaa8VkpJ5VJ/ilIb9Qo2PJ3LylIrr/0204oM2d9ZUXgFC
lWzjQgFh5vKXmHicJV0+MlhqXu8LZRT1FHvRnBlBxOHgUp0DUgF2l8MT8Jyd4ToI
FJO1lfcatSdMKBVFDfowxHhK3xQRlECpVWBjLwMjP/yYPqR/62+5ecBGh8rQ+6dC
CxejijHuLPb4cvLSABGn++n/s4yrk10bMoXY6d2GKuBb6zpBtDclYY3yo77tXalP
+ZWtZ1PYj6I7msR9yLh5ykKugYe0Uuqa8TGg9T9705cLssgKO3GYUdOWl10VQZbQ
CGWKdlysJyYSDF1HYhm70DFcKM35w9P/grMdrD18LDycPitAXcQW+J7ENhqg3+A+
HSOHXqygmFgsVBtwzfSS4sQYKbIHRGJ6nAgohzY2v2cd4z1LUWNsIqZXmRDlF6eK
Lywj05LR4oI5bY5DmknUBFyr4dwW//XlIM5XITB1i8Q+y0+7yADM97dJNC5Ijg8h
1Q5koQszQGUnnv1iGX4JUJ14Q+2PspxKt/WPUocA2TYUbIutHxjp5HpYcAr4LosG
Q5FnMmyneCMTAFwwjyaXb0Qn/CzGOwUspSraALWj8/hVxbNqoA0Ub/1AD9Q/gLN+
h+iJsgMwVgr3iUIJR5Udux556KRS6TvfFHEAOVF7it82XBMn3DHOiBwhBj4FYN4S
mq23UPWZ9I3IKmYnzas7Eix6mo0HYzGlHZsPqu7yKRISEtCO1avZPWLWEenk4Q2o
b/KTMzG0s2YqzNCWth+BZcGahk0VKpvdx1+7X/57bs+z4QD1nRMuFS1tTrAGYOLZ
uSgvYXWl+VYx4A8w5pfhHQ9CJFQ7KaJPpi/RBaxhtWYpDy8Uc5JDWa9FNv3iVMvG
oQ5ru0IR90f4IIaCbs07PBr+tG4C/6JCEWsR9hKFl0FolGj4cNxJH6lkI6s4Io2b
b9jKt3LqFawOzuWOih22LaVp6EcG7x7OQOAGCMRNHlMjQ72EAG0f6vkfF8LjfcX4
ecZfPeFh+e5v6RP/NgEcn0M2XU5OXz5HeBCO8P5wVH3JiluCenytV2adLCuWXLa6
4CJZ4cL/GtEpZxyCrOcLfQ13sbVOSt6OGSPHUEAto4ARU8Wa7kj9isQkSFjbWQs7
wofX5XF61I/p3KCGiYQR+wGPiNyDz0Iwq29M0Dwe++BBtbC+O2nBeIMzjxjbW80c
+wcrb9jQns525s9Y3Xp5TLjJfoMWJLzn3492ZTIdOLEM91WsAkXNfJnuz063EHNv
3Jq7ZgNKMuDAh4uHvDoRo/9tVpssTh5Cm9JSirNsnPXbEIPupPFOdDHE+Lx+anrc
fKAoJDuHHS5BQO6BIu7/yS9wUjp4HWmsVW9zFjrlNQeMK3m4dhspgX1otSR+Q6ll
vbJGs0o8cHmGoMqHpDGggMQW1WtXrlbPCaMDe61I8mUiXxP9OwfqJwmuLOLmjJAd
eaDk0+RnyNTn3EhgbklK3mRfKujEaRjDA8ubktxJCPiDjg0sLKUxRchmxHhrd8+D
OBTMb/icKK5HlkMDVPETJA8oU0qCKok6FKHNlZUgIrXeKxsTgJTQUwhWPtU7cgJv
75EoJh1EGWj2uDm2K8Lg/SkN2+dG8HCMMump2xouY4ufATsbW5gvekqAh8nk5OZn
EGVb+U7q65Wa3IBrnwXEOJH7HRWEvcAvbb24uuR0cX+0B00D4iBzecky80BLFxuq
IAalwAwk4YTzvZWejOobPX9fYwn5w6Uvjj8sR3KUvth2N662oA5mmSSwS4XZ53ZB
VaDfFYZGfimRWRAqnYVh+ApcNjmCWvLOBQwPM0oDSAEIcKYy7C95LbAfabShG+Pd
R5/cjDyBwRriMecRsqZ3nmh/zy53Mwu6TJjQh9/TRcSfri2nBE2XzPC+REQ5MWBk
COVNI30NgZ8b3r5Dm2SlQhKYGHZ6VFT6DmG5m+lpspsVxEtlKD0CF5Jj9Z/iVNHl
Xx6MUoobLkWFnANpLybjqw5zpoagqzKK33c4Af0zYVLHKy21HxKNlcJyj5ZL6Z7M
ccY65GU87NXZzSFsOilurqSJUERjTi+k+kFwX0X013xFvpHSXF0gZ1IBdla3HHF8
jUCAxO4T9cM7sTRQ1UOcC4NzLIs+9UVdvBD8RJCs3BNSOhEvXsAf7gQ0DzvNQZfi
ZANvfBxSH88lQC17D1llp05qzw4n/cnC6+j/Sgp7eHfNU3vFMauqQof5ARVTHZxf
Q2AL+1JsC7In4Z6oqxM7mtCTAn1tX2ieA1IdkPqCG5Gp9VoBXqCwErhXjK7NvuDZ
XH34GS7JmlYk4RpGSvCliIhxJ7Pa2FQS2KIH6zIabgKPPX2NwqZLb3Nvq1hgbKHl
NDaha2rNq8N8uUXxbBtBLLxz5lowwy29ryqxEi6bAcfQ+tFNlZZX55pTsXxwAkqS
UOZLI1XvSEMIzinVU3DZnvukAY0az7DHz8yj7F0Irja6Gv/4lbUhcplwsyz0EQfM
LvipVr95Bf9BmqhKJk9NZh2ShhrXFA5UEy8PPFwZdFLZO/2GeHTu1y6j10CFEjSC
jn0dSH4nHmbnt9WlG8nQfpIZKYGxV3KAkPdTz/A5u5BMNfBLkRWjwJvOeHj8etGv
7PWJMzqLMXNXJIXhygGr4mXUZwQuNV2WRS/oAqvLyJHHpR3+fuL0abPNEvIV+B7K
cyPz69I92U5Ic2sG/bO39GkV3///JPHhpRi4XjKUZ6zbHd0ZSPsP9XHNURGmbdZ2
Lr+z3DV5o/d5zTnlZ0hKWzcL1IgtOAFacYBKi+WRBDHDkwGgV2+nYuh6qRwehEhc
doOp/bEHpTAeKNs6KCaTUp9MLLH0RSj+1VC4wxzi5aJTKjharC25AGzDr7Fo6edu
4reO6rurTMdJsndRbZ12wiFrZxQwiz3+/Got+cS0lCiHfPzUbzfcFjat/bpsAe2D
sGxGONCnh30tBLzdLPmcUnYJKuVsXNcLQlC+qH77a16X3IQf5fbyIBNXFURhiy3x
S6+hPEbz7b0716mbpt9tZ6XBx2QQTcRY4+ScAEjer9DlxItSLWjanvx6vDeFRk6B
+VcZuz/MIteAeE/9kj0RBaZC01w9G1RN02p1GzKvieVTUsAI+UfVS8ptQpRAHLpT
ugpvGnqVIXdikCSgWowudVXIfGOlA20YoMCLbN7lHvd8AIrChljZIl34jm9NrMJP
/bcNr/Ehf/jlwexP7PSXZbdVCn0aM+Tx1XM+5RtLhdj+f6sTcv9XtTvPmw+8TwKw
SUn0dPPsfflP4Phag/OxQAU3FXcRjFwmMGgrzGt4jS9abPktjlVV1IQrEdzeyjBy
mmc3yU3eub+/1I7+f0ROOnzuUn1OzJwf3DDRhS9LF3v4McJOWOHF4jz9c9N3HW/t
EUX0jjf/Z2NuaoTcSzGaIz9+pK7qI8Fb+63DysgKp3Pdx/Y3Tk2k1x0ikRWhKLld
kDxckdAONRKWIRobK+zacUpnImLNUj7ymUOB+hXqGnJDVDsFNjSTYHEQ27LHjjkr
CRQXZ7ts5I1ReGiU4StQudBIKg6PMgFa3VOUx2Cs8KnTjQRR5uSl920U/2nnI32i
/kypLghsSVFJzudVfa0SN5MCbUgF2KwMNy/uezIz9NNVc2lNAimSaP8Ix328hzFP
kpzQ+XciS7Xu42AO26o+Sr+dMH7OxnSC8hLzj9AjfADQEkXoeU/3elo7rdz6vCG7
PI1pkqtqP/7GG4LUlKtlx1UP+BRjwKDpKkwt25bqCXj8NWlW1wwpvdlGerAmLZzp
nnItBz8rdTkwRH4V7vvXpeS8zjcVVInTl+9N0rZXEFE3S0wrio1vlMxCGhq7GeTu
prhqwTvU56goSV01bVLKKMPtj3I7tH0zS6331A3Bg8eCMFcl2hVNptmCqqkNq3Cq
mpUyh9XlrLK3WCdfT6MsxPGWL/MGOy7RfzN4wfC+eJrylYSLDd3xByV0phi4mf6S
mMSaWBuc2zQWVdnZfI6rtuVwj5L00siyoOHFC03bZfzrABusEXoD4h8pGQS11L7m
C07A/Dpq+BAKh4KVzz7cPEax4Q53I4C55kvZuyXc5JnYX5ybW0u3LhjTWy8EveVE
0lyhbZHFLi6Rg3OO9MFzrLlknR/1QGZIyslL7MbW2uyKpGYM8IS9cm3w3VF2fKJ8
+u2eqXcXWSdC83iRM6RtMQg3Zseyn55V1gzI44tZlarPKje2mKu9rj7X5ZcdoG6h
iWGZyHkwTTEZUZ9UoBPUzYllrzabXAGdANvNp5v36RyTJGohV/aVEspiWORy7ofl
m14NyAsgjt7cftH4q7Lpl/5jP8R3kvhbG59JNIL9lY9Cm2ajlYU3iIhE/icKdAST
FndPegac7qewtMf/Hnp5xbs0PTcm4qkIkp0XXdgXvT8vgGmQOJkeGFal/XkzUmyO
W0Fgq3X9YDub3qbOOZOTG8Fal5CSvHmDkgnTSAWbobrfzf2sje5jaGaga8I+ewmA
h83+2rI2nf9Fd27xrlzxGoedMeBlDpbvGZiKXmDGkPvC1RmtCps+zHPTAcWZTwMo
VUqLdKH2/vAu3h389R+0rhgJ8oA1e1Oe+X/g2I2pDSklQooSEO5wvKvKKBZ5gCMi
pBDo7wOdPrm1pdH448lVMhBfz3cfcrScevkmdcObTTYUWyV/Vof1eqtzUJ9NWthZ
N/2gEYHab8BamUAI/0jXByfRiTz1rhXSgZQU+uDO5416mRm7LmWEv7Lxv6fUZeBP
CdnTjeucugzeUKBeUD0COhXKeW9hVxVy37yhqkCrSf1kOR0VXsj38YpFwVy/C+qw
cZI0S79MC7+gGKo5Jedn+dbuyM8nFoYh3JWh1Xt6wPjR07GPGY10ONk0Gse2ifWN
DHIn5yW3uLRXz0i298wF3+1OiR1IEa8JXgTKUMtUrGE5xLcX6DhuG1QoHhVRG9si
ZUdVQ16Vfh3QkD7Z0NzADwFgRemb3f3y5Ocj4Niil/94bi2CvJZ47YA7ownEkmLl
23dmlObZklj3UBSNF6sJTOinVC9kDO2hdCruOargu2pJwLb2eTbexlpxnGqm8Dwx
QB8UMK/QdWsXg3p45XhvzLV+jOzts76hqEgpIuuZjS7j/u/T/FGvxz6aEe87Hw/3
62gKRo3iDKBYywQLZXc2zZcWLlxIIDWBi9a1RVYA9a+AGmcYqqcg3FuvlovCQwy+
vSIphE88aG9wfj1un7FeE66LuJu3kvFZsE4gE6/B6BvTUjz1ott1tZHJJKDxmxyu
QFAYqKgxLTpsJqVh3HMtLUOBGOMBqwfETSxqJSH6x8Vv0cSUojwSYCkC71yRBlf1
3PG0Nd+9aRE0F7kWn1zHYcFzGDRYAbYRAPLdiVvfzM+bcmuCzDXa4qer0iQW8xVl
awgais6eCHrk/4wyxAZAQJcO/3gNjKQUcyImbwDDQu8CWLKat2qqMeHd6wDe1TWX
o+c08o1JJ1QuweB1cFJa/2TT7QQCfbZjbUxFoYqZ842fjMmz9fvmq5Bf/qiTneD+
NpMjAt3x0e/l/9czMT6xJ1aVGAW4D5y04CQrdGMAblxD9Hr9xGuqWPuOjVrexK+7
hCs/pFmtBPNKyME0CFdgqHRnodV0U+WXI3Mk4fWDuMIbNlCVpLI9VnC6e3HLeyFs
W4mg/xjbUOolNqwXYSWYpzbYL2ghkdNgOgNJho3i2W7ijxD9n84T+0leJuPAWkp6
7XSmtB9ANaulzrOGIG2yCcltcaTFkRaStpDJRrANEJLQ6/L6meu4qHQsQSqLQxZl
6Be7iHHGE7GyaZKEYhKrBQRKCCR/yNXhsJhxkeGoF+eAn6szULypzaW5YMoxkmR6
LlUZ+rYAQTxvHcXGEyKcaY2IOEjGnFZLr9ujr2b9kRaW9m5zwX34u6fS0QYCjj2U
ReXdpvjL+Z3sUg0gyxrH0/6nlDpNQOxbZYNAgFHRObCuQ4qDanEuxYDK3P03mtH1
Rid1sG3St86kzPDHSx9KV0uczk0Djp7UYlE588Rmq05hMZ86QGO2xh2Qehj1CkKn
SHvWCEkX0Dq3gwqEjPbk+G84sb8zWdeYB1aXbHQLiCJ8tERL20SMgY2MVF1WnUgD
AU1v0IaT28N9VmFK7oZnyQEiGNslru6OhCLpvjZqTKOHSDHRhW12wxIZzLUdbmDL
HWsgPKeIToljfdr8QIDRkg3di/PfsUfcWwD8+xjvlrtms3nTMC11C/wTEUfChwyc
0gnioswI9P1uZBvFiimARdfPuS/RDqZmhbnYnWUOgGT4vgoVRLAjIGqBNaWiqQPe
LPEUEjklG31pxbWdN70xtsugAuGmxAtZsnlHu2Kla/kto/E3iTZW4ExgED3oMgXi
GNJ0LF12qHoekCPylG9t6PYAu/0xVkD1h1QU3GQGPy5nif93aTNG4mkDBXKe92j6
K+8kH39seX05o/Xc55O8Ba1kD/6SDmbrTjbPCqYC62gDN2CfuK8NuKsQjJNbPfjC
cRGPPEUo5aSjq5E9MxrVYeoOZAk69OWtVM0kjFVIuCL9+BkaXoViuxOjz+oxe5fb
F+876XS4+0EIeVUePYmuA9Vwf/rn0plYaILQqLBWPBXR77qAPfQboMlYzS1meod6
07HGVxE5IgISJp5r97xAzOeTNRXrKQ2Y/MfyFlHAWBSUVZqJoXl9NKmnsLkrdhai
R3Q2u6737w75+8pDRDZTqAQAFqVEMdmIJcpKV2vbk0KFc0clQ6JEKg847LyQFGrM
vnhP77QQVWNIRDPwGV4hMclxNDXXtz/MPARpBZqu58azsql/ewXsKd64Y+zH4PvR
dwUOaOF7xViiSWDJ5GAiteXpv6mZwBuTsIonnUabgtGaCbVVIS+lwCTA/Ap/NUlb
NNNwnmio1/IfOeZY35pFtMBXoqyS5Y55lx0jTLqu+wt98Om9GkpRKBWSEtd53aZj
kGTPADRs7XFgF601llagYCN+c1GvoBM7EzFIyPPVfmg5qQltmWlZBkB3UcdfMXkt
4OtGBDIoZXkvERv0+qJdyI8UOIPQsmspp/OtEvz/vclkTRPfU4K1bQnh7Vv0Jgc+
0cceKTqINgJb3IpJTCQSFaDoDptZXb8zBaIomenrcHRDcF0UAhDJSwmZNic7+9GU
06KGQNejIf0ksstKCNA/IURFYzj+8Z8hpcodWzCrc6EiQXeg/YpcdeXuws1GxGlx
7c90/rQH+u0KjjxVmkxpBB29T8akNp5c5XtIjW4FlaOmaWW6npnlUifwB6hiSYMo
xKQrw4UxuGOoNqIHqwh47JRwh5pbjxFyxQk2BAg9KZcqL8YcYsQS5CKl/xdHoevc
5hRYTRDbIXdzyTGrrQyhudjMHvsR4ykqjHsmgG7P2SBK6E7nduurpLehFMjJGL4f
PXVRWL+DcDeY4tjP0jQolxeiJljDP2D5ZTa1zkC53BqUfdFbrAdx6dqiDoVLKxf2
A3VPihWsMATZNVDStORMYr2Xs/8bILbM0+8poXBplGWq3/sHI9QLKih49U25ybsP
0y4Rtv4PS5pfFTm6krocvtHQ6lp8GY6+9rT3FX7rUQ3Au8b7PCnvRs/2ojkJOFRV
OD608zV6AHW64GuThoCBn17K8lzNAL1LXvV2D0ESrvB56GKn2j18sk8E9a5kQi4U
cHoVa/MUY5UepYIWBjKkrCuN9ikB7lNBhm9q5nENUodjDLvVvGFOTKWwTgyUFwOS
vohVwGfPYbfz4eS+QGuHLnN5S7UrbM9Ee79LH5F0SP8yaINsKGExWsp5u/tuK7zM
dqhdd4bNnEn6MnVJJlLWPSUV85ZU3FEdJoKkAT7NoGsn7eRToqyT41hRgaYKLage
2MP24NZq1l8Ls9VR9F0Be1RN7rn5IJcVmfuaOw1IaM9wKz1JgHHcqDNUcfYwSw2g
eLxrzk6brJncd63ZeqLchAuVK2JaC670fYWrs2jV6icCsoSGNnZXpRFRX975GiLZ
p09CFB7uH33JwHUfExsSYBmK+5IEsdISOSXfDx4Byzv5HaAJ4i+nOwQ1nEm3sKvl
SGYWrDIbtGMAH+CccqkEbxSw8Qx1ZLJVgH4h5rB+sMf5QnmN+H2Nc5Wr8T5WnWAm
lipaiNatGL6IPae34nU1fup8IUG3vw7JDBo40JaMA7I1+AALmP0mYSoNzxDXaQyu
r69rFKOgn/Qs86dOdefHGxEskK0A5JKIRdhxff15NE9oldxuWAJfQmMWB4+6k7TF
vvG6HMK7YvFD++fNnpbnu0gdjsV41AD8D4XKAgKzgepztvLkA/c8slNSuNMoZarH
sb94Op9aVJ6H7Fj7NKB6O02EjdjdtY3jSIxduqovxH5TeIFUzDztm1d60X/IZhXS
wOdVr3qL+Yr+6dNYCYcJaKIaIEO0qgN9ohu7KozDi1DctABTsr5G0H8kY3XSIen/
sykS1AsdLvYYQknx9X3wQEgyDSwWIRkJMdng5u6dV6yS83PNOm0TUHGlpQShJ2o7
C+pu+V472Knyqpe2eN+H6S/KwLcnvEbr3MSU9VosMgrGbFXYvQXYmjMG5xvJqlrT
17x1+5CNHCdolzqCW0NLdRpPFl1hDKiglfvivcleiR/XDDX7H7t5BFLwF5EgxNs8
obS8/OO2eM2UKIKUOFNZaJl6IecX2hwdK5BkG2rHbgB2/SDdk5JHjp0cRO5WeHQ1
1m0wIDGpfa0EaqEj/eZKodQAuppgF67cAOdsKho/yOPfOpP068sjHeYpuFekGVq+
agk9g3M3jwBCyA3nxlcTcnjAkNbiCVnHrXcOaYyQz6hdEFQQuOi7VkvWi+AcYveM
3KgtTXZBovur8VzOjJehF+yvFj115+A1gF1RAvzGHj1l1q5jiP6bvHvKQAIgML0V
oPNH1bKvb12e7Yo3pM4U8G5CdURakQLyfbh4lybHajmJ8plvUwAwhKYHlnlhFDFe
jQvlvJX1P5r8qfBJiF3HaSS822cgl+Jy6v8dJTJIxZYB0oos9QhzYUCt09W6N3W3
xmT6L5BggDMjU2VIJQgjCYRF4rfURLjR8gsoe27GepBldu23Xp/q1UjrqT45t82A
rpIAqhRNS02KpbDJfN5dnKRXjdhWi+igBk4J4OBd+fNn/sVk9Jbbm1fC5k9clKQ0
fAuKE7TSYeINbQ8TfbTp7xafAyTcUKxvMGLlXpQiDthSjMPUT95OcodMmoCgEj/z
fNrnGZQqpd2QjPXs8DNqT+I2aZ56EOIfjqz4Qk7mrPGK2BeT+Zov0i0Qxp1ulrLV
KzBhjuaHkI/vcFKV+Qycv7FqnPQYsmkIDHSJOT9vOc5xJfNvIbL3gWM2pw1OouCg
kVeKmQQPBwde0UKtHg1h0x6S6VTmS+kVfLZE2jp1Hx31FLAOgAO01EK5bZ1OlfS6
T2HT77QFqfqZuYyQ9PSOK+3TRzmgDUEJ20WGAbZ1Zq9iq/pkhv/3ocIzKByVbxoG
83UZnyF27Xu9FUjUM9PfmmXxZYncyHZPICHD0TnBd6icHnZlxMtNXeeVblGVqtvp
MhDp8E3Z+YKllnZWsKuc9qQJYDBJbcKBLJnGrnwloPi7XEpV+WPfTgIb2wn063ZJ
s8CPDUv01iiv5g9PG3cZW3crCbA95kvSwZvdXJK/gojQgs4YcHOLqzAtSN8hp9yJ
otHUeHP6G5aqz1PkX/i3jHRmlG1HxUv124USC5qJtHtO2FtcXNTs8VurTckWrQH8
eR8UuHYWxUeOvRHF0RCKEBO9l3l14IBtZcH1PlWHvNAaP/npAj0c0wrQWSQm7Tuq
kEajcobOFKA25H+vyTbA1itjJ50huyofo9009GBDm8pUrOq64YRs9zJ1cFD75rtN
6DnddkHzYc2SjJp3DI/ZTFtRGU3NkD+10gkx/rJ397Oxj5bzAIcNZer48f0tnugz
gDAI2uYzDMG5UZG0IqT1uJqlu1VINOkAJfDhA4FFYJ32i1e5hGliSqGS9f7+ji3f
9h53m8YuqISHWRYr/kCxZ7UqA9GlzsRsyjwbTYS0sZXD6ty5UaWijenrZqlhI+Xh
O0WqWjT9m/UQyr8m1oZXXZOccN4B95Jn5lK2Ezv/4ZOsfz4AVkRz3AqcvTCCRUbv
CmZyXLUWvem8cWjJKzQex4sxOaiL2OLaa9ZrEmGAjYsQQhPTGRuU3jPzLAI1+UDx
0C3+4WjvCLqSeWdJreyEYZZL5w8AdDlorXru7mCp8VbhMknw+/Ixr5dDserjZyUC
RqxZE2RdVMrCsfYiF+uNDPMH0ssDb53y5aJuUCbF3Tn/Le4o/ASwUkWQEO8UWSbQ
SyaBfb9sH2rdm9VMZ2Rk+2J9FVaI+rHM3rIwhSvTdHurpXRWiYWCQR7tPXItYx3/
5JYs4Yci2ery1pEhaW293u3jYpMX6J0htMqLXK9cd4qkWKMhP1X0mvW3BkRL+e2Y
jBx76dyoVdFigWpKtpMS8yqOxik6y64iuQAZ5lh5YvvINokge6AlkmElWW5yeh0z
oOFDCkVT5coL4b/+2uDMHOWa0AZKYI4yZoVrT445e6HbQjblznTdeyZuUTRy8CyO
/fFiLWvSkyTQ+3fsZJB9z84JdbcNDLBWucuAHwGKQVPh3cNKqX4GLJkNKX5ljXDI
bzq8KGcSpdgS/yrTbbt6vW2AO2wmeep7mYGowAo6Pok9xKo1cqPZgZUMQlu9lu6h
j2J55m3nwjg3nLHctC2ATJlPLGOpqHINLnBb/F5OsBM6orHeeMyeOakkt/7KFldr
51aJAJ9/9fAtXZ2TopOUf42B779M701ThzWyLWnbFJMooBp32qqQ7drqN3uQRtII
NZSIW7kVBVmHZxE5IvZe7Iq9/NIkzVeNrneV9JTZM8sm2g+wbOmH3h4aLLvo4qEG
QHV4loTB0NoQ3PEqf0dwx1874rLUYCYQ4Le3ZDR9qPhWSTt8Hh24fPGynUFBhgdi
C576GdSa/DZNWYa6Pubi2Ph0AJR4t+0/ZZv/9oyEjZdeRofaeKD/ty0mJ9Bw9v39
m3cflI9FEOYwZV69wgfm9BlVnmg4q1G3MtFpZpxh+SK5+oMvcNHouu8c/X/J1ADs
PY1lqY5k4vtMsX+4AAg+iDHOOHhSeSFJmvFpTJWXsDqGwkqDIIkzZfnrE4BFNBEH
RyMMD7QE+djt4U7p5/N+mF2ZP4bmF4i1BgleRT6PsFVn4kRQMlRUlOD/LMLzgezR
0OdFKg/TOr2OtZXnaZ1U+5E55QJk9rn6yOtsk9bwTL9qbJ8P9nK7QJ/vfcTbmQON
sgY6kbvqXbNg/FH/NdoXl9gP1To6ANRYbsn9q/9zksjN+ixcVvqcdgRtM20Uep/8
Di71eNrgk6tg8VFAZqccvWRCa6I7R3dJsLvjyULqU867Bjxw04p7UsSSkrMVGjcX
RNSuIZkfp2GHm9nrrxwt9klZrGAo1qGsBXaeF4NlMmCpMGCxg+xhDK1QHEdzhQ4l
627wmOu8EGzn2rzSEoJBP9UCxbV4k6Wh1KN3zahWsQSD81V6MNLFXdV5z7qX6tZg
uxMFvCJ3CgLf/xWNFXTkLzhpk5wEkzf1hW29yMRoYyVp6gI5hANgUg861cpFIvce
vaMAp71/EkHGdq7SaWrvyPmYrUtX+c5cjFjGLRk8dEuqYygBPW8XmwKuuBaPgjP4
1TJDXPhF90Nq3dXzBhbmWJUtAzwUkJytoAPYT2ot8wZOxbzog5RcaAwCl7Z7bPN5
h+nHNeaTStHy+xf87z8ndhd7+rNeZszai2RNv/4MDC3IMTtDbt/hIY5g0jNokAha
NOlloBNS62sysC4zDltcSPjDTGt+KfQ0zwvV1VOMszZ7VLr84cyPzBeC8Q9gMqFE
YsKzR7PLLuDge+PYs/fHzqyFRPlmE8hR4vcAOLfnqv6VwXhDYph2Pmq5qbB4yThc
DpGwjkvMwvicygWG6wKQNq43naSC2Js39ML74TNfCxTOAmmpaoSgvYiOYcEF5ksB
ssDu6Y8dn7+Fsv1t8LI/X//GRX82/ZzhxJtqjzEz+rlT4Sn92pmubIDNb7Q9tvSH
9u4VgpBKb42ArgZ4IkEnBlks6vecmJ/nxAysL5Dgvbes1Z5ybfIdxWRS8xcCzKNN
sW8ctkxV3+wD02PAtWGg6rdAswXP7FG8QToO2ee/tdV230udY65tZjpXLlqEP3Bx
Yhpqb4QuqBRRKDphfmJ60oRp1svty/bXyDTJ5kHJAr0+LJyePzqECBVu703uanGE
bz8VY91RJoPxG7PASbJ+Swdni6Vsqag1jIMBiH6QqR+v8KDSAJ8wQY2WjpIouDko
0I6DrMr49Vs5ZVPglFCE+kSBjpp9DPYdFg96iCWAbZyMVAiI1UaGzaAI9H6gAfo9
uK1Fd17WVJGxqi9fiTVi9fanznbKeUEYWpZ5eXmSEC3D8Jw1eoCArWP2uSuComNH
4zlayIfA7ZXzyXpqeiEaaBZf7cntEr5+fj+nELuLlz2qr76S66FSn0+FZ+6T5cOO
PWU0dTrs2oBNnLVOfcgek5fFeTEh1+YX3Hmo1eQgUeC8A323rpSXyY5rP6MIaK5i
oI/a/i/f0LaLDNEp/TGZe4yghtFKeblGXQQv1Wv1HaBPonbAMqZbcsnhJeBRon+9
d3M2enFQY+HpmlcgtoDkdKioML383SBAksTIG7eMu4CtxWVOvvsC/RxOhiGbplKT
TuUTPZaIiZGl76UOKSnVp43gfOiA6Cv2ERZqBcjevxscmX9YhEzh090Wv3AVRz1z
Egq4RTK3pVg+MG8XmB2pqK6A1vIEKNHXzfYIwS7Vra6atPx273lg67U78o5ue40u
SRN5+LGVw2eySJcIHJKkvwq/qSM1/+s6lQFuhmANqFCJF6b4q7bL6TJ2OLi8I9CM
osajq0DSSv2H0CViRCcSLJp355opaoy6Bf7S85V1L2Wh0Opc5UjP82ZEvfoq/vPr
QZ5voqZ9Zpzd/h4wTOK19mMPd3n8J6rOIXs51hAcDhqbDQfy8394M/RsvN3x5jx3
OBxJKASh2uJuJvAHf8+AtU5ZGkM9t/DX3ZwYHZzacLrh9pMDyNu28l4oxMdXjxM0
6IScgTZfAHIuD0ik4xtjW6HOFjpiN5gefkV+vBbkYDQyVbk+h5+ybwdnRZcY7MCp
+uBwJy5ILfaS48KfPeyPRfqWOG97XZJbpAl5oEyYa5dKaDLKVigswlX+mJ6cI3TP
44pkp/QrFLL+JZQwk6YyrAe9nt8b/rf8w1n2iTvVCsIx/KaDB1uu5exCC48X0Uo2
TvJx/bvKNwbaq/qL6+J0ngmXMq9qmpZpQiF15FEMVQGYNB3qTOGPgepojqdukVjn
1cG/CKup2lXljA5iBcMnwz0MY/MDSQo4NlyXMYa3ngnv/7mK1T1lM7sJGwq/Tm0I
Fu+SWKZrXYXDeoqcVUA/qKSLEAAKom4f4IUoArwMUNzFA5rXGEnNjKgwuVJmUWir
jf3IjwkPndChlpXhFLRSzRyV757zisZTerQA+85AXEx4eBWIPJ5xQDaDbBkEL6Tm
I9r9d25CySl8zSbhRvq3GOklayHfZnJFZPkcQ7Fk8HbHD+XJa6Kvp3DBTKR52jhf
S1QIzLf1F1KmdpeFV+rZgyWkpeIZqPA+O37unBoYFfSNELI3STLV5H6fTLTgcfVa
ELH6PP91MwWAUTWJw1rjkmtjziuhu60WAhZJvY0xYpOu3auWog+wzQMYlcihE5z6
KeK8pGJ51C7aKOoqte7nLeFXS5O7g2cMzyd+6R5F7rdJcUL0nXNf/s8aKuTbOJR7
UsQIYjUT9uNOYX+Mf6SOwIq3jOBPKkT0I4Zao/mRlyewG2KsYu7H3fRIGHGVEePH
eXZfEyn3dZkjPkHkP1NXpas7WkFjA0WDafMfW78mxhnCGgwzQgX/AbkA9phfs3oV
PyRy9JMOsvSt1rHi1nDEm0SZX68HjgycP+CM0iBI6xmf5ZdpPFfqEaziv3kgqEr1
NwPVIRfNXu7rUS40TDxp6e64sMFT9e8VF6tiLcgm7EqovQ5tsCPGsv8B1oMIofvW
2r7ddAU/Bz9yRFtJpXtozTGAT4ih8Uly1DER8ekZbQoEr6G7PB2L8Qunfga53ejf
zW4+yvGjhSoE9UjsDPJ2DnutRApF2VQ1cV9Mw6wJ4P1MAPtk+YoDsLmAmdh3uLwN
3thg9Hic6CWgyUOQsk1j0ndA5A5HopSg2mpaGoinZd1TjaCz8uBYrEUVDaqYswHM
9fv3hgDmk9JuZRZ48F/LJUztp8XksjiAUCwg8bM8priL/5WoJCUmvCv4gge2Z9dg
BW/nvVj20UUau4hDLhK6urRwxh0+NuOyWl2MQogh/0U+9eyw02jsSaLbO4Mdt5M+
YVVPU9erX1kGpjzteFipxEZ9KK5wBvif05FVWjTJE7ZTJ3MvFpcV92z/RKo8BMFP
CH/3w3kw4SruF4j5LVFCzrJpa4j6ZpHI8/KtwaYISWwYYiPJhAxHRES7hjOuDj1p
fuNIe9nvJsdfUgeUzfb9F7l7FcV4TWGvLyAPS+enmBaNfDRPAuSB/K7E2zmPriv/
VBdoEt4UmLFAnYU0GESW3dF3tkh5S+cLDRlRIqN+LZEv21Ocj69zngthwmN1iTv5
zngFxalR6rCYqKwCFXclEZOAY3QpliN62V4nK3Wia3uqm1fuEuBx6GIQYNErMS84
qETtrQi1rv/7vjHlkeEK/YV3mRCKHdDqe+ucI2uJMSuI8YmK1fS1Hb83BmEUphCl
5pwp+EeC8z9NieLq8OW1WVFxrWbqIdsr5MJweXPbie+zdT4q/dqm7FNRXRWprXwD
i8jcC2DZberzWTxzR9xI9FjOc81wNby50+YVda0a+eYEFz1ZZoxKYAiIxpJamzHd
W19voZ4pr+R9k79QH7sSrsWFcvfN/tCYK8TdfRBGCpyGj4a0d/BmZVlh1NBNX/Aj
TGQuoD6n2lwwf2eqDuTrR35pr33N49VeQCX56K9TO8mYlX4DpaJE9+vy/Ji0IVuG
dY0xJKgl8ZMPWxyp1wLGgffWy2v8m/dmcUQuT5A8rcmRiL+KD5w07u4p+c0SuhDS
TaWpUJRqRtOpbQP2/KrbK/LLOXTCiOHkry6f77Vt/MJLvERtqigVMnuHeTKXK4c1
0GzvIGyl8qfesUL2Pe1jtwhOrylph4xia9Q/247PVez/HM9LOhMkddXil/O+57OX
gvijnteS0f4wQc8f78qoMPpyC6bG1w08PJ7yb34F5RnBfj6WMe2LXuDCZ9Q3MrnM
xeSY5ZH0XKYUBuVQuVUlTo6/LDODoOFKV9IDpnBiY2dC1nZ0IjJ6RQ/r7P2iSqfs
L62Ym4l4XDq3axQs33Rsj/6NA2jBxgv8/1S3ntvLZesp3xqz10SpqmnlW0gGDEsR
+6BBHWAxAwhioJuNGlRLYLGPoB6tkL1mTiXcAT204+FMsGrmTc+sMd5P28Fi/YZa
w+rGp3n4IpcTWmSM0lW/e3BYIsPLu+SEPjGkiBLoJH9QqY8fTaDmH0+8knjzX1OE
ENXsNYkfBYRbz3X+dLqd+9VaV1afeGKllfCI07C4EajgAtbsKSlJ2jMapvCbvYBr
Seu/LzvZ8RwjrCaZ/bspp/lTGEt8pmdpFLTaeg1925srAmhEpWg4nDT4mTw70hxF
rgVXgBTrTSnigslnM+elb1cpF6aAljmAJWS2uIWYGTV85dioJrx/yy9RRSQp+gLG
rg2+hAj8NyRiBwBYxbgZfACQPoF4qmGLMTmC+nKj6PPxtAFbmIgrGGWBgxxQ5HSc
YkFmjC+VJ5O53bh3Q87ZHfXEt3DnK8E7JIfV1K3lgqGrbGCM9OmvadufXPTHGBHk
ErMFlcGoIYY4DrDDlYL5rSPxAafo+pYgrGsGL3z6NilYONpjwyP3zIaHJWyo8ssS
HbCLqSaxKFWiTh87/sfy3XI+4Og8ht1+wzOHnHxidX1pyR97QtETg6cyPlL90YJL
/PQSopb/hJDiFTe+MYdFA3l4fKs4epnfx0hrV3TgJjZQ543fyo5DvrGIpNMLbO+u
I8kLwp0t8jGesKVzOpAPupm5hwP7IykWUkbyFsgTGs9kUvsdpeeto07Na+3UBEsL
KjRui3N64CHr0RNQdTGQhE114v30mLU6TxgQoA0k4e89+mVyxW2fX7jcw8tlKfWb
e535KZBtaPr/cK4MHSzqv3C2tg5OfX0bBPAcqtNU6jiCXbTa6g8FtgQy9WSfyYqv
g7vlRnyvXT53SDYdfoiNweXzAIdNiOM5Ni1S8CY/K48etNwUqQQ4qFecGc6ex8Du
VXhWczpuTT1fwu6Zq+/FX8jOV2eF9ud2xzm4hy4crxbNlrQz0sClDtfZykKlvWl0
uN6nXq18UUFM9lC/mox5YL1siUmXFA68LBN0w8ubhEh7b4n1E/j6a2R6TVfxPJxl
hdasDeXqQU3mrE0OJ/iVy7Ryk8vIIzfeXZppK+3lsn4dWKoAA4dH47Mf8ztZmXi6
UYtmkxyMUoIHQvCt186OEuY/0u682vYA0xOfWGYxhHcjsPiqMLVWEXKCjGqfqpIE
78sKGVo9loFf5duYfjuIFj/WopHQ8aqSN/B1Pynhr38kKsBE3FGJpB1g/KllEHiD
XWLC+8zjM4MQOrc9RfnVyQQp0qZpPgOZK2I9nHy8C0pWJ5wsJK2ZCJhpMbbWCsvH
bblJUXVeOdAIlFAavWs7aJQKpRchCkuX5bXej9bqRjHSCrqOhyi/lUSsHNyp1CPe
foIPM+zbc2+YN/Msrwpq3JdGykMHvtnSpwu2T6CPiflxa32leLZF4SCyDphLSXrV
jnQybqM6/neqSensFzqsUPjIbDaMaYLEVYxwUGk1wFQ2fmfP6EJHc2suwRveZ0Dd
Vr5T0a+4Xepb6vThJaNKSq/APwOIPwlzZOWX3eeUt84Adq5cjZUUFW5m9ENXj5lv
8/1HiXgJVZSqAd1neZW5rugSF3IFVmSHJF1UU24z8grSialeIxtavnenfnvU/ZyK
VVaKcDfBxR7dPH1/XbADAGnFVPc4OOtbL88sQvteefCLjYlRRJKQb4dWZ7igSNDo
40QsT8YzX8K9HFoswoIpPxAN9DzNeLjrX+HKK+Nka9okOV52kLQnjujUJtuIH3r2
ppxhTzCZEJJVo4sPLDV8+KpamkAIkPp6QFSXhnM4BgT86bRTOVDn9+sbUM+65t3z
OxgWr20K5KOaxfmGsUu3rXX1+mW0TEBtFZOWLldd2KEISdnLxMAz/H3rODivooon
yBjwjFJsl+UXWsuOQfrGNEOKgjSNr66/F++SCtEPV2C3bbQU8+2AGwLD5RrfsNed
YhPyKas3dJQobqMCyaOsei3Nba319PjsMVyIuO8bj1e3qkQ9O4v0vEvfPdtznlhi
qaDJ8lzvWem3bCqVnyaX7R/A8VVnrfrZEKZPLD+gfQaiItYLXXoyun5/YUnpZBQ/
gsbnimjfKHPbIf8utz5MVL/xG5Ko1ZlaeCArtdwuYqUtBn3MHT/9YlSyaVfYj9pJ
tOFmfeduZtOVt5CmNfvgRYm9tG5LLyDU50k4BCUT/GolmAnkfuIiR8ZES0icn/TS
ImgTN8lex+7thF1V85ctFjXXGQ1i/X6cjzLwNojjd1H5EMi4XCH/3stGy1jOvMZS
Pq+iQrTb610WXvJloHU1S1MKOTK3LyTjdI61p4VepFrNIcghlX1pUTmXOq603YPK
VskeKx1zGkFlTwQvmc55orq4PZ/XSZ1f4oqE5qc4+To3ajlOteS5d0JwfIxjkEto
S9KebBiN6XQRWoHpP2wgXLb4BPgW9CzglDHJIxLHj7EjQjTggSrBVvxl/XGiGTLY
dnyFOeBKnyhsishWTVtUR04p9Lq4qAOFRlqQ5i6NCwm2DSm0xHwv6uRIE9UAw0Rc
QxyB8uOhOJcgZP7fDxSsxwWyE6zLIW5ZDfFEKfsq6zAS4UTdK/tZQGvyPUxtrXUB
0n2srcjb4HNeBcsDUs8+RNzO0HKlCnzkc5UZ9imRTGlwJIcHImOQ1XK1hmCJYl0l
08ymVknTeMDw/5odGJYL9vxmcRUuzY6XRODpUnkSIor3gcRNLM6IHgLgA2R1eVvF
DW7NaXqB6ij4r127hkS9qB38LqgsaVH0Dri9UEu/Rc0bchpmK1RNf4p7Ev5Zg6Kg
TYF1tgJCdcB5T/XsT2FX0JcL3IpvZAjWbC2gFO0TcNFukMM4iVlt+PkbpljYBF68
pLluM8haAjAxafjOEeBI6ArIyyd2unEy0W7Gtt5msRjPznGSdyZQhsVLZ31Bm/N9
izfFxNS0V49heQiT6hnFn3+rQfXVM+hHszJqEbEckK2LkpNw1V6pWCACpNbk/HH7
XP9jycp683Np2QrH/3Y2sy3MbuqIA5L4xjIPSlS7BO3qnMMsPjWQ6/NR+hR2EBbK
Y8Tj3hHYv6jy8kiffKeBiDeV3cqeRjJvJQJ03JKarhFky4/niGELFMGKZPExzZDP
KtvWbP8n5joAGLe+RQYMAWsr3Tt76gIFaf+e/m3Zne4J377/XGe3bFctttUHIful
xLJN1U44Yn19mnLb8MTAGEUs5wYEL1pcT7XjQYCtl4TW4OWkJ0nFbrvoS9ZlwnZt
Zm1SwFvFxRj/u/J/DE5Gp1c2EwSjjZhyajqXJinMtjdxlqK9Ca+eHgDhyXbA7b9H
yafpEeW8UO37DB29pFMBwTLdn1lRvIsvou9Sd4LsVLCScX+YZ4zBXLLdUepvBdS2
pEV9RWXcUmmdc9gjrKGOw8vfR6dVNY9hmp33r6hkIOYnE70Oz2EAtVmdzMaIlqAb
dFSda96azw3d/BXu8Kw5V9gl3UtQmYfnh2obCsBbi9rsmI0Xcu5HgRKbaa8GgA9M
JIHlF2P/0e34cQESVQxTZkRtwwqhQpuBvYzgxyB6iakJEWRa09wv4W3HuXEd2AbH
3tzy3kkrOWv1YO0GOvRRj6wVHvxaGoR3B8i1BZ9aJaB22nTZxATVg/2cx5pTroox
3ItvqU9JHFpvHtHV4oTHnePzuZGlYWRioCP71ag6u3/dWjlydiTr7XkYwVYb0/Y9
x0K2lk8eY6dan58aCtovRG5EG5s1/DhL/skxgAZh6I9w2/ZcPyPoTmqyfWWWLdoL
XXHz81q20wmUoXRqgGApGbLgrsW8N+0Ht0YHVl5H/nKy+RUdWk7vdssyK9RLWD/M
T/S/ABc1WVLmQwNSOEITeMliEHA53jaMcw1yyS2+gpSIt/9o6cEcP+LIJjc/GSuM
4xpZNLujS2YLY7vTbPGsRHPeCsmVYBzkD2kCZ82Rx9CzwSSRfV2zs/IB7BqwbO/O
7SuUolWGCPO1YlQWUNVjF2bieqULoGucLn3Fyhfr9AshsKVhPZlSKZPzEIKJ5Bbb
jUsZz/ltlCha2CeNFYDb9jX+Aebhq2J78+16LrgpAXvVOSbE8wIcr0Q8j/60Bp0N
7UjiXAweaMZH7ox39OXGsAizV/EfGg4TnhYL3Roup0HdoAF04j8w4lGPDj+8pbdJ
ik5/NEUKUStU3yp5LFLWZpB//cbwYQUuMG2wn04kMFZzzgWlrF7GL+34J9NRJFwA
HwCwtQeEcZzmV7a+URxGTqlfgdoaWZqTShZpGSvU4BcJC4xwPueIR03dorSFTRfY
Ril0KioFU9jxvL/cq4LCCsb5CwH9sPzN1CthFdzrYkmvgFtiTV8/krEf61tI3Xla
IC9pe36OcwphqBSJUBPLBD6AY1U6cZ77+uQLjDzmt3f3mddqxxmxSWud6G3lvhRY
2iOGaFxvVhv5AiVB40K3G/UJ3r2diMcWWbOm9WLiBoy0UFSbswihhbTqojWpWeyY
e2u9n3zDZ9fGceZMc0HJNn8PiiNkYUhyw6zOQFVMJcMOfwIo9yBgAdO6GU9A2Ave
Mf4GkYrJwW1y8auN0FF01HqpL7huj7CBxKK3rno9Tp0nqEv/2FVz5I37kLsJ23CI
ZgBM16bC9UzNhMkMY8lu/WI+ohy9LOLN4EByEFth0/RQZMxtJTaw5tneqZGEzm6r
0qxRg3a7/J9zLS2x92FB3ZztvH9PXoQelSb9ah5jm5ype2LEzttq193ddjKrmxpl
cZgh9aRl1hxQawLMfBtjbjLJo22S7phmedgkzgXM04HjctsPAVgcJq1l1qQmgcld
cx5rOnMfRIuMVBFvS0z4kgogjiWidiQWkjBIumAa5c4zGMYQ5M8T8X05UOWSe138
DezBSBSovSQvSQIcogAs1noxZ8YTKLwtS+2kaHgXEwfEsrzZ76kTZqXU6VgWbIY9
vWjDKsJQ9QK43MjS5BreWP+jH5qGi9nPPYVTzdvgQr9L8JGeysA07Nu2nxQnJMt3
p3IorffIWwCeCebuwhCE2LysVm3qWP1u+6BT16S7GYFA+mvr+oJ2saJfM4GAY4g6
YaSJeRsZORN+AaYi0SJgjme/xuzGoEOwQ3pYwx7McpB+FYbDnMPaBTEYnOBjg3jF
Xy44Ujq2jkWt3PVx+kQ1pIKtHqGsjmjJiSRVITtrRwGgcrb70ZHeAU9bs4RXo2r5
hxT7Olo4opfWAh+sOx49tYZFdLqKAkr7PEtEF051Brjk2KmQ27EHr9LJ1/V95GqO
2uuXSZq0iiGv4Zvqq/tAtsJZ0EVZSHJ6Z20lxtAs/qGzudaKpQD4yj6n+ZqjwIOi
rLa9ylgywFoAWDXWW+VYTODfNiJG3pvmRVJHT5reUYMRFmEE9stMLuPKkKCTfDVk
WEx9IX4us8jDpdWYHRyMODBPr0Dw9A7QFwB9nXlPvXNAUJa/kYx3EmkS5814ebRO
KbxiOFHu9sjydYoOkU5/UeDUbI/S0ukZH4Xa5rfS6xVnMRsr/KN7gmf//J8ym8xK
4Veu8mFtZ/m6uApJIw40Lsrb0OLn6Eo6B+wVFzIUo8JMWIw3x09tT/PWiuyfGrAL
Nx0Xj4bJyCRjUH3knvS4ZbQLQxy/pj6l51eiK+WauAm3y+NB/qFZbcq0gs2ng+yu
zWnzc/ekETYJlh0kE9GYykgdpf8RUlKzFMmhAX2duvJCdm3VciB4i37dYb+1HRJ6
+NgkTZI7jEu0EbnJI5MQpuCZlvFNtpISnGEU/qwX7sltuMDkU6D1PUc3Uh2JPv+U
dKe9CjOFu+T8djxHXPLnKTOqN7fsvvpCDUI6dJZZCWear+3aMyf4TTQcQ0GbLzvv
9M2r7oxsSz9QguYqQxcWczQ5+Cj4jWekperSOJzz6c7pB+qml7B5buiW4owUwKUk
0aYoIsDJso2kzRrDHbWl7+6/Wk2OZ5s6t4xJwH3cXxrpTUBfxlNiS0S346Omh2ai
dtuiB7Q/uxyAg/WhzYt6CBNsmcOB5Cqc03rMvBSNNT50W+E4iA+5pVbobcrz9R19
rbrypcbFBlBxKybb5J5qx+QJbAx1NVQkA7RHUdYFh/gOuP57OU9y2VGVXDNIR4Sf
FOtuPJnqvUCLSYfcB7Vcimx9q7ReYYiDRWLEdA9Ru4aJ/Qn4pEMZxZwHo+WpS7Th
CILbAG+4Haf7yH4ZaC0KqycVRxjudAES/lylYcdSBVhCr6/6TO2k3LdugJhTdi8X
9GVt2kCiGzbPJCLrFStXaG8CZWoWlTZ5nUqtwY0RVP9cGQLOPq1+r8WAPymOJlte
s5odFBTwRgsaYSh+WAQeYCsaNKJ21tvjM8ebS7G3Ppi5hoCCT5dkaPyzxjmGmncZ
dQkv17fXMB/PoIAPt+KXuF3z4E8D8u+m5ZKrfgvLUldy7qE41wXct7KliuJOuElV
4bQMmgBypsO1h76689sq93D7iylYC5+XCCgrnSVcZp4YN0HTLur4MfhmgWxvl6Y/
f0I65nL2owQEt5YYeKPX+zFxICqm3xL4jMvW8ZOAD7JSjYpPNeD91IzsIMhb739i
3lt5u//wR9TDuIH1c2paqGtiAj+zNQdSXoGAXpkO6BiLFFa9eiM/dYVvjzdOAMMy
xMQS/xeLqOzwGn/tOwpW2sK+tnj+2T3f9Khb3PnB0Sn0+b6oRuy70yfjfgyyApeo
XkR106DoRTTTghQ8n9dWNiiaUzb/gcZKI0oA7Xlsc7v8PoBH/Ma5O1QTJJsU3ASc
TPEFCuESS6nhY2Y8QLSUGmayD9lBPONmITEyuOd2XkWNFHcfRS2dufcyMo5Pzase
ZxczXJhxEnC/lnQ09tQU6nhU/YDDGKpNA9zEz1SX6hpoNMu4jhX3p6MXfXVODHDa
hvfgqupqSJoM4KdEm0DUUsuEyZgQFkxaeVi2w51M3mVLQl0YtmsBtoVtXJi4Vzp3
KGW61I4iw/tBdFb6IwdcqTtFNHcta1XEpwRC4pdtl+9MtJiJUENWnId5zblQBT4f
RMCntESvGgFTzJSRD8cdR8AxEXU6hS+krIY1WUTt/Irew09iBc+baJjOpjGOKVYx
ZrgIyguRMjWC6vZLnCl2tY05WbwhmlqIGjMutScIaIH7wU226wyiXnX9CzvaUUma
oYBkWD7rxKIUNPeeaw6biOciRjYpK0UwsdY4l02vQ4OzOdxpE2PWlT2SanJLpoSg
4alDZJRKRFh0oMXhdWhI9TySzCotGYSC49RTRjIqbpahW9JMBHDiU45uVzmUnQHK
fshQEpDQKo69lGqushz46d7xVQMY9xAEoho98213EDdueDrr3Ulr6Y/HusNyIc4J
LhER2tdr+8IbNOjxMOd01Lbzyesq1ubCBo1Ncw5JFgzyWyKWj7qjzL8stLV9fUqt
lat/6v7s5h/RSghAlw0eRvvc6Apbyu/Xz9lWHR33iQIHp05G4tQYIpIZcijlf1R7
O2pcJMNknNi7UzUMr1UVCL8yfPtqLz0m+MGi7iF8mx908Qx2SHLQNG8zFbgS6JXt
IXAE7w3CQgozvYi63QXvN8cLp0ZPA962RxTrGrSJekbKViV07TJQXrqJkB3fDsCq
Lvh+nv7Z8bPzxj7AfG0RwPwBh0zYfy4wfxpSBGm3bB7rSucLIfbqjH9l0B4+9dYI
1zSgGIjIG/GKMUhzaA3lIAxMf4J6SLYaRnbwpV+s1qpedYRMH21vl+uTKQmG/KzA
M0F7bwWW1I/xMlUOUNL1mnUUmMgfzkiB6Jhk59VfsSFX2L6rcNmN0qott/tSMVqg
l/ZezxFIKl0k1PFlj4veggzfLbp9Pyr/kmSO0++2EUMo9DDsPajo/e4wUoHLffFu
2IYVJG84zvAnU8ewKlryvNrFSMMGt50Evsqxv86lhWtm9oI6Bnd7w4mFcqhulYri
R6Dmh4HlHD8AxH9w/8Zm4yArTBK8e6OvPOWES7TNcwdOA69wiXYWuD1x4l12rMWT
fDvERAxXaEF24Q9GhX80jmS7Uc7GG8g8cYrF5/EnyhNrT7yQdxTmUcXX0ZqgsomS
40GSg7s+B0WscYR6W2y5fCoZldJNfjWUo0Mtooenxmmqm/ZKTOsddDKvAGfU44Nr
xb3vwQkhkICPVeYorZRdYVjTA0aXmMJDdzqMxmSSVqDBsNx2+E4PgFrIaMI8kRuO
BK+oQxNKrXsKF4KwfKDB41PtOwyYV9zj3nSzaOIdgiU625Z7NqPe/nsA2Kki0VQX
R7Y/vNL+HQJV7TeR/V60M5zCElC3+mJ5THHSpFL73AVd7lgxRXKL7JTJmiaBTGsy
syq9NVykwUr1bCya0+Ha6TjPTJuU2Z47eGC4c3WFbwafF0VRfaev64ilThjyzw1o
x5FKRa45rOxcbfTQUVvCZ2cXFBc/K3liZ27uLXuTfvAOD9Hu0LNeUdRxQEcBY2q2
mqsSLfWA/pLbog5M9ZYnlbUMb51t8pK0UxwBWQ8CnGhq7p20RGdhofVfJmh0IOME
EPJjFtZbqftFprAX2Kxu0dZnSZ2yyAEberXA49x94QDzSZkQeamICustsSUwdqxD
lEsKBOr53tNrKNz3JKci/9Z0zaeHSEtPr7m0jHo9AKVDUZMSUfnYo2aUFp3nv9A6
iT/G82rsbAMUnLSmEvDHEDHAXtbfExySpr8+fFYLiAe7DvloIBjqhUHLb7dP2jPP
gRdtLBLYQwbLyKczahyD9a7CLL23hLj9v4W1gucJbJUoLtk0bDbBZTcGLWLgAdXd
vUq8zlZ7zqxRQecPNZw01AUmpGxhTYAbp/RJ1YvtBeqwr3to7RlVaBhAZZDRfQ9k
qvDZbhpoXvXbljxogUOh4W8jvLhoQftufwZDIPQEvA4zw7xQZt+pf+xYYFgDSfyE
so7FZt35L3O0EsB20IjMjrRP3AGEdmXnlQ++xInWB54iKEW7OrJ5M6JkB+tj06RT
DrLE+0YHFmLQslut719XlyebbcmwiTSYVE7zB/8TybovA9JwYnbHhAv5Tf+juqlf
7qCO9rz93BLMctaO7/fp2bs8r9KUQeCbppcNU42nuDSPNBdXdwIi8Od8yruybyc6
x+SrOxkUPVoWknVhSusrvkCuU7UqQjeVTsUKBUbUHtBl+jcLPDhnrQ9BdrG+JKvc
xF6A4setzEI4t/HxotB5hkE9v8mPUJnoDPeULwUovBs+a1RPLImrEu/Nm4RRRp2r
x/i4TqUuDYJyw8PmH09XvPo5wqgYI61g2tIQJ8MeO2ZntTan7x9dI1fSqCCk46dM
4zUkApldjHM5RhkOzisAqWf96AUiRi8sufHeGXPpIvUf6zIIiGLzeNgBy9QiDhgz
hQoOoxYEhv5NhOiMOVxxc6ldHKE31JWhUiPICXpc5BydgBbLwWqujN6om2JjETlj
OdAZgFX00WtvcwuGsoXhDS/R9/YVrWvkW28eveXlugm0EftKDffagaQM5Vns+yf2
MuqlkzVe0zwGAIagxMeqjljocEZ1DoU7VVXcEau0+cjhPj1C/FJULE/JTRyEUSKR
p3WrmmutvRAHqfan3rayAf+JIAOUc0ByR1f+vfHHqJgpy81GIPFrfPSVr1QsAE9w
sMsqZK7JeihPlLJqVu1ZqdQIcs1kPBNjdDjJSOVgyhlm9rbBWab0O6phOCk3/7cM
h60UVmnm0HyX/mrlISBbJhSMeFVxa90zn7+0+42EGOAb7P7/vb2iLKXfMdw1kQZg
6p7ANTEYejiCdZEkTMfvVGaJc998phSqQSyVCigUNHQ5XKtl9i69Xw/IJr2wPDwg
PC0z+guaggRVnAphip1SiVT6X+/Kf0k898znkDguZKVP/PGYvX998iILg/bDnC8y
spkW0bmRBPpfv8C4WcI7vNGoCjREsbr7untnUuTTHeF06mmD35JPKh+16aeO7mWR
10Hf9TqknS3E87OQIdGVgSsFW8md9GB42aos+WgCK3V50av+M1fvlmS6Ci443cy6
UzzpUlNjAm5xtd9xehcITsFwGN10nrzHbQXlKtzwaUtUWOsHDFs+0NUGF0ssM+7w
D2XbUaN70Ip0AwSicKVbctLDJE+60PgdrDMXdFgMi2/ApsUlR9oxSpfr/vgspSOr
1h3bVIqZ+9NwJnBYhpPWlso4MAkzlZd5Hz2kdsC/m5WTIqVKa9jXdZfxd7lOjXfD
lvfE5H7wl5N314UTe9Xqe9eRg9XedOkFhwGgPqRQpjKHw1dEm2qMZumGgxqa1/Gm
1I8OhTOCbPjGM2hoqcE0vHnnT4QfcVx7KxGJUzERmnEnGKlui245v3od9hah7oDs
Q7M7/aDah3nUuuUUxaoS6ElbzQvaXYCTXEJZ4zAa3drjO4mx4cexSOvYY6dyuX6e
76Swbt+lsYsRmeHkQEoapXS7mx7R+eg1KVbgiRw66KTl3Zv9ZIm4/oQNPlz4R/sq
RPh1MakscT31JTgPoUNJEZVbtPYslTRGo6jXZTlN/5x/7HinW+wro+8ThftCrA9R
0vyxnu89KIuQj/MjGCxDVEdBjUqVWMuZwUL4cpscqWFtUFI/EqrlFOy2q+VRioEW
5ibD14Fb2bn0k30xy9ZYcg/YNpe/Vl0At3MjhukXjN7vUd36vepnP16myJ8DkeH9
ARkKXYtIUa4gyKRc11RNH79RO3G5U0N0L6/SghMoL/OZ/iUhpHqOLMxW6eKM8kzz
HuQgx51Nqi2roOyFuM8+sUuIpVHJ1v2tjh1VAC404OTXAKcoPp43SIJHLBDtXLnN
t1c1V0r1n8vODbqiMOuRYfMaUatj3CTYL0R1P4D0n9ufJhE8fM16ERbqFwZZaZW4
KGh0p7LJv9FsZSROwF1ph8CQwhw5gqbv7Mi60pazDX19BUn7NZfmpYu6yK9cOAj6
MctiM3btcv3hr9fGURMBiHwBXxiVJy7VA3LxgWLKtyADG52zy4RjEBxviDW8D4k7
Oh2y9s2VQZxzBWm4LbC+ibX1Xi96IVUJtrdOkp++BVIKCj0K8kYm4DOhYfs18QP5
e4aYcSt5ZR+XsVBdONET858QY2XtDs9qZScGI6yJgnqLbxhLN8bGjPfbLBirB4fs
qiM5aEPL1yxutkvs5BcBWqwjkHflUwmuV2QZqjnKnVjZe6BezmNbeI16bgSgyc0W
KTH7EePlVcktamrqsJNUUtjgsmgpcadG4Ms9R80WOPj+WUqDSdRCRpGn71hq6N9u
+sOcVBcSMQhN/tI//R5OpH7Tf5ey81jwH8HtWp0cMxqOv9iqTbZRvmm01kgV95ao
tE9/BIxis3cIylLJj4zOTZHhRT6Y1tBlULVkBpBNJwych37uNvuJVY1UMGaChpkh
VU4eQRN9DvpPbMG9fZpuEmCjBFhkP7JEjdsXoQJAxDR6jaaKQDMF/RMSB8HmGcqJ
Jr9bWdhlL8wPk2HDa1bSWrUaVuaCny7drLcHB/+hu0yam+tqXw3tEbQvpfDrRShy
gZJpzwdcI0LHxcmFieVF1k2jvQmz6mJN6EJe4nLktTPX+3g1KzPFLK15kLpoSjc7
44b84AMObcOxUeMJDozrhsSGiiG7XatD+WF/xjV3uEvuA9BzHOQQVCGl9Vi0dIhP
SvY/eooVjHggeC9TwjH8bSTs+R1nS572uicmpClFVMu+8yLIUKtqzD31GCjKdUTj
F9spwCOqOAyJCTCh5B+g0jZYBm++5vbaHznYd49Wn1kGeoDlDuFeG5OycOVgqgi/
yKQQZkhtcLVZb4xK6biGLArT005WDkiUSN97xH9e0xM5mazjKEsVAhvzslHwqgv+
CAzt7TFBLSvJfivAJQUQpbj5AA+yBUNvZ5sUqbKFhesFMNz/jqLKoVDGjjKHbhwV
+pSDuGhjXX3RtOCf49mrN6JJQeD7/NyBQCHgAI5HNS0sH9PdOZFN6nrE54z+BPl3
tY9cOjQPVbAeAippZYk0F8bkT9uYV4JcQk7WjJNSJldNxBlBgqy1e+19Nd8VabCG
pDRP58Dbzxmqai51xQuO/jESvFp1u8gBCjTbZhIuiT/+bRzpECp6PtBWJDL6nY+I
nBj5i/ftWNEIOlDh0HGAWtrmaOoKXW3sZrqOzhAAZ6vjAA94n0LoGAcYZDn4ajYH
pqATcZp3RdHsAUBJgX29iat9ejMjvR7BempUzh4QyY3N2MtKJlmpXV882vOIGmDI
HB86uNxRPj1AdUZATkpAsCc+Qsst3z9Ohk9yrSeZuoyMK5DcaXJHthBvlAB/r7XL
HI9r3CQCLgh/x7Bp1nyHc0Nduq2K+Ko8ZV4Y7MnMH3M3hOkFlW3wQKgEg8r8p7Bg
HvxxTv8kWY6LfW/pytUDIxz8VqMcyJe6hZnDXnyKnzlNvDnXjFyM2o8HWrxNuj5T
I84NGAP1qJ4iDzbjJ/cPG0zkwUvaDpZjTr/h3OuOpqkfzjvUZt+b6BiwiwxB/Pj4
cn7aX7SAnrJnsRGpdWsAcfCtqCqwpBGv44aJxi1egviY/Aa2cdyDxAuaZh+Krdov
oeBdzw6CTOWD79Xdh6W7gvyy/QAwT/yGIVnFGwUxs3/XmzhG460uMiFUu6CL4PXT
ilk5k1wyLihbL7YvNjXkZ3Fx7UwiT8fnpK60HJoRAKfAj9rg020RCB2y24tjFrT5
qTG4nvFLex0oSaG5xDOgz4OjW91Q/QJziSwoRe93vy5fAt1lrr2bPWc6sOPpK3np
i26VyPzQTOkZ07qgMHPBXb+4CZcdKLcl/m+Cc0bWG1wOEX4Xhl408k89mzKFussU
WHHpknfrUHR4ZdwqL2R81se1+zVNL/1PhJ9UiEjHyVIoOLLMubLqL3T9pDGZZwLR
T/5Ncj/+27Dd380352ftIjnUM3zDr+XGlO7vRovUtB7UDQYjjW3UGlmVRB8xkUe4
CbIaa6Icz/7qEagV0MpUviLYj0/KpE30EQUT98bwSY57vJQRKr/0UbpIuQPrKYoq
ofOru6M3+ltMHd05+cMRxdM0CqHZThrZFlsPIhPF7IFymwfwjUPAbfv/LUjiXbsx
UH/inu9SDiL9UOtEwlt4fulsm/urHwCwbpypG/I900vERpvBY8JndvcucUbSU4wQ
0yIusd1W1ZwrRMtfpUaVTm4ztHBdzAjij3UOcj8lKiK8iyaa6xGvD4gJQ55i7OB1
ZIMJyQ/Hae6eDWWsFb8UEc5eyP6q3DYNWufO1XUTKd0eJPWOSC/WLS++OhDaJIW1
JM/INMNZMybDpc0+wNP8VyEjYLlW0XyAolnu1ifZBdFlhF+qt5W1bfoqLd/KaZ9y
DL8zlKoZ6poets2zu7flYO+cjxxPOMCn/yDXGma4+GHlkWTrwzO+uWN7hSbh9MPT
B4imSST3leEErKBbuG1mYBouRhTg9KUL4CCCoNIIxiSa2+5wKcRTbTiaoswoOCEO
TUK391AW0LzukNsteGIArbZ5PUmEphSC5Z/FCTBuq5rluOErg2cX6HjITS7wM+Pe
T6RH5zgWV53G1sSftslbBY35CNauj/QQVvpc5fB5z5j46TqRZ2k4MlgJozDrImYi
+JPCEhilmGVKXYrymHmpYA8EkkjUNLFSivSArC/7j1rQ7G0J08aJQx6ldA/lroSt
+9av8VZdE1ngrcaa2xPF/3OkOjLTKk1aqsRq57gKIfCu/9Hj4gzM6hZw9v17OYjZ
z1PIn3+WdMboaE4SdB1LNW3TXpmOs83l35621LjQYK+hy43Q0fI3qZU3prU52V9P
tQZcpmxRSy4wTJFhl1qWh6vX7h3l+R2QG8FCM0cZrhTO3t/rv3o1H2C1akM8u+ZL
PJ8M8mUojgeMt/9YDe0Q6jEv0sc4WliN8Pf6KRuMos8/Cmc4G3mcpIxsjT+8C85R
Rh0Zsi+8egWaW9O47HdGcTUNDawpZ8YDLzBk3KgrASE1UDb95sqid0RO29uXLsO2
IKvtm8ne8Cq56RhvSm/tWFcLHjtCdXgbhQxNj+YPL5dMshvhCucESjJ50xe26S8+
lRqh6nEWs0GWN2Q7xOH+9P8h1fHtiyqGJgGl3/D6uFUwhGwj44lDWLQrO/YlCM2r
FUEVo3oo9AME7FHx0GsLkyYJ01LW0FiI3kSpL23JGUoaTfsXPBGyot4Y0JgVMBzJ
bf6trtZhjBjpP5RB26eXgR2f4Fxmk6PrHEyxvZe9yXg4d5BlgkuDZR6vPCMk5QUJ
PEV+EylfV+PPn1PLx8urB+xjZbuoFZD1iff2hXpkWMPk6m+sdFgjRDe+2vugFK0p
Vili0daKCgrPMMKE4G36Tf2o+/UTJqsmKb8bYZg9XVOuFHH897lXe42RTmexJISC
ZVcSYQLXFlUP1OKGn3846YIhHOSqQmfw3+Nbehi6/ORFXVRc6beyNwAR0K9doiEL
NnjD0ResJnQXa6hv1elvg+NddKCcHWjk1uCweS7C5+ODrO82G+002uaEfDFnBbyy
e8w3m7QuLTtaM4Htct6jduGCD6hFLveeJEZ42tup6kaPNQB/zPi3fPpBnS4leezs
Qk4WJ4ILqCeiHS7ljrap2Kb9Wl/5fee0xmzrnvca5Bhe6T/SIkHrvqBzAbN6Ks/A
NIQP3r57Vw9FqRdfcRA8JntnO0tkTmsVidM80ECcVt5limioI2HOFEJXiS2b+M3O
y0lwBoNq3o+idrvVrQadUMTv4vSNd4/W5InFHqubRadCO+6iY1eyp/B2M/SMMpig
P0UqSGvFqUgL2JXyfyqdp+293SRKNYzM4yhXRym8L0ZRhiAcqQIpPFRdNp8AJGWb
1WKqm3behqIX2CChI0k4+gLi2GKc3D6nyq8Om+HrAos4ZjPlao1Rh0kauL6L8zr2
Fg0r+bGD4qBaXy1sVLj15cSSQZ/ZQ3mKBelj1VIiCKaVi2SmwPpegvcIuGc4G9qm
qtthZc/DiQRLsVHM05s/vKXgt2M5C3Sf7CU7P1UfkA89IQ97aVg827OkFYMEJjxn
3IgrgRSVEcP9mPu3LxSsDcrV/NK4A3IgG3t1J4MDs1BcmuE5cf7cy5mK4MIqkhxG
aKxhU2Is/rrYLgsa7d5WJUXrX17ZSrDU4vVtbHxotxSUnOx8VDCYF6/OO/i8+EmA
LCFCjV4B9GPaRCqBCNMGCBilzSqXwHSiBN/gRA4eEvysKq+D8HmbQnfFegkDQDzy
JzdA3UKKgs1VF1nuv4fF8Z34NLE3zeatLraN4TFP2wo58P4A54b+/2jYPxmWNb9b
ba1Etlibe3stQL3FJTG+HTu6i4onWShSs+O42zZulGv/+D/iUl/6plORwIHxrWSb
oHmPIjNpZgTFk5h5TGCevPYV1gIhR8SnRW83qtKkVsnq1V+GnOwEpxfBiAKOdEln
9wURlvyc6Gs0n+IRT+P69iarK/l5loupi40B1bq7WezPUgmUlKa5PVoWunkSsjC8
yffoy2OhI1e02SRRVUuacXnJS+UkLkiScErxi1Dvq3AcJUBgFIeZ6oXYv2XxpmP0
0SMGyCvn1Q6sELX7xtc/doRLsgibq7gk1uLQrnnsv1dKC9yxdllVnQ2u+tiMg1GO
n6nVFspjJprKA7b4HEFQP0vGCAWN9yKTAXizdVQWH6xEmXXkyHfuWQONmp/c6I71
JyVvqWkGy22HkCJ5f/jZhW3FubwqjrZtoCeByK2XnvHV6fM6J9R+BqROAt9+75uR
z7dxio53K7/I7n4CN9zddlMOu50cGKaQzrXA4Ivp8kBGgw2suyrD3Ldj8JeliY1L
NS3rYEsFcjc8/8yMul0VGUMM2Q0ZXJYvYcZxbefnxmBbh0nKk6R6TilwvstlBHVM
r9OnpQZENM6AKqGdawfSCeKSK49oYzF6Pj8dBuawx2LIdXeF/aUgz/0XMEwujOhd
n9FBwPosXZWYj7TdBH5l3hrMaTaszRvNM1esWZOWOLy5A+dU4uod3EUKtnE6gtDd
MuiZTxkuAW1ghlf4EDNDNcS9C2ZLLf2wkBfCogr5VkL2Sb6qD7j3KhFQeizTQiqB
AUVRgw4Z6/NeSTsQ8/1P3OnA/x2OW8IeCjU28QoP0EUuQPoTp3xYQK/QJj8afDZM
iCrhLBbgfJiRvbB4Pr4gE5pCD+cnDfg1k1EIzjE1XRgMOVItrRYRNSk/tOLC/aSQ
ro/MJplKQUlQYu55ygInzc4CFpgucte1lEOE2ZKZ3wCsAfH3ipJUvJLi31RlEjmv
KJfJn0ULLcCE+8TKXvy0NDNGGfB+X8LmrfU+ZFpwAPDf/mgEOl7i/KEwSIg+t2PI
R5J550AhJ7vChVFBPuUDBIzCvm3STn1tRivv9Ej4hV+CfD+XlkXtzDJGBwbnXliR
6xoeqr7A8YWg2OkwZ3jopEPso7UFBsAfX5r/YWYy5vlonuVwEUw1VAjkwCZGfSnp
xwjmdEtVbtZLTAaj1xiJWKa0os1WP/T3ezKgrcZZ9I4YawEDKvIympPwdz3BtI/E
dCsUGgEgiCzdGawoJpysp2uZE3wirc64JzHqm0RaCJi5x3GQK/nEhqcpNn1PAbOS
lmg55r694L4vs5Fbe81K3QxrDaiItFeiZ7DfyozFGwtXFDntaGbPAZm19U2Rd8m9
cL+ggOKnlw0ZSJvvudFxF+0gHSUJP1uaXvYUozZ22wHs9uamaitX4f18K8Zif9bu
IpZ0EvtzWfMtKw1jMzURnt/ZXk6OeNZRpHJoSP972j1PQmcy2SC2fGGi/PsgRZ8D
boKGtMfI2IEmwgqr4iJGEWP4Sc+M+8Ge8ldJ6yFKmxJ50hAAqy+IF0/prEEE6nLK
b0bm7l5oSTVUMWuXtE4BmhROEdBkbFeO67uGRrjexiLjQ5JBtyVw5J7Equ6Af17w
j5ivwYmNaxyRFDwBetZc1qmKCcrr5F0vlp/NwqTDQJQEVglZBV9czGWszrHDTuYY
sib+Mry2FGbl5ZY/t/l0y9ODU7r2rPTc4pO6xP3FVzpwQefck7fDiI3UT7WaeMU3
DumV1C4JYalN1TpwCTtrJzTBHJ48hWQ3f8fwtbJmsGaoTs3OaT1aP9ZIdaDUGBvy
P+x8EwmbW/aVF/D0ajSe3E4hObicSWjGdPGjmyfOl15sQnBu5r7YfwxHRy+KfQaZ
jOHYcsKwzOUnHRj5C0En7Tuxrew/h0ySY5KE/849voHlh/grHkPGA3nT26dc6cxg
7RHuE8gr6C9qXPtMhMb8LWpr4Nx1RyJE+F4MsK84nQm9mUUKXSh1cwrhnZHrABVF
bzSlBracXb0uOzPuoklOJmPoL0jw+Ze5GbOr9UwX+xglNo9OrU89uCQWBbSsSzhs
tiUORNy4I+1sJiWpN161COduF07HB23End7kUdnqhIL35xQGNcF6CPQBX7S0Ujqy
rRwdpfJqDCW1OxvHR87DZ8kcJAKYZn8ca2dNt0K1WVcSRKBky/LFpe7O1X/ISWmS
aovDTCa/AQo+SRvQbMqWnjWtvEfAjB9Qi3zWFOQb3NZarQHMohgglw+6OntkEOQ1
liK4NVSL4G3YkHKAnx56GGAJBwjN30CWGsOeJfyzMGRUOYh4LCif5nJX7sX0ma4V
zM0QHQkT+NWd5zWTA5Lpb5wxpjgNkpkemBXDfAWnHUMLOjxFVfJHa35L5QuYEnzs
mTVXAZKm7VVwRQk42qdIEBqXPRIVf2QkJYvPu/7VdNDGqliFURr/tqPA6T08L6HF
pfxmsssY5lcb+fVJA17C5mbmoXQu2eNmvAwP13hy/7DDdraHG26hgtTSfXSjEzA3
v/0Q4j7xfmJFTgoCsjD+m5MojaqWNb5N2nn7af5IGBD1dzvwtGQOhVZ5Rw+ORkmO
O+pWO6J60Jmadxn7P4O8MvkpC0gyK2uFpibf3XaH2T7pCRVrX94FcKtWippSXcE5
i9zx9kWuPpGI0mfg3wrDzKt0IVMptSXYWjTD++Ra1As9T/XZs2Fye/SoVzgbfDz2
PIP8ouKAqq7cIdc9fjCQ+Pyx0W0RhxtCFk3xi+39VDR6Ak50pRzcZLavJc3gHrSW
F+agJYvNHE7Px8yVGK9JOntTcyWCEbw7SzIFOf1GNK0AyxTqAuW59dQDja9s6gcw
3nbtF/Lw2OvVio3uL/gnU3PGJFAbbHY60Edq1/jOgfJReVPm69hx8gDlCMb3N9uH
pjEckTOZYHuC9fY4WPDPDXnBhUDmrIDShznaRfY/RSW1jNscicjOE1609nmgeSoE
fNMRWJs/Y+VNwu0KTDnKmoeEXFQNu4uNoMB+GJx/b77PfRWkupPymZrPBufuo0Fw
gzsHGbYtm60IPhX25fld03oU64QjEGkCMpH8je+M4bzaCjVRtGJiCMgXgoQaA6jx
SQ4dh6Y4Qj7QJ8gkz01kZiB4VzYhRkzCKYtPtl/IE/OmUYSDvhTnKCefi09KWUOY
NDJRLCV34JsZIPE4XsBZHaDXeRhO7b0gg7UvMTkj4FpKlxXs3sAapcf0l+di+WT7
E2od3ryi6DKsDv4SnxtKn6eDoUZP6BdVEJY86KIMf+zfLUWedIjigvmCBhsfPUJV
MJ2qV087OXP5vO6BthVPAzeUhgATQGXP2rXoUFLCEk+tzTZIlzTzhp/MTuoWMqbp
gTgoDaLtdmNSuov+xzuA4z4BPd9NbLtIYEb0nDqI4ZRNLDcazIAOhWKsA+gmi8Gi
d8RPZCn8GO1KODpHCgVg3jkCxUo7XyaMYQgj7CeaE4jIyryUswV3kPNnwNOW+Lsr
8D3yYkMwLcnk/Bj5TKjeciJlFfi8m+c+I+u39lNdioEtUecLaL1gf2kMMskxBEVw
E3vtBpxMbGJuw3S63oG/EjYTy1HocHd3b99EmEv7NcAeRudkkGsD8xz0inZ5YehZ
Xg+/2dz45T/c9NTE38XSGWC8pAjzUSQ+tx06EfaK3a+T0urKgsUFRjhr6HYm4kkV
ck4RIaN7aROvegWk895kfz++vlNVOVVxfd04BGIGqWXynA1iJYQdJBOEVCA6LgP+
mzMotAe2SvHxjfAzHKm+K/4yBDy8F7bjwmCu3YI6r20Iyebr2SD4JpDLurltg3CP
QfgER5A+BPRlNXYuYrJIj9rOJb4SP58mk6ooeGccsunVNHYitPncdDP5SJPNM5m4
6hudZoR5hDgQSAw272EubCGWT1HFTVdVs1pCMecva1YZuufZLRqI//uQFK8zI+l2
jpAJoCaais0Ki2ocJ8sYmpL3djZ9dxb0E2L8PM/Qi8ngaIUSO2Ce/4E7cPLl4pW8
72QQK5EeJc9Dk2o1DBZjTGE8myFfgAUuB3WiD2r8yuG2Bei9/mEY+KMVKTBQoZ/i
PT0aOXFbUOd/tOsZ21KtuxkxAsCNMLoi9mosT7QTdSRG54O9jMs33gE49HFpq3g4
JjVKi6uOXt4JxgBDgWnH/Y7mz8LqbutN7gsQwT4Lq1pjIcoCIeN0vjr2h8AjS2Zo
jF8a7rRM6pob2qFenZPt8HoGvfPxpxvXOdazQmMyMYne93zzJOGGeEqYmPHRwk5d
qDfU1QJMAujR+JiynCepiuwTqIPn9jkAkKFAtDDUx/C2yk3ChB6BgsEARbszTksH
AWXhonLL78JEBBOm6MEjUHTCHLMkV2lmljxVue32DON2s+K1X/y5PTKQhm/pfIAe
N2pcl4ijm7+8ul7H2Pks4sGFtPjS8z3LOJWtzPuUGpGfscWAFbJOscnnnDnO5hAf
LnaNgSJ9ZeZvHxP9G+JnPFNwOJ9TDs45FRakQl3EdLexfTM48DEGIxXMh1iD+wfM
6SZ8MmhhqI8KHPB0kMPP9EuEz+0kH4iGPfKpS1j0bePCwBtc6Xho62+TZtf/uGAU
3ygS+UL/50CrqvFsSP9lV91yuf24bAp/2MDU23tqlLV2XWSGnz/qKmXUzzuxi0zY
f+wtxQek1UkHI62cwwIO+kJvt2kjiCM9NeRjg3lz4FsLKpJHj9lzB6xM4Zdb5HvD
tMLgU8x3iptHUrwilWsZVpdRR5luEwSssaOGt3N1R7o8WZhJPSeKUBv6xl+e2TpF
KHtcjJTXjlPPzLwn9CW/heiHlyoAkC7jnZ9aHenIyIhgSqkHskv1+8mOY/9kV83/
eE8k5YowoAtwEwXaRNpX0fTVXFhraWlPxD/DXEzrqbkHogVv3+/baReHWGtocKWH
+quRb84PwXn4mHTqBwadRnfPBqr/Auhb55VaoS/ofktH1rnCYieKJGdNHSV7kMep
QJW3pRTPKvaQJoITlo2PtdKp//Ewx8ceG+g+RASHqmCLJNi/h1mYogXBniUayC/s
5TjbMLXoP8/nlgr038hWnQrY6VNfijVSQKVwwGoPgfLCzXMcPS8HnPKdNNMbB4i+
ccCbsxnCjA5ROH9Q3aJmmpirysIQ/agpN/9AL9cNSFOS83HgjPUKFMK6XmGnMXCE
r2AJFSVbm8X2MS3xtjIIRMqdPGsiF7VRxlIJjLH8d5QIN/norDOPN3Kc5UNf4gko
r/5pJ7e8/oTFr+WVYd93zBgyBepgJY0NB9HZpr74E8z1ZuSstyH4hA5OOdWme0eE
dEMjdROGbOyZ7229MMRT68gnmyC6Z0Ehew85ItUJtXYlpmTZmd1C1fiHke0HqoJz
3cARTmB+slpyHb2sTfq2L/+dEZIouP5EnlzPJpKg71m05TN3JlpcSuO+hE2RFYTu
2OZre7QbovkY1AIq5vFO+PfYXMtkxi7Vk/EJvk7i77OR/2Y+KXSV5ulyPI6FpTpe
J7kvxOaZfzNrVn8E+c67KB8ZMlHqyR30F9f/Tp6J9LKQgqa86VxlkG3k0rj9bkHP
GdOBWtggRtP3LjTPkEhcMURsUEtk6nKByVMsmKqz1mO4geZbe+COt6t+6XU/N/jU
f0Ap6glCAkF6LwbuzILRXfbr785F3dAn/PjDrNNVUjIn/R/OQQ3hxx7ITt5XHEss
Xz2LTrzzFpLSphdpykWG2HsYxXQgRAU0KvLIIbb+YRT8V8zaThXvH63W0h48L9Yu
zECbFJ1rVDGP1CGO6HFYKc/8kVUfpehG/K2yL/orSYSVw6NzetL/G6ZKtAg3l0Pb
XrvUx53EP8veH6GfT3AJBqIXxzYWxI9A1ls//jWkxB6eJKtjIpkPlHLwjX2Ckquo
VaGr2U5iEYujX9qIOXknns4iLsUoeWn0w61KhXMUFNr+OGVlW3fyl/8W8Ar3B4+m
arvMe1FJEKx/A08Gm71ntQ70k9nARW5Kzm2mwxxSBdTq1NVdZHJCN87evhC3IN+N
tjmZHlsVK1E/FstvCP2v3tvZAVwzt0+x1XI31gkxWk+6pxkULLzsPu8UVy5LjAfT
L4Edd5Qgq7FKl8SkIAz7H9UqxSQq5/ExyVT7ubeLx4UxZMr15ArCjBEzkQ9nPq0f
+HpVAFGU/kNF1bbLiA9xsDn4ghn38GrzcGAFDyO/XofresmHBu4bzIEOOjDlk2EE
/tcWA/iU0WaF7wrwuBvbvL3ORPe8jq6yrntjXFFNexjtVDwcXhAWSKOVl7PfvYbZ
AoRA2oJ1WD82/wM+5Pg0M1i20XCg3r1JziwOCgjFuyKoxdoUH34GqyVpfT1cAYbo
XVcZpXVkGtZqbjVEKV/Eu84Pi6YYHRbn0cJqEopkRhbLx09p1ln+WnAULWF2rspC
MMoV6jHyfoOztLeE8kxNMFdedJzIX29JfRR9tu4DIs3hilT/OaYSOHHyWkbfZiN8
m418J87d+tmljy6WiWP/+pqYQNvkHvdyXXbzYAYWIPkN48pXK5p++4BSMlUdtWqV
vp179cpR7rbvmqFbDtWNeE++Wj9VbGR0+CrTv2guDJViT8/Vyc7OfWQuoM2W1f3Y
ePGjzIhORhjRtzZzo5VMGE1hRQlEifbL2gVU+lTb2j1n+1xEu07PLrFgsTzAWW0W
xnLFJ9zBq7HBkTUOiGbOrXLos2oOcT22om9mcMU/YLwH9uThgS8eX1DAYu6eMUjR
he9q5pznT2JaQcCZlkQKdWk0dYDqqJeyD7xCQiXxixmJR2pNMUTdeT34NhEBbwjW
wZbWZ+lWBzu571airOjGIMBqGDHNFhTUqZuRY5cAFBHY4rfw1epHLd8LHPi3x3L7
5jjt3OUsnrX1KPYjXPPSoraIzeKButspEHMa5hVImWvp71mfhYkKVH+3DXkERLVR
gk6UvciKxwkz56MFyLB+aGjg6abVIExZ1qehwjr5OhNpSmP+wY8syWE0KBNxEicq
PA1TP/lid9nBuSvydSoily+TobmkBGchE2MfQA3eDr7avsrTd8SBiyUcaCy2a+gV
UWOX/dyHKuUL2yvCpNrGhvLlv8JGkL6Aqx8HtVDMDeIPnhSZHJWB6xRapdDhZPUw
vQexkgTNEkZW878JFEzcHGTGMM/YlSIOO5gtfYsEBmWQ9NxLNDOABi3/+pfzwqUw
KemRmKhXLbr1j+VTT7UvXlM1CYy4IGmPTy29pnhumB5kXC4EH25jHIgF1thWGrMC
zdwwBcLD0XUZUlHTp/q68Yz/hMnMJP6kc+8eom6W6Zr3HUlH37Cc1zliqKuwLlEh
Y+cSY0rF/hvpURZiR4Yzr84DU7SBzU315UdvIGr5qFF2TLNHHbnctiLTuIeOvg8f
ikqnpX/dHliDboTNJpx6xY0JbqfxyDXVeCRVwb1D8EuSrYYIGv6ixJ1RMd3vHwsa
EmgtNFxhKNiYCnWlceYWsaQLo/pBaE34fXmrbFU8yDc7Pmi7eM3ZaFV53Vd9qohu
WKoG2n0oRdu6bHJQ9E4T50jTlSubWLT1wBwr2jN61tTQn2DcA9Vhu/9ioR/yvtrr
CxMas9RoBEq3MnM1LMoat/I5vxziDYfaBe2Oy7JgzbrQl1haWb1AaYFJ7kX/QO2f
NaAD82g/7ROtrKjsq8kvfbXejssbui5wXCQ2C6VEuJAKNu1LDs80JzTilxJffcUg
ipfxf3KdCaq9KdYcK6JRnTkgMU7q3Q/rOQ/w75lFwP0NNnVWjm2j/Yx859VrUjMK
k7lYZOjSnXgy4DPRDOBxJo8S4t+Fd1ajSknLFSnI79mluzqecDy3ELsyrowQRE49
uXlNAjUuld8+HAV1tYgimcBDocWGi7oqTXZvQ0gMj3b7Tct0ddKAd0UuYn8S2GUy
PWqIa5WoQfOuik3E7fIhcLpr6fzciZvtDJi+OUciaegu+2BrVYuGvLu0bfCIB55j
ivs4hER4igBsD79X3C+GeY4FzcNAci2ahzB6HvchniMqwbRMJhn7sBcpfwHZ5okx
mn2B4DYJhAwCrrAC9GJFOBG/593LdULdiQ/5kagJDWr5NezNkGHFoPWFNlpz9nT0
LdagOpvx29sR3ZD3i/cXFyUglWewCAap1YWoCkVTkjRpOzeifUUC6fadd/7qGD7y
TSli0Yar7h8rVtOz5CFGh23jCZIROAmKzpkQWGldjnru08++7Wc3JBV/TgUosRDC
jyCUXgbBULkmul6Lc/JnDhW8LFERpyy3Gjjdx+2bK91ImKccV/ZoKBajpqFytqr1
I2J8lrSlEZSYdelhhcE1Vc4JK2+vHYdk+67qSRNVcaaLM8N6AqWNOOirzwgeWK3o
DILgiENVsgiqcMXdqa9v7jp+e8dKCHQ4qjYM8++dMJCssdnlNERFKzKR+yWiEyee
Kh3A8KY47KA1qQu/UcV3TvCi+84IsYds/lc4Az4DKB5joefYAOu9S9QfGme2cv35
C6gIAuVqrNBbQRNyN/Ry04FUu4XiMsBvcku9fTyU6aRfteel85efBb1oqMwdPwj4
CnfmqELSLP7xsF+9bgHmAueo8Bcc9CmYlWwpB0g51nmeyvPD5wGZb3R9GGxcneiO
RghivGAtJJHAyM0qjtx13j0YWWDKzF4M/XCzJZFq9rDa5oDzP3M2YNB5+71JS/OZ
6LiQgjV5PWRjPBh0hM7JN9xaynVFcOEG22KgapcJdfTKYejN+RRtnKjIONggAdKy
ytKkA/bf1F3WSRHzoiVl0QnPQCo0/1B95I+fyV06kIf7Nwl/pr7TkcUErWfVu1yh
mMD2HzSWvopQiXQDQDKcc2Oyq84raqjqxibw2W5mYCBUfkE01RNQNOR5YW896vt7
1NHXBTsdwKZCM8flMWEezYSpWnl/obuH6ZyChWJ+soeswZBO+ICt++hH3qIu6AAO
7laux7Sy3yKY4xGMeyWZPb6oaY6+wZZz7arsccOXixAPwPf3Wi74uqKFsleqDrOv
AIKMoclhe9uem0eA3vFdTu8I82wcwV5cBifwnEJu1zFDUagJwwiUb18EI+/3o58X
jg97vIxuPIbul/wrHK9dqjgo5I3VgPHWJRhpQOlmLWat2xDCMLIgKvcHQV8TKih9
c54s4lzQMA1ONQe6+OCBjTTKdeg+hWp3L6a3TkS9TWJu536UIzvRQzBGNaEwrolk
Emgul9aCLU8Jt5N0Um6O8rDx/fa2E21HDiAV+9Hqa/oeR5VZrjWcpR+oNqC1Pc0i
rlx9nA01O+afSmQ09eMV7+NJE5kDowMidn0OWl2x7zRYbCWnu8djeAbIpbr4hJKm
3p2wq5fywxjj2rs402mfN2utahWwRwZL/DUQakkWuuvTJVe8k7rdnXvrFXacFaI7
q61NaNU0KXA+4VxKoALreCDsNMd+Pjs4hn0rWlLTKce2M6d8pbGJBmiFMf5MqZgc
P9qlIG9LA4GgmGsz2/77qBjM47gV7pMdZyDlXIQDnbIlt2r4nogXQ14zfPkztS7L
/jwSmFMWUH84UaZ1ZbEFfRfi8k6r3em1zPJz616SXeJ/wZidIeRnGGwl1dbJ3jqj
8xfVhRfyK1BRl09X74iWwKP+DEdxowRXM8x0/Tugphfi7yPqOsMNiWKYTv1d3Uf5
dqwoDedaE7C8C8ytmaYCO3ryqsCM0nqlSeTszA4J0sscfx6UUcDeSJbxglFwQJoJ
IywyJbDTfrGI2LPYkRohxncqy+KcG7cvCeOxRf8knDj5YxWNJOu2S8aWU0F6fUJV
w0IMZ+U22Qo5Kn0I6k1o/sxBBm9LnSUny4x8JT331mjtc7udhSnBrl3D+wW6kgO6
W7LhTEdgAmoixuZiAYl8SSeex6ykGZNGLOhsS6r7CqlEwLFnycGxzk+LLrrHrTAU
mSuNNxl2wT5U4IlS/7B/ynfP6pWrj22DFSGxe5YBonJRiPD9KcLfIsUynyVJw22/
/gPOS7H8EUa728FqLjLyLUtsCcEnySyLOYGbh4Oe4CKQ6Ym588b+mUvQkaSk41tB
AJJ6jieUXfGFVmdSPRtwRL9JOb+FHvAx8mMnAqnbVZKwNZr9c0/tPjvn1yUyV0E7
7FIyMS44nlBYjqKEQTUUnedSgdXVpOMQPsai7bsKsTWWhRZpMYl/iB+EPpUdvebE
tKLw1etHtkhpk136kR1XwadQliRmGQX/sZgK/8fCmfhQABHboi4/WltPeVLFXxvp
Y49/LSya1J8+65NNaSDatDu4ai45t0voAszNRwj294q0pQH6icbSsfSOOvjZxInI
MuDg6XhtSaVxXvMiLMVOfRZEb/ca1ipVAW4ykon+ILT65SQYrNePaLjfMrCVxyY2
X0Wd8czKtNxbPBvqb5LTcNY6rzqTL/yn5Bw1r3NDG6QJ/uDCh7DRLHqOzJGs5RUZ
i07uDj0pBFmxGz+Xs9/EImS3wXs6wQnjnoFF6llzNt+TOG13cnHXZTTCJCBJ9bAq
YGUS2xrVyajP/XX/kaY6bHR3Buag2sHishQeEy261vtvBJSKJx62S0ea+8pS2Dui
pmo0DxpCSJG0aFovgAFMDef4YZC1WOuuDVw3+9u4HLquDB/Ab1uaztZAP2iS4mFo
+G6D1kXTNxMNplKg5d9zPgQ86kFQKipJeKvtHqu9Csm7cqulTLluE/B/OIJXvkVA
m/za+POk6+5xSwnEe7thjkst3mDHamyf6EccJxNXS6buF9mPqN9w/d3EKXzAI6Xv
y2kD2KTpeWPpM/lLoMd/1FKe2IWqM4cZn6XcMBpxt89wneZNleW6baamPltWxU3F
InA16ckPbM90zhF1YwAxMAMvXLm5LKt/FKdKHCRgD6tbHu6cPKWk35ui19ZYtmGr
sC6hL3wJSfZqX3zCmUY2nE93OFsk2krgVF56r8VMQGzbKniuJR9VWTMkiCiCDF1S
VyeicXzykfRIbuHC447uerVr7W8BPfL08Zr3JtHK6T9oY3LTXrEfRKO+IgWTOP3c
F7uLLF4tBTq5+cghJqpZ3fJHnlEdAWYw9Y9ZuVtHb765RQLGLNPzzcaQsvDfn6sP
W/uol8oH3CkFod2qU2tcOH4UDYfvOgN5cq7ALFv/oBvZDQNK9wT9BbDUuSgQXgNi
e9Sk2hM4F7f5TXLlkCz5PmnjaqrtqBioNSP/C1KtSKs931iQz6YNsJQNXnH49OnN
Nn574OAdTtiRM7+rKRVug6tv1qPQ+XcyRnzGE+CuawMMl0Mp6/lon0/CIdGVFS9V
3/muyLfYjSE/AjO/5sxxpM5A5cD5tVAqyKhYny5JBe3r6LWHqQIanVJlys2l5vha
Jx1fTkI0NW3/YydsbEfZcKKlrezS+nzFIfk2JsBWh4iEDsPa3bZHltNk7voDu2gd
0wHDqhEqZCRy5/qze2yDTvabC73mdfbnhgXK6ksWkE2AAE0CCerSk9aWzGrozKYn
CsXn8iO3F/KdvC+Yfr1lry7t2oSiq7oOK+5v5m+OCGTBf+perhlcgf0aCw6G3akK
8U1b13Wdx3by7Z6MhoVdnw6aGidl8ehY9Tp4NYzOeYKpNJ1I60O3cThRiw4fF36o
xipEAyM2Y8WFUd0lnggVvaiPoukMopSk5YpgCBAdA6EIeeXcdFH2QeQ47NEF2vdW
I4OIAuiWY4UlNkwjopm3afMbTGEt9RC8JxYrc2zwlw3e+EB1TrVE3ByY0f2BZqog
9ubjNj87syD7lL+bmNzGCZB3PKMk1dthWXWOMyFU2ronWdt8cY/rqFDep233JuTQ
ekGjsZHEXkrx0OnGHUHnzgRerLCXukqafVfnr221+cHHDtKKH0h4VkTtjw1p7icz
vWxShKcgpp28PYuNIt64iWew0TkuuuEzuAZHeww3QScEvaUUACVSD00OWsjSYpfh
jag+Mfq5/akNBkySAOBAM2F+AT262Uc6H43A/PoVPwPmxS+7DDcahpzZU9jmXfbI
SJyj08y4K0JPjFniO77zH6HR7pMICJT1XRZkKSYz7KFuk7LlW5cv6Ks2jWmB6SVZ
WFd+Ftv9FFu+L7OKjnQceU+kYwmB5SuSRaiWmYMic9u4u5REiCx7HKO//x0m2YAG
ujPgHHemrJALKJV1Rd2EFO3iWfzeRoP0ZGLr7w53xaL8KUvjy6rTFoHjZhR0XoPd
OXIt2491bf7LgyibVSL/ZH5+HcOyV8Wu+O6uH5NBekOmsM74JXBJldIBR/GYCIUB
mXsX1SkvRohYeEtt/XFRJU7Q5O9Tx5zqFMoPBqYXR8AUW/P4B61SvPb1sploRtah
zGX5f0cV6XyMnjPAgatcXlmskN68Gmvc0/dgHclSMyoej5i/k6FxbLZcYSeS5WX7
8vMfAzKc0gs0Um4hkSoJdxdb+qJetM9zHW0SqjEvS7VFlADmP59DIvy+uLliyaKc
dyOWpUqX2UN8EW7/XB8oGyPQBnV2a0XgdrRDWns4U83TZrh9yeONTKXCkZWnnkbd
TWVoVRc6x1Be7SQcJh/O9+3pN9fY6jYajEpLqBW4qpjSffcMamD/seoal0mvO4ie
sYV9mA9XtlpFL5YhpJe9zMXB8XI5OJGyMdC/4QKqUtS1M1hIRrB69dq3toBZdBld
XkHr5pVdqQ/USEMqj1o8czTw2huasBWPd6RatUqpdKfkGleok5LBxnPrxNb84UCQ
RmGRHl7XecgiMP4+saaTRwVXBU9smZMCHyMrNR0xbOCNGGiMckbatUTdgxa6+p4+
IStP4ibi3zMDLSZqL7f0WqAar7Cq9mZhD7rDevmTqSXRa+CXMqHB4gYCEQq38u4j
ZisoVqWt2/R7UZqq/qoK9StmNCTT0oRZEmlop2TA6HcGMzTbZQRvvyPu+RaJUun+
NJCqqQ2o0L9wYcbMLvMR5MQS3VIWSRqY40QBnTP7QJTpXDhgdxe162xGEQP+0TrS
LD5JTb48PyF7WBNuI2wa3db0m491e4A+BMhFiScBI23cbs0pgYQJX8GFdg0PAkEP
pEl+2pF4fuxfyZXI8M5lN/ZTA8J6CzvysH4h/rufrhp3UyKwvpEn0NkPNzKg7STk
VX9dkzBHvJJggW3IFoMPbRDJRhTEYNbGXjkB0+91OmfEK5REiM5tbB9ufUabZypN
JFxTK7QBybBVbdmzXoUQjVQuu9GzSQo+jFfrYRrLsGIkUZf0mUG/gtz/piHOwASf
mxtb6Po280gwPDqkGgcgeWCLPkjHQNOf8pROyd+hQPqvALV5XUtvie0RoiKwQXqy
zo1Avuz/BR7e0YvX/oRsIqmnLcsDk0nN1s7sWYHi1vSTl6hhsCJ5CKK5rcH8Roxk
+YPJYpBJGZ4um0fk1cTi2X8OtzVoi/3bhzLBfCFyeZd3ALDSIysltOBkE6xAk+OO
+q4u38mEipJWV3OCo0ElikrzLqGa/hcAer0HNQlH/MAEsg/KAoj2R/s/kj0Nlk6G
Eoqaq9eFFdv9ZGyffE6TpRD0SFt5EihYsn0S97T3JA4z5vAgBUwhta80K9RqdqTa
PLW8hfNA1nIpDVm7bFy9r7sgDzKNmWB9kjAKXwE3C0WmF466uQ+00s4Wu+vvl9rR
bkP6FnnTTEYEqa0+z9VwPotSTBB8amMjTARuwznUJpFSu0es618eYytuDFvlECTu
lAGio9fIkK9XeE5Fu28xRrN8KLb1ij68u4vZXP+7W5ZA3UBlh/tWvXPDfjhlIyfa
/8mk9R0BgAv6ajabOgT83UYitBUVs7Mk+XOWRUTNNu2h0HelRyfrw3s6PQK3Jjkh
/uhguPm5FRVss/J6vsCbgNkbd5k6mBEV/ZyLwvyyxbdstJgVuKyH3J9awkJ2o8LE
Iv0ajArZKB+Kc7hjewRvFv0WFYp4r6qBioiHZKm4VXxqL7ThZmFuOtPZ5BaXLNfy
Qr+89hQwW1JLDWdc+7AASWvkYHM4qaegd5UpVEeytSE8sqPIn3yi9t6JGzPGRRDK
MqfTM39b6r34hwEvsZiKiAoKVBOssSH6KDmjFC+4oJm1tcZmwZnisK3mzFIQyH/9
XX5OrVx/VMdJklkcrHbeN7IHUUuS+IqH0+hJJ4ea2pTex3LEpnPwlL77rdZmWGOR
5uCLn01LI26cxhlfRdN0jGvu5wI2S+glS/34TnIWbCycrsag42qsWnkQlcyfy2+s
sDVtepxnxRpi5R8CEDGlA3Sc9RnVMgrF8dxyLAY408vnDfH3k3GmNWW/vTQm8wsf
j11X0+4KWxTqIbH1ac6ut4wX9qYxzLVHyPuY625BlKeGCWBO1hUMyrXEg6hSu6b9
L5jYLdYwvTS3jeOqfveyTCiGTXF6v6d/P8rNkln3msuTeheqA9UEw2TdNsuun3h+
o/1ybN4I2KaGAg2hk/3SA+/2vcdRl7HZ03wEq2X2UaTwLaMCfO/GAdW3D28nfTPk
8PAaebBOBuMFU2PrLd0eVarNAQLb8kf7u+scTriKX4pxLz5U2g4220q13nDO1Q7V
BPskGyydHOph7tPZ8A+mXSjEIxT+U9jicP9oL6n5SaPOwT7K8cmNJQsG/SUFjkvb
odugClliHXYsTjY03joZ4K29oDlPoSIUCPn14sgl3JY1lSe17PdeqtMY9VdZA/FD
IdtTlzw42Btz2+6HO+zTdgPmAOLKJq2ZC3/1DBpV4nI2dVQgtKVqaEf1w/hPFm5l
XtqSEp6YecBX7jNFUqVoScDnK6xvt0OXMsYhqudq1qA2T37nvxgF3cTOgSJexYQZ
SHKJKHv7Wxn/ilu5T39+hK+Fcx6j9XqgvHsXTkneed5zrjFlAE+aZHcKy+HM7K+X
l9oJuseCI95DXEd8prkl5WdMrWvx0xYgB+reFn9s2F2fBIARfmyoK3f34trsuy3b
qRlgQJNS3S4/EBEK0MCTW62LtjZ1cVgjNVt0X56mLOosdmIPHL4H0xaF0+14F7+D
5GFJLK8FgM/r01BGzpcKUgRMr6IGc8Y5Tr1yAjMHvdF9pKhbhWLsfpKYSAwDitGm
yS1SD206jVmQMeHIVs8bBs3iZQi53nVqS2DrAIIP3vA3rmlmOXwlT5IxUFvmyb0a
SMltOPkMa6obK7Lsk0jLaDH/in3JPeuqt0pbZRxt8PXsFGind2OVmQ+pNqukkfn3
dyYJShiiksyWzQ30z5IiVGKeCF7q/dSUmq7KM7lReJPi4BMjntKvC/1OK9lRLZNG
z4hFp8RM80Fbc8EVMvmkNMFImpcfZFZw3qz2K3gaLv1151VxZSBbtllZEVoa4qQJ
uk4l+HDJXr7wdhBoE85gfje7gzpkdMewrNdbhtp+eGCf80IAh2KhSCSX7X2C1ARc
SUW5ZZOHE2nx0eEFePssUabxZXa2JbZcbMklKJCqFMsVDKbyldOsctex8mrQbs/j
ro/sqOV/BaC80Pm5ZfcoTP8Xr5l45/mRfu0UvwT4WNmUiGbmkZlL6JiJOiQLCG6Q
8pVvYZUlcVfqQB4f6dxfqkNJEFOzCELCNBMc1+oV2eVNYrSNcDBUh2OmkLekULBC
Q/e3S7RbPKh69EAfKB4fe1HpTPe2ZuW+D+0NyGQFp0YZnzwMgjvPkvkYqTUz841D
mx3gWJAYhG83l8IisYMsPHOrIBwsIrM9C1X0dEziwdbolI2bZ68pBUYXtfJoShJT
3/uYcVe+n/8a2Ns1CiK6F/VYCe3pTqLwSrkBp1AV9r8gB6ZhdQL8mYUD4rhcytzl
KG3aRc2MnKKT0RQPMEGNJP4/oA8c4I0IwCJg8ygqyjV3NpvxVBWhFOLELQUFdmqG
i1cRzQKchFJzwdR1avdwUhNWKM804N8HtvJKYjHQ0OOOeZ0TsXuSPLURHI9i2bO8
OAkoqD68/BtlkjQQifn/sbIiUsmhjEb1+gd0UWmlk4uhdhS0hBNfSfKzTKzs+g2h
RuK6vs3plFePBSFeM86i0LRBnZ/7j6QS8Wpw9Iu29l7b4FQnmqS5XZqFWpItP9qb
Y5v3qRI5SJlJ83C9XREOcis5v+urwdfXLilJMNR2V1HgMmjGinLZNGw6d40oneqn
GtP1HCBepE5MtWZjRtNrO/1YZiYR/D2irx5yUrYiivwznr4kkXHZ6dDugZV6WHKt
pFURm1ZIuFRpRSicNkr9T573wZtlzXUmKDoblxvLRKpswkC78She2GSqZD+m8Bqj
pSKkPN/708SHQvwZx7srdWj2/G5wD9Rv4jPMVXvb9QuyhOzIcmTaxdNiHdb42S91
mH7gbmfCBbEp0Y5dS+dGFwrZr3E6CxQZJKzWKKhIPG+h8CKQgU5lti2agLCjZBUB
n5P5EpfUxy77d7UGyuG39hnlELBkQMI+/wUSeVbxTgkKOJQBN+1HX6CqUx42gUkg
gVzkBd2LfguaAD+6aaEIh6hEbLLQQuvWjg4Mi5mMLi5GjZiMZx4m2eqM7bbwVuc8
zQNItdmEP1jKwglNfnlu+7I5C/ylyXymFXsKQ7/71PvouYPrlvdD89oNZcaW28Ye
AclmNJPNzByBEOdSKPuVM6tJBN7NkX8HzEr6j9n3HQF0wgsKmoq+hoZypDVnL1A6
UrEAJCO0F8RwZevUIlTF8GlXxAlsrBprKpID4sQJWgjL608AQV3SntrWMnNhyv65
5STBWFDHO34aZ1oEaWsGFC2PRL4CUxvcdFAekLPOTeiz7zJBuIeLXlwA746hk8eO
mgAkSNFLtUyxukBe+JoVEIk5CGNXpM0/ZlDhkyIUYjxSRs9yoEcW0OLToPNZ6Pi/
nzB6eLxfV+bEqJfO7B66Iq44AsEWcQHyhcaIietb9whKdvB8yz69MgjliglAApxV
jhOE6QYTuiQ/v7K48sEUwFxGD5QSpPtrY3mxZscb5g4tSsquxapDyN5clU6nsaMC
bIOopJfG57roFI8QIV+Du56M+iHwYd0o3KcVYOYbV+JHZxDIavzxzkQc1iGznlpW
jMTGlRM0qxIbnlEjBpi7RJS6FddKe1Q7FPh6lzY28BY4TBMc6sBO94hAHIhR8GtR
Rp5KbeOIJvO18d8juNbB6A6mgvFlCtlRcPMKKV7xblCqL37LZAfMQiCja8O8Djpw
s/Kg+ZSRUmN4ZjQzrlofXi1FZwyU79n4F7f11MmUsqmmgXPvnqRNU1mpNCdO6qFh
cFyj/+sSUxBeZMqeACSJT0rda32DyQCVg4T/e8RtSFjvVLt6/Kl7TH0gdM5c4deA
c18Ud9J8PPjcjBEW/1YhC+EAWnZKkP/my0mE3EzFwUNT+aB+q5b4zaVxT5qQhKgy
qzJ6NHd4yibvb+UVd1+1uqcavH8v58/SUzKJJPtsP/ueWFeM0hqTSXeRllwIawtq
E8fjsI2KTwIIpzvxWRnk+3FYn9qVTm2yCd3y7N77HBxfssahkeh6YR7GvyBoePSg
hGpca4yHowgESpd/bicQR6bk+NLcxHgiy+qTxIugp5sqE0Cm40xn+Xr9v1HF6JGd
I8+Qeqg/W3wwCm1/SuwfgWI0XyRNXFHufL7kx68HeiQSLoF1eGihjgKWZTaoqe1U
hAzfhr6ePiHoBqfuzCWT+o6JhGj7jTwQ4a/Cd81zJBfJ9Q/3YPIALS6aBNQjt+qH
Q2YKp9fzdCPBXbLXGPt+NyAsJthkIe8t9EYpjxdLSNn7Em8sc2Jo6hQD9aXa9qTE
Uw3W1Eett+j2KP8sICpPhspz7NZXrK8PNdAWsY3VN+3pRqeBpM2ZQgvbKs7Gyn2R
aQnUiNO9g6x/xhd3dAfXnRKKYA+IEc1PdDZjsGcDyNCKdf0Q9pNIUFsu+4Vteg9Q
vOMjiapzhDY+VP2bCwdNiKU8ERfcud1LwbqGmEFM4Skr2ikxlHglN69H+B9p/nAf
tEoXjdmqsgK9/o/ewHj8KUwLGs6p7uqNpwjtrfP2yRogNNe3hh3prZDzZZB5osxK
v3kf3bk54uQq3/Ph7+aqdRqwSosGbo3lWp6ethMkOu/9uj5fYdGkTzPjgse7F5Eb
4pNfSxSUZXBS4iw2yH9N6TkG7BbTqKFC9qHj6vujhZUPqaZMqwBy1Ngu80p6wQJu
DBQgbTWhcEwOm1XcEPpMxPhgcJuOdLOvOFpFIKc4EQo9zU7x8ISQ0nwSTAhR7Mmu
ARxdcf0E+/053ua9iBmUTApbplv5Wfg9PUT+5DDwoRfGoVcUxVEA0bDm6dHZDFVs
7HIS8jlhx1fJqI5r91S7y92XsW8LP2IdwH8O0E21fkQYcS8BHrOO2cd+hcEek/Kr
tEuivxLLYfbOJ5Lzfc8LKleLRMtxhcQJUEHw6/lep5Wq+gI0dz6USRi+fp0HrHF+
sBOHk0JRgA8MQ+gJXVbif4317eHMUG22K0PJf0RJavtpr9KnBSHuFxbVPTCYkgwF
gKyGDndFEA0n0KV5rj1b1LPjAOxtjRSM5oTJ4dxQ8v+QWGOL1OWRe4ZMbu9TIGDZ
bk9/9oai36ZLqw6kgK3SJVB+9FYxagprZL1EoEjqvxzEI3Q0nPEuvmK/g12wUBVW
G7VDh1FeCcQvxZYcfXBD5YafTbQJ+9aWhVf+Uj0RC5Ly4KuMxNFMdnfOnwqsQ8uE
xbM8Cv87+mcG3Vqf3tZkaKzYfQYTrHd2wIP+92w6CsAd/2L+JGGV3B7hLvk57TQZ
zIjoSfKj/ZWlbLzGt61qRSUh339gv4Xtla8PhdQWRogDvJOjb+c3fiKC5K/BE26C
lYI4gsR3seNxQhBMOJsOqQBAJqxl+p2RPNcz/vQnYUx+7KZujciJ/dRim0YCboN9
hyzXtTcXGEJVOSy9ANpcBuazOvweXX2CUhBpPANZLNUJRGd3TludmkwC6iGFwoO5
cYn/doU3dpaEkgu25AXWi19nxkzQS5EfhwpzbrBDFhxBNagqLY/hzoCga7WToqxj
V7VjCneujcKqICSD+RafwwgTkD0PO8nrmANdE6ezzm/SFN/prguX/pqmgKIlXLhQ
GEfdYWyyPg9+6J1jbFwcoOTukKr24CaabDna9hJuPZI4G/KNwcfJ45/tBFw03JFG
f9rcGPd5KripcirO44gIOeaCWlIHAfM7pc+ZZkM44BZROBIe47RvKX0SRjLB661R
HEhK+IUrffzZ/B2P79NFBPZasHkcade1feq4RqkV5FMCzCxDMI0luZDdI1HFYQmb
OrlZGpmJVj0WUaS93+o0R3mYidlTttmx7QTromuhjIwawvaDm6GXjiX/8DqhqEt6
ViKtdxoKqlVaXYC/SPsXvue42+MnBgvX6JUNPIHFtjG6LftX4Yo3DJ4dqKI/usci
hZsvP2Q5VmUQXq0q7i9HOovsJZOYYYx6fFIM/2NHqoCNRqASSf+AJTg2n3Onmbfe
DqcS89PbQJ5irlHck6Epae5vxZX3buhVQS1mLwg4WYQLEBwck16dKyxUVHDv1RqH
/i4gXTlkV9AmuLEVK+uREiPpOghxgkrWQn4HdFLwpXcme0BjDTcvA3LBRKQYgWvy
x4fK5toFYe5Qbwbtl0QguJDMVeOhm+PgLkUloF3Ih9jqvJ48fCM2B4PtxEDFFNF0
+4lRKhA8e9M4j+C92T2tmOKhMRN/9xJcMDb/WMCZkhg13waUBOw9lzhwT45JWVUz
sz5WjRKFMExXrmi5X6Zt4nzFJXKT6vO6bugWVMbcAyA23vfwpVfKO5gisKr5W6sF
W6SwUbnBXfVtbV8CC2GuIMoFhiNOo5e2KhfKj9k4K7xyScoc9mgAgXP/ix5VFVI2
oDnFCf2h7CSAfgxA5xKuFOb4Dmn/oUr1hoeIpQqC86Fi+9yqvZdmO8fBhtojWXN8
iGCIAP4o6THm6XLncMBmMmGeHqb1CefU/xKD8fY6C4iUmoJO5x6kUSIyw5fjnKzg
330/RY7WjMIbSN3svZR0iNemLWgDNYc+KSeuCd83myJWJdXuWgihzPLRrpiWxtVA
jeoCHgEC9xG2SkYpvxMhOORZOF5Blq3p/z6w+GxDoBO213S5Ors1apfwisTA2CeZ
vQPIhUmPTc7NPy3NmyJ3TnYxn4x61Lkww76+Zp312SNuJsEEHsFoVYW1QTY9bOyi
sfPC5xiK1zj9sC6RsrR0ZdLHHCGH2XKZ09MuwHKoLkaBSAvSuBcfqzNNB3M9z5lS
P00retqh+d/u04HvZonwEcx3azLNdGxWgIvrcQoAJe2gecYeETEEkxBe5j5U0F0j
CJ37QWlCtkQUnqpw4x0uy/T5YApTJjNaqwXfT9kDDRt/WddE1Zyq5fUO2GtqQOKX
VbejvneKCAa03nFTi++dGxq/7ihdS/FC34S9MmzG6CPKw45PqShJOnFUV54hpIiU
gA0kKEM9gprqeAA2v1ILa5lW8F2WUtqRpNySrT08CYXopIwuPdgsjH9kT56oxNd5
APLcQ0CVYDUzkolmAQ0R74p5PC2OIHk+I8VswCnpDd+JjzZszn3VQUpgzgnzYBG9
Csk1/h2/9ratnZzPrz7pEjBYJbEJcgPUKf0UHNP6E3dOk1L3Sj2a/Q9VfCzt9yyU
q75Qu+M3EI5+KGDAXFkw48MxXnXlWRr+ke0vaRSxc8cPoMvYOjiKQsf64SixjxK2
zJqX5CKtj9959di3Q8+4nnN/KrdmPypU2Iw8dkWU3JNkdHk3T6D9Lm81tdj5/Qxx
6+kx6eHGX5B30NVLMxxHKGqm3CidDTOlwDaBX19GKsEk3g2eXIPz6a9bQ0jhQaW3
iGfMKXJmzgyMhZAnA1BcPzHCvtm6G8EddpNV++7D3ZxFsz7rOrs5GkcRBDBp/4Qw
ZlAenTBEAzhp+ImzYPqxAo/pdHW7ZrMO/MJ81/fhSYmVvmDv9mtvrJdm6nWHYFv2
DL/r9qpReuka3TQ3fe5MpGiCTuL4cgEWx/D53k0Ct0JLD4+g0PnMbLCOclO08f5w
i/qEzXQaClGWRsq1zsBR4sjL+qj9k9DOTty3QGGpZUFMQ9KD0eVg8/gv/AU79mgS
17Vn4hYbf9R/2zwSHw5elS7bPzMwAmnwk8wmIdStS/OP0V6gjDrjcfH9RquGCb+m
IRSTD6m0aHmDAv1Y86O9CRBuMFbgsWHqabYcgXYRGUJwq9veiNsHx31kZUJOPav3
eEcVxclKf7s60cI3yUVodI7QBbA7UMQB87bjIbNtjbLcfBVfYt3TujptXwP+9rnh
k5/VYC9UnKFj8o/uSjnbnRY5+w17nxXH3P2LFtUwCukI7pRV7I/3DUAEG3oTqVH/
sGEc9hA8nyV3JVHPhmSKZudpHpK2CgthfdTwfNI/PTrmBqIYSz8OlDDsUOu590V/
mWDuDeTmC0EgAl+Ku/CHY5s5B1XKPVHa1NabaOWSXWnP1Ne7n4cBVPO/BmEYutFd
i4gFy4VYyOz2ikANgkCvArGp01gjmZAok4AHyWFuOPGploYiX0r12HiA01FO1Cdh
Zx7uKJVz6EpxWUFGNZBJxUmBJAKw/RiPXODBAKPfdMvRtCe5LtBD6s3I4IeBRijr
ZWy9tbn0k9gRwBTsSrVGcQD/9fR/v/kQNzzb7jSuTEFjlNbpaopC8iMf4lFr2M1n
aUkADv0W75Rm+I/l2fZjddKAWZN5+JnezTVxfG22ImZqNFK4R0t0JJX2L2Zm7Cdg
u4avrkg9izeULiKE9Evq6O6IxSfkPBQxNFLVz/LTH1OgSP3PKx1Zc2+5KTlb8/uk
Xj6QK5sWLKonDDg7Bds+mMYBYLW06OkRC7EC8j0xH8A7+/jOUvhkFTycrC8daTNg
6nbulY5Vx4MNhQ53bfLJW1ftuFgsUBYLYKYEsrtXXrSDqNfGb9w90cQSz38d+QDk
4InESbpk1pFOwWGP4ET1xyDN8yQ6VleQi3ctn83pwyvjv3Kq5RaW5FkEFc8okl1k
q/lgRpHI6c/nj8feo+JH+k6bUHEqzBweZSLBfaRxOpDu0JXzDmLcRoqZNfVlEg7f
huaQ255PlODKHxYmYIwLegobwBc3eyAD/AJaUQkknnMMupK1sadVeYnUM03wSfRU
lPpqpFbo1ojtYv/yx4LdgXN79CVWARu5VH/zNIpMs5Y3AB+9VTcrTf1gK21pDXo0
AJcSvoRgJFmCCraoA5PRr0MHEr2AQE1Ntu/awidiJBf3zyu+60YiPzDDDezl+FdT
2pC3hVoKXBP7RpTi1Aa28HqtNh0+QNNoK0v4jNFE7jrRTXWo+1hsdFmK4wlaVVwi
BE2QNsExyZ4Zx0fJAHGsc5DvOmRlZDsu6FYjh3U58953i27nlIJXX9RxLLeC6841
QmpfKfwCKauMRLFeUxplQglQW2dFeYrsH5ldT+8TojdjppVjzC4NaqruHVxFGpGK
ZvAraIVEQEp74q+njRy9FAaAQbUAVKNpchYIsJ+VZO+eLC4yo4oUZZIitk+FFhjg
MzuF9KRvBIsA8a+awGbfvab5khZA+972cjDFTGPyFbFK3iEm092Oc11++VFPRnLQ
k8vXAxgYVw7fIfiOf9RYUOea5jdx1y+E8Fxr6JfJLlhWBv+Lwr/fArz8gtCKLCR3
NaWBcfg3vKIIYeZcxmEa9ajfMJ8oE8G/AWs9DxXLOPzGbdfxH6Fpp4icCeFGeeXb
yDHkeWtIEw8pD9C+s4cXVqFORJ4nzOl/Xahzl5F0ZXTc3bAm3WtQbBuv+jvO7EeQ
uAdSTKWF8ezzUsgs07QRlA/cdOEQ3y6ck5WfIysW/t7GNxsuKSRYcAiwvZa6KreR
vBs4Rj00knWuhkbYeLihjdoQRj66mHSuk/fdgM7D7U1I7UWUYcrSAcWrVBKVPOgn
WyosCntpBXoesJe/QxSuT/xy5mxqx+9QprK2+3nYMSOoXitPRTddcwgYiKaykSBH
eJn7vtKZmr7VKlBsiQLRybB5k3MM79ATlLMsTW3N+R2HIYc1HtfPD/gcXBPykOPi
7goKkfaQBEMeQItnQhUlSo+6bq9hLQD1GWAn8l4mFYriu25l9zT7Bn1TWQ7KQt5j
IwXA8YHc00D8PGKQEruW5UlIBPwTe9Epa9FEG3DOyB6pudcHPSUVBmTcLnRtmCjN
dy7qetmJGd1kuMr8OzJh8sCREHVNEGisNBMlDFBTMxrho9/4k8tdURGHRxoySOj3
6qhprzznnB2kVIwCugtOVOut3neVDqIX5I4YE1dvs4ftKgbNQONvi7irB/3erBYB
9QiLrvBtUitcPz7c/d26Z4P/vZz1R5HmnAE6AcfKGJrvS7i56BSIgDEBzpX6ElgE
GcRm8lAUOwsc0ElYBWEgJNUMpRmXX8/Y53WPhakbJP2c0FhGqyl0YXY8G88yXH2A
NxRRw1hd/dP8kyk9LkRAjb74xlcNNlySMc9MS7/AAEA6dK4X1xejJww36mI4zi3T
xziwSKjtCzmOr5QNPpkeOrD2nljnmZGxZVvVzVvV4M35WmpmbrNIUG0xxRh5mby9
VSNncwbqHOIU7j1KS7jKOoPXFdHr1Fc0T2bbdjeuo/2e4y2llAbSy0AlHgCWlTpT
e+bbjHJbwNGDTS2f2RsZl4D7pZ7oPM1mUZ1zXMzVR5fop8gaBqSOePbVGajMx5ZF
iEdepuucOAXR3Ctcnxjo72iMmUVbFgRD4PiTC6OI6BrJ6inboN4H4K7PxIg6F3Gh
Bu2C0WFhdAPPMB0UQmq2Ny4XQY/Q5q8WIWhu41nEI4GgQsB2OYFCjvvJcC9uu17S
gCvBWoH/wsO8irTCFaj30W0M7bFPKeJOXAsfhcvwrvLYtUvIE6LfBaPTGXxJZmY3
+116mUfDx22nvUnpBccAM6nT5qFMkFDvshNKyT4O32EcKlL1566d94/m3rQFas0Q
mAdv2PvEM5HwrSXBAhw+qrqUCVlnVPz7B8WhYS6XI0O9piFWmvYAy82nbXrkxmID
aVq9il8vtVoTuTgpPuWSAnNYbk45ZMkAUCSbO9VnOKWqptbsGyvSwEOVf86cTI/Y
KZybZ13X1uRk8mzGLrx8bPLq6w8MceZ9orl87uc6FHi94W0sFDjvGY5bnSq+vd6h
siezhPdNnDzgiXD2UZvfj7djX3uZi5Fne4iMUhZhQsEvhX/lLIZJU1yflEUt7z5F
/algDU8o2A6A/Zm/w6h1LcCglWFF8sEpKlIjL82tIdBgeJ+XBn9bYTZVtuIV0f48
z5bqqW9PGhEKKOn77oAd88RhQ4S6zjayWmRs8IhrwnmM9bgb562h2/U/PcU9QIIc
hsvk2VhcJkhNoKYRwIccDlrRs0vSR+3DmpnOthriY27FqgW2MJEwb0Bim0O6Vj1H
RBSLINjqmGSJaHVq4ZQor3Bzgxs/7MZO3QpTFlpVBBR6FdPsvvBj4IycORLq7v4s
GsHfkeDNYwTb1/zfmH1+9DioJjlXwGmdf8pmxBLzUu0aARoO6UBoLlem2QzlhrLT
rcDLDmp4M4hnoFwkOLV9TelB5pPv9nIcIpfNDlOwtRDoLKN7A2Fd7c2GQX9mZJS7
yY6pRPlt2sfnr6P0OIhEdvUuwnRYLxANc1w1BSCCXmWlLdKgAUymc5OwRRHT22HP
8wAEYPyY6M6J3/apaZUOx7du9ejqw9IzIRskUyYGxoVcPuwKItmclKX9pgljd3y8
mpQjvI+VvcWZoYNtCivJsbqaAcWTVu6loHSFgQzghzyRhFz5e8AvBqAWuxE2em0N
8Y3RLmer65u9oJ5V/hrhNx3r9IPqeaUjtBut8w2kqIrRbGyafiEHlgAep9T/E3f6
J7Zjue98YBJg89k8SHtDVk4z+hfkIMrx8wmHmQMh5oJpWHTb75LdFq4Hp4ndP1uE
BzDV+7ST1KBBqtMnmB75XddeiKDAYFLkciGV+hy1IBsJw2bOlwYf6ueUXSZfBrt1
qqLk/FrHeoFklRWZzQu9sMUVV3kUzEqZ+iI9RLBJYnc0fLt3R60L04295Ic8swQV
l8TSCBYq2B6AFMax+P6zzVyz+fbGHkocu/EhFGo6aQ0bK1KoPW51/t87W+5r7aP0
yLtvrs2Ohaf3cTu2AvPL/MWK9rSnp/8IeFxtW37jqNYjWgkCEioTyhJX24ciLfr1
Cd1DWmhSZRcnRTYlsfUCF7sSLo4vBWHBnZLIr3Peid89+XzHwiU+jVSfK64J4vdK
R4+rwGw8SvXM6DtOUc4+wNEjZrs+BEozvHm6f1I1yK57FxXcdZqy1Nkd4tlbCbD2
Gff7eA8i9suEV4UaazriV3/FFM3uFdvt08QhR/bcYKiK0fcexDL49SNSA0sCmda+
koYAorSJduplmegzRMucHOCdEy6i/SQZWpkuuPjeIsD8jYdjpMTjYpMOGzKuDmLk
bZ2zbeEJkdLu2P0R3lQCJaXbsQEBU59/PoMds4LrYQIMT0ygrUmt72XCPwybnSWu
8sVjIVRu6U6DwxNjwyT1wLXC1rfy7iTP/8Ivpg66lunYqXEIuyuUEKzp9lQNdQO5
j7VId815dgrvKsKriDTH01BYuvOuaeq1pvUtLy0KSeHt4Qu+wDQ2syOZaXF0bQbX
UD++0qETSrNTHPNWbIbU7gNvRx2/PD3VX7G6xnAYtr7CzdumUAfQMk3F8wAPzqBs
GUas2YfdAoBofAmuSw5kf08pcZuz3CuM2XUncGdw+Kv7cYLyCPXOmGV5WHZD1Fyo
peskBi9Szn04mjPFh9kxrtzzcDwqzbrD7CwOvqYVMyFK2s/y6ynyt41vOkTQzX8k
mk740OiCLZ5GZloGCxR26nrHClaUuh2gmua2qau6AKneML64wnbsQ1kv/Hj+wijM
odr52RRizr9gMihlCdzlitZ1BfJedZofsXVwqoE2GdTZAvus4xsvMP3+WXvwuDEf
lIsKJvPIrGWKOOrAyTyMLNKD01rgGKF1yIAcWsVqKoJnjZwt4KhMqV6V9dFhHg8i
N2aVPLwxDpWoZ9tOPi5MtKHYfbZKpefsdCXTw7Yf4eIfLPP+GuBMYDnzMHQrFcsy
8atWrsQ+mRY2woJtVW/eQRHpLTa0aXQIEYsbMROijm5NZ8tgs4Pn0V0FbdG+S1PD
vIj9IaXNGA1QbXduLkTFyoVGAKzajU2c8D9Aq9GcThO9bRAuVbfGewly/tLj2EvJ
qDsJggVzbnjlOchDegAIw2l/uIc7m9cNN8gejU8Az40rUrgQ1BO/NnmGiDAbLHUq
F6v5OD9CmyQG43UZAOvNtc4CKrlH3vNB/Oc/UJwFBNYCV3ILyPM5qwDsT0zcKDB2
/cpVGOcumVjOGl6jcK4ipuQ3YeobOh3mkdwmAq0LJyW7LgRyVMjAQzB5ty3OHtrs
oNy//wlwMjZyeejqHxbCI3XnwESUKORUwUTByub+7pfWrkgU1JvlU6AnJkhHWNl1
CkZlAA9iw6T8g0I2xGtpNlJ16P9J8Y21Dg6JaoAXatemZH5hGmvNlBDrkecJeM33
/2W4EQdjaSHtGXR/aQyF9pbdJFliSgnJVcSCxrxcSeN6RGkUC2sAwy+xatUegtfw
0iZhu+AiDp8z7P6Fl9ACctumL0B4QDv/X3RNgeDnQQ4n83va/zPIAga6hbawoQR6
N4FQNvTgw5ar+aoWv1fyp3lJ4CGGOZE8LQDcV/dGdlDmf24Ods8jdFkdRhb8JVE0
mvAHtzH31mLhPp+DU+eijhtWWlZp2f5TdvB7yRWaKMWCRHyEc6bz9eQgC2oojGVD
19y82Oo/lRgvKRtVSyA+fJZukrpJ2Dr4MDvfWfHJd9urTIIFQ7dPSDcDvfINpXGm
LOxz8ZGftpFA/9GSpyGEmbNr40nnFiI3SXefapA7fV5GD8kOncFPClxw789rirJl
u7OGvBcZxtDrFLF/iyW+hC9Od+n7HOufVNN5PNAkLEyzlbNBDw9RCq+8Zxa1Qe7V
7RDBa+vo7E7d1VU9qm4BHkK9QcdVLfkn4zR83NQQ63AmH50uwgqQfaNGnNEF8AH7
UOLA5iDwEAvaH+xALoZD6sVyzl62geMFR3CgxYHV4Cp3oOxm254Y+QkliGbRyP/Z
rjFcHjry1Bp6PsmReLVVFDM0jKfg5dkHYNgiyIqAZSPh351IrTMBuSlDQj0iTwYM
hIWebD87yTCYktzDaLmNitIN/DASeW7lMKZObKddNW/umtMLMHBF4rg5PVDY04S/
JgmKO/6/O+Vg42aTF4ejWDaTvVIs30P7ygbGK9LVOQlwbQ1zebSF2qoRnPKPdOrY
LBKdU+qWvIyZ546aRdnsSz/yO7juw+zwRXU4PlRN+JQhBtILVREVAM4Iqfw8VQ1o
RNU+RjXR7fYVGFkCa1SsLUo7fCVkVKVD8Rd5qMZMZoiXTdpwu+3+sxyGYlTmSZ75
Yo5Ql0irR0uYDDJYs8i7sxyDGGI8gHalRES3nLuTPCnJeTDz+XgOUlmZCC/37/4U
USw4K333N6txjkeqbBY86YJzhBzkcII5I17dkd0Hgc+K2X3IQXrk3BwnsDCW2KC2
5J1GQGEPjxMPQGMj1xAIXpgG5MRzn3bBWzK7y/7hkfv1lpzhst1NE4EXHAV0p2r8
OtjUIkSV7e2SeNMX8UHl5X2qdrO7i+OKxa9jcZTn+2zJ/EKWFXxzQKiX5kF7sJ4q
XM9OzqkGs8sEE6Es8KJ1nGFHiRk+JJOvjFFlPkJ+JMkxOGWPASPI0OgtKtsOwvSH
v+L6Fy8r/zzx3/oM1sW+XP049tP/rRcO/NPXK6YvwASjrmtOhSe3kJ+TehZ+63Zu
wb1tKSoWZ8BwSFokRsfYGUq71VOH8/iGOuqqYjOAiZTKFh9SOSwChcT8UDiKcnGn
u5oO4Jku72Hk/01oO60BNfTjbSq3iiAGonZ01jzLBVF6eE6myZ0sKIXZoD3gvTKp
xQDRPN/jj0mQ3lWFVihuJYRxhctv3ls9Q+RVInRObx+Z2gFlQ/IDLDeiRnMVzg9A
QzHFlDI+QA1fXHvXTUYRNc+xgMqhqXt6u1Fi91IK6SIBkYGYPic9aJawhh02Dpvo
UeO+YSFPm4SqyKaU8rrXMlQck2nBk/Yx0YqwswcrBrbXGLZdypiHGWPye4fgyAOY
eBfqtPXAn/51Tmbuu5uiRpr0Uppy+zyNwpABcATmrT553B05u6wLNXAQY1xetcRn
6oZUoDp0Rm68Mok9BNroxMBHLZamtfpCDst9UOos8gdWVRxmmuoVKXUfqC2gCcYV
Z+rVjwJNWU0f5TWD87zk7CzWXitAUbt/ai9nvjP88eXlkoCIeXgyF78/EYHdLv//
yTAcFNSF/V2zwXvobXir0BnXLmappU/LyJgOAdsMpLulNNzk/VdLN/y4YQeeW/MD
7QBpNh0mGy4k7GG1TZjKUYVBG0/Gj1zT4N83agWzRGmpYKjEXKxcWmIKFWnzZB+a
lFiFUZCBn70g2mo4Yy8v7c/bX10VYqAZ4ohLxfxpTrEYxsP/jUsCVX3hImxTd1+S
OswcNK4uwLLCqmFYLFcRdstaPYI27CyNo8EmdW+afYzszpuof9K54HdxF9mAHSFn
0nbh1f/nlctWKItt0lBHuEIcYBGNU71JLYqtFHELuCE+WNC/pYs28zfTfa4onVIO
rI76uLPmpXJHQcTo2FzPGqfJxorXlHT/vN8Mc5+S9Eq3/gjEsiE6LrMSOPENot3e
BeAcRd6cu7djdhXYfOBn6AAHOkOi+E62h9w4hajP45oWLb1vKIxrih3xRZev17xN
YlbRp3yZmw7osxU7oIAGWoABhWjmUFzGWzZI2w7aW26/f6m1YfmAvo8soE+iB7fy
9WlyRmHfMV77a6z1VgtGaUwg12FQRRJ/83vrCn92lRbP0ZjLW1r4oFYiUF/qzRni
I57UxkrKnBY/s8TSYDKj6Apn67/9XeLyQdDGPDzYT5coY/q25xIHOfwNnU5DFDwa
iOWDhS7ZQluSA64xd6xhQglQ3o8I1r9kcHEpTzCaRDrwHZagS/hFdRkYBwd7e8+w
93+V08/XF9EqaaRtaMR7aqGh0Q6WGVzq3Y3w0nlIeib/y+qkVdOVGi6YewSeM+8f
bn6ihMHEeF0HFyUmw22QwxQWal5GdAWysAomDJXt7X1U8ZW6aDTYkoEO3MsV4n/Q
DLeEHiO4Jhb6Psr+DBC8wG5d1d2RrRvwVC2pjewPzcDDWbzSpL5J71rXy5XHcxa7
5BpJ3sq2LOLEdccNp8PMTw7M5zTTUhVQ1vQTNUYVp40GUKywYusXXwx0i/hkpYyV
/acV9wHhtT1hU+nfuc5rdzJitz8R32wIsCZiAVufexsb1VBFxJ1TXs5rsLMz/4dy
hYz48E2FDg/PIZcGVUSGGtQysE05ydpi4zUXVyXCjFIhIHs6/wVjYMHf6t6l1lOL
w+GcuwHHgWfjVQMFwrLxDL54VamN9x4jKGwpq19ZhXlQlIajnORnpd44KdYAoQwb
S8PbLRCpWK+GD7XzsdpP6kWgs9Tn9lKgiyWgD5kFAqQnDyreB70eQwjDi7eMau6c
Bo4IcY/ZIZq2UnJnXGi7MHsC8DnUM8t++6ElbOo7dkr+egRxfQIBst3529PFWT3x
l0/+Qmt0BPEwaK8uDHmkVMVl9jIiwZg+YQSU5VWFpXDc1vZaBVs0T+zEIbj8W6Ws
2pBQ+j9a3RD64jP5id8SnwUQmzRsEmj2M1obMUrD4+1yskoevpLo/8Gaze2npLzN
K/jxXj15hDyrarbXzKBgAENMtL+4XoRlwLrdgP3oKSMm1UHZGjEy/Wt3DwzBb7gP
uL/NRjicGwEwFDEqNfbRm5NMIT9EOtgeCkZs3yGQwc/9/0n6K5bygauqDePjlUhG
PpRt+azUvv5TOr0SyikJKqJucfAq3CSXwzer+dMH9k2p44xj9TAfseS7eebPZr6c
BZ1F8a/PChRYTP2js3p2vZMmpc9+eut1dj84WiK3M7xoBnq+N2IMkJsD2MmXSDat
Xz1hBZ+UUU9b0YEgaIdCgPplDZIXoF2I3U2cA/PzOLdoQKliSkdnjT1TkP6jXzkl
g/tpCljU6FtwVC2SedR9ajPrQxX0SacOnQXJPa5wGkJFalDzOEQ2HfqveSbT+rIZ
j45QIBGOZGtoeOSSYlVRqhGSnXUQl8eNntuwB6cygZcQLF1AO5xHMLJGrruof6Sh
Oekb9Ccgb6fdVykuq8M/fBjvi4iq91jxcA/peP6sWdzPpc331UJ8svWAsS1mTNKs
8Wj7bQ2BOScqvYCJBmwSAFLJDLjvd/MFv9NNYpw3Vpodo/txDyMxGNHQjJgQvNqG
1JBgWOC0by964y7HgsQUzLBLuGsehmfNu5wX6qpPb9SssHFQE1UiAU9FrQc1rxwq
oDjY6nzxUntGbKufY4buzAchrR4pzm8nCXJ8rmf1uUd5ibGhR1K51J+TIGf/vqnK
VcATs5mzqWW8yTXqhrZUXQBqd4rgIiUWtWWajdzRTb4aO/OBjuGPEmZMzUj6WLeq
EVAfdOrBiBCaN/YCkUQjVjJXlw6OSlIj11OVw3b4hrfp+RfuxnQebSX0bb3XlYup
vjFp7yuJFV+zqqXfm/fInFw+J22XlgKQXHCtsJsMr380J7JOtNt/oKpOn+GMXqdY
9u4uK7gmjgY9kGlLzbz6DUnfr1Klp+G2Ju8MgHzblJJRMci9B6T0i/QTr9rotmrq
/+zUu4rVY8jd3Whr05OaSgb8bv969ZDWo+J6UFriiUXlRvWSsblek5i7kHYWMpzz
Xu+5ecmPEgh3lRxCHDG2uk3infiTslys1Kvg+r7Qp8PpL5/aF+pjG9Sx1OpOvYZD
V9kHKgw/lPJss2NcmITNXhvcTyrb7yljsIkaAtRkmNsy1YaVjy9jh/CJJMvYMCmI
8NqWL3m5TxG/gl9xmu89jXTo0TAsg44IYAPembFesPtc6NB74eEBtcQCz5zxiLp2
BReH+y6MO09Rsp2p7xtH7lOiAzsCT9ZrszUo36O7KKLzLTeIAmChppTO7hzkWd2b
fy0Bw7Tg8wKAV0UIjP9ULYO8SVFkTVCL9bN2zWggp7Wma9a9O5jKb7wkwD8SdmMM
CrEsK+LEMXRomyDzvo05z274pVTPtKcFhVZzxGFlt2340b6tbGtsXcudTo1ZjeHc
0Ru9DJhCnxmVN0s9AWpAz2j2xh6TKC8dQ8YJ5B2DBU5EuGFfOoL5E3igGsSujrEm
jVqgYzIV3cvtABnRlXtxH9c08VhtAhf1EImRVYOl0wkGg44ObX/cQZps9bySMl2y
thLEirzl29adqMiwKKpcgbtlRTyBwW2SyGuRdgeSEhy8T03/auk/vadlGaD1zfsV
RLi04KMWSgoLhqNw5Clva9eMwgilftqe+0WRZ78gYfWWfXs1hH1w2rGh39sOOFj+
e0DJQLskXbutlC/3Em1uHg6+hv2Abs3PwDQgGimplAIHGgKPmAfT0QAMO8r3JnBP
N0ZWc9aMGM6XZ9utQBxCREkzsv6k7XPIRBVp1GvK0S78eShy2U6ezahCRaNXLMnB
BkDllz771skDPaE2GhWLa/lXleE+lkR/949xxMuSJJbZlasAg+jnCbmpWbTjMfJg
mm+0WKpgM3NNC3MihBIgqzhd3DFOMSxjVUaWyCSjMEbf1BP+a5XSsqScCnAI1+7r
C9fWGKJ9crrUs79Xy1LZ1ojJ5NLqBcnRpKJRCOAz1cyeuzpY55VKAUP4oT+PeZ64
Y+i64PTLmoFJMWfzug6Zvje1zQyCVVJsOf450Cx1uPV6CcSWaaxbzr9UHC/jzzAq
my2eJoapPi3FH0H1v1UY+/fRqVOtUQlQGZdn3qzv3q3bDDTaJUDJc0Io1yLIUz8R
77q1zquuP/vo22l3kFBBN4R+guB4GkTW7D7m/Q5//AKTn8/irXGaRSYNxufE/ivr
jxVss+XMqT9ndgN/ryhyrz9tFNbJZHe5v5IGd6ttQZfAuEr4qUbj42MgvODlQ3rO
cwtPMOGwkiVtqxVHCKU2KMDTHgDrAnYC4YzoLYye9UbyRs+TCuhaZflXvCw+tOU9
TKRRcOtMOmp3CP4gT4yi2KrICivg44ZpbRzfrMP1uCsA7UW6GmC23C30+KWzq+6K
mLwq3OaMpdGfMLW/QnRj11zWt1M6DZi2w2gtFP6W18PfHrx493UhqBDMgVyo/7iv
uIZ1HwLBMyiYlshfHc4k62n1KDRF4S013UIslvTQe7vLy9NpTZKT3fTsO9Cg63mU
JkRt8NtvTvVCvqRvK44hhgu7LooRQ1eXQ0K1C88jk0a25fKKSFXF1XdD2CB/60D6
d3nlSsO9x4SY7bUVky+aiDc4+8mynhz5p0uD3KbOgefho1OSGK5vKJo0sDhwZKbN
N4DV5FzqsuaRFknX0TJQG5vWFi4gik7qVwl0vvodDCRdYP4V2mAPCCwJYAkzreZt
DrIO+6eI7r4KZv5XykGuJ3h5HUwojwc/zmEZAN0tkMBPGATj6aJUYqJD5W85+DCO
VWJj/nJRk+j/spl+R4pWEEdPuUO8lWiFYp/PpuI/ByGJbnpAEf0YlJPWYUrTqisq
XNOPdCjvdhseCodimNHZMhpwoi2l5C7hzqrwlUUjI/ILZ3hq3ILgcSJj/O9u5PGd
Z/Lx6i9ZBAxAjhqMwYWz3ju24rmBByxfKBasHcop43VMnCNrRmOeIPIDF2ztqgw0
zGKSGorBDdFuMxtq93f3YCOBcf+WPfjmKOETBqIWwoJWbKcB3lNy3As7E55PnAKr
v72CnyoCQmSu02q3pCmG1lpq0N4cy/phKux7d46ydbS+5po/YDRDrHzkRCY03FD2
IF8l2rBfrkZxGyZrtsyhR4UVJw/q1kKRCDqWeSxEYNrf0idqWxPWnNdmsqQKYXrG
jB539k4Xe6kVwEGmcR9NaKbVgkiM3eRKBdegFn6CP5bIt+m34Uz8Hv7j3G2+rR76
9lN/Ttm63NFQ/xfV3XzmbnMUVzWioHIcbnnFSEjsoiR30wzovqwn/aEhRsrmDS5q
OT6F4vtSs+ujQzuFMEpwQeOXY3aUDmamUmHBOoq+EzssiGKgv/xdBUBUp4O8K5yY
3HBw+rVsWcvXsbHTPNQ8PR54GTQ6qiXZSNFqg8BhBI+bSefvfeSlgmUX8E4wd6wu
yHNriJLADHyz2XrIUZ7SQlMotj4VIBAfoggudf7Cftx0adx7sTvLPs6jWuhcNba0
goikWn/s3w53VJrluG8L6pD/jrjjXqD8Tpe4TI4HojjAXJuWfRFUAVIqdUYqURyt
DnwtY6GsRTuUwxYEI80IACP0CZWhBfGoXkLrROxfYOv1GO69DQEQQ2EZW5t9ugQC
uR4Kn0FZR9JL0JS2p0i/VWTDmUbEkoOaYZ1QPD1J2cCe1/fLBHt5kSGHi3iH8/d1
KmrzLf6cmzh0Rj34U/zocZX6M0Pr3bUnZF07a3NGZ4K8ECGhHiENs68iP80VQFVE
PJIb3kOs8yh0Wgq5Dit112BSIne95RiiEK7h+v9F3rFwkPVC4jdDuNN5NjM7Qi8I
TcVHYFPN3iA9GAx/Nd//6Xp9faceOykoDyAtzB+bx3z6WKSrAgRzc53PYAbGL4gi
MCsghp/Ud3wfbkrY5Z2WrcoP44FpzzB89U48EF+d3UWs/iTLr2Fyx/9iDtv4Js4i
aPYdo1lHnW9eUGv5uTd6cTlOfOnf385vtj/HVm3xxqynsWHLsJGwIOkU9mT1GDA8
5sWMG1Yas6w1dNKek4IPC1EEVjMuwL+vJaHh52Fe0FURzx7/975NVt34ayklM6lc
5XqGgpE/alD3dwyQLUpkonPEZN1rPEZ1g4h85t6iUy9mfzi7k98JI3Xnk3idsK+g
JitgDqKakM/dsd03CSYMgoV6O4l0jT3E7tZdeiGR2+2ae2gPN+7Ptb45lUi9sdqJ
iHWq8jdmYM13uP2M6fLQQU6R98iGsSoI/luyYKUvInk3ewca9sZiMJGAHMd95Ghm
KSsFxvffZlwr/3Qcd8F+CcFgnwJsBycv5BJ1YYmmwAhknQme3Ri/CWc7tQ55+KVr
vldBFeJlUhEBJTPXcU0thU5n/1HxH6cseMaYfQMHzM3+7II0r+TtKIfStFAZLPp3
r09Iw+yO56hU8c6rMGZOyHUeWm0/anag6WHWFIw7qGO6vGO7IrmXnJ5yrY/M3gHO
JXHcJNej7DXTWMfG5ZD36hkFBR/JWyVrG2CR9FKV3S8iKlGzTWyCNsG7V7aptxmT
mAwNW0zqsoH3LNUFgVuGrszKuFYFPFodMpITGAVzwaQcKHUwOExOiw5d8IeC2czx
SRyWdMkGroZPTYhPi7sFvzggkwaPo8T3sUHYeNq5zh/I3pKw//TXlVXK9MsQRlFL
+B0DD90RYs01mRhrlFNDSsGzPqk/6wq8qgWo6d1FdaY/+iT4SLThHBz1QGeQeOf6
hSiMW5cugnZqqk0sYGktpX7BhajxASKEjempOPfFkaNFa0yAWaZTHFxgVf2qoUIP
4z2+ILRMk5MVhfTUtOtt4HhZqhGYwEY77KB9wSHcErMrMMUqt/F2/P/JNOnbqcki
y/SadXoJ/+vbTusR37WmSBXLK4c9Y6jCARtc4PboweACcRQD8NOQyfKGmFvyyPEV
dqpBoZzAyVFZFqeRDi49K3m04t8BEe8WMU/yFbq8jMX+J0w7lEPi4ws6s/D9Cv/e
EiAFbVSGK2b9OxhT0JnIxd/ZKaGoxKCUQlgt7FyHrxacUiQoXNLL23HYU0VE4XNb
XkH51qPBSDv/4gnQ4Y4zNpXExcx0jABTiDx5S96ww5P92CFPLJlf36jAWKFgfmyA
+RfHpyFu8bJ+pguwrykryBFMV9pVgAQK9IHAf8CQhE4PzpIPuQSmGAS8DcPV/xTb
b/dJxR9tHdAxanDLl5jjeYSyRjtOee1DaQiMIKuD7XeGb3cN0Vl8PLfKq0ebYHrP
ALVMuH7sCv2oFis1OtUZPbyIQxDHIVyv+41BQHahJ1ZFx8DV2lxFwCGo3Hnoedld
Kh/OS0IxE9H50rqlPBny3XO+gDXOjqx41OCPfDPx+hlZ899bY2N3qyr98jSS6++m
/2NV3oxrpeUHLJUUjaOpZ4oUxjKl81w+gnifDBHiyz8iF1khTlMhe8KxceLb/cB/
sQB+JAHkpigs6GgaN4RtAHeKbwfvICrUat9KK4iprVeuaAbbR53l/T9OPort1VWc
GRnzewRgZqtN4+uw6JoNNcsyHXFBPM6ScvsVN1NPSY8rtQ9EbUT0ncEu5qh1AImn
kSjvG6XdeXWtU48zwXPmza4YddBRX+eD3e5uliCbT+IlWll60QPO3fAqT52u69ld
m6rUkS8dLEFvNVC7esOPlVnCw8yPFs6Dg87M+kJ3jLx1/puVnsy7lZFT2WKZV5/r
i8RuW1Ap8OYmpqgLMrsrJXtzZ2khPbX4qxcSZVPm1JI41hdDqKnBEoIaqboxDtDe
uXwtlVbSvOuEDzHDXZHL36adG+cd2xRHl6p/VT1r/nDvQ3+NvJZvIqlCvXIEuSEU
QqIuT3Yj1/aZErsNv7m92WFDCYZgA7mzqcQ8W9UFn/rbGQbUwECJ1+YpEYYpWofd
odiPrTgNn3oeuhQWyeVBrmGhJR1Co80lXljIa211Q07Y8uVLstwH7LcuSesukw2B
09E3dnEI1IqpEyqPZpvusrt0rxr2GItWG8Bt7c9MtsQoYBwFDu19rBRzGQau1UVP
XCxJL5zemh/BmbvqUFgXsMKUiJP7qURr5N1w33vMdNHSqOdgiTtCg0TMHnOAbDrN
wQV5Vzgbw0kPtcBOCNK6Ru4gy097TKXUL64DIJPjdbUPyzR3rZCmICZhwyPVeM71
g0el7HFy5uHsMS7xuH0znIjJI40l44/thC1PBTGIpTskq0cB3roIZQrMKfyFYSYT
g9jMai9okmW99aIGDKHJuJqJ2sDo618AJWCu4xJl5H17Rrqhrzz6i/2v0T3rzC7r
CudEWCPaTo8OhBeQVjt6i6PASTZPjMIh5qPXmmdVXEkIN1MxnR4tjPUZBQcYvTer
hy1Udc970HAncIYMsiZcN/GyNf2vVpzoh1RfG5CfHZZXG6Rv68m92mFYLh0VW7+l
dVwMC4f9+98BZ67uJfJDUzvBHdwvT+ryeEDKqAhsgR3PJpEmG1dAim77wTNuw7Sq
4W54GQWXTMokpMNo3+pxb9DlRu4Vv5+AYGYcgWCf6XO9ZlMjylhZ15tDanUgCJFP
7rKhp6OtMcJI2FjthWLflRPb6nwowd3eh4zAdS9RwkU0RPbBD7fOQ1HEHK2rm6TQ
4ypVWLMg9+ui/D8JUSur9unsHfTy/HNyIK+OP1ZuEC9YUcgkwS6YNSlbt7lBZ3/z
KbiuvZiXZDzgjHFy8F4joc0zc3s/+5UvlGu6tozqDP5D+pMNMVwHcHkNzJi8Bhwv
Vv5Gd1AlLxt/MhSNuGzTYq0bawqPcEL9nxfynm+joxsBTWSWJHclulJ+OaHNJyN4
4kE/jAbaJsbC1PHVk2UAUJR/04f2AtfdFDDJHuDVj22/vD4GzS2d0WIGNuWd2R8p
m/xFUE7T02pmagsOYx4/5/NuhmmaCgkxiMioC6zgmufJPY5F8GsIhBRXbJ2zBbia
rgdFNamp54rlSdPBDdp0tn1E6mEo09DNnO1xQOcHSlSxYx7l8/+Uwahv1SbxjP/K
xRDmN075AVLeyfADCJwX3K6z1lnzOfyT31w15jPqXj/urQzLYswcz+sMGEYlNt6N
/5izy+ZhxCvZHNqwDsMPweGhpIdE6Y/3vAO5s3ki+StJDKRPpuksjUn7D4v5DLo3
0jJRzA/D6J+IMYXvfgXOGc1499qbiiAeMyXtEvQqT8OKYQ+ON4MzQsHlzf70pPLE
0JZv1fyeRXrl7kSfJtyXy/uWsmPhv9m0IY5T+nA+kx0VZ+zIkfrgoKGJ/6cmqzny
BFkELcIDYkbAi0GBNFjm/V3Gg4Vw7XMiTDi7BWGDZtFGlv9SptiP/wQqVz28+NAN
zEYK9aQEYYV60wwbs20lP5gJvWJMiMagR3aT9H4/bqZ7WdD4LmVDkiSIPl8hRV7K
mZCmNESyIO4JFCR80j6MPHU9W+Qp+C02UEZG8qGRu1l2WkKLmK1Wwe49rwfG10im
JOtJvtCpMjGL5BwvwsxkjS7Fb/vWmmRBAcvu4og7viNtLA3S3JSzVfp0nXXS+g00
rseYMWEYCD3+nRsfX8pD1xVobNT/l6TxtQCNizWKge4TBuQTQvtEpnQt1VVqDDO+
vExuEiROL724UcSbUTYbS+bGHyqMJXGFXk7SK2nwdCVj9tW8+ufO7gCCOdwa7A0c
aYBqeZpMej2snbeDVGp830VXCg5pOM+Lx0lYbD2E7iY6MN9drFV5EGY3dQTTl4IN
WlSW12TsgVJPgxJPXs0HnWvZzS9ixSTyqIns9bHDq0ZMWG79boXLusJunsDqESGT
q/EKCpr2b0w6MxhAXgORw7RCWrhXWJsKYMRFLRSHKgT/n4wmY7bCBNGSVNWKmh1w
Jx2r0zrQ9JLpAI6E/yPKmPt6QXPPsK0KDW+Mo4ndOX8TqiyYJob+yNfijeDsLgtG
JcnX96YMsMsJpzHsao9bhYKRujZ4QipHh5qQxv/rD3pMZ6bJRIUWg6llfOUwVSbu
SKk77LtCn6rbm6T/inJlgE6NDfsNdinh9iltfBPWLYgP88ikHZPHwgEXao0q1+F3
vfth3C54AOp5MU5EKaNyOGNwpSByb17IC7qMRY7UCw65t033OEPVWSCDuyT8KgA8
i7F1uYrLPgKqvIJ927KyoPwY8eyXaSXMoWmpAt/vlR7PQabX2BJFU78gtFRoCJ86
oLv8/6y5dioQg1AftuNiIgm+TrSOFQf/8cnNtDQ6NYqvmg5USen//BagjqVn7YlG
2QjQHbPvHaH14or8v03SfRMg/bitCT3CnPgEfpwxjnBMyoEWOavPAJgvFYXxk9CY
XeGKLmU9I9Cg5jCwTdmT35gtX0MbgJ91y8qlCGLh+WcStkyFeyQyPyCIDBlomJT/
8X75+WQVC6HQB5kQ+dBOIj7ZmWSJbcwuvXfG5StKmRXPG6xyAo+RUtLRSMWxFoc9
2Zs+1dFQ59wcW2EP3UdTy7UwIcL79HXjwunPmW7PKGaRbDmBnK+qHIti1VqUy2XZ
/X357exgZLmm5pfhT3eIVs05qaVNnUYLm0zuZ8NXWHAXap7fmclOZh1Am0OWoWUH
MZ+H1hkkE5emxZ0MJQ35Yqdf2L9KTlg4bC33By4cI+/LRvitY6BcPwitbS4WlD99
a9wIFuHwWhe6BDS35+QGong9xxbV+/8CswdFW9kiJ+lpIVBjofH5AZKog3+fQS32
8uzrFGjhC0f3jovog0mCczfUpeUVwO5XYPhvp4nH9LwwwQFYKdfCJw0OoLh03tdK
Eywqxn2j9BWFWlrT/9Ec1k3FNP45lAN98bIT//j3Ab2NZ/fvucX7ZKkkU+tynVFL
1YyTxH+tS1vg7NnA1NVzsDwUjy+aYKao8ktwpxMnPjIbWwrn4aJPkQQm5MqqyR+B
OYsmmYKZm7zJJdkJ0uODZldARtQakHViaX+TvCX8W1/JEgbEJWO1m8adliVDxfbh
/n6HW2mh6DOOlnBgfZvHhhfE1tzzAsHNyAY85NqEl1ZncPHKRqyOinOEtOyGpwuM
2/9D1Kd0Kh2uK/hgv+3PrOl2dVe4rj1V8+VHmwz0THHN5r7XbPvmbaTJ6rmV8P4Z
HnQZRyE9xzeXJRXqxMvUWwANYqYUjTcrXcRByu/AwbLZatyXNKFp4fl5WRj0qQEu
Cp10o98HJ/Ln52h4VLa7H9Zs7jMAkNJtf8lX60Foa4RZopeSLfPRQJ7KXq/UTMQo
nK6PZpoTidQgE+Rc6qVw7+OEAraY8UHWD2F1ZbrJAm89/PAzMRAu/B+VbgSpO8+X
GFGCWLd7Pxz6pPbh513Xq7NPvPAo3C33qR2L412/XbUv8ByQBipYQuBCT0yLciV4
Tdaj8oC8k1yD7fmQkRP6JQXeJKXdDpr13JI9t7ZQOW4VNer+p4Up1gvOPQEzsrbK
i7cCw7ok1LK8LQlify7/45r9DSrlad8Gh5O6/dAmaeqooUTKqNKrEQuthlGHo9MD
1UHd74aFYfv7nWYjvPCbwj7khJCwguhP1o+EOuHed1UgxebfGenlVaR54XuFcZI1
+xXSrPsfszkf4f57/M4qu8TZFCYU+vGeVUL6HY+3XkSi39BWJkpiYNbO29hRLwAZ
3bjVoVK/VQaPrUjbHa8lM65A1uVy6GxlKyLjZanK7JVjU5DRPBR3SbiP/biInrby
Yxd6CiSPrYk5dMYL3URtu7+3ttaPzomznakUFUMrdKedsdcCfWvn5BJuXjPihnId
204Ee/eAxGojcYhCHz7URpVCfWN+VTIUbGRRCU21GDQRQwksXUKSAtCkLERqfecB
Nz9eRZYwZfB4jTJiNLbisdOUe94mOvieSlDhl0uobm59ehAn5lu6xH9HmtoscfSF
G+94k5eWlhCEETxrXR1/q/nZ1NW1NkZf0sWt5PBO95HbA6Yf/CXsdD9FbXxaVae+
um7IMq+gWrSbGGhyEwc+4eJx4Grg3ImfusSV+be1pPP99lYeyHu11ocJAvbhNSzO
qNYC2d3fynuvww1D6poBuuAd5jDpvKUZ7TRn+n6bSK381sIkQ6cILj+To06JMlA3
3zRy/Hcnxq0tS/LF7kxxiE4H9Ydxh600OYkYl08TWojGN4F3+b3Vdaw46JnX3tnC
zyLBqAMeScNHaZ3AzJ69O0SQNSzTBttQpR6TMFa8JiYmNDXdiZ8/zWXbi41A4oFJ
BL3HPZTBjcYunbAgZEPyn66eWCWKOsb7NeqzkczzZcRclRBgf8SX6I6Wkip1b9Dz
af2eRGwevcai71REOsgu6lT+83RwjgvzQ2BaG58Ba/qNKqdR9w/oRiPmp4RAheEf
qDaiGjcEIRggU8ZBy8Itim3u7CyDkPwP2Q76y31LKAYeelU3d7Y/Zw9UY++UXSaM
Xa0i+8pXRAprwM7mjX7Nen5zhyWWkOP+D8A6HoMNHUhuRF1Ne9UkkfIMiBbSr4ex
6sOEUJMVC8bbVxGBQ4UuEBdhTGbWh2m9ufq0WdNKMnbjVBFPfOJwADHmTKRuSR2f
FqJTtxbN0rrkxXWkBewc/0qbgGvVxrxWRw0oEpoENe1oiXPpjpf4a95rmW2tC89N
LajGU0kBMUWnIK1EVZ5g3jHYs7oNrHoKVnYkgSaTEkX/Lc8SueUdZjiRBlIefpaL
WG4Zx0eawyp9ROdx2g2JX2EmBHwhy5b/jkwdgQXE2AwskU7Jnbdorzsim/8GnjRS
GF+79zRt7d0h1VlFwKy0UgzK0xcePuRdEckXwkRwbp25tb0Zu5/RB5CPjCzbK8kN
yf52gUy4qQ1QUGkpbB/BitFNqKOh2kl0lHB158msDW0I6V6wpIc76WvZyHlbJ1UO
7+1XTmcZWcIfgyHGlJ8Sxk64agS9l+7L4UuktNhXkIml4enDZofRRMiuM5uSuMos
xKf8HDiZCgF6xfJj5RWMYkOyh+v8vesumd+xGGhGJbZ6REjUdwF9q2V/0M9+TCET
c7O34B/bigJ3cDKcvQ82QfrpRKi8mpX6BxDH18I/OzS1M/PM5PEOh/W0sh0hSgNi
/mSyWDHWnR5555utbhGm4EhfB1SB5dc2E6AzfzxgrVnC7v3DIo/JClXTDtIp72Sf
iXF5FaPFD9FHqgg35uY+W7ahBZHuI/YCJI54agj/1p2rzDCjHKPNQ/FQUHGoC3Xt
EEhvI+M4ltp2pKWFXnX6zFEicbC3iZ5qtCfxWqXS8ksXh37lZCs+xvs9Rjp8IVKO
6aw6+Iaj2PnLxk8a3pyEEN+6Ud++uziE8zLCCMuWGyTdYZIeD3+6GdVHgZGSlzfP
jgk9tY6z2AZgABr8vqCQP2SQowx8iFrGeCvX1qSisRnEeR+jfbtjEdTuzm6CoZG+
SkoXzIbZKpdFv8+moPW5j+8m8pyxy26i0mt4+042s6uBJ8dFS6yjbHc1AHOJekVp
qaBJ045zRz7gripKDTjyvWtit83w90ANN8+EiuMfgdNwAZ65msslm069B520ZZ/j
fWiHkeOGK/FzaJXoKg/SfVPrBueX/K6uBPN1vvS9giw8ivDb1AS6m61yuenEh9th
dM/F5plq6axw5Gx8dmNZDzZKxjFyEOX9US+8yna7C6bbkyJYekz6iJr3jwpPDObp
iqF27K7W9wI32wXWUgnpsxeq5Ttfauh1F+eIU4s/Kb4lv8UXOt5s9oGeVPfo2p4k
uVqH501FJ6HZ5XwX9gFCtu+b/gc4CP1sSRfZVR5mUVUg9D2OpLv7SfUnLhlZ3RJm
OWcT2W7drml/ZyzTogLBeFl1UFp1W7WkDR2/0JLl82HlFfTAfMo92aj9DX44nYMJ
x2U7iaAUp8dqes1gBtrFI+2UWoOYoCMpM89evS5ytPnfAGA7fUZH3EH1j9qBXxIj
J7fkyJkl/XyvCAecAddOAk0V/9W6Zd3vuncRri317V3aiGYHQDbKbqDjx+KT0jx5
bl8nZc+o2y52AMIX2kxw5HwAlmYLY7nFRxjLuv/k1ZADzpaihJD158xN2myQKJv4
TICetUunURiWvdwdKKn1yXApXQPGgfpVSJ9nJjix/N6Ri107cxgX9CP9LyNmTnyi
7j4O5V5I2JdaOdXNtyICqieQ0Rov1oQ2rEhh85d7uoI8fSuWr5O+4hlrpIvHR+IT
WuWt1uPGQ69zOyq2zMb5dXgR1OoK7TCHlbYGeyAYWGh39Csf6C7lFe8Dr3I5f8fA
aZxtxJdiQsStHxxrcHyLE08GCnx6KK6mG455oJCoQiCVJOnGSt4qBnbp/njmneYy
nbqsMgH9+6dKkBUKhi/AC9K+V6JFQ0ZucxnAHV4weIfpm6zaBkqTtX2U7tLTZAh5
/6C/LKj66SIbBw47WUk3fl+Xdt4PTKxHtHXoobQ4CvSAIRwSWZe6Ahe2syipDUF2
iHb+wUh59/IAhZDykmX/JQOwXjQopFUdkAYL647BQQExKdQyon1NM8EhJARibD8b
J/n1rFQDWMUtPfWBbxbKLVb3zt9RnZ1q3J28+8y+ZCl603NQwvKPahxXxHeu08P9
l196lJy1rYGngXh0PN9XA4xEePtUopZmrcgIO8eCO0gTuyuwnMWHsfoc3APnD5vY
PkN9StOp1H288FuC1DCJBv0kqW5/LxPQj8No34aqGlNIWVkhhS9+SnhtBl6uLfRX
NG92ddVxwC/fuIqe7WJrN8x6jv28QQG5prF88VsovVEFjiWUXyCoTdno8qMEtCCF
N4bKEC/wKobiocs3rbAemzWn6hJ6UEITt3wbDqrOtJ8Uu1waH9JV02KIM0vao1yD
i5xeAFzrq/v4VbnlW3ZHSdIOaPc4ZgmJoFQp+sizwmbuzPPw0/qjlSHmj+r6r351
hCbo+IBz7owVfQ/he4AlNe2jjrX/gJ9T+0zWGBadB4WlPuX4NsQw2eamT/ghxBFY
IhhsC4fO2SPHIZ4ZYV93JUWwl6XfZd2O/APPepj3JGpBIeAUste0RFGZ8kTt+egv
Ff7BPkeJFQgwAvn7hsn/nj9tF4NWq/aQ0gvZhvnzvk43oIbCRDNTFjOTX9/xrFLL
PwZF+LrIlvgj60/YcXeqUONqXAuVm5yUKWnAP+bqLNi7UzEiioNmwMuftBMZtvt5
WESz39NC40J7WZ/cEYoUjQ1q2rlVNY5D0m221DKPCD5Ung6jqK+EI5l8+5D/cpKj
0HKMOI9r6u6IgJU4HLS//M7EKEVjTTJUljgtOWWQtAh3Kq8duoTs/t/DK2WNAcMi
8juIbkgtWwQ+vtWZ/ipPEkBnQSyJ5HznQCd0xduTzZwC79iPQ3EoXVYw5Il0yH+C
7TzFRAbpA9/ZS9MtBWS0VK4tw7zhHevrHHNQQUgazna2kRs47SncFwfDQLZ9zj7j
PEu5qiQuB4e2wndSq5j8K/XyRJ68fn+Cz8ja4npdHQMVx/vtAjqWmWWIeASgSV6r
Wue4u3R7wk+nrvoe504cyJjK1sxyeW4MOibzzRsTzWMV3MgiCku6JQ0IiXFaii24
la21cmvD4u8BH3qHfqxdc6SlepWGq3DmWGVVDScYn0hcwWub50t4xsLW5Y2R9Yop
ZNlf8ukX4dbtrCv58QIMOgZgwknvgHQKtgx/8E24Fyawo33Dm9b/G/txIEDjdxgH
tEWnBvzJ9audW5kmcyYA+J4aVE98JpCt4LRVpWWvE3nNx4n3dAytIklu6XqHYc3n
I/U6c0MOfuBvCRVaIeDf/S6/yzvVHmsn/GpyCPbhNmE4baAIlA7stogcaTHALx0d
KmDBxPVKN3cr17eD2iPuodn6I6c+s9/6iya81m9wVMRcjk5fjsiZd2NFsnILTN0R
+qsDcSoZici0dWxYgKHMDePHHwTId98Z3sYSNnYp6Y/aiO+e7TRHJ6P3AnjZ25mk
b4inhy+0c9lJyRIDS8uqL2Y2Bg392tjGLj49bMDAGXPP/oHsOrHW/Na37GEH2AMW
oeYk+A9BkG/n/mH68mUQN2lAf3MGlD6WXgO6t7tvrA1CIdHNAZqjLNb7viTtfsLn
afewJRTUudJhtUkyzSXLj6lwtDMYmYxM2560Yg5hF8ALTd5Zv5Oac2L8RNFjuerf
fPmnVT/rLUQPlzydbjp9r6+RaouxEqhZtkkfgNwqWuOWIUIi6mhcGFsGCl0oijK6
W9nFxeUNAcW1S92NPVZuV3rk8GQZ4DoHlf8F9dD3ArKLRkjxNJ34LWZbUEYNbsop
GkCcf3WqAetmuvwIIwh7HfH9biwSciB75hvxsVLFqjQXz2n1zB5e5vyVbU3mNYKL
P+dCrJlafNAz6yGMgoofxNwidnyPDgy7r+P2/WLEm/23Uo0kboGBVyBhc8UwU1Ac
bSsnCBq+P+3cfvZZ/QmIeRGKnWMKEGaXzWAP5/gt8JutB9oLuWAHjS/9bquQqUXn
3Y3WwLrmlFcLqBYQpRdHT4UAg4T1miZgJR9tI6m3cB13qdp3cB2IRFL3bde1DK3z
CL1EdS7BWR1fsbAxkR/ERuv0VReAQcD3/we15zrTJI8nYCQQ1I+ZEho4A3qUwrto
zOeJhchb7GRXy409hMRK/JX9aYhInE8KQNWOeBYYzQzk9gP0f+jFihQq95ykb3wm
pzBxsDFqemlmD4mzTUu8jAciI4s9XoRN4z58L0wPQDK6tVJWWZdoG5ZephNo3NAf
5TLcsnvfLHuMVq/KwNM5LnIMpr6wtuR5AkpmWcyu8tATBJqgOJADlEY0TJpy7Pju
Mw4/StGA1YcR/xCn3GVdsFUUBouTDHnR8j8gVw5T9VNHmdf0v3vy4Xz+qYRTEfeq
UuX1MgVx1ye+6IDviemGXcFBwzyvamylfCDeMOqbr+CVCr+brCldIMteM2cvXOPt
bztu+3+lYBOjZZ/N40omkkBmg2XMBgCrOdMWajOdqoFCN0vVxjZHfX9Ip9Ph8Fp1
eas74oamhzZ5rhjvmfCklz+UQXf2daVTHQqO+TXQ59XGcBnpoEPDQ8ghWhX5CnBg
3SPiOtfSN268O9tQWYKtWLcoZ3ixpR6ZLpA6MrZj+FJJBBHJqOzhedtbWdoiS1qK
v0ScVlG0dCkmxrV5z78P2oXkciw5A9h9g2C6lksvjkplYexK7g2vz8VyQYUp/PAQ
Te7TLol0Ufy5r36cG8VPcbXejvF1xdTgqoOONiwvovj7LDqmt+w/bbIK/zCnD58C
O/PJPkMX/I+/y5HxXuqS4FyU7YOsbjCBQdXqh5bai+qu5DsvXJ3qSSs29SzpTgSj
pjCu9JOWrBMK7MqAxxpZfwKhIIEswcl9dViqeS8/Zafy6ivVHlXeh2ILw2apq0/o
BQgFDkspA55OyJFa54idoyLll2qsTfx/lxy/ACMkCL7nOOsxjH7hjWHX4bGZgIxs
c/qxeRXvY6Ly5Xyi2I/fJ8FUwOv15ni0QEqlkJXVVS8GS6eZZosY9nxqv3By/Jkv
CSaON/5P2MzU5JZFkNHGuFHrMWZNly30Bho7BrpWYjWC2+DFhsPEliuUSDlnAPL2
Xe0vUFCp48tcyXEhxoRitZZyeXDPEtAWS+NxPu0T1BvzcGyN5iZq852UGuxHTtsn
cEuOV2D3mUOrSAeXYf5DCANft7tjTvhwBh9moHWWwWdK9jnbpDal/N0Q7mXUOItZ
P0RQm3AcRS5PS0tqCYDrtbVhGwnK2o57VeFPCx2d4y/bjRcPDt8+flBKn62MLgaS
TAtx33ukBxjQ+5Yx3tY3T0Rp5IZo4OT2PEL4g214VMbCure2SZxV2wbtb6fIwaTx
HIjnrdFYuPiCkVDFMK4wpz/PAmCCcL6Lo3+4P0UMcFuu7j0k68f0yITRSJzS174i
GX0klSqwf81eeapEKHgIVb6kgzW0gy5DgFltdFNVAd7Rf7hJauoYafRIFxt+YMYp
9wReOOp53mO9eJNjx1OK8X7uQBBdC0Qoqvh/j9ZDXTTGUO2xT3H0xWydIdN/2va7
6hmdcy3vq9CLJZRgGOzMrWNIEUz2av3N8PiahHyvilV1M17NaAIQn4Iuo+T25jbJ
1WKDAYiWMPja078CfcFRdNG60GU+CAY2QzYJF6elKhBe35qa/Fu7KdCpW7fPrRo/
H/mcwljFj4EnTVp3R0Mxxbwkrjk2bcxCWiWKvovkGBVKf+isvaiWDiEOWOc3K6iR
Y8OK45nTG1HDEyo0i6SJ4nll0/O48d3ZCT3YSq+rAdZXLyufVvceZrGdCjwHC0Yc
sQTuvzlqC3DAr2mcgTULHX4D2fcXdSAqPlbWUbrQVFODztPSLupXvpUlC/NVevor
6FZFvLPCr+UoWniRhROjnesLPe4Ij8UYc7g9S7g7k5FisjuaPt3Y3plRBNJw6IE2
br+svYEPBqevt/uvrUhZY8NxGQ8bLUDevdM1ef6MayH2LCkhBNdgyEnH1IaLm67s
6m0osu+INItngnK+hOvf3tRs9qzpw4pcoPICx05w4Z7lKVzvNOPLGARvWU/vZqAC
EWA5xCJ08VWZ+V2typ0RJd0XQxhUCMoNF/mY4w0UAR8z0rpBVvbuWCMSAxI0wBUt
ZmAl5muFd/m45IHq4ri5allRfA740z7f+psWUDKK96nnoDUHKWuJhzb6ikj0uXJT
jzUUP1Scid5Eczg5h9rkUfmkZtHZ5YbwsWDVvJYLOHNjYLrCw7bC9ULvkVnmVsvC
BOQtmvFB3SZJax4+N+UTx+FZdqwlJhWq8SbRvGnVgO6P4eDO8xvt14RyB7KTUesF
sB5hrnHrt4q2MBJv6udtZ0Wn67ZYWq016MO9h9VrSE1bcm9lRyf8gRp9fX+VJ5VD
tNwTSBNh45cgizV5pD5MW9bCAeym37Bw6AYy6uasgKBuchQqcv5WcQ8XXvhM/h2N
nFIqwb+qkLiGthS70ktCNyrWPnXZog8gWBTDs9O9pHQlXkR4f89V+l9Y8D2RsRVV
gJmbgAtxlSPdw+NrreFSeOslx+tY4gHbDXj7/ePoei8t5+Zt7wRFhedmLVkuYg3h
23p5SD5J1q+qC8l3Caf2p1OFrxu1kfcvgXEEcFlI5LSxhVF40RuifiRpP6OPmsEb
b+cmjLqnEFFwnM8vlptpp8wq8N3VrKlRC0BN5XpaHXbzdX7GRRlt4wOKVq6PmNd8
xQYzCzxMeuPrijPdDRR6igbtS1X8IHsKx/8URJqHRQmUc5fJidhnbliw+UVmXCq+
dog5/OSre7amN3zGbduklHXYdzvZ+4mE+3MUAcekh8HQl80MXHQKr2CGS2GCYM9Q
doFnPG2LoaKmsZQKJgRtnmPBaXzLRoD2HeYY5IeWeeW/eFNXjPeKhsc3cvLlNKBL
4Rapg0ClKsza2Ui3D7R89AwE+w3AWa5QybqELIt6ojjORvStdaqQ/POuf+C2xvNq
bfPyek159P8xQ9HCLGZ8SV6QlCCfjY5XDLdAJY25T4k4GvbfWR2aCaZPz2z+YA3O
18wSXf28NjVbH4duhqr1/rqmn2hlpuwnWQ5TEPwDaByZwfigXhnuLWI0OufSvGxh
SPViL+7RiP7UrXrO5m7UMcMEehTmD9mbXTeufe7ASQFh86d9eLTKrkM+9Xyf3Pgd
PJBgk+AIEpBs64ZR/NaHMHaKixWQMIlUr9X+8LWCIu04QCGimwoDEgcTz5x8oCmE
3p1fsTnvECTUlayPowoJO4liRVkEdAdAUPihTLeoW4b989lL4e0vjgmJJnuPEQdS
kZuNSjQGKs4BCbQJwkrVFGc3K2/ASeKsa2zUw4Aeahb7GOyYTUU6aRefvhvC1S/e
Zf4Gne6zvgoqzofCeTxtGESQu3oDr1JnFuaxzMMcjthrCSQwhaiNfgsQUtVlEI6N
LudtRu3GAj/W+Wr5hYA7p4Eyz8yzDRofHrwZs3dE6nnS9JawMqRE38afHQb8P6+f
oUVonBl5l4rikJlvYn6mn1n9TE/84FDQbt3ujkCxm9ZejPgkcN6WdaV8OjV27taH
cdDXve4Bl90mfAm/zblTmv1EP5IPLxeR9+zftf0Rh9W4G/QP508P5WjtcdsBtLTz
sbtGXvsP6ZOnoty0tYhxtyRvRSdx5hs4Hvd4dyvE88xY07HZ5Q9L67HTHX3ViD3r
w+4HhVi27oXyYGf1eenZvvoMFWMw/bDtCDUYHlrv+fRkMEkTCfdLQDzJFB8cWe70
n5dvKqfrBcMhn17tp+5gduYApl5qqztq6YsgsQCg3oCGv+aYZddjucMNEz41BYsd
dpXF65cY4halqs53Wd3QPgbZCM4gpgWA3mNbbKzRZ+35PMb445Wv4YNJdZm9dfku
gH8IyyIfUWeyBM/R0od/4E8rk8lDGrCtwv7hFnSdvYRo0+dlQRspQWwsfvg3yoSo
iYaoLJBq+Gz3WEHOc7refyHOefR4dftQ+cRwHP+9z3k1xoRTlqZPhc/C5KXFy+4M
vHTARHreuXtH2u8h+6fbzkd/NXeLVwMWEp0RkEFSTYpxRInhzelPdjOWMXhqzDHy
ZaFMbclY/pzwmKsP1T1IoMpxn+GLVBMTTEzcp/Ac4ORC8Y2VooDyQQCrzCuMXDnK
LHz1mnNukWwN+okEbUS4BOet5euECuaK5IpzPqnjwKFnb5GS3TigWOcZ2chWXTWk
vh7aAI9ESAtiJvPtwozPhEciwPAoAhAtEwUK+k9/+68QwvqgzYqXTGeZcoa2pSRE
Vcokt3zeQBaaOrP1vzhZfKdZhMnZrOPNua+Sxipmf6poqkLHRKQ9sU4h20psCQy1
N9zNfrZXZaIJdrfSekWwooxsg4P7+ztLBBVI5AYLTICUlWisjLvFaEQ7GESJ9/47
/9o+j018GQT+sZchRv84U/NtQ8+ng1f/9T4kWXpEidnmGccGzw/2BpKjUZIWakmY
XK/JFSYVCLiMcHg/TPMTZMCyqOsz1n/2fp70lSZ4tipUcHCqYWYQcF+Q3E87fQXG
+s4zJMHNyLZEm6slHT9jnpJNRHkoveAEAiiN6oUUVSGo9My6ZvlGefibkSES2IL7
ywFdPTM00DLvfVTbHjwFUTRaJguLGNO6lOhfRmBmZvIrt9Qf/rjCdVzTe2H/5JuZ
7i1blDF+PYHXhea9kNnaIAeM3jbIRMQV6kQoATFxYVuAzeIMprLp+cbZYbblbsL0
KyMFMi3oR06tqds6vylYVHpELOZprWPc329VtQgWngjSAdohTBmU/SAC+zXPissB
saRqYzvNvfrtf+75wz6+HPU7Fma/LW1jqFXP08PANujGRpOdBIp6Nfd9kb1uYSNK
/OLwQfcW792yRgogWBStIrSv8SOiWLDqYatWBxlF6oqajDquZUNZIUERc3VtFO/J
20OhX6H0fAYQAK6Ri+147yedZ4Q18AQpm1TXcmSp7pZuPP/M+HB+P2zCb0cXDebb
KWYYr2HiALmO6reF8jD9hq0l86lXSOmHZ1GMgWx0M+Ye2MvUu8b2b3ObuPVZlh1x
mYpHEAhXX+y24+3LF60mhqGp0V/h4i0kptkhXCiZlx9ATMKkC2QrDCYfw7LVom/9
9yKm5ehsb091e5dh3nMk0P9/wcl8WoJIr4lLivNBs1TAGKJ43VGLebf44kphrRTr
d4v+ZpOxCWKOOitKxxe2hT6jalzNZQGkyPJX24yye7XSnSL5/BoMYfYR1uAlthbU
RZ7E3XMHFVA67zckXHkC/tK7nGYJyLTlpPqZahrEGmBxSOA4F7XocoPP5WkO3Ulm
ohbznMiYGYNCREiW4VljpYkVFBMWknwaK/JLCMBOiI/TRB3AJpQuwokQoIteS+jh
/8IM1unoEpdKuGfYG6EJko9Q2tLoJh2CoHl7gqNQ2XkU0D2CVYW84TCD1wC682/f
kcFSoZeVhZKbjfPrGp2YgA5MQV/nlViUtmrpeC/J1OCNgcOXb6mpNH1QdlkhKP5U
mXAxNnR81U07Sdm27YolUbCc0JYbmniQNqp7yc7x5uclJETiopZxfm7hX0wiX613
n2/lpbFRZyScgOQJ8DqHtp9/HOtWpPjNxPSmqZBF5MMzGkwoHHAMJ8YVzQP2B3O4
1mLeFQ4yV75a5VXHL233gT1L59Nweyh4epSaLOyVs/2eFhO8gMrKgp2LhlNEKU58
Lcrmk3I8tlyI4fkGnrjiMtCtEq/V3izxT7MqpswPmYNnRkj+23H2tLgPBgvniNiX
svA9bV41wjr3wTbehiDqe8Xb6em0KnlZ1ShEwyQnuTF/kWTqxgZNSTZYzmJAB6bt
cDBPRdpVpk8sL0SJzKyyRND1sZNBAuuihvNz3XA0mw3Fh2zFDt1VjkUaSyCtWh6w
Rxy1SUo8cfQerKOz78QfrognmajXk8tjmHH/yhVgt6cH8RsG2nQmNuO8LCaLkYel
iflZIGl7AK5lTr3k5NFkG4pJ8HxdUegZisMg3uAJuSKsY3O2fRYu4nBRn4vbWJa/
PIZD7RLimV4UHMHxrtbwRTARYtuRWfk/ZykRQ2/x5q/skvbGHY1ADi2pKcylr3BW
xJYX3DR1g3k+ed7Ke4s3U8hGkwYWE9IvkRHaQoR7TgcShZoWsPXjSoFbZtoO9ur8
F6SJs1ooAUDxUqbFE1FHfV9vPD3PuE1cuhze6n15ca/Grvj0fDvt1YsK8qC6I07A
DE54xzeR4mzCHVv4H8mtn0uH4mKRLFgSn2OF6MLXbsFOUSt+H61lSFyW1YyGunnH
DxfH9/AsUmLAFSPTe+ZEiolStmYSez+OXayMPEQBVV/uieYHnp5IgQ/0QRGIOtSm
e5C142xeZBPj/Eq0olp1lh9HtiVLawUmr14Q35/PvfqLRSQZvS2HY6l3rPzmcZdU
5D7iEDz8Ih64xxUoXpIYRKad3XgGzCmMO37PBNI36on4cpBZD6Wx4g9UHXFsPEbx
F/npR8gh6RjfmbQt0aM2j5igXqRJ7F7QxcaWs4UNTGcgMDIPlhoe/eCTRfBo8nIz
YGKEdUapLt1XLzSr+FTjr1/+aPl46kGl9xhNK2uSehCvmr+UjEv+LM8GU/XQiXzQ
88lYL19adbKPucjSoorK1JGUGIGsLvQX33xc9VosDXvTlnEaweHdWxBUf7tQ9DG6
bPBQpcZIhqllbHzAZey3rE2GmAAJMETyXt5qtOLaijvqbvfl9qYho0S5SHJotcg6
JMVubIAVEpiwTjpOCcPXbUyANNX4QKb6rMhoun4DnDmG6UqadfCJhPUVFSF0kwiB
EXCJtUejso41d8a3TLsgDgsXWW/bcrjdaBlHK6TwOkPvhWVyGKINnZS25WhegUUr
UnpSEVe0h+hZ1ndTFEsGLbz0pKn5sBUOJNdWQgcGzWvLY8DCHJ4m4MOR7Y/DwOWU
jHUDxqeZ2KGl2BMdo+Rc870/YpgSkiQuL9KyBtlOBST/vIRV3BSPdSq2FgNTaNgF
/HlmVWd0Tr4fSvndVeD4HUeaGUGsmUEWdbQUDb1iK57Z1ZTjA3KPT7rgvB/fS8BA
e/7yR97gVx4Ls2HxHr5c1sO7Ov/F+XJlRFZ+GaYBW4tDIaxRneasZHte03W88D1r
rUhnzd6lx9EI+/A7/nJXu5XLFm8kKGoMgPxPinzLeRGrdmLhSUH7/bQucOVCNnvU
69Mt6917DS8I/vdTtce47iIj78G6WydjKDSF26YRl1pLgh9T88JIMfFy+D+/O9mE
t/4cknKpZIVTma/CcBDxKfVepoxj7PxSA6rzmx3pKan5NbHc2FZJctxzKcBbj7Eg
jWn1OLz7prMeS8+NsBi2kmkBZohqrhyZHuZG7GJm6gFpsj/J8DN1Gnpf2D+94325
2fLOxgi3zbHKAXadeOoAQzzxLoKJXj0vapsY/wfHcdHvirXkswZ0hmWZ9tjAjn0n
tUlh4qOQX7R7af7GdkWR9VPxPGxCryFAxeUdzoMzggBo4xJ7bbsXXCve8dlLMZud
JiEQIl3yOQEI8kyBfavt3G/P1gTllQ+SwyqJOrg4ArG0d24dY3U3ybcrjiymJ2LT
cB3l/YUpdsjqikX2i/SK/IoMWorIOxsqZl95Sez+jbltwzcf1W9ooM7Kp9JEDM3h
6fdXHiJY19R9YfLOvX8dODXbpGdFH90/joLihdu3mMPjmyYjQZwhUVRv9OJTN8QX
G4RiRmMO3tBQFEILm0GfMbu8/ABRHJKq4ehyn23EyobzVzw4SIE+2hJA7DgfseX3
tke/ekF1TL3CjULqfwG+ujIujvx+hKl96Mn0sxGNbbimrHhMtjo0HfMLIYTByD22
DQDDPNnuBDTW+KGv9ee23ZHNxXahDGaLGrEbiK3RZ6ljnprOE00khpMzKml/eZ1B
kEQx0VAAW+3tTgKcZ+w8XMwI8RlvG7bdusXmu4umWpAwHmvSdWm//GsrGhnCMf1N
aKcDJKqCOA80aDZQLLQqW5OodApPxTQk+Wsp9hS3P6ACI5Dddg0FTYomxQ+/NQfo
HbPGidDVC4/X/hcOg7PEIjt1WlJeRa9QV5NcTIxzpdcrjXbna/Wn12hVjuDuqKFH
2BOC+dotrfauGK5cN9/hC6Dk1fekNK9i9gj2Na9fATPD4AEReJ4ZxaiotzYB/oNH
38KdksYGq2oxP4KDUkDGxcpTvBkNU1+hS8UsB+Qtay+W5QWul4MoZnGfhG9wnhVi
KJEG9TrCVtyTEUqjpwRUtTZOgS3v/Z6qGhS18uLDDHLbAHdtNvbw6OO9o3OO5vu+
focrmDF6KqOsUwUUduc7bM9dzO8EH+/S4Z9Y38VnwCV8HKw+4B1/66mKITZZ14xL
xx8yt7pZINnNS8rVk/umMAYHEd5lpfJZ31WO/zJt4Rdq6cJG+nCG5WuJ77ZzsY6X
IfuJ6YeY15Km254kGw29YSWe5dWrAf7xrocis08HNWm9CDtlc2eGFxkX8arWBFyE
94XnmOvMq/KcpiL1k3160dxJViy2NzCSplI24Ro6QZkRvyjtyRGzdQMM0KDJNd3Q
BE7VqJRd5fJkjJm7gY7JJIWZ3MgTe4hAY+QOfsMqkb/skfIN0rESrMNBMQso37oG
ecFocPCA/KTk5BR2g/PmVE686LTBrJQrd8NWXK8Va8Oj8GxTzNABtCv0tlyEg0MY
4qyTLSfkXU+k1yx05pqiKBbzokD34Vj0zyz7MUPRSJ0c4WB+nBT/J/1e/bs/S6Am
jYaUmX2ICp7zhWmran7hhwUgE1pbXI/DtFCE/9h58eI1rZ0hTVN/7NNuT236F+Ym
8ACqMp+RK3KlJib1BOhl6Yh4ekRbolD28RwEgDaatjfU1dYrWzSgaUnv15Iub/zF
o/0bJBelbnFbeUGdQ9Fjl/iuIgUNf6USNWvKXVEP049xwU/IrvZDACTCJetVa4la
YU8X25ereXlItK/HLEQYBqSc5fN2IHNNDYmQFeqCmM/rdxPhoh89wISSWFgeNEMW
AizN8Ep36q9w3X+/fjqA9WfQ1ayHOAUvv1Rc48MCl2UftmFBSiS9PYZMM6OgVGrz
+2FpLOA3czYvUElslk63PEHHmiifv9JF+aEnWETKVS9COJszJOT2gX0hAENBOPQz
MJ8Uvob8JkOgp1F0vkoC1f0cZp9sFJV+Bavqk7ZHNGHmsCg1zK52m5iWbcLiEwzw
WwIlAicwmlbU1PAaWfN7i+IfYMZjbJ9HYlaZ8EskzJiBX5hjXpZQW59Z+FzWO2od
DHGHLAZ9LxaLHU6GVoqejgqb6Apdkbyjh999WYOG0GRjRxFsc10VNjuPpVTbXXtq
cnK+iKgzYj/ng+ICO/lXaQK2bNV7DcEwb2KNVWGPUTisaicIFn3IwsFbAwa/bjHV
UGEM5ZKfxCdJyUeanzUSeMaTf+/fFTcOuDbdefZLI0157JR80+XaITFb80xUT74n
qKOX6gwcOyiHBj/2pVA3fsR1m6Y/EssezQ+88+JvXF/8gJ9Y8hZCoA81Oxz8CfZw
8TZT0oyvIlJOsSwYSqohYpsRSvPoRrvr7n6dkeO2szD1bfjq0vU+IxrbVT2Qdgbw
X6KxHOoKLitLTiii8Vcg/I0u0/WKuYqmQNrl+WEch0T6grgF1kH8VJ+jwsOOkt9y
XIPH72rxb34DL3Gyfn+aaAWXOycrpEKCsxm9AG4rjcSmhfURja4XLhS0LxAtj1Bk
u3eaukYnxl1c/9FmF0OlEjiAKJsQTjYn4OaFJXyd8vdZFb6NXA36Q+4v24J+3bex
3AwbXPf5fsGW8PHy95eI8yo9mOE932lTqcEBx1qL8qVFFoD6gtF5fjkdOJytX3Hg
XyNMJsDUy7RcNuCXmmIvdw8ICudEHP9y28iWN+pi9je7vEj7jPAkoFD6nzOKoIiw
wM/acTwjS8Lse+JVPWTsaJVxHKn5Rb5CWfHT7I31tVHEGbCf7WlWcq+uQex/qg43
D/i/tcLMaXEAaLe+fE6MPugjwn0zTDG9/04viRewTvIGYkCFZIdn8ewfb8ojn7Y7
6/0mLhL5KpfPUWeZY7ZoeJayIR4yF1jaDfyEsagXB/7SlqXSI/LGyY1B3XfIvIs2
iE/8bA3f1MeSCqGn4LuGPNa23ruBE9o2ccIDCXApasrojbc5jSg4MdWGSBe6UrkD
I2jR08YVl+hKL94CUwo2JPfrj3Ef5BWhy+dsv4WIwRfOt2ej9RCIOfJ+b/4GOmyP
WymoN+VEmHJom1m08/mmFgzTn1RZGSoFum8it+5wvO5rHmmVajS+ngEgMPyb2V5y
VvtGuxff/pmg51rWY1PS8JrppZN0nOX0iN87/+MpxQGlsniQeojrGtuYJI2WLRPs
EAMMjbR2nA8nUUzehn3zbMSk9ks1PoDCmkzkYk1Frvd1qfKVqumArtok0tf2LUAq
ScZXZrXFWOY0LCxT5hbk7swpcy91cHIOobB/j+Li6sqfqBpz1PTGy4hkkGB14wLp
fwT0SLBPjbnWLCkRmGDvt8KB3sM6hAcxB7GDZ53UE0oTLR58Yw880sA9CTjxsdVy
Yahppoy5XFPzjHzjQqGNhabMmtE6BjcSDKsVWKvwE2FeTxX0AXS3n2AoIBdZrpAe
BJ02EiHxvcvzirJOcqWdGPgpkAZxmyo6MNj4g6/IsMtJuBOi7IFgdV79VoVu2AlM
fwUt31K0oxlahi5AI9/4FvRj8YRFgOhAFktha0YNcuP61RGL7Za5WpmB4umupwJi
vqndJMweoN5Htgjp5b1udTUuwcgq1qsn9AYzoCm7sjDADKScIpJPPmcNOEKIK5BT
8bIMMDQKSxRtx+QpWr4ne/hyt2Dd9K4+4Nz0nG1piBN0SJEuXn0puffWj/egOkC9
j/gZ1mm/RpK6JEx7KFonzLPGhvMO/4RMTZMub3pGxzc3PvlMbtQmQ6qB+GkSXued
oVIGRNJJSKniShoIuw9eCqExO8zxtd12jKGlRVqTQvfpLWl3jZPcIOjC2nrrV9Wa
de/F9MF/AA5Xa5xsBLTDfPMmMlGgsZQFD40Fh+kxCKI0uck+Azoo/AFKiM+871RW
Uq9c8ZlduWYh9LIVgn1BD2xfJ8I6br3RJWdH6DVD0QN+Y5Zaka7/EDO9LGzAYdnj
oEbYxWtdDEfvdhV1O0gzrrGeWKk/rtCXJ3e+9JnvgQVZFCS2iAUgvBSfaYafXScb
FxnU9EMSTFufIlqF8apSyjv979RSzuA3hrjl26PHfemDHqYciRFWddcc1PYq2MrZ
8T2zVuo7ydMlNTSiSaCfDe2xbmGyPn1CphIh4PPbpCdrdJEd5aZDsZ0FdmyTLzeg
tF2qNSgUWXZV0AJ6j0tgT7njw9K0phn4VaNEpGVkqx7mFXMsCLKRRhvCEfeIhLcU
qC3GIo1XDIDYDJy+zFJyQFuJVM1NJB3Rtkz1fTb42WaWASS/S7l41Z85HjTIVY8j
7M8RhGQUSlABMqsuvUCPMnNC15R+Hx0K+LxYoRIRi/W015Vm3KrO+xy8+8hzCmWa
rAoDBGiFUpWS1mAkqMPQ+MISlPXlFAKlH3CSdqPNGhix9uEVs6AK5mPtc3/OHFjb
+WW6qZSGB2G/YvjQ6Kx9NAL33CtWBMVgv1HXHkxg/qKB4G/jcSaPodV9WJDHYrvs
pVPPR7yECnATOQZR4JP5QooVakuwM4WNAi5zNaqKwWkb+FsJWi/nmxerQSWCqKeB
rzpL4YWvUZ8Ok9m+VU7PMRu+ZBUCV793WlE5U2zCiAb5ApphgEm1iEqaflcVtST4
dQFnUI/bhNaUZzGvB8VxCDeM7/J+ceefw7bZqi+dzbgehPX4LehkKx3ImslMsKGe
mNyL5th6M1t/F89yRkkHK0/AUcUDIRxNY6f4MfrFiSDAQ5aKOyupcAWjDgujycpT
g6j4M9DjJgZ39ATODl7ltf/5d1aEmffKHrlHYqhFYTWFzDTUVeC9g+KEApvxdRzI
chpXJLqie7TS6h8FVqFvEbveKRVFJrG04qG9TcMioSSDlqUcNo5pB8tiCKkNWmJN
14cIaWpUNiGKdsDsDMg0rO+ZNOoHeobdR8svTsqpdop+0gfcGfzO4pn7UB5mflRt
ABVR0n8qb3otdHI/86ALNTlEL+zJ88Nz3fL1mxqOYQbQZbKRpB905KRFj2VLoar3
6FZckqi5VRi86AYWbTxpgk6iNaqJc0WWzIW8qTY3zh01X5reNkQiL6MStO6yFvaa
27N0/2C5Lncl6muCqKKsX0fsZFjgRb8Qom8x4DFOm/mloxasjclzz+0ml/G49wcw
GWueYKnxWdjYnb6Ss5RBrx+ULGjzfR8yTGSx0sgVmmIgckr5K88wrYEz97KFuWuC
Fz5q/hzukbgV7Oc4O/u8Bq/T0WeJ+bq1Sp/IFSiGn0WTpGfZULRlY21bcFemY2Lf
zyolRJE+qvBBrQtcAETwzvd70qQLNOMBrtFZMJ9lTte7+kcKVtP2E6aHGOg6Ny3W
PM62fBv+zVmqSjiy2mDiwvj7X0H9AU0tuuPCd8lcNdP9pACc2Wy+v7561Nh9Arr2
wH3SjZO/4tYqvA17HsDXJ8bDXWExKuZrxRM0l3KJX1BObRuR6x1NqO8yblVJ0g11
f403DuT7O6/Fds7t/SQQ1VD/QM8DDvKU8+32/AO3WWjryauBPel8/eR/bO3dE6w0
G1Dpm49jl3OK1ca2uOREWD443CnLdSEhDSJqUFRGMLixTLxjs9oNC3D2Y9G0iadc
bQrXcToTZqZAYDxiTPMx9W5BDNdpEV676/ba43d94hhgyiPnPRLjUJoufWzFwV9H
8yzV7ES1DMOMNdSS4AObqgdPfmJl6/6nAuszjwBW7SLV/4nt0GomiGIUI3EpTK6r
uBAoIjE846YmYL8HCkSgFcDLtsZPJFCZk6PuRKfF64OvHJlTtXtl+sleK/wNq64C
YJrQ/CuY33EFzk6FMj9ULicynkcsCQ8SeedBHb8UPW4vJzUeGgmkUj2hI5nH1zZa
wi8jFnpR8TuDeYHDgAfh94hm8xvr4tx0yPwwHZ8XwnZ1YDKY91Ix1Pn257oG3Tvj
A60KAJ1EVCcY3xUdAznQsCgyiLetextouuix3Qhphn4k8Z1kl+j772/piEYM/yi7
PsuQieO/6z+IVLqisq3Pvm8zu9R6IIPpy1pgo0QwSW/8Ld7vfhaAZui2HiwVMo5Q
oE7HE1/iSIJN8+efGUnr7h3bT4qJB055TWaWAa2TrodG5u6el96FdMwkY3/QOUwL
rfEbjVHtrhiD370jBWNS0NscXS7+v89hiFU7hD7ERDvdhJDL1Az0Mk+lXtsxqIRu
u7JGejYExBxQ02hwHA4Q4eke9DOY2IVK1F2Pudqc/BycGIfLPKnkSCLWIfU4eOtM
0WKBjnUaqfetu39wRvezvQENrn87e+ThPHT4EkaBIN7/UKtYWmp72gB6DTqjtMoG
rL/B1oru2ODA7kT/n7BXovG+OMvQMm51HCyFtU5sn3Ll2fkKgLD5rrj1lMuf/5sn
T1Bkpv9xUuVTbktYeh1RYJXcGqEdKZz7rsO13w/mo6RNc2XSE9C9kfLdT+iQWrNb
lT26t199kykTu1JZcDhAR5pXQxDw4u6wb2ApIa1Ty5kJVHAwuwwZ19lWRdwO7qW5
vjD2VyTL85/B4CV50r8dekoUBdNT5Qs8iUDzuMSU52PaA5DrQ+QWWVApURZ9BwJx
Ib0xp8H9hmxHw2dFG5Z1i45au0Nh+2x7SlOclT5MzfUNtY0rxkBZDKq9SOVoPOBN
uzDyR62SUdYT//mueExZpKSM7LNz7eUne3dEiY1IsK++yK7J3d3p034d1gH/jqwb
abAt4yDfJ+1oCzEajC0BIDnnETQf22pJZpRipcI6PImoth11+GkywDnL7J1wq4UQ
oztdgEAHdSVqEJlsVysUd9PZJ4RD4tLpatj3eQvKk95+7dqmSHAyVVDSCROyFch6
Iub8ev+4O9Iso1mOAgpXgeEr3UCLJD4gBSYe9b5ZX/iPF1eS/Hzhr99fAovBgMXG
JjpHl0GUMNDkHpSOVnqJy8JzMcAyfufMC6UpLrNo/qV+exvf3vn/nYDfuvspL7nN
QwnE2XIB4JmKeCNcJAeHV++K8XP6nHwNXGi2nKh7hwGNzTzJSxPnb3euTslvfant
cCGxAIrFTrat6iHbRrWlPYfZT/8P4UJ4XDZ3A2Kne4+g9779QimGUkjwjnZiFbPb
SxQkIozq+kLqw3ROKUMJrkX2hc9llrica60Nsf9MMUk65R1BntEo6s/eZpojGrCa
8/bd86LNJxep7BA/gkxLTkmp2rf+BTOESPMqMye+kImgR+dEC1LjycnCrz12uXXp
9znxaMsfdr9JAt3d/7HFHgY1asyWIpGaX29NU+avJuz2mbLHdTZKyldaOgWlsn5l
va/VCa52CdVOQ+11dSqu7XM29a71U41ZmRVCoQv5ieA+YtQMI+kJ9nI2HfWwCP0q
aGydio9THsoGycw3v0t9gAT89bw1Jq4wyPaub51VfYdROwKz/Zdnw+NvJ8g63xmj
YuNtmkKBKXhjsymN0ygDvhFK+DRpZ1TyQoYu/bsScbi5p/Cg1X/iDpPPCTvSuJPl
WtkmqydkZuiqxWgrWi/a5AJya9X1vs5nhQwm2P+7BiWXVtrp9cEvUKw/9so4eX2+
vV9gAQeGwVCwULIIdvA8MmGvbl0eCEWNvfCcd/QFfoNcAT0pqRvFg69Q/QntI8HB
WkFCV604soJg2WnrEPfWzi1Zz3vqtLBzcgQAQmn7ScvBEDXLObkDh5cl2ww4M0IT
EFr2GPAFOAJemLIUGE6sYlp3yAbfd1lGm/iT/dKz6epQtm7J4UgqWm/LHMZXtAUu
1BiJHAPEk8V41gnGe0QAagHM/Ui5wMYMwi00KY4coKD4pCKp7EbSET/0sNOJc1tf
m88rG2mnilQ5kJg6yw8MMp7UpqMPheKWZ9sSyh86eoxAXfW5L8tceGZRHIPQtP8r
YRogg/Asmc7VRBik/ooJPKEkE6DEV3kQ4QkkTNO7hVNiJCiLoA3D/hLryYgLXOEw
u5wA6hAm8AzKstpkq5Bs8WJj2EJClr5wM3QvVNwVmHWiqzZj8WCAjL0gvaJEocBW
4JDNGHlIET2ZFxLhl8nYx/vBzZKgudtQJJ5AHxKUUHd4vGKOCiri1tQ6pKgKpO17
e+Je5mwEphwdN+Dw2Hd8neIbOD7rV4lJTHs1QjEepYFiG0CpKy5JrLdQw+3Wmvl5
gG3UcCLhPF2PfRIkY15kWw2cNF3lLsVXWGXhxWFcopbgis5W0rvFH4qGfCg/riuG
BwabxuFJmRkeUmfdvyZpRi8JrHsdNammyM2BlzAZhEVMaE0/bNG+FHFs3nq/x7a1
UwGKa6AU9EvthPIzjyGgdA3QN5pcpQGjYzCta2wat4S4zwlGeU8A5SzmM7cRv9kM
KHSZxlWauaqWG79TJ0n9bFvgOGysdvHHnSCnoVrdTsMCNtfkEQOE+HIBLZDERDi+
vMnZ0PsSdVeTIRypwDIw07uswyxo39CtO2EvVqUVKFLlBSEiuTKSBojP78U6yYkS
AFyvNqPOMemtnf0zBULGGEIZrTPE5H4X41UHf4Q8foc8HiQAdEpFuujT3aRvjf96
ECtcM2OEkNduEF9TMTC9mdbCA3G8Yw73ziTULF7+2ShX5OeEoE/bafrnmh8+3x+U
X+fUMK+xatPj8Qv786Bjt6iDO7b2ctF2c/+KrvVQG/5kyweAk+n8a8m/3Neeetd7
7lj4YAsidUcWwzOS+/5qymGK0EERNvob8f0eT4E0j9C6Ctcm3ztjiVuRDFuULr6o
RXpAeOUDXnENKS+uz1j1/cPnrmTWVqx/HJvb1YHbCB3Pc45VWeDhA430OxnEm0L6
3cCOoBTQazMbpKX9+GS3u8l98k4qb6ddLo13ABBAZ3dzEdoto6lrjdVw9ujAmXJI
zKNf1vj8TlHmTdV4n8ngam+PlSGpw90wDvYATZn3wVExvjKBOP8Mh7VgP9TbSLQh
xWHtOsvhLaBJXv7WKuk6HBypciMNK9/Tux5KEIB3CXBjdl7P135reBp3cD4UygpD
HHAebY3rFbDtRliWK5SMaPpZL+HaA+Mx5gKO2xOk9GR4C3/ch1ZZESk2ZCIvn2He
1qiokC41RPIKMtgLwfczL1air+TNwazak+3nBpEQdPY80He4QhZTNXSeYqI9gNOH
HIQ0IxT8ZSoV3XRGbvylWQKKdyJF61ZwPGl5LS8iurNVYm/0iG5o/6Z/yMttNtHM
V6iyMQPRiXxXrZpq/yN+cxlNrqCzuqzkojJit37hzbz+mF5wXmfye7rJHDV0IP6T
j2hQOnh1rV1aGMFySPVIB3WnljD3cIA5q/lBCb6v22e1TP9UuLPVvnMXuX9URNRs
2vpyTuV63HkEXUKWLI02RoIYEelM+e6qdbkyZf+FfEzFLlhWH/yd4Ve1++ZekY2t
MdxR8yAP6KW48v0VD4OAlObPv2QN6NpuN37PqFy5Mb13D4nrAKzvcHiyRdRNT8T6
vPCUZTDMYE8EW+FtyTQxcoqdod4C8OyULn6Xrq4qhYEs0HlN96Ib3vVA8JfTnTmV
qvifmmwMfmqYSbtjP53vIDWMXDqwnsDj9PL0wVQj8t08eRQV/YPMGmK9kRFqkJr2
gJ4iqyItDPUE6qwZhVFt5PzgmHhZucaSY8qRP8W5zuTS1VKRLO/U4AlB1YBZ68Hh
kZYw+FCb+c8XtwPqWwB7MfUj8EG7WokHKUPgM/1+oJQBjKfJdP6psxjPRTEbe7uB
G3GWXp91fpya1xi4xazsfXcGbksCyh6yMgrEtOJ4/mObwczgQH28pBPuka8muDAB
wb1IalnZRRdQJJNXWMjLSoMqBTFGkkzOegQaoGl8+AEu+PAZ6HNtvFx0DCM486eD
53e1jJ8MbRv0pUYfGTmx/HE8XJbUtLz9/BPVumChr4Ktk7Umd1L5TdL+PuexhGTH
dILA3aLELLEYTvBSzKSfn8q4F53RgNPOEqRtKZygtadOgfRWDvF5YHoIt2h2/aLv
gVgUixVzj8O6eLaPa0kSZrr5U2mROhKPm2UMQLisush7Fiypk8b7GKwFB4ZePnOO
2etXUtS8uVLO23PlKkk4OnThlSPrmarMnEwdverKZwtC0QP92LaidoSfgVfhIfGH
u24n/bRMedSfoPnH5T8+n2qAJHIa2dA7ywaaE/flnclfTHuYifFtHWEXtq5HYxpC
wBFriiBZYdgywTEe5unGSKdXINbnz6Rpv7+O1ys+q2/lLSGslqf8CEJVzfLFZ575
9FKvf6bbgix4JAS4EX47dvxWMhCcj194lJiHsH3WXoOIHT37wj0kQ84Tm+CtBzet
8rPv/+3I2SLJDgPQeMB6tnJ0qrn7pCATIPxeOL0K6YkjfXBEZb6wTIufl87QaA3x
MHBaPEx46PSpHku3XhIvpr5HQigrinURZMUTq/UqmycEshuoUfolYtQQwwXxHaxP
SqP68y0TVr0YkESNQ8NMVDxLfpbIBKffzCnqNs5/mlv2p5tLS1XnKU7fQaVEJzvI
c8jEPrIqQKUO2a/CeQjBYPXd3VcRlF5J7ThBeW3tLd+94tlq3AQYsQZ5lJSFD/wE
GNk0ovzEnpXRqgtQhvFp8dIWREmbIWDqTphCMqqoYfgocU7WwLfbvHQT8u2+rEqg
QK6DRjFFH62c9AHwnFPhCkGIsOhhRtq+3QQFRAvGLfgWw31vqokZQYc7CRbaKBEd
44BI0rPAYqftEprEk36nF31ko4HdbdAR60dSi37sqPVvtkn9azwRJIigdJYU2Wk4
SZosU3+BEqgYlO/ZrfI/UW27cco98PyGz5UhS48BuzZt985FceRR/z7WKCg4buFt
VK+zRULDj2j745vdYNnmLHHutigcaBctcrLW2M84O/KcqpIH8Alwuhzo57ohLsDW
PXBS4fzjemUzAl9j7yzsYPTFG9yiPiASONTeLxdOmga1mCeg4vr+4j5phepL+753
Fz71dCQbMpO6+2nbKkcQSsAYBw7Sh5iiFbNNqy2YZoaB7EHem2QSc2sHjIFOF/jR
+Fmig8dWQnCbzZnEJ1zAVHj1ONq2Mutp+bSLzc+8Gu1AzimjXZDW/UxWuCSAUHWC
lGOwxXpHO0kEfwon4e9nmZCelooPsYkpJRM7t7CtqYyUSgix1cSwoWMOW9B9whfU
XgSJ2HdCdWPWdiOqgrLzBvruY/1AOUeumCCMQNCr575WbbyWftT+hZAdYALVc6Fk
F0yya6rDJlVpT42RQpHPEONydvD46TeFVBKBy8zVHHNvM2qEBgkKKD6jhfTYlITC
0YWhGqX8vkJ5Dwzzm6dNPsCqXCtjGtzKfLSo0KpoCxWO229PKq+7bbGTcP/FImAA
TtteWSsb+l7mIW8qvyGDEGdKKleynoUyQxuXL1FFWQEfeZk7GbufCxHOw1SsCjq9
viIU/+nyNIMkymoUm10pvwVruOk4gX8rihtxbItYKpwRqwqwS/+MsQ8hTPAxGo6R
/nlnHEEGF6m3uQFyCRfiIlQ8jtQpuQ+CcEhEkhQ3k8z4PKoN26toInQnA6WXut0C
sTPGVjHctk66Qk+320pVKE18Jm2eoVETsmtihohEjk9feh+svFysaQcHVf5fyJxR
D16XeizurnMR+FMdC1qxx5CDefRlQzokKd7Q7hPhB+omklIGrnZTstlze5xpxyUj
2WzLYjU0CqZgPakf246rz80z6lK76XlNLNCSJ8/cv/wMhlMs0jW54xnL3WFPQTYJ
toFZSZ6CyT2YNu2B9eK+/LiuO2AcokkhtBrmD22Nd0j71MNg218TkocWYumd0jMG
2n76LyiWXVsp3QOHnshcd7byx1TONP0S6njuQSSFLEnueMeESpPsYBGtT2tvLWs9
HrsT7fVbm+qwxW2Puc3hJ6qh1kM/z7Jff7Wwo5GBN6hr72aP4JWmO+Fvu7rU/f29
WHpg5CC5UzCCApC0XynZEDE8AEFC3fz1R26/EL0OofrreSRnyYn6OLOpFUUKjYVc
o3mcca3rMDTRNQQrmw6/+lYQ+jMbmPYycdgMn9E4Gt/TvugvBD3rslN2r2b/HXo3
Gpy4F7hyzZjlLQBOcNy4OhO8moZbmyapjDb5lK0NEwPoyB8KzJz43sV+usPkOrvC
Jwh4qsBoLoBzEiEpwipQwNOOtcnv/43dI5+LxMZgnvll2C8B7ZNEckKgk7ZFTIQQ
mEADYuJh8TesMeCmCIS0wC4nSclzMlmPnrJ6fmgjXxYgqCMYYyLUAA2wPkaj3XtX
Y7lOCFrZ7Z4N0dIqoBzcy//Xp5hrJCDaqkxUDqnEjPzgudUtZTG43xP2inhDVdqB
e5tpR1lY54FfRz1Nbq9QzhgwjvMEUGC6vDnyccNNyoPzdiP2wVkmWBUYlZMRkAqb
L4u4MKwd/fpFlFE62jxIBy0Hp5hsMks4whYld7Eh4rIT+n5SM/BP/BBAwjtilnz4
qBdL3NZ98A8V2EWhLoX2utZtYxT3RE+FuvfZTuX/Cqcviz4wOqBzLWNK0+ppTmSB
g990dvDdYPoT73kWOfpC03Je+pOsRX7Odo/vlJd5FlG+kERAsTEDWj+wTtl35byp
XiDjXeu5tMEDxyRPs2107Ay5Px9VNM00LuZPu3MZAuaX6HGJjWO3vjmgw14TM8aL
cGx/pqpbOQPjKJsP4fJLOBUo4mFp1VG0MMukn9SVddS3jM2ad4rvM6a3Cpwb7/+1
iy8JpQWy5x4hV1cFEwfziauBHo1Ea2TN8BfGa3lhxSKnRTWHZ/3TxY/vLOv3r/iz
m19ix5P7JLHCSe1ZVc6Jnsdvg8eE3uNHlyRrnfm1/ebDDap+JLSDNXAQc6u1BCw4
hIVTrLGOs8RmyPJD9lDSD9tSCCaRJiDHF9ZPZb3ZI1WI2xRzFFaAG85H6nGHPsoL
aT+G4iBd+gzWs4lEW7L7HbOxkCdWNab6dgT9PtzjMWJwS+kYE40iIn2Uw5P0GIgu
jbT49JtqPzNY2kquRhDQ3/rGKi/GHLqKtTiQbtPL0FWjdSSa6a3h0UctnJDWMlrn
wvEWgKq+EEzBb+yeCkkHq+vNlNtY0zylvRPELlq1oRJmm/JT+NqEHPY+WA5AxkaL
3VyqhdpfKZHDYG77YqmOUMulJZHaSc7VptqHVfE+Wp25SPNIwfnqv2A4wsiDr6Xf
l+1SqZpne5GMEVTLF09oM/W0pdlr8vM6+FlXME+tLcH/s4VPL+tajshumfPL1X4+
+WMYiM5zi69CpGq7IwRbNZaBY5vgW4cwvtqA6Ed1SxPhHVpURZRYeLGnSmNoARJk
RSHkBe/tESEQjfxdFLRv7YZkP2dhQHJnq6yQWl922RK29mK1FemaYdcJ6H5yGmzN
Ps04WiYUKTW3ep0wOU+J2ZdIpbcmzMUCPo4Qi9rcRrG5lC09LhDz1in9ZzzpqQ0v
6X4cQPLcFRW3tiHiIeuUMBSNHiBwCc8TF46X2ZBI5Cc4azwAL5LEHiV1eCW3Rb5M
YgZ2gj42Sxi5IzWLEjd+2Xn10CwY9bqVFbkBMRRU9ILcaiP6eihjEVTs4EwbWq3C
Ys/SwvUAvyoMS3kJMcdLedW/Unk75VPRsw+AkN69b6hfO2qx1bUtVlT6uYzAuUre
a6E7rScbMgR8ZbjHQYeuwII/UxcR+tPFU7firP42fzPRQqJLAxFz7a10vpWa1bYH
UakX2GWaz8jdUQvXHxeVIwRqdop0vWI6EVh31MPqqwQo2yoH9ebySc2qUlKEv8BV
MTyh8Eusalg2tXQolAUh9kcIutnj59s66LJKCsmkJFwNyDswZd+DUyHZS2b00h9m
hfVOlmq0UPRnSlNIpgzBA8yR75+zeiqia+wwUCP//V3KP/YrO8p9F1wwe15P1rDW
wLi53PCHYCJYQUzs5TxUeP2qlRX8e13LcHlFxSOFim/u5GWq+8hknEKzJY+TFx/h
2dfMyQ/Ibetz2DmbX59Z5t32jA+I4ka2ezG0SO25ANgd8JPeZNq+y+YDt/ZXtOA+
C/ydRhwc08UNemN6ajHBhHj9dkjx9xDZ7M6M/aygGnP+xL3waAptc2hrtrZGFMDJ
3MIJbaeucJfd8plDIEoa5AGS1qrZjrcFWKRxoZRq5bOvHauSBB8wAuPN+Oe6zVtN
r2ppw5U0uEHA0Ea76w+eimhYW5cSfwgojV9Mta2BevD920UimIRzlUJYcjZ/xhb5
LLgedOvp+98Gl8IpZVGtSTima8e7HParLVx10eim6S5NLt6i/UKyLo/cW6Ae4n6x
MuYQYyMEWADhMiTkpy4wJZgAMn6L1lyh+Q0Lgv/aFPd87fT9hxU0WE7MLYeQPI0b
VbpO9bkG3xij2QzpS1jJER154oDgTE1TUrrzzLByctWRInwjLGkCxuTsons02QEI
EjHNVlQ5fFJgs6LFi9LhqXQ0VkTIV2jNyJhjso1/c/rw/JwJlNDh3fFIbhjNqjlb
d8iV/AIFRnBMnWKzxIajBAdgzzW2oWb7D/RMWOKv+C204i4KvU+SbrTZdSF72QQf
++sWyNnsq78eNjGJAUjlNPvgFL3G3lNl7lkk/EQWr+it+uiZrOvug6YrwF6/i74a
M4Zm0qjqBElFKc2DTj/90MR8i7DI60z0Evdkc5mMCqzS43/SVy0x3OX54/LKawru
78loUOCBbSZBjukmemgejPrc0CHchd+kbM2YDpW+0MvpuP+7uE0wsnk44l3jZ/cI
OUQ3ExcomlVGszWZOnWuQTvq03aK4i+k5zoAy6T5Rvn1hStzfbie9KFuHe5I+dCw
CX/oTiYggItIfvcqH09Hv6yQsW5lMuw3JRNAemcLwYDiTEqkOaagvSkXApXC2ynG
gqeeACdXDbUMedIaYFJ+g2VMI4/fETss2oM3bswPh+B2VMu2azqXO5zT9KlJhsYK
BIuMkXN/3yNLHDNm15i/dONveklt7VnxyBIfx1kkGtDCbGuck/o3UYtXBuRZsb4Q
Wlx5x+T2vOLcDCUHn55/NGi0HOCUkE23zO9Iy8I64UP+79KPZp94TgR+J+KW8H2q
WKX0HXz0umkcspXwGa59K7jOBwG1DQ4Dq6i4M2/bLOw5sUsqOiFy/Ukzmbg/iG3d
ZyD1ARDXsOl7Pz6UvZxme8mhVyi1xt1R076o/G4BM1FmSHtp/c5I3DCYxDYE/kvE
sh80fnAFoTkg1w+eCP4zNjX9PlUoJbXCXIHiLzVguOw3hjQj5vhfYAL6QGcWGWf6
iVQBmQF8EweCGWnIM7FyTdDZArm3ny0vX3GV16FW9lghJrxzi7wkgFd2m5l4kGH1
yM3CTYU8Z+xNo+exFwmwGGk2zYVL2v/nVNPok8Ie424ii5iF61HnUPqtGN84DiKB
aghg9OP7bS1M/I9L9z368dEFAOK7FPvAHZshszhVKs0kBKCaT46IWTMvh9uZV3+g
CKZkkW1zZkDY9JPFt20Ay+MpsjZ9P5/Nn2looUPrmBQHNAeXRfZ5zG+oixcXxeGZ
49tW52MTw6i3lgbyk/nZobGnsrlj//V7ypBSvD6N7C4RAZXw5raCabLSQB5Q+6BY
vAgWxEnqYZ7Y2Hd/NBFOmhOg66Wmr/wr1sj5Ub4LXnKJU3ogbUlPUKglbezX9uBf
HsEEQl6IZiN4r6uhnQ4ZcZb+QF7nfYXkcSTqtp7xcEU/BeqPnFthwH5XjXygy8nW
4p5c3rBlxonDQogjEYZV4ZSHIJ3yry45w8cFZMSdzlc8b9X+CqNqygBlwIJb0wpc
mxWP7sAoCbzZ+4ML9toBUXe81tEAbtsyAn334iBOuwCWtJTFmxsQwqoe5ashEXE8
j9AMdMfQQ/spg6RvWlXK855S20unUTkAVB0Va9jBJElLFI+o3qliv083c1/6/092
nWpaC7eIpKT9DNoRtxLcS2YOpyHcwead9/KJL4tExm3N61k+KFWz7uj/jXTdSZiP
P6QhWVleGn4BrKqvoERvIXctZCbrpDWzX/qsA+06nGrJbl6Gri5pF316cbg7BWvw
8O+ODSaj4NdLdMCAQoAwZvhABHilRy7/y5uV4an+kkNTNq4oS861s7rlE0/o/ol5
5V6ku1Znry7V8liY4CtgmGZkRHvoeGcDV4dTJiYPxky36cdilOc0h5GpOqwb3MAC
8eCxpZDiARsnRHBpEMw2F13Ya8YrYts1wOYhqrIWwqJ+JU5YVoGvj1KUzIYz5T/o
d9GOXTjIZcRVGDm/J9A3Cxp+gQ12AOQWcMM+rv6KrmkVoQ7tJnvbpKUzMuQWFIRg
EF3X6wTlzAGjXCt2rzBS0ADc4GUv5lQltKnyn1j7nWu5aRIYZt1o2aFB0C3RqAt8
Rf4V0XFFIsGr1Ox9yV0+jlAHMzBMzP5JNhbtxQpi+/6y5OgCqM/Vq/Ljn6W3YJuq
FSn0nvWM5s/S6WImGVyUakzs/MXvPxIdinWgKlyu3uaQGWkLB6qhKO+o4PYK8QBh
rSdMz7klyS34exTPiX0ck2ifNP7Xnu/HGYV9+BVxAxn7SK5Kuord94oe1VKQGzij
1uvZALgw02kQMxPq/pZWTXPIQGoQGKKhptV74LiS1niMDtGh6I2MZEQGjAuz+S4L
gEjehpMrUf5MJ/DGErRFtP4SrxUBbtoCMPL77DG7NRI3+7CEk9h7utR3sMc0S8gA
/d8IFLbldO+y75tg2lWV9pO5cdL9+SeV7nReSQJspjU7whZ9KNHTL35+tZuCmLZq
LdCRrYIra1cRS4lF8EAfc52ia9cloe4F1MI4b7x79rHd/eRrGCC4mHxaF310iWgq
+AcsIiZ9/Xpg2sI0M4fy/r3mVNOuV4YeKCzYrhpizj/pcTbiQ14ZtEyPhkziF2PL
tv8Ui7zzvgkkVThh0jzT1KW5yHG8uAgyEH864BETCZDXdpsRi4Nve9kxk0rKla2Q
ZY8L7oB5GD8U1pZcv5gH/POXq44aKHpThdWJTuJa9RVK0/lfyvFWf1SXyLZhqKGb
iVQViqEqzWsRYWRRO2+fJyEPecG5/dywlvYK52x5u14VIrVF7h6GvuQ0Ws90poTb
b8v4gFdbWJZ1y35zMn+SBnjSxm753WS3D+aTK7ijLloG47VKDe52L/zyfSUUc6Lf
SeXV1dWod5I1XfQCT4ZrjzUgwMwmaRhp848Ibq61PMgFSS+L4cE6Wj1aWyOGa9KD
+O6ydr3pJcnHuUzqsw9KbJeTs4cdv0UfaMCKDz70YMurDjam/oDwlmsQsEjhT7yv
LNAARz7qLsLM/b7aLcCVOURNgx8tm58Bsxdlkqjli7Hp1KwfDomoNUHxKIvWsTV0
e4JHLp21qkB3TQLDz85bK/ZcbaDwvBaSfhwMpwc5JjKceDa5tUFKWqXh6Lzk9op5
1RUbwlum0SKWCqW+ykl0smLPScOqfXJWGi1FJ85/cgILGzrDMNmQzGYA508a2SBV
09eiko93Z0cwOZwcOP6DtecW1/nAeKz2ePsWNGGNQDyga4Kzd6s7smFveiT40CsC
zPqzY6Ww0ECAhiBKKY0VuGJfjv2q8VfWzZUAoiHzVSuQOO23KMBJE9MnT3PP1F5s
QzHB8mDSFEimqScB+8ZZyeovtfFueSk13SFRAmaK7m6xMcI+838IKHq8foaGYT0f
iJO01g2f5gnpRVnBGUxGhx0JnX5v+N/p4hI4gdjv1oCBVl4hIUBSB19v0oJTidAO
SFYQXzyRd2Pj5bDj81oj5KYnB9g5UZLQNo/gOiH6KEQj+E96uiWeYPo+6/u33Uad
Pqp7+IxpT3EhNExe9iAwyW/SUvoAL8ZPFfKo5AJ6zZ4tDx2DmpLSTbWrbUd6hBD1
wSmrbXnXI+5OKepDgudvjyr+Q6qM+384YsSBEPgcKiPTnQAWHfLAiKJG9IpFbrXs
kxcDEY+1csGadecTbCwEbanGph8bcPMCWf4elXIRfxDmRiziU+xCfhJkOLLCRK8C
6VQT8D8Tosk0q+smi9rJ+MqOyf/e23Ftns5noN6jJUidpWhsnT/pcORMrErZMB+k
Sg2b2AZ0bdigw1dtLRbE3oP5TQ6IHIiFr48X8aWlX9B9TQaN5Jld46hoeoBh1rFo
FCk+3Ye0KQqO4vMGSD1iqP4yP2+m5WN0H22Lv/Uwvpkm/W+FNzjUeOiA8P89e7PC
qGVIvkx26WIvlSRXX7PpEiIYCbuRqYtAT54RtAVB81YSZ61HTby1oWyyaaslPb3I
gWGCee0YWr9cNBOrxBhD+Qho1G8cNzx/S00HrEHudOwDnv07zJY8aENIFFaTZM2k
FS32RoaMJZrG5sVSPqb2tyMok2nbxjHjj8lZ2On1blc6rBbgKRKKVEl5uQD5TQvu
+OXFQRTGukWptmEpU9gDeoewEJEEfhrRlgEK7OiSBTlyYwMG1XnlRpDWUc1qbl4j
Gi3EBRcvAiCQI4Z1AuFYC08Z91yQploq+5ZrO8d01BtrRMo08OMs3j3lbZiy4FoM
Q9ZrzdzXea/spoCN4Gh2ZAbS1qBAJKZny/7JWin0PX6A5aXHpiiZmEr9qZMkkz7V
Jfd/BK1HiyefMZWuYquHRhaiCF2iRRtmrdpoqb4rGB338eumM8E8fnb7Ak4Mdvne
YQdlsJ5lvLF6gFn0GtYjafLen966Rc0kmvRMw7WpynozqLHJpKf2L+Udi+LhEARn
KwsOemJjxVUGvcZEe5VsNMuwnwaaCe7fRk5B4O3AlmW11zju99FqjrYwZbH5QUmn
O6kxa/ARB8ENOGzd9MBm1Qlrbdcis0oLjtgbH8ccPEAZwmMc/ZfdSlcmNAegEZzJ
QWctT24hC1vsMxEQmHbo5MkeCnoVQkF2LvtT3N0On/SocG6An6q+ke40fo5HEMGO
+RvLyseYiEb7MeXbyPPJIUFTUGzNAQLYKuaqSpXZL3Q+ogGAC4qu0QdeCEzMI4Fq
9ApzsAP6ZIvnA6DM/IdYs5N5RvcDF/OexdqonqFsm+VcJz/OGhOL6RmYiO0wZLiZ
fwLgGU+EA3hKSmtIj2NECUOzhPDaTmII5T1YyGhlCK0gsOG5LFGgCzIYgswP7et/
C+6H/7GvGWkQztRrFG4u1JywSaZl8fr9VAR5RqhYG0FFcDbYQxVCjhuG9wXOaoU1
aNCEsrSQbcM3KivEF3hKa9vWQa+RMCcYmjEoVO6LmkVaYah4UmxwclP1VBvFpBPv
P9SLABGkG65ZEKWEUJYAt637qNc1ZlytJ5LfyuH++i6ZY1yMNS7CnLLw2lNDQ2FQ
xLwt05FhfM1ELaZC7k+s4nxIOpTo+y4WaIDPOMAVv6FIqRQiUB5eEYjHwAfIME8t
cXBdlIaKQNR3x4cUKeVDU+UxFiWPnflWATlXw2s2aKdmdUqq60W4TTGCS5MJE5zN
M6ojexhL8TZlYSQ3WcMzaBQLjt68XXl8suG/x6OOhc7yeNYt/r+ZgMjB0Bk50slW
Ah4yI/KosTzlpNKMBNng2JY2np9iG2bMafg58No569jjDpulftF09A9MiMMxvwrI
B7xJnXeGUHe8wk0f5MqNKE26xxcYPUG/tQJVYpV+E/VXj9x/orJs/T3R9ChjeJ15
XptcWX22U+oLG8FxsKbfgeg7nYiAyPksbJub5z2dxCWTnxufzfZ8LR8ZF2sMXP/f
sM0NIK77U+QNecJUCN5+WbBEJfEEVOg+MMrUJPsp3H5BkalQJ61x21BfWTf46Km6
Q1IVB5QE26EHYg0soE9VzNl1L83DVfzQqhBY5bkTOIyyDnnlAsyfy9mppgQqqIMs
QDzRlLPLsrorFTTwp8APt9woprJQK5ZXJ4e60JWZvKDFRNqg7yI0VJI8DmqTpHmt
Ol5w/GFbsdMsiC5ka43iCGOxT+aea8A4v8AasanZpNGVAx9aO/kcNyltLnaMJ3eE
uPKnP735dQ5UWz1SLXaTCY3GZgnFPPJTbSOVj5db0B/DiZyERxyxthXMpMotjUCy
WcXI4rAHMtiz1+ihBu9uw/8Z4lZXWnxE7R+pNg1fvirWF6facoRGlUVyg9BNqm+w
cJeXXZpM3hUKat8loUUFrPg+FhQLGqbrD7dH8hRPw+8ww8Yc8AKDb9VwzcqBKrhk
IAcEYR6fM+OWUHFvHmUBWRYVdtMFurbu8UZCjCGeBRYBqPuElqE4hgsauuWOrhLk
dV/K1xe9u5EQtdPSqVSnS1VOxuqr9Ai46lrYSQZwYdjKzT9gOa5ir4bxJjmjE65O
6OcDUC/w8u+xDQRRp9MUzoFmjnbSIljD13zNKhS8bpyJWpiswVS5um+U0x0x8Fmk
4OZL5HcgPKmyHfhXlGi7Ngr9ejxXkEjjP+kv0uOZhUh1vY0PM+Y1dFQS5nAfgbZv
Y9JfvYGWknd1xQFvL24vEhko9McA6UP687BcDWbMxWRQrVAsXs4X9VYwfYukfI63
VRGH06VaOY+VVXEuliQGT5M1kQn908WJ6vidJO95exyPG30x6kegkpsH5qZaYkGh
Yjv7LRHJyTZfEJHdGyysqNHT11k39Ru3mlzqvxMH5Bet+EsvrlHaZVS7yOQ3Or9O
VrHmn4+oWRZAAgbpdgZzKjUJTulFwnHZuv7WT2dJsz7TjYd1YwFtxd5ieOYEbEgk
wrBcyLI0Fzw83cS4+2iJyLL5uuvfhNX8nJryjPuOvOLk4/KRDvXviXtyAGBlZnZA
bISIL0LGJqsYTTVFXkdrCcAhbmmHbfFddJ/+Yj3p7wlQjHyOegIBSvMyxd6U1iFs
eRvNvKYHDIImtmxWkEQtiOx1BPnKxMdr7ggPpNmM4j/Y1U+V3kfItyksc0X3PUoC
VDT7mjmzM1IE8sT79n55wCCtaVm8w7JDuUTGdC+MfBkpAxcL8zaQM6EoioxLcQo1
6fiADXH2SOytrgqoKPtrIIbP+wGv85ie4+ThCvcfaW8ZkdN9ut1MVeLc3bS0mFF/
zgib3GyY4KCQiFKR2bQSGGXdAfi8ZJSQ++eeGP1LP0t/WbfLpqcYawJWTzJ/7o9M
q8hvifFsWGvpgaTYkGhSVnMLwq7TFFwi9NJM11rsHhqPK4FTE/z+uMGPfRPvbge3
Fkgy4n3Mj7DCoCIkl2MMkZZzKRZWwcHPXrCA15Z63pisFdjSPzr1oa4y/WlSFI7O
m31nkvon4nUEqDjUNLwcAk2BwQSoS2BfcqfynQcvEfdEXjYzTD8zyv2UhFHw4aQX
R5SjeoQrbtuhrmDHqj5ZJiyRpMIN8iPUmf39d8QoSbYZkXfpxvy3qpTb+kxXNHML
FZF8LyX+AVOMjV/dZqyJk9n/X7W17Y7BIISJpFCxe6Cdfqq9RvxT0YpNtD6BDYYO
BTfuEXihUnnI67zWnT9U8riNjcaOM+DsmIgNEkYa4q1Ok18mzHA3INyqAep7vyZ/
eoLn5fLlj4zDJ0HujdtOI9qYAqB1TynWM9uLCcqFuQeeYSTzjnJ3YBn/HCTHewVH
HSVzvcX9tmWIYfssUmSMDhhvkRyDZpedkFTl12+1Y9t9EVtBZ6Ixto4Ujtwfgcu8
0cX0/oohH/TOCWU49av7bdRtT1ncIO2ykuRS2APEpcX9McRJz9mDN+QWV1GjEbS6
KmJPePqUtL/6SVKXZ6d0g7CI6H5mAAU7lyoEKu2ivndJw8sZIT9Ta7gA3g0K1ryE
BFdlR7YBAPP+CONIFcflsPPyDaXUwXYqY8Ot4+JYpZ7Sbsb/Cx93tMb1fWP+UqLj
3U5MIajASrrzTU7NJMdzRTftvOPpXYtci8FsfBpTKO/VRWn3s/dPEARpctWBMO1E
qq5Ps2PxNUuNAjSng1jkN9pDUMZUoAj5/smkh+VfHJZYBaXpgYz5Ei49qQdzNho6
d++LB+le2bLfpXOCwuLF0QFfZM7FSG6JIs6WBAUhYhfcmdYwGJzJ0b/yExd3Xb8z
ZQF773l8HkRBYTcPRC2P+MdkTUE6yB0Dk3Z0JTWItEpxVJi4A+q09CWsmvdrBvgF
KVbQsCt3Jkv5ziWW3yMs369HxAo7qzoLy5T6/IekerDYAHLCIp+f1O20oXSzeW7L
JVstluM7p+j5/Yxyi/9Tu7tbQrofpsN2jDii3dXpYKrvo8yxB007IvT/WNiNKvZm
U2A/1ZgV3HltBiogOgtBM0llo3gsjmfuUlFVK7BK4G8BXWUaVvIyROl09bGj8DBF
p/HEZb5wf+T+KdxzvZyHqD/X0/BsT/F4ga9CMU4PRMdH9g0nsMklHB0zakzpyzM0
knUg5barX1tbT6pR8RvsfueRfCnnP36EnGob1GEFpe+gthzng2wAt98skj4bmyiw
MBtLoo74Otn/FwXkY20i3YqU/e0gprQCtnU3W0UkrkCTYLi0sA6aOE5x6rdvOx10
UJuxRxXAlwcXjgOtnM2FPYlg7ODDWzv5Wp0WTTbNk1XKN+asTKUPpM4FJ3zZDmIP
F2x3YNMDcaSbFPxjfNVtsSufcLmVZD3LjYFXmYAXG1UR3cjiC9EdvSNNW4UemWsx
iminXMt5ywhfWek/+sNWCj4vVBVjt4Qf4YTcqQVDfX3Urfglsp28DlQx8RwaRD0p
wyfE8op07J1XdtPvboRDqgeuhbhDhVp6glMnBQaXcZ767dH/j3PTeHap/sjg1nG6
sXu4kMvaMJirHDUQZBRdacdLcZWt7/nzb+oZlcwq5EtZ+ycQmTxhp2xhGz8+7aB4
RX7DrDMkdJUKG4NBFl3b9obadgFL+p2SBgZxmwkA8/0wOlBcj/K5/5hOxvifwuyg
HbP2bGSjoa30+H1RUSpJT48jVSF0fabYMPqxtDZWwgfSzUNFlRIiWTslLn55n301
CTaxaFEox6eAqw3a7KhB11Wmuun8b5bxQM1L2L6AC0omcbBji4qxv4A/kyxMXrcB
mGbIBrE5E/bt7kFGFlM7/sq56Aw1eds49zhcQmKSBV7Ce9DzHxNgziFyJC8TmGZw
G4STqsjZTIdPILTkXZhf6wSYGQK14H0EmAlZ8YDJ8J2Nrx0r28b2y8uJbbOdIJs6
2XDcx2QDdOElDtuHlLWQ0s3mwQnYkINuJVQ9eDa/YqSKf6HSUFnhE60hkoYrV5+g
L/8K4LBwPVuYkdTSbLFqFy1e8j7WxI3DeBQxS8ZEYHWEs5G08KO4VfbtexLig6F4
zwprhvlAlKrzI60DMeZbt/JaQKAdo9+C77jxYZYjZw03IizMAUnEk9nb+WWd8QMI
62r2o1QR8qJmnkE0tVbXmteO3Jujd4b6CCWKnLXa1UtpnUf6s4uNBlJkDS0Ymy/n
92haE03LKQYacbDdI0h5j/F3bZA+sjK9Xux0a0EibE3wXED5wNBGSJDpd8hI3htW
x3NibOmAGjc/ypmgw6N+puG2yKKNoHGzcvtudp5MoLl0+S30VD+fbgEB6a+b7JuY
dmUL+QlyMTqGYe+oRuVD4bRTg+wm48rOga4noV+qt45fYwhgQxIhkLnXskMlOKo9
saS8ugrnVmlRZenbhYBUNr4yMpfWhNO1ygDdlUTqcFLHFYxXD47ePsKkTjh25l/A
6VMKPMkWA2zS/6ibe5dpPVeJIBtWBNT0ynPJrrKgKBh5j8XICS+71HIa16I7LJdN
nfLA6szbJTwA+EaEmG7KC+CzFiQRo5EELjnBAlhxteDsH2Zm/zeQbXN2Wt/j9lXX
V0Yj1Z2mP1GEvzfze+Oj1KKEEMrBIOxPh4rEwkG9eSyIcCuAQIxDgoww6M4HM9lE
CvQYghT5mX+kNAgQcW7ucweBmJd76C48D4w8rr9GiGceO+vGpKHK+hFKMa0Ty7Wt
sh1cblGUO6GB8twmT3KfEwK03YyDvF/RygjHzs1FLWvd6rCbYCg5uu2hIiR0zPic
kY5o9gHopNNXrRCcOw2LvxzNO01DZcVGHw1gOs5V/+IeWu93SThLbIi4VIRo18gu
cDqmJ8zZpjvBpKRNLxc2gFJC1WYbYEHM00r1AdaXncIMgheAorqNFdk/saJwjbOa
Pwj/K5h6/JszvnTun23pf62e3ZntMR+OLmmVKythidZaIy0KDsqYUjygmhb/55bF
YRDb4axdk6mVyYtHuVNDUwCq56aW0Vm1I0EKfZ+uK/8Sx/LSbwRHR+I2MgjelIU5
4Mr6SdWG0Fvby26T/S/4rgnqZTKwTwUNRpmYTaNdoNOK5ixbvF2CPf+h/iUDGUQo
7FjJVN6Vp9NsgAgGGL+Mk52dxJpA2DFKEUDFOQIkHKZ+eEsgLWpXeGGs95SGwrpI
HcK2PbAlL87fh1bthlgc81FOc4ive350ANPHwjNB99Wp2GtPTeT+uMvxUJm6v28O
APoAhMf4SxJlw3n7m+eO3PrYcV4Ag3Ugrr01oGz7bj0eEDbTnv1hkwbu9UyHE7Ki
LiHnJRgzFpLciuuee/rNXt6zCQrALxVNU7q/NHMVT7gvle8ZyK9YtLqB/r1V2Eod
nOGyKI09hgUoev4k2kZ6GyixMzR0d5C/kcDCgFfdrZIQ6mYG5ZT26l3wBKTFxR2u
UdmGnymifH6GtiuGSkZe6Dhojer1V17NiRrB7TadmV5OSvPvvLyc77AtPpDiUCIB
Q6ZKp5xpW1RuadXkKf2WPyvV6yuqBRV+M4npDBDIsL48uAX7ERqT4KcYpYKBy/h7
eItTEgvxiZlojqYV1gp/8PWpZh+8FzOdiKHP+dXrko3+7F4dxfFYyBAVFaVql66A
/SVOfTnNk7Hr/9W44ur9bl875fKer3JQjk6/puBxfOS/WfObxJYOSR4qr7NdY0aT
is2WHCq31f8YmI07EIRCASWprWCaALp6kblap1KfdNBmU067YVl+lo42XHsS+idY
wnJekW8NE1Wk2Al6qdI35P5l1OS8J7iveRXdknZy9EFNHT/3J4HJgawq/SuY661l
Zf8fWvZVIsQe3skegysx6dyplT98l3c7zJCPfyymXQYrQ9+2vAKIJaVccE8DSiXk
q2QXGUl6c2+r02euYggeylb4tFaTIacUtTtYVQM2UR2kzrp729331ZYZP9HjSZwX
yEQasY8bVcqBJy5dCxbccL1EXSgGDt/HkWrwYg/OyzjjQoOycW7u/lXTMwjOFMJ/
Kyvvw4NOUPUyt0rw7fvEF34yAJXT9OI2Cfd9f9FBGtGMKroWA3uZ5zWn8K882z9i
99Vps8iUr9m7Axx/FAZvFJZEkYbV18dnBjI/01lQrFpjbYO10N7QzckLAdIOUxs6
/+x6Z9VQZm4X3UlyQTq1wHsLil51st9YQn60UZV3vB66Mbc97wl+Jbui6rMz/KXR
REDfxn3NQDznAxf7qMxOpQDUzMaPioA/UxApZKCBywFIfcMdTAJE1F3fa7XIlNUo
rqpt+j+Fdl6elP6nnjGK04LfAhMiWZdx9pBaiht4yF26RWqyGmILgFGisNh7gebO
VFt9sICNW5Nz38E5wOPGnu0j5nvQbNUD9H+3Ice0kTyGJzGzW+hwibIqA9CzA4yR
CAAv2ny9hWkZZiaZdGQQ8bXam3RThRqqgRiRAXN+xgYCSpHw9v6Ex8tzNxW954nG
ZX3TZbK87nUEcDcrQGKdEsijLFRk9+STyIuSX5hfLo13VawVN18UN4/ZIFmAFFwh
k3kZh/xh2JOBdwbZz5RPF7uHm5D2ZMXNqhpG2ipdk3yJ0hPQGzRaMSBTmRQnhCJQ
Uzlb8yXL1hdi5Ca19tH8Xx/tY5s5GkuzLRVfb1IDaQsY1Udwb6M0MFYz3f1zLDMs
8BmIK00LRxOzgKvXpMIgOJql9iFx5jppdZ+D8PjxyPTqnMKNfeGCg3UQvwGgnPSE
I+X4FEgBpyCfMtncX5jhXpUkFClr/gh8477k3mSVaHAZsDjrHE5nBl58gnx8uUS9
4gA6D8q+Wmt26YdxZLs5ISgdKvwBlDjK0U82nHhykTVG6CRMlsNtvC1R/NHlV32N
X95Kqd78QtIlARwA4CYfosqFtsv/4bLAeEOqKJ9CFhNMCDMFbRQfeqWDB/xVi0qZ
p5heC70aJGDKIfWoFSG00Oh2aRa4M9B1UnOUl1ipaE5vpPs5J9sf6Ji4DPmkl283
K9VtKZs9tPZ9Gr1rxcuJ69Q2DqigsQgiUSxAOw3sburDoiw+ZVQsCcawJAUJIUOT
h3FM0Plli0VnkylKd7qplqdmJi41gmLhs8qpY12y9UDoXMdnv2bhGYV6tSbREmBu
478f7Dfq9Tdv5oHSB3/Awz6skTckKn3Tsl9XHxhqaLKgLhpXLsbhh+bMSLbnDmmK
ZzwOByk5S1VhG2uc1f6YhdIU3XrtdBAxtMlAVgur0AWokL28bp8AyjJP7llE55+J
tgQkoL/8v559wsR3l07RptcqyLkM46cQf+d/YPAUjYwPR3FA22MMLUAstQCrtq3+
CT+OGwAXMkFu1CboqMa86V29JjCJEgtW7upI3VDao3J7JmdzbQ85mAeeVv4fli7L
irtfD62gYQXX5UWl2QYDPaHXvVKuEH/0b2VCZxrRlxRNdusGvRO745SKWo3hCEEM
IEpnVQfaCSgoGGdMaDvWh/i+aa+BQLeAh7WiZhs7ZpllpgtAC14pAfmQymPNP58u
H0dHu3F3QFHcVzKlMGGMloB1VQrnFdvmVVh36yKe38nQqmi1yHPSCNeX9mv0BdG/
CFvRoQx80NflOFWHygJfUWkD1M03ojlMnN2wrIPAOzrYe5dv9KevkKs6lHRzqitr
LZwEi1RUS5WIuEzjyfVFIHsxiksgUEhLSxvdUTuld604plpct3IRzVT/CRv/9Z51
6Uf1vTCjJJrpybNHkG8KdsJb0syOqqzIH+AFLzrHG7lyj7Prs0z+Bjz77zMHmSPR
dSWPxTtYc7/FnKycbE01p+k0kP8NlAm1QlOdW37Blpl4dleO4rylwX2iOe7bbzGK
RgqJIzZLguBcoUYjtL/TOkwLAH4BaNU8vX/6BA/4yyooEyffwSBiHURqc0TNcIZM
sgmxeke6XmtbH8GPvFpZPgdSWaFTUDot5PJ6zDqKY+yf+DkQ8AVYlXH7ZfBUxyDa
n+0fTMKUaqfo7JOu8GcoZou2UlgIlnGdt2Joc4gqrFxtotkvpnEfDzYAmK2aBruE
9f6DoLoWEq9QqW0Pda9Y5AnRokP+X0zwia7DEjqW28e3h7Uw9TJwUgt9U6GkIFmM
ce+vhrTJ6VQYQtbdLr1qYDYR0BCZDkPHUBsmM85z/u3Wgzk4BY+BAP84hm4aeYK7
UGWCLUZg/vj4uHeW1sfgX7scLhu3AmPQmbIuD1N5fPgSID6VQpuNB1fRmhsFs1fP
/3uFVroPy1IztfwxBkyRvgKu9O+i27YTBU51aLEoW+wXkla9NRqyQceJS3chmene
lkdaKjP/uBwVS0N46pdR3ukFaX78174qul5Bcc1+oc8kZuK8b6WNhtXnlO2qFg9Z
C+JuzkwNEEdXhgk+NsLtByghwpTSVQFG80AKcxEY1fBNzWdNIjgRGnzln5f9m/8h
dPp0QJynk6XAx6Co5tgQZ2Bw6jdpT5xXY5CBQp1xUYi8qXsEoUFj+A6+/YUriFQA
as9SA6JaB/+X3vQFeDnF6CDKuSNIl5CVYNraSlMPt6daUAOT8/TiOqFoKcO8w/1S
6yC6vrr+Bz4/OLzxhdiW5/jNvXye8RNG5oSKoTIoKA3JmxBM82Dms87aZBXdDT8C
mZ5z4h052YodKiRpoNwdlnln6Kb3xKpnZuHVPlE4eOoIMBzBgnKPJh36kuehnBOc
6z8PuzQOF7HdS6HkajJ8wfwiHA7gLvPzPhV2ER7Uy77ayAeE4cegD5cTq0c/czwZ
50Cstwbur80jdKeDlKlzJTqimSFsykarV1g8vQ51kbDSndtHVz2mCj1GcuRRNKmB
RhAGnC3P55heMBkse1vhz8um3HT76BW7dS9xgx8NTXcNuk42WvxoGFHapBNbxC+p
y/YgbMwSLr6VfzQmHc6ScyKk8uzV9t2/+YKiSkbzj2D4DMP7WWeU73WhXx2B/Q9B
lyb3GLNCHOi9hNDkMoNy4yjZePy3eltv0x19XmaXfn1t3QtQdi/SxMISE7AZaCGW
r6PTXx9dVu3tFCAbHltXs7IlVl0pbZtgsy8WgwihVLZfTtiF+Wl5V5mmnUzziHSq
ZBXliULffkZqxtaTQKY9pl2Q+/mEHnv4C+8czSI1ow0aHtFwql+NNwy9zHP1A8JM
+7rz5sPRYE0dTQrmDKZ999UR6T+M+/ZCsM96IzB8PxiPDzayiwxcpBuFIIDZrPe1
WBjIt9ga6fOuhvYgRhdl8Eh7pu4s8uu+gh5Oe08pNzskxeC5Tph+dAdPfdFpdUek
N1X1YzVN7ks3CmkIfNSVy67GKDT/0uEjt7ZFEPUIRBbZ9kVzJgeiMfamhmGaOhrW
WczZNVBVj7abetBph7OUyDC+Cl3zaTHFvZLFc31Q2T0IkoG64kmxmoxcznWeYKqB
vHeMxuWm89SPqZexCDOt+TGSHxMUo5hhAaKyrn9MjmwhVQa4ZxapPJo8iDkGP05o
scGVGgS5ruNjiEtmDGNHqG4WvUvMUxuFFBaQEYOjRChcYiXNfo0rnozxgFrxg6a6
lxdWYNYshHZW6oCB4PMOs2w1to4gYZRhq1iLuU4WLl3abPVVg71aziB/dce7G5zw
F+P/Fij6yJekn6Fv9f6zbbhvupYHggwVcznI7ht/18QKUj9sXqZmUWPK9nOOZezA
vRP+KY3VxaxKef+VrPRYma3niXReveBa+lfKC0A7zwjsWqjuxXnmOXrsNnABlW5W
UYt2xN2BjEaKRXiE1TqeCEHB0JnEccANB/VG6X31C7+qxcuE9bd/fSHYlwsy6FOA
6WK093Ydg8U8wEecP2/IIYLp2K+i5fyh5/IAyJ//h4Pa/DozUIoIHDSEkhLjYQNC
ff0lOnuYzDzRcnVLD9IhoyCC8Lo215LFn3VJtCAbZz5y4vLFY77O0qBi8b163Vps
4twWvjwYtX4/xk9ajhqlsJebfV/fMmxUZJqrQ0+sWERt946tjDr53bkb6Zqf5tDO
++FTnJQQuZYfqDNOB/WOvcBWNJSxQqagKVeo/zp+sCH7G4hKPcnCwSwjSS0EYwQi
XDrCsH4X8KBIPWoNZM/s/sbBCGOwbKZaCriaQDqHo4b6Phu4cVWZK2UCKwbkZ5tK
yivZyYLuEU9x2GF87doH/z5Kb47YWgBPIdmbkc76jFLh9fo3ff1Cylvya6wVHO2k
5Mzs+7JoVdS8PN/XrfRv++Rzckj3Cewy8uZWhM4ArVd3zmYWqXCQwHD2jRMvuiJv
0ids9RmUIicSBeBiqIxSKI9q4VmtumDe5OV35FyMDvV6LmMyVUn8/hkRpenZ4tv7
KPi0JB5KJ3vdBjAoKwRry+osKjAL7nwI+MxWGa1NXd3LVa5eQlPqEweNa5VX7SnE
hUwx120eCvGGvjQUfa+pywmaxetPaDZYp1G0qUbQRR/0/h7Poee0u7tm4dFTc7gI
JEsKoAOXmsMbp07biFPRyy1hPrxr8n6XGr0GkT79IU7b5Ch/5I83YpIArO3ZDHez
m+ST7xDZu3X2ESkK63VukYypcYCrGk3BuAJzI3umycAIeKLOLCQdDDsTrP9wz8m1
nPhPJmh+D4DvB9k+alqnl8g/JLTiWBX8gVKpBn49RbjDN82Ke0iqOPfU5O0jv+PU
L5obgXoZi0X+zvqJbEPL7JhC0pMzm6ZupiodW/Ss+0ugF5qmDSb1T5/E4QBLwn74
p2+0n2NioFwk/O5aSA2doh4blzmNNG5QcdHQ+lWL/GeihPsizJ29nJm6GadIM+/d
IpxDVKsn0h2a2k5caNL0D59TZ0jEECj7lxXYfOwmmWaT/P+8NoGNIu5xwNqiC3nW
02QlHL6xmeiP1sLWZrvHHPtgQ629f/Sid4GEps9pTTeu84+vX2JNR1JKE4FKiToJ
NdhJ9JiWqfcEtKTcTfoOlPlnAMZYD8AzMMFpCLCFQtOrK+RBetD5g/qX+YFQEoUg
BY1rqZcZFd4jM8FrvtKjzF5EY0kNVuQ2ZP9lUeW50g8CoAPDiooAT2ysWcbIkixR
FFFaLe0+NbkOQGpNDguO4YERdO44/3qnJiI5i77fn1ckWwduWyLDXM3rGZSRKssa
guHZx37skGBQRkvc+wZr1CTAipOKDvRkYCP9iYOATcdri9WUUfkzsMhD8sRGguiT
vWEfxiF9HAkCtSc0MByTSR+2/lqxtrY9qr/KJHaIoOudlA5fmaIEK1hD03QC5BYG
E8yTjQhySLH+oV7iafA5G5rzcvFoLKEMUlxkH13O3+UA4KE3sjIByKsPBQcznzi4
y/JPilOLwZvkQ3V2Yyo2c8AmV2jeC8qcX6olKujSbbzu2GydFns+jwlTFmi/i0Xp
0bRozsKIMKdMc15NIpxFDRl+NS8f56+vE5d/5tzirLTSbCHTWtnzZ+O8al6r9xVo
Hoi1B6NY/GLbkKh1KPdKJlP7aCJliB/fjR913z6WiOM2Drpd4gdml/Y5rQ/u6JJQ
SSmFugKWaviUOr0QwFsdt9RTDX5IdwfNZT6c45JvrgiiYqvFI/xWM+lgX29nn/Ba
s0drgvpVaoqPxq7k4y7zA64O/sc5rSOSDslDQNm4q832u65zxSgn9sI08mQL2lde
CUy5/bcBCd4vZPq8L9AClEb3wu0j9ER50RG/it1gtiqJ1Gb3hoZHUwIbvJGiL0QD
rnnSKWUKkBbOG/EDWcs2icEKLwlWGjjAoJG89pWuDf5W2cKt+3Xq0wOxT7EQsSJR
wn42IjR/fKxntDg4uGDtE7H0UJbZooBLdo3GK19f3v7TqlkSmeX5qG5GlPwOb6Pb
uG5uKSKUdvHeXiKS/cciRG+gkM+EsgPbzryCAveyW3bdZjAeLtRY3xXKvnuNSYhK
P9FHoJ/wobRJ9+4VqIYDF5CLr4v+BMRoA+jyeDPuIp3+TSlNqY5vp3zgL2vWTxTN
WbF9S3++zrX4CS00RDLKS4QWjBVtMvoO1oiT8cE/Bar+NJA6GzCI6Q28oaxUzKLM
E0gKz8ftYOXYKKBvJCQnf/RABZogf0jMIvTjChMG6Y9/Lcnx7i08nyXVR6Zmh5+p
6wtVKzXtFibAqlR9gl21HwmgPK7bsX8eG+DmYmveMkQ5/kX1XHmd/kKpTpoWWGsS
bn7j1FOm8N3BT6p3O8kMRPjzKttYLccx9xgnMPpElzSdSZe7tBuCjLSzqOd4jQhX
xKTDokavAvZyysSNGt0Uz5ozaKgLLMnbXV5dYH4Fkq4Fpt01l12lr67DolusHHrR
pbGjsITovjqv+U5V6VSaJA1P0Hnz2wn0FqZr/IuHW5A8e6ZFugrIL4bO8Rumht05
odBwAI/Z2YIZoFY9kDbk/G0Q8BxFYB8xayKHyNy3DZzr0H4GITLHcWUX9bZbpMCp
2/geh0PwNmLB75k9sdjeGwL4WQI1BmE8ixPlE4xC8pDlHumDJEZ0wVqtuAH6C6lG
Ea0UVSSioT3ZHGwEMmbhFM2JNbiUmevlthX7UtglRshpspNJMEekqnsq8+sPWQQT
euJTgV2Qb9U7mmzsh5nq1Ve6JDnUAVc/ApBxU1yuvd6pPVW8TFWHUvzIPI/4hlyO
WiQr7gQ8YaSA5LQfW6ylPUn7WZ0ZJHwNeumbErsCsH0bxMAsdZf7rN0OFs4Paz7j
IVN8DK5A0UBiICe4gfyeOg+noR/De7D9PTWNlbZH3yD9KskFF/tlDMniH20Gp3g3
tQkGLstf3pGcpgR1kdg+jg18SaEn65Pv0l5zWYcQjxolTySbTfE2+yuCQX94cqT1
kwnQdwO+lBtKrl3TsLwFOvqRpWQjRvv3uBRMx+VHZsYGuTXqm/4a/ixo6uNyNsCl
CWALCEJXt9/IE0b1OuhKuco/FTVBoFsvpSa6X+vC+ENwie3vYoy4mr0Q1zUG07mU
thfvsIYRdVBqYGtnk6chmgoUFoQmlMGcdANlnhKiWDIv/RqXX9LZMrzjZ3Od1MLT
+K1xdzUJ9aIRjFWPt/xAI447n4TX6COf/xkMz/oTcvH78Y+0NNMyy45C8tkKWMKH
v5VJ6I1TEDSfaxZVN0NSZGmjklu3QXcHxjr1zL2goUgN8j2tDCzUP/x944oYBFP3
oT9/9ozm8VlRzz+uhUsnw6W5fIHP/aOrn0PNvwSJKqrTB72hhIFPEwY5RVpD+mvY
+obmqoAaZESUjXxuLk+qAMWF/UTgQT4QkSE7MA7XLIKaoMFRyg3PaAUQeJ8fz65F
S7zfldtC3dxq222glyHZnXYH4hFnnlrnHyaGyTQ5yWOI/vWbcByPbnKB3vapf9GO
L9wEzXnqPFB3RGOHTY/Bd4vvMIAJcgVBsBLfmc1yKdhVvbVNcV6BH+/WRIswt6w3
T5VgMxfwxv8NFd/lNiF8bE6Hf2YNhjxedFJtQc5ahC3YRszVYgmJuTPGWOlZ8enr
OPEYudHAO6AiWZ3dilJPi8dA6njYwKcKWANn3AUwQ8jnEhKsQ5CXNuqYZ0L61Pbr
oDQN8kuYUnin2mBS+677WZtlGVOab5cxml4nk6umyc1pOFXN9p1LAfPv8q8tIkvR
iuqM0K/8ZoQhISkgAGpbCkODeOg5Lkg3NIGWp/ISuax8ibhQKilzVlRnlNgHr3q3
FCUHlY2/vwkF9oyDGYfygwMMA7Y5pGJeaDqrhDg6T7UxTnLPWA0D02X0nw2NMaZP
8+WgjXdZHgMZAWyP4h53Kwu2cgYzDCKCnoj7+Nob+JYhZ1eKFY542o3H/me5xZca
NNZi5+1u3gsu0yLBjq9ASW8UqFtUbkHb6LN8rLdUHRzgyphSMrJwBPePpoSesMS8
a6pwLl28CblIsZEO7QRzJ/K4O82+Q3Ps4CNE2rOo8Mqbjum/xnJsfoaiAnz5/cHZ
HKYFzCzsTkV1Qve11Mc0QWOUJHcyMLJ5vJINLZQzWHsTa/9gMn3Gib5lcx8rq1Np
ndmpVzCErRrhMssgC9GRLc2f8ROgs5DEGO8+0h1HEBYiORjImHW8TBMgpRx7HqNy
G4cszLdfJp74IbfEuVW5962V4hG7qXio68JriU8VxnK5cYlUWT80pyT4h43Q2xBd
C0OJLmxCWsigZQjsZgruF/7chuPna9tysRV1svaS588i1loU3tqiq8+BjssLteT7
3dhsbqQeEXF0BZWJM6/vLriCYBY2sMeVgyiQ6yhrjhu356fdXTJKokDfTCQi3Pf7
OlhTY3AHHiKYxtnpZLtMhA9Ef1jYaN7w72GfNqVcpyJG5wbd0jeD+Ru+C5dcFd2b
ietV6I4B/5PlrCV5GFwl6ZzIXksSHWc/7ouS6hA0SxqG8FPYIofGvx4s28HU918x
VBkX9+b97G2lHB3HdF94tO24ESa8K0+YoEYkzoK/5zNeMpz0G1jIFECPBf7EWil1
lS4V6aQGg2H5NT8S0lvWldgRPNZUkPNtPQS053UTF/xxnOPVRzHT99xn55r7NM+X
tuGQNEgw0r06WaxWeXes4BQFq4v0esLPF61F7yIqUiXIkE/M7isXJuHJ/ZsiaVS1
sA7Hi00lbXZVrhPCGzh3kIWjhTjSzpIU4w97U1Y7NSlrr0NSzVY8FnXidQ0CoeKZ
WG0uGaQNGCn8I9AXW69oo0lvSQ8ZeWMF9EatDo5p2XjXZwGJBwMHUk+Uoqq15EDp
X3FZUM+AkKsl/KxkZu/cNhCv5SxNL6W2MI5DRqmfZUdJ13KrjRf4FFtH0wlYXMLT
8BkIZr58YnuBmBPtNm/dZr2ETCF+LNp11aEHPMSKnE2uxBRJgNRbyYivVrbCNZVX
mTl63D23rcNNmc7+0UcEA9ELOqPA9NIJXQqIU9rph+F/GrhdDB+B1TQ1xoAL/zkC
ULinHvRy6NfyU+UhuQZgFjG5cDxgAT+iZSKBv7zcJgtIZl9PgCCFtaA7nKm2E9xe
L0f8nexYuRWNEoLDxHmJ60kP5b29p93zxYC2GYJ93ArNf7jr0Z1mmApE7KWyavIM
yHKGH2rlapraDswK30o0AfIRR4I7oeyEl7C98ICY6SljAybcXv5xd4j4D5leYl8A
VxXAZnj9/EBRUOFJlxQ7cfgz/stxzJs1dx6+n56pJssCquGZlyeQlwCMcg3+hE+a
fPE9w5r7u5bXdYhCVp5sm+beUgDJbWHwlVPfHvZIh2RXJdIod3dBWbyJkDddNM49
W9i+QmL5ENU2QV0Nu/0spcCW+megp2DBrrtT5mF+yay9lu4B2D0/0z1ZYvkZIwZU
T8P+5tc/pAS1RLmmem+Gi5kBjAOwF8EGhXW17UL9w09bsbuZZas/Ds18Wivz8sEu
g1WjqAwEH0RW7ETthBNrQo9c3ftE0/BIL87F8/0YZvwfNvPEp6oOueDD4QjZ9Mtw
NAtMQIDX1+fAz5EIx8q+u+PpJJJtaGzKILYCoorBo4qFF1v3EP5fdQq9DI1uJV4Q
AIrGsV2b+vTZJlVeUE020E5YclSeSUPgYrGMzeQCIYKYMTqHRAI2e/Xtry6M+Afl
XyhPAGwPpQt0auzZkdG35ffjFEoBoRZxWbJy1jbctRwfXz/vd/Ijgvp5Q3SUkhkd
MkAmXjxQLDECqP1NR2hWRKY5J4+v+1hODNpftKb7HKdU38KimuOqEQqXBwjri79E
Kp9+D+//JVhUSKR/xoUDgqAPL0joV72CcC1fLridFT0mkwqQN+maUnK8mqR7SVsV
hbSDtNGT/j4bMXAegeHp0MBFYxYVNE9A517PUvJkXVydYSAAuFEHXXfwsv8PrWVz
sVPmSwT1noWuoKEQUgi/jdtdzzbHPZqRjkdxYToE76j2EbQJYuX1s8OwYseQiaAg
2t0ygPAvu5HCbHFjFDgkDWf8RTwbWgeHow7XqXhZ42YE+tpkYg+h0njeHUWkVI1y
A99bRPemiec4KOHQdg0M96p0lWYfie0sylr1y0x0akt7ewuEkg5Iis+vixI8e5EP
kX+5TstagD50Mpk8vUslTETA+jlxb0pnlj8mhoywk325+TnpJFHT0/ZepHDhs5Mt
a4k4G02ZukjPURQgF/XtwI77ZluWPP6o1n/Af76AL8NIsKFMsllYFE3f3E5PyP6c
OZrFvgF4jZDEt2iDKQGT9o5eTpBn+um5esmTJs2UUaOHXxs3FaB3gKRQWRPQwvTF
F39rnYsX4h+TyK1zwzZXWLfHJfZ8Iw2sCiY1LOKXZIO8Vf1jjsT0zIRKz1amyrRu
VqJBz9zsgruL/x9SN9K8K1zbNyiF3fXwquAHqK0w7m51qWK5pQ0ib9QSJedNw3MH
rhFGiv2eKsm0gp52doA2KgurBS4aWt8+2HZ04ZgxiXFwMM4SuK7DM7n4Ve8ygO0h
wwEvcSz14Swx2PCsI+bx86mPfX/EncH4yYSQQpoltg3DyhElBWBLg4qRsmbDpJI9
BCjplRijWt99xyE2xyW9axKpE/qZPiTzn1nQG9yGHVqgIjcGPmyk1igrkO2UZ4Es
O5pDCn4msOCHLzxDTlqOFI9fhrTiIktad7+gljCgq7T5sDWSV4DL+ksyXwQYhr5k
q7QPOGiGxST60km8dM43FzT0Y0BZICh9zwkIp8BpqTDpOCwKFPwLEhAGkANOw53E
YUWuFBjewYZ9YBOAC7lukxlN26A3WduclD/XpSkXpyHMXzAMPZJjPZkp2MIq1AuF
s0gWA6WpPAcssHy2I8iSy8udtrqwPD5mzfQnTo2Xnlk6amVq5Kl8dw/GOq6tCXAQ
3icKvDjuQy9yHaHR/T7vmoFkEnB+/Jv5WMpMjXAhn+vCuQYV4LOh9MBehH8dvrb9
wZnJ7lRitY2DSzGwmppqN2iXRsFj/tTSW/ASuZoxqmgsQ4ny2Q6OECIMMXK38oFR
/yb8TANgTzwk/T8+1w4Itnk62T/V3BoA/o7p9PkV9xBn/Jz+4Wt99bGhlJCn1m4q
MnhYtFBqPRk/1AWklocakbA90cpYOJw3fcK8rGoS42qWyLUgDg46oC6/Nu2Gn7td
u1Hb2TcJSAmyPfYreFNOzMjOVqyyuG7kXaxzA+OlDyTstDXeXd9s9fuonyl2oeU0
sIinkv0FgoQwRnwJ5MVea19AUFdvD61AkwTeXvrOZZ05w+72rmJeaY6AYsI9kEP0
bcij9Lh08+SfVtfIsu30u4hBjt6t+9srfkHjWQaOzl9pqJxc86KoNxLiZss4/xLW
BdKWoUJR1nuVsU33c/FTNynhqGjmIkugLUHaI/xCUby5llIUkezRVrhVA9rAy7sK
E9yL1eyFuVM/hBN6qBfbzMWkci2i0np/1EaWCQsHv64ulB110/unyfDB2KxXYUtU
dUzX0pFFEmKwFnKhCVwAJsfLr1xx808v2DUvJFS2WUvhAuVDqvKjeo/gXRfYeIn/
LcpeJcCi08dVLl0FwhAUbRG7uaVRgLDxgblIsyBrNxBVHrbA38BOin7yQggVGJKi
gNL8MnjOkwBSVIKNIKHHh3BzG9cWwwkSEGhIfJOzwix+cGlIBcJM1P3fL37cTQMH
ODN/265R8UvZjnEdbksICFJi31h/M2GQhz8/YCwHr4tpiaa/EBiS46h/czJUYfoy
+Oetw/VEPr9wmZK96XZf18FzJJiHLOZ2afefDVT4F6zB57/UuYUljn/9hAX9g/Xi
FwkH2NABxMVrJHDbBKN01fVBDlmcuiZoTBuQYd3KqGG3xnf4VqoEte0t1ydt8H4J
oKV22ZcY6rzd/7MYnalTMkT+aH7VTdJwiKULeRkRx24MQG/G+PHpQPNIi5xaNK3G
vIsNnsy2k57DCQ7fA0DYVoWGBMynng5+/CGu5rQkO0SUzwZu5JetePPo1AKTGArq
cH9CS1OynJbNNi1+rBtvNiRq95zVuLO/Nygy+a9mYDrK1aLG1TpTW30t7P5/dyYH
q3kP48nh+MYb4PWMQ6YJ5I3yOLFou0PURNI2qBJk9LnVt1XQRnw+oEJ8iABdS9K8
qybG8Y5XX9uuFhZ1wJZa7kgO6jtEqAaTy95paJjVQ4EYeWIkRt/RVXe+tcX/ik5q
bPZ1Nfe/EvWe/yizshEMi0kXdSkAY/uJu4zhr2EireiJ5kNhkyebsl/u9uu7NJxC
kuloW6BspqJMgIL5gyczfsDBuKdsxy0FVG3f+w+Ggu3cs25WZnF775XroLM/4pjf
nPOi8BixYIwgpLcZlDUq0XfaF0wkyHJbZFyco676xD/y4Q38eYGtEnCPXj8ROIbj
EiTaBEmYfCUYUGUElJqoXCtYWyGT3Dn//af515AJSfT5oICcYlvbugXj9nRSAX6Z
svz23SnOPDLr4mDdJ7o3qeRbDhP/GyLzRslJfDE3LDigu5xAqLAh19k0/Msy7YKI
/t7m21PwTnSSA9qgK+azOWBOS05alqN15u6WEmXVkVU+Y0QV15ulcAORWgOYWL1P
KBGmOIxs/GLkIcdx/0q38DQK2FJos5Vroji1di/HRxR42K6iSKcoEwIha3VX4AEX
maZR19i7MQZ3ZgkzWQCvI0/xocIBX+dnVWH2wJBH9M0Uv0Um17IiXnfbOUArGhyj
EPl2XkIyVgrGEkUmBDPHYUHtVQASCdfKC4L2vMPSq/zHqat0EP5ORSYhazstPPmH
Tz4bOBBmB8tXLo/kD+3GcoYW4rv36rc6LD27mi5FxQvJQV2Tgx8KPJ2NHPWvJTtS
wColixbEyeypdM5/ScU3tqHSci0goYj22b//x9gQY45kW4qpSIr3Jo23f86d3L5W
KIK6emelRXRHnymKcY7KmFYelBbQDDWEx0HC135ddBjVmjgdgLGdgl/Io9LNvsjb
og0spJp9MopiNhxBvD+YrsDPdmXvayKHGaA8xyDc9yU+S1yC+GJXDtigeVODvX94
EMMSflqCJYI1dmA19/3xAwm8Cwpar3teWNaUVJ9c/sC0MwsOdqaw7a0iN9+1z0X1
OvBefgC5jAuZ34ZNRNesGN4Pc7JcSb4crqPRRxRie4Sr9LSFZTvMhvafP7Ktwapi
HETrucGrUtwDnOYjIOAulnSIonsR+xTj5FgPtxodCqYOMWrnb4ktz+NZmvSFLr1u
NJnwxtDx/O21FjgTRSPV9lN908PHCTGpVPUFC+q7SMOvvTo+xoCShSPYpu3eQdWQ
OqYpwVpvFkbvMsPbahhE4ph9k7fftx9hFOJnz8uUSEbDYyya/AdLXOldQRQuDk/z
Mk5FJ92ga8eOsiYz8Oxh5kObj87tDa8OX6P3sHo3+zq/yA+qgs3UAHtCJBbY1+tG
uI0NJJtVH7bRa2utjCSdy+3i6si93C3nBr0CaSVcvwT1Kif4PtNz2HC/bB417j/F
td5ZIovqqZ3ulSJ2daSEOMhr8zqQHL+nNOasNzfyVanNt9zoq6VAgSyXGT6mU6tq
+9fUXreIy2iwzHsArx2tPu79DqeI9seKqErETMZnxoihpm6CMJQ52IkLa4ULMvwQ
ZRZQuOO3CsDsjJXZ68N/NoNSaybJZngz4/5PECOy0js+itZ9JD0ikH0BWHubrU+D
FukF+vVd5hMe+bwafisG61eQujvxJWk+ymCsBNPTWi1EIhjTBeXoL9v6vUMjb8uG
fJGCV5OrFXhgzd1ghc9BFF3G+Qs5KP57jaksRlmHXS0KpTMZGwvOk2rGQUxegBHn
fxJ+hbfjtiWmG79IfKr8rxTEienup20TH7enxhiIS9e3H6fcl9tvzqD0MWJTSB33
7Me9qm1zHzuYHR7y4QNdUys6PFozQPQF0Iw2tOCiLFhJpkUMUIaCetn7GlUZ3rDR
mv9DMiMmLUrb7kUNOYA7LcB3guG+VvOCHiWKxRfZ4QnvVE33D/EJybElPZ6CU021
W2ZU6RskNto0uFIcO6o3y9L+29CMtf7I3HtxIx14IQytmW0naC8aDak54i3fWpan
B6n/i27wfSd/g1qio5efPfXiuLn8jUyrNI6XTvWdyh4QJEMxoF1cjkt2gy5Z5kAh
qfyPlbolQ00KbTkNgHtn/Rk+Ife452g7fKBgGAa5DbTAcrcvGnbd1ydq9Af5VKNO
EOFEg2E42Wcorpy+SrkqJfth9vWavMzTjV6WvtreAPnucl4CHlI8sleVsXzO9Vwf
r7370+y3RIn+a2sYSPyO2AVZg+hw0H6I58KjAw1Tug8NIMu25Nssw2GnKmnT1fZ5
Tp5s7bBnla8gdvuXNTui4VOoOXHg+qrUnIp79JxWptJ6sV5kH896fWhY6Z8L7RPB
9PjFeIbsIsbPes6PTnA+2fN44JhZJbsvGRKyBioF9fhp0uHoOu5azGrCBZiF1HcO
Lngs3XypEaO8NnKpNqW78N3aD6f57Tr+Fm9XvQFivBdz08rAEDUM/p7YsMQZHUMd
Rl8RhtifPAFGPe57xC539OGsiDKZ3XoIbOa/Y1tn4o7qkhv5PibvzSIpuJBWcx+E
iloWnI4Kk2BNZE758JH9gEGv5NteOzP0QI4vwMUQ+gVsdEgffLXxGePp3LEZvKth
V6QKdsMtPvDnfr1jOJPkl/ulPRqvfLSlmLhfwjyzps8x/9tn4nDV2vQoCzSbaG4B
j6l8aayZz8XLC55EhJzkAn0QK75inQmzscBYN/yHFbEhI2cwA/RX4lhcavWYrGb5
7fFkN13fiFUnz+ncZ0ibeVs1JmhRTf1gFf6T50QOF5AKtuenZR5d0tRVYnl3DgbB
3bo65L4VRr5Qihknbm3FenIdPTjZfiNW/EN7kBG4bicwgN8lZvvJsz/ZQa2OxDpI
UOKh9pt+RqzpjeFzcngdv6Bsc3HhoYeoGZdBssmVXf59aK+FSsGmPfGePyeVSWrQ
Qn9NpfwCvoFdOD5JkZ46V5NAzyOMkS3tMeu63RKbjA8rxd/a9rgus00ksaqVzn/9
/hD1P3oVMWtCUtse0JPzhBRMSKc/TYTG7rO2B2g8nHFwZ5THBvVy/asiQof+hPjX
n4R6h0ApMBk/i5nDS6LDtZAmYxj8DGwKR3FkYriks8X9PJBI10uuZCuK20CAhvXP
8Cw8mQX3ykBok0eI36L9qYyBwsJEdMbgyyUMn5GAYJ9m2wzGbwpT8h/GFHHHKmLz
F/HVZITIEWvnPmW9EJHDOigpvvF0zqrMefN3CeXbUitbZW0KdyDop7+5TAtB4HnD
lxNLvUwpbtMFLARB/4lVxmhq3g7llz3s5HO8E0emjpF5/ZUg5rym4OoTLiB/rbiP
86M7JxejFdy5fkjrHSB+Fy8N2FYNqKKYnwaxnTu3h/+xe5wI1MkN119LhvWXzx23
AiqFLcOWDl9OxTRYriR8Zoeq/madL9pnG9XuCvEakHjT0Swoy6LVrbafsvTiEAlx
zNpfxKptKdaKcUbej4lCcDJtEAfr+rk0nsb70jxyuy0O5zNg9KRZgZZDJlP1NvBh
FA8LhDwk2IpFe1os7rq5Rii4TejqW8rVTtPFw8QCffRrbMLygBqVZYCUpfbdbk1l
KLlomOKMgYyYLm2yU3n+HQCbyfySSjfwbpkQhB9+0qVmNRKUqyPdC2+sullPoS6r
jArFyN7pbp7RupbnK6m/Whva0a4wmYHodODTZb+oCQt0IwYRrp/LNccjO3NihBl+
ecyMPIvr7fwjEMxUeX1MCj2KCW928PWzcaE8SrlbVc8ZcFqCUC6eeXYr/6HWuH4i
HJ+bLnyBnsTNFQFTIlWQiIqGEwPlP/zG8xO0a/jiQ8f8Jh/aAisTUzNoUlFMQJm3
+FoUsACowzXEHBA1XIluSsWS37G/T7D1wzTyuJWC+JaJ2gUMWxU/5PpsaSj9ijxj
dC9rSz4o9mRnSF6ZMvHhEhh3+D4mpEfL+VdrJ6BvIo7PJ4rIF/F5kDs23GCJ3f7v
NTWNFdQg1vxK/kIC0LgIMDUjzNVo/4Qzan/QTuh7+50pNY/OMISRrpyNfxvgW4CM
cPPnBKsZUOHQ3T+N8NY7KD0udgpUZ4HcYZgHmSzUE/baemTG5qh7ctfX9GOzO/wK
oGX9uJU4gyuonliinfPSr15UW0jM9NJo3O3TFHd+GrnbqsBMU85RGtCXkm2SeM4q
ZaD36o+Eluvw446vuf4AVMWW77/gheiafoDsLixHT/GGCf3Xv6vtoAOehcC4K50a
cjz9N5b1WlxgacMSIzclr2/I3e2QYhGx5WH0K9sY1UpLvChI/8o1qxSQobsLxyHV
k18j7M77a2JjP15K1nI3uLzBA162B8wXVxCy18kcvj1taQZtFG9sawMD/T/vUSP9
t5PKy8J9PR5wDMWvXHLNIbLla9ujXYsBtIaG3cq0xoqAt2FgXyqNB5E7MCciY5/I
rinBGfW7EckK32jT8K2KtVW+2dOBVOGy2ZUFaddwBhwtcNdFM7A48kRcIc5vHJzr
c/DNnDa7x8dgD5FvX7/mxrgQE+uR68tA+2cKrCkyircyGzcB7F9crUp+xzabwEDB
lmIiHmCqiZ8VRxj6KiLJL0SL7KHjpLWz94gAH3RUG+ZG3L1+ALaFusDDVaQKFfv0
2Pk+I+Xkz6IOCSzz7+R7Pgn7N/zPA201WIbSk2BMoVdRGlJbD1erxsXscFcvIyUz
Z2OsqZk4rVhZ1MSe3aEb2uOcepdA5yydxanWATFAEBE5ff0Jtdl2QIKT7lQEFZ5t
rOe+BRM/9EbPM5G0nAaReueqL0c1plrCJmSTZkQ3HWvnCs0Jv9OH/73i1dmcYnlg
8tmP2e9LXqiQ/UfTdKq7FCEFc6lVcqMRAGmKQMCyCsujV8KiK370yC8vUeO6d4fs
3bIv36oLzLY2gyuStKpamkO+0Rv897VKxe+1aqEpy/Cyb/uQ94HNDbFah0t6Nnu2
VkLMFBokFdsgFGBiHnYAz7a/jIbiINNJxnmK42SagwT2oz9VJFnlLZhbHi3pQscY
NQVHTX+rx06lQ+rCprQQ8pixQ+THACuDsw4DAvc2dx94WnS7fPuYRdXmZCjG3JY9
Uvz5hf+vN4VXc3KNWU3aAkqV/xm8L4BryckBr6UhpwrwLGO3X/FDJT4Aujs8qfF2
67pyI6cnxgeC9XqXwCnFVf+1qjcmeogrZp6KD/CTydE12DuNCXV6xnQ4/s5oAVOC
AG+sN9fW497WJ4ohlVqJdbIpyuaVwaBktPIaCPspV/RNJVpWhH0uwF5U63Obgl7D
mic5zRuT7iCF+9wM39xjU9Kzc8BKaAnkg46gAeAcSmcCg03HdccK7vo1vS//imUk
lLr54ZaqqbRDygDjvIzVoLsOEAUwZrGrkQepTz6tdZxdgtXq9qJvLcYnp8uM8DBf
SyWuqcJbup495swSi1uf9CBbKDmKd4GZoaigsdD8A5QJP7KqEC817zhJucielMDp
sTYXpALeUSNTNOTc24LIUYfXr+9qt+Nw7Gk+KEDQHUUswuZ62Wh2IyIoaQQu1mT0
GSRc929CXERTg29Q0XUuJXbYDdibg3fOLeIFyrTwG66TRXjdN5P1qn8Q5f2YMT+y
iODRLVe7vIdCPaSyJUVrVg69oRbeeMvPB3avb/68pYIVnLhV+scS1E9GNvctCOmA
syFKAdk0b0tMf/O76/OD2TBppuul+i98zwpx3WLeW4IleTSd77BMEDDKvWUNHx6z
HdU96KrwyZgRS4aeU98E7Gy/dXSwABVG0A0sAUe+uA8lrSyD9INkpofoOfpMsK01
Ak5JqfkMHRAinVY2I2ST+6Bc+CsCwqDKP5wOxb438g89n1MzGgyDPNBy4SCTQznm
3JkCtGuxcS6+pKRKZZY0AOfkb6BWe4p4xJdrhRsOOu9SUABfkeXz4Q0yJZpmQiA5
w6KYl4GZUKhcyBIL0KoR/P7GEfNg4x74BK4cALWKniNOiRV0h8Ddljkkx+e6SPE+
Z8rgrcAcfShSxp9bQ6xZpnWU6N5D5MinZnOYF5gCm/tZx4Y/410VQnAGj+fBscs1
Vj6cMURL5c465/BvOPZ+aupiynB8iskEuDmmiqQyKt+rSIIR3buwlH3CriTrUTC3
5JR5oZj23kf75WiGI4i8N9oBsvh1pgIAyxBe+gGM88O5nzQEXPcTcaBCLQHzBRAI
ksWuV5SE5zqA22Vt2SaS84ZHcD1FCqvKW6rDcme+Tu1omfSV8BACs80SAQ5qQNK8
xkZ8m8m/OH6ZfLXAQcT0CIsDNFxHf8P7Jxm9pjyiFk/nz9eJ/LSXkIMXqF1ooaL7
WPimtFUiKqAreBerRLPxfHcihbTT3Vf8Bd5gu5TEz9XhldPoywX+Nn3DddoYn8RW
ljvgMWljy5JFpzKtJgqn4PwhlPFeLsMpw3GFE+bPE19TRybUqtTNAV2uPAU14Thm
jGHwIQWOQ77ALI8J+l5HxHXX5FKGzDsGwiUoi5ZFhHg5mZy/eTA+PtW4ytczVp4+
YfU2cIFuctmMHQEpR6yjvOC6zzeU/YYJyaf/zfR+LZ8etHP62Ni7SNkv2ksxlOew
XraJdta9EOGqQhqoA6tWpFm5dntrH0aLI1GPzMF7mBFjBR/Bx5REPQgjud11OaKP
zEbZ1lFNt2xHWW/5xQDZZX8i3FLwG+vLu5RNtGvKJX95JQFXMpcRK78Ix3zdpwdj
rVhdYEw5tzFFsIn6ayPc1r0lkkCL1cUj0D0iEEj9TxVSRSmSBWnNfkogNzVRbPtu
F+01i6BwCaafdOqhpMsIh8dd/TIngLJB3uAdECttPx7P+i2k/4dRvVGiRM/Q3lzC
6yHfH7DsE0Mj1QWMeinACnWNgmfmqJm6MNVB3NhCPQQBmGkupqHmWAk61/RQ6OqD
Zh4PDZLaa8gzwsQu0p/T6Yvo3syGa7068Jfn1Z3Rxls1LfmT0DAKLQDNPC462NNa
icfklgEwP2N5yoix2Mk7J5HrrXuTFQX6qEKdq1Bod/dKb7wz5QJwEV3ulPqxnwiN
0a6tN41m4iFNDpWymi4n5gVOeECFTGMkD+GH1qJ6xEfR/y5GWEDk/9QPNzt7+0v2
xwvm5wPZ3f17KHroBrZIkhCtlf0RJNPOIm8LZCIGTCMw4EF5WvF4/QPdd/hmXtUX
3bWK6T7xTLLwCzYOgO/HcxguXPhut2VLnQkh98LOb7sQC64nqFkJvKSdLPtJzOrM
OoWI7zCAXwHzaLMWn6Rw426Rn8OA/iBwMx9JVpBBW2efgzXPl6uU3JwiYDtfKNy8
L5+5++cQRgxQXrO7NwtSK5XCcB0rHRS/FSeLJoG/GUKTH1qNHO1Gxo1lgOMfaecq
A6XfZmKlDL4NkBtbq7Kh1qfeg0nS7EiB582WTBMzcZCdCzNp+HSXZ3ZA3c6lEEjP
d/m78NF9TF1BykStKwm3XP2QN3bI1PeAa0n0kBq4vn6FF2oBxEjPfk7Xx/XfELpD
kZUgDdBTWep1doszKa6RvxKan3XyTxj/8Rn6bpY3+m8n+UIlivGDcKM2q1yWJFl6
Rgx0rhUN+K/9vz9VTzK5eqleH/qFwWcK9YOnruXL/DPIjH5p44DQYZq8LAzPHa+m
lAM4w9on/Y1rK3yuT3/IauNjW5ebXgAOjLEEHblDdtljHas3EekLC/oMrWyVIr+A
YqhXVflBx/CPFfSljWSThCMvGwhjFxlZROuOjkpNB1S9TStGUdLbmg6/bIT3grRH
GcH2vjCuyIAslqEeL9mH3BSNcwauT9WMbZNorHn7ZBgY0T/hkHLputj5dygeHU6a
tT4eiS2p7+ARgQmKYSBrREQtChH/nyRPkjCyWWD7NR5dw2tLFAgkeziqvlKrk3Sp
aknI1I6l4eC5whlj8fb33wnSbwv3WbxjrO3z0FTNmdnAzWE1OaWfDF6/jz5MG5Og
ymmkNU0S65aXfXVevC5eQEghjFfoF3pcTi4mSO/OLM56FN4ylFOpnGyWnWWJCE58
eqldzi6p9zeKIg863EMrY6F8Hw6ZwiB/XOt73Kwj/S0FLtTjAmwi4jKSfSiERCWb
sO3wr7ty4kQOISPY9F3bhRmY22xjtQdN74dENRp+Zn0Pas95LPMUP4Nl0K5hAKmP
bGRR7+fXq+j/VVLEJbOH+Y5s15Vfz0PIQCBoTvF9Ao9kq+wIhmO1mmKl5zXm3Xss
YDP8RLyVYnFfY7jZ3aubHN8OFLwOhQFF+At+DZjGtmrvWazcRdDgW/4c2SMT9/oo
Jp1ssdq+bqmfieaN1DBHPDkLRPEhcwkxVZPivKlfPNl5/6Uq87RrmOfkZoF3moFd
piiLRkug5ixmqngAdk6E3ZNEsHDqTqLTx8WpDpdKDse6Scw+O2NRAWICBJ7X+3W8
o8QHhaQGmXvEj9vrbz64Hnq9A6k5T1RQVF8AUR/Lcx+uHdHOiabN/rAM9SdrAM5y
EL1/R4XQK4eIcZkUkdMXEcFrxhAKZ2zFsgJEu50o7s+1E3rBrNndMUCsPXykifBv
9wjjzut4mlhBLC1ZwLqynIjXPAm5/VMSq5ZhYq0qf+6TBd5YnUYwo9TgoKYiUmYg
bfMdVppmZMvaGtaAZbbjWQBhNnDbzKzyn0P5cXtdX2KbjPeuUNx46FCq4KFPeyfr
m5EorXOeZs+ZhrwQ5fX/YieMHKeOnLLXIuV+3v99LD5hdcsktfb5HmbpsEZV6Rcz
KYn9tE/onmZ7Zt2rPULAZbnSQKebQ3HPy6JXjoV6CuLvGJa618aPztSf8HoA26WP
Vg3u/DG0QKlI6i3LKyhDXKtdKYjQpLMEkEZvBbcBINTSIgzSq23BzQMSD8w9T6xr
sF/uKnGduC4OrqueHAeyv+Z1057YgDJZ/u7qZ9aDWQPR9Lhypgp9f5DRexauzqEB
sQh0zfrHVi9FM5CKL6TH8ytFFhOaOSx5+s29mz6+eSOo2ujqkfUuqe+OhVREhE5n
Tmh7PPbbwmqECzaqTaph+jrKSoma+bHZRTQggrdcvkTWQvK2J1X1M6uLZ8DBecaf
q4Xi88QGUcrCgMtmbpkiaXY28DWYFRTCyUhMemWyPjcOgY4bP6dR5qcOejmh/UIg
XMGzgacnfbIh/yLyYzkvDx7t5diAmfFoqh5ZSckijnWOT4dUgZYTYO7S+7ZwT9Ec
vZX9rmf2OTe9Y4w5H6IZkiUCjwA75JC5xQfFz3WBKPnOPz8cDdj9URmVgRg0wo75
yiXfvmw4rg6uHH7TN+Sna24hUUIsaXeoEg2UOmRcstLdBuSBJr4yau7C1WqX6YBP
CKhBqSfoRi3qhGRiv3LD4ou5b2YJIVddflcqXW+S+X6LPKv9LeE2aXY9q4MK07ri
oZbqMJyeaoMlqy3rIxGttdRxeSg5QkKxLX+77504sv2jy4Arl1jbN+1MzByxlBCk
Be/i5XH7aouzGDl+Z8qc5Vu4huiOWJOrSOtHbL3zR8iUiCVrDn2LfEQXdAJ1a4vS
u/xqhbbhkWjacCQqRGgbbkiTFwfZRrIzKpXgp8RxfaqoicwAjHEZfh9Zq/Vml2Yp
YaodH7exQMbzbTFmJUUkOoeSWJgRwPwXclYwIe5vRU7nWEXcyvU2akWTJyAuz3dS
JkJJ6JWiC99kGtQWYfp3usmBCdjSeUcf5Kxekw1Ol1r3v2+lbK1jfgewLDeEwcr3
3vmo48p1QPKuBPbie1UDjAELeMxBzH+4MWpNze6peGOICzSrcr17SS+XO8/ej+29
CZNVqBPI5yat9enUp3m97xLuNLUvtfrWGAKKhg4sPhnmkhHHD6AbsCuSbZDUqHAb
B+V4WJjG3oK8Klnyz+htZz+wshKim5QtFnp9wBYqGwj+Cj0yPrJeLphIeaTdXiNH
rUhnswOyy8mjFAky8i00F++YDCxa8HnyKI4zFpYYBTD07fD5yN1LOCFsIoa5Knb0
DChoUY4mJiK7Xij5oh97hv0/tMCp1U3TKR/hsA+AtLEloDUrzxpTDqPabQr543/j
kyaZlELJb6OJBsDvpkRrSKadxUdd+DbEwGh/ny5ll51AD9IzBWpqTI8W0j6L73MF
4eC4goHBWUZ8gPjW76m5VNqGWvm9zJHq0y4fUikw4f/XjvY8TQ244JE+Qjq9dax0
eJ0OD3M+uj7mxShvEUpYLmD5yp41DRpfKxKEUXu9nN1IJ01nqXIIJC+s7Jf2o3Eq
VOjSCKeIUqgbYn6x0PyH01qwQ3ONE3zbRvhh43dm2Uh/pmDb8LM9GCnGHR/KpX1i
nkLRaMseMEcyW306FwO1lHQB4L4m+DbwNzcPzHrNO18iUO0SmKcuaRJqxk/eF/DD
WehDH/Zd+Xpju+Fx9zP+RyBvd5UDMe9jUw9U2fLiEkgK934iIdqIkn7PsMjOJeFH
ao5BC+5SUHLkO26nOAVGkPgxSTNQAdWRLod2ksALHZEhqSr9IDccQvWIDJILEdmK
iy3ULSWRPUmieZUOp67lN/jXHsdLTvxsnzxj30piDFXFaS9lK5VswDZi+EfBlhzo
04/CIdG+Nj4Rom6rfny97OSeEAiaWv7D0/+6lVtVUXBecb3jvHp25W97j5SeC0JY
1QLb/dVMsuK1h0fHAph6EIUE77fB3si01pF/EwsmOD4Gpep+XNGiadITZPGHstnt
C65NwnFkvlIJ2n+13Y2CfuE7NKT9Pclv82rrFXrOlv2rPaHDtEjCZHYnZfe8B81n
uoWmH+hacBzDCUsCz36KxQ0i2YDg5cw1C1EXYPjBwXM9A1bg76QBvqZlN7e7ywg2
Xl/hXCRtLtz6vmdXQIAEQeJyNpwsu8iXQKunL55i24xwfkKhJ08dmEigZbINEzhi
BKlJQm6PUEbRUW+eU1kOCkIWYIyyGeHt8DBSpDqcRnuVM852DZ5oFDOB3F9FxjBS
QPpl/hbPIzS4XV+r6rpcnLPvsxNejOaMHv/s5nuSL5Du82Ym3qzcCo40V+g5KJII
m0O5CshFrfb/+3T+SAozuLpGtyJg/BGVfnrTXxn1ahkFfcaOCcHFkAnnRcZfJFLT
kCJ0m42Q7k+CePZmi+VtZSaKZy2KADc2exeWn2b7Q3ZtlFsex+Wruudmo03y9LHs
z0F1aNM0wgB1OMOVbhwdfkRChG112eJ3FLj8q0gnWsbNia8MqWiFIGXfbgqOycLk
2ndFBo25ckf4fVy/ahkSqzth9CbwxhSn4/4xuhv/rZjc1TsDAYzHz418ckgM5s2K
pMOCGXeUjdXliGBdgJjMpDAPdGg03gUSgbWq2Rv/Qoq7n0qoSlmPzHTqk8Xb5Z2Z
QtDcTxjDr1LNY+qxBEsiePfVQoD7rErenK6CWF8GcC6YloD2OiNjhBR17VWqISRQ
izIDaEzz+eyvltT+po6r5oX5rGA772hMOjzPQNci4bbsJjJPltPeH9Lu/dCmWBNy
4WUH2l4M9weFWOS+mk8kbvGtU2f2exGLyVWxh1N0CSmaspp4scyXT4l30W4Bpy73
NgqbemSQOmQMid6gss+sYsCx1RQ/03HCIhiVLV4GhIs1wSlP5jeAfIO8tlZqAmEF
it8gUJJD+9sEpmeCa9n/R0BcYiP9ICQEjt8Njv5UfjCFKH6yZ/2VuWxjbvceG7NN
nLz6Ef+z/Kk9ZSRHYrP4/m/K3kBPLEEjga9U+qGT9gn7/BMZWkKc5OYJT+0hkvU0
UsXzbT8PBDTy6EbNW1mjxID9DuGiw9AnwgVEJjyycJE0rRsv5E/zMcHIDj0Enrsc
cwIpgvbHbtpWE7Cy8pZsp50pW3wnQU5g0KTdsaOGeIepWyt8w02ZOG2U5IhSetjl
8FeHqKUCuC7Ngp3QEt2PZh9PWCCVcXOzX3j5RCjVgkeNAaWM+Ku6riJe53gK32vJ
yb+9y9eQSVo9G6MNcYaIBsqdYY6iOdoLr0mtgaiYVREZWHzddhTMW/QXc25jqRod
Dxb9k/aj+ohGTbqf9FXDKHgqdVMGrUlnl3diBfoC1DqBlynTnH1FuPJEwZFMx+Y1
ZkCMNEhKZqLXnF1UGJRLElrg2y05X4htpc8Pt5dJa+j8E8MJAYwPwUfPqHTiqJlz
RPZR+6WYV8/RqfoNS9X+dhT5z3uul505U3e3Fs04LB3Yc6BZ0P0tTS8OvlYI5UoA
dJ77JfM5qfiCyjiEvPjcXa4Qn6fh8lQwNC3+kdL9sdrjyiPVdOEowiHMVbuqFb/S
ODsB1fFCa0CHDaHkeX0g26gBQgpaFzM78Vcg/CkHrxDueoORpNkYrdf9BaUpfkXU
tSrxZdrg25ZQz3mNOoif7aG+HfXDg2aO2e0EpQes5bFGZWGfGmiLX8cHVGQSpeSo
B50XYqMVma4hOxulZLwUOGb4irzCHZvJaSzHRijMVI6ieyO9o0symZwHnFzOMhiM
kyiwdMNCfCbpaP0szN3UrPh9v+doxGLp0RH2tnsVQR3aBQQoRLAjdmIAfgGgXHfB
7iw1dfWIrnNkvewxiOb+6hvZz8ivbOXQSRfRxyoBoUVjnf1cgI7/JI5g+zpUdS6O
UxlDRRHlukuOGIGcbiJCcsU47H67avHXD1HNccz/7F9Jy0gBF6RlgeOxcAXnfCuW
Wo+XhmDg4if1wKOcHyq/lRvWeyqnymAtaDC9ypCjZQMHQxh0Ehp5OQZS/zXHaqdZ
zKX02CtBMWFIllcOwl8CVVUS2fFMHg0gm+e1FlrSATchiPip5ci7yw+x6bVK6tz5
Foe3BNILoMYCsgxiXfHCWq8NCsrQZWuMUbojfpIhfz33CT+xqweDtkyTz+U8izAs
hUT7Yt3CBzL8zoDoQHq1w1GzZLb0LydcafdzAnBKXDculb3ovVH6CiEisZjQRNa3
gtOmW1uxFAAEo5Qb+5GQL86Z3fMDAmG1x7SZmiUaCedLgTH8UYUVhKu2xDoxakjm
Mr//k9eaSzzKAZmOXYi0Cw2MFPP4j0O8kp01xV648eTxVMcBVTc4BPb42eT+RDqR
bNjxDg/OwFycItTiwskXjPC+MffWNDJ4yLx9eNKgNty8hc8plUL5Grw+NPrJexqe
NZXqlebiBqHvHxNecNKg6HpxOBWaDWL5xTyZyHvbniWZKqhDLTy6Z61LKWRQsj3H
BKlw1+hlU6DxZtXiUJclulu7pFpISKxTpA8ouLseEDEQxZwwPXM6yjDYJd7VUflO
ty9X8+L1uS/q2qAIycOor592BEXC4JqAbbNZaxhGjOD+GS94zhfJdyIF4+0s0z4a
dErurvB5CXUeqL4T9TGqe2xGZ4yJFF2J15KLHuaTezxMLpK9iZbzCo5cgwOC7qnu
EgEGvHxwygXRJjIvYfSVNqlAeTKtvsuzjybDYZFavN20XR58of69Kq/pDRrods1O
n97rkRaN+l0BiyY5zT3346wjKYZLvzSl3UU/kph3OO+riXb143LuXHhQ1D/xNDrf
ffnkS9nNZS4LHxHvemYN+gwrvgbzmln/8Q8xW2gX9WRKg9H4cU10cTptgYuaYBZn
daqzBUmeAOEbna7HQpeeHlSEWjKIBoOirB8ZWfsM2fjOhrYEI+day7cTPu8uRkP4
Z8egbuTnB/LVyN4sp6jrs0sfulTU8iPfXrMlnYSrYaWO0Tgcc2OtEZxkUeWOJVVC
K3rdmnDSPChJXnrZo8iIzy8LNgvUqUONDixswiJ9FL62VhnQNV+4bpEZczK46NEl
MPgte73UYxRFRabVuV87xNkyIuyrCk2SwNb36Gg2WEH0V/21zeERhDw05cEL34Ys
s+q8NOlh1xe3vITI+Hmt30yR+x0A7XjGcrUR/SFTE6wSc0WnaZUhNzUN67mvZr9m
egb3zWRGZiAfxkbRRWQJ3kZOPGZoivR3qSMWS5EinQI9JEEdF8115U6bkNmo8xEs
O963IYzWgvvwIiKjm2h9ktDkXRxlFg7lLkSjMHcD0SCNJbPhp+cnViJLqkiIqOUx
mC+Nu+DOGDxa0HlAD5L8+4n3ycYbHZ5hnYOy0SsyPlGE4D2pm7BBqyUuSdZLOoln
t7NoUSe9XN7pqrGlpBen4eJx5BJio5xz517J9Kd0DX+JeLpqigDvrhb+cwmZO9BG
ec6sX1Mv1OeITYXyPVK9fh3G9+q2/hSUPHtyHYrcihVWBaqaZN3adKycDvCjPpK+
JtIEKfsjLS7QXaOS5pKEA97PzAv9B7LvDMVgkR5/gYDD0MOJ1enzq8EzawtaZzPv
TwQDXPCMbJkBDXN/fhwJJwYfIothpU1c15IFFs1RHwCmSqPyqMRjKu1za0rpYh/A
Ksep7RfreXb233TND/boM+RjEXLaDMl6m9HiEQtjRDtIsGsR5usnOcyB8HoMv5DI
RMaMP5o1O3FKi39/6lXSr2A5s7QHg0Xu42J8OymojSesahLRZ3kLnARXZE3vX1Bb
8NHVI1nNkFYSc3UIiBRaUaStngYrgGjZqwkaiOhaz7HjQmUYPONhJpi44UYBM8wR
wJtCi/LRAzji0NuyawQ3e6svyvitj/UEGjV7Zc8ONR9eYub2O4KWTkw8wBH9+2zR
Ug1Up1oiKCihnYmzum5MCb2WC4CT7JSuRBn4et2rY0+t/6EezMwfMwT3jG+CPDW7
S3R50twxzCzKowPvugXKqa/rfCg56RwP6HwfF/R/SWpxASL08TkXNmpvV0RwGorH
bhz5AwDPmX7RcHZrvlTVseY2H0GN6JB6j8p0t5RKpCxsU2erqYmRj5LdT6J2naGK
xlHn8xZG2gX/zlYZYDSK9kr3Ir63VtRrmVzW2vBMPRfVsclhmHyr9WJZePsyVstu
2MhpHs+OnrFP58C/KMGOVe0BRq6pWkX06hbZGLqdF4b2zjt2gKVBpA+4f7Iiq/ME
euSu8dLlbC1jGwCRqncK1rElbEsznlJCqdW1n+xFT55D1gOFgPWGUOGLE411iXlH
bPjv3pcuT1VQbbdXUgfO7Uq1SqPZZNSZwORjczHX3XAGuLpEWjB72tStDCGGYbJl
K3/FUE5DPLYL9aEp6UUzi61J4wY1SyA02sdrbAr2P0XMemCBpinkP6ks/Zyjl/Yz
XSVf7DZinuviKpmZ5T2Bv4NjYbaKiWCS14144DlEH0ehwjXcEvb/fUk1xDSIkW52
xUxMXf4/BlwO5ermqtF9U68ZJ9M/hIoeEO/q82Rq/EqeHVMPAHrzZWOCXLLqCHHi
NCKcd9R9e7deydM67wmaQOIy1KM9ybAKcKRwK1lcIt6tM2e/Oj6YyDfX4af2wMgn
+ACSNm2eEiV7lNQFpQqOh5b97aSSQsmiBBaYCTLQAW+/0nkhzHZnt5VeZ331A8bW
y0tCSeX2AQsM67rI5EHqWkm34AjvISYL7L9sO6YzlxEc/yNvIlIYp/C7Cmn8XxTw
YPG5wZXxp89wrc5kI8Rv/OwtU6DbD2lHeqH+i1P70bIuWkGjp0EsPTrKC10sHeRk
pafBZOWRRMPtfZKvbIWlumV5ufwaT5Gr5ID01A1jfGc7HApcGtRNU+AyedQXaeya
QPDA76kWsshySOam0Xp5UnGfC1k+832OyhpaGzxrPWNtDybJTUM/v5jdSsSgOngI
j/cEBbRkrCp02T2KauZ3/lKnfkNX+6mTWVyW5PVpKuKr1LP3L7/PH9tqUAkn6epy
dmdnHcS9j37zPI8AMzZ/P2kl7JsrSd8D5iSLw9O070UkrVi8h63n8IIzu2etEyYc
aMp7S5PbIy9zpQxVQVmDjRpwagqn57GZ2EBNFFAZQH9EutKwMfSwpVl9scSXmQTf
Q45dbQ//KbhgfaHdH8KrOBLPucdEJoAgf+AijQhPIKXNbL39jmobMbAmCHp+tr7v
5UbkVu4ZK8dxGY8wGoLTno+AfsZzfBHm/9EWKrJ8zl9nUc4NFKwfSOTSmcZxl8rC
m2q5/XiszgVK9BqWsbhJUhzJCyrPTA+IV36ErfBdigGWb9p1iLDNJBzEwS1MsjgD
m5NUQqfaH4sIMmmQlMcYiMy2wRXeD3LJPW4jgGh8DAZrko+KlOhEbJrnxtieOvvU
0ZoY8XFISUmkk2eQskKgKQMAUw3bCOcqSFX6+ZsNic1QckrHL124QFxX1dPFI3Hu
CPfxJ6QibabGXYI3qeahFZ+SaweEOsXrIrAqF2sEvIt7qui3L6sH7w3ocIrmpeL8
PzgPZB5AajmbqawCqzqE9zsDVfN4lAW0ZKTCcd5K7gp3ukG+BD0l5XBoxiy8HNuS
/iSkugUFxU8PTKBpSP8s+Ql1iz1c7yh7sl/btVCQwl7Y2fkR7op77z7n/cKTO2VK
qfEwhZ3YE5yPZvIgXPFByzqzaSseEAcZtGTsaODrWNBfU+930oZ7kEG8dYBRPizT
IeGYNZFJYGyjb3eC6B7s4inVZKJUy5s26Wa3HGdIGVFO0Dqe6uh6K75Bfdw6kWyn
HPm4FYT+UbmuyE2VgKFJH1UV6z5ljbn4hPG7rS4Z7YJ3EyQh8nDlhijx+x7w8RLP
7uI45y/uUSqLV5bml8R4kCgUukWPeSDRZE4NkSDwwz+wmzALgKbHh9XR2BYnYTvH
1lDNz4ka1nYOwlhEhbLqIyt4jc3A2sPQNUKlKcq9XvPmn8Q4jhSv0GWROSKSad+2
rU5oEzjM8x3XtM/785jhhMPmYA7UogpCgDl2pzjaXUtRrWcbjelnHkhxlg515FJA
7vbOn+wRfhb3HdOrutD59OKlC1PxCjulrFfdpsiohVMkJTQ3fOMKqlwPjyQzheLW
9Apu0WBk2hY54Y2wtnr5hSHbww98APlpXOQsxx9pKGGj7bnr5uV/xljJtFHCMRYF
eWALHV+j1XfXV16DgW15xku1pkoMKeOzgNgolQVu6B7wnIdRuBVsVCILGfJciSqo
zcjJIvgt2ZcA9DFA37ybqMbTIoprM8lXruBCp+o+2Xxkor8NSqruS9T13jG5fkdv
IHh5hdvjUfCyX4Qt1Adr2WcGAdF6YJ9q6zOZ+9Lf2+wcUrBRvkfVDi825UP+C9Dn
/9DhlYJv4Q18mM8EBN9Uq4hTDw50KyrRLrk+nBiDUmgfDAknBHEYOaa2r/AJGKkK
Y/5TL1uCfybrngieOYmHxj9HrZKBTJfR54M93WOaQMzlR2dBGLarkSiWtqkT+IZG
ijS6UlE77v0YZujG/saVjfVxcTbp/AJ5y8NNaR9FHzenmnFDgvsvT7FoIAkM4cV8
2uuhrO4JY0txVoXiods37UQj9i0TrxXI947iXpVEIumdE0IRCuj1jcm8537vqX6r
STavgcqqfZC2vNsDo5WHkQiFloAAufQbyhbXbHBrEzw05KZz66JdOB2kN5E+jgkk
tYwtQdAogRr/8ladkkaalmuZPKrVR+rKqlVUyoZ25ESaFaOV7r89u5huQ6nlz8ph
zc1Em0yvCle7a0M4xU1j6HaxodNqt3AxLD3RHMwYPU2QvINAkcLx7NC1ywLKMplL
ge0CkxBS2zxytEr29thDHE4ayZH4VazcJpjBRsfE2wMpt2A8JftnB7E2tda0uZr3
V1D7N5k9FWi2hAenMRYm5csKGBO3b7xfrW1nj3W6Z8SRYskGCQgKYyCpGzaegymd
s8OB1Vg3+lKKXDXOUt9TrRJ3u0Rl5MTA3pB50SoPXMLCQwpk75RuPRz/XqPOaH5c
Et779UzxfHQdxhxh04btkbmINsRqRgqFyJLNtU5kAbJuFKwU26pZ0g8BEE+JdRvK
LsnwhyRM+z5sZLEUd+nYLVV6hX9N8YvfgY6VSotXzFV/L9785s6wLd6J71ea8wvl
xiuMVHeislwn+7zRzTAdhQ0ib4NOHsOmPgAWeNNyuwFh1AzYCPauWlJUBHFtA/Uk
9wNIxHmDLut3AoxWZpSgQYjAdMAobyRcq997b/6MXpDPG8fjVRsQna8YNsOV5Fi6
nTZIdYffJcBYP4R6hdzgp3WnSqax6thlm2CGwSHdvma0AFe3R4fMdotPMh3b08Vr
pqlzhMUmMnllnrOJNxU4HGd8fp/a+n9Uo9iHWxNhVFMEJzF0sOhpX8g/YrGXILhn
VidwoZxwF3EQ7440q1HgGo6M2Xb/nIo80kMUH0ZXMmra4ktw1orEluUYdtioLwCn
74VZSHOTlya6rUC6iWcwUrsLX/pNlzeS5AbsOzlLYlzlt7TXfD3BvNx0MyiVaL6e
NqypcpOQoO1BcaGIsjZ5Hes+muc7YjivR1DmP8O++8hwzJP2Y87de0dWqC8fOGA0
0q3PPp+mJy86lo697PIJ3SFWPhwYHHh8nc0h4fz5O3KPOQIRE64mkbSqxH0OYqAr
5UkY5yKkGAFRWu+oPlaMD2SHsH9kdduZjdUDj3Fx+4Gi/1iO81rgtlgLPat51L2S
2AXD9LGlmqBHbOgT+7WC/W5sXZTR92VKeY7XwzdDf46fFGy2HMQ2OyO4MmurDL79
FfsRRVjzQytu7XSSRYWIManLOASuQT+bsd4nI9RxcKGQu8HtqSLo6dTIEoRszt3a
PAeILkzfuxnLtYospln7KNCPRVRfPP/6S+MvutDXWvQ7SUAaVMrrQ1h60v52CX/K
KH1EnhT4HYDT90jYaMvzp8ByV9eF6MBB2uDhNEef2yWiHbsNrQycbBTk+agqGUvX
wEhMt2bS1cPal8lToLvgEYBkyGEgkgkLbgi22cZvnopsw3YGlzUFHnN2NJeVfEQ/
VG4H2ONqTkYENRaHrtM+YbG7+xvLJS/F1qMO0cUfURTZkOJCC3fHTfNKkZ5lARjF
hPQAqaUvsEZ3zgRnTqy2tjpxQi1qODvcF6u8CrmVJEoHgDcCh+vGqftTq5Op/tns
f1mxJPmq0h5f8yY3r90I/coWB1DjokMhHQPdfeWLE3xfPesT5n4/uiKQWbKTmErD
Nh25E2Ah8+NO1hDnW/N7O11J8Gjab389LsaVFfW2cO+1vnrIm5tqw8OvXvxcvexz
yqJg0gIk4PlQMqUnEV7mO5mvvjyIVtTTdZkinV0hR0Mes8u9X8Oj59uvse+/IHRi
lbA+lWp0LJMDJpaOp2bKBI3jSnpdUNIaMi2Wm7G9h2IYKYtCs/jkf4kO7jcOo+YQ
WcPtdzzM2QS9k7nUzIIhLSuiRVlMkrrPwubdggcD1PblRA2cCPIsgWi4MHZbCpvU
l3HRTgLMafDxYjFOXGomb8/+sC0PCIYmVqrAYgj0OLx4KStFbV2hBouJ9c33lELu
wNwP8U9xHoYMM9IN38QPT3gP8IQqKoX3iHswD46pij7jJ72VIpljNylWcACNLYrT
6hYRYi2aSP3kmGe/ZQHLdHZD7F4Cd9ZT1D5x7Kf8sg8w/nXu5ZKo3u09SMDMXluT
LpQIhmRggFbiBl/XSi2QIlxF9FSOyDwrqzdixFSuyEqx5EFbuSNnaqFTIBqQZhjn
h7ees3DlEGkiZeZpDXi0WPiW0k0ZOWQJCe9ggtFMBFHGm6CgWbc02ZNRNekC7fKQ
zuTVKlroOpsLNmO0JRAch7cilAFEqPS3r3t3JADXJgdvWKJmgmmJZSayw2A8Acet
FWYOeeugQjfNtNPrMAA3hRE2IGOCyapECe2fviQL2drZ98l/53dr2opt8hjeFwOC
4wbUhs63hthpgUAaT0MujIqs1ylJZns5RphzVIKdGjneyv0ePgijbJBQ6f1YQyvd
dUEstvFpm2axjMgEhJ9vSFwiRKQsbzwr2Sjw0/5YdrUbkZX3CBPNuGB0QX4HX6L5
4Z/rmPUsxDXHbRrsIy/kqia3NIW+CrQQo9C8t6g8LCcfpHX0EljcLokGiMjpr2j3
MApiBkRRuV5qkix1GORUxd/lxqQAYH2E9OMIzxa6JV0nnwI4Ov49aDRwTlC1pOo9
+JLRlFnCxVsLccf2Ukph0me0FnEg3xi2N3r6liNJIya06IoALrPMTz4i4slyEuhl
DZG+QYO1Tg3TkWpjB9X+AgO7qEOi/zGzsGdcgiPcXvb+DydxjEpwlILcomgYO0IX
V4Errx6SRXmma40OytVOyQ+Sr+PHDvM8JIDt5CpBe1ZSWKdemxbUIXTIDFR9dUyC
ZdcoH7q3x9hOajmN+pRWsrijr0LNuYyemf+sP6vrvzqJZpXEoHnCh+I/+WqRR0Ze
IsWwr+3vZFnwGv49Vk2e2OGXQ8wVivt7txDjr5bMgdnfgsm7EoqrxU6z/oznVkNR
Sy9Jp9DzZ9i3oDeGOkUZOFy0LodK5YCJ3SBtEQU3M5G0xPRRw/75WsHn+W/3Rmns
4Hk5nCBhs2VBWbLK2ra2I0mKRw8+TcO9NTkqEuOWeWLuSI5HlDWN+UcGCK15wQEl
BXAF+ONTdxD5WiG1EeBmgiTwmdKaxhKeYYsZQikLsckuVXw/QHwwQuKAIN+IOY0N
vciGmdTTvCvJg/pLhScp9n63oVbZonL5AnKnQU6r+4f/lsY7PYNeW6B8PLFWRxns
82k+7NQq90dbvTOaAdKWVfpR0yDtS/GMxsksLBEcmO2rMSiNPOyqa2eqQ6uvhDZ6
4on/FtKWtWo+E8hAsNVBf8hKI4D+yaycvEXOUhK1eful7Ns9CLpcOp7Jl8VHUiBf
gn/iIL8Mja/oyScOKHJaAbmmMYxRWbPXHeUZyLNyNHr8lXvUICRBKHFWBFanjjlc
At0EPu66g5/6IB73CjtiED2bh+993gdVyF1ww1wxrt2F66LZoplgA+sq1QTVL8g5
JtdW48MoCq1f+PIgY2rDPMsHg4jYeNcUIMJGm5cQbxKm7WNATN24A6T8zbvc1MF+
MK4DncGVyx+PCmxJuYMrEtkCXXTkqn/lHXUCbw+BRvoEfT8Ryqu592+bzORXJFr3
3H2oY6rms16WGk2YOIVLWo3Ml/ZMvSm/lOZt+Wu6WJnjHteknKiN4cW2AFAcK+iB
A9LVJGM0wqhDj/fYMC0Owg2khllzHP5P/xOWwVLXBzPOfwwwXS0ZFPxELft3EtuQ
B2jhCFk7Ambjzr+dM4xjUbPBtoaEUS7sJp9YxkWli844ey+7p9i/Hpp6oj1gm5M0
VSJpkR0VSxjpNXkmP9BPjkNGHYMCelgc8lqRKrpWfNfjioBEVhhOdsuOKE7jFu9z
XY8RbsxiGjYw4BnsV7h2W1LegSM5XE5Aa+n638ws+tEbsnw4kfiV8TvyEBQEdhZI
AUm0omEhTIhO8vnqKRa3tJJuaLSIgQLs36cTabh9UdLQpRBqXnobcPlSDPYTeoPU
uTXTJ4WhGCEqTtMtoyUh8db4eMrRCM9aovu9V5McJ6spgGPecAxXcFI+TrVlR7qn
2ZNAOBmOVU4WqHwIZyTrDMb59N6rJo2DwSUdnRQyhn5O+ZvQj6MhveSRhdcrquOW
xExbYOz9gUdO+Q36vRuoifZd56gWUDPQUVKDq1J1jnioAhDqGJPZRyPiqlchxXy7
QF8VchHkkT+FZXy28YT24KGN8xD/3tuReUsd/S9iq5FYRwhV/c6sLsFwICpJ0xOV
D95xj8LfKdiX4SclFjf2nypfrk/9uJ6g31+darQTJZUNPxIk1D6AdxBPeoQLy2m9
rJs6A8QyItYLl9KKVJgcqi0IIteCRFlKnDDDmR+gFG3Inj1CMElIAl1rvsBWtcTD
Pr7Z7YAdC0nf/DAcUon9JBaYu2w7/V3TlDHwZ7xNYFstCoyRLdxJrjaay3fTQugs
z78wC03F3KSCwHm9IHGqzJoJvGNt+XTtZK8n0w12k3NXE+2eujchs7cJjRFWNvkF
HZc39wLXsXqUCNF4zox95qM1rZHHnCleHZrQ6Z/AESpf8u4049wygy3dLn4VcMJx
7NIw87IxWkdAO8be9rG36b/iDoh5F96rhHH9nQTuoysVCq8+efA0MjZmQmkMEa1d
5wpZDMkdkBE7izhW33ZvNa8bB34Rm+6uHykBTrMDR1iTaQbs2MQB6Rpk/+zlOSbx
9upDFOl2FAG4T40QrB65ZAySr5zgTemhO4Kg/DJUeI9/64JPZLwtcfYzoNjvK8RL
HblAk+uN9my7pUHHEsE8iVbdsiJ5vaQId6cT2JTzDbawZxHDa9qFePSCFgQ53Guy
hXDgeWNhJIaL4OZI65hAImZrTOxtBt5LYvh6q2vJX3XhJTHco0hhR62Wv1IquihN
vMSFup4B9U53nMToQOwTJ83WoYbbDJflyc2WRXBja7hyQEpsMBFQDK8UEnVfDMcb
4yfzyyCQpBosewchLRImRNbwyRoCWqof1pVqH4ElSIedx/JXS6+uhJkJz5Cyxejo
xpmp4CQqAKytrgDnGQiTJCdoaFstLMjGJVJk2gRxuwcvbLtpnhgv2kDU4shWm0e9
nGP7IYLc6xzsR8jim+WkluNfQnbM1iSwZkU6tGA37if3gB9F9ZwJamiiB9QwxsYa
KTggXm6cEED94aC0WliUDhN+TZCneTonK/Q3KdO4VppXMKIUySsBCztmHm89Tv2X
w7Z8QjHeuLzXNupJ+BdI9AhXtAQQ9yP5iuhZ/ufHuAqNWVYl9QlSXcTWGhY5ZFZs
0GPb2vDsZ7VcZYnoAAZ4W0Tn9YQruv5KeOPKKl4A3R6IMbe5lycaS8WjlJSrwktS
47X/RERWWGsPIEmo817OW62Seil4euGZKuEyGL/DLJ+vRO03jkGkVjyMSw+BhHIm
6QepKNWPnSlJ9+UAHxatlIB7Epzg+SiQg3EE7DiUOnj3HXiLMrYzmArFCG346ZYq
vqO874BJjRKnj6WQKAtKadVD8d7C7o2zqWSAWYP+5nmGv/5ypQyVOh/GoElUbYfF
QjsqBCZ2oTH3S9b3+Y0Mm55I2OK/bF3FDqr8xSMGu3CRn+blHzEg9QhiEiINFENs
+8d07V5YuIHd7iF9zjvoUbI+/gxJRUjm+wSkm5spxeKVcQvmP00+b9AnyDbskqDM
VqKZ+4B6kq2NSwAsRuhBw7TxaqU14Jpm1OWkz7tDzk5JF9eKOFhK0gsdzaPDOIen
0Byz2uLvhHfxbhbg8QR+onyGnSLDN2Lu4lM+cTS5fsFo3OL0pjrewhv/dYEPhdCl
qp8A2SgylrNaQX6MxkOWygl/YZvwwdvWOOcqrQ/JBLZJEhA21xLw1zYcJ/6k8CkN
li8G4r11Ig1X1jUf4fuNN7GwP/VGsshHqa7d6HwS5trgU83j8V19Sk4fWHh9wdRJ
Gk/Quuxm6a3k8tXDpBcuhZazTtb0+4mEDn2XWnipm46cAWQZt8eqeHb1RlK4aMUC
a3tjhNyDBLCrVFoteNvEj2xX3hY8J1M8zAVssn4SjPReBzJHB8InYkG9a2rRth6B
JbbT3ZvCRGmLZ2JtYTiyDzu/J33uPcOqpDZZ/eqNMqwhcvmphHOOq+S2b3qqp/3g
9r7RiofMOjTJa7on/3nWsqumulCzK8WONjMJnqw6xJThWs6dq2XSvRTlXu2yJ0bI
aK5q47sOc7YpwynvySHMYY4POFLDP96tDWrg+BNOg0g74eJ8A7uB/ZPBwq+jdRBw
AA4H6AgzTuKwRnS9GYZUm5ZyDYIdLk++f2hrKa+G0B7qboIz/l0OrmJlCYWGG6oW
h/u3nhknu4NotyBm5kNlhdxcu410pIieQ2TgyMf1SdvllDT9bWF01kewX30xjz5I
HgxR2Fz15gFKAzMeg0DAlSrLUBe4OQHFO9iMuehNqeyTz7nZKajUqpMKVcUSsVQ1
5VL54QWaLNAF9hhDZVd8UNGeHXTSq0f3AgRBsoap9faQXy5d4Kzcrpw+i+38v1FQ
RrWIFIdMiRlqPujfiOTZI8m1Y7Ab/Cu0cZLNtMqif9aF2GtrOPOsRkXY+KdlKSrI
xQggStK1VJOKQ9RpnCyHj6+OZaEM4PrEOB4GCPu8QaoAh9Z/FeCfvWAk9w4D+1a9
g9uyubENg/XNDRo/v8u3d2B0OaRoJbZPvJci0y1mA647rDBTBErqQjh7hVp1my+Q
WTlBpoeQNTnPS56JePY1kCVKEOXnBQG8RuF5MnYaUkXR18xmlNfEQ+g7lqkPjAvN
n/hMekCt/4PNDs4SxqWR7S2U5wkL4Epc8NBokqLqUg2omG63LgW/IMv/3+hAVzcr
jwRUd+1/gQe2joG+945d+grNQjlVlmw9hC/ByHY9xmwZjk6Luh5bv+jz62V0bIWz
W7BlCuEPPNInadVdN3gps4cTOJy3I/eEkeTssSr787u3s+hZceab3/AJcwiAAhC9
GSbok+ceI+Sw3mnfQLARQ+/TiKgSMkUsvwwps6JAPuG4xJwwrxHPLC+9dk23kd74
XWs2ws3O5sbDKqCztrQ5QDAa/ePyMOv9kZB4uRIvHHCH1OWhRcz3WwYXtUE10+ky
YexLlS+74aZsyaYDgoxsm03xLhP45AkHRmQx3lQUVG498Gdj8x37hBjvAYicLqtT
roKx5jNxeGtyB/1Uc/Nu435Li8N3TBzvewnQyzV15ua2hRG3xHTbUAV4JeF+Fkro
bvNPhSxNG8HqW/530ecW+5VyVxSw/BYwiKKBCtid4EvHiiYMxeKJxY9mg5c1KXr+
BRjVUiF9NSy+TdtLRGr74SsJfbkC+J5fH1ypMT17yqIvtHSs9oVlAvbV7NPtPUk7
DscWiM4rTJDtrw+5h0lfEf9Mxc/xQ1K2JNmbSp0fmdmq1hB1TUK/FziI+5nPUKX8
HxLtRvHTe+CAYAiQwdL2QZMat5VFAI/ZTucaA9Ry8ewt5w+flmVs12im3mpLTFBJ
beqvpRgpd4qAwTWg0S24nxgEGQX00B7Jy34xwx4o4ztIsC61ZVb4alyZuHNYxHUu
DTmuAiZAMmAp8YngTxiDsyi8rQJsyY0x863OvRIbHfUg+j00HcoO/t7dvy+g9LzJ
tDTY2odS/YQ0gSOytqXvadg8o1TLBfnUW8PUmzZ94msW5qxT848LNa6Vi5x0K9U6
9Rd3JVzjLKRNbUFw7leZgFAwXG5ISvqvq4hy35O3oq44tESp8LWhqlEDoDDSsRyw
i7/5cFqB0A1i8DzjsyykT+sTQS2bM9zGIfanffrIiaPSTU/3SX1Ka1Ejk1k/rkBE
T5MZUDAv/ii9x5+BuAZB7SwbUOZWAyQQq62GnIcPKLhB61O3OJfgSRE+TnjIavV1
HUTObwA7I+gfsl8bbpzs8rXbCp8RmwHt9AH6VYQB01HyoVZlsXSrlruq8hi02fMa
RXWbjsE98EIcfop8GcZr5ZAG9JmLaLLgnYo7QL7L87KOis+m1pC6501wfxZdzgrm
8uYfkuh0vn5Kg3WfaFeVpfVADXWhfPxXlibf3o5gyNcr07yujBwK/T8Scm4lwNl/
S9asC+JjGOGg1vde6Y3eC1PZf9wpfRRH7TUrD4qakXEhSzoKI4C/BQA1zMmObMy1
kvAl2rX7HaIvJIOBeMvQU6xbziWUK4UsxZIvmWq5i4FA5r0svmaHFLbEG903oTK+
s8G+OYVVBzMSwgYSKwm7MM6S2ui1ljdJQ7gGKVskbpmrtvXG3u9X3AirLKL94MCZ
kJo+PTwNlxj0SgApXwAe1jj/PI0ur9Q2uvZKPeSrWH02IfcISU89xSR2binoHgps
YXAgemF+HX+67UUKeAkKH+1DyMFFYJLlPl1MsIPfQ/R6xRhVgCNK3ZLA/LFEuZKs
2J3qsbMS/HSg0i/Anq+7wh6crkBvG34UH2MElGSEnT6kxm0Ots3O/FPRVWmF99bD
e+8rnKeUBnwL7UvDCnrNTunB6iKeJuaiV0ICRIxygqBk4p0Ypvyr3ZBDzqCBQ1Sj
JxYU8z4TZoGyYh7+4DpUgmLhIPg/O3ZF4vDZV7qM9c1OrYc5+nlGCZsNQnVpyJUX
r4rFA3IE3IcAWgp7NiYvvclCh5ym9LsQCJFEWlLrqm+Hw8LdLDkrbYVeuBLQz5v8
XvpU3wTA7yzh6PIpm9QC16Dng8N9WUmnzoR5wKJVX4Qgf/Qfnc433+gS0BQEQLYK
ubR+z+QTFhecx2c08XgIvByrTMAHyistHA7x/GZNNgneVv6DnwTvZtr2thJtjk2E
1FqRCTJR3de+VXaOFr4G6/8Vjr2XC6oexSZKBlDjJjB0SV1Kd8rjyqK4ONpn05Bk
h6H8K2pIEFk9lsh284uitB2e4LUCNQsfFPP/iHaPebm+9g/OR/8aTeKbdUsLg8DY
n88p8Sse2yxEIQHXIXShSLZpT1XJZYOS8x72YtiGNlhxapse4oZ/pEinwA3PuYiR
FGkY7ItuwkB0LaniyJV9F3ecOfwkZc0QayICQH2ue0M69gsSPXzlqh6vnTtYuEu8
rRJ5taljwqsicoAG2ULfkibl/7P4/Ik/HelZU7r/0EN7p2dyQbAddfLKac9LTqUH
fUcToos1dXvuBFTQRkZEIG8+oay5IoabmWTMSz2si2VZSEFFIHl3+aFOliw+gzG7
dgQ7YrUVBijWDNADIGlQBlJxOJHd+cRSkQro/SDw+G3AQu4QvUx8uZ1ng93zbxhO
P3wj3qyyQg8tkrKy4lyaNjRrO7m1KvafKJIsbatEqaDv7sDBoaS0hbH97Gy8xHJ5
ZC8ZdXIObB/wdji+96RU6Ul9wEgVOf8e36ixqWBACSpdqm8mtbAA9B6hlMM2d06l
HjTM2flD55dQwNJ3qFI0PwGZOHfFlrazg2LQwXmVZm+CQYFSrFmZTYwHKj9CASii
4E+53Ex+dwwxbY4RVl3WTQ0yuKzD4BjI51SYCs0oGUIKWdPa5+pnG/hdVKLrOKRa
wUtGgR6TbIgQUBkLRZvEpvDOCxiveWpnAdNijUbjOfm3OeowVllZ3hQcAGVlTQR2
ep1L0657yOgw1vCg69pgnlau1jfvikxHfHoAazaAnxviKBFpLeTNFsqOcdiChnle
Ni1cQje/78Vw86SIs6Sxy/J2qq19ZbNMsW0u9aHTkQrIGV6DoH6/4mkix64YovJb
GlsHukBKu7aLE5fa8W/1xI3PRd4diUhSQleHvH7DttOf4123CBhJvQbx1Q7Era4o
7TDMnVKK3KQbRXkIKBd4pbs95fWH9Zv9RrENljzZGORoJFnqFhROJvTQ6KEfcfmj
OjMWRfxaj4cD/oqMfMOw4KmOhKmuYe+m7XtD8RXdByOYmgTi8aS9PqDEB06GL7Yf
ouOUfsh9WrQtUddkC4chmMGy0iL4DT2FOI2wdixJ8EteVLyNZMMnfCkrynVKOGQt
zLeiwE8Lew+eQ2Nw3Eg/TQ8Z4+PLikmf1MROMP0cZDTaQ7RmxfP3ptAiDXC4I/Vy
eFLRZscCfnQPBgDEIcAdc4EWFc+pZASFvysFT9Ot5SSQUD2KTg6jyt9LcR5e80Hi
nfdNM+OfHMuRckyYCx++W9N3ZVxZjZqxEzyomoPNBg7a1ce/xJkUjDAU7RxB4l7f
h6kTs8HaWcv5o4/tlk0aQqrl4po+hRRu/YODLC2LBmEsc3AaG4YhWt4KZUH7SQJd
NhnV3bQ/hLK30XDiYnCMWTUEV6WAoIsMOc71gsy1gKVSzDuJjlbH1GSKcQ7uVKVQ
4ip3yW+cyGKAdUMNPNvvMdh3cBaMbpg0jS6QA8zIPMQSrPwS6g+qojq5B2lxNB0D
LFPlsJm0WQpkLNtcAae70wJtH1h4l6ZTNtkRJvPepZqgMlHvXPjoZN1VqDHoxSVM
NLZMaG+C+0J5exULKbMctrNNCf3bAbYv/4GgSlrVxBI7tq1B2gxNER5pyy3sEUww
uGHVm08AOJNCpODOgMTpyMggyZfj4zPTACAVhXc5H5cwJa7StIqKVe9NtL9pKNIo
Hdv0ocClEb/6Dc6ulOeuZ/ao1Il3OpO8ox7N6vTmPyFQcaeacrVIzl67NOg8lGhW
CYK9tUQSFvRfIIUG3a6SLl06QL2y69gVb5e0k1Tw4JUGlblVyKgCh6V5R1c83YOg
Dn9i6Qaibjtvfma4gGSOP0gMA91ihD4xsdCWzeneGow/1C18M4d0yGL6E4t/zqkB
u/HL9lS3UBLTPdTr9EM/dgV+fzigaEH0hE8tvhLO22ZXZCjWrZ8qrDyIxdj9+tBo
aCFrFsb4kTki2l4dl6fnjSLzV8HqH00Bt3akH1KvqutUpck51g5HcFVtLqnWZF7q
bRoKJwjddCT5c2K/3bEu0Dmn3nLPf7ZZLmuKW9MLxDZVAk9SGWAdSlFG7PDxalsm
BqfbW0WbkjjZ23WNlkMHFN3hPjRuDt6wfT35vZRcFiPh+IAgg9VeFRR/1dbOmUQO
FNSSqq+AxkM5i/mzUnfGrgNusut/fgSTF9OnRi9bINcVMx/ejGD/cndOqzlu0yM4
rjTy2sB7qJVJ8K8Lx6XmYLmG1X3VSOboAnffZh6WLL6Sxl99JNUj7q3G5rPEJTMi
FEIiH93WmQeKHiH1OETwLqG9pxLt6TrQchJ3E68uWmS3Kv51aztpI5FYD5Ii59wY
Bj8c+q0yHHJiuYz1CL2EFeWkpvgygfLTEjQ3HLdCokQCQNtRmxtV6mUYbrojoFIL
bhxQvHv/knxDafbquaM9yxGvcJL60DMNa2ulgRFcm7r48Bh+Kaz4eEHvRda+UNHg
mC76jQwgKw8zA9loXUv/8XTWRVCoq1h1bxiZCR8YcwdHvb4Cj9s2tieD3Ae61LEM
s4GQX/6eRoI5d8FwdNMUBBL+QL+AXL05B0rdiXaOIY3v1UHue7cpYrGURhGbpeOk
25jMX13KfI0pxl1sArcpFxg4CfqgBfkoCawzI34/kzSM4AAYzidc542haalcohJD
qzoRbVQA1huPwic3IJEHUI3f20kHy85tF7kjpuT7E+UO1pmG0NNoOEHae82OQPQJ
nBBE9LZTuR0Mxs8OtJHcfTCWn4AeOlyoBXTWLLUJHake0nwsM2wxq8mNl/yMOhIP
yRRE4RJuH8rUWpMAif8BOxYAr6scp93PG5pMi5bShfA93TEH9Q1+vCA7hJbahT9k
NBXa6NsIV1zXbU8ua9yNNyp9B9W3z/VQ7X55RbYskdKh6FDMa5ZA54dbGz5Bxm5A
X+YkZGf7rvYhR/GD70+NKV8BbKQO4aIxEWfFurHR+LKNr2jGDN/Z3NU4+R18YInS
XFRthW6N0RMkVd6zxTq0W/R6PjHkxmTtw8qSAf/qkOh21dPWvKyOYenP+HRxHUwZ
FfxNhtuUi35mB1HJfukeZNH+L5DjvoPBxqCfUR79QiWg0U+L4fu1IKLm6bvivF8D
ASNK62adC1Oxg2ujFMiA7TiGmlHg32r8WBH74mpPF1LGBKV53fWZ/qE3rJvqo7nN
QA48gCJp6Au+osC0bZyV7ouHUXE8NOviaaI0/y8PUAYlQA0TS10DB3tct6/LMNk5
1s5mbNtLUMTUfkj05+QAC9u/xCrBGPOIo9m0Y5Lxh0Hk9cet673sEdo9ZO7JmmsL
mk5FZSyaAKKoLBiS6R1KPV7tRd9j2ZbKdO9L9TeYoV3TuT4hQLn96s/i5DFgyGKQ
gweb3fsCOVKPcFYtJvdZBEWJKdMf7Gg4YaxI+TYhBXZ89D9q/nawbwOO+BjhJAax
AVVU2eJd4CrKDTshdF0fy7PAFpn/nlQKmJkV397zXnYKgnLw/JtXvlzgXoWMI2vu
bwp98cfaM5Ib17F58IwYogfbehN9EHMm6cLLu4mdiWZr8GCEjpghqjF4jimfe++b
LSrsLzCx/JtD5SqHGWhl6VGI+8j0XLl/GCjp7R/nz9iSCaz4qeCaibfpBD877+P/
7jfJT6k2ah3+eYNXML87WIPOpE3cULXPkAjT7DlG0GiceulOlSpVreDti45dsnur
tebKCSmsyrJHRwXMQXoC8XZKkB7vQC8NOSJLOlpKkdLLEvfZX47GSKu/9Dz13M3x
u0hAidWC3DlV2r1bKQQ0DVP4gxF7PfCaT87Ggw+poHda+qTePaNO037FO912Sd+Y
+pOKoQDEPsOJoZj9nIvvwk+lngi1O0Ph28yk9RYTQQ2IKHchlLoQkoS+d0ILkTGf
sNMIMEyfcg+qJWNfWENgMTuSM6fTjso8dFQSz3/sgxfoH3XsKtwuhIGjNv6Qz/JU
sgeTlysy6hPchFyAyBTMS86k8cJFWs62v49CoOzg31+4h2eMAIZgqUOjkp7e+ED2
SwWY8wvgvDsd4UeB86l/Y3tPwkQFRV8bj2Jzsc3aMhD/eIBfsCNNKfruj+6gGuAi
JIZRp3wadkzuE1rSbr8b2hu5JNlzspdWfPxDj2QR1e6hvJ5F4ZEHLZGjt4zpxmc/
rULQ080pGA2ArqO4vkP9+/iDn5Eu0JKy7a0h87U/ho4iJHkFayYlxwNcyo9ziK7K
PXlp/K2D/QJuOjVpssbgOCP8nxHRrHrhS3oEAV351Q4ikAh3mSYi61GltopkGRiG
VZ7tWyylgzAXyApVfXYvZcPIxbD04NJ0DVpptBEzMQsVvRzem7uUtEIWMf0dKw0l
3hi4qLwAB3NhZZe98ZJjmfMmmaUUml7/KPcW77WHzNhSwPNgSFNIBQXQ/fdSHjNu
aDLQOVcDaMXYC7ql+2M2VjYtXI7iSdyo2LRG58AfwtV721LSmLmdjWez/A1RYNpJ
Uxtxo/HZTzBP2X+9kZIsk50vC/5m8oSa70FFREAAF/SSE4p6IoDHEOuJJW71EtTC
AlLHilYZq+/1tzDkFwxRGZSzI2C8fFF05A/ZQlXO11vHqALiQWedA1VJjvUycX/Z
3vP9ZBMPL3XttdRRE96ExxbhQMpLL5vpck6ZU8delkW0LoPdJhAFTxy3ioeUS9ka
QkZBcHtRZpDWKE5KpPUxiwA+zQPlj2p3XJnCScKSC9iyZH4mx6mVmfdqVJr1sbcm
liBNYb4Db56w8vrhU77kfdv0dSn5mfoeJvSoH9mRRPOeENwZYE9jSbCrpz0dN4sT
ituv428QsDcPTR2GC0CnJEFHISaziN6ImQutFFaBxvAcN/GnC2XEZlgnR+2cHGVL
DDzeFBu/ec/LCmQ6kJqJqiDfWtnbQtCWE0WvbaFyg8SdoiEAFRhMGYN+i5NvoJiP
nB/hxgxliutXFZuolWbjaqiv/UWLpgJ97F4Tl2AaTKAyjO/9MWzZnuwgbEE3lp+U
PY0/AnT4Pv5EhlJNNoeR2f8VGWm9l9R9NMSTZVm/fuICBzFMuDJMPIHoIoA5KCtR
AOwzf984OuB/hwnUoStWu1u7HFd9S+srthhTLFySMnqNxL6TbUK7l4MsjpUDlxR9
i9SxcY8JwK+bYgHDNa8+X5nigaibA/yXxnBlqBT9vnwb4K8+qb34OJSPOTlqvZRQ
WNO7qaWwn+Naag5hijLs2/kbKNZUwcFfFuC7o2Z43g2QvYb67LP+GMlJpH6hE5Yb
eFxplElcXak7XNwuAcoblvMM3vVNA1pqUdtHLNc/bUMI3BfLMOokw9hVR9xiAGBa
rFSh0fdtFDfMENiEggpmWPIsP24TgMeEdyOQn5vLeJF5rt5KTG+MPGFLNprQAQ5Q
UmGadLy4vxYe+5Euw/wCwkVdLpXpDdrtoKiD1s1+GhG2fPd2cckgOcT5gfKa1wjl
jJr0Z1zDYtMLlshETy8UfDjGmaf6gF8ihTfBs1gkdhkkoiyDhLHoMa4c9c3YGKco
yKcw4RYxdmdFX8IAHppgI2uLSSTQBNsfHY404jTI1jFBfRk2IkxMlmvHNeHHRRTy
bF7VxpaBvt8g/gLnM34yZQyLB74wNhoxaS6m2lg9BeGrHATl4u2GkwwU63dvHWOq
QDGuWv+jW5BugkjXzMrHLQT5Rv052r5tVVAMpUWHq9/mNNyEg6ARFRr2nOat2XKt
nufhxoSyHh7Lof+VgTa0WZbZXx63PYfF+/ArH9xgnn6PXaOhEEUbWHQmUK4HdRLr
JZJ9AQFVzQs2v6QtzoGYCU0w8uBFmefFQHIdFHLDhQFZT9at7e4j45H2zxD+BTmV
rPrGUx6k7xyS6wRx2eIGdB/ewy8FNiNT1sz3oRZyMhh5Shcb8vAdm/0NwBf04+Ca
/FY4O/bzihw55g0XwPQPb0dEVH3m+VYxKPfzMvBI/PZvK9fhoJY3JMknQmCOvJxd
BWVRC7vLzcL+NJkIDxu+xA/egfR6FLSDv2v5jxJ6BxY/yfjaffOxl1+iKcVMcB6q
qt8gkDN81LTNN8CK5TdrzWYOaNmSfsRqH6vfazqpbnPhNDy0EVYAGoHR5yr3Hng1
RdwawLqxf6JNpMFHBmtJdb7QI+l1qdfiHKmkRYy+hZ0ZturN1WbeGRkP09z8W3Ub
GxDcjVFXrBXrxO1HLcwv5XrghE0GSSk7K2+wVvF4nwlLwuMvU1bLoC6VULKYKMbf
Dn//Ez9bRs6701YHe4RyQiMTIZij2b+x3mltQmq03+OMM5sW783fZ4aq44C4uBRx
Rts2dqulM7eZSdkpo30l1LuplKsuWWu1JuP37fTucv9I0DyuHrpKIIHIQoIpl477
XtLjyoflqTR4LJpM9RDiXFXzd7peTXDCih+//ZK1Lh0KNaGGyhLAhwkX7n2wR+Pv
8+YRkfDv9Puv4YGQI4yMUMrjrB7C3xhihwKU9owSkcK3IpnM6d3kde9eLYHYG88Z
Vap6fwROB6GQWGx8R6d86Ba8rRhxCxHM1VMogMF14xKDngoa2FYnkauTEh79N9qG
HSafJJeiQnFyYm6p4O2Skqb9fxXhNsdixcpVZpQqJb7OpJ0nXQIberqQeErI+U0P
bzspKmtEtHqI4Viwqmz4DqkWKgFvUDpLOvCbSZF6MEUnpEyDO6xn5zd6y6SlZBa5
XdOSVkUJm33U5G9Q8fI02kw1R1nnbeYHNDEclUHAnXF+uMiwnDA51oGG78dZ3amT
jrcvOBhw2ZDe4cH+J1flKCDegXDbzgZZSoLwaKOU+JMXtYjFPAcn8l9CJTR7+juO
fQrPY+nMyBO4cSp6JJEE+yody3gpTxFqXgKltx4ik8YmXzxrnO0d/VUhugrsrxvd
K8odE/hj9nE5SoQ2P9xIpCzvn1mCcmo/7CSPJcF4u72FNpr8OVScH/pZIYPhx2aS
9Gt29Tii5FH3nGjdstCNoRa7n5Qafsdy7CSthOeK2dZFQjaAGZN8QP6BPLyYICld
z00VB6KjXcr+p5jQWyaEeY3WUquctNDe/mBdYqG7eeb5XUagHMHtvL9YD66HZs8m
nscH2pr7owpV2vCUbJkn+7xy1RhBRtXoDFIYcCjEKcJQCcRH8actfe+3PvGQG+6u
GXKrj99fC9HCYlua03sTCUluj/HorNC7ODcQR1Pz8+Uyu+TRy/8h6e/+9UZcFNsc
HE0T/2su/aT6Kiu5CX1+nF6TbOHjppN9u7u6cRrUwVKduPcQ4AyQH0fRNVi52EOg
PJyElyU4IjKtUT8WxX1V0aOjUmkhPMKtmlE6kEetVUcV16AjMspxmro6BC7E/YWy
sjKBpRIhih/gqztfFRE6oW4vPVLzG6cFlE49g1uyOyzxjfKxoxHGzVaGFk61RACb
KsvLKqrs/QiMeMotKey/6PGvGgNr9Xo9sud00HBZeXJUy2QJQdzBwAYQ5OS2h+qv
ZWcOhlp5T7ZApzd5cZqcSUhPnpCQ3R9nwHesuo8FsONQxJ8rUnWu4PxofUDElyWN
VQ8yyD+eyY1r4cRk7lsanIXrGOtEOuCBlvKObCAM5QVK1Hojd5JRYi7iOwo7HXza
8IL92z+KwaeVXX2yEBCT0JT3nm5b3wt24Z/hzcKIAp9yVVbmcALE5uLHt8Z4ONj+
LzQ6r6YFRN2wzgS7jYt2CPNs0jN5qJ7kTvfhxMUyuEnx5g5OELwKd3glF+6lmayQ
1LhlOwUgz5YIjumImWknCCBMKnRsl5HWJzCB3OPBHRivvbimZpk19LjHA5a4brgJ
W6tDlAPKwUQfJyjlyhoBgAztVnC/hp+XHSeZx8E4nTlk+/VI7f9VVbM/IHvH0yuU
PR+KiYTZbQhvzqdPpYi1x2EEQAJ2/I24pDX9mwSZBTBIlKUwrmPLmRbL18Bn8jFF
5SWZV9uqCeNXKyKogA5YqURbpLk/qfZ2ilG/zXAf/cp9DGfXxWhehBG+QWMYcHkR
X9UWhSF3QUD+7H3Xou67EFsykEkL1gObdOGmku7GQQ7BloM5Ccmal1gN4gfJ/r5r
Rj7PtIIz1dfXREOoe/8aycjS92PHg0FKQEL12Z0dgA4Q3BRVxy4llX3Na0Ouz9/7
xu+DeG/wdhd3/40YWTFU4uDWPeSDAgoGs1Cv7T/lfQW3oq7mo+DheO69M3Fe6Huf
tDgKTKedPKJn9iayF8zxFlj2jnMxUC5IsFfmRPe0uRxawO/n8dLH3ovqPEVVsSUv
XE53qKLojYZhRSv1l+MaLCmWCyh+DszCJMqiSb+6K5WIIIlcSOlIyrlPmJsYhiVr
jZ0r4kPvHj5dQO+JI566HnjUcmbgiMZ5h4y3rbxro3tL4pKTgYroE4W2+xMX++cg
IiDx5WIqvu8iYq9nEgH3mLlInhwqpZ3UWnbZtfHdzd3QA74h0bqS7PmLcpfh0eHQ
K4oS4+RQV+k6t2KcLYoMELwX+EMFfofkkrr9SB1vstdJzE/ugiLX/fRmfu1OG9Xa
KOxc5yPFRKhFfMmIUnL7uvLMohhVbJJnXFCGqGHN4K3rRO6wxzF0PNGhJTGqy0qK
vo2ETrZz5DrvakAvb36RJSg/JcyKa3LGJXvqKkXMkHoMa63uBqPp+AqwsVzCIktx
2PKQem6Kw4NJ5z7cgXevtfes9hNVWQryVU/hCXVvLC+He/ZMQuwdLk0V6Vl4foCK
UNn4FwR9/l7Y3L+nXTkQTUiBWfMwgQFZs/uu9L9dqSbG9RAIwzcr5TgntiuSAzIG
wGqzoBT4+AlktB8h6F+B1PbVGDYf0jdULMESIikhWmlzFExLZvogCljWah09sB9I
4HNyrOASLtqDOoem+kwl66HLGHqvZiLQBxBpaZGIuOEo4tornKaQCBZ6oZEZ9Lz2
XGRnydPQBMOBE3XnyBE/XkD4lATAiWr1B6Kc5ZVsOqOKUJ6U1lF2WrXFKUd1vORH
Z1WHBzGVBPb04foSxyIpgN+5bFQ8dYQan9iQ0MJOZbSs9gWa1ZHZ1iT5N8eBO5f9
3IhOCrNjpX7ho6NMYkucGfUpdVmcNYiJWvAgoBBhc7xhYNiW6X8CSyG/2c346qhu
23Zp4SYKJ/6hz2duvFhmKTP5a5StMcFdGdxUNRqQlTSnEWcibwG9vyJWbZBLIr16
KPIby6zFnJC6RnjqPvKtrKqUxhU2AGVZV0Zyidk1usp0ND2FJG2kA1RoQ5DiCWCq
u3WlXek3DJHMDMAk/wBu/RbS7hRyamfvIvHGqnSPi19XWiDZaHNaGWhPMuZ8v+mk
XAsQVGgjqB8VE8tv4kPQUFG6eajuoa2HvthKxhcMkTuv1JcfEYpGd+wmDqoiO27A
GlzMr71hYQoOPJhdYxQibLM5Vxp+dyXJ5hiiPVL5+RhsSQguiY8Gnt0rTc7gx1X+
kzX70likfQwmSud3Fk9v0UQDlumIGDtyQkq8dc4nG14yDyGbjzvuUe1OMqezqYQ4
iyhCqK1hIPJmJqQmcbKhw2vrrHPOb++tZKQFo4r8kO1NnIaGDbuhPRrEuwrhvkgn
LDnPm07j06ShCA48i5uQosun6MQsAN4lDB7Q1e/619dnpL2yCy6zvDUFOy29yRhF
7zsQimkfp8X20n+eqY7cx/86X2YCkwpW1lcXbIlG/nN+zzAjceyr5eoEvNKcDNcx
UBCnTZhCYIpPF0XXdlCh4SDfR30OIr85Bd8JB3d0R9J9juHnWlfD5AXPI5uU2iSS
T0up5j+9unr2BnOGmYIbgU6bb+RzjOjw5gPhQuH3Pys3YpkpNRGFEL5zySZurG00
MX9Pb4xn7xK8Nu2gQ192bcIq7m3Ojd2JQdJSbG3n9roeD7lSvzhjL+ieA/1M0udj
LEP+tWI0j8xSvIexIz0zlSLvQOVZAs9KPjERSqxKHJevrQBrlOfb/RhxKmmsLf7A
SRJaisk0H0gamSCFxjvjrdMQq/ul/VxWxHYmtOgdd4FRQLNv9aFdR1KmIVAA0atv
XKlPPa1zJMjsb0w77OkJI3JGIJSLHXGbzMPg2YyMgYDv3L6Ry9+Ft9jZzD1UiGMf
DM+y3uXI79Dvl5qShmwIC2VjivkNhdZro2dCcNpm3+p+cRp5qI8GkF9ogvAJ7d+J
I8hJQQ+07dBpuUHl23PVz5zDWTHl4QD72OMmUS5m/VGihAcIke2WTLN1E8deEWQH
oiMXW9RxxYdmWxuKyHu0SK+U+Is9lsKxLysa6fbQIDIRuL6U62a1qtTEEiuLOGHZ
fNKfjKVAmNRHz+bqltLiUe6WgO9tUdLllpvqyURDw/czPte+el2GPDIsRdHbYqPN
GZwmTmZ6K3c+vtsngYy16i4iYNKVS8htTtJkMbIxySvzebUI6lbB7mQsXUfGbaNi
Nwp491K79kEwuHqIEXXMc7J8KAb+X4rAnmbafZnOZO4ovuqERQBGcFfQtV7h60xj
6bvNqDCxPV5NeZZfXaYqLIPGYSQ2OCR0sv5cDDupFGuZZHorfPn3yMmDvC4Xj5dl
creNElbX3vZKz4SgwaJHLASjeU+nra0Op2uClnO92pRfVfQtL6sHq758ckqMb6KB
f7dyDw8Wz1dNdSAelOirllKlGM+UhTlD2IZwZv97jyOGGITGpXdxbAHVFWLhthmI
CubeJmVivKj/LstP0tBJkllkQ7oYrEqhPYNdU7ufwAeUGUW3eNg3qU9eGgEDz7pk
WxH6LwHOQrJgaO2UBoFPngE4475ffiqgXcvZyJ3Xc38H8128Skp+8iLOP76GUm0H
1cLecS615dLXWzI1bgfsb5R/sHVHl9mL8GTPp4iRwbd5Wo2iYet4ndm0cYDLw0K0
9f6XDKsqe0tZrp3yfmvynHLb7+TV2defTw9MrvNtBXdvcnHMvLb55o9JQ2p7SmeE
D5PSKmH1iiiUpQdIpbujOvRTt7RAcEeNbEGpAHuvgNOOQVDlIbpSmkBtIrgpxTO+
X/y8QPV39h9gCF0ahr1g3bPdDlUOxcC9n/ylN6xgrHrHbN56tnt6IqVlfGArKEaE
0UkRmlWjQx188k9U2j2CXCMtTE58za2vj1u15NQhre4HMaCNKWY9dQsTf5AQQEMo
VB1e/2+W2mPd6rupW2IF+PRptXbGvhjSsdyD9E61YLmr9au0ONah3u9ewjYLzVt8
8+aG8Wc827GcVx3BPrMlTZyO5yFe3UYS/tZ9I85D0dHOoC3bZRkw1kqLxdn4hEme
nVMjK7kw1pjOXxG6imfRziNqL9h53CjdgBYOHerPzmOBJPc+cIX4ICh/IkGR+1iV
Uk/OpEImcBWEv1ZQTUkVGQFcPLPlRhmiqTB9Dwq45hyvPVlhom57xARcfITQPgBN
NK5osHhWuO5/YY7CpdmNyFc1VZia1NtLImBuVtxJipFhd0Nk3O3FbO/irO0EwoNQ
OUCg1QPy8Sv2LG+DoonoWea85yUaPzt0VMwF16H3gpASEBuLlLWG7F5bEzWFBInj
sc9jtxMKm246sYztuXQk04NewA0XsDba6AZtz3s9QL9vN2ysSiMRMJ87d5S/i6g5
lk9wskAH7FI4UtwKAAHsTVaf7YZKD4dL66MUhtSgbqQ3BbQ0QyoMIioccAMJNODU
mSTrXNdkgq30Ku3CohAu2Evow1R3qLwRQjaZ94L3aEXyURzOEPfSoT59ea0zYHM9
NDPWJyjevEGn5RPJ0k1mqR+JYdLkJoXqAFXWkz7qp1tx+hRnhNM1Gq/JS/z/Ly73
SvIiQ6lijh/3aYKBxQXZ/3JeyBGrQB2VBNiQl287vZowjeJYUk9AnqkoAjUhP5d6
lcjtLR7Lin3+ONdoL/V/E8Zf721vrTeSp/0FGwuwRP235Ztmz543sbd9mdQoLJ2R
26sK2zE7zakMXxf97msHdgQ4D6jBSD4AoYNEMT8oE0/kQgJIMTrafNXianWtg9Hq
qK6a+GSYbxVSF+goO6mNWbKqOxeujvw5SrISxjt9SnlPext7fmFV826kS/XaCz3m
c+YyEjDK0dBajNAvCm9lbOxaKQ366DE64sISEaRP9QUWs2QGeQfJAMxTEWdWiRx2
xaq80NeIOAbkP6K92F5meC4Dhp4NtTsddRmzfAe1z21wC6RbVaHiQ3+ObXZjZgCF
22dwmynvGJlbBBDJgcYN02LERRnPZrdFaN2qu7Djca77yRZxVQe/pLK0iFC/bUXx
WrpbHdLsBRLg6oixInrS5iLYcflvINI2h4kIsh4YlLQjxeFvs3iCUPUcU6uqlITh
WzMT1ENBJJULk0OG9k2+xKGWkMWPBVGfbQE3tK0FsjsIP4CwIycVel4Uwub+B6Ib
pyo2dpqQzv4nIBenpUW2SVPMsQheSX8IzcuhzT6nxrrzZuqttNRhoDUv9501a+aZ
Xf/qHZpu+D85iBJtAaEuNegwKh24CQMOds8BblOCGm4NHVQmFousm+o/7ylZqRcY
IsDlgsSfdRzX6Xd4IjV9PYUK4x55Buv/tUfbmcmr7FQy/IEi8eK84h2c+aJYb7VT
uANPAO3lEcoeUp861LxXY/w+vYEvrh8LDj7Kt4QdmAz5zgji3MhieGyD/PWbG0Kr
7QFk7CKLOfLG5/ALt2FLW0LH03QsYet2fWwjmAzMnAw+Xfv7om5J1papw2W8Es34
uu8WCBwWdL5JgrylXlPE5KBi/GBdFtHSc7KBl8vd79rCL3cL2o1VeDTtr4AvqoHx
hc039bbWYfEGlFKCudcsdCTpaW60IbwgvFY7/IIF9Yx1ikxXorstKVqCgdGpOqrk
hPepq8NBtZg+dbOIyQBGsZeU/kHfHtzfLpGUzqAp7ZmE7nEXLCkftPHNI/obEPSr
KxVqjqrtnolNhqXX4G6U+DtqHxrUg49z1ZR+zWghCP3ucGE7ve8x3z4fNUaCdk1j
b3tHuBI3D2dTtNtKGnAP3kLOFg97YErigLLc03h+6SnNAYxZBaElhUgKAILRLvTI
Q/EG5p1i69iuKV4pfMnY8sxpwoynK/97L/8+aNRRQ+PX8+MTu5/vxUjUoLx+Ge91
HQhltAbmt+abyYL9tzhW/7m7k1uPcsXujwqfqJJZfnlRXWuYYEqQcinPUSC4MSTk
VaXaU2DjySM98zuN9bXlYmhNpma68seKIqqtcY33Ewm81PXVXiq77u4O/xJY9mYd
MWLYWG2Xv1q/VsWUT7mkBVmsTbB/8WGCyAjLePvRc01U/DjKR0l5MiChwcSTB2t5
fyeFZKiVbRvJdDSSDw/SH1emVJ6goruGepSSBFIbmLt6zLDv2ux1dnEEi+i6vbTD
iGhJT205KL0wpPa4zl6fwlod5/4ClS8AtQYjUU/X7VYdw2GVnC5rQz2x8WxLx2Dt
t0Isx/rvcNOIJ1Zr9uUpzWQqxTbFSnn6oWwIw0XlPHHq9zJ+dZj3WWrVhRA0x4vM
KwD6PGDA5F1+5/K3JQKR/A/jE4mY06lvMAhokWWXJl726MFZVNbBnNFilZoeizfc
cR9kWn0JLlzklLhZbBSov654GKWJJymF7KgT+DWcmyggXryctYq0XHSg4nWR2KkR
xjV+tO52Cj4MrUPgVozWFHCKGboxOSOuI1KNs6fU0+MNqL3xByRB8Hx/sNWfDa7j
pYPNRE8VybtEJFzAQYLIPSDdidaWDUNaJZS5vg/6RYcs6f/4TCxpj4RbTAhA37Om
kazDVAWVKRjeMdx3sv1R3Ydsmdk1TfYKDwixIMC4DDES8sI3tdiExnShpbCScjHw
NHJgOXfp662kUr94W4oDImISaHB90UQOxE0LiWHeiY+87y+hEDJEa5fPE3nhRMd4
Sd/uwfbkOAS9I8rhYmAQg2bJVIwWXqp8MwV+z5p1aGZI42BfvdjusCypJp4Uz2f8
D3TC2uQHY5hR5l540QaHRjywVlAeGtYrPdvulm/pTGKtfMvkhAXCQ6d1nvRtW7BY
411hy+uitjvEwj/ETEDlymMasho4JDPDTxBS+xvGFPdygvtCfX0Nkh0Q8TeK1CCA
eD/AlEXKmDIKggLG+drhnkafNE2rxsTYK7LeRiGAmJ+WUCBnlHFjlaH/hoxe8Pwl
4X7sb/Z9REEBRMeF7d/STtxsquEsgl1cK7r5LNsqZ9myDMnNzsxwm5W2jta1h1uN
GDc13ev3uLJba+9QAfRpTXIA1/nw9Pjdjo/NLHCnIs0Ufwud0TImTD24wLLOX5vn
IAF2voXb6r6Z42w4Hc5IhlV3INsfd964U4ncY7mNJw9Zj1m4gyGuVEfIZXl716lz
of8ZNmm2HF4ToLMw2KDwf8tiWsBzeoOax1y5xxQfv/kbjZKvN9gHqmgZxz0kmhuA
bJgYTj7f0/3i2YVnIEr6+RU2Bg3j1+HoVKspRlg+YFp+NckRcXmqAycmI3/KeBX8
aadWYEllP6Yv6Xpucp+OFRkNbgeuOr1Xabok8MWVSYP6mw3Rd9KiWIQBvR0CsJ2K
bkJO8SBfQk1Co3V88DdLQQJ7u5nbtWfn9Hj+vQ4ydRD2vW0PhL5jNKR8teugt58R
o5nIKrcqTnxLIUz68sugNu31ZrIuUdYswGEm3bRW2LoWAzWEZ0+RZ2rz08ENrVft
6KcvcXe4uDL8+rvWyO17XTQq/gLqX44QZtu2i0TaS/PtMTk9SFH8rW4nlc6aDdbU
KPoTwt+zttqiAvoZH3Ms9+VggS/TfYIwDXI0bUfvN9u1+ZBMsu0hZ1xAx6BePn9h
GCGLHIO3L6EAcru3iU/dvq7R/eIB/ZQQLubR3D1F3EgfKv/k062799XYeTT2cYng
ucSBLXm3M1sBlpDmDxL+uanetj1cMZxEIjaQyGYAXxENicpeYP15OStcpTk1+CuV
2w1BeIVyUx7eFHS3IqkUYaOE3NtXGhjrOaudBWh2jJicZzpNEWilOOyPajGXna5F
iUMKaiflzglreLBDNUg9Ao/G3nD7LeWk9f1px1Qs8/R2Smv7Hb7fNlP5g81DR5UE
jINRsgGRj9rIx1RmRSyxIRext7K4iakj1FAskLmQ8DnuOVp+ZNsN/HKLmPUu3B3d
X2aIuhw/XJYBurkv5JE6EBqfrMXfRLIj/+is+65u+izlChLiwtTmBnuZAxr/iQUI
sLUZ8FfxcRzO8JzpHwgVFqzdU9a38OnnLO2jfSPhMuFXW911TzauXAsMI/lB3D9u
y1yrjGktim5i+opY9HL3dMpggo0PpZQeMuhXyiSMSOhsiSO2S/eRZMmoAIvPGvqD
eeyEywWqCshM0ebyM2WDhCuUOHogTzLU8h76mCqgiT5BrRiQVAbc136TloZjGXgq
Cf6l5ckpjZVlyFRc5rmEpzGW1EIEuFfAfteJatkG39i8YHtzWu2hoFph/Aaaxl9l
MSCoL1rCgmsp6P7KChlb800l8A0WN8yEp2GqRY7Z76nfsJjJqaTWQiw4FIuYcDj9
DDN8InW7HIOicWPtUpg/MGdorEAktHawnXVwViFOZYQUr0MSwJq5v8lLqSb2VQjJ
e1WWeTvpqB+QPDnfwYOg/vG9DeLfDsMhlL007rhGxM96R3RSKdCSK3clgBVLGv4N
xkrsPCcNjAeOFUSWwBmVrdIUE0kQTPkQ2gXZYUx13TENIm8/Hhr4i5TTAXdMAEw3
+w2vaIUtNioHgjCpFraSE0JgLtVNsd2+xxWwiMf4Vr1yvRfWGEaabqD3DQpe1xGE
Omw+3Rc5g1BkkrMJaT06z5Zc+v2ZqW/xUMFKdH6yPn5ZrFMQCFPKoTQCnYt9UM5q
frGU+x/J3dUiGHsO65GsYjjpZM5Vpm+NsoJLRUe2BiZ+RrdUX9AALErqjwdqH9fy
1c0LtF5N5xodSZg2wqQ/UsGAETEGwNcHGU46GkoO1sUKVkM7ByKTs+L14dIWBeQ0
mv6cSOLU62UhZ7dveHQFwsHZj7prT3OjbAs9rWWUk8uYha8eXfpJNjTzXxB0N6TQ
aYZQOARa7FQwA2g+T0SyHmszy5s5qvF5HvLUq71c2jeHOrYCsCJ+Xz6qTXl5/ggT
OapI6Yx2XCmD+cgkO7Qf0/5M8cWim/TkH5aMUnbtzip10o2N24TKxvVWfzIOsMhx
Vpm1idvNCCh2FieyhtWgmBzPpDK4GDswfljOqY++ELHKLi26dAvuSkVHRAnJf7Ki
ZcMei9mqcDCt95Bb/9s3KKYOcMvib1kUibwp3K/LqfvfZwb3X2zEHBjCgTM4GZkQ
HiJGy/CrwQ5X6dr4BFBFSiR8aXqnzqbzc24xorNugZEd5UlkYJDtqk5wHIqxSwQ3
auJrhR1l9E67+gmaSTD+MFVHS88/2+pbCNAHqTf0SHcnbhT9bKyDfoqD96uJ8KBr
UBljyMAzLzNk4UG2y4eZJsp16Mfgou/JNB1TZ6mi7UYCMLK3XLjgEG6Wlpt/48E1
tyyX/aUfP2rv1OfqLd1EU2TVLQq+nfl4/Zz79K0Frn7eyACGMSaYdSgS2cDv95H0
eNKyELmIErLtDlurX8zm31D0oPXuh2LMAJpNKSTXT/xz4CDM6qd6MLrpdxluEW1b
oqKtNhtRrlwH/VYpqwPuokm+4BAwtvlUMputeUIAB117yFKdUWmlOKCZ/sdqMAC6
SsX8wdAEkvjfHqc08Qf4Vjpfu+BQy0vUh1cfdaBBPGbPpYPFGaYpczdwe6pyo4bj
4phPmlMj05XPz3bzuD/VbAG9GMaCavX6lI4SBlDhrCM+7UZkBOJij9Tau8CxNCym
QTMYU2z8jAc6fHVSx9UjEb1PCPFCbkYGupDsjUPTv6ZCg9ll5IaaE/oxT4nRIIrg
N0TUYg2PFU+3Qh9ZKf9pLUJsjXcDqbXqDgmhvpSFkYjzKfRoyttnXpECV+1f791i
uAsoqVPvSXroAtUVrT5/2fPniGRqO9HQE9LGD4hWfZYlDTxPlndHcYOTV0UQF6LD
14OFDiQq4LF4eVv74Iuk6hyALNTKsSI50VzqaEIzXT12MAffrjToxd9KN97csc3C
4vRh6iuXJg9r7MyIhIlo9p9g19tmF0o1lKoI9Q+48AldJ9NL07XvIiKF8I6mBfUH
C3rhorumO/QEnbYzNGd1B7lD2yZWsOa8+OUkUc5tGIy8X/Xq/lt6w1F+rTBSNhbW
HuedyzT3yjopxKRuRS6UIBj0qR0maQJ5QZ0CTNL7I7spc8M1XT32a11LVEj66gMq
Evnzz5jasWMt/tvcBjCPdEMnYe6Fz61LUx44lAgy/5PdEsr6rM2c9dDe4aV9WAvH
L+BrwI3vh6YEzrg5O4pE3PD7vLS0TReAlZwjsNwJ7jUSQgPMZjW7N58LA1hs9yn2
qzw5+dLUHwUxrMIR1JJAqED7k9F58pjfQ/rckC4JFlKwBJX84jQhvoKng4wi0lF1
jBeiBp0/cBAtNHbm7VusIsVIymBlgDqvhnIJ6L7wU9wAYKoD5Ep8EoQZU3lo9rn0
z048ZNj+gcrXzp0ME52A/cSSghLn/P18XPZUYYsw/cYVigM6daBjTgpZOwqgKPhe
wd0raMsOq12VwdI3t8VA80vCX77vMSnJqQxLgNi6chlJZvvwPFH4GMjpjQD2oXbq
k3Yb5LPeoPh4sbRGX3/OZ02w67HBcZQitR5Bm0HZQ498R4KNEuw28eOXyHSUDLOs
k5GTSpgQWO16lHwm42rmeSIMNvn4FpgW0f2Mbro1LHsla24bwYOSZo5n74BW/MvD
6dBf/N3IDC+xlBZTykjEY/7h5w/T2w5dzWkztcemL2qxyM05s2WJlNgIsygm/v4C
ZQQY8J1YPkdGXJh4KP56yr9Ri8i5NOutKAYbCbj0KLmIM2g1W6RWb8Tptip6v7ev
ev/90gGo0maw+5rUYap6jdUZAxCZ2pmIKfieEps9k1MRSlKuyZu4CwOBjh0MGuga
d1SRN8BIyFUBVavV/hY/0aqbwskJFb51MvRJMZbvJ4VOnom42k2kTs+6xozqqF1v
bc5ys0AVmqXDRsEk+P/OmUVFJNReDU8Inp3kDPL9ypM2+jm7lm5ImHHxG6znrGoP
rr4tj9AhXiYqj8JtBGN2ZZvqCqAIvu7L9x6ki/EU81c35aY62lJ7NNhysps+EOTg
WQFH5xc6BL+XFNv/dgyOFBUDMsy/jxC8JlGCj3xhCHNlwRbyGqRgC593NvyApUBo
6m+0phj1ACSFKOm2012NFyBbP9qQEraC7WDGROn7oiuQ4GxKB8xQ0bmZtGWLVXvf
7blNl6OsPes+m3EPAmGsZHMUlYHW0JXg8nxkXxyOl2+ABYEys9E8ZQhr49BsfN5Q
j0zPzu7gIUiKuJ+gbctgXMcLu7IhQzYewANWmMHwAl4bgiwgGqNA7rdl5Q1wAlfo
1rfEN3LtNbJpbey51xlfUlkhqG5Z3IRoxLfep45mnQhDnjo5Xnk2QMr9gBIUazdE
Rck4ye0j2YNrfvkUp2p5Hd+Rviozlw9uSDFaL11LBvsgH3fEs4nhVF0X36WZok4O
SY26f/g11x7gR2hMJezklN7MfJwcysC4Pht8zsRo4DsO9eLDSfNAQgt5CtA54tXc
c5YZhURCmHaOZq1h6nyxW/g3ZwgWnHbs85naAWWREcSx54Ri1yBCzLjniv6Khzs2
KGGOLid/FM2Sk8NLGqHgchSQJT+WEJ6pmfhX5CkNPgVe0FpYCGGTz4v7wRp59673
ZBbwvkXoV6tD/1iCkNb2DWiqM8SePsG1hn1qq+s4cmHxXVNSl6APbERGnjbRNPXr
HBdT3ZStl21PHaTiCQiOUqzqOoKEbmPd8OcN8LK7qg7CGqVHR5013/0Bx4eGplcE
cFBZ2yiFIF1UmkPuaBlgRKvGzEYhyW0/Wxm7Wk3kTlb+94KJszrzq31eGFtv60da
qEfHX2KNWGsGyuLQFfP9L8HjUE9YHK+GxZbsq5cjCvXAj87LDnm8npn4KHGwqRx+
nPDN7S3oBx2SG58foVcrGRIylFuPdqd588KUPIcyNk6ky8vo5MaZ/vOFY8yIM13Y
0xeIkdoyP6QAR0Cx/sEqJhBdjm/Fm7MwUNy/3XDCrtsH2jyeCxtLhmbdVknA7Uo3
P4/Ex9Q7NhszzmV6SQC6Usb2mxKlxbQhD/h0qdwINUzm5STAlueJZ5nXSkf1VLbs
QmwfrLbXCYjy/SEPPcfUna9CIiFL9PH0LbS01b77G4ZeIlUyVkTsitnQH+ypu6nz
NdZSKqONOoYZO+bo4YyWJnWdeF/lZKqL5pGSv4Lc/wl0/jaBCM9QV0/NneVxjOWx
HJJVpIu7lzcsGMpuRNu7Pr/S4j3t6UdGl7cWn6tHWTxawLpjjvWS3N5ufyi2eoob
MZhX2GahDzEwD9EdjF7qQiUzvowqliprg5zVNL8tHnA87yQS0wVoBHuqJlvAP4UI
GyR19s0Jx179iQkuRttY2vr47YNvewMFOCmR8ovDtK9sUPqNmEZr+42iFgr4x598
QNoaLLNnVcaYdMz/P+7ri1dCB/qBko0kZ1MTbt/6gr4auBXMxEYIHB8AVPBrbTZJ
IWCTx4JwL4jWgzrbZXLgHG7ANbVG2miM0yw61hyLb7vh4Cbb1VyQlON/c/LApX5b
Awu33+LEBaQtd/PkG+LPv12JKa+jc7EMQWkP27DRxUdy6EOMTF4oXcgIta5CqaZ8
TKHlsipn8kUb44nV4WB5enyDTSf797VUnIu/4YeAKjDxzD0RtWc6Wnb+elk4fQgF
n2tUIG5UO6hxlOeCvwIhcwPAGgmVlkeLh4gXdsCgyeQdxOdJ0JlYSRT0bkAo2Ced
RrEWEfPGGZoG/EKnhdbpjyPeFpAJd7V/Vx/t4SmEP26f+mdCwLrF3LgmLry2E88i
tihAPhB52+wo9XCTOcFY4oatNL+/48MyMkCotkYrOA3ND0UUSLwl8UXDKuvK7b64
XslkdCJBxbRGO7hDdL1SCJMGp6bnTVsnij+Li1auHIVndtKhsFDRPzCwKdf30NGJ
hqtC6PVCDVbtgyE5QNOzrvoRy9OqXVGk8ZpZH+72WuXPFuIgcc+1lx9TX1QxnXOl
EF/69jSOD0ja+16/XLGp0zOGCc6VYYCIUJ8DtMjX5KXjNLtc8WdohKcpoHx59S9p
oGQ7DEJ4LoyTmjJkW6o/Gv/leRmiZj50ryaCfLMrW5+0CxGkXmxt1HWRZe65gdwx
yx07FSbBpFZ5+mQbWJ1G0q5wcKCGfKRFwP5LgWA30x16DPrTyyXSvuVJ+s7WYqD5
NJXjmC7cSSAEFVIBb4DcYAzK30P0E5UT3TEoCdIvj0rmLNfonhxD3P+rkaaoYs3K
dZUtMEWzThi07xjPW6hJ265HBxnlQ+vhIQjvcR7bCMl1QWPIRPsP4m/x8/HefMoR
VyJB+bEq8Up4Pqsx3iltL/a//+ujcM2yeL4gCkE/5VLJOU+UZ9YWzeu6A1sz0S26
bIaIMrlpVaqeY4d9CK/FSj0uPBSCfaHcom9onPli2RdM9biTS7SzbbaMh6wkj+I9
ADyYWVT2pY0D11c2dEgl/uBLiQ43FwehSqsfvTp+q2/0ip5O5W1B0O6nt8tXhiUG
pPzN0nYLi/wnGRqhIKivth3Anu7Ogz1oBLPdY1fetm8pXml2u0nULSgahCZVsNBq
kyI/W8y2+HjhN8Kf1v5uNwvAgFI/Hy1qwx3tvI9+G3scWzjbacVzRDoM4Zx+cMzq
rKTKcS1a51jVbGCIASQGgjmVlH3iXaHCNiZpCIFT2wUcXj/d0CEXUABnQf12VBww
FUUzwHjQSPyOoigvJmWg3KxWGy/VzHIhhQ3aMbj38GbE/HB8+1CYTtfbTqTewbnv
XsNGkDJt7Y9nw/86nMDO1Dv4x01IRnbLsbSx/vblwktBjX1D/JlPP1PXoJc5vVlV
z8HzmPYGau1eEqaMBZ+WfwlgMCiQcfGRspLA1rJSU5CvlvVXHHG7K+oQJbVe9u0Z
gaITRmNrF0LoUTdM54X431obgzjjjEOvRjiyN/Lqpd4ODi43YFUYt6km2+X9Msja
MOUn3s7ATZdqW6Ry49vOhKj1PHipSCXcvB0eE5aJiptVAQX+Kyvh2BHjsDeJJT3X
ecsV/nGDCUVJtUx9OMtCRk9DHpEmAvhfS1UI4oco3QB3SpB+XZe2uxQEzWk4odo5
TUpgpoZuXtm5ZKA9BPqOqfAjCULa+IHxxl2cib5Aoawd6y/Hr0g8GIUqAfGEt3aD
FnjeqgGgxJVJikBtrxDp32Hw3OOtwTkC7eVg0iXTFeR5gUQaTl4b/PxdI//20G9K
zq0orKqU6erBgkzcfplda7zyEYPa5v1/MYER/bjBlAj954DYbrZ3ufHcHzqUrEhQ
9MJ2BjBtwPJ4ecQkHemCbWme8IlZfIwM5wFmRnSQHO8cysnQ2vQVyYc/nIIY/hrL
UmsOwrhtS580hHsl7kFPdfCEPbqQ4S45SqtYMUqEcgFQuht7A7Yrs98ksDYvXUaQ
N/1siRkSiRe1VQP88+wodZzNTXTf28Utpzq2FRssyU2vYRQL6fiCUPA0IQUhAxYQ
H1M2p/Gmd9MmZR+5ncHRFsPrS2CB9wR8WedqSo44DJ5hrOihHaLo52glITEppsKn
a/v13gAwSbjC+PgehqPH+OcwrV7eDujqCrCCk08JJg6yZn51l8k5nE2p5q+32e7d
vt5j7Gt+ICtyMOKigDfxyWWB/F5HtVEfCry3sejty3SvwAUCzCe/ha09jJ5K/CNL
1EaEXVNl4rCaS+HD8MFwOhcNdd6h39bGkji8G69qi9Xo5wXS3pGh6y6MjjJlwJS8
lxRMXel3m/LPpp+6N1dLNa2IYawo5rpjD8SXnBNCl606MHWYZCOQzCTrmR6BVn1Q
ciAg1AXNINFBtC0wF+6UwlA+WMceGT7OvyZhA5sRhOCSyDETCsP3msnM3DO5CMn2
dGQqY7/LQgBk1ykpkD3bNgozDFtW1ReTGurXZLKK4gFLZeqTHqAB7IVYPFFswQIo
y9x5cvF1ICiD48FO1vaUcTm3gp4YbaxaK6Hha+Wuq8rTMPVh4uuHdrhExYVYgTtj
ej/QF0UoA55g1yzFWYxv6huj75OeXl1QyeUQGS+Mk7LszBZAMn9QmXZ9meeB1wG7
DNwWlxCYC/edNPwzb9KbnbiZ7KOpgmDDrZwXinQ7D/sIdIN1CChvjMVBheHXuEDq
zCo6tqYiWWQSRkgghkZMeMlYOCVKtpgVy0IOk30iUBfuA4zcAmH6WSv3pm9xVetq
wScHkQYgNhxsE7vRcCS3TC4m5ZNRBOsJoSfvkqGEVijLW934N1eldErW3aSY1hH3
9ahvzMicYt4ZCWz8UIJlc3+JGL0J1D5abNKynE7aLyCkfyDt3oyFjBx6fZwXLxHL
RKxr5JvwAKaEt3jOnQQqUMypLJ9nUYJ6nDWSmZtPhpKV+gH+8RlAoe4OWAnVNtqK
asUcztSMttlx7RMjKI29AGvAusP10Odr/5yVsstKyqCXbgLvEcxYnLNbqMNy9JUm
5fMbDu/KKBEVPQmpU3NX2/Rl9rrKTgkEIie9l9dHbEiZX5LPRr8HbvAlBjGxub7t
/gK1PmV6m7IGsedyMN4EGQpaOLvVpBMl7zzismC2X87u7TJHvU+NssGTF+rNnyD7
xJ/ZWYwmpNsWUmwOz5rv8DSpoZN/FGlYH8O56yGQYkPzNm6iwwsn66weYBZpJrD+
sKCEusM4l5OTkyTNri1GWXo6lrEL1NhdtaSkGfr4DskDCW/i4/CzqpQH5Z/9+5M6
edMOfGt9ReVZkAdq9cf59gh/YR2ZerPyDwXuc/8KKcqI1VnsP5/xuyXSQqVg1xz0
fESw0Js0sb8s2heJv9++xWNUn45gI7YUc5orRIbn/TE4suu1xK/YA/IBTbsIu55N
P9e4dIXhnIm97ogwX/p2HD2zJVxQfZtJ/UTtratVPMgrW1N8nC4U9dKhncSSTJQu
+oVk90DY1ki0okjJRmIdhEQpts/0P4ZajsXbMhiBpTBzJzPDFTqHI+qfDWQgfAdv
HKu5kY+B/Jg/J3E5uE/xLio/8O1ycPdH1x/6y4CkENksdw/Aoxw3lPcv32IEOlt4
fnDwQ6LTpffb0lge70Cyj+4EfnXk34aj8TI6MIVAXiHxX9c9X0OMXzMFEvC+KF2C
JiknLqT4lXa7S1zV++IyIcZMvT5ZpzKp8AWuE9EzEswYTNxO4ooGgvzgvjcie1d3
6NOrCkf6MT6uyh2NroEpEXlcvlP5ZUB1XKDT5CayJb0hVJVYVi0uxIZI4KN7AIQ0
bSHh0TR5o7UzgUNdkQzEVDaUOoBOR0hOx7PB5aa0TyILrcvvC6HF1DZYB7Mcf2C4
djXM4jKKtLLIiQgYCUQwynXyI5VIj71az0xSX1eM0JqUUlaPtNriuoiWCvgdqE2z
jm/2BV8YYdTn9do9l+/145yNJtwCNjDvLHlh6woQTcOexT3rebF8ercacYJ+uqy+
yg4BSb2kVz2ljS+S2VcIb9pkB2NBQOA5KmDNoOwKPT9dI/VRYtwLM3x5rmIoBEt6
c5clLs7vy6mq1v/LY3h2IwmiQ9fbZWAJdHdcjOW/aMH9PEdBL3xNbt2k2JaWIWAl
DNEWc4+OUDN/KUYbB2zLsF9FV3Lkv2XI/a+tnIalRMYNYQvAi5cbqlv031jsST8B
d/3PyvPdnD0ShrDr0yN8Z9fT7AK4pU0DkZtd5wEe6U8N8a020TYCsbdStnbuUx+3
PoU69ZxjxF5Uxk3zklauUFnmiQr+XfJfdXKWUie6kYAk8Uk5/eoDRDxUMY4+M/Gn
OWY7FQ194HENb2MIjqggNZigH2hjSvVylaEC1gZOeCAuQ2qdV2RYIoLSnVncW0BC
oYF4GhPGTewOAKVfop53yjPgSYrxTegQPtJtRfi/X9K+1kfCk0qdUzSouFMwkiHD
gHWqrD4vyMP+k13e35Q/NLsflha5edwBwUj2Ih+zYlmnIOnw5NlSe98MeFexq0eL
mY3Zdcxyc7J64QKwnCwKk0cjdurcxvSXjWrvESdhCme48czLt1W0NKYC4dLPwu95
uX9jSIMnzJgTSGXimD+dDN1pIdIdVdiCAZf/tVA5MZ8EoraXulp/xybbPZbbZa77
lEX/BltKY3ecLN8/xA1toM5chBRacpMGD86Fey+f0fIWGtntMo3+kNZtqHPcfWbB
1rfODCSO34FJPlAEl+8u86NYTG7BfCPwItDmxe0/6SvwlqhcFFFv/rZ/CcXNP4yA
DCJ1XgCjibMexNAlVd1bFITY/b96jh7hasifhwrir8hOXFQRLNeXKoPrPBZG9ndJ
/TMf0UQ66lYTxZ488liFt1y8h1ekapUDk/IkdPS/2pocS/f188WLoEvGIVn4+2Kh
viraB73DlG+i5dR922hvKdeEXuphAw81k3VJOtdBCB4li/UEtUD0s0aAw9Z6bcmu
628iz1u3B11HtYIgru7Ky9G0f5ZBS/cTYuJDPYUlDs6WYHS0UQq2fh+dfYk2aH8s
1oGBmUL5CU8bbJ5aIyXWKB728sQmwyR7lAXa1fA9RnWzy4qeEAjiYpoFfOv52sQA
N5dahYoRTTspZ7JDHCC4ueULu5nbjP+/h24CUFxkelnuDSCJRQpYUe/YfRuCeK/6
I+4kyCz2Q9995VyOaYKMeS4aAuL+a9YoArvKdCbwuE+TgoCsQIXNKu3bVO6ZSO9R
gDEin5aD515+oYWsrPEvoVp56/VgvDWeToPiUl2WkTv8eMdRhk/7PgoVNtX/0DvS
QlH51ipiWuEPv6+BS4z3s9L9T6HuyKzgQ5TkA7kIu9xaiXhHUCm5KhVJREItSzxR
utdCts5OdGPtoXXhoS4uuDWBLi8fRKNXQLuPrJV/LOvjcHeQNdc9K3Kge0KcoeSX
T9YeF/7ZOBXtE5J8C4PDt0918ASuncRqkeg7jkvF+dOJ+UioJ0Q9quPMfPQAjtSM
NEsRBew9ln8sr1wln43Xkn+gI9SIhLW+D19pt8nAIKjRMhCX3VmsLr1MPPNsWKV5
xE5ol+XMyZnjU1tnVSwE+y8ftnMaeYRKybWAX/mtimEpEceqKI1cXji9RsaE3ZS5
yIaxe6AgwLxJD40UNZuw5J4YFF3qBC12OTdtdk2KNj6T02gwJ6qdMB09azKMKv3Z
SuXmFsrAZVsRkM5DQc7ytM5uwhRzkU5+70epiLvgkStxKj485Ps+zn9FGjE+L8vn
zIG37A7V99wLfiK9j9He9DN1ZfqiymBLgHBUKhF08G9ShkOLEej31BziJJpaVInL
RhlwDnrr6U46rlIDYip3o5SGL3jR+RqH+UwbgW20B63BLY8v2xXiIpwozWp8TMjI
7CBaw85BkwwUpLd/2DyuyuHYhb/hnWIyL+w+3PGjSC6zIcDe3EFof7dkQnCiW+9h
sTjxBRXUVt0xU2N6ucV9sozFN/294Su8+Cl2z3Koqp1/QwJ2ZVoRm2IzTpD+FIvo
8ylBlbPA+Or4m5RNtXT8/k7ZzOiJmW3OGImWE1kuXvu4f9J+4zCT11CJ1EdNMRKv
EPIxMauYSY5sSFfZWW7OvXzW5UqnM9ZTu+8cmgf7PC/b4lgXrfZHg3o/cYYoPg2H
aM8gf1ggY391Ljgmx3l30lsUbOabZ22So7bs8XbSBtBHC49VOtU9DlCnb7sUyK1f
n6eAUKoN/0JYfxttTo1d7G7il6A/EopA2lz6mnEfFgbO4OJ3Z7uH5h+3ROW4wepi
ePTsjKR37RhPU7c7cAaULmNaFl2V/lPB6Rd2V0cKvLKTQXwF9zGNUnL7nd09drL9
bYwxdEFWxph9YBi1fPA1fT83G1g3SOwIgazQcHaQUZxcXHYIoxcdgqQ/9C9PKUWb
k2Cogreh/R0pWwQPI6IKHz7+oTtu8BiKjxt4SJi93VB6kGhK4xEnNDrS8UKBT5MD
91yIkRfHuB6wTnETdbnv4/yRQJIXn/1y/TwJE/+Z/kYemYCnJDxT05VwjV5fxB9J
/jfW/kXN2dGUhMP9YtjP2HFpnIopAugDUMjONxdjk6y6rcY8whuAbbKvYlAMwEwR
6NzuKrgEzL/BkC3YaOkcHDCytviSnxEqRvmrO+TnvMuyQSyRXUvgKGiYKJ+T4Ou+
Q267COT2XZUJiaPApr98Tm81jSsRVfo7rfuBIiVYppGknqmoQfXLmzvgGvnq3kYP
fH99/WwXuhNXtyPTkUdPTHMQXCgn3uCNL6t9RHxUNkmfoCr3zflT0y0fh7cS70L5
jwT0HDSTbXkEvZI+YCOcDAKdj/EUV7+wr0s3ornCxMRR8L3WBKaauHKkEgmN22gA
DZO6AYu54o3xoC/EFsy1P825LJ+OIG0QJarVD5XphnIIq+iAfIKfuHIyY1Mlq02D
hHFPGffPFRPPEnDBCzLE28o2btPUKqX2E0uk0Jrh2StdteBB4oLZyeVXL9iJ1h3a
ZIoCW84oy1LRi4wT0GniIk9u9T2p9l36EceLGmixXt3HowgTAFfhlfE81yrinp0e
TQ9fZuqoWOKogAz+hMh+qb8G2T6KQQZe+7QEOW4YudribKuCY+74NxtvlAYvvCKv
RkZdwSCW32MG2dI2tgOM/znBkoXirVfoOzmMDDeTxVSOS7V77F4IwiOLn5dbG14o
+Tpa2RbhxGEci4d0Egp21NpPRnL4eeunXuWVjM5mFDQrFPL6Srdc4Myb04IRQYfZ
Ot7PRB4vg2WNLbqrAXIR+clFocc5Y0Sk5DwK4KiL3NulkGvJMcZjt0IccBIC4pma
QcEHwbJxDG8Zi4AzAFXsD/2+HriNQBMIXRhAq6MqRMmbXL1VNIMRLRCfvK3fSbnQ
hcLZqNIulISbwn0mFmECwNZ3f+nzD+GbuCEKNTp2P1eBicHBTusdk3RyodoDSEbk
yf9CYwumwSycSowxEoxnv0UQqVR1Tl7REugksi7GZthDXu4PK8bkfejF9HyZKbVN
s+RrNqbKWYWkx/9XA/YvPZBsD08OF38Dd+LLHdGeDbGg+ytqMb8sKDaNMS4PsP6Z
dueu+Cggb0VJ1c8KLvZp0lAN3Z9dHmsKDDHYlwpLpF2GLsheaThTB/BvwQEMFGPh
JD6h88M9YPxyCzJPI/BAkzZOtAsGVmSvVYZCvLKMxWhMgvLsIoriD1QL2T8F/4lW
EgsShy4yBUgRb0CeLLJF7uI4xIslwtehWKDcU/WUf+jAkZW1ClFUyKy83I47hqWo
aHgMnAeCfitjlAnXfsY0r4uBtjlAhgtjYE5WF3fEKX5oe7RnreggtNLqox7YuzoM
7CPH0Gb75cewN6Z+0dVghSxru1oaNXnpl6rm3/h548J9BEwT+P46d6l/1uANyYum
xO0lxNV9Iae4BXb5JQ6vbKP2uNaBUgp07GsN6/u04M4+cUV9oeYFF1Lp2MFiQs4R
vc3PZZEjqh/ZsU51ItmZVOhZoB5O7f5jCho8KN096f5rFtm6x/QocMpiwJa3joIx
iO/FmYasJhUC92/GbwMrxgPXo9tMofucJ3mACLtnLvjR13gHmdP6hKjMhFVtlz4Q
tZu/UcoAzGHSvisamQfsUfE+Ra+YeAttJQHNErjJ946RAChXZ5ZK1V5tyB9W+Cuw
IKLG2zaZF93zMlAhPWgOCbu6NI5tm9KfGksloWnDeEzql/JHpokf+N0uSPYbibim
c3u7CfC7R9RCavyy4w/+1XfrJbyHCXMRrUcJN1AJab8Oc3Paic2CI8Br729U1dXo
T+jhQA3gxxZL4VrAx+SevvampfYGwrIvSIr+pAoTLwnrukgOZ6ELphUonbLvoObk
a8KezAw5J+STKl3xmyZNSP+UwxX+oqjjQTnXo8CKhySJrCVRkcevORhUjjva5iRZ
nuY60DS2WHYMVxodXBwvgz2nUtGxOjSus32fKRrql58Z0lQsEuWX+l/g6Z3af8Gz
wIhEtxbajM/eKJ6j3qc2wyGjNHZ9wHP+55sma5FE0UutjmyNsewHSta5W0Fr8dNi
McGNJqqSPVrfx5P0S6EX+9qCTJVAXWle+RX85+jgnx1wbLx0Yp0jDxO/V8ZgVCS4
J2SyRFAicOXxLNW3305s6BStuPu5NPr/ujRIkpO4pBVmpsojkinr2J5JF/dZ7Bix
1dk5nR3EOymjTqkN8kpM2zgzYelSZzsvTczsr+Ml65j8bLU2FIIahRLPowMIhnvW
CdwcUizIjyiPL+5s+t3QLE9m/aN8yoHKnBTtL0uFk69M/bzH8UGZ93lGS9UeT0ls
454XOj7cA1k9SInVIMdcSt9mL62g2Log3WjzEPxTonx9XppYfG2FbR12vEXaik7M
HhX8in3eb6HmyXMmEF7sa8dpmFAVxhtlRuhaf1uS+Yx5Du4jEXrCvRXVF395UYb+
ejgtsiSKUPEiMeNKeQVAO8qw/eJ++49cVeCLfxTxGmVBFPHwAr9kjDxPKHx7vt42
e1CGByCI9R0TBoClLOGFGsQ1t0TfBqwBUyqok34z98LWkS4wAESJ9Ufv8CDizyI5
XXZq1rnYEPi6Sg4sAOLFDunPJgW2sZJDMTN0ycLg8mb+VYORqJkDtgB2pjtuI6DO
0l86GE+ojLGcNPvouWNcXK57rDcRMC1ZVl5+jeIwTXXgnd9F/3L5/su4Sf5OpG85
LVQwNQHg+aQstydTd4k/R+RTcJ88+mF1bU8WzmsO4vWLfg+BB8IUs6tcwPfIuZ2X
fTyLcqyp/tuEGEJxBPVl2ifw+Zl5+gq+wIuXbH/kC+sFyx8INlyb56OnfwJZBCMn
arQ7CNnWcTDU+rPCKmRq8XY2707AdTqwN+thowcst8mIIY+G47kVaXCY0gi2ixUB
njNGozpQRtbNMyjmBb3GJzFuwAErVQmyINo/vZvbNI6a5tYsNV/bz4jz0hLbOMQ+
D7+AyHE8hR/8YPHEOAMYjvklYPFGpUbp/gOruVH80+S5usNbG47jP+028Dma7Bq3
XRI8r9bSWrO3cbeXw/S9tUxC42IzN2vtaBLTpCaybLinxymUxnnBz4sPbdDYvwC1
Thta78y+/PolXMAT13HNatpyvkCssWoZfvKAClKbux2w3xSWMuWuyY6XiXJWt9y7
DgoYoklzR0ehR8U1jkSS/VXlfVUq/ApM5a1BBmW3MI6qCZPlnWpRIQmxcw2FcJpF
JdiZHNLDw7YdAtzPlV8nbyDQenObVGb0I0VXulDRHMPjZTffFA94L61m0A19JswJ
GVFpOnEyvX0UkKiS3PXDkmw/Yhlo1RW537bjS/UCDzTJA1UuuGJJBHFW+zt+Sjyg
jWK9fK0Mj1MukwLdMJd/pKyU5truVNM+JwQ6wN/8bMt2W7S27Ob52OA10oW/o7Zd
v+vM3QLqbikG0/ZNFzngP5VLW3TM0+DtlRbf3hJCagECN1cs/RcJkOy9Z9SD6qPa
sCIcPpkIEBtfc7Qc+U7bcycW19aOW9vmp2yMso5VY4M+ltpCECctLMug6/5ATngF
LRltxaLbeSOujKnxyN5TTM5Nl3HOwxQWr86rqGG+20AcQnUpAXHRLB/CqQvF8CqP
RVQIYFFAysNbBpR9y8RwQeAl7hnYdqXG32V1DMeC20qX8q6pTPLlzJcThSATWRQ3
ivJk0aRkAL+EXuM18BSG+/2174KKW98qSWJVbdfFIHYsKa6q8E13x8327wURyK3O
TIDhzL85LUUdSI/0dKHy9pFqpcPn+Z4s0Hw+7LGthH1AuyXHE8ZNkVShfo17KcmK
5Fdkah6+ApOTb3yNe/AdH1v8si31Lfk+nMqyf4+kOtVOiOQhv0byGD8sTDX990Q1
8+znraugXYFpEvOe+6BfrnjeHn2zt7St7s9SHE8uDIs7T93zi8/Ut7NNWg7JcQx2
cM1rZmqPooha389KZ96EJYCmfml29f955qloQPk9gO2X5Exo0KJzHJDZKQ625hor
CDDL5urZBEXtp/OeVAGLxH/XMvk8TQpmLL6MJeSJL+uNR81wsce3cNlEaknnREKE
ALYDVhxv20gz8YT25CDeMG48yx3p5nDMaGqRUc6MOkQSnh74kJiGVP7fQsaQaS0R
X9pHEsKIJt3A2QGcisb7DdwSL97SqGnTVRkuH6TcT1xsAgUsiSx6SvP14JWj3TjW
EJY1ha3oYOep/NF0forctWGJ8nsjFkakeT0TXkl2sKC3nvZqbjoDXy5vHw8cMJz0
NbneWhXU/Rca7hfCITCKPbF+fidcMq0uMqetwQ9e69jwQ2I5PsfE0JP4kG0ClUGc
BoRlshqx1HbD8BzTAPQLMQGvLcKG3HcO+PQM0Yqm0GcAk2fsJ/bEQs0Rts1XwO0Y
eKkJ7xHEodw4N+PdxhLS6rfcVLosi03Vm1aB7ujzWZ389Ah+o6F3x5jqauGMWE6H
Y0KUtQb5Q7a8Q//Z1vJHdkyD1HHwRN7l8QG6YagRdoBQS5MVMpkYXfdqVQqiL4Qy
+I74agG6Ebw4wYLkT3JfKna2gylSIalNavfYKweQXfMtuFrFwiNvjNTI/1fQwV8m
eHXTnV6bWLWHRucq5009LY3HkXIt9xbuuXISbpg7WL4u40lBMalT65P3oavUpTIX
jk+6aUyhRMwS1IaNkJ4O/ufB56aG8GpQg3lVw5dGSqc/gBh5GjxO/dRD0RLKN3Z4
nvGsDHzFYVx8lr/p4WtbYAVCM4cSJD+2swdPgD7v4XvjZ5bip1MDomiSr32xWrHS
EMZS5CvUjkuu3Zh0oV9rjMeQIWNudNohRTymage5b/WN+Z8rBgw8v2LcEwiCsiHp
oLgcwfD2g+9t3GFEmUt3+aWa9y/G8DIzg65hxc3AMc32z86I8OpekKZF3gStI4t5
VNQ4MfVd+a2as48e3JhrS0oV8yk0DNgOzqf90i4ZNYBmktIwOi38m7DTTPNsYDZJ
pcHVVpN90nAlFLx1F8AY7remxykP66GTbiUXsXDw8fL7dGfab0gHJ3frsdUfIpw2
2Ap5uwwQeLSpJhDS4/yQZgN+b3nq6UlM0DNYv1Rpz5u2O241uuJatTnkFD5ZV59q
MQDYnlKdiPbaliasb0dmGPmBP+y1FGoyoH1EtvGVUL58KUMqlOPoiZakWePHl2/0
7csQBiznvjfNwCWEHrkDK2tz+Bl4JazBeMUCyO986qS05dcsN929XsriFrTSvqzh
WWVTP6fHtoPdu5LT2ffcU1RhgEfP13NlOxcNrVYGefPMsgEbMUBP8uaPxQt2p395
5G/0hqHmJUVgYsNNt+lk9hy6U12mQjHcCutL30Vu4Vyu68+llfD0OmNG3V2jsCah
K9d5oeJmN2pSUmEQJB9dbrlt0hYiXi/OJHT+XuARUBk31gc5LZMbLL3ESIzDVyk4
2yKG9jeYC+xDnUBDeTgnY8qQ2pvwenfqfzHwur7M/KhKbjUe6lgNE6JjZ7GHrmLt
g5vfhGgp4Mi9Z6zOwqUc17TabQyiRNb46GJtp9BOvXwNdp/GnAvZ3wQi7XnPljhY
/0Yg73K/rKUEcdsnkdG65FaJ23+BzGvO3C/CmUFJFtJ5TAjR3yeioIC5o2hTZste
6cf2wSIgqEzfdgs5G/C/Or8NgVQZTSwQq/DV94NFAL75QCnh0iJCsOBcn8IddNbn
wdah+woggeUu1yUy4xYNlJYzFvMOR3AtkDAgUWBbB6kn2uGsNBJTMox1xkH3NQCK
nDzGr8C85SdKRTmgOa8E9IoEqkAvb4x0Zf557Cme3TFC/nUhsRQ7pMjrrZQgnPmB
MhhVEKjYzSia8zQmGV5H6o2BOEf49IHWB18Qh09cHYLVT5OV7O7h15FXqj8fPF/G
3Am5CfFjGbQUx8IAR+4CT5coiDkohAEGgCpIAvzYFOdJUuhSzxS1xsfcMypbYcTo
Up2fFETBPy3JB5VPmh/KqfJjDTg0BtWZXeBvVMmpwWgRKeCdgUXMXb+CL4+Prqq/
Iz5UCOHRTTlo4pka8fzZ10P/Um54dG0QRp3YwHhnQP7lVdr9sZ0WisJ8iCngd2yo
Xpj6LkD0TGWCo7xGpt+7CAH8yZC2UtHrnQ4GE8gSxEu7JMx0jLLqUAoJUQcUUzBf
3pY+Nh9s7HIxHLcM4jUR9c0rOla772uhUWNwPYrM2aIbFiD9gNuwSJiA4ElRHkjS
9ArsVKVjpkH+1EVWkDrxqvEN9iRrETWQwNSZpbCw6DWqpTekWxy9If08OjaoPvu4
w1U5wBrRu4LIc8ypNxxYFLiQE4enFXDBahC4yoT0ptf7xP2nQckM+2ljzAvGagSW
/IuE0tKn7Kydry39YK/I9t8Sn9lPKT4aGPVvm3GaFMXcrn0Ym4HnUMFCDYrm3ajJ
bd6IuRCnlVpZQs7rp1kOr/bXrbtocRE55I2RusB4N8cBR0mGdBdCKhe0aVQ7P0A5
fjcLOvZ95NRE1xjfOiPB4M/B68tUDi/KHjGJw/xmMkR7Fk3v9XyNj+nz1KYlWPof
jlnlzSGgna3THSJEjj5ZXI2EK+j3XySXraNVZIEaEnW6eAO8EDpJ4TS5GfKztkoq
vfEDvcT3bfqjo9UlXfjC9YnkGyznAqQCyYzAbSxki7QP1yyVnSdd4TaCFmuYgrQW
dD+s2giQLGh26uXTQGDnaBRpnBnM/ntKJbrFbYXufAF81aXpRJZjMNBAqJh6mxs4
jxudq7Mm696o6ByglLKy1nksF7f6OIG5PTcVWLDh4O7dJWZf8DPqlrKL2Ht46R5s
c2qrhjcKRrbUNs5FvKorFf/W/KT3xaurQKMKd17B2Txj1MVWem5HncWYoohugzyj
1Zj6kRkta36V8ur458nC07VKaRxoMmOyZYJmgiTH/0BLgjq598Cy7wGJE1uJeU0R
RUY5+JiAw/1sybBGs/kF3myYxu+lvRG+a8d3qXU+kHas7KfDnvRj6BHlo0B5q2Pq
pabh1y4Nalpwl6MYegpU/IW3kzYD0L9IsaxKFIWcYNPP9MAtoVeADVD6WzIiUyVD
wfNt6WH7z2CZdEu34fUdHX9oBWiqiwmJPKIm4+FAJrF55xWFk0rpNO5PSVIMjUem
CjoUejzrsOK5WTnsBnBbmNiS6ppm1TJx1rwexVagdcey+R2ONcRFHjb6icM8qQMG
b3E0PI7fIb6H6ATEm7rjP6d/WbdWHo31Mv7zrVa38lobLXTHKpTOCJUwKTJJjYwy
FYaxI6nwU7dofIa+abka3SMBnvQqdhzhpEn/wXHqombktQ48gEpIS5JDOHOH807v
W14AoJmaDIEGzOenPruJAKeR1aaHeGE6TEfUS3YFRh8F67I4M7TOUy+AnGJ2xLMW
YV0N85QtqHrXT2Ls8STpVQ9nhtajk0tyBjqp/ZGN9XVVKVPeu1hko2rt9I+Et7V5
64Mwvc8MaeKd5Hz9IwzcUNCMYSJo9IowiRxWeX1lRUAKReHT7s8uBNTm7tADTm6X
4toieezzJmur3RYVpjGBMgtx2u5yImNpfGuElvpuE7yamHpxo1zN1tbfU1rzSnkF
rjVyygf0CKoLEsKj26E3s86zat2jziRZj8xcn2mF+dHbcWrbL9NcnDd5LSbpWg8y
ECVRc0IUfuDxBqrBTpQrX1YYeuLSFhrPkNwDLyqDk4J4T2HUly/NDVeWvLZ4aAQs
ZPexgonFVTOQjkayaUPb7OKuMqsgUQMcaDJnODJS0zl2IFDM7ziSR3zRCU6rABY1
BEuFE3IFVCPATNcJrf06CQ2nNrr0oo8LUriPLBydVwrvMnqV0+jppvIkCROb4DRi
OECMGZIl1G3WsiiufxgPnr9lWP43nPzx0LV++F9yYQZiFifVzodhjj0AQ+q64z2A
xdVTPoZ81AJzsz4BVjhszYnQNn6n0r17QTV478bX4ePaNdrXsTrPqM32KhDQ473p
+Q/y1TGlOUd1CjiO7YMBDDEhXFpWMv0IAdDlo33LKquoXcD2oIUu/W7kNKDdOzLg
+AdlyuUB7JjrH1eZqFsVZh0AfK1eD4xacwmwbiw4LJI/kL0o2IkrZ88NvUMDVSPi
z0s8vI4DNnsYhRTmMV2tkAV2dVqzsYQA1GUDZ9IAZUYBBM4BBaPD+T/JVPP4N7Mx
UVDqF+lj3HS3b0ctJlFZMmIinmEAOP9aVcTDOko6Ng3umZ3X3FLQrvRyOIiJZ0yA
2pZY2dR1G/f/0jYFeOA1AuGHWTdoEk+wQaQsnKOn/z0Gjh2gDRFEalfOOwsuEL5e
p5II/24+FVvJgf0aKQfgt2qy0dhCtsP5Lmmc94OJWKCsrUEMNzbwZFKw4/5E+yqL
H4ddZaz15KpnZ3fw1Th+BR9LytaAYDDcTjuzQlDJ31SWAj/md+oDWAvYEbuqtIPw
1cM0S1je9K6zJIhKYYoEzE5KxlGJ5iU6zbMM1O657jNmb7ZB57GnlNjNgGy2MIPm
uac1De2xIZm6523b6wNp7HGk60Dhx+zmr5Jko9/IMd3xiOzhbNhJe9P2b97X9ANT
xPBbbU4xWL1fTAqHZQc8sCkd1aAsmJDHjbEBvdKoapU0KkkqFTI18wLMwa38VL2K
ybKA58tsBxwMrxEJh3i97d6GMHx1q5X8VFSSZbyUNBFfUTE9b6DubVa9ZML0CYiZ
WBVMtF7JjqjGWyHs8o1Q9V0Hple5L3pqVPRsMCT0chOng/iwFGr2yg1PJtO32oCJ
D3XEZw9SCZV+15QNGAclslEHrwLAYFuzzQTebtPbFBJdtPl3W3OvD87NkGIfSe5e
D4zULPfNlqLN45O4aAfh7YhLdhbgoVcUswYHjoeN8OpaHAuX574F8bXhqmBCOuLt
YPD/5hcfOILYCSUb/U11lBhjTGkJqrz3Ql3YGm3QLPlawbgxvcHAZfuxFnrvJWN2
9OcCzxomAQEg2qZCv7YHB3A1XHa8LRy9fE6kCrWXwCrFGdMy33zNvs3B4qp9Um8u
6ltOLTxdxva6zeKG+8WhuPcTSzX8TpcV4j5vmJQs0D4fnYQL29tBWvtogajH31Qt
9pV8Steqm6+tgP/GllS+hy8AeZfi7+jkKaLx3U4tnlwi5nYvQBNDDEqY7qJ8byun
DcDxtaVHOnc647IywkZyKz7EmszAWN1vv9lG4e1DlObVwMQiuS6eelMqUYiYBkYb
IvFFzsdRT6k9aEtLKxJRc3b3s80UQul22+KRJE/0ezzK0VtjjMm+7Z7pSFWUmn/g
0o+36L5+Jn/uJgHOzEflRYRVypalOEWqoK4NfbHZolzeX8BQwQ5ww+CIiQK/oVxa
dYS8im9230usGzgAR1tWrucsm/FbmMP+A/AMn86DYYTEdBaTsB8wcReukmVz2Oj4
nnY3um5e/Cailj1BAVpraoFCmqswH4ELaxx/mQ79N/JbLeV3L3PP5QUCmfCcwZAT
W7vib0h2ygz18OU3b8ulhptMy0O+gnlKJAM3VzbLH+utdjkZXYGgImxBFwImOWl0
Z1DXsxDe3rxW6dgmPDherlbCk28PjqFZ6pH5SyKVtvup+TF4RZC/vtdoWVqfOvfE
Kg8xmulRswc1ShtNP4gs9PTiDsbXKjfeEZmgvSo6HBJJLpG4wn4AXTIL0UBvuTwp
9/nhqpDRiQ9MxeyG+Cta+WXRGymTC1oX8Uew48RJRGUMW9bBLK0bKHM7sD+IZgFM
aLin36gZh97GW1rbeYEF1BsvZvYumEQsPg73YWYieDsZBNoRoV/3lTi8CtKIBAyx
Fjpor8ZNyafFXClZFxJKn7GUJn/U5nBYLEiXJkHQUYAFKUSwVKI1WGUH3fPaW69N
/ofs48TlMUgcaSF9G3AF8kLz65KJ9GheIIKZidqGcl/9yzRKY8sFTUUZNCBJhqEn
48sOkam0G3pUCrZYfwjBdBJmsP0kb9z1cZq0U3Zl3xlvprzJYl2GDy5WfDZSBOFg
87EMz6sxHzt8/RBgaRO1liHzS64NjzlHOrhE3nycWYKyAUnsHIgLDNunvxLF4OiM
bDICiAfFwXFK4VQq8wrW87SbAJj6pO5ZXDRdmXY8HWZv/n8PiT/lWK/eYA7zo2B/
CdlRujqdL5nkACNMR0bMkUKnC9jJCWsAcOrQZQXg/yYns9ubTq4lG/ukuY9k6eqc
0ldZ+ONzKRDSS65AhtLh+uYdbxxyWRu+T26ZFoUwtWu2bBeFu1vlvrV8pLz++BfT
apeuOqKhCs15CrIS4NEjGgAO2IAdz8SvnkYocF73FLxQ6o6cM+WyHQzPMlcjkSp2
xvNOq4xbf/N2ymLJOY+6nsrjb47I5gw82IMXFzA2rl5yXm6J6iQD7TTkV3BuUf7t
CLdFZ9O5D56yjFj/aFXHxmpPo2ZdndsD20NNnQKaWwP4Wgx5hog0aZiDjZ73WdJi
X6gX/qXNtGx8+MlEkCGgr9iHCWxn/Mur5F4bVS6s9SA4keCsdB0xhMziJP2tAU7o
7qcAf5Hh8woWeirw1AWbbmUp5ZjhXYkF1t3m6nIZEUfAZW9B6lpAGyoV2o+yBWaZ
wo8T75i3+KMSZvs35Zi/ea7LQJXTNjwI1R00CdVK19H98iFO5YZDCKEDiRJPl77q
NjND33F5LXaGmEKAf7zlr+sJ5Tlp9ZTy5LE6iKfxgF9rxgryhzPNHttKE3nw14xq
5qEspnnh+tL7hGDnJncTkmqDmkFGc8mMY2Vn7ercBeH2EPcE84JzOSY+94SUg3Cj
qbtVMchOnFCBE5zS72F0DZtylLqoE+PMrE18BY8tYm+xfhv94IvRxME/iKDikf5l
9C7Csmp3ZSs7C1pocbWknpuleZe1r/L196X4T/pqoxSUIfYWniq5XTglyo04du2j
ESpavORxuPKuZkvSlparbzrQfxjVOFwpvH0rrmgxEgB1kZY9UhfgwPKCCjBBJH0N
3jSWleyO2UrwWhDgjdaTlIsMsl1NOgO+5NsMMzU0UgCPXcOjzznyB67wwaAzGl+8
sbtfzxvudE8+nlW94O64xK7VgJbs//3PTUf6z5LZKqPkGxmFFFPMC3u5DpBnb4b4
MnnsCiyAVX6YcrSsXMlYLoSEzgbBxDHww+/o88qxWGSrTzxZXPHCEb6xWhz00pl7
RULkd+eSX2trHw9xkmYhx09wudeMjwr9mDsBYvfxiZrGd3/jkG/gehNrMdJ4Wcwr
CvqsDzYF0L2xgQnUqXZASCf24YIOcZ3Hj9GZmcuMVTCJ5FyREbIPLh9mDBybo96U
1bO1kCXM5iBy2/nVEljGevwWV4U1Cao2ojqg1hJFy4HPtmPboFGsJXcSaB31UCn8
e7chiwpg1pPhenTO6+TsrngyBHMxNMAsXRyJG1l67arX4MQ3H8GlVBz8HoEwNwUQ
O9HGeziwV+7KXojHFjfPatUD2cwS8zNJ4EssTxDW1LZ06cL4dmBNax09EOnx9C8D
e/feilqrt1fgAETNQeC8qc/0+Xk8PiQnV4+eelwFyZ3xEYPaxnNPyxqNtR+X9VPu
A0tCm+Jv0zXpX0sfmeQeDX0dkaLPECipI/YIFavbLpIkVxU2PW1nmz+c+klrSNxI
7ELXs2qzEQXnlZiSMpvRk+Kwkc7mqYXaPmQ94dSHbIN8HWS2V5Vyzk1KS+4P0cyC
aQdvgGOkUsMuu+UsmfNqS5vGiPDzruI4vT1XpHMdtzxqxnUc4u5lEoHhCw/MlE4T
YN7vE39mQojcUSjW2MawtSWWW3EFREM4bt+jtovBYP5D8g/M6UyskSXNLSaIszEO
j9NVjCrS4pAGT8uyxJTIVi4n64lVNp4MGNDxsVtr7rs6JYpQqETcnYE7RNwVh9yd
ZuLL8/TzZs0Y8tVrO1hPOvDaJ+d8p2Y7wzbi+ADUpGIEDUy1JEObyJ3PcM/UrlU/
INVw/d5Nr1bQ1vY+J75nIv09ZVAPIsRwQTMpJybc+J9KC0AGdV3NPaKO7G/v0v+/
yAYUXGRIiVmqsRdgwfAe3OxdDeIRURDeKhLpcmiQ8+ZEqLZmSx4uo/F8Hph4G0+p
lvZjTb47CduNi1m629hobfK9ztEMxm52ctpAN7xEENItyeVBfbkOOFqXmr/sNf9k
5GHQ7dk2ENCJ+Dac+Buaf9+VMgfmrqFp489UvxqCLMq1uPrNI1fjwTPIOHFCQp5e
Z6k8fNiJUPxgupynoDHNDnfnV/D2HAgOHxcYoDNI6pw9nV3EiUTnZ5cCMc2pnggP
3agA49n79Ycs08kVXtt2Tmy74KKiAQ2d/UVK9M+xP5BaCEvuGrBXm6zIwn+8OEqJ
fFxMSq1Jtc/puDVHQPriw33H6bFv2S6/mZIzMi9WsMXpL+EMr+V5ID0vmA/XmWO2
CEFSv14YyzEiund4PfT9lI7i/gifcMFggJUtLKONkbcjpCfOBdd1HxclaWpwow0k
r2PsZ0BBmmdOB6mVpVbQsWhKjOH6QttzTiO95hCGMPMTIEX/N5isXUgje6d6JpG0
yql2AnaAn1kyiB2jZDJ8PjXhIAXdOKey3y+qNQU668cyyM82kPeXTFVb1PJ4rmrv
PI2ajzd2vH2qjyhnB6KnqhhcKSAyyUCwDKuogU4QxE3As3oATrKsIOPTEC+FeK+V
8vjAwlVovSUfIJcreXztIzCLPIZaTRLneuXkmrelz9zooppu4lyddKiNHxQbOhD6
n2eKCSR/wZPIcvsYxKO1mTKKABt9VkeUzPCTrWuNYYL4o4x+EkN0NlQTXFAmCQo3
asXLPKSUZQfUUJMEgvAPEOE22kYwwnfBppJ6OZSa4IJJsijjb/0t1soVQTeqiQzb
E4Zu+cVl0bP0hEdzjP+p38z1cM/uzCEahUTdXXLApHcIX+Fch0pE3QlgcW7gJ6R9
n2rauZJkWGdEkaZPlHwjUuPfAlk/I9yDwW9CmVT5bA0NyORocWkoIVC92TkgCL/Y
nWcPdqmgn837Muh3yW58PnFyCPU1yQUY27+jLVuVq9gwt9bEZlJzDdCKZC5NDs+l
O/5m4WXEla37FPJelUj34jBLFuKKgki/KyK1Swx1zhG1FYEp6HjR2hfgJg++phAY
eNO3AsHp2xrQIa0fPex0LfWEU+habGJ55gUBYtUpSc9ll65jQs9gOf4GWF2vWPlK
5A+ruz1mHV9pHWRlB8PYaHCFbjSE0F5XY7He/UcBYgPLLdHh/ZSZ0GOBI1oyuf1+
wXViOtRm+d2AKitEsfiIgDTKEqw1oiOV92fSFrjoDBw5F9Skgt/RYXQZHPvkkZMV
u/PAZjVTsdAN0CraPNXEPiBi+EeTcsI8hjKrFwfZEZFEQbMOVhhts0yc0+VK8ed+
bIQPM6l2CufUmESqcmsevYhVjmCzgiZWz+lTHMV9DIVzFRmRtM/7w9Xue+oyM3iu
GA9zKSXy8fxNpnrHSwoaJUKLsj63dcoB55dYIoBxead9tuvK6A5EUd0GaFa5yCTC
9vCuUyhafU/M+RToTlRB8skB/8mZFij/1YxZDkWyGL9Dp/BTUbCjTbZKaujUX/Bw
uSV5WNWXziRjpeAWLylgLsXi66ymshSJpNQ1oOrJzIubmtX0fBJM/trt4JYRXCX6
RUm/Uk6j0OjeavRA/qXzLGB4IM3vWlB+H3N6GkrUfT6ybziytsqRUo3wLHaEAjWl
Sv4UtERstWhZZBjW2tl3Gg9hA/slHM66PwSx3p8spfXaHuZaBLfNBxZ1sY4r0a8D
DbSvV9s3OkL6ybsMcCS+JW5W2XMT56Ae/UmdJA5nVwqKFHDxYUaNBRIW8QAVKBJd
6L/lmZDlJTv/g+L18kYWC4HbtB7Tem2c7lZUhPBcYP2/10+ZzOyjYXiz+qhlH2sb
UDX4cQiaxmYgIkML/qbi7IXkyTX4k48ibhWgliwy5LxFe6NWGu8HcR04tnQnwt2+
tf6xewDo2PXLZhjmNtbglnDTtp1qVTgqe8LTL2ZFNKHlLOqqv4riAXVvW3k7fnUX
gbxdGLOYZvESCQPcB+zZHL/0UIs1N1QbgjRuspz36NZahF1oNQuQ6WqwA6We6WiL
2xHWVPZzsK+kQCxkSc4yCDh8KdUNuwHSl1qsutsxhxdn5uQKjdJ+PuPZlG1NS1so
f2OmuFdq+M59VwF7/lUGkf2tiRdT8KGA/XqbRSEkLkl7LHEqDWxka+zf69jH/PTy
GL4SfHUixWBuBAZe0xSY757C5VP6iiyqvGYSv9C6nOVNwPO1wlBDkNFd8jSeo15e
D/C6ptSTovsNyYC6sz7xRHByEl0jUPgcE1W3/GjT4zm36FCA9dCwlTIYKAhRj2MD
MqrtZ8+QT/xbkKhqRDM2eeDzH7TtO8+3x2DbxNCN2rNge5NDLJSySYZCr+O8CG1X
BQPJ2h1ntgnjeDW4LMJtzw3xoQ7pxrhpfq+jKftypuafYS/qLGC0W4vPiUFqOZKM
dGUEPj6rYkq3rZGCvOC+C7tLv1ryJls2fBaTPLl+HJMgco1U6vTQWH2Hv6mAGKxf
05AUDAbVzuWnXyuIO1LuGQUBqiyqVY/GB4Eyb26Gx5EOEr24JHsrHcp6Ox/78SsN
7vclraR9YFBRecz1ZIdWlr4OBPT8CeyPkdtUrd7/F08TGblVuSVEXJYTOMOYgbf1
DHa38LgqoXN9p2g/RxdNwGHCANL+Nx9fXv4DZ4P7STSY67A6GcVKeQkJoptQc/4d
+AMe+md7yzBhAPYZIz6h6huwyZXdsIm9FAi20nHNDguKS0Tjy7uUhjY7WdUZDZ2Z
7e18oUqvtpoJum3MOyje8fDwmNyfeD+Yv7nA5h71wr43wBjrRkvsxl2UeFHISbuw
L04nbqJ/i3OpqmHPNO9tN9awN+Ork+6UOsZIXyfoygNQwKmaEIxI4OzKFUptJv36
r+NkZhNQ7xySpc7XQvHVAGZ6sYlT4AvFO9UTJyY9oHU+O3HpndbxNfWBL64SEVAS
ZpDGNOX8IGSnITtxCgCqC1hU3dutt0SF6W9oRpfvWPdrBVzfrNHRqiZhDdzwIePH
nd8ml6N3Vwags+vuZZVG51sRqE7FRzxIeOg6XTvINOMPtUXcgwVSjejaKMCWnE6k
ab9jKYuP4/n0zixYYOK5ejS01yGCRfNAHa72NzQzTsEavrTcmOWoiRO55+j5TxOX
6dXvAbZBEOfRmLvdG6uOXwgvJGshxA3w6EiksZmwJqARAwsd8c3Tif+EY7HlYayT
spOnrKG0EbBX3JFRtj85bUWsKhO8ZcybCz98hzeVJi00sQVpKAGRG6oxkiXHJzbi
pnYSOFE/Og/mSW7Nc3QviYThXY5/i3Lc1iuqXy1OXOoJk9pWbL/8oMFKSKp6+m9h
BCl44fKbzhM+hZtqmJcY1OBwaqiJR5CLipJGgtlwBq6Hfr2JJyBieveNn9TEIScG
SDf9TJdxegj1SxxRDbkM06dr76Ts5iY/tKoMpp5H65YmA25Lu3qYgv6VthERluSP
axUcj5FghRGrut5bZYYQSswOVpb5+ww3TgVB6WfxfCpQFctksz9I96Wsc0rjanp7
TSTRDlTOLNmunXdZOELuVQ3ZdGHVLNGrGl+EJR9SyDwd//vcdbGgB8rp/Fac7ijM
mHzWwOy0U2xsflCxkmgSz0paHwREndTLcPEl729D/iR6136at5Zmd1lSHq/F46XQ
Gs37pKBWcpYaDXORxUt4B5w+S6iJage4bmP8GA9G0dIlF5yXNyFdCoLFgb0BuRc8
k/RdZs5/+Lr6Aeul3YWcPQQme33S/APMftnqfyUqJKZLXhjjYIYP+TpB4Bmp/J6k
DqWGJIhJLTPhOfqt5BZVqpSiP97howLSydN9M07SisA6ICgvMxK6s1BJ/PBk29b7
LZlAxJTat9HEqApum95o9K5bcPJJUwGfuWnugfy4biDyY+FOtu37F8/QysvI9alL
QjfQP41/rU7yt7NZjafv/YDVXL1cpqGhJ+zBlewpgcrQ1s/HI7jV3drsyaj9C22C
UlGv24pF0rIj19o4XNw5OCTi5HZGteH74227WdlzPKp4r/xYWZUVy+n+odu0nGZd
y0OosFz0dBkaEBfnFt5mmUtvrSctCDQB4qZSEgF+xyt5AoRUUZ6JMBmi2USXCUrX
3EIi7q8ciSEiTRcvT/Ht4pIZpGGJa+zwZZac4xQtSKo2r/eIThjYNsfahtmD48Oz
j9ts/1IIeBEmz1njNrOLt39uKzU1VpdFFUuzeosCrdR4HgcSKbNLy4of6mXoNldl
hpMIUaR28ykpPGuetYlmZnFtKvJVW0n6ncGmqnnZj9xFxN9Y/xS1E7YQ1wlt8B4C
zUkJGesARsa3XXeKeN+kmH3CoX7GxCksOK4PMLMq/Q38yon+b51qH6wUY2BGucfT
6+4TDuiy48YxizJ6KLa5GadgBVD1mvMNHZpra6ySsM1rWMKV0ksPHxEGGz4CYlMf
ryFvANLfFS1ILyzax/tJg1SNRfitoSLtqQOUd1snXhVO9w7fxCuemgxk87Up3UDF
xgxwwWIJ8/fjLrRTyZz48KGQBCJV5umjbHev8lZIGRLjppkjL/60oF2fDvQY/146
U5jXtZFJ0J9ENqMYnBdU5Ld06oDCzqWOyGASGOgI0ewJI7Vul9AP54KhDagb0lTt
zg576lcA2ZKXJiWBbz3dvcG0/Cm4fRI3vbLCXSzHJjmtQRrSuwkOdhxOx5hsmzXB
7dwN39uzEFopNcy7e1BhkQjKUO6kd8Dzty1VO4uLuRunT3RJ3dSdpzlxIGpd9p5W
ypFY0MMTn844ke/hS7F0uqiTQBsXcObZgS1IdT3AuozzoDs83W+49axnJu4dWnbh
YOB2XsQP2HWynPj6FXAVJYKSSBFAxuN3DPmXWYfGR7afyBy3qgAy7zIWbmddaDdb
l80YYOeMIlZxBLcft21ATcMycXj4KFFxlak9Mn5pdXjFAqoqJuZcRkrH6vjX1VOP
OD4osCZtl1niMpY8FbWBiwmEjl9bfWTBgleHAsY/AKYLRLu5AP3YjaLswzQvQoZ1
TkjNNKqWsfJnUPkpsCgpuXwR+zTpdfgWZkLObo58zo68T5fUlopWxaMI+31CFzKG
ydnintdGZs1/UP+2hMl4s1xHchxwHUFrJtHWiI83nb0Jg0BSjesRHM0tbAxI1C4p
Q3yYd7jBWpt0RGHApj9Goq2NO4rsWyiielHQ/zMlN5QhFivhjFDVj/COjPqbd454
nD+dFfI3bovlKTzR6hLhA8j40Z0516nDA66gi3nmXh5ohVNfRjGLvJKf7FFql0hl
tfpCPbBi+j3fxdbtukhe6sIatWCcWjEIdeNy2HlXAiu+JVMPB16PZhYscW65DDi6
6A/UM654StZf+tOvUZynND6Itn2iaIN/viko2etzlyyF3gX/ngc1qG0FwM+5M1hd
Si/7GHainKvC3y4so0eEh8+kcXcDTPgg8EWNvkmFOAk2HTcrKKwDI8AopeTX1Zob
53XwaNCoZaX6j4+IvwtDycCblofzBYmDjXMhOuEXa9wUphYWAvn7LYFQQGsv5Z3q
1E4ORNp7ElTkrAah7RrHBh+a9hgn2J9MZOzATRAAezZvvJlXGenMvoO6M0edJJf/
mVR5GzzBbITyyQzkCM64ls/98/EzbUlIdnBO8B3kavur5UaciO5ZilTydPEPH6+t
yrUXHCr4nqK6CeJWrxqHdsUJ9AgclSmlQpKHOchoF5dL9NKgXeED0bDZCKGPYPLV
Ye3lAPRS3JrI6kKCzPLf1irOXvTi12Mgqym8Qv65vaX2ttnHQR2wy1xFe705kO/8
z7X543eWALq+19MWruealYGUWQ2roZscpF0EIhvEWwRSTPCxXo/c1eRJpO5GO+62
NZQWbGIqi7AFvqE/O762rqLb1bcrbLnYEcwsd20tSdSKou2DlhJ2D7fHRmfQJm7Z
6RS1jkUaZAOStRIVwTnTIIbzUSPHdifEbh9OoKVGVx7dwciOktVyacyfs4BYy0Jb
FbQOzTjfO6YX5HzycSLBK733XwSvm6BPGoGhJrj5ilY0wa3dz7HMKPQz66t+nSZ4
nsvhhQrQVKBCaZ2XDGlRRMKkzBJtUhG86fpIMpYQhmWlq9i9UDnyHG9iQVylSp/q
zBeKpRs4Afrhne87UbFOsGbNfMJhJ6N73/yG0S8wfMKkc7VxXpDdHm/Km9c2tbl0
NRT5+QogjvnvRpkAX23GbD33s1sBg3EkAxszmWAOdH+NcvDo9xcm1H8pDfkYr0e6
pv14sMgD5vgfbQ6cRCfxf21r+Rk8rOy6fptSKd/+YhAiNdB9bnQVETOMTQa9NVFP
eTDcOM1ArzHX6kepCDInX4BABuQV/CyjyMFjtvxwHnU/n7CDpREJ70ZqgrSnb2lR
48VZWEscQvgTcGKp1TbuuF0UQHw6zcN8t0HOHFLEt7ghxZNeRp8Yp4iNmDceYySd
rgVZtRMzdaeahgLV5EulL10xXpxFUMbF40LILk7NPf1RvgQYht96+POvAY9n7QJj
wJNd95bV4c1T42IlmaSuEEo8Gt9zqrXzwO972K8jlFGqKy+ie4UVc6x3niafSinv
ZQB4wBsWBO8Jb20ww86LuhF+8Ij0niAlLAFQVQC585hmkOujo/ax4IFxDYECpMXI
XtcPa8/XaV9hFoCXAwlti1t5IpQGjoWGcHU532pup488FOGpT9Ud7/xHLydT4cM0
LKNGic6QIhFJZ3i1kizgTG7Bcj0HZEmonVETHkC46n4r09UMuctFkP628uq29BzJ
Fv1V3V7/3QZx4e788nl15A38XeV9ptRz7SawammaIGu4/VksCxxvVvy+Udo4UDli
20kc9wv8OM2NMQ0of8X/ZbLvtVLCH3VXJnNxIA6M1raIOfgbudYRbDusCYdmjNZi
EGPGKGROuZc50fvSgyHFx6x7fy/VP/CPz/lM9yq/XUFYmNnqIaNzbVqYJtq9x61H
3Cixe3qzIbGjGhHtzeunIEPSIQq1/GI4pdfzFTguChDnAFKDH4TSHb7HzPMds5i2
AEJ97ouNuuV/AIgbml/5/CLqSzi39lw4DCYrPfImmb0MiB3Zb4XVgJBKfuanWGoq
29gTEnu10H+O/Ru8bQcASNJRMG1Ujl0H37ieSJICVc2yeePUYnM3m8TW5urG0jm1
fjEUU0+pnHLBJBLyDRGLFWjPoLsTOqTErsUjPe4YTWcZOOF4YCfCOvUQNFn4k8GM
IwqR4uZsx/V5bI17psZoqOqy5dPz0FesGkwSKeDPahLPYvuhTJwc1j14berLGVsN
RsMAjqEr+C2X4uqoyEInWyEQCnvKE3i6hsarV+o3m6QtZqc79xcvs1szfMXJUMOL
4GK5OY8bhY9/c7xektFydErU7PMTItrcwQQRkdYQVJiKPgFRFh1S+/BkEvzz48tn
MWmu6LojZ94us1UD+8gAsPF6fy2YZRwUmEHRPfKHbgjf+gzYA/QjcRfuu4Qad/+s
12nWIFN7QH5UcvDkV/vusA4Ts8HnPIVZXYRIOm3IJX/pvwpj6HVbamRQ2Ad2lZbi
nMTn0aU6LWnam8pUuK62VOjdrOsKbs5Rfp8xO1nUZKBmKBjkqCinx1358PEpjA3S
EgdQQPOISgjK9EeRIGzDgdrt+7nf7t0gVMLe3c0ZEWIe/DaxkWddlxpUnQCAH3nw
/wNoHjoOcKMa14DdxS9fFtVz5uGSsp37LM1s5cibxnXIV2pDGlXWWPt2tfRFYE2I
SONMM6B8IQqvddsWUWhP57PibUy7130ui4arHbrJytZnjKa7oAVxmtQv0CD9P74o
A3zNbeESpQqXFG3aTTruoywj0f+9LUv4W1gWNkC84lE1TUel5mVY/fDRRsgJchK7
ChmFVr1an7SGeuw4XK8CN+8imbN8USLL1mKAEoIu2uS2Qkd7Og2xqDOmb9Fy84tr
9HZ7b+LV1vBleqDXRKLmCWyr3WHltT8NgIASU7Dmo9WG9fKAoUlEYtgxgI7cZuco
/zrdiAE9wz2P0o6foru+iNX5zp5/mjNkle0RAO2i9o9F2ILdR33O+Hh6y3cE0VOE
dEWaQ4gAaGzjWTP3WzEZz2ordRg5isXzK84Mp6QVcaLKqhzkbEjssUQ1GjlsS1WW
jqd9PGWaftQhuZNdwv6q82NByAiuFRBXWM8lIKqxCVT5zVBv1A0GBc0HRrCp+MN/
KT2Gqm6yDqvWsz/vsFTOV/L+bDgjcQAakwpsADtSeVPjlVFW7rPMfrkIsXuRZmEI
ocTJgUHDWHCc9yYeLakylU7QZA3XWhzF3akMTUw8RFTyiIJJolpLRIrXztIjhjJy
jICAHCaE4FdAnY2N0noMK70Bx18h7a2AtzpngHCFUluDQSyFJoCQD9sVeOEnRjL5
PSn+Nd4CdYMKIInhV61AB4cj4ztQM3a+X6AX5nzYDC+ljJjsAQfSziawJeTtzFds
ML0Jb+S8IZWEcUyy1N1MK5URWA39swzRM1p68tS1GEeC4WrkTvlpZ1B6bNHIK7sj
MDey4n1rw6mlPPzqU7egdFcRFDD1GqgNaxv6aRAZqz/0PCfJVpjuRL9jymdyysyS
Ag8OyLiok+BreOhUylLHXwStF9XqMdJD9IV6BDExrWd4H4rs+1Zmlu5qDQH/iW0w
LuLW35Tq0qHHSaFBUUhQ5WFNNTsPZYGDRgsQxEcitfSdo5htW6vxSPE2+yoaA4Hb
2dAIsK3tecZgeGcdPthTYFhbrWR01IR8AgwCBN5UfEtZ6fFyVkLW2zg+LD77zWJU
YnlNHEdK/nxKsKGcaixtOrd2s7N81iGrlkBkIS0SE++ov0/NPkwKoNhh0mJkB8pB
U5e8KtmM+VvG1V9/3KaSVW/VfxQtfdeu6dBNoedY7yQsEbWBxeruN/gdRdlSrR5Y
DDQr0OO/a7qbB3f+u40oyon2vdUJZ+3TaHc1HMTHMo4PzRWoU9sV8m6V4JhNULnD
TzfdP0227bi6bdOSnm0UyDcEc9rrzhtYemKDGz5CVWoB0gKY/c1qn21zqwJQWDO1
wY3GBXInfVKOGOVpWAkdisu8GqCfgHp8GyCn7O5SVUaHdqczsOGrXkNabSFpJu5Y
HeKEYkrWpop0C+vLg01DsQ6f4m5DSug6DtN8eLVZavJVydv+yGyc7GTQJgsinvoG
YDOOvRjv8+iWOjBdcCt0LJdiTS2tjKn6MunMw0KngZekux8/Yme4h8OcYAHA2QZf
q+E6z5hARMGgWat0dHeUiWUFUe9EKLpCV2xZl9f+Y7shkKNrjznAGNoTyfxzE02D
u+Vn/dmvqeFdaBWFh5ly0Ym8sDoOpkqiw/3J8KxaQUbX36qhJLjvRoLyQPOszsj2
ce33aoQiOhSd6q2UqsXFcLMbiwJrseSSBu8r+hz6P6P+xAAo94PGOuS+3BIUR58k
N51JLalwb4/LSBdIMLEwGRh3GaLcQG+kBdeJsQkO5aO6V/jtii0gqjRZe4A4nitb
zF6TprbQNKGY7vW7EdhG2lvl1FuIrydUs4lwRRZ6zxqRX0DyTl+TH6YtOPtC2OlB
ztkaJybjtdAn/+piRc0gZpt1MGBUWHLFQijH1/DnwA+ikr3XnW219GgTaUjESblT
wrlDcQawVQBnA3s7UX5vHKbU6tmQ9khJ/jpEBiy8bWYptRfv+Ul2yOWYQQrgpAQC
Nl17r5yeFKyixHdVpZZkYH27BlPWIyDG51Ifs8tfFNji1uwDOuoEWmuo8Y6GZ/Nd
UkbUrIdt/Wvotezeg0ycPlqSsKoPWvCp7L1sgP0EFzLCcnIhnQKu5FcXBi70yWbo
slwFPJvXoJkqVCsHORcSpIpsVWkTepY1zdHhgR38WwaOjfTEZeB5ggZ309T2NPab
90fw4UNB2ibvnfLHuiOGadYybNFu0kByIqIOT8wlFw9l4YVa/eNiWiLRkdJUP8it
KfxT17LRM9YmOZ+4gKrZ5WzSDBehCMt86Xy4aLXJN9tkp5sX3yrH7gxXacluw/hK
uM4qRzbi6AXxCq92Rdt2nWibNJxe4/pv62ro9F+DQFud9h65u5G+9UZcdwrgh42/
uhYUc4CAloVnhq0AwqLarsE9y1QW4cyJruu1xLhE4IES+feiAEEqFv1zMNNwNQlQ
G3iQixVlTHn2JkLEUllFkihctNY99H1gybQ9X2CjvzXtB9XKea9ZUdtRG5jdvVXg
s4wTCMZmFyE1GtOJ47ePxBS68QnjrH6utQJdkV9buGcARkqVySqA7ptobBRr2wDq
4wCWa7UoH9atUgJ4r2iwcRfwkso0bK9KIe1rZq+yfHSbsA0OnEbbg1RoaeQ+UDWx
YZil6z0Rpmhe+1tJLwFl/X98DnrqLVwo42CiDAHwmlFXbtx23uaE/S0Hgk+up10E
b30pxB2O0/2r4uB3h5M3DRzAlqP0jBOFeH6b3mKHZTAQ/hZ4JZ1LkWbvPltSEOHm
HFSg9B2wNTRUIAuTQuQUZnIOoGxJwaZX33znMiGOQEvCWSQPZaX8jDZ67DuoTRVY
42Hg9AhGoxf8Da0AR/bQjGStO5aJ/mc/CN9zt6XJ+P3Ur85LOBIIlGR8mR6B+g4e
+KAbeN0E6qvLRCLJn6YNLHuwfp/MAt2966kxVcnusvUsahgLWUUyy7LiIpX9wKva
dxSpNxcS4ew3HJwRkr4VCK/zcAkQE5Aw1ooieORP046vVDtQnUpaz6zTJLVDZZKd
VSWs36nWHinxRJ2HQuhhxhSFZtlm1ReWgWS7DU5s8pcf3g+MlJeXz3vgwREqcpyq
70N1mPW9UFNZHnyCISKOiO0g2+1A4lMPeDwc1/rybzIIxfLPKUZP9FMRSQFd0zTY
NErQOhU1AaL+5dKM1t2m6KfWY3wYJBBBAILv2DCKaSKDLo8YL7BOewpjYDdMN7hU
/at8HWP9QYJbQoXoO4sRvBnS7/qQiBFdG00xp/lZsWNPFIZj2dAJUOaeef5egjkU
IXtuf5Oz5pfrctbyruntTExgDMd0lLiYm5KdRp1KsrtZkRyMb8d43tiXpBuv9QRx
pxLz15zWzN9vODaVkvVCataupj/K7JjJ8BG2sT+28Y1yv/FdtuL0csGwsv4jgBMH
o7NutpYsqalj5OVgWJqz7/fjlN1AGGxx2VzYtc2OUxn2KHrUtBRGb52Zdii8fDJc
97ajiE4PO7qEAUi7UsLzy0bUaeffsLLiuiotXtfPJ8Oxy0glR1oegJ3Q1X3dmbBR
lD90xc0rsWS8wZnZshMyTHmrqpdWnCNt8o6JuFdmzUwy1zkfskycni0WfNWsu3P/
EBt0XKWI1EQoPrx/HYOx6CsdAjN7l59ZxwI5aNfVEyP+N0KAuljE123OnNblzRLR
Gv6gAZ+LdXrTpVCyMGh00KHypRByFSaUY07uOSPR0DA50gW+Ro/TuGf6W+ZqaO2K
dlEtQ+2MCWgQMRFDSjRL6rdO+x1STwIvtgGAYDKFmAP/8kMgpEA9Ml841dmkGadx
9DNGUaWrnOFiPlGuM3J6Fqb7XykXJVX5JHpTM0lLKh/q/x7R8A4jCawOYCtk8FTf
ImVVMp654YXRoFMoIzrXl0abkHlKkrmflVChQyTxoB8obejki/AznyGeJGKz7sdB
3/iQtQIn1af5+YiY1RnSfRxtqDiRphExD9L9zXtJI3PAXhF1z9q8EJq2DAe582HL
1uf3wvWHTjQjrVd88E23xWViGder+oPj9YipKAq5s891SfXVVb4ZchFSj7nI4Cj+
psMQjNxJsSNYrAeHGvn63NmqEb9aNI/ZaFgOebuNLR7qC5i24pZrUEXO8ElPSPs0
HFom1QiK/5Ombaf8z2DcqBjO4+6UgOlobQMF+kMrRRH44Va5zCBbGn9WQP9/IfyC
XexA+DZ5bastRXYtQTFjPnA6bVo/JK6EaLbHuv7ZOTa1qsKmSF5J2h6A9GJkCMBu
LcyNMTuyUtHJsnC81soiHA5ibU61VNI4NFLtTIjyMm8Wa9d+ADNd/Qqw3hP2ZRwm
ISWG6WGB6i5ad+lfhDJ+7J/hLv397TxO9UzVtH/bcYDsV7E85sl6cUjZtVZdwTN4
sSzIP92ekwqoCvrB5G/eyb1uj4v5Aeb+2DouGikl26gXz3Je3Utx6On3X3r9KUm6
Nz4BEUknq0kHKA6xQx7CrkKvkL8V2q+LEznCNm3UtKccnEzzgtLObHVWeIKIkvii
jgBpLawCu2DjNZD8ri3LeaGhO8ZuQtJyTQe5P9TWEoU5N8SdkrgFWcyqtDSefWJK
7xwHoE/7l7vwyuj88a2SjDK2oYU173UGg5t9g1swRZAj4O0nUZz5aaD10gM1E4gw
oVjpKPH0WA4fTZGexzDA80sls62Htz41VP6J3TVwhwsN9U2A9G7RpTDx9NJ7mg+1
KYeO+M/BakMc0MR0twg0x9aIL/qWgmlVghhqbpgKTmKI0n81CqXw5YiBGiO/l/qO
K58fuzCSsixdR0j6xfwHVEQ4QgNHd0PNCMwTNh/R3lAks071k3Xap5kwpvPFCLl+
L71Zbk/OWDWBF89k7C4mW/Ti8xeDQxXOq5OjKVP7Mkf5qWXqD6R0B3ym0rlsnAKE
zpqFRl1hN/jRFfkIxGMbiuHqjHwN/HMch7wpABcRbC8ZFtMXjX/KmNkxf3CAHaGu
+yZasjed2KjMZBoG6PTYbCFct6592Mm1wc5jz477au8f8oMFZYcEKIVFezv466Tf
AWI3hvUXAann6KsIPz+EfKDHEz7vdC/Ku1uZxBhcq6ThGu6Ty11Cub/TQhXx3lHg
siZRQKm9WZcwC/PdMifXns7KvmKXH00voSMje87HQvUJcY5Dv9oWMfXnTCvlCVgl
VBk8bNAZ0X4sz8HlDgfVVbXymevYKCL1SbcIFYK8tz5XfKngSfuc7/Cb68n1UAo0
O7B17a8M1zOO0jYQDWfnNHsjJNKLqp7iZ4FfQgeoyGwr3bUxbBx8QDSsxPH259LS
cchVqUf0uQG4Ms4arahMqi7lLKgoK3Bgs6cKCoYtWJMxI4r1d8lpYQe5/s/zpl2t
rLAtdugNxcr57iwSTHQSGieIk3mVJ2YrtEhNYRMP3zgCAiAliszGisEnAFFfURXD
kDoRnapFnsLb2zlzki5Em3WbCbA7HeAF3dpI7k+NY+6o7PaxPVGimnSPQGSsB/Dv
EiuFw8/dLNSW5PCAqNSArO+q5Y+E4gjeYH8eByu804crcmPKADnEG9LXIF8ZA87M
lqTFwTdo4cRU9XS0cpVLmqzdkZMLXp2JZV/qr1awcVyHQS2HZ9KhkgGgECHGJwv+
1GFO3NiGea3z7ddXyDrQDTsYRgaKMoWFGX7EgNaOm3WZRT9KArN9yytkZyhwze0c
NTa7rs/7W+1WDFiGBAiFYS5EbDcr3yg3405tbEx22DzaqnC6sPw31afasrBK1eXg
xIwXllfG+NP3U8BuSSx3KfUz5/ckmQMJAGhsaBdn7oETVMZT7IngLaV3IM4H0Hj4
15RLTaBFX8DWTcLbddrwQGWqOTJi9nFdZZrClMFYe1UM7tw1EbM/77LO3IiPqpJJ
nPpjajvO6wZxjjLbXJsQzfFrdNHsrkvttr5Tzfr4wLkSvpsE03/ZSe6uWEXGeOIG
kq4Ey09dGAx6gGkOA/FKeOmSH46HQqxEKCiACazN/+efsBmvYswV+dv6/APf6BmC
9CB38FZiCNWr4uZHkyVpqb+JkK6oRCJx54VeMkSWByFQvcL9/OFBIxKCHgLWrV+m
8u53JG+kYHvONoUf5kZG+zfTY6eWwguZLsSm4AQxg3wdQgqkEIkcwKb/tCxboxVv
/WhZ4yEjVrZuJk9iFRB3sf6ElOoumfBZD7Lc7cahKzYTCGpU/+YB5BS9qViPCLW2
sF2ng+3Q0G9/JnxS/KZBEHsbtsEI6lFVvZj0cb3DdvRNNBgMOY/W4+XZ7CJnTl4Z
Jvc5dSHhwIQkohnaLZZ/aGGDG88GJrLGBDjh0xhlVS8yIqi4vVPj9nVZ8QPGm3QG
LM/cbkb89y9CtBPzafNypv1aLm9PiPzJ31RuoHjYdmTfdrYJsnqMbfna8bVYawz5
2uNh4SWOKqrrgvn0qe6ykSoG6to1xeGRdXwYTd4m76+Eovd+TxhrUthiPWKeEYMX
SmT0KUINZGTiXptaXYoG1mIistYTnxjwYSot2TXiG7O0oeo83HAQ7pKxfalg8wMa
zpeIHjCqtajkqB+s4zRCR9iPtbiTMniRhPLuU61vRX3FgjXHBCtLp4v/TxkAebJw
u68CbRjlu3Hpxobkr+djpV1pkMEZeBh1HUiEVyaGsL3zRhlSQ2a8DoAl9RleRlst
rSQiT3HhFCx6vp2H2IrH/pdQhUcH9XG7r9mYC34BFvjIrfoxSd0xYjtXUASkjuf+
/2+4kF63lHsjVLwjbsc7cDPT5qi9MvrvQnCKx+suy+KvcnGRhr2OopytnaAJNocy
xUyum19nonyyBi/1JoZ+M68lCh6nqYLblU7l25IklZQufphAbcLhgKUbf0CxZXK4
c/w8wy3d6M0zQGvpv/C2Cknc8MOXU+5EM/nvohQ2Dpr90RmLwBHMZrGp1imzNkeY
UN1YqbrYurEFaSiiY2XUzjpw29Z1csi8imHzBqXNYBmZBob9CrUsrVbt+r1oYBf2
f53rtMXCirRBH8eXL1qsRkdXADhUWHeznBcW6hYZ2SNmf+63Xiw5TNUmThzuEpwi
ny0+Ok0ULaQ/oscS9K+C5QssHXPTfYfuMVv24cBIsRJA8IGAI0AYUY7dZbNaD0H+
+HKJP496cGurB+gxRoLli7TeGF1gJeFhz1rKmro/enleXhGLMedP2okJQ0FSumzk
w3eOnCVRMyATtpD6kbKfs+zxL4+tuo3sa8eK1if84NqkMuJyU0gdW8v76RByJD9V
YfuXBW6dtVMTp5m5uAF8p0sG3vAp3QZb6JvmTRTiShAIDNqMBeV9wmbIU3kwnAEY
vhckSpR1XrWLxDpqcnfReB+ruwE7evlFX9WJG7icoMw87p9CH/xkG+P593lRJjCz
05Yhpul1fKOfp60BJi8Vi/3F0z/Dk8VPKlECKwWnyJZXkZjYcXdH4dzvHKC8xOr0
00GjYFjIcN9hdgyobP5FvYrUTYd3FLSoECorl8QrZh++uuEcA87+DeuiPMoZmhYX
T21hYv08SOltrVtcQc0kBcuq8iauShMYoDO/yP63BgIHij7cDHFOddCqLcBNK/gd
mYqAVsBIOv4RuO9zEeGlN8cdN827PkirHKXv6YnOoHyGuZSa1KeVK4L6HpSGjR9+
209NeBUuKofL3QhiMCnV5svwE1QUwsd8cues6RIfxRw7xPYhoRNQeNTA8E44VoG3
wyLM2Ffbk2yk0pckKCabGwwxI4OQKLr8/wbkm0gaxD/UVlGXFFvgPkpsrSge8glV
MttwVf2SNG2iuEpIRox9WM//ZnQRQ20p2AlhCPxDMw54PN39qvtARHhL19+xTHhs
kFQeeVGnbLQpl0NloX+N3p/36lF6Hzrl/TF54A0fdMw0/Utw3HaNsYmxwOnwzebl
jNdMf4kL9y0H7fN2VIuxXFycItX0z7+1oHas6E3WYOMXYs61ua3e2dXmF2GZSxY8
qKGN3UgnxC96Efj7AsYn+uAT2HDhsg36uKJSWnjB3a/Pi6mcT4QiigMhb74U4wKt
tPVuJ4GmnrrA9mPvEJ9npVPJoXTGjZxqibp0mMRkB0uRrm5lIsNFZmfG6/PI4z9D
8DrGatQAP7IfjFCQ0lX01oQnAhst1Q6G0saDo4FiLCAlgv/3pmqMfVu70imR911w
x//YEYenv/XdsLm4dhIO1MP0FNpeJ0e9xY03unukzfgZ7KATmxeRZi2MteX6hESl
vhSZef7LYAF1AYmsRTuQwRQxetqjMmGijVaMCXHLJ5EbAioI20X47bdKvLww6Qem
mzQxzuQgcuVUfcoGQeaP/0CG8HvuPQgl/7vce/DDTqhquPVndEfFcAMbEyylCkDU
4QSeVLHtY4bCT9LtfUUPSJbH+YPizNrqfHcAVoHs98UKkCtR1N0ZwVHV+CGGJLkX
2NbujpxCjxPcYVJyEj2hsSi6zBuh+QpUBpizuGCB+ork/b2jumWJxzrvKnRkXfLC
fivPjla5j4xyRMPZVt8fH7fJg2nFbwDOgpgeTGLx1tLqNNwWcJpYl3QUshGlzwfF
mCVSbGX4Q5OjSNcsAJgJ1Sh39G2nLFQKcdr9N5PW5DxbaewcMI9h7HsbC3fzZ+or
7d6JvNWfr0oKnFFISYy0yOfXvHMLjQs4OQ1IW/X0rcwPzDiP+ktAujrAcisdE67E
PnOcr1pgMZAAq/w+mToT18FiRmsVaWV+ecI87G8RtbeEPmUs0OIy5IVY58hM9l2I
NEyuLsl/AwuUasiIWt66WiNZSgEfCNEE924HQB//0uNJPXeBKFwCOyYJ6Yay1cOa
2ZkX4ZOQk/Q0j3yhGWaG1zOh68azeK7BXSVpk/5XZCwt9st8UbCYkBhYeU7fqvTO
xlEvogV2j1NPg+CUt3fFTuuk+NM57oKSc7ZEAAXDXFjGiEKWVhoepAIkwrcFllXY
+OzJPSo3HoOo1+mlcmYf+mv4nIHBw90jZP7TEU87EQ4j5vv/sQ/8bGCHzmHqNnMU
w9mYzurQe1fePg8dhVK/SrhZCjVysGyt2UwEMHvVzb+XyJzPbLs4044IdBycJYeH
O4Y4+HbR/nOswUTKrlr3Z5W8WP5We0I0kUq/ocIHhNB3/O2NtA2Z1M9d2TR5PoFr
CBgG9jgYcIGtIpN77nl0Rp3hX+xyHrYUXOpmXZuT+HBRPiMR/tFQ+W2lpek4EL0X
zVb5UQdmRvPrGepiFsiWtuq2gDXYq45gDoHDUFd5OdmN0lDKrD/DgKocwNdFyeZ3
tQUrpaxq5QsgN9zNOYb6Asx4ui1MNbwQIxdWL8ikVTWd/A7ini22itJsNLdI0/aM
OWgb9sol1Hfa608z+9OyiuhVqNs+Q7cFvoChh03WAq05gdTRsyLh3uW93b1D8uZA
JdznHCD3nym2vnY/Z+U4wdHqGRJAkHk8Lc0EdOzxjT8PJzHWO+60fwn0wd1xs8kC
5aztcl6O3FAv+XalnJDc3F6DEplEdKcVj9b+NlpqmEZiPCOTBX6R28nrw0SoPx6H
k5/a9ehuxb7oo+SRk5f2H/wz+ES1HNCmNeNZviiaSY09XiRvn2I994PqatEDkwki
19VoOxSDnY/fzUHDCUA9uh21yZ/m3agJ7zamGx9xzdytIpOMMO69dkYbFbWM4SbO
kJCNT5ape0UVIZBZSe2SqVwCTVPIeABzOHELH5zcoUMmb5crb3Vv3EoIP9p11obK
/GMSL23JRKFshczopU45nLG56fO2VCu+5wLA+IXIn0M0ayc8INUzRibj64pl9qg0
jq2jEuEIBYVorXzQG9KFQYbrRd7HfjlYFKE1J8CyU2hrxOmiCtUTIybOqxNFe8DB
VJAh9W2EyoOL25iDYbHhp8B0xkCer99A4v0iEhL3/5R1XX9Tx1z8pXD7lIJpV/O4
D/9aLAP8DCztIpxAROs+wDhqkxfwccs5ZswdY4UBJMNzy8dYPXAFqu/Xa9ItMQQV
pyBIVMakRszoPY8yziUWclsPd15j6DdYExqHFuKmvDM693ijSVlfzCsY5QRy3XSh
AzeZ97KYSobvhxr10HK3OeH+V6XdT8VG15xghPsDnidPO9trNQ8Tjve/1auukSH/
Ewds7ybx2ei2deqpkkunf9o/i9I29/dkn4KPQvtGJTfOxmFoQ75IJWl1wV1/XNLN
w1LZqPWHwUkM4InXhJstqnKEzVPy+FLMmoNo07EbOrwGBi/91aeDmd98Dpskt3+5
sUY1qOqVYEHP5QbP7Yv6YO8hVGWJ9yUHqDJnrqOXAxm1RF2Ef876C62CWPu1kINN
rlYnji09teVscb066T96Q4ObSqP+PSfZJobaTASMIyqF4rkrLS/K3kHVggq9t/XG
Q738A8wm5+uywFPyorsuo8ibm63XA3QhG8Lrt1ApQPcj+ePU3RCOZlWe+6OGe5kf
bX/QupzLT6ketp8JsGnzimpYvK9ctrS3PyvQwXG2FkAYutAeNCFr0vgQOdyjkpFT
SVUIlBffL5aiM/gYgs1bkL8A5cxbji+f9zop6h4hKX+1sAsH0m0+BcxqH1E1hqPo
Oma9J6Nyw4shqD4+ggIi32gdSXkeydNoCw5Bs5XcLiiYbhAJlkMWcxOMc9TzsCuR
s2v5Ejrs3p8fcE92H/IfLfxfuIkHRwd7YmtX9hccoR5eo1uCpkXiomP4EeIvjdWv
GqHwfKuXbmgD+e9sOdMTZepLmXu67AbTyOz5sAFcRb3b3CO0BShN9nJnQNO/YG/H
pOyEH2GhW8Rso9ZTwukZ+QSDoBuZoqvNpdCFZykipZgRGuvyZf5jCDCkzK3ZkcZb
ZnBoHC6KjH20TggyXxxBzLRfp9W+XuPg6lXCFbdaVOJ+PFBGuIOmgfzHs7TjSJtv
70W7+gayMfQZldaTZPu7H3XC4ROaOJfx3vG/P7xKVOkrLe1rhVJdAyUbhLPvT3cj
L9mMclFv9ffx9CdRPLk/GHXocv8dGpDj+vP4FhlH5S+wVqnVnChACYNbQk6gjtRT
PGz0fSVfQZ5ROr0UiJKXiplhC0iDnIiuMU8KNOzstFDtQes55H8Uc8op7EzrEEJs
P+mEUOy/kxU5nBXTUsGJ8aCIP8vlYyxvHdO5zbdBeXxmtjKW915OhI6jX0TSrHSW
eS3vw6sshz+R5LMjD2McuRLp8M/NMMQwSE1FWK6KurNDIz8thDBegqJZ8x2uPHGF
ry8WDhHLn+O8VE+H1QsoDQELcJT/9xuBDy7VX9mrnT78yjeXdWrt85XWcOAviYEq
JXyF4h6b506ce1ePPo0a6RCdCVFp1MkT2qHJkJHO43RKY47tOfQY0GCw3PNe/f36
Y01vM1TIN/6kI3VcPvYDO9zHqjkaB81C+PuBIpcK/Bgowedpd2ls//rl6MBBB1Q/
FS2LipRsRq/icnI71FfrWNlSLVLn8OUXl2wyh9vE636txwu9kNQIvHGDNHfjB2eu
wEKbm51llc7rhvylvgwm8XENE3pgAYv7WNLfHwxSXaOAcgGksjknTeFjPjseJFvd
JobisToPkWkcyfG3csC4E/BlO6lG9W08Ce5WKQw1RxMmaFOwGmYBAlA9r6Sjy+VU
BJqF0tQoGBPdkh9VLo8x70Grfi7rDtb6PflKlUjB/13efebJDTK7OmyISVTv/bBE
Pt7XD14qqi8K/L9sqHPF288LvAvstAYnV56PbCAjUGfRHVhwR07Nu3nkKsSaKmVx
qMkP/XOfWhCbQm1oTrRbfMRdfjyWli3pIPMavYsT4UP7m1j3NmYa6Ywnsl5KX9QB
1ucuijdVWT8KHdSlVVhx21Sp/+H7NdyR9Q2bZF/DfUvktjy4ywKevLfhVXQm9FDJ
6ENVslY6wBlv2z8SezVK+EIJrrN21dld9Q6G2sd1vjHwiYqYASutPzY8d6xueIbn
UBJ7uR0GqbZD1BbfpUszyOH9qtDoP1qehQoOaVByIvU3MY+BcqZQOOcdY7tlAc1P
dGTTrkP4WqWWN2jZxz69PDK7giGXJzxdQnBAmVFvkyzL2aEkv0hSRXoqfrr2Jvui
1nr+73gy2bv8ilgnr+DO2KFNgEIUoBbqs0nIBq7orLXdwE7oDBt0Yp7oXT1WoSt4
qiiB/nWruzL2XyZsyW6mYpYk9ZGoyeM+19+X1s8uoRdfQQyAeKH4Iuo3NxFQJuW4
6CpWFgUGacLJqKbHaszz35e0A916T+rC3gqby/ansSn8o51W/x1xhnuEeEYOiRj8
gegPtuQgIBbpp1wRAKI97/evoHbngLjMvojzp+0xF2PcIGYEHWdUaTDRYSJ0qUdh
F3TsNrUfUxoluz0WKHQIaoBq6RydBenPq4trymTImofaN3eANHy0SAiEl6J6/lFQ
djKNdSdwAu1Wnbx5DUFxqtUIx3Svc3IwtyvKwPSeKkAADY7yiF6ZW11Ev74ck0mz
xEcNRsuyffZ0HkhQUTj9FqBY76Y5rPduiz0D2fZfHETWVryXUJjpDHjM3hIh9fij
J5N4Vz4VOs86MYMmv794B4M6ossaUeDWM0O6lzjxILbSd/UINA2amuP/LkEMcMsS
VibQiZDf1rsd+W8oJCW35J/o/5FPw+YA4CcXZIHfN9/vkR/n8pK9TA7hKBqIZZ+R
rHr5vPxhO8tfAtCE9gM8P6CqaxROEhWS1AeabbOAs7MDnNOz/kqlREgxdqzfBhvY
YRcMglFvfO+9JCydFUIl8NhrSxkCvJ6YyJIHnwOK5+D78vdukJa6tjfgVZc0lviJ
YJT79Yp1/XTx79BftPZ75pLHqfF6nrt1NDWpiio13axWcmRJ2KjXmlx2Z0Yw12qI
B7sSdEjvg0c0J+p+B/pid0Y+Io+iz40rJ8Y5+awhsmeBnzK4aO/ZYRqtsu5V2G5h
gcgWDuHu7KE6EgohYBGylwvy2sZLM2CK1TOEiNFujVibijfqpkLcZCWyYMMh+CVg
isliGoA+XnvaqtzJPr4lV7vk7Oe95HvaGatuQF8zjJoAzMnCnfqKWVJQO6TgA7jH
KevPaRKFEe/vCM+w1RwXqChtQGYagVcAye+B7Et2pKbi1oQ/txQWZdBsLyocLBxJ
ihaGEiPjtBb3HipMkBKB9XI31zN7LXXIIwgPWLcbN4v9ZZ/+c0VQBlqL4+sFebKa
G1KkurBbz4HMCdKytEkwjLK/MhiDEgcWb6OGAf3s5zBjIu3rbpxMJRWxJpikn040
f3DGtLZXaAqAgmxYNrjFNiO0hK12YhQa1gbsrSZhaAebgSmUFo1dCrXCbZhyNhcy
XG9XWr0cxpJHY6L91ZvlwJP9zXkOnzTbAy5F+8mx460eiXMYXqoxe2OqzQSQqCB7
OpmDRchvUxlLzeE8yNN+67rOHmo9IQyaEjUN4X35wXSrDclz3Q0CeaS+75okOp9g
kJEa0hv5Mx+t6tygUpG3tp/0KjLD1/3uAjfChUa52N5RzkJjyjxXbyyze3T5Z5Yx
CilqOsooC2NlZHy21d802FCNY6b4aYF1qm0OYvB7V2rfmlDTZfI+OTHcaOvptH1z
V/wrP1sVTmED/0HgQATEexpWl5yIOME6M6Mcx9WbfUqlMXrWFTAnWLE2Wz892fa5
W1YbJzliRLkQpV/shAd3FGfW1aS6sIHkx5iWY0+c/U8Hpa9roc3ZN8hisQzpZL7o
C07zMUdr4xL6pWQQsj6uUpPl4W2S7xS83o2JnHiU/qDQNV3AnDFMID04AsFN6+r6
NF9/lcqf3qwJbv1Mw5Oi4uVWBi0h/veL1jDsixliR1FKKYXSncjGuWeiAT2jfdg8
nE59xul0X1UBK5NqwmAdSW3Ag39aQV/LuaWM5b5LrbO762R0jgmbS7DopC9+054W
LoO3jAFRyYLDw4foBoXAxVfQ/wBjdogKmAvLjAewuU3NFII7DVcWYdN+Gk7vUuXT
n8j5X7gAt6hrTgC4e4gp/S18gSCGvEmjV+is5qjz98glmtOCi0VnjtRPXKiEqLsR
Er+e+Tu9/cca0v9hd6POqYziLq3s6zIfqekxzq4tSGhEGUxSR5lb4mlqZC0//xXu
znmFDZ9NWtoawXGXLJhYXRW29e3Cn7dhTVfjgxGlXd/VMnfOf6akC0tp8D0WeFlL
LDUOaEiavvL62LdQODaxAdR4z14KHw6V9Pvy9ADNN/2U0Xy9S3Y2zWk1Nz/rXxP4
fEG5CJ0OoJIT/eAa9eKwXSiNoiO5R2e8Yv3vbfi03iohnlmi+76EMV+82PbH5bnb
Qk4z18oSPzYuTHdrdAp8y2ucuMfyqsAckhNOq+SBTtXQMQCsPWEtrT4yuwN2xren
VKw3f5T3vpwHofsN69Z/7QCrzn2MiXEfEd4ocZsOzafNH8lgcf68vCOFfMs+qW6r
9IemWBI8e1Kyu9EYMtQt/Sw8UelfpqCCuE8hZZ8PQ3krj2NefFLZpJgHmEsN1UzU
Ic7CZBKu7vNYDGi/oLeK+1nl4rdSZMzVaS3YTptahgYleFmbHtpmLZcpv19w48SK
NwCUc2LRBhrN/yTCB+IgvS56gi02chsknlPTo92ARSwGg+XVxZlOFeTON17Ex+lB
Qgawly9bCN7mPUWwo11lkl8AB3GQ3dD1nE1aKL6+QdIJYRn7A66s80gqfWld68u0
k/08HuXvwpS1jN8PYZP7X1JbybOiReB0WXAb2JzXcZCWTvPCinAr5eAa3quXPTuL
uQ1MIHMnIQx1hPAB9PTZDgKbSdHCQQsCuX3nocR77l8Ondig4E5ND6TanKplpZ7d
vB5bqvfpZC9zemxj+vvQcbAxsTWgAi869w6vIJsDrXqYvZRzhGiluL/Z6CXiKmhf
5Z+yS8F0arHJG92XCjEnGaOux1GSgTNnfoU9KImfdC5aJAFqdQwhJnnAFrrpCkoO
xl4vf+1uM5/hdBB8wdIBNHjthid5tgg/H46xLZhrXPP0di1Uy5E03TCvkFXULJJK
N2r/abQ3yPDNk2TXEtcG8s2noxH1DXbBJ2JSAWnQpOWUslWW+ILLA0KiNOvbPXI9
gTmWI89xwIlACyztqqMh40Rk7N2xNrSbG4VAenX1GtlBY2+WPuNVpsGsoYCPfQ4K
qGYw7EXQKWsiye+snvzQnAeeRomJdyRA44LYfKW97NgUtsElQxcoyXM4SjpGlPQ/
sLhINOiTcbchEw0coNyTKuj5RgkAm/+OBAAntriY7hGsLNgBX+wVGYcTJA8iG7Vj
q76QEX92E8VuxvxroBhjcPw2KvPh8kE5sFUKCjXpdi89QR/tKlEo3GWjy88oSxtR
xlHDb3PmpOZ/kbXnLfZPDnioZqtFTtGDGAUXkJZmsGpqdL+50MhpiFJpG248qKAG
PfGmJS/97yWAQhVaFjQnNPNvOOI+R6718Lr2X7NO1FXTGO7XFogPRjBYf7bw6klS
XiUayv7X/jcdg9FN3+AR76dtFQBDzcGNVARPSfVDV5ZJ14RJhwJM5CdSbTNcZg3h
rYh1zgyxfAtm5Sp3QFNSdOwgZLlpMaEmeM78uE0Veg1LNE+rbkjL80sMCk8uIVoa
Abjajz44uLRBZk329f3ewdSnY6ax7yYpu96r6c0FoD9y+WUcuC5ZrQNgJCVCaXNQ
/bT5TQ9bUaTUFHAuj4uGw/iRLeYmeSz53WLT8vVqR+JjL3v342WTH0Ztr1Y7r/oi
PuBOuoT2amum+OM5gQuvbi3xA+tF0Yf4O2MLnzEnDTiCpphAOwW09GEK8m59NQLW
AhYErf7fRBMzNEZKUoLU65RFwAjx/uWxKBr30FDRzmNiqIu1hmq4Z54VCp+J30DR
2JwsRhMHeR3A+V+Rh+H6HcdjwU/T8j30rLDTnjEz1xCd6hHpBwHHNwcl1A8lRzNo
bnQE/HjPtjR5EFjBgx/nhO8PMpT1MPkbb5WLlzCJGW96H1Y8XlcO/Ufa0yv/Mlu+
v2srtq5hE+JCjAzFfd/gffqeXjpaPKlI7WwTOxNWAfRdGN9yxbC7sfztpyUMV+Q1
rEQ4VQOVgFoJZSVrSPY1CL8ws56P2QQ9KXYkXxXsfZVokB9LfpjejXq4OBehsP4U
0rjBveGhkmCdLZLy5snlKMrGCaaakogQqUPblyUEWdfDi3ucvEIfc5yPgayMnepZ
CDeS+9AdgFjD00GtXr9Gy7nCiEU/VU7at8Nh0dycfFmmuiVUbmAOlh9DCaEkXk4x
8yfgND71YZXrI2wCj41I2wThgS0zWzZceDH35/qpZ6uRNivgvGQzTPpxKe8rZnPX
A92QXHUtqfW/zuFpufeQZnW1vqkqfVKtSQhekpEKk47eXN3k6DYbAwPDlIiTiRfS
I+Uxem+kxpydmD8MpR83SKwHVQk9a+MgvxAdk08G2jgJ0Nz/y5ewznR+HLyAQQcl
DnULjfpVXi4COCMVa19RgFct4+9t1d0AN3bk0VZGEAXmGsysqgLtwch8Sua502oj
Z6Fznl0mT6XDGWYOI2nzrLGHXqE2xt16s25op/Xw4KsP3Ykouqia/0ezO+qFZTWV
gDtp92UD7gshKZ/2shEzwDUQ0xMOozZAGKHUWDJi89aoXXIhltDzBvL7r8cmC3nY
q8MHLuBs/n5/57TVN5dmTeRar6JnYSXb13rcMMXKg3KFZyxlN+SEQVaDa2SZ8Iiu
G/Dg73AwLeNOl+qXrS0YkwAnKuUg16ZhTi4qXs8jLw4Z5FSmQluZ93K+Xn55Yhga
uzJg17ChwVhqEcFcO065QzRC/9vOhOAKZFaWEMzkBrgEGNbS/fRo4i9hqOszi2Dp
1SBXU6tQhIk4LaICeVg+Jn10ICydQtEomvXcxdJOhAJ6wdCi8v3FWpzYa0g0iGnX
2LaFMDmxh2xir7v8kAEtc/FBHkGlO6dPErUgdGK8d5sUdk3KOJOwTvIE5JmYLgGb
mzO0ukdxcRNxyvB9c8LXrBaHC/sIkc8IiTQC0zw3ZS0tLWoWOh6MtrakpN7Z54AV
KD3j3ZnECvro6GcIrSJlGrns0vRuK7EIpwZe6XGMqcVXluey59uFRItROCZDNHEj
xEbjooCQSk5nErRAyfdKB/ydNUaIOoi9e+yVuyvjG6UPfFyAC33y/nAuovS/Z1VM
P33EPl16isSKx5d8VybPJgC+1z6segWjk7Wf90fJrhoml4VBh5hssRZzSuUKbeCB
DwJsBA73x7r3uvwIjs+ElbT58YUc8DRmFJmrMr386xd7ovWL4CO0czuDPVzQUPNQ
ZPzvtZK4ZCZpwz+4FqUSKWG279AOlicne5POH7LoEgK+QuPvmRylF154JQCbz3vo
AgmjTxpiZuPvhybJuq2iJXj7eG6NRIdYuBJH/epd4CQcmSQV+bZQ6n8jwVe+72tL
nUQbKYKQg8H+EmV0YQG6PGaHukhgXBKrZntOtKsORAURV++JTZ2Ibq+GYCMdC4j6
qh0anWfwZXTlk8PoUND00GJVGJTdQvs2ZKabzLNmX1pepYyzmthbJOEnMIC3O68m
MfSFBrD3wFxdpWO9wx+iDlV1yXMD2QBRcp4nj+f2gazQi9freYKh9fSgHL1qw8kX
H1X7wNeWbWVplqwUrRUcZaSpHb/Pu/aZcxO1ZedDP8KHxi0GA6KKzFg2XUoIfStL
rqemupY6559Y4raAiVJKGRUKnR7ft5acupG7KC3ti50YcM0X9bYOMf2IpCOseXta
v6D8957kEBKgDXdiEFIhvRjsvq7F+WOR8RSwsrX8mpJP89yFIFs5A78rYWtuJLRZ
nqi00tgm357DuHDWUBpPkzPBimt2Vdrlyw7RP2lhONj/tbLhwJ7Vx+rMVvQ6TyfB
5Pz0YKSya9T424i0XW8Ui4zo7iL5TbGZeoprIJSyhzyAV6nmkMQwq7ac3uHphsCR
ahbf80y5AfL4emrj3fatkJIuufx2HTgaFFNLo28hjRlsjTnByfrxfJeLdl2edg4p
IouPR3uAhT5Wy1tSCsFE8/Eurx9dZSFnJy95BmR47HtJU8eZz6v3WeHChhICoAkw
7YZd0RaiU9X2E3LZTCe04rzTu+FAAy+bdsF3OmQ2Bnic5Zn7tbxKXYLerktNjsiT
yLu0NE+iF5pvYKR0tYPzvKOjtzERxM2PzFXaSS+No+2Ozks7Z0l9NwH/ELtb+t9a
BmLA0eTedGQXrg5H6iOX0cDYlZzCJNLlkVk3/AdMIVi8hDSWPkfOlokQBGsncAun
cOlogpuIDNrHITYCCWOn3WAw8AbbmZ8G5nxhXVcgqt0hKC6zC+rdqwmmVaRkKZ7L
Ann8sadvvDmbC3Hgmg/0YxSx5+bxpxuvIIhbSvbpMCMKAVJpITgZlTg+rlYw2Awj
35fgYdq7HWKDVSGQbbOCmvTUMQFFjdV3zFrga2MBbuCel4XtSVTnhjqp5GvAOblG
qVH2EmAw1OA2O1PWFirmMejV2fLXZc4VjW2+gYUwuryKqk4+eMqXjfmAEp3ScidA
ELtcjLRi59heR4nGDYsZMT8stLFG5k3sza8mZa88v+oKXGEnNtlIKmw1XKkg9of6
GEI0gatBhcjutli6XhX/wiBuyiFSTovPsz4ajhggfXoiVHUtnkp4Qd2sFX5X/oxJ
Rc7MfKL2Z8SFq2ujZgkMpSR9RpgoHz/J4vWAVr+pqNH5RXhYURhcnKq8k4NyBdLB
RIgl7Hffva13eASt3054CcLBq0/rSd6gGd2P//2J+l21ab02v9vPv/WRzNcaP9XD
KslwsrSODFLS7TyTrqhTfmGNLibUFY1HXJS7IZYIHjMSNrkl1TPw9yQSaS9E53MK
7CbMKSrL20Zx2nMTNR23XZSwh72kQT7llCUnKHNNpnby2rNykhxeZDLR8qxHvNre
UwoJugUoB0MDAg5NYQDBlbdZ/QkFOB7xaCFPTbn/TFe5Pm2PEGKa5jlH0NAgD5Yt
MTSkLQjwJavlJsCycQmL4qdqfAXKzGAtgwzP0sJ0gVSUl6O5Xb3xe1ZrMqAKx3nt
+DMzWi8KabPWk2X8RtSItYjSmh8x7kaF8Je6/PJ3pb8rrO1xqxS70h6GYZazIS9E
YzX2m51Ljr3BOI74pYsKZ6xloep9brQjQSdigIeNAD/cB6ZJ+PXSkqM1xDFPD68W
Lf2fydCRFsd/soqnn34ptQ5xGsYOYzYfJ9EZe3LH2nOPj7Y4ZakhcJl+TlW3DyeZ
YNexsOgeEJbqK9L5jgZU/IvvT+/XknoDsp9uTtK6GUoxKy4tuFb9qc3Gz3weTHSI
uoKo90OE1oRwZkNVGCDlATbId3q4uwlL/HdL1pYvupv3VAW1nhlb0FX1C7P0Fsuk
MPUhRUSwjHyGUPRquXU6/py4murk29OtCPWemso+a2HNVWiJe7I95uS1flm07moC
RtC+RcxaC6iW56RZKeN+qn5oN5LMcFCIqDHH+q6lHGm+G5R57563U+Z7Lh9UOfgm
RKx0IjEDU2s784QhYEGcNkGZdVYqb35eG7QLprMyruaaUaOY0as04sB1wxeSCa8F
H/c8Kys7lLohq/jdE2iOPwf84JKQO9fHmrtblsAIf9CqbuClPo+Lmb/yM4hogtbM
1Gz//eoa85/vwT61iBA4dBSdINdm2DWTLMhwvrVInazSnWb5CmisN9qkr2K/cvg4
2AmxWDHV3EsTjB2IkMSy7Xu79AjOMZvbR8fzCebZy5ECIyD/qGu/fbfOxFVXaaXc
xzTUxwDhAljOjm9vYxLdyB66SuOxZyxN3xxwvhcmwYF+W7QYW+CqF9QSa0Zniu36
5M8eOe9ImogCAAGkPdGSIxcKGj9zDB0oyw+gC40CJO85aXAxvok6EqKUyqwvat/b
gjplHU/EkByrH9H3bQV2GHYyGNObgJgFMoHptR1u1FxfKWwCeSpIBAzZPJ6Nw4Fx
8/LgAj3MsYx3td2GaB8Z8sDis2820djdQvdnDR+Sym1Oi8AswliJlrbjPF2wmlzx
GSHeyYy+s34s7e1IAiY1kd/oWT8EsYHyJgUjErfNse7QOcfJiiK0InfRJgqK8QhG
sgYIX3Gc8MY86cPIMmbyTH2IqVHFS8aOL1DdQopNPdnv8DdmC6Ct+sBP2ChuYQVa
xpm4HVJz2xbUt3tUIp8LUYTzxrATDMaf5JVOqkpdlHo+wiDSwWI5Q39Roiuk+g9r
oozHhpn1/M+oAmGenThMxwQLIFR50CSbl0meJXD4u5NuzQLl911VfCuR95YwIvP3
pslKS/LcpUt+uhufU2uuwHp7rM5DgPzwFkFN4UmkJl5B+49kS03cAtluPXYo8Bnr
9KtdXZeUBYpATzW7GrF4LHFssjRUGfy5vU6VxPhNvup4LjJv588X0RFfNzPeAqrm
DE+X+C0CVuROhVfWT3IG6HnlKg0R8aAhtgnHqKptNlgWKRuckwqeNGHGhK2i3u0Y
VZ0xtGGBdb9p+GIuXm515mVfqH3U159HfjUlOfRoIutZcM5fHmtFoaZwUe15YFFe
jFR0M1oku4yUq7b0QFFVnOAT7FSfnWfNRdh7PCNaR3UEgFmpRsZYzinx/209kRuf
sau7iJ6Bu5XANyCH8y8gnHtcQ1lvlBTmnDmwl4h+hScXbFJXe2z51rx4DAHoayxg
QJ+6BkVddbhtxvM0Pd62QpqLtOdHgQXCf5kKJBnLlNxkuTI0/Wwu8/KrRHHlEUYl
Vw5ZfOHl70k4dH92s3IecKlQMaujwr57hXYrdMy5yz3NxMtF84/q40DBGAfeDpwj
noTl+yhfeAgCOvu5Nlqyv3e7oB77zUK32fU2yLd6hHe9dIESuVa1YFM8tkAct6Go
YD1P7djm2D5kh8nQ4DWwHAmMjlBJOPHNcEJ4Bma0vgc0TJ0cXCqPAZ5N1lHJf1Fi
465dmgOS4zB+yg2PyXuVE2evQGIzxha60Jk/4gobh2rbAYnsjfouMEHasApDcieG
ZcRUvygpI1uAfGBBfrWy0ggHt6yJu0Q6UsSSy8cyzOH54nxKC62QpVuQZaUvydTz
FOvC7hd+53zaygCHBwgOUytsuySogvxP25vv8Morf+7cHvYTtJu7sgm2w58hoN2F
sMoeeAvKvnyEab0U2l5JGraKsmWkJSeOokGTuEkghfmzjo+Epu6n58ac1rsA4Mfb
9LS+Yn03WUDo1IYJ/KyeAL9NyUcr4K1RlKNonJGUxxm0VwiTqLhcjF/mID7SQFjz
ujwm5w6iDqJ0BF63aGayc+56jx3qwf4JU2lojCnfvUCCKkno5/ZK3kWtEocTG45F
Q712lm7T62DhAG5DiQzT0SQrIhyPnoYf5BZG+B38lp1c8kiKr7uBAk0kTPYmTi6o
cK/KbNBgCHuQVwQRZSAs3OyY3F1Gigak5LyAEeZYgvYM0hpak6B0w4tG3E8Mw21G
TXs42HG9nP0OtAE8C+WYJeclRD50/Ub1u1tIkEbBwoq4zVcmKpCDMwmSgFUgRLWF
Dgmphz60EY2Bve8Gfz6aDDuzprfhezH1m+2jjWbYIPoC4hwc0WgfqNEN8r8PdkUU
d7n+GovXSzccGXgDtt5I9kSRDocIrPd416R9TZ0v25RMQOYWnuSOFGKUIkhbv9Df
XMSED+mH0yjBJmXoXqBIFe3i8AeWZPyiS4olDaNLMws8n1Q45TeBKQWiaIYkg0LK
epTQBu6kSAxsaZWn0/N5w5cjFrH5uj4ZL1rqiB/5978Ij7e6fI0X+CzhBL1le/ZN
JdVwKgqOxyCxGqDPfvB9dg244YCqJFjP0rYkNcbG2naPm9Hn039xJYcEK6bRdh1G
RCZ2zzrBwKaQbCYqaOREZ/Etc7zXy+k+2IHhdL0r/OAHMRu+inUPGsqkexGJu4B6
nzbHe4sSfN8leau5n5ON2rR3y8ygpaUokC874YxXj2Fb/PBES+SeK/L39QRw8dQ6
8ufnu/FjiGuR+SJgTXBXlij4wTwyrAzcTmHrvuPT9iB36PHJk2DCJOP5mmIwiB22
w3mfgYJILBDmZh2jBbM4SMDI+EAUOd+O24KURxqrvgcYLenkp6I9xItAKWooirkd
AIrhFQGRlaViSHKgnkwODAFE7pQZcAfATFLgiXvQC+M6CyvvqZKNwfidxHubfBT0
QxX86YuB311n4I7lX6xd90hOSW5lYfsMxhH0yX6Jqx6OuJnDsUzq/ESch2h9m3b4
yDbGOiVAQE/F9lOVQ6xGPreB3St/AaGSf3K+r5liK1y2W+PZg/x7Snbcd+1Jsger
ENNDmKhWvZXQzwsUPPbLYYplzYuhVNPPVjzTF2qdvDXr+oK9XeWeZOJQ/I2ftVVD
2bJm+PFzSQlsms+0oHMYiwwJiBoe/hcu9FH4tR6lcVHgQRxDPgHAQ0NOissSum35
SHe2pnh4msvnKEJwPlDix2NARfmvSjEVIShHagrGwYgEvehUPowatSR2qk2zUN98
Id3hHHvnMZEriC1VBGfZYq2rDTdWk33ALa6qIiHuZGJ/or66JR/kBpqw6w4OznzH
xI4RbeXr6xNzH+QGW6kB9XtgVG45+vOOmxkoLpUSUeXZymKSSFyLKRPhbTL7Teda
y04JQE/0vmPLP2NXpvbGCOUjeKcx2OkD94GLu1vxTDsCZkPS87rTlvvahfs7M04P
C4O0ivga7zinSQJ0QnGZGoP8PZ0URJ2oATzqsKBh2G96pKVkp5sRYqIFof5Je3Bw
pW6kA2wplP+mmfrn0rJI3tdEs/7RvhmBRXAt1Ybi35qkY4NU4ZXU1sWl2cXt3ChJ
WiFtGZGyOTZgM/jDw98oW3whRbR6xSTSp1bU3xYpn142RHPTB158MJbY5Peyl9Wo
DmPa1QJyQ1GxmsnNsHfIG8yn404otEuvN3pGIO9AgHyKrTqMfSBu1hZYr0SPSDk2
avB7ec7a2PiQEQsJTHGiwscBySUaziM1hf8jjKDFOFQG6VbrQGkIECfNdeIetUid
ffc20wF1gYqdzljC4IiAxxJCVrR8Zi7zvpZrCIzUqW/0U3qaLmkzQCK44Tcy9ECe
nWXoVd/8AQB93ecx2vu5JuyA+0/v6GfQKBSp8Hbh05QEBH6ZRUUm6+BGNdZJfADX
6l0N7fYEqmJRyDuej5FmdaFWkWzqGy44KhdHl8Z7zE94y0TyV6e1tIwVbkEuROvS
VRR9qcsO29I6g/VVZxe2f0bdZN3MBCH4by7v0PFADR0RYsuXh89FT347EjvZTInA
mc227wwkUyJf511UEOCCc3VS4P8//C0Q5X9BVdoDk2Y3oWAyWn/iRMxU9riC8WDH
OEkMskVcGWGjZjcJwHlOQE5f8abm49KdR4swu0gpUgTS218pTmDZ05ROLQSH4nyr
+03uUAMX1zrh1b5nQut2CZ09H+2GMgJD7Ac9PWxxkfGUKyo+kXbTAvSZgySbxOWH
m/rdN2Ys3SXgq/n/zFHyUU1FYOIZh187XwaR6HhOzSH2VdPu2tKj44goT3a8ovW+
7So7LTNIWUDES4W7cyNBh/JB6IC/7QL2F5PMQbv25Ks1RhGL8Rx+CdIsPeY9S1mx
oMYAi8Fu8oI6c+YdmWUN32FWVtn9Os7cMtsYuAPHxRj3Oz5iJW2EIxCr9WqvtsAA
5BV9d1cW963n+8EtAGFQ4+ntEDVX3RpWi+XSNCPSAFyyJwt6zcHGokkeBmuzVnXk
uhmH31ZEbnhANXyKD3wCpqMBFerNetqqQXPs/50RCVh2pE6bPj+GXkLbDBQJ+rxL
aZJL1cFOXdtdIExw2MQnXK3oIl66y1fNdsyRzt9apnMBFbiVMHs5pwjH25rMrewy
stKbCp9q2oKUHstboQb5ZdlvBy1ed+EUgTadrswaxhBaBdsoaIj97dd1cRj/wOr0
OfrGAvmanLQIgQoRecZkp+NyDF+xtEmqTTqx/UV4sENmEzGA63bG1McyGU9mCw9S
7rdg8sMOd8mh35l4MynbZQ5O48lRS7l35MA03jF5ly69c+b80rMbyuCsdW7i7iFG
S+xR8S/KX6jPhx5Mp64AAPFskkXsSiJHY7UD6LqgyUKLGe4gavD7VFr+PAZo2HP7
pwPKdnOpvVZIduKfGfrMACxWsfYiQwqKIFzi2ZLD2KyhKWPZRekiK2erxeEzqMT0
l/3DvIkbnl6CNW7O95FvnafxcMvPoz4aenXMPgBIh66aOIJOcdyDKxONh8iPeDXG
2MQq4iRLcJapatCr4PPdvfs5jQWq3HTxb5Pvd75q+sARXm+KuK69OmgY3Bx03AkG
Jqlu+dK2AqNyUtY9YD0FLkBfNmmLfckruibzmFx2N2AUkEY0HVBk/4YPI9ohsHW6
5/HEYBg93mf5XEK9aa37k/uBIy0/C+LRcy8DERF1H47y2bcXZ0jU/Y5fkrcIMUsV
ZmKdwytVWvAJH+XJ/yoWotYJLuhSvo32lb2OV/E0yJIGofMopq+zV8XZxeTE54No
JMhRIzWw1hEoiZcuCE6nMkVNnZQ8SYJVp28/m6FUpFmP6H6N2UL2/7HVL7kqyfuT
16qzS1VTxVQjRJ1xOjSPPyW7B9tYYo2zeVUII8UFXZPm/MhzzTE2jVl3K/7IffLj
VmPHwdYCA1kaMLxPCywFfh8W09H+4nQPOvhRu/YKzwxiftLqxFFITuI/F081TPA2
AhImmVr4DHNm0OABowIHOoY9eZhk8tLzZXxAWP0e+q4BzwqbEfZcbU7iESQScx1O
TwXiDOqSv0dxxpRz/uGryWl1acca2irLAP4bm4rCYZPnfw9k1D5EszGuA3tqeL8F
4J02uvoP/6NpLFt7IOF4WI+yPBXkl4JT1U12JWM+vSCnA60+mmiZqF5JargyUD2a
oFnPBB0zb01NIzwfpF7wHmnx0xetkal/uISziGW9GAgh3S/PunCpJEoWqDvjDltp
+TsHV5rYXeOj0JwA6GSNMvatROqHVFayp2PJpEaXCuqfDPTj89B8vMI9mKTVDe3u
74WNOKV9bKw7tZySRbXZsFm4wDkaktfbf389zrMe/4xCvr0vHFGNS3Cygu+yLu93
7VRujkbtdV4neoreyuOZuZJ4BddV0g0RghYPt6EslJE+P0AhqTy+9zQoNaOdeXhs
YnNSe6Sp1NsrfdgJn1Y49YEG64iO8nx8AlQkL9D7rBHe5BYn761fGcc33mpTYqhk
/jcc4zyGlmShi1XLCBVV65oGOQo8ICDXQv88NESMpQ9lk9P5gV3JzqliZ8N8CISk
DBaw+sSxxZKGIL2U32o3Jk4b2Y0PJHVBaW2ku4JdPpnWJ7Q9I9m9rjnqkwwaiz/G
VwX0YXfqzg2s8bnRXaqUYTzoQj62GcGx1Z4WXHAfInP9PO/QghHSdLqpdJcLwraL
vRaQs00UoPjra2KSMJV0HHJH6iYQ4VyKpfkfhQhbqi/9qk0A6k6iAaDQ9ZzVx8+b
4EWcKdSXFwcW7lzoed4AgOwbVWh8U19+d2viNG2MIobFKV1UIoM/iT3fP2ZOpBqF
76IueyrZ0IWofQly0sDVETVEkiZjtF6Kj2THzVFqPUtM23HMkLg2+WQXXC5hGWGB
5QspLUstBeEc5tgDtQrMQShERZZMeFlb6GNpXacyjTrNNHoTBz88ttHoxxMOZl/E
wfRWQJLix/EDyrCwiATY3AXZidVm3u5rR5MyhYNJPQTSk68C38odoymKK0vOlsUT
Fw0bCyWg6NlQIMNqG9eK/PzkjPlWG4u9MparVKAr3S/RLd0OkfKrG5nYxW46LJen
Z1FBtY4DUirc2Ii3n+t8R/UB3Zl+pTGEeZvE0Jqlsdyfyw6bQaPk0DjF72WcvHsO
N9zjCztF31WFpDXNbe1unY2VpOm6/IA9gb4SueXf/ZDY1vB1H3S+ObgWWMZREvS1
JqlBOhpHZRirQl5jqI9dT6llT3KA5cEFNXagzfQn9rKTIeGxFp5R1UG/Xs2bfz6O
E3RaKjsU35mVYMzI4vaoqf9+oKDQ96seVVOtsZWQxU2DgylMinjlBy9jVGVUK0vV
Iek3SzQy0d6JqhYkiWdeyDE4GA/KJ8pL5QLe8oWemThn1Z8AHJyTrhERBrlSbsrG
wueaA3SgmdnErDX/W+yAtLQPOaTMd68caBo4VvBA1macHwZdqQmPU0IN6rJdc7Ir
YKAV5p7CWfGCZfC2VHt5/BO8FhK9nL0tlkC8fFs0mrHDlySZlPqD9bDsLoLzpcfh
zbDMCKKr+C2xpagqXjCp/ylPMfd3PDOcvH0p5y/lwWr4FtjKwpaEShesUdJyhW2W
a+u9LVWqKlCCkK2Ki6pACB0Joe3eChunrk42eT5jzi/dCQJ9cQmiKjHrL4Q/KLNm
pnIzXESzbbWz7v6LLjcrW3NJmNa9vX2eJE7mZQUUeV9w5tC2PVcKizOKtzZsck3q
yywwZ+1eqh2sXN47KjaWcvTMtvQ441b5yiJac/QkuZdYXLZ3Sy1WxUJsG03GO+HT
yzbnnKPYjvCwE/e8t6pb8d0dzNcAtdsrDXWOtEDkWF69oPAUxzF4/v+ocDKKW16E
CaR6NMjK2a4gZsnshtAHcBPUSOK2LT501IK+Afz8llQbk68fj9WWooUJqSfaEvza
rCrCdvQFd+o/iodXuXY0UrlWYakZ+QV6yxyIdcb6OZhOpyo4WceMtvPwKlX6vcMK
QPDIRtu/pOZoeg+UViPWsaWNlGfQ/7t0BkEqN/NKpsDuD8mYaIRhBbcWieaYKfca
C6pBnh1Bm74PTgY79Pvd9XV7wixPtNdvE0VNuu/GCT2I0g+3qMeVe2W0DeLQfWh0
Kqw8KWgbkWp9SwS8nv7kzAfOtltYJWfK8y6/YlcgGBJxIxnmGbI0mSm5wTI2m97y
tW9vTzLrfJXAtwnMpYJDYvKJN042zvxpQGVFcglPFyHrrbwUmATuXXXQ7UyZeckn
BoCsW6xk4Qnrf1RdHyb7sF6jD1JAuGzWLIUOphuimvWXk0bltxotCnf+wFgDDWyd
l0EMB3wF0tJY4IzSc7Rknjt+uVnHq8MrVMnBeSFrbiqtEMN3iLGGI1qd+SS0qBDj
fxb5HYN4PLXTf4U6UGZsdyGx7Y2EuWf4qI+9wNsWxkbN13IuAGgwtYivdV7lWh7n
84ObUmv6n3aIRkgdaIeLS0Wh3AhceiakbdayaotRP/fXpaP01cXlgW4/sOgYWcF8
MgCU99sX/o8bDY4+FHVplinIMbbEToU1Cs8OZlQOJtLQNGpdmidPwsPeQxMvNVHY
YCQ8I/vLQFFb2PqjSd+AHxX01qYgrP2TRsFRR+EplJu/rfwgwQkoJmnUa5Rkr2gd
sNw+csTutBulEPAbT8bDFupP+yxj8FrsWOIs4i3YRoMxxkt8Re6QHnr8DE0bd7IH
4222VamQMmsxYiccK1P4H0gWSNd/i+TpUOphNTIeQ29NStOKE1G9IJfzThygDBoa
wGQsjg54noqK2EQ0VPcsApXvqpG9T6jH4SnORScNmEJgUUqk8/3q7i1xHPwfTWuj
Bzs2eakxcaEr26AUlxd2KB9k9IzrN72n8rAq/6sC+bHXEUGdYEnFnD5sGtUfrSM4
Qvz88AaPo4qac5zpVaCEoHP30UKTpgCo9XtzLpLrOcBubKqF3RPet0Q+LZgRpZBB
3wIUpmdS2iq1nnHRl9Rdg37WJFIw6WGNrr3Nz7uzoS8STLpJ6hXDhyzRES9i2rMp
0NgYofrX83X+lMgFXsO089mwCtd5TokXP5c5/aR1LuNAQKq4cuxN1bFeWDw9Hy6s
7CHhQnn6hnLRV5QuFoa8IfhKTgexSku2/cOWUPGQJUBWz4AluoEegW5YRIIrtamp
HNxqORo7fYGM4UNdzVbdkG8lX80Jc255yBJgBn9Rqq1jwCNYxjPrshh9F2dov38i
8qLAz3VkCKDH8lBrtFF2Kw7DXaF/zFRMvh9MugJkyPlndaEXDXjC3PopxYlV1Mpn
XTd+rvDWxKzJlFWpzcAWvTXOWtvASHXz/5Ts5SdKeiN7sg/YGggtQYaQqitp7FTt
7uggNK7XNwDo+c3NUDSF8QPQvcbkhx/7Or21Ig067fZgmaeYcZBBQ7pnc48OWPXJ
DCe4ItFoHNxP9MZKkjWBpgJ1SROqprXoEFVyTzhMvD5zWr/hNYVoCIdKoJC+lZKY
AHgytOdGcs7ednvJ6XAY3pgKz9N0L1ZFXWO1vmJWOh8Gc6K7KJIBVVjvtr17cqpb
8NJsXiXYiqbo+O/lcCTKuwTm/dd25kYMyLFzXMpFehpVlMAM0O0NW5mjqiy7duV6
vwIcwlUFBBUQHPYycoRpcoMEzCwVzOLIXR55bB91el66pHbzYkKXkZZ6redeB16D
Yt1XE/hxk0OARETd0nUwWNcgW9LC7BYNV/3+dghsJ4K01NJqfJ3Y22zz39JyFhQn
5o+glJHpna19xqhi9PkIzKJIDE9x5N5+AzXIvE5KRy9g4mC3BrOPXZWM1Jpsahis
xZ6fl7JeBDKH4Y/ASGDtrzT5FEtU9LwKmAc6bRbOcqhejJ67OddnXrwDi1wu2oVK
hnz7iVxZxDzIxYhQwB40gwiz8zVif3HM+9pAUZY3dk4Up0TheYfhR+WeC9IdygSX
9hRoTk1mJWkyhEtqH4KxPO+SBj6vlA+FEs8GF+PB76DUa23XViqRyAa6lgxXHJXr
eqICkWJ3FbD9QhitViu18kIqi0ZyyHiwIKAUuNU9LbvRJBz2x0mT1V5qFCjS5TQj
t23PPaMDpQ0bIc+PW5LYVJUBh0HQWRkcbTcSoJxkdgAPc6nfi1yQQuRikAatmA34
zPyWqNPLwATQcCLfHVq5JalwYsymqv3GkHcgaB6haOJ8VKUfP1T6Rd5gqaZthElF
L3wpRMWGQ2pmtJm+n5heBig6qCJpO3B9ei5ZoLjW6yasBaI0DWKAaepfD6gKLytN
B2yxr8bITwvTSMVfHUdAQUDCyc/gv01bgMeR9JDcfU4zTrNcv+JV3vnpfy1mMYLv
g+RPSGRuk/KwM+j++ktfsDuzIEDdfyopiuRp3YcSHYsuJZ7P6eX/vC2w5S/MOlcC
xfiVYwvJwE7kyOsJhPb4nquJifnvlkf7WE2nmxts2Y4WL3zN2xMDSUS1f0ySVfwU
Flbb61raIFdp30fiLKr7xmp9Vj474U6U7QQ0FLnIilTHCtYEgtgOFbtL1XXthMi0
9AwCor6/XdBjtFx55hiIpFcxeTJZW4AJRQ2pj3ODQ6eY4mQm8vcoBHy/JEEnZv7X
oxin3xyQY6KIVDzxtbw5EPiszsR8hZlSgQvLz3wMazBgJ4Cpz3KPFujoL3jGIfRh
lbfwnZGZFGEMipKpLMgWrhCI9aaGdgWzY9iBD0XCi87uc31Sv1pXX4sSK9guXY1r
+jw8OEiNbMg193LazlMmc8oOL9Frj7EHhCXmA1OMrBCYsQDsWnBeWSBNkiQPwNa6
LZ64I7zLnrIYfHdBb/9di/x58Qks0WIZnCrmlwAP2oJ+Ttq+U1hAwZfPwWNUaqaJ
4qAT/+5idcoQM+gGX4Nf7fexE7D2sqEQZxot3fwA1GeCiN4gAKo6qvMi2Li+B4hs
U3Fz3t19wlBcbe6eXPx26zQMRYdV76mUszCKt+2g4GsItcLwvVR8CjlbgmhyGnJr
gxA8gWjIf49WCfjT4Q0iOI6EIt0c8Hln6IPomAPugkKYQkDG4oXlroWjnGZoz4QK
aQRMYJqmaYlICs5Ed1HLQdTCiSgR/TeUW4uYlIe+SGU3bcd8Yw6TzxHji1NrO/W1
O/2zqgkyDptoe9/t0NwmwPl9T021FOIGY0GBM4ZeNXknqLCgoUgATWsN8cFzM/sy
d+i+2sjgwIIICbnsRqP+J9uKrYDiyaBY2Jh8E37vjPrlzKyhvzF0n6YgLLtw23QH
6TPOS/VHlELlqvuZG7z4JWNHuAgcA4oVVDRYvfeweYirdoJlLdULnrXjqulVXCk7
7ee8gMzhtnmn4Ry1m3KAAv8+Q0QhNftxrIqQ7o94g3oJvNfml1KOazP3E5iqPINm
8Qk2SrZTM91/LADgrLN26IMT1msRTHL/UfS1iFg4Sd0rYlmNRpjAJl4sCXVe4jSt
f3hrpQTcMP0otCxUyUlF0wmkzpBGXJCN+OTlIlEmjSqWxMpaHcejJbpPVlJ+aY5g
0fKp2SiyR4gL/kZu1AHdrZV6qfL2xgkr66avmyZlbxDM7AfBt4F9NZ9dgUi7sR9B
r14HLbDsIK5pNxQq5NnMdPQOhdvTjoQOpNY6UIGFgOJEulR8NlE2TGMqXTjjpDx5
haMIXTU+D3GCBJhhrhxxBIrb1HbqX86WDYsmnc1pg2qK7mg6Dn6wpUJRg68PcGVo
YY7/9+WwUCLQPxodWmpvLMWC2gdFof2QYYklOen1p0QbRfqPMnXD2DqrMYUiR0Q8
V5sOYf8l1hM7CgdpNY+B2pv6fUuzvqvfR97m80+AxtCBCwd4gt+9jzhV8wqTtW6u
Xf186+mz6ZePVdEtIit4hJCE1UI8FIF//aCVymVs9sMDgvjYxLDGTy5o/8PzEIeg
bmwtISIDsObQ6UW1DH3lMdr209kaB0J4y6uAEU8h1HeZNIzcVFSwJfTa4rbTfmaI
6pJrhD/91kxeYcBwMDIZQycbJpjU8gm+8MFeqZmxejxOfc7QxYUj+L9bZ5W8j4vU
nFaxdiIyjngFyydlI+GN27UZTMnNkGrwdk9Gydw4xAaCvV91b/MzEr/68lrNyjVn
/R7Ue7WMQVYIlmytmMjrUWE+0dAuue9n3+GzgqwR/z+CpkY9eHjHNEDcdCnR8CUg
yuz70TCJklftcbBPMrw4zP8pDnvLiqcibbgo1kXsqrCMID2BFb9orUFLrb3BWDvA
dJGn9jYlmfBF/08CPsqHcVFuOpUkmPYI25hZz+zrJ9JixT8ivmb7OcbR7gS6mmwA
eLsco6c9uHbkaeEfCZbZKI6GFsLY4S98B76360OZhRCmXlYxHuPKDNRY4KuXS4LV
Fsl2mEI4gaSaTx+1DBberdGc6NMFMrniy4MO6u5L12jx6PsNFDvEvH/rZ5PX6N5h
IUW3jnU/ADMBsb7m0NgfnAam9uWjGgCcD7swXJN4WdfDP1UX/DfquN2hdCNE9JJZ
czRCPvhCfWeMqmlivKkQHc4fAK5B4ysgwmL2bQJ9Z+yM49J6osczSEWvAcTxgcjP
5NGOTL9LQqKMZsHQSeOOGvEFxZfW6GMwVN0wVUGYZFmqXNUq7Hk3BqbFc9/tDsF8
abtII7BQNjKT2W7rExvoU0V8PCy8CgruGfXyhSWEukpuMnnvpywGSXAvDuOEgviF
8L0w5QgaSXJkfMuFN1ouN21gdH42gzoUYrEtx/UEqW9/vvneX+6xWzhZ/FtH60NA
zje30nMPPA0p7mUXqNkZjauVI9VykP/NNrAiOAluKJL27HoqMCXf6U2Nglgrgkq8
oqEEJf0diAbVxkVcIy4VOSKCz2RMEKpSvtgpLjFrIQ9QSHXj08mz1UaoaXu0orf5
X3rjUGT2FRfdLLVydozJz+/bcPkCabiF6ytLDO1X0ngqSyprjfTyxcUc7lS5lRmo
j+ivBb6/j7n/ymRCkASu1aX4fkY7kQoeHdUDDKZqfWLvwgK8PQSItkZaPXxx+wA/
KhcU8s7yKL6bWf1rY8LXhoIFOyPQREm0Mwdwf7z2Fa5bmiNTPRbxLoOqY5Uvw3iH
PWdEPqapMqG2RAYwqlVg3cNT1MWE4BqiLghTQNq38i4VDEibU+BsjcnYq97GWFQT
qtMJOghvmX5odZr+tR9oghJMlSiASHTl3d7avHttwZtIYBHzEtW6lOHwMgQxysQT
GdvU0UHD8aGQkM6exTeyaX2fKhnahltPu+PqQ/Z2rFbgS5RwwcPONhVEYid657xO
sCepy9De5OBXMiG9QAh4Al3lExpz9wffj/yWfq/EC8qYosoYZPKQYOYuBZ+P3wee
KQNRwyxx1bVndWM5wz1hxDJZnuquJnH4tYtNXaho6WojhGrVjehovDc2XyAKJ0oh
DpH4jRXAXpp3is5kQ8IeL32lkaDJPR2xV6JqWc/dEEqwsUPEsxmi3kk/6KQGm5AH
bRaLqP9uzBS/CxnG5nsKwh14nPfCRjugrVxrYnITSMbdPXqW6qmJcCakmWVHVt0o
4RQI8/ht6BmkiP4IWPmJX7TcWEAt3tgnCG5Ll7LYKsD46WyLnwPKgN049xpvDUtk
YQ0nU2wf0x+Oen/ov3/xKEt9vsqMgs6Yllvqpf5+cEdsPw1EIMESVJxw7vibiJyD
xpQQRO6GzLmOky41ht4fvmgU4szPYlkHsiIkFRrOIm11Zb05TWgETOBXIdscmo5y
NP05A6usDplKCSPO+VP5dbUD6WEPoi+PV/SfQ+3aOEj4fxA92ogyvQfOKQ9+3irm
V3D8apj1AtffxhUr17TNvVBLbU28vj6j4RJ8rpcCr6+cGlwvn6aX9bx90urMgdPS
9LKJPxg5eS7o5fZP66lt10E8JQVzXbWrcwdLcTshn6YO3nHELbChUIzfz0slNlML
mkupE8muQk5JleErzvRrTM7gydU8yrRC51tepF2QBnmU7JzjuNC0IINgIWSrpOxD
fwdw/N1m79nb+hI90y577cOJ1dPMv/aYYjLJdJApjcyOAjtTmhWIMfXr/7qUj7H4
uc7gr5qO7sACU6vxSR1SM6oMtH2EQw374moLt4XKmywZUYohMc7lny/4ql2iHvwM
wN5Gb0jSGcG4pTsUMmDTxdcPDfIjtrwkKNL4fvluBEnP1KFT13yJA0InMfKOZd8j
N1NYQgdFfBf6mBfrMcsL3suHYbZNIUMQp86kbq0kuGdeXEOaffi38ct6zqI3TL2S
+WyF7QCqEN7tfqBKlt/YuXfQzprsoTxfZOVbrV4YMNqofuFbqjdu4S3sEB8t8O90
3gG7baExN8+4qXFuMARa/lAo6wpFplnIZKja+xaHxhC8musGEcVyzFjfcEjries3
PPz0QmsBtIws7V5OhuU+9WwH3Xc4h4xQJ4Lt5+ugA2V7m7yqnY9wb4YfxkYfMDLS
bLxCLABg4d8Hr0rHAuj5h6IZj1WFZM15QRI5pst/gTlcmJpxWctqI8R4VHYKmUfv
XyAYRSkJ53x0nsGx8qyySXX3p4kyG4Z4aO/jux+SVW8SeP3Ub6QDI7XG8FaOzJFo
AtDMVZDsQG7EZfktCILX4wF4d7yQEDu0z6Fp7WjIZBkPMKscYnp0ham19ME2+lvc
45jovWvpeyfBYdkJ/DOHGP9wvI6mvF4Gy2p+bQLboDUxPvn2k9Di0el/DLiY++IW
7wYmFpp8//q+Ul1FoDHlyHj7xxNQHyLk6jZRQ4UssUmV+aLIB+G18Vc/j+qWLPb4
qDLirbejYzabNiwBi7Buu8zlyAd5iESDHp8u++bH6sIn0BsBNTlOgZymhI4l+dfd
R8NNHA3VIjeaOy5IzsnjXjRJjenxegmxjYV39PfzwTYzx0o/nGztBcyyoTaXddbh
dWosdqSn3TbZU6SNZkKGcwKAqmJibT0sPAwoIRIOnPL3pEs0688GqukrIPJjXMho
FN2DkNYSNAcWpc1ZJKgtgypICGMBlNvCXsTe6Q3t00t9HBzw9dnitJfiVtIREo6c
+GgIF6mdbPBH8QTWtSNcooUPdxRKN2rUP54vuadnU9c84N+EqgCY9g2WRPvjay4M
gNX4+miMroWhw3YzXPB3InfZofCTQ9d7ttcNUQji0XAY46H4PIxMp96o/SfO1fCY
1aMrhzwg+6HGNQt6/1qMdZ0vKJf26Zp8Bh5/IPjmLGjSi+4MLOKEyDlch920v5oH
5QEz0befWLU7oJpO+4D0+rIKDJ9flco2kltxwfs2CfSbRr6x+P38LhkE7LZ782Oy
OugDyzEEZSqgT6TAF+BWMqsBEaQ0uJ9+TTX7GwxpjOnkezTnizGrdQk6MkFuVtp6
AOc0veKKLk2EP3xvzGNCXlB+SMpcuU7nv5arl6aIljqe4YPuXslku0nsFw2yr9+P
ZsEgDXL6YEmKpt8VgtuUpYX9LjaCZhuRU/MK0/aDkByvK3ia7glTEzS8CUZ2h+qr
9qybQAAfD/p+src1bQNpibZ3KIzuj8uNL8+D8xOwdW+l5mjXqLUdyT+iiTGEswov
m/CCNiCztNYIF5FpAdjRHhpee+g3KJxpG21ppS733xwJKmqlI1x3+gpggSxDLZlg
U6TGkYqHqoOGJYMJtGtJYPvOAf+KUaMWGPC6YEtZwkj2JkSnD2rwrJKMuKX4SiDL
SVNAgBB8i2AYhwC3/4a/2OEYFZyyLQwbPQqwvu3k70ZZz70Rsk0+6WzIPbSz+dXZ
4zGp5gDh4l5/DuZBgy0dp4Zho5THDkwLzpeViW1mM8oXdmpyrmZpwh5iRjkN/tBM
6xrE5L71i2rkaBcNDiuzCjKCoaA3wlsWmm6wIYubwJmz7sXAULSg3pnIgXpD9Hoy
BW4YFHT2Up0IaNcqeaBYZRLiQZGlWrI89XPPadp2LDRsC7D2JnFEiBHIsgqN31oo
xBrgPLPhAx/pTvQGBt2V9oypaxVgx7ri1nB8liuJwyRbIHpCpnaFfFAa0SoGz6rC
5tiThy9hLwu0Ou8YduoOERqfMIvBNnLJRLYEkNdTgFYazgqI4jrMhGMKq5gEksxq
mA54hw2HA8quWBS7jnBY7ukwtcGI+Ah+y6apjqifjUcHNv9gncG7jo9K/goDlPJh
J1vAFQ1rQ0Yv5TDYxGMUzhCUowz4v+CW2ln6/exlCemIsjhvXqnvNsHvsw3tIcx0
CnwrAclGdU4QL8597SmxRdJ75Lbhqeen6InH+MaCkl+4vYt261ae4WBei+98uu9S
pzhaB8TNJi1E1oJP6oPREMmOVfH5kLfIcAiw00i39y4pbQGwYGmvSwSyj8Af3KeK
yQihkat8iFwwyOlFP8F9K1EWYK10sHnLHvg/aLXU+qEfZBRn9TnkippMtG45lUAe
ev9MvIk5vfJLsx4UPAxfNSEF5ysjR1Xtl7PvgGF9fFSiA8DSLNBLkaDH7E51wKkP
06fu5FI9EvERBQWZJXWrArcL0Zb/+wvt8ipEvN8kiDc8onyHHRXOw5vprL3GoDf3
HZ/EO1/JiMtlDHeGfVCNbscsD/yzgEHw5wYVV8Bst9n+Ik4qh56HYPYtMa6q8kzz
07rMNtgWh/+Vv8cL4vCUZIPttBJcwEQ8lQqSCmSG/YfBeQW4TGAkQZd+q8TuZQsr
jtMJ5CBjJXuWYtBvbRgbYC2bevt2OQGV1e2Y+oBtNKhipFmjtq4+6w8FeATKvnTd
Kr2iHsx9D/sbS3ngMJVuj67RtcGrrTBWhr1bZVUCHr/eP7C70hVINpLgKgXaBIzF
6adub3vix6ngoPtxV0w8+DlYyn9lkicWOzvrdoA49o4ttRV5F0fxihWoXCLwF6st
84vaV602Hm2gRrDVhmWVcHrOWUFQJTESRhQHQVgIUP1NeD+LDislRqzMRLQdY/NO
MZHQ5cNPz3tJKwmIDkmGmBIGjoO7GuuV5avQy770yd12xFpKjX0IyY6bMcy924y0
GrPqvquE7A9zQfiBhwgYhB/KrksX5BF4buXy2RbPyygfFRqrVgxGiu87l+9S+bql
ozA4fyOR5lOaARB09Ay6GU+gaoUJjh6tlO8mAwLH7VmE5+KklkiZKGAGkQ63wH22
LZtaBOw4N3ZmendNvmwau6ugIeIGFOPURxlyQYl5XgQThSwAG+WhvES4dsuCqsuT
pomZv50PY5MBYHDAKx7ZJnJ+wn3BNHpoerNRZeUAzg73c7mkFwUv840eaiB2w7xQ
ANAhxEk3Z7y3iFf/JxS9BsQ2NWorQl72khO+kLajEUJOv3wB8CoWVzXzQLDXdqG1
4xOWteTaj568jP7Wj4YBWzvjl77P8BgcBfPOXeuoQmFzv6UKZJku7tbP0HhxJfEN
n0OkJjAqLpkZm1AjIyEQlP2Yz2UB5ngoJbryRdjpOh/aMbAb+DBB01sdkSJLCL15
utuwkaBJMvGJS+yN2CVtIKe37CHTCLuteZuGWhEZGOC/se0lMex3CqRAzs6kWFF4
kmtmHAXS/X0lOO8CC9COPrP01qAP5Z48qWTpxCplgWyiqjOuuBElknfixwm8yhep
88feN0A35UB1ekfYE2QTrKQfcboEixE5jP81xbeE1+XnrWzZJFF12Liyo1aXa2nY
LOxJrQKbTwTSj1brF8DdkTgD+K3v94SZvHrQ9Pul1+EWmiLEtMPbFeKGoOyqDksO
bq0A1pgplUgoQrQseOQkJ95B4wbOJNi6L3gsVdHvBONvrpeSAEp0bXksjITQqYq9
uA+PJt04uBHhf0cAbZHnDIXzRSbEm81qouOi8s/GkFUFjGB+fjs8euDqfdq+ajsu
ZxvBbeI2xlGrj9YEOgHFRJ4Z7uMGZJGGi2fjE93kYFTBttEaH69G5A52eHFextaz
CYqe1Wzw0gzQvuvkHELX3CMBCo3tw73l9rT+YLwIbpZdUs79MN6kOBMobQPf/rra
DMduxZLiLQp3V9AypRjXlL9l5SydMsmu/RtspXeEEPRMG0wI4+gUQJczDD5QKlmS
HLfJH4Zpd0xAiPJD26z55qshfUS0F3frAg8aCv50HpbJ3SHZMaB6dHG9phy5psGQ
khndtYlwVLBXyYWeatY5JvecuYV740j6S7vC8eGQ4gU5LsQlRYax+/3mcLHkTFdg
ebOzyULdmWoNWXY09TGk0XwsPeCe9WZVq+ICm9b+hyymYHNksJt+vTCBibVaE+x+
BBFnznR5mgl03gdryifoeS3eLn8P/UANbQgVS88mHZvURa3ymTNdum20xDTAlEXp
WGGNlnzeCxwEiZaoVBrAMTUFaElGQtjdnNo7UO1j9IFrQrIKK9bPs5i865uHR9Fn
I/8elLc6GoZKmWz0MlCHb11gdIrBWhPR4EyvLD5Xkn/qwbEHWvPzmujwmL7FJZQV
0w1vn47+2MoueuWEbmvRYUVVbRN44KzyXw7TBqGNO/vHigBE9nerFgrQsVV53Vy8
JcDdnV7Ex78LKHzhEKe8FxCiZRsp4PWEaGlCpki8K/GQ1JZcfA/rf1CpgKw0KZgd
pQVczxfvld+kpLaCndM7kwVVatxjqgOCF+8pmpo140Pb29cdx4D9iWshk6P0bF5R
nmv5yQu5sULDijf7nIiSHSPDj1NAfjlBQ68akjIzC5+dOJehzOemmIjAuCOYiM0m
8dysNcBf9X29xcgR2wTotYYDwd2S10aiQCTvN86Uc01TddEZIfqJPRw2tErBh9XA
MydmcYEoYo2F1y0ojdW3T36ImpEXkqVzFUHVRKGjr/SJVMLLFjQ01/BTm/jNxFid
T+uIb8LHBkFRbbTDY+zZKEDxuQwYS+z4VKdN4ad11vYVkvSW6OE7/C5mJTbNLdtl
hNp6w2Bb8kedSU9fpfp+ij8KXI0DxxrCaMaVsqgu8//xnMAgSHttbsbN2X4mpEj5
wApeBPjqccUx1wzH8hMMU8YHzGO5ep2WODrkjpQfIKZcB/ewvHhAnE42b/spEYB6
KLhfTeIdIigTQfYrnI3yfezdWDJ6azACZRU4uDGteOcothUAY1E1sJOG8xiLyVy+
XSyrdsb4jA7360n3y2UPjgWSPqrLQsz11P+vZ24k10O541yFtZpC+fOydnRocJpn
RSssdDT0dOWXOobuKFcZG43IjpdXxulJfzHXe6M+jCUVDtehTR3PHrGmzR2TjGD/
HFi267wXOAXgQsWv3bBwxrPWvnScHVQXcX9DgPvM8ZfTg5cSQxkFQt+rhQdZLXJl
ufKgIwL6qwZlQaq8xVtf8yvwbTFm0KBFb+Qsp70tisO0R4wWg/nOIUkrOLNcqtD7
royIzJHn8KbD9/dSUmuzmeeyKnJT5rUQyiI2osxkXDO+Z90zFT3TEZ4964bOI7bI
jFqDMs27mmJfTLSwEFrXXOC1yENJi3VTdlK8Zlh7eYoaFUUMbvV9+Xax3vNF3sPj
tMymC55kHHXDF4LVrJoKUaHqY2Pjy2aiz3iBQJ84TptopLk+9q7nRkrhLQ7UM6z1
bcCF5JbonL7lpAyjVvgzHgHy2kF+qeJ/9N7ih08lSiPiablEWShLxml8U/uFnFsJ
bPUWljrLXuIXCbreryaNOpMzBtbjA8bHIRx7fz2wBblPzH4HA+PwzMd8LykRwxMZ
iUMsSynhX/2A84i7HyF8Fcey4qUCpSa5T0bVzd3BelQdEp1jUKvv92Rxn0IVs5wp
xi4K3rOjq97dc2+jc5Xrg5OsUI9siCS0a5OPdfG8uWZd9c5Xv/ZKlZpZgTRAgITd
Hme/i4Av8HPDDKmrMlBmypPKdyPGNn7CF+lDe2mfjmqXT6PMwCbstlALniSb1Jhl
6tqwpo2rCpl7HlDRa8Is82eWhXd6ZjPCX6PNr8R+HaZv4QDmeSrxkjHZv63CWDB0
zME1oAMrcLIkQCZK6KlHmlIfqpPgQiT4dzfqyMajQklbb9bsJIRzFbD68+y2rOCg
8agvGe7m+Wsgw0k4aGXK3inDlqqlzcu9MAIQlu2bXasVhtYZEwbpvibvM5tni84I
r6Cbf2aTO5ZZB8xy1gk1xvTm7lBjiliHiePYu9fCdrSSblYtq0bXcmdhy/hTHZ0b
9lFvNlA1klAymDOTNDGav6/Nz1eU0MY96zf7527T/greMuQHKSvc4eXOyNXgiC7W
+48t73C+tbG01ANtWgpcHy33FflgWCW5Cyl7mbok50J8WJQ7aIXa+9ZQdqqCtJpd
WyJXncvLjBC0+4aS16olnkC9ONt98q8p+3Wc9MQfrwd/JT8/HE4pozo9hd6126mO
IU/m4Qld9S6B+JOJu9tyhUalLnAPzhYth7T1mfYThxFAfg4FMGqW6ig57xrfJ8uT
B2dNBjssYFCgO5aJ77EXUFNSQIeHnTHnq4nVaMfYpCY/NmKazun+4FddXZmdIRVR
e3Bi2rIme5yUag2KDUeOTb5zWHMOa1+5Nf+JHIhzJzfd0gM6Y80HytaeI7jeYZ0b
lObNicHqussW8aPMS3adfS/Jsnp1A7rifhMZhK14dFKVxhbaTYombBbjIsjfl87o
z33sn9rP6+3FzOd0+x1ClyLagllT3OmQCdV9FoQcTTqAYBb5ZwJRHW6r82UjIAoN
3zeQLkT+g04sluChRVQoEEewB435LUjkXu7i0Cybw0Y6dUNccw5S9svRsMSDgsXh
c/7vVVmnsFwEA0a4DrwjY2fsuhn9AmADM0uZIAMhxolW+kMkVm7yZpA4g8jIjZJG
cj9VU+xuCC+zEJimMbUC26PWbQJxM0IlLU9Fue0c97ttsFJyonoh46LPMw9P+QJN
wOAa4YOnSNEpZJzcZIJRN+wLzr+f9EatlhUbUO1XkaP3gF5zuSmZmoLStUpp5oaU
B04tdGq6uN08obzgMikqb7Oc/99XqGuttpYQsVVDXoUGWheVp05A9sXAyCIh9Mw4
ruDULuv83dJii0Ztw0pDWqj7wT+BwcVb22BI7pkp1dvj7UZm83nhaxBMFLa/Vp0J
q5AeIJXHZ+koWVWwSV9vRRDXiLbC+wcdp7wgUsZU6czeWLBTUpiih2LCms6p1itf
83a5UKvc52GaP8RylukzXz1Oszrk/rjtuW532IFlAK66d2jlI1nfpcQR2dgcvcyH
vPTUClEFM0v5eHgjKOnURGI1dRbu56WV/pgsZlEzLPCsnPDxmY4p4vgaPw1OR1Ms
9r9Zw8oOCqDkpyAWmrffuraLZmHACGOQdeqQutCBeogunI7ZlJsJfM2PLoe0Z8MR
0KjSdJvKEbyrHJKQmwHaey8S+4tnLOO5wM3MgjaOt4zK4Jfn01GeImLgasuvgM6U
LqW90BNJPChKX3WpKzcDP6H0G9fQcUOEg3AyXtelOY3aHgN/bQ/0glf3lSAjp1q1
/lSWwWUTyiE6ODqyzz6qWJz8dR2QOFdv9Y6cPOY8VfCwctqaYR08aqYbWLRh1X7H
B9E3dHKo4Lz+1q5MQnyXBHqzVN4yWUFwwvQy5SD2CvHb967AwdYcLr0xBTXch6w+
Uhw0DlbmHmWn31xqIVF2WM8oyx6s5ipDYHrWs8I32blWaCVAfc8+FBymH8bjRZWG
SQ1yV+d18i0dOyGwMTgf67QZGMxLbvnu/sIpN6KrNnyvo8a2WvGR0O68WmMeobhJ
ognOf8enUo9d702ur8lC6RHHZbDLboJItBycpy558mfa9mk3uFSO0vsDdqf9vdGs
3zGtBoclckJEsorRNiQztPhhSSK/F6mg7Vmuy3yZP0J2XajQVgb1sScU2Rl8uB5j
ituAc03THdKCvBfHqtgmt429zB96euDr2t4/j65Zp8p+WHE/R1SX3YaotdiFI0MK
acigjOX/iBH1EfFbwe0Xhl6qxwR7DXmW6UB9pLnwL+jWNBA5aYUc4jAveaNc2jkV
Y27ifhmFgEL465CXcGd/wJUxCp2z1z1WMTgI4Xj4Nj3j9GY6xd1xxR96kyMx2XDh
mjv4nMWHUVA7MUlvwDDb4JD3x15mIH9mvCr6mmm33msdoCBfzyiC0bnpOilxCZcy
7J/gH8DSzeCRAIsRCJvoso9K4a2OtxQExvPI1vVNL6PNm0yny4aOAteiLyLBXUeY
XRNk3Yx5xD/qZZsDyQimM9LN/XdhDssdpDl19dkvsitYmT5qyiuhkI+LRprQAR0W
mQN03raZ+TlVaaxT/EgFe56ONBdVu2kYqn9e5nZdQaTu3TIC+ygtXEun6LZOFXzx
l/SuoIN9eNDwqf7yDRYwPsEvi6KlDREtdUXBd21DilRKChoyzhg3mUfog4Y7RyaK
mwpvVW2cioVIWSoc97tz6zwraHB7lgmVsaeHyWE9v680h/90vAKSYclqlO/EMyYa
KHWGTzxe5Zw5o4jDwBODNr69jinG9T0krbTntvXxn2E88WR5DAHKA2WlETEFRvCa
MmZxTNxQxMJ57nWX1PoJCCddtUiXvXrQGy1NHokYjlNn5IGd+bTNAZi3kIsDaZII
vLakueRMF+w26ef1yCLfUFbsOEwsIWG/xiHNBXmEPzWWr5OkipbmE5bFiQ5SVm2u
L2lUo2MopbLqSfK4/8g/5A/EcxSrKSde0RMOJBk8dF4cP+HwS8wAnOhNVDqQO+wx
XgKjSPzb0OywdcCmaZBqFKxN8aeVm8hMqT7fn2FzgspOHmYzcYzE8PolHaJZgx2S
69LkI3cUfTxn657+BEQx1iO2xu21hLPIafA/QjWqCh5q9z7F668m7Pp4zliKmSba
cud91SnbRnCwMFykVAhr6W72dfUeXZxdu3TNXzerT59580Qd5rdO2fanp/pQ1mXw
FZFsZ5P9e7Mqjv9jYv5Zjn7LQWiGCKMJ4pZ2mtkRju+6V38h+uw5+r0rnGUFHr15
Y/NXXjIUaemsmhZEVIdCwTd1oQqGwD3YP5Z+0oqKxCYYzVqtbLZLyxrO2ahK5993
/wtQjXud5Nn+CcDlHkI+d0rgc/L6Eu6wSWMbi+LhQNSitdlRZ33cVjPA1OEo/Nk1
FeeCc4kX+m8eZKNqO8reZx2n5EVkmpWYZ92YivkTA/QXMhPt7ONXFqTs3HmI7njw
1Dpatv8VvUHzaaKtFogVnNe4jBDVZqeNMNTaciCNzdQmzUPe0CSguVZnGaLrEGrM
tttMerg5OaSB7DkYX1BlRHZkF/PS95d8jUnlmloHsQ9B7/eLZgrdW0qwDXRJC6jE
aH8n66qs2IwFMRzbSHxrR+hngp5JuGsfAR2PAdVImVY3uNGd3+3y6V2O4j/w/Q8p
rFvzqIP0vldOUbl1MNdEuYSC7g4Str01oMEXlFdvTBzu9CaNNae+rr6Wwg+izeJ7
ACrSWSHflSZfmtJ2peB0cMs0rCQXU4h3nHqGj5aUDkF7bjlfvxhrPzDjTh0OLdns
czGiHe0YSahB7LbE34NKwxYG6beF5DLM4agcBQAs7e6OY9SuNYBDv8xmkAGMZI24
Mt15G4QOfG3cZYK60ZieYRa19SqH9sss/yPMAyg690GlFvjB4zi85ilW7fCDGWUR
IWsi7wIUs25zBQk6sp+j+fsU4ObwpThAC0jKOxHsqV+xg2aZ4E3DwuSdYWjPrQ0r
OuiOICg4fYCMu2NqeYoyoxhlqAuXLb5Ral8462sno6fIT6JFmjd901087NZWWL4m
CyDof5HfAg1mLSpc6VICEGyYa5gOrg1vkWnWrDNmyb9uqx21rktNz3SqHM5O7Ps9
nV3rRp5M51gvTMqB2hJMik1IrV2wUOiSqL2GWrKEVXRaK2OZxpHfQF1i/4jmtgut
5znSPdXn6eaQkpfhnFQgBXe6zrT7KY2HGRxIwcVqFfzHuVpXL+s1WL98RE5XcGcy
nbY6rP834J/04JGYOo+3Jt34l/8u50eTGDkrDWSBFezPN0nAPeHTyGU8ywy5R/lM
eaNsvEuQKQTcArcM/ucnClKOxeWCDKEC0VtZFZ5nrsO5v2wKPiPoPUolP0DEj8eo
Nm33f/3me7HQSZUYl0MP2jTjBCdEIUOGQ7E6be4fSDqGcX9WCFkC/JyAdgnsihWu
IA2xingwHOWUe0KRn/2Z7KpUd40KxVxAoKedJ/gcMG4KjT2uQL/WyTZ/tDzGbf8J
xcEjmmVlux6RIocg2lxSYkIiO75aMpdoqA79yjMso1z0jDOAHM/58UiUupVYm1y9
oEPp4zyBDx9tztUAyucowIEpzDy3ugSjT1h+h7rLA/ZHn/0dbyFaWJ4CQqYjU4YH
PUl3RUIWv2tJCz6PazN4dGiLTFOfshW99UaoYIrCzTewe46KKWzHYtgDHmY3FTZX
jGGIM4v3TG+UpIln4TH0SQt2gP3FBfzimZcrOd8mjciJ4G1Xk7xq1ePOiOamEodl
HaCfWfqDDRApUpITkuoUPvFQzsjaRlkV+lYe4OUdePG0ehR0mPaIRaqsYVpv4f4L
0Wo+fyJgqcNMK0NT+6AKyUgNUbvqGzBqSGqRpYRVzOmJV2qDKFGzNkJAuuhR6E73
DkjT2uRQ6z/ozIuTpXfq8pUh+SOflUOSbQjHHsuNIdrhH2K9lfjBB1Kkhs96oZJi
md48qfcICi4R8gGSdwmy9mniazWe3BUgh8jPzhtL0mVlyvxxdv5Oru3z7Z98yMsT
nWuZWCuvJ9Bx7gInaCywXdcpL6mXbAuE810AVEuvcMRTrIj9LxGHYPlKSrdp7cev
nvsS+dzveSUWt09GxRNEIb8Nvb8KxB0wYoUacB3WXv4LYqExT5mh6sNmTaSxpn6t
T2pPRppJ3QrHWyMlPjStRm0uTTAAlgDmr0NWaZPqYYaYbvp7MvB5QmhETYGivlsx
wq7mJU17BtAYl5BbiDOqB3mHtjarPpO+tOqWCO3IzrOeKZ4Br3dXoOfeX9qYKB74
h8iu5iG+Zwj8TItrh4dtQMsCCaq247RMCL/MPfNEYuCCaDui5LEAMwOFM0d85YFf
ilrYhygVcT6GwlPo+Z2d5YB52Yp53AMCgLtDG4XRWqq/+wgmRBwaExyLB8yJTpTb
BrNCTjR4Mh5/1hjc7dHi6L+SyEWX/VlQ7kkLH6ZeP5i10KNNu+2f6lt31PQHrN74
hvz9ZPIEimxPyw+cWIFHx2jR/YLO1FH/sZyRrYf34LUlQg4ImAr0TNUWD3O2OdW6
X1tNWz/1Oz3L76aI0KoE6QAVW5YU8SSPoirxuKdWCpjkaLpAvpFt268QE1/u8Z3i
XAk/duYuhSGd6U3c5iOrUF2XNmb2AqLUUrTIWPsWqFgvyU1mek8OmDgXx3blFcnS
ytZIiozE3ZyiYfCbH/TPRE1uyZZh79QdZ+Mnc35WYCfgUnGFh7VXuaDV+BodTXzs
emoM7iRr8714p08Ky8LT3V9r5iDl177UXj0TwmesuMkRC884lgVRaPNuOyvB9ggx
3X3ehBVcIigUIzcvtSRXXXWm/1fHIDyRraAYwaElqpzu72+3DnZP9a4ZQcP8RZqc
WvK3JkCi1RJoPfpSFDjqOjsWMW01RVGP5MOtIXukBdCz43l8gNdgKdEe+ldg9/zU
8Wf+7XxEyEMHst2KJttlZvsjLl3JOvrK0/+GHCil1YKs3XOHN1fY/Yv4oDu30zX6
6gxA1tTtLSEaR6ssgOQETyl5o4Dk99vCMuTq/xWZY5lzIJU5TnA+l/Suc8SK2U8h
B9JmAbYxIjwZ21MgUr43J2zy/gmC8+xebn3yr7Sq8smkmU9ywmMshKMC7VJvIjsc
+lkEQNByBHYvCggOjN0X22Ez/+bCB2wIBoTtFkEAI8ZOt2tXrWyZT3LaB8aSeLok
k2qQsJ8ShiAwijTpAs9VtWzxfp/yIacqb8y7zYaQvt7Zxu4mw1QthMwgeV1MK6lq
OYrSZNCuZhf+sExStECOKFuKXk6c1NA99+XLlyGXjByYcqonv/J0D/EfaIKq7KKC
hni/UF0r3kZH39FcR0hDtANDJslM8GYFKyQINs5FxhDjg357NJAjVa28nEvOYdmd
YhG4pgd6HWzWsIA/f1aBAcrktoF8k2euz/vf5569hQzvUSUhXnJX5iVpDGHH43vc
YGIZuusEq3Ra0fMRrMcbqSX42x7CV1U0y+hk5fSFsjMpVhx5LfQhIuF/TXv/dS2+
VkoO4YcO2impExuuF6JtiYG11iKcohBi+JRn0LpDian9UsNg+weU/nBwhZut9rJ/
Tg0wG7bl27dKL9ha8A45P1YUpH4jUrVcF5AkbDG8tuLK0o4xGNQh+OiohwND01ph
3n4fOuBBR1QcguFYeZEYUBRvicR5zH2EwtGgNRV8fmtzMjJ2l8zeyjUq1yo/2j9w
Lgdj2ZhZ6iqpzSIyVBgPuASIXaxXNNU0nUM8hmUWQMEor05QdFdvonXLLIJjrp3a
oQDX5ip2oipvsMnWGvwYeY4IJlLfkEeNFex7HjGZnH2StWEh80fL/aSARsd+a22F
fjTqS7tvA9sEcttfOZqgxG66vhUPu+b46xDopczOYjzeJ00sTds8Xj8ZINEiLS7M
effpAYZme6D2iUw3qJQujktdQIW09Ma0feoiyleVJcqY6N7GuQPtBnh2SjZsNjWy
2tspdwuzIDn1Lat2GWlY98p4F9ylr/Qit1UkjW84sdvoM7JR6B7N4U0xio8jQ1wE
j7w8xKGXpl319XW/lf5fn+w7hQwfdD/rl8qjoXEWQeFLSJ7oLO3yMAhh9p2wBnhT
7cS8lTJrXuIdIQOspLkEF4hpYz4Y8OEjYJqmd1FxoD75FD6jdoiwseaT9tJ1d2nf
pS2fVmegfddmj5p2FYpSDrigrYWOIqw/qjBxOVAKFe1Kj+m7il+5tdDqz+OYxMhZ
jkXMEEkTVVtRvUtBKB8UE9cimmXe6QXGUNMHEU7YmpEMx0iBXjc7S7bXbwcYwH3O
m2sEPLQLtgoSzubYMyM+gZQtNH2gboTUtIZIjG9kfj47ynujJxR0/M59D7po/sdG
cXQQJJv57A+xTF1q9B9x8Z3kHAG5LvKbHPx75KUq/Nycz+oTmjvRlWWkZan/MSGr
S4hMnC83AobQSbe1ih2AcX03xK94J7tU0IofHxJGPfWN/7xdmWBebkxg7RYTQ+j1
n3yq0FuJ+zOXIRpJAAjPMbx3tnYHOlIxpLpf515/+mrZ3mQQY/VHig5gO6NG+IFR
FLjwUiGRyreiyLDH/ltEMBkd3dgWmnNaFn49OUDZPz1QfCESF9VtaifIa4xyPkOl
W7SpcwENLUeYJYbCGucr9lXfqRAsvXAdU1U8CiNV2ynEZUCrJAUjRLbau2xrhwZ+
53uvORLJZwlCAj9ZGKGCp0IDPNw6jlejDxM4BSdqQyUrPGCup6JSRE1GcbbX/tZp
Oy5CKzsZ1ypCforNY0bBZLN51vEPCySC+igW7oZ8b45Alr0NfpSurmx+gJ9chMnf
5UBj9OSZzgNttf5nfLaVggQmzXyoetW3En5e77M3NHJcvqXZDdXRqYMgPY3xk0Zu
gh2RDC2uVp1GBMFYVuvtkL1rq1cVXRPDXuZOwQHOTxcizWhK5dzZuBita3aThhMN
AzR6mtqRwkTOmMEeZvhqlE8rPplvNYyf5G13GRfOX+9XwSHWfpV5WTWiZBzSbE2Y
HfH+aKz3pdJfXnIw9GTJec/GCsY7dhnvORbZ8o4lQFuSGgUnrgm6ExfMHgaAZfgY
YNW5S9HMRDSlhpee7l90ssQmWWw7zX1T3NMIkpAeO5op1jA4fqKB7xQldnjUKVCO
yVJDtSTmFG483Xdj9C3BJ1IdZ6v9PhOCW6UdxnvtUgRvUXHcndRR15YzXi5AwnIz
dm5WKXJCXEaVgaVPtpd0cAcrRZPWNcYrf3/4PFHcMxuq5UBSsJtaJvro92XovUqk
ppNKRA4Ir/yLW/0vFUq4Vpea+XLGA74Q1sYMm7xYtZtlNrsP0NGrL/r3u9NRasFQ
vVUOMzxdId/43YVuQVNubJqIuz6va5OHRITowS8GVhiXZqexl49Ubjxy26eG8xnV
nZIrBvVvTJtxFDwvOOon+EHl1Do39MICqL0FAVF4yAwctNc+VoNjI1IsZzdHHDbU
0YnXlDN/VxABKjVYULhD6KUwdTxOtWByEBZVwtxpPejHh5UyPyF4pjekCLSecIxG
be329tWkrOCRkhvw+UEDd5E4HLD9H/WkOMh4p5fuDM5wAZuV2NN0cVxT/odt9Dtk
VbMiy1wk6Ky5ArtKBAc1xFvI/tE+R53nQkVIrbJkdZXhObcNPLgKkPx0yxvXr58D
GOk0I2u/wZO17qZ1vunczh3tP9NcDYXgw9hpUnEJqGiKZKk/hRN3lO7IH0NGmPpt
d8tqYaTLMu2s51PaaPBWkvNIKupNr4zS3Dw6vdgvk7oJZgZk/H40+LCRLWNVT1HI
d9VapjFfRGuRQElPtDKxFbBEe11Su/UPwh3wbiUrLIb9ILQsRdoYuiS9ogy+2K83
cUVVFNm8/8thExLwwKdngnrIPAQpFKKdQmaPGfPbUwKV8YiHDZfBHUvA9fBLV8jC
i6R6/au5Go+Bf5X+CMDdUAuMzYmIEXV5y29v0L0ek9K4sEAU6+0svQHjMqZA8SMP
lI4s7BkTPtohvQQpdEsYthDFt5R5L/xbq/djQO97IeirAW9NMz4dZVsY8zinp3dQ
LBYebPMSODfbDguyx0tKuy4ANEvZ8raefHFN4nDdPI58tjuvDhvWszQfCh9sjeOr
D4XjOG46ovERRlGRr2euo7cud04EVRHlB/siAAAqWLI3QVEtJJKtPu2h9vOi0pYX
Q8WaO0nz5+qPgx4qha7T0QBazzmdN91rv/RTnYNmAo81Y/hwlw9taTgDzxSgPln9
rK9TrYGrkY4s/XA9DjdGjUM1kg/uE6Z+GLe07NVwCbBEA/Uz0FkxAEdt3GBlV7dE
E1HWtlgwezmHvN5owI4kJxcm43u+hIEwy+fZm/zorwj1qGNGmnwjUuMTOfAEApel
cTgmodKuoH1oquTIH/BQm5/M6R55YrtoLUWYhKMU8HuLvRgVenUA7tvUMQi/+/Wd
LByNea6jcI7tqNkjhez52D0Xeth1OsEPMpPBJGWuoqoWOVoKHNait5/FXXIjegDj
oE+2O5ETu7npa0gNcQClKPr2JcK5204sgMKbRSgmUw7M3dNUy6+3dZBU1RIQkcQy
zwP1bZhb9Qzk9VxuHwWFHvwqsJpyXw83LCLbpKvcSnMH/JsVZzrqfre+lYNyHRHb
mAjs+1I/6hFVynS2gFtJnNyFb+YaJzTcBtloj43HHu3yulhdkYXuJoi+CwSU1WQN
KOvjruKPGNBe/NTQFoIVvDYR46nX4WZvvVOO2jR7aNnAE3eAB5nu6wQrPuWSgfUY
nvK9MfD9Coa97BM5wc334r5XFWJRI5Y0RRdscPZFI5RYNbMFBhMN5swzsSbe+44M
9MChiyRyWsb6nZDH4zSvOXB+08PrioEiUgETO9R2UsGNGnoDumFdC5enYF92IPZC
GcAzpOist5eVAJCy4MNcwJCddp/AnWdK9Uz6fz4nNM6abowMYNReJx1q1x+tJeTr
mmywT+vBijt2kl6eVHVLVoG9zMoH37VPdECCQnPZz/pZlQZ2e5ML6fONjE/Yyh52
VZSgRzCl2Hz7ffY+OuL8qRYeoz1epIOBoQE1Bzt8eChW0noXvKetxXZpdxn8XM10
IFNah8eBCZTH0UV5w1jei8Tb0drbA3C95ToC9hSynAZ4bo9P3a5iG2zcMJmBLeJ0
ARvnNYxOkhKzHAyDkYZqBbI7R5cBUcpD9eJBSYOQW5h6oZ4domWcuBpHUvE5AUH0
JpqGLqmSnUo2v8z9sX0xSWj89GsSsG8NKyrbRphA8Xh4WEKTUNRF+O8Xa9s3kBJj
TNLpTfTAPvVVoATyDJQKl4P8s7HSlOVAfu1KgZCQDrPt0+kp0GJlD8Hw/iOntwvX
0+RpkUM4/qrGKG0qSSbH65AEtcIBAr2AUpqwbj28ZAqtFIxAwO5wqTp3LANTGczm
953NYxj61BmOFD6ZMmLZgx+AZoP6EGrB58bQMxJsFhFcvVFiSNas0qGpu0BgxNhK
ildPJgFK7p0ZxVqVo6wNNh2vUIcjxCjBaCQf4jhCo1kmWlREOplLYk/z4JqIGTZP
xQ2G7L0VQZPsdS2tl+t6G5hNPy4Wp/CNqRQVqMpIQgLQMMhqvgiaAfwKRsWfWIW7
O8HAnJlRJA3k7pXmTCQFlqJb5fN9XqU7SSgUyAVc8IxQMtqFSIDl0rtPxn9tBlMs
3l0i/h9e/YpZSkXVVu66Givm6ANqRuDv/2/bgIF1Vf9PTVsG3/tnuw8aingWBMIw
ama7DQarY+feOdqFwVOB6ruTWMFaf1LVzg2pk7591+iNvVoddGpDpFl5E0Vj4/Jf
JOuxov89l6pdLDV46hjsPLI92QH9uF9I3JA9AnQDaRwPfGtYQHdJ/tkzg5fWALlA
6Zh8U3i8Y3XjgnHTNXe47edKT1rPXD6Cvkjpc6qsaL2mxaRoDAzBMql+T8hz4t7D
gpPmMno2SR9RBs/fqU8X55IsNUg8rKIw09sqkDBOSM7/VO+uoBwuMcLevQgDZM1t
HWJONt4mPyNns+kW7QNC4NVdSjxGrL5FORak/5gdSY5nUz/zRmCjC5OVRWVArgxr
++WPSnrM3TDBlAt29VYHpbSy3N9un1fpJVhx259dv2mJsTIZ9Rx42vCmlkMfYKrp
Cv0stEnJ+JGGAMe884YXSMeoOib9B2l1ceEdwU3HC39nhcv1f3QRAO4BofEaMAAN
M7mF4Y3XlL9EQ3OEhjH9Aw2ltTvKWFbED4t2TLBsrSBAju4Easb6CU8gcQCcNIIw
AT/RhDAtiFRPm4hto1z5vESDyxc0ZRfCBYNg5QtTY40nSvF/8fWM4+OAkNNmNROC
rv3dlPVW8x44JAcIluw2OyKKs8vDaGhemj6NZb6E7WXnJoAB77Js5LXbyvXCL4wr
4uCo52WMOewgY6nzdQ3TwjCotD86RgRdRWgWSG6sOrtN/upHrn0f+CMxZtf+UaN3
lq6C3J9s0gcjw2tF70L9HS2ZHJSCCAc9gR8BvNsyqEk5wkMO70FtqrnVeZ6bfmTc
Hke5DiQjDmSyj9p6aCT2IlXXW1vQJ/6Zf8RsB2+6IaCz2BR5bgtBqKsVwYaQQLiL
YPcaE6T9RRj96GlS0KHhs6bRpT8/fNlyMXjcruQR8sU3zLkZdTBSKVXBTgOiSTUF
fjUjdQ21NmsoIbISN1b1dBwJYs/IKRM0GFkEetMxbYp3z4UNDUX3bX0CA6UocQKU
dXIMmDQdvvVruoKkKqi8mi7Zv6HY52Gep7RUhwnV+qwB3IE8ggPcdaBMyPNVPp1+
3x4HXj/57EDpV0doxNtholz17D0ML+oUSqc+EpqQc+qdolhoW5HIYeKHAFyaR59y
M4fzt//UP1d4i+1KeoqELxqGSpg2f2f2ySPNxHbDoFqlcMCJQxle5mlEbGh3/LhY
WL2fqVWIJpZe18u4xZ7Ie57JlGhIpZvnBWtBocEh8JPwSeYkkzpxiiHDL3uqOrsJ
tqul6zbQhwGJaKllZudoJ1IzNcMvFM/RxoM7DnSecouvuICkvtE9xpdPTWMx03rX
o3nSjTU9VLYRakc+9IbZa52nyuBZKzNPj55yvU7XX3lVMKW0DVDpnZiWGb+Qt1ci
yqfF+aIPKcAuq0bS1mbo618W4EpTQb/CSe5s+BJXahQN/JuXpDB1W9ub11UOXAS/
bPx3IJLBVxV6fTRmFHKpA+ChhmlqUNqDm6l9FiK/wdwY0QBzFIHyfh9kW3JJwZeu
tCPDRwJJoU0cqUI3MQy3xwkOCAwTTvuG8R5eGUz7nU65haHJq9twDXBT9qNuLzmu
pcU+JdXYEPxHSOd4yOu8V9qdm7xLkUArgp7Bm5SOTYlqRmKHY5cUyPKBwNxm2eNS
ulmGsPB+9IFYuYu9MAQwRcPDsN+ejA7g+LlwS2G2z1bLXiSECfbvIMkBqPdJ6n6E
h2VWRb1E8ZKmUz5hKgucopoEvcdq7qW/iR2tcnzJtk8jlry06BoEh6YyzkF7NLGu
l2ME37YFEpMKwvzAUt5Q3OQWSByTMH1kYfcvlwQuu1hbzzCYm3NpVEbxKyOPvc08
xLD2FgSC0WJ7U8jPHZFbYQTTGIOt3+JSCR3O7ug6GybyXIippi8bvGnT8MY6w4HR
6mPyExkDhtfqIe/EiRQQWsWkrPk/vAakzapPnEoDEePVaqx3BxHIU9vHlFL/JlPg
C4URIgPkEjY7sx8KECl362MRBCj38oVQvBCBtKNbUhpca8Gr0fnhHwXGr82b0+1j
7EKDxdyanZE5DHQqsfss5xyh3CG70NTCi2bUKdDrNUtIqFnAV94viDnndq8125Mt
HMLRtYlX/+IEe3AxQhqao6d7i269QEtXmkF/UiC6Qvy/Qot7idtc9scKQhxJaAbB
YlWW3tUfw5dhcJrFwgcdzvM14mxes+kf13HmxT6TRTGYnpavic4K6VIYo0x+/v4U
9Cm3EWLQldSq+wtM9y8/uL/xzI8QXsnbtWkm2r1XjLRkrCIv4ID+k6SQG84HJNOz
g8NlPCPLIezEZjH1ek2IPxp+nlySJq+eQ/uRg5LC3tOlOjHmHs5Ac5fnvGvVkJOv
lcfhZfJb9DQLVZ7wYJGQqNQIo+TuCiBbPcTlZn12nF6RUsKYavFuoP4DFTp2M3uu
zHRBcSXEaGPByU6kZKGUSEMs4zBEgP7nuMiVVui3avt9y5s1CGOKY0rfkCIrTuSo
TNeHmRxrdTuepAcSo3nxqfSOFncCKrNElnQLHd1BcEvrah7BI3ndcOFOQFxcy5j4
jpbcbhGKO3kfTOU3v7WcsEH/nSJ2px3ae0strp4eEKYm6lLHP+Kz3pmaxPvrGNI/
5r4fd2IRq9Q/2fHL8N0RTiHfU18WSfbcBDXcBxe9Ahmr94XfzKs6i4V8AdMdnXRY
xLYG+5TceNFGKB5SENPkYtk0T6mZkocUkaRqfyCVaLnrGAVgIXK7mkujsX8gbNmi
ddxu/05QRCqIy4hNT4d6iWvkBcy2aQSrWSBvnG7csJCUQqr0CFn4SCBLpsKZ8V+c
L0ZqEH6Jn/o1qK3G6XQpK8Jr5cfJBH++1ezjmasEY9/fjCgSJG5/UYkCk81f/dbm
Wl9IKrPenty9auZYdFlFE4/9ngKSzvshC7WfkggPxBxD1SlW0NtWVIOUekDVVBzy
5mFY+9jewzKo0b6xYE6sC4TOOdaFo0wuTGOOfzYYYfUaqPdqewInldXj966WAyvB
d6nUgz7CJWl7M5Kb5Y0Wnc+l+qUPLHAwvIFGHAcnhCM5pSz5K0KRkecN1oQe20ri
/JeJgtZx84XgbrfooROWZmaHs9ZJgFOQEtvVhSi797xo6JAipC8Q7TmLXH69BdDi
T92XadxeEz26f6rh8VzBIUzoWuXu5KWwf34bRlfWverDlYFEF6Ox0KzOEcuEpBPh
EGuGkUmR6fgU81QE9VhAox1qXb3I43wM9L9/NyR8jp8i2i0xr2v7jzmqJ7TLZj+7
sgUZc2P1DyFmD9GGHM0nuRdMbDs/VcAYhP7wkCexOK1MnIrB9Urgre7LZooRvO3j
CCQtfzyMfZeicr2M5U7iO0ufvCH+hQ6vafvNyVSr6f0CwmU/vg7oTM9OUVZ6NFLN
xAxLq1yy8CFRrHjfVtojiIG+4h6todjTs0yNC3f15yhOUNmkTfNkdNEaGshzNOVW
y3pnSm3W1TxFJmeIwbxLeBxdU+UqloUHjg7kbKp5rxj7Uo9XJ0EUpP/mo3u3gjdx
SmvJLQu1/C8PBurC/Q883ZEqBoCDxijQxh7htXIgMyCvRmwzRBuwxFYEQib0ImMf
oEfczMrWTeo8oyyd+Ja+wFa2buCzZioQLzVjG6/3/FYaXMoNIbWQ4y+gmRqNxlIO
6mHyPFTaWxPjYnyGoxS2/hbUe5Vcy7KdveS/qArqHUFA2ZZ0HDFcp19Go92QKDYJ
ScEkvDxln861KllxiV7QPNDf63jRcGc3iy/DDRxk4YuYfEYDPjZrGPIqS0FG2epx
kI4jObE1FbfRxgLkn6AUbO7BL8WnVKogL0XhIRtgMtJ5fQE55JZqWt3irZpi1btb
y4CAVt46F9W0ytEsAaRShO0TBJJNlSNr28wFa1H/9OuyVnlJQvvQ8gygOUZ9fhRS
wY/+Og2YRCfHlu2K2XZhl6/phrrnI2Bt1BbZmU1pn4wxUFF9Rn+KJXBsOlYKYz7N
nf4r1ABCevgnOdtwYwDDGgWB5xdAEFi/0ZBBTKwzXmK2ViXQ80wvDUiXHnF40BDg
0V7rOwTmf0WWdg39bQcZGsySkTQKymGWjcellhtGkXkGXgZap4YFVm9x78eKkTKS
khj7qp/sDzkp7ABABRWjQHZHOyjPehtKBQzBImXl3QTou1dekKVXT9dWSz8X3Xh3
HXzcbjcWchcfejKIpwv0JETNIfdXjFniii+hvA/g5WNzxoGmovnKSa+NXGM+k1LE
3JWjNut6dwP3FUk1mCoReYe1IHyqB2MKYh0am80C1Q5XPwvRmNvHkbXnxh98Thv+
4JmWxvx/dWjy4uRs1l0lJOw6L4vOF9K/fjc2TlwmWinQWwbL0P6L6cxC1i/UfOhI
hxoxnTbz/YMpRWnhLwM/BAae4oFuRpIjCJkwPzPyyKrvAAxKyONp2GCVO5Lb5RLL
vrKzWD919J8p5s8GFloW1h/XpuGX3RkVtmx/r+OGkh11YmyEIOpX6L+OQ/q7QM7h
PvG0Oem1lN+LN4+rErRNdxibxZrPO09fa/9eWdUitODxsELg3An8GtzGC1VaUx8n
m1STaQYb9//p4eYP3lESH07Z3Gf7Qg5jKI44n/qAFTUaXEvClncaAI+jM3nEXVur
2tUX4683Z+Iiyl/GAPB85ZFxh/tH1fr7fdJf+ggeQ+GsZpFIdy8Y3dvGTUxE1TOy
asJZt5N4MycT/YYf+YGMGVivVGx8pNKZ9+l69uof5wFzuEhsEhcR+CanTjkHi1PL
Dnk4hXGhtnypn83eEt6vnUFlkR6Jf7vJeCYfFD7KAhbJp/PxxBFNhciC9k6GzeEs
Xi6q0rftc3dQDFA/dZsBDv5uIqSSTH0ybt0LffFkFjDUWzIPseshqBkx7btLP/qZ
t7eUP81KH9S6kUtKEcRo+qMwfhqdfo3G4DcTRqUcxhQ/yZKXNAv1qN1kGcNbof5Z
PggNtj7wdP3Ug8iCQgtTSdNunoqw4mXbCOITls97zibqvYL1EXg7C3ebS6t+tCri
lgrlM2uFFY0FkgDLr17aTzQPGBqlfG7QFFEAVNN8/FiYLGKQDaOqSmlsHyuJL47h
7Rws2oN/L0nb4fiWHOKiHCsnKYYtWz6ImFIPSk4DcPh9dBR/j+ubjc7YUlMjv9Xj
4wLGgcoFBBn+o1tfVT7TNUS7Glw6t1+e3QELvg2lgpWPJWRcgIlixxp1ShleKcPq
y0szXsESArO0TyFRO9Q824ZtwiWrG0s8e1uWYXPARnXqgt1hDfWIkDCjtftKfIB/
aYvthqs/8MnVohPfziZjA4TMU4PZMXw2ssFgVekWUN8PrOcyudnpy+vI/Qzsl2pT
PDGB6qMcEoZZA6OeC3170UDWVWpx06dUZYOgb8hpYMM7WELFOkxrZjsdY/FDjwNC
bFOHlpQ9IIbtKM96XyFUS9hcnzCroNlEHmV0t5s6J9LJzdnBlKfpLz4OpKrXNpz7
7ok6uFq5b0SE+NVaIRIUmFxUjq1ZVWsXB0xrIgK8GF6xYZal2akLhDJANfLVM0k2
tp/eAngH3cVEPB0BZVUei6eOvNEKDZinkFFax9zuqwBZ06XKtpgNZt3CUxMMbXEj
Ksk94AcJnyMyNVgz86dNsfl54u3ljqZrAPYWB+FsDuzfpMjJMDhgShtZChIVC/4w
MdzlKZ46XZ7SVXk//JZh6yODD17g2c2aPn/22u3Mj3CZA0GH7m1FUXzaFA+Mq8kn
wACJ2xSU0dQth21c47TGGcYabsnUe/S9+FAmpINxmp9y3uO5WecDRWZxQAqjH11a
0HftuoxX9If6R4rpxMF+nbsgLZ3cd/0JrWfomcCiLWiOTw84+jq+/aH736gWJ1gp
oht+IiQx5eY+4HPzxzkGa13h5J5679JPGdIN8P21yiENHYBJRJtdjLkn3WPgtVf3
JLZDJtR0Q25eQIJel2kzucipvPZ0jw5YUTpGIuGhdGGJvVpqbqXx7MjFiVwEFOis
5Ovx6/bvSdqxw1PnQpOswhTes+kDTehIQopgFyDOh+bdr1sgE9FLUOEl/XzzrLAa
OnjmrugULvNTOa8wF69Hdw7P/qdnXANeVsCHVFpSjIadJ3ta35avyJzigD+VFPtw
2wr0x59f4Oh2MinAOLC3OvjvqDgs5NIZYo2aaXhNoYKffYiESEFvXiJvKHrriJfj
MeWNxuJUTQyvB15exxj9sntQbB2AFzgUjcS+h91SGoB7X+fQGATeLbbeWgORGnp/
kVZi0crei8etNmnsQgViTzdkbrgdIFru98Vqg9Jlqyscr1sbRbHhY5+xSNmDkUk+
y4+DuY3TuNmmMm+PxXGvM7iqpGzpsE1jrY+sykz1CrRroxUS2UuWRMv9cuceW7EI
BrBJDDFEbIepMs5s0dKU/EmRwpRSolHtMlsqL/jBgj2nNlmOoFOZ+ftsxNnmwZ2W
D3VL00eeTJkNTGWVewWj8tChyUAtpgMW+TAmeyMqWkH71OCIDqTmgWsKhHzzSwmU
dOTmtC5orElDWFYM0fS8GOu0kFIl4WVrtCw4B/+8bbPJCgZRsRQD0mAxYX8shtwu
0YSXlrEdTTox1JyCpQ7cxy9OwuR8ei1LLf+GQFRt0V1Prg3RvbH83ftzvJbVRj3h
cpoKJLb+0cnNGz0LTtLpdVV3x3oxZLJOrM3xAzjXLDvRDIE+UDs13nmJ3tWQqGu+
oQO7NToR+LOoQMjPNw43zrABlW8TxNeNlWFJq1pvmVDqs6wmswqXZK+RkEIbPPGg
RyE9yRU2GpCaesWSHTqPsCbRIL/uNBBwu5pjDSGIsoEyou+HRUL0AeqCavdnTjR6
AHxBfJqL0QKfdQEumEp8Kt9NnbABZ0Lt6k0b5zBAOiOdArqHBK6/QU5aY5UlTdEK
4rK+8aQAjJ9KfbEaBPWX086hKDn5rICQXCRWaTdN26lbX0HhvJ8hZlSLQVZ9dVw3
yc1ZDsM55YZ3aeRXSF4Nj1LUsGSoAkbbi4IpDsuYcKvrdWkhTtynAi7fzPfR98Qo
ofwZk5ybKRnR8VJ5RyWvRdnmrrowKSsX/yS5Zsc2Cp4HowIXXa4Ax+3opaawLGcv
vyzy7zWreCYqy8aq9/q23lk7VgxkPNyXiGIKUmhX4VLps5lLrMioI9eA0To98/eN
eigc+1OJBVZlxmYsi/3TLPKAlyrqBvSjpkxpXdNAOTOjru491zqfcyU8sXzkd5kl
lyYmCPZ5wru8IgzY/T+0kZy3EIbeWhaRy+nOII8tlmB9NWCbLA+M5D4TI6R0vicJ
zeJBLQnMwxe+bRobwkPY1OD7f050+u9pAPjJ8jaP1I6Hj0FcNhhmcbzIDngxU66I
zKt28Wvwj30JQWRSs+68jh5B8avmJi6tISlxqxdSA1R3c9JHrkhdDatkat1k4PIh
16SqE5CI0FHxpc6JGYVsLShCtiFSz/l6l2xDDhykoEhfXT5hzWt4SVHbi+K51BVg
AwWrfRVZ2tpvmaZkvLoSh5CUMz3mw1SMIvZ8y6foSgaJ9320PxYXzHooS9bonINa
TwzOPMA3WIjTYGgJTV72wAYbJpkFdQ6cIOK87ijwdrV0FKLld0icO/WlBe9PIWBg
Spf/vrMevTEoO95GOpS4RdyMM3uEAp+zNcWhk0pHfQ2m/FVmJ5qMOqvtrhq4nHg0
7+plkCZeqRJ9oeVnhl+KGfwktaS7Ain/PJt6aGtW9KpvEMBSMIJGbzNFDu2SXclR
hdz2/FTt+9SrojKZCN+43lR8rCyPvnzOv4XNhoTDlCjhfEjI+JaHpoZ4jNOistYh
LMmYT0UIIYGq6mzgyR2Lgt/X8/w8j8akVyLsPlTjwgCHOi7pW153R1bbgeoYz4bF
aL2T0nYBY7opl4oOoWVWdTY4/38HIt6do7b/3fpXgPAMYnojih74ecZkyraqaAAj
IkDyqbJ00nn5Nkeep2sGNjC6ZOxGZWGOsFbknKVIcpw5gcDZsx0zFFRGxvorQRfZ
Dy7M6ZrvU8GbE/fxC9NIyh9kPYWFqYFyXQLdkb9gMJwWfCHvOn6S8e/+LeTYiHgV
7q+k9Hv4XKPR1AhbJMoIzcxSLorFCqGpe3pJTsqkWJYRpjQRXrmavTGPjJHkOyiO
CkfOHS3ggI0kcCLHd44kLSgF6KOJNhYeFmg4YxXABQUMX0pwgs8kRzv8ytXKXE+Z
sP8Kf2NBZARjigeIjcQRzdJSLit4q89zJh0tSyadGhZIq7/CJq9A7Iponj233/EY
nXSTpxYIYH+L0by0T35VV1yWvKzxF7hOjmA0zqQRMJRrdpESIyE27i3VMLrWIRXj
Uzf4917puJCuS4Slbsy8uDFwB3JwDX2w3vlx4OAxxzbTKrvseCRBpTbvHllPezxT
rJb5kTO4EpR88SNTqZ7V9O4qN/ryRRxaH5EOaOk6BUU2mtSy9cy+l5UglD8IzE9W
LKnGWSGhRF70YJdl/Xcvh9qsOo951IGcdFaRlW3vfzEYaQxZfEGyI4eFNb5p5ieh
wAhX4jdSl8/a0B8H/ua3eoFm4dTGeW7WWDc9F8Zes2X+DNhfDS3vzzlHCpKvjXEz
SclVoKKkxZJp92LFqc6bdfIE7/LZ7CEc7qksEhf0z6SfHJ6aKLUQffCWxhdoTN1H
fP/13PzUQGl86ycBwUsSIWtFBApcz0GKjM2Fmm31U4so/1cYui7vNgYdTVsFTbRu
4mFbgIxv4sl9CXa9x/g1fPweWkpVDsBaxRm4KXQJ26hjWGa+gl3zelID0sMbgrX3
++RsNOGybqIwKJ8G+k8+ZnnNUT0uL/2jOM7ok0efHKnjbheKg/gi/C2q/3uJJFxx
mI5yWlWks1zHR4y/R09fTV2eXYJG8A1gacNk8ruAb/xERwe+hpRIpEZTh9yty2Ew
1oXWRTfJKxoaksy2L5mUyaLQu3bGQwLdhyJgoN0IeBJnuEWNz9DJBEmCVaEjP2eu
v5IPJ/IZnrXNOnA34xbzdFb6dJ2QMH5Xe3hX8pXC8xtf1cKa94pVJPpuW8G1D7ST
0291f14LZlj2oKHHN5rInIoMOnYeU+QkAWVmB/psFZ9emLDN92/39lvnDDElvrSv
2NR9AzjuGBNl76EDwMW+w2+DYX0J7365eQ0G1AadstT64tkjb4AeUTD2KKxciek3
YcurbgBgMfbVkz3BMbUX2tuy3KM3y7zMZeUSrxc+0LHVM9EUeChxfZxluWIIak70
9PXHJqSlH3jdPLbRywhA5HkoUDHPMPfT6AaO5+dIEpPaOgsMt0pGI1xKv8Ke4Y08
lwEc2hAo0ogezE+b6N8tSIlh/6/GlAnJPPJtIv2vlLElkfyU/ZIwysRNPcTPYMhd
gsmfIUUoPce55IqdqK1eVIAYj8PJbBYZ//s6L86stNlB6JdNU8QHaShy1wR+otX1
DO7MQHzJKVwMnnqR8ucL3QqctmkR+h20s/MH13oRlhPjAZgwbkMnprYUesyxT2jQ
93LLxbJDN15SeGNrizOlfKNdY5Fuek3uNGtYs1Ge0sh8KIZ4+jm1lpcrVtPyWqPL
k4xHF0dJ5yUXnn/TfjjU1JuU6liGLoy73FEzLVQDeJTui3qq6c3+9bo8wQl15FN6
Kcf3k/sj6imY4ISmFR/xtdMQKEwaZYsaMG+6bg20crHAm7r3Ie9oAmjJhLZgDGJ5
981ky96dNnBcFPOn3P+ZXVrWnSHykRfVOKjiHcurjqHgj9Ts5aW/ce/p+zRoHzgY
70CcInh8kghix+dLU8Stmbn5EZHX0vImMDxfNAbBEO3B/C8phEmrT7vXU7vpfoOY
k4CuGeJKxkBMMoKHTRK4TIkDec75hNkqOQeBQDv8a46ZI/T4CxBpt/JS0X90MVye
J0F5pLgBbW3nWcw3fxlYkmC/MSc3g39DQ2xtdNVAtw8xzwi9n+al0o8mnc+Hm7Sk
GIIjJ0ybUmP1/pisJCOAWYqthxCbNlFSdEcoZcC2mTvjkFMHWhYIZ6N1lYkmuVTc
FAFVhvox9ZqZW5N28m6IBM8IjEssa4GLqm5Ursrk5cLHCZhyPnFVdBSokbxS2zAO
vNEDz6XDDpO3nckjTSdpXIDm3sCn4/gIoEzCVwisOygc5EmGI2DLSf+T2NkJ0fTP
Iv15txEks3yAUruo1WWaDnf4bFTuJNARpY7XZAWPZcvDhtWWHHguuy1eYGsrh02z
iXt6pZZaSNBgqVmiqlPC4HvgBIbwSOyMHdWmjR5mZVJ7wjwZjJKX9kAruBSddsQa
R8ueOmYCkgW1IelsnMUD6CA/COhU8iBVmYGSSipN6JdKjfP9da2sAV0I2kZKH5Is
mNZe4sgF3KhzKUIwtx0K/jsnuo6dGtmCsGz6Zv2KCHHlllBhGTPvcCYm2ovgL24X
gaMwdWayrxEdc3MjVRU9tWTpwQxRzSX36e2PVLA6xyG/RkEfq0hKqBRl/zgfg3th
g86iKDrKDlAJU6VL6CyI5rXx/Fb4rI+RVfxuK8aUwpiT7RWx67UyFaGYKk3FjIyO
7rO8liros4t4fFjXuFd82q26B9vo4/CB+dC2leV+KnZ5no6xLPONupnxXFel1X8v
pJ9p7s0tVAk1s+HnVlvdjAID3+pU42HqH6m4UUtBRCnktLrVo3ACjFg1sBL1nCAj
1JwbaAVmpRqEaSHGhZDFk7ji1Q7HaHtrPbyHZJYAmnGW9QaK0ST0axNNnbmKGOf6
tIq5gOJyAOjPfLVgb6ZrsAKUAjVQ4lkTkpnawPmEz3/pEsozVdAecXVY80A9eA4o
pSHcJ3X99U4oKqiS1bbjC1pEXN3Ubg7PDSSURKxK7ehH6r/OY0EDVCVEcOy73s9g
QbX/hp5GMVunzafc1a/G3/8P9QaPfl1QnJ6AiZuW98XSnsvoBMzInhECyuxBrQw7
lJsYlIUGyfHh4Ge1vWxsMl6st1VMMw84/0HbZ8l6t/IEv3Ck4jT0Dbyu5SEPD1lm
8NqE2GR8TZkUlX1ZIgR/+P05fC0qf00E25V/Kr5I4zgylvn1FRkQTBv3ojkBmElW
9B6ucV5+smgQyhIQz4rvU5ebj1PbxCHLslESF0t/8O59EuWHSjlg+SgXRf4tO6qs
vBDMTzpWYhwuANAbzKH1O8ZrEhPFZuBhbZ7dVXmXgrNQIRm+2vP2Gn8/IVRnpfI/
dvKuCVBhYseW49CUmX5SCAeS5UzO62+luG74bQvewczAKmPjXiM4pWVbJmeGsaUl
vRWGVDCnOHZ5wolADpKmhn/un2LS/xn4OagvmENm9/mfwM1RVxtWfVl9IbXr6i4x
YZJs/lMHxOput/pe4nATDrZByTQAu33yo1Hxff1ROpUiivLiKZIWoM+p/HJu01RD
D0Zz2iqhBDVwBZ5lx5SE7RAXtGDcUcCK0N5tUyiCP+6dZ5FgzCo113CnCci36zcm
mgnSyp3RXwtGjyFGfzGOpATyV85UoI4iY4LT9GxGH8FuRiEjW9dYmnX5oF6RxoYH
PRkRMjimmYshTVcqGBPxFgTY4PPz+6KqH8IwSNMsfa0cj+DF7CwwJkaSKXQUVEWf
t1EHvOU4lYxR5XLVZCe8gL8LAVg4JwLjkfdVFjCeTKpIEh9u2HzpFEtnzX+KBn3D
f6Ou1eb0O7PkmiqbW1L6JgZt4jLO+r+bk93hzbW03uKJwqqyRIVCNVpa3ftDj+Il
U2PoHcNvuyJmw82NOVuSmOMpxd+kHrNrs8I4kyvIx7BV/n/w8T/3i0CAdDDexMBV
kXqWRpIEyJb2xXkT8hcPLhRtRPia3a7z97teeI1L9ZUGe31a8pC+vAWOWOnp72mH
7NvHRo7zJJTldRY0KYUw4BqdtUz3tGdyl5IYSPQsOaDnfvB0ZxiN/komFzI8eTNH
mkphSD1eUZXjbbUejBmxLTQRP+w5DvrAIKXKEmJX76I41Dao7wvQUfHmnHFuyKdk
SUR7IftO8QeL6RnmC/D97rUs6As7lbBqK9R/IgXQb8pQmTTVBLsTKRxfIVv33BdL
p8V0fm6SHS0/u3vpG4ok/7KhuS3GanGapLhvTxbuNKqMQ4S8V2+iK6k5MnvdzUD4
0ODJTocBJloVfwoyFfX4uc0ehalx3pY1Y0WNQ4h7VeGQD0fH+2aBfEat2GdKwg56
1yOL3KoLZwBz+iIQ/wyMm8QtQhdmdZPl4sJwl+xfW49lUdUYXR3rCp5Xb5SDpOSY
z1cRQs1hXzTrqLZg4yvw+6fUfxqsyMLwa15vHYTjX1lK1ulHZyB5+LI81+zLlHee
Y0rJbmk9zr3DvVk9bP5UpAoRwcMBfpIeWN8G6J3n5stplepFtoUEL61DKy9JKmOS
mS0MXVQClLjoU0wboFSf3fQEuIoPXwgsqPrYAVHCDP30acBKO4ayevhqyp4kb3ux
m8WRM90Z2yWZoMVA1u9w19wINqw4400gNRA+zC8b+IHom1qmA53asZhHQnkQ7Zw2
O/pfIbxzEZ3YvQC2nIAu9+Bz16plhz5/IN8Hfmqnf++BBxXGa3KUP+D2P49gMu9j
FmMxWX3CJb/Pngi5cbPkmiSZmFtEe172PAjsD6FfLhNIL0UE+IpF23UFhV8lSPwF
3cDRKRlUTTnOIcfxjiPjrbAZWjnSt07YkGNcdedNaQ2NZzA5osMS61ApQfN1KtUS
QLokMrpsx7Ai1xP7kRK2RDzJDOrlaC8D/P2zYjRNt8JURvgAdynfqrZHJbZjjIZ7
nNCcP+dbTXWmNsRy5uf/XstcIbFcFjfE0wa+3FbXFZRUufvl4Q5axtKcwpYl9E5s
BhwUw2puIWqjZv/knXQgJrzhPYPCBfrRkmTvbsmT1vQQAMHXFk4/cYcLDq+WLuvo
0PZcwJcPbwzfeE75yYqdtV0Ewn74ndlWZzKIL4/Xm5faoMUXGyoo/C7rVHI4AJEX
z+EFd5sKKRwbxU5vT2qQriYJYqLytq4phxbL4dPEEwZgSWjWz5jApjf1P4qrGQfw
hwhYYcZ+RioZ+DtMEaDzzBj9yxHgNSFBrJKBS+t39rfBOJ9YucxSFPrGLrqVwgas
eVNpT2OLXUNfFJ8Io4M23Lwp/Ibvl1Tohai1kSH2XWo+8Sbl7mwK0XMNn5c/IBsz
22ukUEP+9zPwgVN/YhS8uuyZhnp5VsIprcoQ5tRMjdr8G54qe+xTf9gBeAyJJUAq
58dagUQmeWQ3D9d+aqX4oM0FLX24bV3EzgwDFXveTUUxOaDv2IPBLmtZTrugDqxw
4AmB3nKpam1bxwItpTILAZ5xHapJ5bOKXnSC0xL7VLHMM+CiEXla0pynyzbFNP9B
FAsPGF/hFH/lGxwDmw4OuSyhO0YVZi9XMLTxb4VJJG5i3uBwdldDvvpqzvS5HUwk
gaAVVsW2h8sG8+JHh9bWergw/uWZWqU8cs7oMtn4aoUPJtx5CkaVn/BjxrSmQ0Tp
7M0mt2MmIUhWvHa9gOyOFDBlTA65eQgT6FgmRFLkVi0IAJWTAkAliH4s6G3tne3S
fqxQ/on2GaWUuxJsUYy30oD7yXg0AGuFQvjWc2KtXvKW5FD44IjOkh51/RrKIDGE
tcOpjN9qVf0QH2kpvokIhpohgqVpoSTcTX/DNl4aVNY9sx7csiPX1FblEmjZVkz6
FreCzLqy1x9L8uJ7LHEqrpqcBX0tlX87hM5WdGXzxT8HoTj3/yey7kKiwFspgYqZ
g3AJaREw+765gxXp5ba1rjXDNaCfowTRX5cZYnR/9xU7dFNaaZL75i60xAvCHoEg
E1IytX4GrYlx9j6BtwxuaH5JX+cWQBLk7/WzsDaNo3PN8/uD4NmdGo/zB2I6yd44
RMB/x0TkZoAqW7v8sIMjFYRs3Ny24TSPoDu8EAsa/cbEAtV6RNCz9FLIhjPcfW+X
QTP/bC2MleTX6lIyiC0Dk4YAGP28OmGoomA6B/h6szs8sjw7yXHcRj4cs7oFxGl+
FujJcq1aBLuN5nXFFcItEA83foZw8y8JphiZUdX76UPU2pT6SYuNTvjVjM9N4iLj
Ou348U7hYaGkYAwbdSFkpw0dX/4TtbIyMchRQVGQOsoTt8yUmW94Hfr3LvMn5WLQ
yGZvxG9CurnsS6zBC2mLv+eZpYC4kKCFNfXiBZjLE4/tap3IzU5a8AwBxIPEvBI4
UKM1ZhCGBJBFHUZB7rKLP1ndH3vGZ+I+/Z/Ci8MqP+cGR+OwAbDnqm/DKnPiskMH
ZFlAkcff5gyMMyoWPxJbAzSFSLxoQZ+XDvmPMiPl9d0g1jVKcMw/kpnfS47DfkTr
VbAXpDtNUf0G7jl8LEFwsYW0A1Q4ZgbJN/2Te0fMaPw0Eo9k8Mb0+hFMALqyJspM
eh4y2PgFJT8w3DNS9skwMLqEkbwPhjdzI3praXy08Kf3GEmoazqEOGWb1Byp36Zf
p5YTSEbKZVYdTLULhhoNCyNBw4td1uFBliiflN0wo37IZyogJUXZ9CPAQ3YC+XdB
rXQHDKkeuzfRYVIjR4z2K9CfrVDeyvl1xWwQfkyF68YnEo2Fiu05TeKM9khCHIxp
yuizuorL0mJsr1MYn4kbbc5aP53/Acz3HPILlqdzNwIj5a7Fq3vsMtm1oGvsjMt1
L/wPAc0Jh2DA6MwArVClFjWrBOKc+iaQTHr8B1LTpDhhtMES3XlJnF5X0QBFIBSK
GV31E7KY2jXyKGKVttaRsIAtLdKEgfXYhUvCf7FZ1ZKs1UEkx5AuvRzNO9ePh0ew
2fkrPnv96GimDWV40g5eE72b39WQaoDSw1bLOSoqceE2K8qEBkdg1fVHAsNivSjB
ppo1xlTqwMUT/zBBDdD+inRob7ZAfmz0P2g13Ft13F+28c2i/92iZdQHYCTa9xC1
Dr3cXY3VgpV0kbTwHDgBEEEu2V4/0W8CN8MtefReX46Aa3i2NC96d8dNkadvfEgg
Oj7dGKwrRaLiTc6hkxFJkKyK0ytvG4/NYmGbsx5I83o7zAEaWEySysZUunvmoOzJ
rPBb5925N6WQok9R5sRLhzND6UliApnmCoSpHaxe3HiH2Ciq0vqFlh02yEAWt5rW
I8+VCgMJ/3d5Qzgyph4tf6FLfKvPXBXoR76+xYamQftFTX2Y1nTYlwJntMaorZbD
eSMT+MGVz+jCG+w+eto+f8RfoNamxtMpA+ds20L7McHQXJH+/iEc35TI6KbJUU37
AtkXnlbe+47s9nPd2bjjGVZkUXjy0Om84jqqTo8faLkon7vWZePiMJK38zQF6gfn
d+3SYz8LSBURVheWshqrYcCvCelgX5bfGlEO7o452N9/QqcLoz8Z1oPKvrJujFaM
QiCseF29RD0blwEXoevyotlxqCn8+NCahAfvsfpXl+o2ig+lctEyDEktMNsOaJ4H
xzKEWrayPkud291pQNfrJGMedT1ExFzbV7dmdsJDpolOkn08X/Tu/mrOt7TkbgQJ
434AKL3G17G7BbmizJ6RQEbRi7ymh+2ZA21grHOT5WubVCRvKuWyNPjziDMeeJJv
ezpCTQNgniVBVK0iTnl/fLWdYt5on04o8Qvm0aCrrxBWydmp3fB1pGR8Kv1U+u2t
+Ac61hZruPEJGp4U3yNdNPYGDD7b/WtBHXEdgWzOY1DbCfJGnPkdDIxp92YiXb3t
KgwJioyzcLWIIwunp9SnG2n8j9o+WDxAnWlLKmA65u97FbCbJo4naH++81AByyW9
6BEhWV9mmIVMR9KogZyM+cVYX5VvnnFzP6ql1m30/6jPz6aSkvGkaH7QiKbs/6zN
/A/Wvv6AQ8HLOTuhq+BXrvRzPelaS+uAasUNn444c8PzBh2redM3dKj2mhpmVSYu
tODRou3O4tmBmq9pIn8p1UUPyFmzV0IkAQnKmwe6cj7p9X0Q3hZKqJl6uTVCJ+fi
PBU0kcJ2pMGAkca7gwdKAj0xFuvgNRTz/eUspEn7jKYbLGFKzJeg6I7jhP8pxDoS
4yMK9+heyrjOyCYDYqKUzgMia2391skOt4RUgyQB5nNsbdcO5t57zsXWd1MeE0Lf
xHSTUSgwTftmX2FlKlZ+PpMKaCI7xnwyEuRwSvc/wLmFJj0QzloknU03/fWqBlSV
w3IgXGquevTESh9KIxbSP/TKZJkECx9QExGStmI952aIdfVxpuUv6wvHTHpJhTf2
0xAq+xZEGhozPZEMAa5Am3P38DN4Iiw5+FFiQz6c8pL/RWThRkusjffJyQSkkmIX
brmIampWkS5Mz8k1jhNGA5wN8MWEZRHeD0oX5Mk+n1r491z3tBnOJ1pidanmyBcx
PhmU79XLfaOt9koXfXucFWs+JHDrAqPUkQhs/cTIITz1DElpHbwNMOQZUzzPOFAJ
OVJPtVdjtHiNSjjbCI9+CvRHXEwniHxTARxz7GF3UnpUwjlc/osxERhGl/y10S9u
VBRBiT/e0nB5K89JTJUf4AL/ZU5XVxqd9NeIfZo8odFw7c9NuuGWFJ7g6CfuLfKp
xbECLRXqBtsP1RVAhEK5GK8Zp4arqFEby/EnX/HnvbBmFVvZI8bQ+F8obP6F/mEv
cWp+5FFTRPgM0GOfJTG8XQGm41yxra4zpj5PXjh5IVrmXjTWxIVCqNaSCioPYC4I
COMCeyDMM3L5wsOtbujtCMN/xlTjgWhwLcu2aXGqSfLWzq9m4uQeupBfUEcOTrBs
bSUh4a1GRdkWQrTjB4RIgSu/40sUK9NaZCsxQAfKn5Vq7z5gyLRdtMVjZPCynJJ2
IB6xKI+du4Wg2LXHiCtck5+cBBtKulFb91VdDp3//wnEulIc1Ex6c8RpXe7Grv8U
9yr2AzwaKFAKPZBBM6AKvLku0lyapOWUtqnGHEyiOBeHLCkKN3cwebGhq2NTUA8T
/qtiGlp36G0ndDbyxRusD7V8vJAGYPI39VABLh3QANLLH2C061ocwmUgXBhXveWc
KnQjQsLXpxzfuGM0yYYAWIs5ij5zz0yLnv01SVSrzoKErlk79dN0vPeQky/6Rcrm
nRUz9mbw8KQ7HMSOFaCfWbTpWXaeLrc+vaT8VS1PqE1NG8/4ois9KTacowIuFG36
EY3BZZpkdZ9eQU9abkcnFaf8SJns2TvGx3uwRhX1HovXoqzaGLozfTwrfhXwheA4
Ij7+kKaOJuENK9hCRYsYXwW490tn48Co5UyKFDnQ2N2+gXfvEimPO8p5yI00OGxB
mozknIxTvUF2nbFe2AjefVLiCwrN5qqiMjv6HZQyv212KszS3QLy75+Fp4TkG64C
D7T5Xh7WmOtaJoqadQoBvviC9XDa8mFqsbtRhFL1W1VwLIx7qil/u7KmdbvbIjtp
T4bZNAo+VqNgggQrEYxRp6eqWGNYCVxj7KKGxIZgyb09iNN/xN7CahL4oI21tDAx
hVXJLiF8T0mgnpySuxEIxzhyoY5nOOswCjKKTnVS/90BX4lpX+1jAl5ZSJLiv7Fz
BCKeLp5IKPVDextRfw001g2lgfIqb2uLGpl6OJpvp01sOWblYqEzlK/E2qtGHfrU
V446RZfjPY83GvZ2oCOvmV1WFb/4mICXQzoQsMkBBg3hxszUMLRL40w2v11zIm+7
ReuFopVkSjlQE3/4cZV6eqPBRMpdGInfXh1IPcn14kYYIW+sLIt03qbGxM75q1NB
VrUpmFW00Y0OuZW9Npr5+MdHYf/Z128b8xXuuO8cFanX1AQQ851mVnb7qWIld3gf
hm5AT8XEwu78gbCEQRZihHRKqxbk210Onm4H72pOOmHzWolsO1zqQXEFw6xxwfw0
RwBw3wuiNo7o787LMAjdTugRIwIokdvut1pKTDNWyl/+/JD1FoeeSQzVk025q2w9
/eARFBylxz3HRQ48Ub0VpNXzd7gvZG7kRqm5kZeYxw3+vqRJDuC4GwEOL5K67HIg
ksbwsWBlkTHGkwY6xdfKKY4bw/NDmzRpA81cl2Jv9WxkyiCPfidWts2VcJ4Bzhk6
qIhTt96hudjuUHrcot5ZWosGMeKYtxMEZCk1PF5Ko98RxHygEr/hS4llczQ7gFsG
uKaXb+OXL/ma+U6pjHNg7OmQZnEcN8Bw34pRr7KRHZtzuP3EOArHJirCSdzsRjaQ
kPCVTFuj9DGjUteRBg+/tgimocTFPT9olnrA5ISomif5S1Y1fY3kvNjckGFC3Zfu
pMkEt9ecwsLx8AWuWmlmQWuXesP7YKBLbJ4nRmO8CAcjI/NDV7x5Eo5YeYnM5fVX
xRzZb3hvrwd+FPVhlIy25lw4cM9WGGBAhrreHW5rS7IUoHnhgE1VrweBBbNsFtz1
bfFa2nf7g4cvwxpXJpTvT65QN6uCvfH+/DvO4b8KIy5mmMfJLZr/iQ6CixeiTPlH
JR/TQ9EEqXtmXTAkgcFAMtYlBWubr4v6Zf0HRbZwvyln0yKPtyox/9C1HareaR76
qRzY8OGzjoGRC/tX3QPvbzW+7VCJcwFKkLQ9bkgb4bMsMW3VbsBNU9H25Jo70CLW
TQGwgASQA4p9PDB4J2HNIodW7Ht/NCfPN2HZqDE1yenMzWKvuqRD0MMAPygXkj6g
/bIdlWgVd+glWIL8rIDy9hVnhl4C5cB3C2j6jsBhcBV5OAU/cNnO4GoFy8rOPLRM
zMS3cAFpjzloY5PZAsbSfYGm97s28opv4BV5Yigg8SwtvQkpR/Z72mNr36fpLeeZ
bFXoazmugo00jA/rIbDCTeHdsoFBsN/+smujmeOw7//xpYLJoj2XQIMHl4oMhbGa
kUtmxSUEWWqjUlb7jR3hmYu5k+B5IVwLrKvKsxyIg7V9kGn9TQaTOcnSxmx0Ldnx
3RfhVzX1JgaoAlUPllFcgpcCemgRvv4BrRZylzR920hvsUUWYePrpDNyAZqNKMjK
nkMirK4Ke4L17/nGBet+GJcu6NJhYfDUeHGHo9+5z0/Dct7K66makQpPhVy/E8gc
vxyW41u5oWWIYsnV+Cmb5Ryat7h7PREL0xLSxbRLXfUEnVyMCE/U6ErnqeQ5CZP+
nTUild1ddFY170yCqYJ6YQbvzYVlL5DL7Oo+40bsvZtHVQkNT76ESgy/2gi7JL1g
mSaU5qK+KKBsNISD1xOefOAbbR57RRF9VEyxvfG6pKFjpG8hNNe7JdMXLgKdp8JP
2sufgiq1oyAGkj5VPD1734xGMWXE+kdWeCGJe6oThBJjxujVs2K2qGNDykZqPbpx
vmhi+hvG+WZuyqz2wqLrk0tG+zY0YJM0asp1gSMvhOWBqQFF9CVF7Uf46tNLYMm2
RQ3Of3OG/dWngd7Rd2vm3VCDHDxXE9LduKKjMZCW1L6NG2OjFx+AlOu5V0XERklR
i1EmPubMQ8vqBY8rexNOXPoQyDKOwv914JA3rWuGvLiIhnlOKdB6Pek/4O2bBhkJ
0z2khur7S7Sv7m4NQIkYggam1FLE2pteCTFiY3unr2UmzfTbKnn35yfAEQCD9h8h
Bu13behR+/ZnsGvLDDzB8Ke+vPdrVjEl+tqQjf0oZDwo5GEBrDlENYKzn56TSliV
kAD2hj2tfx8xTSmuQ0YEKVZ//EE536MESPSJWy3B6BeaSmrkWkhMvVn6Vks6MSpn
axw/zjbaG+S5xor9WIsTADyYKPSWJyKKnXrqWQtaAuOoL3oJZyvJ4dL9lEiFuGrK
e/kODPC73ig/+YYhuPJou7KxIZ6nQSeUdJLEA/73WYs1BjhtulDR7M6mK0IaG7t6
jVvGVFSFSO2ju6W3cGDX3SEI4mxDLVd5Ysz483SBXI5KOBXvzmiNfDSaTlpOuRLG
D53/0FgtzR3+giOAeSfS4BRZYoW5OCVhWUX4gGNBVMqEqJQ/7XZf48uuLJlFr3wC
BGhq06eqoItyEODsJ6NAm6g9OPErLF75INeslhTaLYqk4SfwajTBv2fzRdO4qm1W
qetNWma1QWg018mfdAr0W8mu0VcSzv+Uxjee1YBkdE/UuOGBxZfVV/422yXTbEEO
waJhI5rKiVo96uwsGlemcKTEfgOeORfs2d6WTsF6gQSPNkj2t08gN79LNQUbkeXB
2l7cPZer+4Z8QpTTlxc47NWrbiiPNmINaf/cGyooXrDllzmWLSvKfiORVzkL0nNW
6r59jHnc6IqTiMbgsVWqOhmM9NM/B2W7vlzJOiudJDhslK+DFJlJfMYP566WTOV9
4YsmRbufqumqI7xKcW7AOglCDwUzqtfpJip11fqUxRVtfscpq0CwbcUBLTdtTFZK
No0IOdPfxbX4DKLuDNDyNSdvMXb//4NaYf0Y9aElnw5EZPozYfWfvVzJW3gYTmnM
fqF+Cx+b86aB8m3wR3y1fWo0OSxsGUTQc5FEMm7FQbZ9liSC6KNixTzgXY/6Tz4+
yICCAAvBCG+SqL6QpxPEmMQ2WAl6ruc064ic0Ui7Ob4BQc2WNcRFitjlxCqWEfyH
TIrQH6XK6U7BqwH9DH3oPgBsEG+EqKbG6WYI+Uw8312zKUfd+/L9oovFjInkrcYg
cDYeVEYZ9T3A95twTdPLyj8Ur2v1cIoJXI/Ax9Rh8rsriaagdhvsk8JD1fHRWSP7
EcGO/lmhAcTvXRTUklJ6gNhlfRiISLwdpIoQu1xpvbcsEAy/q8TCjYOFEqDvBqGj
YLKRImEbHiM59Pxa3EHWyXrKyA5IyfnmIYWvW16RgIiziVqazsDG13dbeQmarI3U
Ag+9s6rbC88ZnjUm+WX6qlNLAmYaEMr1KwAxEwoc0cbmyozrS9rLG8U2t3ZpYnv4
PFdnf4PiOh5GknaNPl39SUwzoUm9UygmXIjWk7m5tNnDlZUr3ByPznwaVJQllsZP
oGJatpPNsAyLQc5oHhurA+j3FHoCIak4zbVWzjHj1eQvh1Oi9OUKbdLGCNhLIqyP
ZDWRWChKYqnYufQ8lmbzo2i5NKT+CxaZbO4xw34FsAwFrWmwWGFBA5k8+cSVh988
kjonpz5c61XChqzm4vpOkLA5EajjUwNWcc+GC2xPeOZrpZebs1P+snzbMBLwu5hf
ce84kzMWfQrsmvUY2vIyr2p/6ylMcdLuttlcwOGDqN51fibxbYloq8mwKlAthfvU
sX2HiCHz9RRpWJ63tmulYuyUAxPEL6RkTPgoKRBGMif8cc5P7dqWl9FnJ87HCCh8
pziwJhqlME8kiNajH1e7qi+9ElRjXRHP2uKTQEc8zhfvJwfzOkb3STAIxGVFOK25
Hf1T8sgRzJys6P9FroSJaqM1qPjBRwgX5JMHG01gj4ZhvdIEkaDQmw/c01rnoajP
wW8AwCwEYmswSb7lk3pp5pypgnnZcJ8RvbxuHTquEf62Dkj8oiS24LQdFxK/Ryxd
iYauoNrd3k1WIYxsLoFvvuojS9VgQqtYtoi9WV5ji6WvFeOOYK9Dm+/LLkH/S56C
7wsZTKIQBc0Ofxj8Y9s00WydTZVwCg1AipyCICDIfeBK06sMhvEvwnVpFY1zwrGO
2tVyYDdpBdvfR7Gd+WDt6SjcFbHNRUzpeJ3Lue/5DHHNx+tsMjefv3SDjvYBRA/O
iI1nxhbw7CM/NZrZReDAfIMGya81kfj3Iv7x3zcjANiFYbIFMC6yfyeK0aYm79Xc
p36FtwLqdblrqHmJsNFHcpkvPY99/UJwNSXVnnJUrTyDcWqsgdKWRUTluwbBmJgw
ivg4/kIZ9smBkLf/HGORRsRL+tkLyJ2WOn1M56sVrfYvj8qLLolbfqas5EfMLdL8
3an3WJXvM8C+a/G2msBw2P4qMAHro58cbntDHTjGv+Fv41N5XjfF7yYCaebhsCy7
A6qc84hKuhE+gmTboyd1Gziib/qTobuZb7IsvIz/0Z5q2tap+K9NOYyEnIFYXy9l
86eVe/G/TuM3deELBpJNMsyyFKuf6ViF5d6c4+0Nq8E6VqZwLx2pqySPh6LAAhpX
mexf8pgsKRJPUEvLCDeVN3qTqfg9LPPBaxLfJt6DaNwuClGcpWsyRVK07+OAmCFU
UZ2r8euSl94Ta3+ae+VAYmv4LNXewbgJGCNUh3jNfYjWI6TUvdVRzbnF1DBw39ui
RWr1ntQ1t0Y2QzJRUtHmhCFEWBPd6aTwKuHYq2bJT9TplRLPolc7MqE/zMh97oTQ
JgaCBFEKdRp7dnDt5Yuk/YdUD+mpp/ILUuGsDEyl7d6GGY2hjQiiOAgRQxvd+yOA
NKnfbEAi+7BzzDfKfgMfhIc8jM45Xt7jq2GX2baTHeRM1Wtd7TXY4uSd/gbkDsOt
ISgx+qMl2rqyJb++V/Uw2X9tsRqHmnaXxQWe0AzwhDj9BRtY5+nkIrPEwJh6xV7W
4r/OYK+D9kklRoP5YCwmIbk7FLh9eQ6yIyH0KIDzVmlurtDZImIIHSdx3B0qA3Kn
3BpeWsPeYXRkmxaD0Vu3M8x+wT59gMsT35NUlayOy4IHzj00LniuUWxUt5zfPw5r
GXVKoOnHcuNP3D/oVwZlcRCSIT/0k4rOepMysBgEFoeeMV6QKzr7hsYS73eUvJIw
1oFdyBsLW0T2CTwEMmphDZHialSjI37MAnKizAl1Ben1O2rM+xnH7DItdqzAoEhj
V0lJFZLB1BwYFMO2rE287Qw1zIsQ4YeRXHZZMeaUTdh+9cVUKRIFo9yQ/P9m5a/M
AjqcwkfU2rhJvso1q6ZBWsr4NZsXg5/OWC6zE312Qe+Jx5ohHa2Pp91Lr4nKjkOw
3tlC6u6k3KOP5Pb9QQA5cCL4KZq4Ge2SGcz+5syLYMCdsPKf1cejCv0gFQLiGJxM
saupQ+YEpyNfc22eJCqfK2yo6H3fffm8fvOiodRGYWG03VSaIOH9TOrAjGJSgMMJ
NqnjapMb8coOGnpCv/U6AbxK004mAm1MiypeFDPRr67SO1dbWUsyNiC8MdYJ79G4
t4g41ZKMqWX2gOYyoolScyTsYiZoCEl9D1HdPponkcW7lLVQoQrhlg/4h4cNKQhw
xZIN4JbM705G4ZR7kYyyKDYpAnKRvvJRz1OcGiWjJPTqRfoRoLIUpxHPuZ3hE/er
8TcJ/jjEEo6xC1hFY2OaF9eILreRNjXiwSw93qT/z1vf0i+fom9PaCHk+gNFSbBs
D/agcHwL/goDahr1+in3tGu68WCiWb3sX1dJFfUai31djwAtEvQJpBx88cKviBt9
YHo5DRntyWontQ5hqBvwRWoZDTLDIpumbTTGUNYLI1l2XMpyRx5XoctnWXcmJTtN
OrfBRTaXPdO+1qhyGlTm27n30a9axX72NiAbYCcp7uGcBqPLTY7WK7T3KxBuLTf3
vLzm29LGsZfNrb+SvTf6RZjlWbIkxHyvAua4GJ7lMKBx4eT662s5pehMtrxJHTRX
+skNBmrRDfsK0BKLQmYfi32slIR8FUqgPa85Sv51seSZkmeGLVXs9l813ILn359e
z456CfBuQIJ2ymoO7eTGKzdo/62R9JudcPmhpRAZLEsLybRyFKdIX3xRO0n4oZPR
6YEkl3cE3cFCiqlam7ag7/PFyET+2EzTMbiHiqnybrHsHVoV+NyLqC2EMZ9LtlQz
VMfdgy5LnZcvmeOd9Yy1D1YHHP0s6AuTmSJKy2Yy3FFng5/wJVsmimvMhNvZIjY6
R+FrWSArvPKPBAp6j87/3UXnseSoytaAJt43UbieGmC/fsjEDPnbxjyqFbcOkHwY
G/V3O8EENlwRdkmr1DibD8Xc7f2qZqR77kj5QpwGv23s5wv+vZLnJzQES0KDdzVg
ccAa3NuRP/IRDYo1ZZDp8xdaghXwnXgmF6mNVJxnc8RlDqA8UjCyZhgHdHvNt2rS
S/x0m88ClMy4yfWSWWtXDvlkjM2BLoMpdNSkR98XfSP3s+qQ4DwcPZ10c93Ibga4
1EOHqY1zuVhnRxbA3Ohtg/vfId+rgaDIwMlHw9K8tOP4IJprieY7UcZiWpoKMCEY
AEGg9xcSp8rEvd86TIrZRaAifvr6IMzI0CZa4UoeNrejHVJQfHH0FVgyRzT7SR+M
+GCcTlWbhFTYj1faZ0M/hl+JP5lSBQEggIU4SyOT+0+SPF1FasLhDmk1ztf6eJP2
6agjpFXGffJFCF5ZwnIjCnGsNW/IFaGaXifTUGHlNfS9wUqUKuxcOg0Xc5q3/sfU
+CR8YyC7j0O8MYJFDswcw5RQBd6XwgmfOoFrMRmUb8pGOKytZOC8Zv82DbG5W8aB
gvV4IK6RU9jY3asR8OnIbUNB/PTiFOC5djVLyX0kZMAPa3DLoaen1CC1ewKWbhqI
xtMvZUg9KCgCiwS5BWVRrfF2yEVydjXYkITZOCOGoy3a0vIanXOfk1prDP4xUryB
Ig+1V7SwYcBUuFRdez4qTEDLHsTDQIlKNrDa/Mjy9BTmP7MqOshKckGF9K0H3lyU
r8m99r9zmHhSFvN8GWSyG39c8P9tq/S+Vhw3ERsiOB6CHxFFxj62eelOmQ9EqnSc
PtR55hIbiy7/iFPuHbWLP0OzSiEv9EAABQz47Epj6JH2gaZSUW+HS+LTm4zUQ+Bh
PabmYSPyax36Lwmovz/ZmUTgUOm90qLjX1PZYruar5UCc5D4r+rAqLyI5NjvBUGa
z/1PMYJTT9JzW4tANlN3KmvQb4e0X640FMzK47hBT5pjRFu5ANeWxXaMFLon2f74
lkXLcu8yy3KnW8rp7gqmtneZ1ZPeHXIcvDsCPfvRxwN9PEpqEesQ4zouvIn2lKRZ
kwsFu/nD4Ute73l+YtLQNcvJrpsvtAVqmxp7hJLxwlGquqtoDTwCQoAelnJOV1fw
DxuCZKfE03lqIulXih4yZNBykOYKXNlnvEi99ajtarHu7+18+4PKAos7ptVJ/g9O
bq7myXO2quu/FlUlZeKZrxtjw3m/2leWWl7ecXrOHtoTUiW/Br6CzjmpVrlciWDf
BGClCQkSZV3OD+JURzPYZyzIqhfNFxw78vbl4X2S68qqvuDkE31aafCc9vl5d1LN
fOXks/CPUyJ7k3YrPat5pLOUufVRsvLVwFFeWhJmj7cNMz3To7ypjXlwWNKJOXjN
d+8m88CUI5ekndg3d544V7ZuPcmuBoBTIBh5BC5N4RHx1eXI4Qh0hcgUyHmnF58S
WFj6QuwqEjf1Go3oBEXaNAf6dAsBMF3RUuLFajKVivgjDCtca5gCNHUusHCbraCm
3aVLNRgUi+eOC4GoHMKUTLicLxLJyUBk7uBYhDtg3bDp1p46M0eRw7OBhfADhnPC
A7+7UcyDYfYvhh51YVgy8/A8F6D3PHcZdvbgtCEBdZo8ufgjENa/6yJk3ccrwQLL
Y8ondgqikM7Vh1qb21XFcfOrTonef9T0Dj1nf4z691uy7dmjRgp7rlXZCwxOm4Rs
C7P4HUEWk1FNveNo7H2i1Hv/M5dv9H8ViBRmfhUFtlsmUBlM5afMx7Az/ig03Bl8
k37v+WhB/Kin2VoWXsS0Bl8ND1vTFVL9ZTQlFEINQk/xLYQevoDRm+KBfLW4vnt6
m/7n9T/8X4d4AJEqc8FnzhPUw82igu76yA15X++d7Of9Pdu3BsVts3C5dg+yjkg1
Ba6Z3RkunTo0lCHQJDZ7jsGEDrgEcPI0CBsXH5xxjyS2nVTLafSrEqlLaN+F8OLK
BhPXTEzdUwhId5BtdVvescnHWK22+vduY/6YQBps40kiUTY/HeVBQu+oXbF4ZQ8L
C2Z9ZusiEcADq0Jzu3W+CR+PPKi1un/19cFmMmdiWTM/Wm/lXQ260n87FiXBIKLz
hUEmn2QpoWWQbeMommlsUCnfEEFkYFqLDxqNo+E2R6ZLjXZus5WsuFLzUnPjPMVb
z6ZHnfGkkzKL+OeZQWc1qiFqtul27Tf4HJqNyTiJPZ0UAchzlFOZqtQFtQm0VFcd
XKfkuVriCr5AWlDim3W1leIytQ1GLO/KlDq7YvAvhvZzdzkVO9/Q7Wej+Cn59HFP
bTgAAHMqMjD+DNKrnNHdWZaz4fhZYzlN1Kikdcr7jM/C3E19fJi8KJeISo6VTJhI
Wdefbo6083Cauc4SfwNDw4KXDalut84P1Y8by7zUEDEuvjvU7mq5kFcvSoLcKaPN
oOhAE6jaiWHSa7ksrsN0PNmRolpgqxi4BR9ZPXOk7cxRnFtz7aPjjJfXul7jPMmp
lFyu5lmTKng8uUvbtZMix3J19BBwoZ9v6zdJCy/khdNM6pPlN9kEwjPzqZwa8mgx
Y91IRUl4M/3bJxVPwPMCn/wkyO2Pg3QRLszhXYV4rUxvXUFUxxKZdpSTgNU5g+Aa
hmTawDXXyv8Rxt9Hb4isY0BPsYQXVmwBCUM5qeA5bTsqA04OxJWsfA30DrGdE7n7
r5Xd2ZUMbBGnQG9w9GUxnCCKy18G26Af+OtK5Si1HqngYt394y03+U5DSOd0lQbd
kimHHr7FIu37Cxgl9XqhmCsehnK7EXzFyW/uGAAaDNijcGJrnCqf818H/eaVppLO
DvOseFaawKOF0PDYCj+7LH5AejZK2Dqt9CArUl4IxOcVXRIiIquLAxJwSFKXpFBX
QuISWYf5YvPE4jQShLUqlhmNCBL79rptT6ix7ZB0ccmPWZh9OwVpUI4TVp9fQ21e
Q8VdWQrkZTdj4tIHeH5fYSr+XO1ZBsDfKbgz+7+jel0jKnMwtDM33R95qRzRWNUI
gIqGfIWzUx6L08s9PJV3uV+Sfjqb5LUYLDjorvx6vmV0UnQ75aAcK4OtjfSu/teE
NONZvK9qakkqEHmyXRQa3amKbyix/EcCNor8QbNSZe4/8nPQjp4gJ3kfoJxkDYii
BGyZuK3LbBCR674eGIaKghHiY/KDHMraakQnOGio9GMWc3kZmQBFXb+9YPG8VtNg
kYp+rLyFldC9Lfldnin1Iwbsqgh7b+LTCJhmruEB/226Xzlz/HtDgI0/k5x2ngrU
64kQsYcNlPlTNXPZ2JN1C2T8WWLzF6J/5sCF2dPi96vCqEVqcukSC2Hc6rgaDvju
izg6/AHLXzvT9rjcPbAZVorUPB+KDo446QQP/+JorEAyhUSIclVQ/xQUzCtfwqWJ
TnlOf/bNfeCMRaSyVe9NcnMmfteE1A+k07DjQfblih3q8IbrvIf8WLJp05tAEpZB
kHmSHRw+Ej/IxPEfDf5RFa2NHxCpzdhzFajm9is6B+6fasirYN3mveLXDGNEHWcb
fu/dA5JpGcveBMbSxN6OrzgQc4bNOfZTLjQJ9IZxrrf6exj4pqaYHX3+dAB0yzmy
KfAzzO7DKGyBKreBcK0jP3PAeidR+3002++DtTlleIRApEpIYX9aZORYY1+KcK/y
0v7LybPRJm5BaRPJqMnQfpMQZA2xGHGN91t+kDoMnplhHwqBRW16KynKlq91UgQK
KZ8hy7ek5HsC9fxbvgjDKaAHRuWCcxNG+mFUpHR+YLTsYYZux8CF2TtsfNpjA3vx
Frq8467iLAhQdvZ8tfHCADUvcmYXB904aW5dew5Q3u8fLt6/FRnELzks0ZxRpwY2
fQ43TfLWiT8iVzXPpwwJnAUwUwhwIhS8eVBwUp03l+rKoHycS9LrDtDlp423Yr26
eQ14bqgRMRNiLupObff34h+EKhK6/ZI/ukEDeqbciMZTcc5rYaq5/wyDSeZLVk0i
4FsRxY4GGTfUM0Rd6l8WmsIPFbr6DDMqg0cPC5AiPbTyizBoX+Aye/Ss+LSYDUEV
hjJcAjOzS0CQiFgy4IKfsj+X9pZtPCS0Mcnka4Y0WhfHmiiduNp40uga759xbA+3
NqHVBvKgfg/N7rtdDeE27rj+p+JaS5mfos+qWLUcjQRRWV3UzUJBCGNgAHh7cqTj
eDCruKh9NwWjbFyPxu73xjnnLWDmuvlrbCg6dQUuCZWF1XBgqQTjUNb1S36H+ZWj
Gh5+nGKUlu6K/POlDIgOsqapp/JawTufk2xs+GVXv3aTjGywB4w/YvTB1W8iI0iR
t+1uZ6HbjS0+fA0QEB0t7BJyG75HHuQ0GLAyzbEHq2nBqh5CBXr9RDHYYxJvFyl1
4IiT8E+9ZEu6gYEsQ8B5rrMvR1sokZcwV9B8MyacjLE5iwW1QX43GzAHQY0FJLe4
rp55zpXqDHEG91/Xq2SHJL6yf/98bWEXUexUj+Ec+r+oKsAXkRfESFL6MERy6Ekv
uEdDZ3Z1537CsLnP/ks7Ziv+oSGbmjwDwkZUxBqvtKsq0HIv1FDX/zVIZ8TYw1QY
9h7MfeiCbyc4RdCo+2Mr/c+IQU8rUxrGcGP3wLAvYZl9QcTnK3yew1jGSWOr4oyc
V5IcyWrTg3ozM3FBtgkl+dQ9/20RYa6LAljn67YxByA56couhpzCtwnFM5W22i3X
baDjieMEsJYkgo3J9RFAp7CC2oTpWk1IDD+oHN3qMx2jkig6qikCekW7mEGpNt4X
ErLNwfqo3CQWADKA1rQYlPTZjH6tewe3PhgqwBuRfF6IScSTnZRpws9URmxBUEkJ
n1VwChdJ7UTXJ+cKttIFGBv3cWfmWq6o/tTtNBe3MAzNb8zXCqKLbkwemSDzLD1w
YQiw2Nmv+Avn9m1lJ9affgaHytyWt/zXgxYfMtX0JNGbu/11yx5YbyjP7NS4mKn/
UebGuC90mzrJf8P97oqk/wxhj4EjM8vn3O1ph5zS5RHFoZSgX0ayo/ZEzF2nKfOX
rz3jiYoYo+Yqf1ZbqqM/Tlwf51InMZLWu0Jbhkff6wnlallqxX6GfEMbUbtjYg6Z
7G4GTij1yK0I9d02/QbTWDUk6gj+E74lq+DbuUT/5yTq4dch3SwpsxFFCXvBX3UU
u3JFUjGlwHzeICW4JJ1qT8md5xrfXrbtjYcX1ljGr4mSMFyfuoFnIEOKWnzxpEzh
urbv0hnN1BucnnOKsq8iPkBYzTOs0DDR8Xp8eNvPjz/zw6gNGHauXJrlkyiEgUSC
CzOqC4HiqJg1NsQYMO2+OnarZ0MiM+Hup0YqHD+/Z9K8SzPUce0XeZ9CJl4k7bFO
opRVtHQQyxriQXKuGsNAozAGMVOFJ4H2ZE6tLU9r6/ZdaYzxjzTaq1AWAL9p/9tP
bJ7pYpn743fc0zAak0kOd6da+Fxr2Q5YOyJ5UoIWuYXi2aAW5wAffnflvs7Kidi0
6RQblt4YkxF5/LbBeYkgrapGsGnmPLaf20wbu4nwM8k53mngW+VHGvbjv/Nqx72j
GiKxSnHoA2aLK+rTN6pyKuXy+xsjY19ewkTK+K3zqyM75AMojXwcZnsYWIbEzkVB
kNUSO509gnQts2G63mNVuIo0ieRggtJdNRvilBiOWee9bQvJDC7i27hyrzKNMdxZ
hZamU0eonrD2l3HGKFeLbW66vrVGFJ5TrBa7aXJnbB8ghRURgxuIlbn81kbvNRHe
NBQclKcsLynfomXcjUDVSgvxwXGSXEO9QinPEjzgwnxRsOGSYF/C+J1mNwY2J1mx
wehLZF9EKg2Qe+Gay8Qq9L8jnUUJKmopa36unROoTTMD90XSHZDiBlKstFQqujF5
FRNlER3Wbc2nTjXkKfN+DUh2rfHQwsXrqslpCDvFnr3pzlFjIt+qcV9s2pV9i7U9
MJV897mK53SbXd4Dj5WPZPcKtkycE3kQ/T2wTXNFWEpHWIai+3rNSfOirv+yC+NV
LOk5xfx/FNrKa1X+gCDy3Bzs/Gz2kSbxDchJG3wQ/1HPtW6tIJuU20LWJtkqdLNX
ec8vvsl3AHaMV7tev08/kISpRwMb4iojU10RU9eVzqi/enYiB46+s6i8dRLL+U8D
JdUzjVBlKhW8hRFY/k4BHy46FICjQtm0CuUIP7gwoVQiXZm/mNtSHM/t/yVVAU8G
rr4UxHbvbvuvdg8PuiIEUKKJWqK63u8loHpUh8SXIFKVzyuThPStHFnCwk23sIQh
ckbDECVYMUgqzH4YLl+rhsRN/rprF6zysYnfaOua+r0DEa4hmLJ2fBinmH0QYeUM
Dq6ZMg+sXYYXj6Objhp4oCIQ0KJacyUtavBdzZcKv9f2Z/VUezojWzd5X7plYi+M
CaZuVV0mmZRju1t/oogA0cs3GAiUrZwkpXY4Cs3eV+t3r5tnVqFmrYe/5xBzQ4KY
EZWwqAWUTIrocqCczg0Q9hmgVA2AqIcy4s2tnaAI6c20BOWZxtXrtfanqLpd11Ux
DGyt3szpryRCw3/koYzy6uDDGlhPHzSh58DfkQHH6/pIRu/A6/NUWXqTxpC9SdrG
XM7QBFHAn4XKD+nN6BUN4KN4o5G3sZMZs+OYI15s6hH/Dfr8MI1QBrk3VyqXjtd9
k3H4EeAwgT27X/6guTEg7EHZQf3LaGrrX8+qW3C2sakHjMjNMKtZT7WXU1UbSjbS
GGgaViQmL9rjlCGFFnjihSJBkSxGhPPk9N+PXaafCjRlD3xQdI0DDryP0KzY2JkJ
ojf3Df8g8rux58nbfmSCSqTemU80ZxzltPrTFkJ/vt0jGPI6Tlw5lTxV7h+gXx88
NEyP8YqE7g9QIVP7zXtzy4MedwTeHKfsRrjT5Q0FADbpyDXk4KEZopt6JMB+0OZT
C/zCubp2Ve/NkW5utuutoOfrh0jzJ8jkiHbiORBGVREs8rXnKMfdCqIai4zIaN9p
VgJL+ClWR3ZmA7cjp8E4vO6Ko3uwEk7pTiQl3r2IbWoDANJxKDgWCi99Dh0djI4t
fx1Xki/mY1ehPzicZKTIxm/Y5jfkjwvMFFkL3DWPHV03IXK55xiRy4+InVEIpupd
xgybZ0aqchepy3hILfwcET/gFJx5fE6oofUOEwigQcwF7Q6nz+r6EK2plO+joaGO
u11pdFfOvcQgE0GnQlfV/FT+3gOOWYQnPE1ai3neFI7ce2iEvt3WabncfWhjB/xB
FNdtuGzbfYjl2BCBs8cidV7uX7ROH/U8Rf4CHUHJS3N/6fDwLWnx4v9tTfON649V
7Iu3yAie9nc0RM+RyTG7YD5oMafDxMaJE9ydRWnkgi3KvtnfnUYhKWBKWyTbrkTa
pqkJJtQ8L9ecMAueFQqQi2P3QWhEkD0NM6E4imGlBdEoIqFLWwqmn6D2QSEyO/YX
Gnxoea/sZgBQznemnnfn3oVkHdaTJKTc3Y2i1c36POa2fVInNtayObxPattHHvPi
gbVmq/FJymx+fCzGMoTBS9ZzDb0aHZ9bPhLQ5FrqnmGyWi8wi5RwKcqFSlksi6CZ
JGzzLEBDo9Yh0KgS7KzXIsdi/JDgdANJunWW0oh8+AdWKd+plnUF/aze9lfsJWRp
HNwodRba2RCByPE0V5/3boQp3wPdLvug5rqalcp+eKOdIkGWb/D16fKDMz//BE44
X21JW1pMz3isVJSC0YMDExtFNLBFL+XWjoagE1xhTWoapKxR6YElXceBF27au7pb
Tt/eGMX9Ez+dXMlFgsg7C905ySidllvKXdQftICH1uq1jcy76H+r64wzg9M/MhNc
MIr0k94xglPU8dEvGNVnZy679oW7s9Gf+6g2lfspp2a6Nv/PjhyEDqoVKRCVEsWY
WPbUiPOyqJ05DDYKtJilHnI0UPTor7skIOLh1un7K0eosPfivOct2acewXWAvHFh
PBwOWf3TuttddctvosrLGqxphEvRBHOo9mgFgTXkpJAVFAFjdF8+LOQt26qdsQt0
rPIRVftjTLDmKUZuI9hAp3MYfiBQkCaaslTyR38VqRULheuYS+9zQfb/k4AlrX6a
1zNAL/c/OcjD6ahY1K2XwNI2kg/aLmMGVih6JshuP6ntDRIXQ1mOVUPt0qiVQEHU
4BLwVQI9v3Y9Ev7fllTt/ENdOVF7MXuzuI9EVap8llt9jtcr/GIWFbSl1e9Uiijf
G1unHM4SUOjG1yVdnDDFCUGr9o2Luokv9Ujwv/3rgJdzzaJ7qF9AGH2x1rxLykCl
luuVSOx+TZywWCUu3PuHW7obyPiO1KHYUo61Ub4m+U1QKz1ebF4gDGB5Qf68qv8l
CAqMeXi6xrjySvZdoaaLddmFflsBFk+sfYSfJj83z2km8mg9yqEhSHwdjMH6CwBx
YbrFRFbnTrclGwW6i1BSs7/J3WPUPMaKs23H+PfYybM8gRfonHnjlS0Dg1ppHkYR
KQXNahO4JcjC/nWTDcJ3JuSJMn9zApLWzFoyjhLqzGTjklLzsofoRp2BegAOKNYH
x7MuJdWnOm06jGJZBX4TL87wmxjb+XlPD+0tMARouAvup1f5tKH/X/XfFcAYQ89R
O9gh5/FDI3fuPQHirOzus2AWpLCWi0O+9yTb48tk4IIygVxeRSmfhEtjrfBJuXaT
zHuwr5Wxs0yzM4KNc/qLEJoEoZ04RmT7mj7fj51kV72GER/1nE3uC2y5ZA93s0oj
mwrDS5QxzI4WexPity5FpV9Gxp/ROhlfGKnePWUlsdsELLWu1jXhAAr1AkEi48JO
WugqyGm2sy4jVpM0NQzPB5W5Tm+thdmKEFJacXWetJXhTkALWqsZSflB5a+/K9l3
FqM4fWZYmpCMSj8O8HBfYb/80uWJvQLbDdIVAF0SfkbQhD1/wCs7ZDo9yHMb1mTX
3+jECj4lVtmX8mS3duHX+w4Pd+0QcXIAdu4X6rRshzJ8506MPB7fMRyVLKLbgw75
oYchnYSr4gOpBakXdMZIN967jLyVJmKAqdloflFt1CJVgBno8Wkyndgkdvr3uKyx
Hnh4sCmYmS0quAc594f6F8ZkGNI8ywvNlDn52p+I+00p/DtzBidbD7oDb0OJ3AwK
PGPpBzezH5ZzAYeCGJMZQ9N0t2alTjUQNCvyO5b7sa90PiqJg/Q50MncsAp6RXRp
Zv973BwfdyMksFCZRNrGzmZ6+6QO+rKZQhOPMURwDGQPdx1S7bHSe8I5MLBjSYpH
nYyU7N9zcuQ3mQP9VHkJbt7DhqL1sWzJSwtYo6/JOGYkEef/mNi+k+VKmoiaF70W
k6fcdi2+OXpaYaJiG2Ido12OI7jqnyfowvmpIVRyVK5NiRGolIf1n6hwUI28YZdk
uQ7cKJY9tJAeBg8FyAQLf0Zyg/A4i4eIusflLkkvHO39YDZ+Rm/+LID3JRqAcrEV
2S5NHsNo8T3pvqt80zfPliiOiKCJMunPn15PCDiZUooiZ7EqSUu9sDt6GZg1YMwb
zegZbK9Q+Tf5pJb1DC6sqO/IcCKxL6iDa85yRDfaaTUq80L7Ll8HCaDCzoeW4Ocf
9gTcXtGMrPphKeuWlkErCucnLWuCpZthSOXVZZ5bwRIrj4Ji2w/H07F0SFKRLzMY
D7O7oiCN79Y95uyOPeh5rwgqtSdlURyiVL6hhaE5CtgaDZ3zN0Ha6LIMQC0wegY+
z1lhONWcZPFVEdDBNIroE0j9dTEC1G2KyqLHl7r8ZRywpyV76oPl9QtZE6lfMzmC
cYL610n24Dy0rafzuY+BRacGslIyMZiT/bZDY4BPwdQPLR2alUaUCRE3hENzkPjU
pZCVXaAZf3nF4ml7oBx5Rd6lmDK8/UoyuIKRH6wNoVHVAHG2z+4oe834Z8pY4ZZw
JDg73CN26CwW2nIX9MSXRxdBdrzeCQQCLq9Hu9rROzvWhRjcvFYWhDrWzTHqZx8N
niGP7MRDL+4PMg7daamKpaaAyfIryDs5PhKvLpZGCCTp9DU3xzp4uotSw/crnuXu
bK1bmwPJnZVRSkmyvG5gqXvUXaldtrHi0j8Z4dohfTQ/RZDYye1lBCq79d/cx3iL
u3Q77nPSetl79ZxPaXNfXPlEae2L4eDBJttejT252x5eK69QHBPt6EyuhntljFQG
2nPLwVxVR76+1iQ0h+bNqRJodhEfawVcThy6cmfC4MoqdabEV1ichMMp/EJ1CsNx
eQYNyOlxkqI25f3O4Qp34VEjmUvxViNzDkM7ojWVqZRq4cxV9xvvTj8RzUCdL0Or
ri24S/Ghv5W/d0fK3M0AZIi8jTKnNy3dTOMDm1tSoYLxKaWoH6WNIeh5/bpsKTmD
Nm6VnfblTFKjdRjyVmK3CDBwQlv7cUrwGSZIH4/9Bbe6CrUbV4DIX+sYx+D9+O3H
zLx9RJWIxIN/EjhArqb8OMN/9aGSdcdpE5dugQoc0hqkNTP8kSrZHTZeHbdNp3gv
/1Mr5BaH1ig/rfKithuG/yO0bxuTvkm0GK4azw7/e3NyHgLXaEblzLNdW3SM6ANV
x5ZpCwo/I87tTpS7rbcKMvcxcCVItX6e/cbxdtBAiBRs6dTe3VCync01Yf0MC6q9
1F7v8LaO69UYfF2h4BWiH7AzBeIKYNJkxuwuFMy/nd6GZ35eaTCT6zXjmUqa2+Uw
oUFUw7kHsqXjXXg2ua2HNA93QyZFJvS8b/gorqTA81oilYEZEda6ZBGKVEjhCg5L
4ey+5r+f0/S2noga51PJHmP9h4I0+VE7/a6ye13ILQx9PqQ+fhU0RgzEFd//b232
aBmubV64m5v4GhIkjeMLy5Ha+F0CX8XpceH6+vcLZjEMbipbQPA+W17EpDyicahu
yy6BVltBTXSr8pD02J3Dj0v99CF7cFG/j+mEZGvvYAT/wSx/j1T8Gk+rQ+aygHSJ
XHnFMC5YyJG/yv9+nKJiW+oyoHLLMB4HTF8ZbXk4arvfjrviBqwgj0fodBou4a7y
lBW/HHeSJ+jaJLYqaimZkqpJqn7e15WoMPUdivuGGT4ZuNGvURSp3P+CjqPeXD8Y
LNUYxtLptWokuSDWU2JqEMPVpZaQ2HRFtPanzTDqJ4R0KelW8jZ0/GZqgyefAt1W
ZFDgkbSDFd8VlGLrBPJlCH4uylEqEFUxuxpbcijL7IFWofS7lCxOcMixNPjOs5f4
QEa73l4emDmP5spBG3wRcOd4+SywnuAGc5HFq7qQv59mt3wQt+gDmdNvV2KKwIoO
cpkTjd2sgibYNk+gkUbTLFFdLedFiQe7m5JhsOQ8nIchMFzpgIVHOTJ7sPk17+AK
XLQfpFJ11T/OicvZQrukd/uQBUI17m4xI/o7VYsNUmm9aSFtUO3rmEe6zlwTG0Af
828fx+CX5r5PRf1MagoCNTC362afuk7/fWrJWL3XGNdOkXN0sg0JiWJhZ6Ugt4zK
naKL8Ee/GqVMxq3ehoGKjEl4g8btieYhnoiaAtGEEfLUzklPScN+AbJR1yHhmLzG
vftCPU8VgiGZCm9FzAqIf0Q88fHt7wzSkQs//7hJURd4f25SsRWspgfIXXxxqxYv
aGFVEV4OEgvzGZElZ+dMaruygTsMKhNG1VksmMPGuk/IwElnIDi2z/kALaZ1o3UL
ai+G7guPVt3r0JNk6kuqpm/Vd4O/jTUd7iQ0jgqWFXWJPok7vZNeDy5cvmI4zfRc
+cwlIugGNS/ga2ptjeGp4Wi4N3xgVM2p9JoPV/fo7YpTYK9Qy6mRLPsCFEOZH/Wp
iUnjAip35GheOnskK2WRdxgS296G//scr4RSdZUbb4VBpdHTVtYTNsQx7X5lRt+N
rdTf9DhHA9XBVjPdC4f7EFV2w2Vc4ABQUedhq2pm9aUkPzlK+Y3EQ5yoMzQ7LOQ9
R8rHL5bYAjSXRmpqsphZW/+lqgC1/vDc6ixraCyN/cN98acaJ+MpkmAlt402Xv/R
f3ZaAuUDKbkdacxGZLki7YrHtjCEg9je2t3hJUdveg5YIBOs8izGxf2PAiHK15MK
mRkhMOKJ2llse6R/GocT5jWdf098fyIVMYBL+LSPTRZloX0hg15ImA7XHHC8JO1a
CX5FHLTOHowTeUJOkv0sS+Qar6vzQI2xj8qo9HvE43leQXyV6G2O22oOfLDsNX6N
p8u+KAdMEAvlu08mrcH54LByGXZQ3Ml51PouqUMWMiKP0Qifr4xXVi3u/buzcn4G
llyoNLwrVVktBBr8NZsbBE+Od5YHSAbeYEzGCzwO/d7OL28ICLRHQDA2Bj6M7k5V
DWMrtY2gSy8nn5xh4j5ynVnOd5eE0GCbBNmoxNsvjF9KdMhU7nEwrVsCkSL3tiO0
OwP1/R3pKYyEy+EQp4C/su2wP+6F+862mc2JyrBNK6l4RBkyYxZ4/QMkQvAxYV1v
oqeCgeQU37pwRwdLkgKX8Z7kv/EDMmSAgnDLSy5RRpHWImJ3lQWoGl6GF7EWPtBe
CPYQ4JUcrdRYdpgNOxt8hSoWe2RX8cIazmk8S7HKLnTtTL6ESJB5lzPxRO8S6Jtr
IiP84X+82AIshC/rcSkQcEpyj4lUdFjcI3LazIaTUqxEnGhdhua8FOFOiD4t8CJy
ENXCPDzAmrhgP8uZbfSeOxhmdrKHdOgNS6tJ4dbOmfsVBnwvYSWB8eJznlsPXs+n
23R2fnEpfvEys3TcxMkUUtWfKbqx9PMBC0bTOmYDaGbPj2dWYhhCR5DdAr332UXt
mHBMlt/tK/eB6MMd7YT9FrfrCq9MVTZbIByCay/C2blhJdWN431KBDf7hos6PU+P
kZF5RduSg+H1wGAIl6sLQnkKO1DNFXTnZlgUNS1zC+kWVMjxuzEUwqRv9X9XTdgM
yFvF1x9opGp46N+0Rziwl9/L/LNS/vZQt8m5/r09PPjGVUGGAKkFSMg2UdoNcF6x
TH4fRGd1whWXJA8hKtbv+dAnEVGe8Ftl/oHAG+Ehr4a78E3/Hd3GzrIKX9WEp8is
ujSs8yE95fmbOdFk3fsdiFwM2LWwRUbQQS+7Ce4I97Pd7nvkdk1hHDNynsvalRu4
JjB5UvdsJx8bXe7mOZqAucQRmzZO56EPEB3o9Rubyf7K6ckPN9NRkLw4IoQxKgIV
6oFNJ5aV2Naxx58JrAHVBerm2wr/8dQu8KcUKqPfPb/B+WH5ycX3tyEEcbJTBT67
7Z+6hovCh7wGCm2erE4aSHm5ORWZxSVRcZBoKOmS3FXgGiKBq5qOX5fyzvh00FEZ
8ms2asGsiqqwRXmx/51tzHHfnfaffPlBwjqnLfUA7SUBffA+wPBMJlV6NR33uHAe
ihTm/xUgiEt1WybPuQaN0E8pKOffRi+ZaU6c4SoCYfDkEmdtUTfq+h1SXHGx/rIN
qeecurTsVeAOd8I0rC/bOqdTQcA0tx1fTCbV/iO6zwassR8Sg/C3CCY5F/C4Y9of
JUTM/aV9RwReNHY5rZwGfDaaEN1BBPTyVWOT7oCP6Ar5MEvWf+EnGhmRvZ7M1Cxc
lu5wvgJ+1/fZsyh24lcHDkr1Xga2ul2NOMXTthJxWE7hetPakDGoJUdejeUsJmiC
bSdaT0FDGmjwHyucXM7EJ2Zp/0lxgNAHhMbvZBbc8SiHQ28i44i2Y5er0GzgJyL7
tk65hZAGXZBJNhmN5mBrzHGToTnVMDq9WdPQI65zihMqmBDXiJKMPB7AG2PeEpE8
VfcsgTlX5HFUOeqsBNJoagAzM8z0NdKu8YSYPIljOIRxqrHu0tJafRnK7X0pUwc6
++TmeqQhf3ap0e8YfLJCC+tY5aT2JXjNhm5vKcX8yxe3PR80BL3qQ77xIqaufR5h
5zO7NjockZJFBGW7LPe6GSXRWOL1dEte8vWTXj8HIgz0GOqYGeMcQFkFW2ipfFRN
Wp5opQrA119mtZsvltKuWIJrfyxrQH31/5BPzklxRpdF4MvQkBfBRsharajk8hFl
qQqBHoNPbnTxPxrrGilPXLojxzRT3OyXZcB56ahZKFfJqxh90+eqqEZqVmEuEHuZ
WaqJ7E4DqlT4R0D7oDiLfthcAyIp71nSmFout0gEv1oCy4NvKWUsu54uOlTYVcrl
zlkvwj92VWasawloXiju5JMhHHrEeSQ/P3wN6VW96LMdxRQAguX1DNWQ164aNwvh
PdIQapLOnQqzQP4qaVg2V2v3t7h/NlRUJeUPzwzgWMZWvIUdVbu5VpxrRJN87oCU
w/NttfNNYF2A3i26SYg83KPaWztEFf1y+IIMEd75FCiwmDQ3Z3Io7CH2hGOJZeQI
ZbRbI9y/5yGvoRZ8InmFFTWqZ4NKcxo+aB6HymJ1gTlimQKb1A7Bbsp/tjCFCw8m
f5Nctdej0BdUINHYhkgFNW2y2KlGeQx7shnjrCoYj23Agi1cqDmz16Ysl+6YMe2f
DneolcjqRGqpBgI9ade/wtMJXLY+wUmLeWMPB8/he9Uv8rGEWWccg1z4Vhxlf6Gy
U5GhZcpnJomINq4LtXsdvoVvReCh+6yJarDGjbR78n/J1WO9W7fwJfTFGefsrtlg
uOeAyQf04e+HPD/et+wg02n1wKaKV9CJUkDlyqHcf7orITu8+pJtuxD99Cr1OP+R
27MDUzUN6mnNXAnTPUdWnCM5fLLSM0c+8FV9lfTa5c9FWOKfVTnuQFSJbmEKYpTf
QVd5vZdfLAM7/ef18dYjMXCmZnyts2Vf+YLWdQYDjWC3Saoqkx9vUfal2PMz5WM3
qias/FwKmzzD65qxDVObwio272faPDaLSvjyW2TRz1+ekICNkUw/ho2ZHCQ9cE5T
Q9j2Jwy5xP8+R2tMRMbEoWVviZ+yg269VBlOPcEhuFveJpN37MO/0f4mkVENIFEb
QeLQ9ID/n5JG/rSCBLUcQxwFQwLQKnxSzqnuNAPujWKApDRcmzilyFQQATHVCDY4
XXk5sb0PJiwmJEllfB2qr9LSzXnLDNaDJ84Z65NMYaIf6AIMNzjWc5J/SOUIBjy0
8uocGbHMrZ988d+4k6KiVMOXHGzWibz/8s+fZ+VAe7Ih6CE1jzDGKBlDqq/s0A+Z
HWTZCZqT/b50bJD+4TXxvuc7auEawIX8//+VGZnWDLCx/0nxhKeUfpXJL1r3Y8jh
Tz2pe2jH7t0rKqM7TUGspdEpeXQiZdGmmcmd4WHfXvp5sXDU+gaZcmjcH/KyozLE
bZQ+KVcDlwLq3ZPY4kPhS9odaD4kB1vxvJwZv3i9/+hvg68Q3Y0NkVI/IJgc44Sz
rbJkMbUSZ6o6sIagnItvytnlHw2oYBwG809OsLZ1iCG1v7DjfA0V1EouPPJLezDL
fD8dVC/ww+x/V9xwazQk8GES9bfW50G85ssgSsphJAEDvHxDLdALJzMjYwCqJ5wX
0vg39kfzkOiuIY7drboRQmmOUMJ+/AJqiGhRyW6T4EgeEctEn9nxC+xn/ObOuqfS
6hjokdAh1lnmMsYnB/GXlAlobAkXpv2zByd0XyGAcp2H1SojPsoLkKG7iFP9R05W
wa4j2Ubb4jbSWa+TliIcblyCACcSqvLSb022YevI/Brq3i9D7Us/CWd3ZYMBAxzt
izz+fN9q2OfImZrUOSmTEHv9xfwT5NkNIUs3g+BlYMUmvCfyKYLkfiu0+2rdYoR/
a1lCpKfOH7UeIov4FFVW4pmyQI9AXRHaTi9MnX4my2owY54W+cuAHg8jmngB9pvv
ONXbWFlIesZSCKqdPldMkPQmyMy//sDmt7qB8qKo9K61RHUQAiGcxl7hfEXVfJzB
fYF7hPJ854SE4RGghGXTwOFmMIhSgjiewXEIuczKOjB1A+WwNeor8O8VuDDZDceM
FP8vgn3rpFlHCa+zoofstvvr4yAzmwvNuftBhsOFGYa73disKI0jrN4ghfHzY7Uc
pyRut546SDHQVg5MmZvhXnmrm+UunGKFgf0E49e/s0GcSLPDzWFNKCX91676CsTU
n1qRUUNEOn5Q5QpmTxnNQyTfN+KMYZxMb9venp8zaKLRPQmrgnmkJZM3fmU/nshT
uLarW/OIDcKnGQEyUVEFrCFXS6nr5TvL40YyZuE94dmXGUq6svyoeaX7lBgv/FQf
Gsxk9TvPRLvyT15PUWFIX/5HaQpOkmjAAXaTRZTBPS+bL3yjHLvw3a3RjcpxmW5C
pJ4+gHyWPKf3CdZ0oA0ycHFU//Gf9jqbd3oKvLzQ5kEDnS4e+Yn6lgCRZ/IKDQgh
i1Qnt6jVKrSbE/QkLU0LXEDuoo55l7XmPs/wzGwgTeSmLTrTxFPOCCaYGYgne5R2
dCnxgJvgh8xOXSqczrE+PacjAE1ZAppqvNoKBUea/0xSR8C3K6ToedYWNlwvXP+8
co2suGAGrgfrEaRwNrUk8ICmu1YczNXSHc4LQOoygLOQm0Z/t9O5EnoqFXcI9PI7
BzJDGd9l05/S/W5wTuVq7gr+WHJlZq0vzbeTf9v8BA9T7qUnwwMMhYcQcgdX/7Sf
43qTJy74E7VCBSzw+ZtHY6U1gYsHOi/NfiAnosJCNXE8zoWp4JA/142ZG/JazcgZ
KHX5Rqc15SLiImCzUJQ3pzUFocSPxYsRDDJP/pATW8dzYvN7K2hZ7THg98q03fV0
OJyvPPKdglynkRZYArgW9cqXq+etdO6JAqMmdWiT9LKG7iGfJ8WyaC9p+/KqvjPD
7YL51weWN7T3UAbJGk2QRf1lHNWIqmNUmrg+pfdMnfZzFQEMNIOo4GadnKAiSRzq
RuaLBXMMYdEgc4UL8LQwyj9eI83NaS8pDc1Q8+BjvIn/mgL6icny0Aphi3i+UVzT
l+oFV8Wiw/wqaobGjQVTse/RjM1UArQUZhVWKjUxqo95N6JVwpLl4Y2fM3E6Ublu
4G/mZ4ylUvN1+3u+8ziNfIG4dIv3m4rhBtHQKnIuSV5U1+PXtLs/VigJT7YyAcqj
3MAmw1PW8mtFfjOd+qGNON8iIjaRUplsyudF3xmVYfOCrE3nEFr41YkNPG/jYe5x
casQLrSjSWk9taegd0RSh2wXmCXn2Dk9U2FVLAux+1bYa0ILZKOoBrB/bz2CzdqS
vHfk586Ch+KGFOo7XdHDRvgaSdKrozVOxv7vV3ivyhTx7A/762Nr8EI4yMnAwMi+
Ztq8iH7rtlkWIdVqwZ6jEd47Csmy64jvrg6MiXOFtokTUZj2k2O5seT5zAybaZTD
GQB+EG5zZKMmYy7ujpmgfIFgsnpA+nFDXcBFnfVgccpnAOchgqQ/cEzsXsql/Akt
zTwuTW8VskDIkUkP2nvChsdAu16JnLZAIgrcnChSoyLpmCnRSI8/olPpk/wPWR2L
L5FjmnFwui7ddXg2DPUzbUDR5VO27PNUdxPJ11cOan2WftJaeaQf58a3dkfGBne8
lI3e4MCqUSF15uwoBoohGfWSh0QP0fMrx0ja/dDL5jFgoLHN8vdIhADaGfcSt66r
LI+y48T0TYjrc+Z43XnK+1r86X9HQ1DkT2NNaSzna5j7FfNERW/3dQ00vrZWyd6E
kNP2XuJkx9H/+SM/R9nUlM2k8kMMTmKVzJcqQ8v4b5vkePTTFO9hX4jNNQaOS0Wd
+JoxL4/Hg/ZY+C6VMYr8Vd3txTuDxQRYaFQDHoeUZbsmMaVFV3oGKz0MP+LxH1d9
rmE9oZp1o8MT2mUKyW+0IO1AfpvFlaiIRryZTyY2/ndgjfzJk1SaaRlx+rxHLGdm
KxRcqgBQ5RGCCKzaH6nsFsdfi2VxNZOBvOMo1ikWMQmvKePdEMAgvByXkQCGXD+T
6PLVavJCHTmcUdgrGqO5AVuX9mjETFfgQUNbf5noY7YF1ea7Sa7jF7qxCEEoXFA2
06O3k0aTRcaFk9MEMHMI/vRol83j6uN5OEmm8ChCzy8uwjqfRPa1MczPzNygEokj
0EINUiFP8bV0BpBV6bCX8ex+6Jwh/p8gu3+iJxnMsP0S7G02VUE2lhJ67fEqxpAk
IOhz4YkoRQRjLVCB/4MbbvSEE0SJbK40FboCn7hfrYp9TKx/wSsC0IcVahkZBtlp
+gHxsXtZ6mRfhU1EVzPnXNGCsWRNG4XvmoDkov0Y9gnOAQp4bUSz1wWEZRpdzRIy
LKNbVGUshs9Vu4KaUHUjfkJtyCC+W+GwxtI1mkFxPwyoqwKQlJPPfeG+FQjlFsIK
a+dtmpOrbaj6ZXM5juR7O3qHoaxoAPTFyF2IIyx+5IPfko4AjmLfFMO12Z+WOoel
kB4eI0IrgEKQa7uwgeo97SevQNfRZBVfWvK4NyzVRb7K8hKCbn9FIk5C85MlW3h+
BaBOJQxVY420MEDv5lUiHChaciNcMcbGI9oOpwnebbccrOTfEEhbM9afTJjjexW5
3O+mlvVIRBAeYrsuwgzrsJJLtxzvAXiac3/FFfbxhVVLYDdxUHpmRohpIYCJC9uM
+7Nk5unlp6jt7lSrF80VugQKODCocH944tx7Aw6H2AbNYYguBoPoDh6mQZIvAiG/
bMJe4qHUxTILWOPdhzxDfoy9MhFRRZA0+AC3/yPkhSvhau+TsF27c3P2t0V0t/Ey
0ci+GbN4J03PbO0wdZROdsGyme/jMHK37dgo947SGEbmmZeC6bqb1atpBZWFHNQ8
MzE3oATbCkiqeaNx4CAD3WHqT50Egh6nJ2gItkZW3PlXjyYhEgKjJJW5tOhZY2MD
putPE3k3GvqflOI2TkwN0MNBPciUKpDebZNz5xGJmqGbaLFcjVXuxwYSgJpzkezb
DCkg9XzG6pGIL4Uf+b90g3coosIT4yqgX6MiSZCotY0TJ2+piTXrhLQHC/21dF/Z
DHLhwugZmwLe0t3zNfZICXd65LaH909TMP+d+Q8XPWSZPz7ri1hkwY3iGdNOQvA9
ShutPeKsMw7t31dqlB/ibkkfxyXnuYPkWenARlxq9Pbl8AyPbrT93MbHgHkEkjUa
d7xtvEn05KwBjehko9YF3ec52oVF5D8yoaBI/g6BE6F/iZBgQKBnNjurfsUv/77r
lA7KNRL4UOkEq329YBqcsXRDoDLTpFcbeIE8zULcPkjc23bQlcScDm8D527yfcZV
Y4BOwcIyH+aJ5BQ7oojNUd7Wbexc8vLbY8bKTo8HHAXQxP0ijgcJDqJ1encYfG01
FiiifC/uF8vHkE7xV+IqML783FlzPrizq1SOwwnIbv2BEZKB5d/K4mUq1egNNOOP
hQVjGa2B0ta3FueldVcu8QiKzgbWleoxBR4eLtldxxwxhLQCBeX5wAn5X2jH4E6m
YG/zEOb6C1Cc1ruNfE734qGORzrsciUGv4Q9Jlc/Q/nTWQaS+U6M/yRpGD8j0Ani
IfRhsl4/KJDlO3+h/5cKiYPoXy9R5HNh7CISEMa7iSWxMlstx6ycfpiuT3llTvWT
XYvTCN3iRcVEAWkpJZ6tRYsr+1SIljxzyt9BtOxnaF3lx7heByL7jkLvWmD1DtbR
WP4E9bTiFp7n4M5iA1BWZzAz/z/0M+XpPoY5tCRrFvyuYKxppdOSroTncQV0FzPg
T3UipsRsX0AqHBuvSF3Pz4HIOztJSuIRCYnz2il6VD1P0/Fz7WKVF1nycV56o7R2
lO0LRMZErTNg4dNDe39WBF6QGtW54cFUZsgv6AfZdYnInElNCXsmWF/jqXZXVuI2
QBLSbvceAP8Y18+ED+ikrYN3DrpWvg6RvqeeYwZlsL8sGv6C+Qzq/R9OZXllfa8D
X4wZo27nLy6gcqP4EN8Z2vDaBn13TTV4qZdS3S3By2XkUqGDr/wwdRuGgZo/KxZR
TdXEMwsYI1rKrVUuzGY0f1MfKEKmlQ61t0Fq5/DfCn/1kPrSK/LkOf1FufJsElmP
HCcZEkXueBk5+pMNU2dZZy4AJFt5TLC9tjHRVECUgoxm4nAJu2YWP0oP8gMHWiTW
zaTtOrs2thLAtJdmUYwqYFmKK+xEtqOCtYMU3vOtkd7PeCe6mv4OPrN8hkS/EwuI
ehQiCbRD3noBT7OHWILsJGdNqBDomIEEN66JzxRpDMX206/df5UYw9Fj5Q36fBhR
AKybUwmIJMVN/2bXabu3xTkB3zydx+WuGZXUqJgRuvKZSkNqID8v/GQ/wyKaJQza
DBwQ8UHXktzLVoPOWjnzoXLCLIl6Am7KJTGXXJdMwvdSoLlqLhc6G9g1emU5Cjpe
ynlxWVcNCvsXsJXXCMY7Kf6fGL3Leh1jIxJ1LlcC8A5R08HYFzt3EYAiJmWUFLAF
kPFLDqFD4qO5INbpsFFbFKnoqiMk3Rt4rXRU+oyCkT1RfiPa3HaKJmBE8s6spf11
UU1nN94aVHkfzmu+Xw9FNjc34XMobdjLs9kF5FcSoqQQTir1fQXDwt5FAAMaEvQI
vD9tDNX0ap5AVWWDro+daNYYEzRHE11ZJba/7db3vmdiXtFwjs5igaqhimNJRb1N
nyKeHzHPvgN3wUNTtl2XbLksbq7fntmYryD0uOrjsmmg8DyzB+mocDJj55LtPTXg
fiSeE2bZvqVmerYa38NNktT2RCTMQZpNBVPYTJ+on6NhO7yVk4wXybp/VV+zJJgk
3c4UptZovbC3d8/hXsjhnWHcRTi7JtQhHwr+XM0fybXOYXIAidhch9N3ii4R99oH
EjGDnwFEf5ZsLJvjnmnPklk/HmG3cVBvxhRF7W0MHidZAsCQLFOXJkQKl4qcwVss
AIgezbrz+rLg3KcK5bh/IPnVHOqLz4jdpFp1tIOhfG2rmDZhHlN4xTKEYGrbKeJI
Kp6NgGF+34Lnlfpb6i034kJGwxRZUknM2HRXPETCGjnW2xwD8gr1Mip9hEWp2ScW
a0NN/ZNquZeMrVtmMkKcGtM/mI9EOOrZmTcvg2/YMeKTPKWwBWwHh2v2svGApc2r
/UZxCWiOfD1t1VsBpncKp6fCrqipr23J9F643zScfnwLKKPvE9CALaT3/kJ13lru
/JuvW6XxRHOCrXl4aNDq5e66axMWyyZaP82HFRpdVvg3eX952ypEq7WLZ/vQFWUY
s0kx3iWufEyqaogiSxaIAdbYZE5LGkaLQIEeL9kRv5Aw/kEB/KLYIGNXTuOQ3afH
UhJ/PUmJnGJn5afXD2Ag9Z5bPd63jGmpmFJJZN6sy7yB7Pb9sd8b7b9zwlhjOHBv
Pk0VaFkVI3XCfJiSf0QywSIKfU/4poaO0cvp1hiXGW2k/EK60DaugLXFaTWeb4cM
PFlcoiGxHItBhy+wnA+1369eTXMPTMP38/2ORxi7o4hFIsMKTi9NNFNMmdeZWBK5
WYlzgE9wGam3L9bbHLBw4YCkG9u2fS49Mz+aUIUAXMkoGSJ2coiKVAtMP2rRoEEZ
jIhySoFSdVlKKBgKUt5odUsk0+VkINAS9v6t2JhzKZJ2JNnApI0BAPXgynTc5wsz
BLt6ks+NQWuxRHDEkmOtg8p/QLehcBNcEWihzQLFxpjniBe3ToTP7AjLu6NPK2UV
/3E2HD4N6QeEsiKeiryzyQ18id2VIy8pzCAM4uPyl4XpSxE7qlNsq19RthAGu6ao
p9vK4t0/SXXvKOIOm3y1oUFbpJbXGPjRNZMXzpAJNlck/CcE2TsVEbR0QA72X8Ru
5q1ygDOlHoD6q0b3eqhZ9gsVSsTVsrwJLbHvip83Zkf8FaYc0VvpNCnSyNnFkwVn
VS8wqDdPtevzuKhBznrS0a0XwRDBC/iJYMgg93CYSmN6NKiwpEyOswHEvTHYtYl+
LDi09OUARlrTubq3E9ucfEa3WBPKtauD6Tivth6JrOVZ2jjoOiqnYn2idBw2sIsI
10RvphG/3PxXalqC+6WZZkgiiO83yGtR0UEJPM0a+f89O5y4r9ywXm4DmVNdo90+
AkjdIwLwSPKYAgdxbNIqP9CuG1pNu12/pxBHwW00UuXOETUUu2DLkhB00hiIJ66K
s5qZyRfMSXY/t08SAPdPLcY9ixWxQapm74/12mF8mmFUQ9NHK965cPNLJodlaowp
4WQp3wmcUPpbeXPhv9y2N5BG3h4C3jcH7FRDGQi/n8Ph6RaRuxai3oAlwen69zwR
GvYGbgHHwb1owod3DViFdBTOZRKymUJu6J8KgxxhuxkdC2vOeiWUSNJSMqwVvSbI
U/9aYZ0SBSzEfdJoNPTs3My6sZxq4MbDQWDkMxPuPw5gGI5lmaGcKolQg+8unapx
uiIawDfeGs9nay5AL82kXay71B73YVKIzhNtjjbtvN0jeArzyt9yXTsC1l1MwI7w
FwjGOEpnBIqY+6JCp9QkQtEl+8XnlJf5OXYqYe03NT/VPJoStiPajZ4ZnbcQr6gO
cugBoCJuJ+pKLGg/Mah9DYIasT54BXh0sN4lYHaQOvRMBxLctXhfmGaPKUQoOY9j
j43uNVvGpzzdG3ur1y0Js0GEAR4MNH826DFs6u6bHpVRNw1YWWf00bDX81eovOiT
KrdB7ngZbTVTGWHTZGh66DozV7sz/6Qf/8a6bE+74gNiEqgoBjT8fhTSGC4m68tG
H6kIwjQMlaZdybD81Rwe0rgwygFJiHCqacZlKs344p59/gYtbjC9QtFrkPDN7gzE
B7YFspFh5yj2WN8WaHghjkfS6Q7qzFXPAm/s5ppPibcWDqoMMeUrT6oTE+7cTB0D
WbAlaR/nrYpEgN8xPsEJXzNq4WjLOstsJoydTqvggrHK0N4UftunJlvtr7XNZS/k
ZPtd53fDAHEJU3L7LjrJs7vzo5OuKQi0syTkh9nlHtEJVlrqSoB9QtAMSjt46/Rq
6ROzosFv01Cs1shLdjTi+OiLr9zgKmsoMV9vxI20NrmEFqefMtNyoqiWHhQrCzLE
K4Zjslpd9/mAPP0Gnq/OkSVtpMuwQYjZHFIYWVf1HEDqxvFKNz9yzzFLo+bzTsbM
pujFsoVk40vwyg2UFRCB1szCN7AyJKiucCOfUTxTvdwOyJQi9QrzdXIeG03WTRyt
c0WLKTCDK+F9v9SrRdqLzoOHXWGh563wk1pWxl2iw8f3e/RysK7RjgD9j5FFB2aH
4x9LvMvfLFIdJQh8bFTFDVeIsi9p/BhQn94V5dQAOkxV2p9OsrftPGDU9Jbja0x2
Fl/ai3v+GJa7a0oKvfLnuAvtAX0yjRoKAKEcdXhpYBCU1aE/QfZ0ueQPCKBLQuLe
4I6C76879MT71yb2S4MliPUgne129PfC1ZgIT+p574HjsaXDvSmjCSRNzG53296f
0bBCMRHo4o/jy7zf/pE6tcLyinXJ9NyykHaeXu6w2TBv4t+GXUm+OuMSN4TAHkcu
5lfGx5x+O7izPOct4pWy+vxpqpysw3HYXinxJMeVt5IxvWBN0hollU9kFke7ibMJ
b1jMOgGUMvmS/d4w6XtNMXKF/vmGcnrI5ZKmeDSt2vL/2BWFc72FPGfrsw5YwnKp
+u22peIc81Blk1qEvvWVR1rulYyzeigSvolMejXZu3Td0VOVaTXAAutsFibjeO6W
FoVljhb0gfplj94Ia8GWUy5Kwp4gVvc0Y1+2a2XF5buDZyP/yuPxfTxjgXPp1xWQ
jvDDTS3BWuJ+DKonXF7HegdPrDF89BjxQVRzGiZMx+rWd/HjzreMcxx2q9cFN0uP
gVHXENUmDxW5DVdpxs6yHxCVqFgn1tqwO9EXqoRLTsyHNkE8LBetwqVT0AAtPw1M
6iD//MaRHbIsEDDXO6U7QRPm8edRHojebWo71Vc8xAUD1QE7os9G4rvPP53gacRo
1sCULZ8rkl31MeEUa7hTwhtTaxL97yG4LlL+M23w5InHibu33vIsYnxaSQhYxObm
3tPPQ4AQ2v1cPiAw/P3ClIwS0dKA+Z2QOnBObbLBhvB1SzHWmeVk9CWI2OIFhZz3
VQBo6zJfPREbCuNBVAkgBoDMToM41y/ZBxVG8k2kSj12jAhiQ8G5YYmWSQgrPTcr
Dhtrrhm88jT6+T3v75m71l2WoOADLngPjZELEeYh7DqbWPfxQD6YZZhmuIWyfufX
GriVH+7unDz1FFZ3Q2soFKIyisc85IyEDfAxeSujBKR7HW2J7u6tzh0748FjWfyM
W9kjpLyMVS9NxG1ivPaWUbO9w4g2zsQCIccLh4h1vJlRehOy24/5WQHhTOb2daaT
wZC/JGD1w3wbwzw3tph+xmugULIYH/1BwFvi8xtGXHCowqdX6TPG3w3gyemV0WpL
nrDME7jpBbDaeRvMyDT8oKgCM4kxrCHTa/8UdI3ZQggxRUUvj9o9tbObz9DLHF2N
SHgzWBtSIzmMiE3NT+doSZur7q0G431lQAz8IOJsMaD0AzsxgGd+1qXhuUPIb2X2
P5UHliWVfpLQ6daio8jQOxMpBN1aFK8jPhHZSI5JICHp8P8qQzS4TcAH59wdOKEm
oRq+TYQ4oaoSM08tq5BmTgekKysgRH9jgIDaUzVrTIedQQ4NP1U+KgGmgAhiqTIS
+So/scE3GmZcb+gd4ThoI3VTiCEEcFdTahh56bCQinTaWRR+e4j3fYLytVtcUO3r
AcTgGqXcjo3BTNylwcg9pEc3lZIRTiMhp4O1gDJ4kOb+B6ChZLEqXsJYUKQHC1l7
EOFd4ExM52VfJnVI0yQG8AaKJOT2qMox6ZwaICdx9eXqvrfPOIPpj+xTC+3ZLPIV
kVIivD2ChppwjeXAVd0zQoEHIjUycMwvp1i58czPbhv+GZn5p601UC2gPMmaxL/4
8Cu/Z/fBOUMy9cQhU+E4nkkwMi2B09TFDV2BJCEZuZeqMpQfsj9NArHWJkXm+hLg
784IpQNkrgGhU4VupzUaJvNifAm8rKmhpAIUoy+SM5JS7i+VAQ5+kjLLaa+uEkNS
GVUWmvhzTPc5lK1aGpuJYoMACXTT8WPZEz1z38xuED762DibP1Tpro5PXk+l7adE
ahyaudj/iNhi+iVOAKcE63oANi04YC8vV6GfZSqQDRQdw3eLxKJBwgOh47g+J4kZ
rYPqXShoPaOeZS4e7pDDG2wz1mit6zL/biyBlNioVvQzot19xsj9OzWN+D9AHU82
O4xkmE0enxcaKP9PXCGcopZoXJtl2E0blDQnBXdMpp/YfovKN6wLCKfc8GCBTQxC
VpJabzoAb0uytE+lYbDFE2w9p6Cgf0OUv+xb89UTzstN/4PlQVAnrp9con9GUspI
ptrrc0lV52qnQCqtm7N4f7G15OIkYVXfdYG4LqiCgrxiu/85DbVVsv3tOVrCDfzb
gUFrS1CT2IzaypPhRynFVGhTB70S8nqGJC1KmzRb/keWnLmhkyMPki+LPPoMpWKi
Rr3tQUnc1s1VTMemqxAp0ubBPORKYsJXCRXFvrLtfGy0KXlnpGs/hbzAIUCmWykN
ujvdkuibw1MHr+xdoWKEtUOqswn8o/NHROEJk/85jLwbaU0FwNp0l5jY6QxdwtCA
UIoyUV/4fsTgtOepBOQ8hrj7MU6g66RLmiVbsUqRllW2EPhNZcVZJWalKuezK0ZL
bvC4oa/5a4vGZEXEFKdTIUnM0LIa4VtiiO4JoLwSjn7QDYmp5++0HwBZSNbp8zq3
O+TMzI41CKoc85kG2yPhs/ZwkPSxxS8WMxZ26vLDcUsGPDqqr3TjK7dm+3UmciqK
/6oWggOsDS1/GRzAow+uqeNouFhO5s9NDsOAAsQOXxUzIfLYQOVqAdS1tt7dFDJo
zuF9+lpsLCsRaws5bDQHMwqSmagLCuE/Ryeml6QLiNrUClKGxlNd31KrlZgaXPju
pfbPh1AitxdBvV3WNv9tP58KgkMYt8aksGJsvBbdOM86kUfu2B9rmWyijoUK709m
O9jf4nj4blLaBhQPsbYcPqAUWLmQD/VQS21K96t7Kmb0FixhQPzagwuA9v9bepK0
zpR0EZot8nkKqkw6R0VSA9uhH3DgZLNDjvt0W9PwAiT1slfqJ1bN1NQ6sZprUw8K
YN3Hp/893PXBUUnu3rrWB0/+0N8q5wA+uPq6SDbEgI7ksI3vPN68RMCq9TxNqzgM
LDJu234Cre2Hn6Onn15gR8ra5RRmeGwamY4dTOKJaG/mSelVa50vPYB0sob1vP3G
Pck/EAirGHxMy98PIlIzPBNrd5T8qpbN+/eZBBKCTq2ibI/SDA03RhTZnvfNjnzB
lgaDWcp6xEDc3bHYMtHgDPXax8vWrh6RDhadQxJ7NwDjKOL4SdXaPz3AUv3ldEEG
rJ2lbdY5iurpsDaXpXLzOdZp5BWjryAYCSpZtEYTTdDeiUdaxjobi8OYubp6+uZN
S15v3HfLEdvecqJK8kFZ/FJiN3oC54uekIMhOej+BJdiTR9SlVP4qjjZzgJe/YKn
rHct60vlK5AyH039hZiyalgasBYHUVUaNq+gLoZ53Bhxa62ogjisRzpKp1fHzhj8
b87w8eRqvtkO1icwEwe8Ow+7B24j9TVw9XllPyiwm0rxe4yOBzz3V2XtLndPzP1R
pQqZLOPT8XomcIgGs6j3/3qDG93w7mlaVKbUIhTQLXpak3cq4xiRSDyoWzVqPB03
lUaUeATtGt3l1817uZmuienSYkWfaNKdPVUdQ+0xN5BVUKJNvHi4INuOy+LdHyDZ
JHWSoawfHPsKPVYMzw1GZN+eZ0/ve2B+XiIlaS/oac+jwjG2PjSfuKv02+OLYcuv
xZ6fKOFpC14B9NYjrNnbUP4viZeYsMlB5gz8Lpg1ogTyzFj9ElJZMCakEDirV1ru
g4lPhVAc6eoqNYTYgt7xwcPIFGeZroAmKCj53ksntJbX6EgGIg5SVFhnuwnB+9h3
vyi2jvM3gp400SNGamKU6snY0UrWQ1HDIK5v8LcAsnZTlLencOo4eVKGoOPZuejq
Tfw4uLDZCJlRYeJg2etkaTGMRwKiXFXbxZrmm9EHihHAPyasrMyia1K37nC+UxN8
wmtxr08YRx0fc4WDj6oOBtnDDFW3zvZtVZu8yPTtxXKVfz87zyOwrQZciWUyWVIB
gDnOflWCsMb3n0gX3ZN0tLeVVof2/GVURPTCwortKl19iuu/srRfMkSK1e3VJUet
gEjpy4aXzXShZVbKaYHcWynlI4I1w2no/TTaSTJT+9Pt7NJwa1iPAm+dqAQ1qIJQ
grVQ0pIg/yRrNj3VchPBAbNz5PsTytYXFEjzjCHz57OcefD+wehdVxYxzEJmXWxP
sDK7ltrHryfp1dzRMxtVl49NoPTqfxBnL6AP7nT4FcgB9QTUOEPy3tCqKmN4hyF4
RcOGcdCg7aF7NvOciuSCMe0i4q9kkovi/3hNwBR1HVWluN2q4WBn1Im8rkByl0IM
m4dKbyy9iqV0SGJwumEs44we8EuBe4Z7LBPCF8MrfOZ73Qu1GqSP/sOdf4OHH4Yt
cmwxwgXh5mUjK/85bVz1+nVsCtODVmtZ3VP8ldSkcWhKkZ/yBSWFkTz21xXNVmA9
tz0nTHI9ENNMomCKD/pg2ZzXjwHLcxw2Gf8kcZVjye924oAhCr9aNT27yfXkaAjc
c59LEbooaoJVc3tcifDyWjQPxiEbGptLMzKtEXv8fHkMAV+jZuTm+eRLahRn6YLP
26pejBt2vZB7AHxWg/QMg71w2mNyn23CdCdMn2rSFMa9A0CixA8sHHWPv18VDMPF
cpZspiVjrfpmoEdo7c0G/oyvNitxNEAquJwxzR9m8Rb/tfvonzkz/X2mkNxHZHpS
9HLuEZRbezmBs5lnRFhx7i80iktoViBDIJIj2Cz9cAkiPgTQEXcWoIgWqGP6cl7X
XtJ3A0A8GYjrgnl88A3orrT6df9n5UhMcqhQY+cxNl2pusFzHNq4zkZzG8qKEHYq
g2ngWWhTQNBRkR/u5pXFUMTPu5A7ZbH9y9yIDaSe/N+fr96zK2pSzvLIRR/kUQUy
aTDMhqrREtuzyTphOoQDstIHfGuwuZTw6kGsUMcYdPFjWkjz93OeXu5wavrDpniI
LdMuWnSyLG6iHDGkluMOxL2+hx0CdNTbzZKRQKwfegcK71GnOureYSvEmzkIHz9c
W72mRoNfkIMb3x5fsnosTPJlFUvvGAgL5LS5nrzlyAFt8DbNw00o3Pfyr4Ng4KHm
4h/f5dhdfGVsgZ5by+9JYXzK2mav4riw/6FZCONPNZJofXDp7eY7KNHkkB+edo7j
TEW4R1bpIP0PkckEbsBD2GilAQZqy/z+nUi3PyhEkYlzkI61IiiyJSNEq8z2SCDg
OJvR9gpHoM9cmC3RIQ/aWUXSMxojovPAM3GPnNl9qLXRuU0vYqylt8sSfpEiIx24
UJBBiKQJoMDwsswFyaLkIsS5liD4CYML2s0du/pr49I4hcZ2f99oxtUnxDAYeRLG
ze6pDQx91oDciC8+yVf36DmCNy2ZbaJjGa1NA8CXttmSP9amaCgwumkFyytQ08QB
lj7W3JJY3w/fFfJvQ+MiJ82FjHwAPYhcOjGOQ/q7MVzNItGr4ysU2OOLSsmxiEkq
DNMb9O5JddEZBdg7S2vACfSPeo11msZckI7clxHiSm11MFJaq+/B22+402ok/eqh
Myerh5hr3vDtFpNdTO7ARaptoBGKlj9PFRCLddb54DdsZyWDtMUMkzWqJjHFNlCE
DNh10TEExfpbjWxf0zQZvAOZLtuHG3Qj39Lk5LcVEytq1pmAeznL4IZnUMxi9aLf
RNJo8N4cSGPHRRXj0lax7qY+NDU6ibnr0YKZ4TDQ7K682zo49T+EthJ5XkcuKjEi
JiGRQx0dwT1qy/7pIqziLdM1YK/chIsLXgGrxmdMdDCBqnESwT6a3nA52wakTe+C
irsbjp4EdO70zNo6Z0wZghdGd33rR1J3c8DwPc2RYsnVLJnyOlpOgWpLw1qw+2DT
q55anWYMIB0RQWOsFKPnopac+NBewqsg8NBQqK97tM7aiNnIqQJKuEvGVhXyLEOS
lyhfBgH+S30B2Q+6weuqKBGgWk2vhuw4C2ibUnNeXRcNlcJzPcEwyk5X+xre8L1w
wZBG3L/CCbDWZg8L0Vs6ZtvuTrrd3svw5ToNFfjHcaTBeK08NoJRWNb6qbqmIrEQ
2fUm5KYhNwq5wcqhmdMc4MaHltqaEV0N+Fi5/ChzWqY/7sdHcilFkbdrxhIVm4HF
p2qaqQT3z4FR3u00JDyhNzNZWYsUFKmgHvl6jSwPtgAuXj70AG3YH4vfJSxAM4Gf
qsDeXULWGkcFp1H33/evhNXxiiogQ2YPnRzMMYqtABMdRd/Ey6lavxkYCIZJwOWC
43PzwL6nXgvs+ttuA6e6ujRBgpX4C6ReR1iut42WlRBVeZuB+PT17L7GBDF8931P
kFgEQaQkuro5c9WKWxia9tgZwamh1vqhjhhmxKdgPM+lL8hm+3hXzKXARMGWwIcq
WowQYqmAE2tekUb23loeTeYtLOblJQOvNeohMyCLeZm/8i3Qa/V5G3nUhD3zEBEb
PpV3WpRGe7Ya5SrBUP6u+yR3qtSjhEfmplrP/8LvHbWacKVIalLqfp6SI7AxzPC0
XHAukzMhneLhArjXUq7+a2Ip+Dm79oLtI+ppyRWHxfCQImokeyqhcFCRKfCuktmS
kFxe51TgxJbodla0sfozoSl/QYhdcRxSval74ZvHHH60ImZh42Lqf1uR741wOY90
UIhsgFaimt0Ga+Bo1dpfp0DLAyeHxszGgHsO0o0P3DDua4KZcti1tNzRGGl3T7Es
qDkNN99EivnTzuEfZUs/GU6bPQBtIVOZo5vQMaG5YJ230LRIjlVTCe85emrCbRQi
YnwAVBlxJ1kOOP9URceK703h8nRA3zgNPFDK+XtqJuTwTekYNQsdsh4FTScvbgQH
V2t2fuwyiBXDG1HPR9YEdj9RmH//H4U5sBnEcCtYbNujX1neTqpjcjVDUxtxWHsG
4nG0anQJNmP3lGE49fiSg1nudUXdRog1Zl7eV2v4qar7BrQ2lZGi6Ant7edFOZ2f
WCYgigysZaYQL6HYLHhydH0zyFIwfGjZsX16dIkVkWkErP7qFUxyCl3wnOmMyIIk
LWH2QR1IaxinLQqLtf3vWJgPeyr11BJv0l5vzdGyOeqJ42JoYbGZOFHHBlHWBx85
1Ri752LzEuIg8s9nS5WxzLH4EUB1ZpvP+3k9VVCCotURldCYFYh8tXuj00X0HTId
aZ8bBUD19KJbhKj9x3f6zrG7nfTjQHqSXyalGXMVCwChd+3QVJgwWt9azcAGrohx
njASw/sCQLtJburM8yDXSxA2uepBhc26GY9AYramwqoAdnVURsRJ8T5JlMD0e1OR
z/7i8ZKI84b7eEVGuvJ7gCBpBtPHunsK6AYqpp7Qt4oRfxiIozg/A4m/+bfrI11A
ZPTbxb1NvAaP0mBwa5ath4EiJ9LsXb1I811cQL41q78uJ+Qttd67ssArbbge2u+Q
JBrvUO1n219/xVJiN/5FLHssK8DaKmHAXsJvPKTPkCd4d2bE4Ex0//gZtwt+Xgpp
yB+MHY5DsChA69apwidmhjKin5O1ZfJ9RtWeAw+3CoL8wR2azGNzwaIb7TZa3a+S
il59bQEXf387n8BNmtdAX+yGt7rgg8rq433dGQqQG++tq2jNIn412nlWJDlZSVm8
YjQs5f06SznGS6vEzm8Syy5O/hJ/i4DiL808o4hwcIyb5yPm9jCUfgm4/8vI3rQ/
cDAeMGm+Ps4aUk9ApOtRB1OBe+ke1/3EpQyWUNOA5k0wA+aMIgzVwJXsWW/YpHEo
xMePEYcjFVx4pwFkp5ZcbfQ55bihonWnvr1tKP3YSlLa+qxoJTeA4Ni7OAPGXhSC
EjUv7Bcwo0ZKD3MDyun8WAa2W7klKLBISXRMSQKaSycIV39vCdb4+DDdGdgChxyv
6+s0/zLlXRZbiPNyotVGZq3HMDSLC0ewYgKJKfxabwdF0/plX3DYdAufLhyx64e7
nXpOnCy+z6DegrrOCM07FKEdK/y2ZR5dVkkoj/WCDB/B1AY6Deg+MTwvtlC8L5nz
ZRRFxCZbAcUuT0+nwpIBQF1ybDFOJUMi5O2XrEqq628bsB1k+GvxQutUN/oUeAEX
FTMQ9J2XTb1klY1wF8/0Y1qNS7rkvPTf9FLY8DaM5E0T8ez4FIskv9WKJoNp2emR
MaZxE7IFZpKJQlO4VTgS5WeQmhxb7BPMzQQZCyf5h22xa09LeWBt5hfRJABu5tbg
J+rEsn3DIs47B15sDHXWpVboBRwC20PWpjrstnb0eK2a49iztYt2fBO34QYQO48y
F2NPAT0wEe1Ny2kV2q6mXnTNpjb4fDriYAe9kq02M4X5B2kW/QX4lL7vrERrJyU7
pKE7W4YoLSTMLSt1PujRdBPrCZG30kH9J9k2tZrLHgeRan1jRaWtROydqBW3XaG9
8bPJQGaulk+5Id5qkGr0+1W01WWOsboIRJyJymnnYUPi8U/0Uxmzm12slkLgHH37
4J3FGWDNkVM0+47ndP/GU6Wq7amN4IyfqErEgCkBgijenheOmy8wFXtOSksigDK3
Dl2fLGMl1BxqXNCfBOJOBOHga/m/embsQ1Q/NRB3bLNdAIKouZZ7CICJaBRF6P1Y
khuI6sXStOnkz3E4fbUgYzW9h86TFoXwg/jAvQYcjDfH6WEp/WK+14STWyx4wS+P
VnLsDp0KaxcdPgNeRFYw4zSJmfUPO3LdmP7OkENjpx4RmP6BaY9mroCx/f57hOti
pzxNl5bDC+colpkezUVhs2nXOiq5j6N6bJNU82KYN+Eidz/8L3nBE4WvJbsxRh9S
5sc70LjiMMyljQ4Bs54PDJ4Xhu4E1c9ZzITnUYs9QelM/zI4FoKD4AzdKT+BEcbi
1pvJWc0ecW1eGmzLa0AGS1ro9VaE4LACHwvHQjDsQ9XlEfKd4Z/jihFAsBdMCV4j
MkwqP43b74n+alKnTwbT+wUBLZ9rMNHT/YMaohqD4HRniEVfOLeyZ6Kq/rQr+MpJ
dwKBfv24OAKnnTW3QkI3y9b1OYPFJ0Nj/W/WtPE7icGl8eFzAaaVbmVTQw6ubDef
/yD/lh9Q/78olSo96QPbrnwZkIkAa2mGUxzw+R9b9vQGO4zE9Q9xWHd+ZU8nK0VV
C+wiG8WyvAfO0CYDyV9q1m1kbYGSZKQvgszLlgNf34v77E3h3fmZrT1JNZGYlRZz
qAYiovdF6jSVil9lhRghmctCmtFfqQgsjGQ2ztCENQ0ZZggmcdfoV5YuO6HHkIs0
6Q+jZc3SdtLORacQQCEpCpD+T8q/uLxd1oihyPviLxFvAPIabHanpiu1H3thxIXH
Djq3YF3zJWTcIi+pC3E9ChAa1iKgnt8JxEOi4yCBtVP3AUX8DfNyMtJkvLK9+Hd9
BE2eUr88aK+guLVtFciFVBP1dvlvNG5WilbiMOlAwvaxgNDuDddfrUz35hpOiNsp
sktd/e+ruazHr5MBJgiaFZKD+XQEiBentYGNOKNamoQd58z3PB+W2Rx1T8n2+tW5
w+HaDRGqhXKcYkRsH7Z1+6PsDz+deTwb6Z2puS6usrh0Ol9SbC6wRmiy5Y4j+OeB
SFE8qlE2i4GwDFJl1JQHOZvaZXId3S9mT55PBxKw7w/fHwmvpi/bAQxJabAbCJGY
ec4BXlDWTaNuljEdHo09Jix4RKmUxlMA1RfTsUuf+eLvKX9SZyaMx0vXZdm863MM
NnZzAYiasC8qHJB1uiz8tlBT18HzEpdlqVlHo85RFhhLOAIdO7IRi9TKIkEJh8s5
wp07z8/hCPBzT/zdxSbWSSKcCEJPkV+4Teu1TbYrmB9ge0KHlj5E84fJNaRiKGDc
bKO9qfvyz8UjgwlRKK/Y6bPjD5n0I1+pEVDHu1d4NnsPLFNdRB8xhpv0LKD0kc2O
M3PFopPoFNaWsZkac6fDKZAEA3wMNOY3za+5OTVNP2BhULEijluK0xBt2sEo98EE
FHzUxgL18l1zlX+YN3eoYjLLCSWVEPDm+uk797UO6fi1tiuVj6WE8rp01/i6cfEu
tfFvzgcKjK/NeegKYwp3GmPjEMtk9dkRgFY47hFBhl3hBsra2kSZWq5YiYMljFXo
ekrEsXq5S10V/mUSwC8+z9gsWn+cRdBM1bSKKeH8MZkiszj9oGror1g9FZ4sejGJ
wd6RF6bGhScWL2WfmbDNPTfe2sMrgwXZXTpgTAZKmOoWPsR6ANcr7tpLRxH2TT4l
pJ5C2NN9xAhGUFKCRelsUmhEgS6fo+YK5t+u/8D/is9ZpaW2CpODW/vXUgZWd3h9
za2cN5uYLTJM/LoCspKXzKuvYXSkloTU8OsnupbnxswrG9quEBjAIeQC77n5Hlcb
6gyu/+05VnJWb+LRpJBgakzFwxT4u47ZEZgL6QRejZmTEvWOOO1kA+u/TTCnmob6
6M6D/1SATx4rWmpeooxB7/9J43Nh0IRi9Hk6bcWdFIMVd7RrflPjBrCwP2DAcyVo
aXbaDyitGwAKrUe0e07DGr1GIqRcFS1XUzx9f8PP3pS5NBcXxYUDs5hycXRlPPUx
hY69shZRMz2FJRX+nMQ5gxEmYldNuU2MxdXnPzUWHRpCg7yHS+XbC9hUSErL/OAC
un2SfoC3KDsx7b6e0v8qw4jbt1Zmoxw8lfXy/evbh5dHXk8UJ3Rp3F0YMLmYtzyP
J2GPSvBE2G3YAhgWOT5WmXrkgibHtEfELolH3MrFRj/mJo894jQ8YVXFVSsWEsPk
B04saYO5NJaOJAeg/1YvFWRADsV45GgzjxFNBPPlR4XtEh5yMdQY/qVt0xFKPc8R
an5q//vYE5n8DU1As9TMaLsAOy5l+mDIdL2fMBKF3pShGs+4tIV2j7jb0QcnVduh
cQKF6XUcCOWvWfM8PWI7gjjXJXoyLG9rmed+PpS4bb/y6MpzwQgKm52mGNKDaVKK
gNSFRrAfJbwvJV2ATOD/kEGNpqMbnQ/bFCzk8DqXJJ+oWQ0BYGL2UqQ8h8RC3LUX
nBlWLfgAMKWqWAwjAKPqKSBYdRvUhmd7MDMJuDl5SV/lshI/HdDDC/YROoBS91W/
06O703Vr/uY+Kecz44Mxer8e7qQ3JkBVCqzkbVSuT2H9gdwU3tVfJ8R9YOjptnMS
nf3mzlkck6A8Xxkb9mjqn7yZfj7+5Ll5C10mpee1Fnd3s6Lr9bD4LHy5yEbOKrMa
d/Dajuo2RDyeo5hgNo/x40e1P09pBw3ZWLHADFgMvzs8fG6K+/ikl8zVSTrRhnrD
J5r6LSCcB/j7ef5cQ3GUepWvAt4+T9CIP99jxSRiGYh1lDLfTEojzHsvRw8r/OsH
RwNAlE8vpu107hqoJwGAtSReciMm40wuvoRCjwH6TAw3AKxX5TNYJBi6ypXH4j3A
ScmGo8f14P2hbhsxEfCoNAY1+WMbHro6QVkIg2FFblQzTibmpR3oIwQrkoZbQY6H
C7Uy1E+0uka7cgeeyKV89pFO0vkklt/EajsoTdZhXbCgMtlAfoEO3hAN2l9RGuN9
NYJh/fKkVdrsbCQSVbEjH+7zE6FSyEirdgcTSD6ASRUFf0prxzxcAOOV6WFGerjq
NYwTM3W3GUCPzf1Pq+JlgKG9sBGu+60kJfLBwe+olaMv7nSsomf4PZpePFa/qGn1
HOQK74iPWFbN+j/gQwRUPKcr+lra7RStwgltmn3Xm6EZ423b1RmUGV1tEXf5ZnJC
CPcBZDczqOk4fj6EYdraoWHicMJFNeLW3g1lgq+RyB5E/Rme39H5rjyVeuS4FCSr
16TtaIvUhgIZkFIKHMRG8zEHP5tC2kvi3y9SEhHmB+yoZivDu8CBZiL19WXVa8iX
u7Y78lEe3zHSZXxpL2F+Pd29yE3C2zSlCs5PTHs1sj+87a6tqiZDDmhlNzpA1+yg
j+P7lXQcjGfSlc8gk1hoki5/9uMHC5jSKDmzvVSVE7lV2kgU/eBB8Or+u6g4SHSY
Ct6EKner8tT5oxwXMTQyDxDtZSs0roWzkDGMi2h2/b555F6rVBZk6DOXreAtAZaw
TqprmhZNNT/Q2OpFjApW73GYSDiJ+TzGhIvOR7uQ2afDBmQcjQ204rg2gthJ+0Lm
PNnHEJQdK9QJ0xJLPAIjm4brLdxYOuNJB3Cei7Pgiqvfbi9NT5bpaU3JxKZC3OYl
1fmt4cmsbB6lsGTPjnfrx+udWjg2zDQ9M2uAvOfLg/CqBoNfHsbqcd8f6UYHlIUl
7ijMCzq6wVW8UoQuG0JsEy7Yiqmtv8V2cSUiKcZG+s4NNhyozs5I+aUMsulJp/rM
W0N6gi6VD2DfWW8JqdKlQseZn1Uo/1+vrAefvdSDZhIBr+dDc9pCsDyuzQq4ldI7
4ASYpfZXxFZyQ/AzxKOgM91c5SVIrdOgm9GCyQ1CFGhplGjkIy4i1AzPrCMLHVWY
3qGLp8NvSf5lHRP1q0RImXezMa1lgtKdsmgYUzFpdgW+iapIX65hRoqrDKci9Grt
cdCvHUk6ECyZZ+R7g3ZuixaY3hMlp4UpkueFyvaIkzHkfvwIq8nq4P6tWFRyaCGf
ETgRdA2tOaHXtzWz2iBGyuy4iD7W01uURWoQUy1KOLfR6qOjDTB9S9NaRI2lsXZB
hlezs2J1y0G2kWo83oNG3Mcfyzh9Z7vJQS5lJD2oOzWHTTBDUwjs7jTZN+4XTwXR
KX50q58sz0xGC5pB+CYbBsbtEN4Kuz1B7f7R3DLxUS26YsMRkX5Kmk/8ZRDlYMAj
UWQYncM6RBmbEPQ0K/lQ/CDE7N/oegkOJxG8h3+lo5Q1uf1LTsAmo6Nu+S9MNMI9
TLHlx1ERM9UIBFb+st4P1o05kBhsvz0AJIscRke87IVUuXI/SawIz/zBjHt6cHm1
xUMZHZ572ffQmexgEcT3Vv/I0QTvD7gdZ5XwYUqb5BqGQYPo5xBXj85pUE5RtTO1
BW2F33VoIiAKksc7X1ReXEeU4L9zAe/q3jOJ4MSRWghupeDeIlnz0b7aHEOi7tYv
X7qesrEwSoYm7Wdvf2weGc4fP3ACtIqegBGj0pq5UN6WZ493WlRcRC8sYxD/JGjy
db4O0ZL11eqy9L+3QvYUvm8e4KxmBIWr+KmYvMETI9MXifd68n8v/Cjga4g31G1C
O2Tufdh9A4y5qQhZzT95eOLDW1L30UXG0Mllk7fI1fdnwQpWCSXq8t3gdgGxgHRL
fAZdLsoSG2JPSVobMVt86/9oEltYWFzHBAKixw1YiHDCWaKcnB0rZsi0Wk2EjDgL
duDxL7mAeI3E52HtNemimRQX+R9xCObynlne44zsbud7fOlRIjEM6WHE5uvha5G1
56041MCz4KJdPN29g8C3AxLsjfHs/8lCwL0PNYfDXoMBQQt67v3IsT8+nTTBDD/q
IjOFP3YYmjC/xDtlLrY9UK2isuNhftqxfjyXtFn9+/4BfGK2+3mNsqJhJFH0iiZT
+WC3Nyb32kVnRP+s6wCHLUKV2I3bYrsx7Ommf9RfKoOMBu9zVCJ0c+Lj77Own4DE
7JUn2wIzfhS4YVwLQfjOs0Wik9GsEG6xS9iejtTcADGE7g89mcRrB8MrozMR4X8i
+OK8YGKy1AHy/WA8WuLQYJxHGx0fhhZuAOVGh6KAmRXQ6pR6a1lTlXW5NHRrz+1x
5KtpkRfPjRbj1hSwMecdGTHfsawwZunvSddnuMtIC6B69khFmr+AX0KEPzPfXR4H
jg2IDDN5FyI3CF5PR6BFv0xLdFKg53A1fUf39aHXBGUcZiL1hAJmfeqQ0E5az3vm
QlRgszyZ0P2EVQXDpIMMP37n7Aay23NEdwyfE4HZKeBqEL0iZ6P0zVtcXQH1T6Tp
9BXTCECiLc0pCtBaixuZx0T+B/xMKnDkjeIwifoYt5jHHljhFot2RFYzI3Yf6paE
mH8mP51Ki3i48q2hWQs9WOtS3sZbuArVn20+xaUxDDG1FKI7Mt4nklMTq6sEDfNQ
moRb7NaWID+eVsU4JUoq1wIhZwm65FWnEmnIJOcl7SNFF8AtOGTlAU5IlpLhWCNd
qCrDzu6L18+iQlfIF7B14mQEBHMHQZwxVLp2FUfijWLOsdHPFC7efJ/1lFdjyusJ
k0a24iAGR4vm5cdSOKQ6sMoqy1/niQqpBGn0fHy2mU3jfY/pSANEd1vOW0U1eSZd
x73i5sEcWOoKnlWwmrc2Jkt2/2HUH5khSruguMYJkpnRtx+xUgI0s0z7MLQaxi1o
DMsebkB1VELISzIkzxgzxLWuVw1iW9+wDg5qscmRDF1mEl+mbjCQDdzTWSriJhS8
z2j5jqyolmj29MLQlZyOIYiYQLdTaWbz5yc1AhcP7dAR2z97ehBmSd/bTHWgV4+C
iwvE0qv6vj+qI0w+WAaX+/qwcpHcU591yCC2mj/rTEZv7MrAJU0bgdVW+McfnJe4
zRIkfo2d6EAaYRZsxndj5cJUsv/7jMjHIh5XJNlpOKw6NzSLDmX+40y0QG2GGIMN
zsVJ8Nwj5yIjP3boS0h02xilRIQLs3bSCWgA5Pr/wQwwuY/b709k7jP1l/aucBsW
E+7r+Y0CnAwmD750qTestqDDFvERHinqXPRmexMO/kLRDaZq3CS07jGIRkrRHte9
BelwrJkH1nEvisgx6yRtJiukYdrEd5loXBoNMwbP7BO3/ebbUDWlF2P6ovWASQ5O
x+3QUy3cHFZVnN5FeK/zOYbELkf+YBnZxsiNBfDxx1tehJd3qJf9/i44NVMl6qmW
hGXWo++4qTezncPDM+6dQgyYLz9Ko0o2nDaAnPP8Fdxz4yq8eESJO7PbuGn7Rm/Z
n8+TinnferiKOFPbUCCWIg4xHVRr1uEfbykk8O/rymSe33f7DheT7R9BDh4Ifq4F
1lgDgq6kaRTye+mQBadFLaRr++EGmWzdiQqjL1o/DiskIFgPMVzC/ePNJwywlez0
6I88uzxF5ZxghDuAkeakziIkxLcjx/G7C6Cg0mtUiv50d1/45QRZ0v9oNQcPfgdA
ERRVhX2JqCJLCQJTSu0VBd6AgTbCO0KoXfQAVJf7ASmYAtbgNI7s6GyKkrD4LGob
6Qom2ag/j5dMRPXCaT/MydA6lBEqxAw3XA4V+Wb2cLdY0b5DVVk+I4wwYSHDyekL
nxDmwKoXqwYEmcm9gBkMR5TgscIDdRi2w04ZWcqj8kj56YI0vNEFaBIt6OIqf4xL
stn/n7BsYiaGqUh0fWyPGsOEZfMMRHLVdW1yH+AhT0itN5wNNxUQAobff8XYuQNG
HUd1+2nUjFXkPUKNALcJAP7XghEg51/0qnlLzrvYLABjhc2TUXTQhVIie6Qem5Ew
Sm00A0mvYgkp5Pel+52wC2sm1inQ14rr7AkqczDEQDYYl5Mfgq80wlS0jbseIdgP
ZmTJNDxfC6y64f9dxVL5OYA3Qpewva8bnzs3BwcmKGKubCBm51C4rwOGXppb7d9S
ljKIDjQDllC5gVpHg7UXMd4VGbZLtOvDjok5r1T0FwL0KdvxJX6jZ130rqMy6rRn
WUuRCpeO9m00sjAFoqIF/LGfkTPXn7ggYZNR8/xvjoV421Biat05xJjabOU2j/Lq
bCUGouOlmaGpDVGDbgpkOmtHzS6sjvIHl/PThAknbjol2vItWuBCuFDV4e/yi0yb
u9TZBjRbk6S7X+Na3iCNiPomNjNz5ItFjRwCKC04bObb5MlEqIqJrITBZlYPV5dm
EEwaA+95MYZYC9dGCRK1WTXPF9j0FmJdTnUDkFQyoVGBEywORrg0icZOinDcuJNb
DCwj+ewYPKg9lpbTmPGAgeg7Bn0DRGdoLW/7sCwicyXGIMTDzPtcML51EqShHHGf
0W9nEdyMSSDQJT7i0J4cnIimMWbQ8qAJB5K9aWhgvRZw2HEiXqpPF6mh+U7+XJ+L
+DeaEMGRrtL37ORikEa9OQ6l6rmDOolRm0PBt19IkhczGpa88lctxOPBinmiQIJg
Rn1KvZpqjjqZAfloZELhR2awsK/FI5qK7eFcOLAvuwDA+QHyXDyS1L5GFUL7AsEv
XbgRT8iYMtLFSWBYu6euyD27yY11kb4rOf34iCInxaSBEWmjNpO2WUBHEut/W1e/
aY7o5H4YKRZ+la9hJ5w7DTJdjBO9TZ+i+d7DuTYSHZaEA+f0IVEybRDwuGk2Iunh
IfAOkrZXk6EU6Tjozc9Cmg4yBfkIvqP4CjyTzmu5pLDWXw8/MhLCU5dcYtowC8Z5
Nyim6sVXIp6rX6OTXns31vVrbwnzeozjmOZ2COpZFrjli6rbyKeprLHraK95vW1y
m0TtNpk8EWAcKdAoafhvtWb5Loj64ZX3czzO3C7S/YNFi06VEohvmyxvMXjvNkqR
4fM5A/5rU7qtpXr4TkG5sOLpPyeK+f2z3lLc5ULArbpOFfhx9lNJA8z+L2VxiKfT
+hY8LIAAzQXyXLP924ySjTSh1sX48mBS/9vaImqcU2axCkYU7mc5d0DuICH/DBau
t4G4LQgz7KjGeXqJuEFhftp0VH5HKrZBRqJap3j7D6BkdBxMKAvbJ5k93/4BEFXE
vbLeJ96E/OTdPVg5Lv+W0WDnUiAjmWJdsvheDM8BBc1s8geGgn2wlOgCIMEf1sfM
gl/zE0PD7d474+x4O7WCjjKLrskXORlkQwUjWztMMC+Wr95K+0p6adRqWIEUhWf/
YQZZFOL9UcyArYcBVm4Wuas2f960nlu7kxA54B1xZ0Zelk4lYUplESeSci6q0Wc+
U7AYERvTHI/8xujsz2RlNHMDNhjPH89DyymK9A57W1dxn0M+weG2rZ88FuRtoQNj
XyhL/jF7Ww/QqmMjk+51T8b4EUdkqKde632NOPAzEpPAulnDKgZyb1u94exV72Us
b7dXz8ivQjHHq+//qlV8aW2Injt0Xk6fctkRYcHqY+uXck7iQNAPdEu6g1rPzpqS
f+XKxVH0NafOGQAr1NiLjDbsekilWCi+HYz+6ob0rAjUqsbFmfKfdFaFH2ztMBJq
ID1tXqffpOMPNBIP7m/qFoLVCfxWX44CX+atLZq+XBJQpHiAJ8iG6jcuJ1+87uRn
8eqOYPiVmTDOFThtXALUzPEKP07LwfPi3Wu+wUO1+lb2QYf2ft26vVUktGMwu6+g
UaLXM0Ypg2p230941FFtl5Uv7GPKWCW4AkF2VpVUTO+oTTK3HD/J8/6aZ5c+llJ2
P9mLHbm1eIx3l7K8x98FAnvg57G7VXDaXeBewgdKVk9UKQzeq5uqi0dMAjYlS4BS
JLAMrmRFtFo1EVfYAai1o8XTIUKl3L3xuOvUrL0o07g+BllmlTQOoEoQsen/VSNM
hbY3kQv6feNmPAae3iPQDsKBgZGyh9bSIBJ5ThVopbgTTK45ymQkItH9ga4dwY9R
3tXsfOz/7pn6T/ViG01VlqsDJDlKL1c/MgJR5FKQSG1+GT2xHTnkuzBOKMPdeto0
2Dr0v49bvsLgCdR15MqYeHt0VQqLzp3lgoCFAIfBp86ZOKhpw9WDI5In0vRitKuo
YXTxVbxpWBDCuSEqByS/1yAQ7EOZ2pfZHFW6D3P1CQ0TkycvJ53l6I+cj5QxBiqN
Oz+DP7UURrkUIg87XdzAIFLok7WjRGy80YcCD27Cu+A/+M9IrQ8zu47HdgG8MXdY
jsQoY4f4cFJrelyztV5Q8SLPMfpLQGi7aZFB5Xsdk9lVJgfw7p/hkxhxWOMqaaAT
Q3njq+7YnjWD/zbhsCziKlDzHGHiejI+9mcbAOe0fH7DesBhVonJp0ppvOauaAjj
NCi/zDVCCaX3aPXKcREL+0AcFzPs1PQx43uPcjZ6IUBf87ldJxZWSjN2qqiSieQX
2EvQjZLueCgiXDVlL8frvLZnPbic59KnxLraz7cPKF+DpbPfVNedej0fyd9DI3X/
hCEknx8FbeVunNzlYBDRHCCB9TYxWxhDktHS5zbmw6cifhGByjQGjR8ZqBPiFU1a
GNKkkPAXAsvWSQj+RbFgMgiLeQzrkeg35uofUuEJpGMFWwIg+LBph5rl5DUQITKC
FeFAsWZKLSyiT7rqg4D0v5EsnUUDxbk1mXOvHOcZ/zoflDW+PGsfzXvxvNDHwDtQ
Y6HbfmR8aQD8klbrn92xD4hoAPkj4Y8hF1r9u2T5xKG0bp+Wdfm5gGJOnsmd6alB
fpMWOuWGUrsoXX6M9LhWRrZ37ydxZ6ed7GgzlmRr9biA1/EFvIxXrKYsHt1qRgVb
T/fu8o8dHONnxVmEeX/3ciUWP03WJ08woD0Mf8TLk4Xyk23nohw8l4+0/dVZUfVg
bs0eE/JXq5bhh0bhalS/m5eLAhBTHmwxsH+/OnM20bLVkcLUVzNiQv58MT3flD2j
EpySDZzRbg09QC3ZM8G9IcBjKjlXudjot2SKE/vgcRp4dJqNa8pd8WB+ujPNY5EX
bQAvBOt5czgHIg3Jq27vg4FTCVf+s6oLH0qsPWrs59+Wkxto2P2U9TMhLQJfEOmU
oGzfLg2A9E2Y2cD60rFVrtOokysxVGbpjk3YZF7gNiH3MnCwbO75kh7aAB1TX+pS
1I4nnMCz1nx/n+sWnIY6EGX3ZSDYfiBfnrLkxJGUoKumCbCIlMOGOiJYXdmbmZhf
vdUbVV9+QpvkrT5GsHklbL3TRKsdXGcMGUgt2iEQjplDfUWxdCNI0YGvhKOAx/Vj
mcfdMXAnXtkoiXKZCN6t5LefUIl/yblk+mGLSLPQTRUDhQrMahit9Mx5FhSiMhm+
TxtVD242u8vIbLwczzr93vBzRrQGyFEz74VVTJzLVG8dh8xNmx2tBEiDOMhytLj0
9bm6D7tLc5NQwBIjZesQoPvdvCWSB4pBfrjW8WFo+TOpiWaCw2foWKrIeqCouJCi
EhXBo40e7FdAcXQOSTp0AFgmDGDg6FvIo3Tp0eTrIFVP9TYE0pzxjZsJixHgeQQ5
lDSJ79EEC0FNJo8Z5ARU56ZNFdT7NWo6eVRGb7XVOmgM7OzU0BP5WBNEPgoZDdk2
Gyf4gW8l8Br8tXbktytIjCwlH1VM08iyZpdegETLCn2XhMsQaUvPIXq/jPOvtgQ9
1YEYPgKdA86pSTFjVIaPdsEpPNyVWXyNO+7m023RRL4qxHR5QCZLwZa6/c7LCrxi
RYIlPgDHGO2u6CTBRwlgBnyJZheRolfqbSGRFUg1kLi6V2SJA+YDoT9Zin/7oQxC
snE4d5b2kQMZUMjk5CI9sswhnpKwCZrNa2dNm+nINBc2YIoGtO8dsBSLhI4KN2n6
2z2ciHYbTf0eNITMv/bwjTuk+GbW27jebua2Nn8NlzbrnoAL3ms/GimktKu+e3S2
So9MQcMAzVXjT8qk58yNkEJmGdZIEAH9CN6MFcbrFdgEvevaPQtCz6/4Q3xSudCD
P3pGMfHV3MzShtLb3tqn2r73si2S4adoaNHE7d/tJenN9zeZpeIGteEWl78SscZm
kjGqgJfxCMV2uDgwe53E2rok6H87e1GzKHuNJNdhVImCJtk5AGVJOnaWMPpLgiX6
ZbZtvDr613wfVUFit02gT6xqyEpkCRalO4t+INzHnZTMpRiFWE6u4jzHzw3O0GpK
xEQHK1OKXMLj3VJEpNPEuyx/YLC3fXVG3DetEdFcMiHVmfD6FnskUo7qbOwjGSn9
yO8l0RpCT0mXZNWqVJeb7aedkzXooT8jcYm3OYoT4D5iav3CaDJBHPBAM3kT1V4K
KZusZy3bh2r+HLY6qB9iW79EN4cHOB3fVMoIwoAiWqjJiFgARKMBS6dlCv5Zr6PY
k5F5UEmvo+Vi7+eeIeXA2I7GVvbuKDH5sBxYbC4bOe9qvdfO67NJ3O9CBbGWVm2H
jxky0x0F+pW725+4P4vQ2QuNiWeuCvGBtjQmbijtmk/fIrIDLYEz/XPVyg5RcYUt
WAWYYYDxbLV1xlY1I3j3CNo0yup0WBMC0fwB28nZU0cV4EN8iFemRa7ZM5pS5FrG
MziSqhls+iTrg4z+HIWjh/zLDwBoyxbpxxTVmGlEQ6r/45vUzxrnZOPv7X3RKxkW
9CL5m2yDZAF1WMUdLCkApodmo9dt5qvWZFHdm76y2aKUqCkC/A5QxVe4Cr7Tvpca
b0Rn3Q/JDMqROk8ZVFlBR8V/xFX+oDCy6BPYCg50oipN2jf7/E3tuQCWSVCm2NMk
oEU20JlZN6I4I1IRWvil5o1EGBDJXGqlYhBmnEZMND6yBZ5IhBSnL9JXjr/HUA3y
mu1UFAJO8RlKwYoo7zaGRBxQ0Tw5F1f4pV3eq0zlM8ugAFjKWCLI/6infJFMbDcE
ZnbLuX6Iqw0PF6pRvHPZ2t/HxRxPUm6gcRCRFwayeYuVqDVFUj8ukSwPguBsm2CE
2jmCHXjbTN/wdM5JDfFqJ2KaO5SCC6FqBuKX1JamiqxmsVajcu/rncuvfJLOGcrA
aUtQiD4gAsL+5+aCLXolgFFzUrYO/igIdsMVMFgc5wXAL+S/dnYleYJqQy9qpnlH
CmxFHBuaNSJeUZxERzhGlDysQhQhyW+nTRf+JjTzW3Z7+WPEN2cTtn7yH0MLGWgA
griXLO0TAFLAoDUY5Ejmn0zy16ok5nUwqp0FdAm54Om85znrmEmf3TY1hean0eER
AwmMlgncGJPAKNltspRZoIbh7BdT2usnpb0AWLQ9ZmmErdcAQfF/DOIbCxIcNbQa
GhjqbZDuLrVHQTzbv3DC9ruj5vUcrG17qcye795WiRjDuN3yjz7XthAovlixMitI
TccsPC3x5Qv3v5LqhkAnaQCgXJX7j+n0qTtRgxAkruaaYw8oRcD10glCcV836mO8
8zW1r9A7vOqdsyreH3KvDHOzBCqOAfTdaVVuTrrVb1pFvAfDtOIvtJZAe9RjQON7
n61+VfaENgbdFnjP0IQvYT+vwZLRPaQYq7aCC14IklMa5lBoPqY4QL+plz8StR6S
e833JstR1B0Npxc52zcZ9eYkGHrZDfhH8OzurmiBYbdpPHS3Z59uLCBxqXnI8Qpk
8Dd0L5v1RWzawaH1YNAFhi1zKiAsyFAoQyIyElWyBLVaXEA2K9Vfa9h8ePw4ZakA
iVT/P/Rlib18Y1IA1w2kWSO6fP8ZGk3MSuT794LOfl/v5sY4Mj8sHo2xM7ezMynR
8eDrigMQC6+cUVRVnGBrciu2us0EofVNiHKYJ9DO1C1d5ufdR5KoRBxueg501zv+
XeoZOoXAqVlNN0p+rr+xz8k+BPZ1nvg8SpH+Qa+hx6cXDWOfSea5uXhEHBrqzGN6
RZ0Vr2ZfW5nokwXHaf8SXTII24tORjsvXC3MEp41tcRDp4FVFK66LUsDSAxH2gsl
HIohoedq04I94424pIwr4tQeSDwCAgp6i0gp9xk1BlUmvEgiF9P+0NLKDW6F71vo
riQIa8wduvEZ5lwrdNnZ7zwmbfSkXH1sjM2tlnzkg0mAWFbpJ+wcAEM5A8gGWdwU
a6HIpl/ZwtGJw2BnunyKehz1Rh3o5sIXM/HVlzTLCKMYnHgzGkRO52sJMZ83ARQO
XMubEixG9/0N0CZ55OfzbVPjKE3514fEDKzV89NqyK4AokQRoYjF8nAZyR/nIfoE
DhvLapgzhSeGOXDCNqRQfDGFYO6uwpzLd2ApKnJxppAljK+q/YkZkwNCIOYIuZ88
zpCFnOgZSjUWDjX8Zx2iQauVWGfE4J77YGKEFGmxFGUqxfNVEEfB5ysuLWYdNUAY
7uxGxNLr0KPi+nXsfe9uxNYlEj/RQFQ2FZ2ARPTu60dZDN70FnWc7wTbbkGv9shq
4H5kLJ/TBIjNCKW65GcA71dH0QgYvpVIrFYIRNsKkP0eM+dmepDxMvHtMmpK1Urr
syEp2kIAih6VrmOcFGsFz2K/oo0yHAs/8+epeySF5HBNj+zGwNkdd/Ax4VdH4xnY
QygSv6dgT+p2r+s/q+641qf5AaUvf/Lbb1rxRxLGdWe0IFqsxcOfLtntPM+xlbSG
597USzi8UNxutgZmbW5IB5sKdkQzox2f4r0QfbGLIdqRiElI6eFZm64JiMAuBtHw
E+MXKmB4cF8OByev9Sk7LqS4Z0YmSr+JqB+hZpqYgSfKMSdhOpppj0ud3pkOmLs+
g/Ag9zDGauNjvOGew7wn/P5xN+vhj5B/6vU/gMK7YES6ihZvD4m/agizKQJR1PNA
nKI9f27PWEMu9Ov2CT9LMPP0xkQsYiwhsYsxwFpWnOKAYYG0fZ+QGwTpfllXUUbv
jPEUjrhEKFLN3jGVHj9dgGcDM1ckhUimRSNZH/SFRBdvsrE/VvjtVm9unJBMQbKC
ekdCiv6kWuH5UzViVy7f7GWNer85KQtajnDYqODOLfhIwsUxrVZH8VSOTwjdHoZq
1MtUtkfecx81lDw+zO6fHBJji71/07hgkHu/9kP6nxnhFBUQV3as/4EhVGno4mL7
1dOFlHE7CA1fnBys0EIqHYIzUPptYv3bbyKB0dg0a4rSQD7GMQUEEWsAstQQ4Lfm
1PTnniQS1GCxj8jL4KJ2/CJN36VGtImdtzFzMoDHbsVjWLOvBgg442hMr04Ieyqr
RoqIEE6XlcheZrNL9O+XUhbHgDqsYpKqc8plrsf4w3slXB0ZWuGDyTZ3z/HJWQ3p
LZCojIIV5+LsKJvCY/+pJvDq1NeuXeBXBzDnguhaps+8XoblM8PcwoQ4enzAJNyF
eru5u2OaEv2FTnAhpZoLlyR3Ew0boGX9PygssipkIclvdWN+0js7ePrqlX0ZOiXl
KSv1midwwotRuIZmuQ40+Mats0CAmtbyFY06fA5kgTreIJuFpV8zspS1tdibm78z
ruhzm3ZUrYs+6et7HGDY2s91nRXTd1G4Tm5Wwq7to1nN8mx39ccJDfkLybHIEwGP
bFF+8b2yO0patbbQ0enMAQPYDWtzX6YA13nbN2j4qvtY+bJ04s8i4xlbfPgTDqbN
goSdzJQOP+QVDLATFzzwirr1buydLJN3xX+DUq4NPMjpYRW7xXAPp6JgKSxcyKXb
5zOMBTwsef4JV38nRVscGMtSwntpS66Xxfo1M7DkJS9qp/tvEDmfDvCKR5+Swj3n
dHiKmi4eZosQmT90hbPvWnWVVaG76foOYu/ZSxpv04qEqjJRKwEbleR2tfRr4ppe
8tXrowYsvR0lbx3HgRkUnOg2FKQzaNj3EBLbDOF0nF1ljo+yELAt6FxwbYVCq05W
fRFvZn1ao8f50rcYpA3ea/EBARVEmFJBLJXMGbD3IAxRkynGjGreu/0tpJWdhD9j
V1KED5I2F7lQw3qEAtkLBZrWO88tX8vvLVMIFJR8ug4OxppqQ10G7h5QnsQ3CZEd
0PvU4pBKghAnrbsaTIP+AWp1SCKVNcNM5uBMS5QXkxbwjq+MnQJyKXzR9bdiOvet
uvuwCzh6QBfzIXGPVXlKmAo389qTZBhd+hCtH15FYhHnx1yeUpvQreAtVuU1p2Rb
RLhtjGG4d2Rg1CafP5XP4TrSAKWmOvFyr0BRUNSROnMw5+vdUsbpl/7MOOB0iTFT
d2d72UXO9YTR2QOisDW0bh4s8i9oYst1fnkD3GESppNLlO9ecQSFMXg9chvvlyGI
yxG8Oj6jzdOibPmbjqVLBEX3QU30zswzkw+EzSMmHqX9kYDghOG1SMLUHsTTW+Xg
nJff0MAXh3GVgXWjQGmZSxbWX1wVZgsQ0z6tvhnWWb+2IhPncvNfsoKDdzOmEZHO
/pEtLVxLa2wWGUoZFQYKTlSv5tPFE2V1SeANSAqCX5cftsIE7iJ0nlIEhmQ56BeC
sZPinfcrWf//Xzixv2tyKo8j1vzuI+IzSyVNiQ4Q7hq4yd1sWPvZ5yo2i6T8wM7Z
i5zv3JJNl3qUFhDyAUoN/jg9GzNPyeD7HjLnrOMEXDVyR8ao5SZKEkmpZzS4pWK3
18Ik1q/ZA6Ls27J2Qgn08IUoXe4li9xC8nWhQdn6eKSCaGvZdh4iqfb+oyEzyor+
HRQzFLyyOv6s++xzXW303p0KJGi+9Yb0Ul6DQOpqM73yv9B23qImbsewCKQqxQrV
CKi6SzwndKQcQY5mkBm5P3iNUEB4VDO4JvfzEN7/9O9nkTLh/cWfqfkEpKl/FRbv
mNCTB+Tqkpo4aJfJwAgtBg7t3g0BVNFEVX0mhgBZqqY6FgyG6cdx5HihGONgWW64
UXvvbx8AdUAvDdBEeid3IbrwEpDJhoEBmQAdNvfrkUDOxYB8Y97+TgwsHKoJUzEA
o6fnjrNKhwbS9pA5cIY81nKrSgrbBkhv6PXdtLNXM85PmhP4u2f8u6i1pZSJJ3D2
Olo9TMWIWz9pUvOIDAR94j/T4nyi6Uu520FHjGVfcgU4AgkqJONM+g2jiXzHzoD/
wBpbA+xlC2XRmTPP1PZdeEQSDYpO+l2u3fYvBoGKDquXmU9VV+RV+RfhB0JZT5ZW
0tRsl+9gm6hO+Gy7hGmHGVojPQKKHkQ0XapjSB8J6GrvEw+F2M6z9xrw8DLb61DC
LKlEddblqHa5rzjExhSbxv1djehz3WTwocTXlGhps2DlIw6JDNkcd6iodaIN1cxx
YGr4eYzfen3vPFzYm/SNJ6VFfi+DZUReNV5ePnt0w5OsyID1sJUGWQN98/JpaIim
WG6jF2yCcE15YOCwoOxZRF0uAuty2vcwwxawRf2UZqeKjVMRtvhbWpeCvKrzEE6+
FBaq2IvDtccZhP4tf9QCE3u6m/hqHoab9/cqGQFtxomZgxT+VR7AKnP7jlJZFCxe
jCkKtl+E6ATPrnrw2yvKU93mGA1kkM9fODmoM27PT/HDBDrjHrWtrMbzxiZlI51z
lyxNv8aplXUGNmgpGbUhsuEh9fQVtfzTihivjDHv7/3F9etdqcuOOMMCdLjqv7vL
c3tXPrQGX/GqQwmfav1pBh7KklT0VnBcV6yZ89xmoUSbKjfjkEdA/ffaEz1JpGj5
q/N0iFMigm229WHVkvlkroyD8mp8DHZPi757BSRtYDMewmtOGpPagVWFIQUXPZ7K
2UFnrOYzmUXw3fFTzKNHr6Ph7BwmT42/W3lfWoRHzyg1yvdlAG4MwZCRaTN0iNZi
KU/kYhXLYkmgcP5zCu6iZiJCq03LbtOt+XFAxs65pxr7xwvngVDN3T/j/ugONmBA
YlzPJ5f3hDjH2lH6qcobi/cC2PoykkBvBLLk2gF6NBHN+Kkl7QFtR5yzPSWh4UKN
9KfshZsA9S0MKxsToYXvsQFffg8O4ykek2rcw0E7PwtsLof7kmqeDRH6vNgkJTKS
kxnt+X2GiXQDE/6UZMiGOysarGHBV63lVnt9HRZdNVuMvDJnh+Im5Z7Lpuek3sqm
QK0ifI8YgZyOy4SWdBoa86eWxxDYuvejZ1uxLDaUYbDoK7mspbqurgTCHpdAFkcw
xrOIBYCeCMvHEgyYN/t4Czg/gOzR6nM2hISylyRLqBxuFGlGJF0ce/xMxiq7nJZ2
Fkg2IocxQt/mcNi3aXLVdWzPxxGLmx7CZPQcW1uV2NRjKjp7fuLjuN9PIVJxGj5/
GPEavNc6/+tuOT4QEwBxo3sOUfsFMM6JlHtP5vWruzGZnIV9vUsbJKYH4/vijdnL
lwk+np8A+aGZp2o5YFwwfJgfxvwrj22Nh3GhKlRY4QhpruBb2ac/1/siBoNxR+Oe
Gez0B58uyWMInzvkOYBZScbGwHfm7gPAPTDinPZmxOSuW9qXO8wtGit3gH9klO32
4pep8nZMQzZ+O9NlhChZdj//DxiEFJ/IOEaazb0cIrqss2cZ1fLVbEmqFUGnEgr6
VcjaBAifsYodxMKfzcfp1qQi3ZMSbqotFErf5z824qtF4NVYst3Wkmr4PrtkjhOx
KUCRrgsVsIfjazsKvEjMWs6GBvkvKfpPTAGm/Xv4lYBotqsFBaCwErrCZ1tBnajw
M1KIhz5QIeVobCrsv6zrNrp0XwK5stKdEMy8r7mDH9yglV+PY9PZz/led4k+tCIa
8BAg5k2P5FoqdDWU6ZldZ41L3TYupFOLR/2iUZqwv7mk1yI8XmfuM+Fa5RJO96UD
ava/GJjDSPVH/t292GMhOYpdEQq2zOjnKbNXlxMgHfQxNLT4ptnsAlA8S3kHHdxS
yWZQrH1egI5fS2qj8Y43a/nznh8u2XvEwNISB2h0yaUrcoyMJVsjP4EMriNT4o4Y
Tr3vfjxHqWNoHIjRwcvScEOFYkZVYhMIdMFpqMQ5atHrnk0ovwc+UaWv3+3M8zVP
dA7vjAgRD71pFiaQql58ZUyGl+S3fzy0bPkWymscX7yvex4Mx4vBPb+rUALDcel8
HwWdfRFDtCYlnj9a4WbZL6tsCaEZPDMBQO6LKQPAKTGqBdOnI/CHYcQfsBAqwqzR
sVGeO7DcxMtXqiK1uKqI87H9y2opT0p/cZW4bRFie4AFfaRcn3X6qV8dGurGLz9Y
o5dVB+CLKuYH87+tfYnK1+Jw5ei3jarO2u51dWWXncZo3fuxEXT3KGz9RzPlp5iF
KTAmBtX3kHMSQUFkqcDSIYAB1BezQLeB9nwrowSOX8v//bMSluouzLbJdVgzWbj6
p9oxH4SskVa53S0hrDbVYG0JPU3olLbQzl7x1pYEQQCuDxrIbt9jE4v903JruiOz
ZvCUgLDf2/3vnVFiayFEghNMP1L8kVFHal+CEmGlxCGQcN/PWemXUFAvY+U14Ym+
7qaO3eYY7AdcJsrCvcfo4+00ELU9uGqPOHOnkEXcMMuhVqUU/xN70Du6NsOYF/l6
b/nkClIj2ABFKUyXw4AIwK7uP0hEge6wJf5k2isYWHoXSitdyq6FmLdhFJfOs9Rm
c9u0oWeZRoF5LrA4zFu0h7UlMvb0YVL/3Tr3U4sjAneENhMQhdDzSpB16YyQFJ0P
wgusoPbMg7LaBeqnHNSSn5kMNNXuYMnPaiUQ6iH0k5bAjuS1TT5jEonTuXOym2zc
2IOtdXoaO3YG8NI5yzmC4uvCJ/XVbK4QNmXdKlEYjJqwmTMNhoEOohCtNZs7UonH
l6gMkVX8aVs5MKBrMyG52hPWxErxvx0+yV3+9wioaHX8DfYzymWRnpkjuv3VuVZC
GnCkPo3nXgUdrvU3gi0aQXQMBZ4bGaVdcRQrRR+m6BCo7LHdNCDNY+ASHNgqeFY0
uyXoursiqJQWb+93SOJXKVxrLlC0tpTOnUrqF9luZG2jhwUcg9rKyZiuV6gesOCO
lDhbo6ovB93UIT3c5LyEojZrGtqTqzq2f0gpQke81pa0GYZmYloVhbmwUnmlNAtj
bJ7W1dM/MTLKHbJwTuu1znzDn/rYWTHNULiTV15so/LSXnfFzMWST+dDzv9gKJEX
5OPBd1jd4+ccmTa7sG+/iOWpyqh4ya9/e6sRYWH7NAFo/CPaaNeCSXrX2AspLLoq
XXeufXOkbzhgN2wyvXU5x3163juO7iy5TY0zwPXAYwBgcnrJtnj7+Cyohvf2W0fD
0fyyckLOGnHcBl4SytbTQ08DNZk2RNS8AV6uOW/TlTGEx1KvBIpMRrPpdJfLr26w
KDYf79XLYyNr0co0wlEsrGHa3pkuw4nfcv3mqXEQeJEAbBIUe3/p8zWJzlVTwXa/
Zr+cAR3enD7plFSRd3IaaoINdjSKr0bVIniABxUFYsrrmMDHJGvs9vABDtSp68tY
1ZR16lcwstG0Hovlze5pwi4n8hNYZhZRgfxWALjabXvYiE15o4p8/5EWUtHKWyBJ
BOjet+DxaR+Sh2/4xTuN+T22H7Wc6u/W3FSK70ddgPHF8OtS13aMR4JMaEPYSAkh
0ccnT2KWhz4AwLFYPM0pGaP5UDwiBUaYNeUzrChaHEh8sR+g3Yumg8USt/hKaGbi
Dof4MvWEYIUgs30tf1K2ENrXi9IeLUdX4vY0f0bqTuMHFEAMnfkjKhrVTywCF75T
qFa4p5d7VJ0Rq3Q2pCBGLmA7rD8CqDpaKTvQtF6sol9fkvY/0UyyhQjALd3O9o3T
2MKxAsgtwolIz0juhQEalnSaeCfBjpa49w5lOcGxiPYGNYiD+IARsuAozlLACbHd
m2msUEEB4Enzf3kYanI5jtJY9gMDVHdZag2LX/xJHr8624VoMGrOnBALhZYVIIea
QmzqC4wL4VE4cyXqaVwHSLgDczPrKc5a2ew4aBsJv32BROqT88ESSMYPU8iSuH/z
ayqat8hOOirMsbkG8mPTSJFobqP9JVn8i5ZTwA+qDqS5GMclQyIVVNgavoKrbeP2
SasS3b9myyJabs7KpeY6HHBcdcMWxE/zk5xcA3dLGUhmf4eApWIln4gsy1qMIS6+
UAd2c9E7qzOFoe+Mc4kuFJN0r5b9S7JyWhRx5TDfuklM1Z5KIAnVdawPmYpsL5TI
xwc2TpBsKphbo5ss2X/T2pKwofohIWoWvtbJNBR+k4NQYxQ+N9Kq1WZVEBHvbrCo
F26XN6gnvhIk9YtcJgGlOr/owOA8XrgXPKVaaan1YaZtTc+Z6YiNfG4bdFYs9q3o
mwP3h/RXZ32OynrnPB1D+/w69A4K1WYqmHg8YtLvOMkHZ+2v7uuaDF0Qt5ZeJ7H1
4OixxOF83fpiK/JliaZPLwc+LJAUAAYtwuyY5FcVsxN9+Og6N0bKZah+ScBYrUYT
79w95kFCRyW/JXQm+fLtmw9xs2e7ZxsIyeAoh5mSn/tTBzPbuAL2DWIBe/2YV5qx
UOCjhUZNAhOw1BeOMfTMuxXg+lAmNyTqH+bftWaEFgJvQDajyU8Ae+c2JEAhrjhZ
/D5aJIqlOlku2LqJnhzaI1oCNni8U/MZm2RNn3f4rToJYuJAWtWCTweQVbIBDc6D
goB67lWnr96mZZ89J3AK6HlNIjHFYJVV9ucPnLCT9ajVGLVtgJIm4yD50NcXn3K8
pm70Te8awWXApnQE3Ek3K1jsftEcgE1b/YekSzDlVZAFWlyaoMjOYdQZjkoVvEOQ
sAUel6CAJD9aGZEbYz+1CoWsjNEq/D+uoI5oWH427pQ0AnKr7CVhavKYVltV/5EV
ZkOBOOg5kpzItxkA3TUJZCIIa+zoi80NfO6ZvyAGOvpXpm6aGpRNIJukzhqhPmHZ
3YcyJqdgoSFYKRwvRLFcqVuhArvDJCMgrY4/3i7MaOKDSUgVrjJ6WjSOiivbE/kX
z0lloGm6aFeJuZZFFBUp+oKDJbu75NShoIG78vDZCYPl6FDA0F74kaQxBNm8Ou8I
u+tgjy5xVK6Glnz+nsx9pkEm8crRKeTLP5toX+MjZ74XPHPIvT0ztCdSiou/lQnv
ywTWDxdoSm4hFBVSVAHXYWylU43Ya9meEx+urNlM7scKti1o58GzOgllBnEuXyMe
jSr0CRR4Ld87z8CkE+B0QLed9MQHTRnss2BN+GJ2VrmquVRQvEQteM2inICrjMyx
bXL3oGTx3IP59xhYQVXkwA8FoAzCJFu1S7OvBeBAJizRmKSckVNx8bjEJx8ODf94
0QfP/2NqaatIPbWJyL2BYvBaPP8ubElc9mj46fF1jTVbXbttq7pb6LBVWTWv5XNK
IHrvd07P3cuQVl54R/5OMQUbm6AU4VSsFLF7yK08ZnXkqDkxIfnAIiVVMZukmDXM
3hpTeQx8Sk8iHBoXeVEuZlB6e2twJ/vPmG3aLGGUp+qK/NcxtyErbQxQySo4/GCh
H8eS/E0tXZcAO0Ia2oRSFS6Ko9P/P0SPNJtg2nw3nwoZOUR5dqDgmlsqUQ/8hA0A
n4ny5Mlr8I23GmCZ2tyjMK9kMT/l5krxzb157RYtF2EnQvhSAckS00wGx0H34y0j
ioky3sbYQpTo26AKaRWLuodIZZobZGTZYeHEQ15T5Q7/9Vrtx7hc7Sn8dG2T4qSY
vYf9e61PedjXoyYypEPZpIr9CxNjmHOMjaWWVXC71qLlgxe7t/ulw1mqqi8+DLwZ
17nNCqH1hvjMDvBeiLLlxWYWNmbKw6u/XBoRhkO1VKOAM13ZeRXRPlROGxNfyFPz
Jp6kkOvpFrG0jLZAafFAQNi9oNjU2ojPPPN+hdhMvCLo7KXyolu8OlHmIZ7+kH+8
uHIW1WEKZ+8T/Y/fGXU0Xhn693ks4zh9vv3ovTzdz13B+n/IifMs2MSGZDu0X2xs
Q6FNoOZJRMS28zAT0LhEUfszbilLTpMDHCB2tzXwFIorTLiSBEmes2i+2AiF9AjD
A+uGvGnx6v23o9BSFyyDWle+HSMCaEq/sEG8w9eERKLecp79FTVf+bJ/ALp6+yzh
Jx1yael8IwttH5ciuqkrtuzPgqMT+ixJtOexUb/KRs6MuBFlwD9u3mTiTxp7oqwR
quUFRNXj7I+XC7ffDbcLPMSvs4UfO+D8PCmBw8W8ukcG5r8RwRL9sTOWz5rtF+pH
SR787AryqgNnI2mjYtfM2+igNsoBMwt3/bQ/f1IAoXDL6Stn84nTc11kNTQ2Oodf
31QloPG0fhNp2d0W2zqQWmft67EZvqJjx3MkH4Wg/NsdvrojnoYHzyr+q6Yf/vy+
7iuw+OnKhruQ286KG3KHYZnJkbUl1MEbvxkcJncvyZuBfglPk29EYfkr7Ln123dr
MbG+hZjLMFnXFd1Ag/xf7jew/AiMptYRzfua2D0IcipweIRgKByidQyiUkyrmOPL
Dw6ezqh99Ssu8X3+ZGTuFH0nKsOxGvG+J9BZnxaPpPmKIpU+d3JqHgV2q43gs4Ht
j/N60nZblShAVJAyi4+cvhSTiUSW/eKF+5Efdqu2XcPul65wBkoiH4iVKjdom77p
WRCt3xoguqjCAsyjie+d02Xvez+v6UzTiQH/oqRPyfLZ2jelL5j7inSBpmmdRyHZ
L/0C0FRpBvMm7oHL22kq3dwhKTqxQCnyue/uj033eN+ITHrKZfkGhBDNByT4T56Y
UckkM0NPY6IYc4+knp17lOm3wY3K6NOaMCVwk11eWBnvT0rPq5JGWxuJ5ZL6+OGz
TUCsp7PtVKjUbql0qjd12DV+p37cdA7ijmoEtfT62vz9u8qaWR128IV7cblU0lqK
0VeSQYdT0mz9iwXG40DTMVsKZfCoBNnWzM179TTd1oemzHtk4F1Chgnxw3+9j3Tj
0lNgn658EtJcWQr3XbSkXgD/7xi8g4QMCC+Q1zqc0vqJakTr5PDRR8ZHc6ikI0O7
GNqGKThaeiWp/i8Vobk/HGXWmkTHP/m721GnUcQ8GhRPoEi5Y1RIh3s/L9Ff4LaL
UpOZxKwzAsWwiMqf4ajfrCsH1xwB7AenfTZdB9VkEHeMX1B9W35ZuxYpN1+gNlJu
UnjZFp4i8Kl68cz0QjCy831iOxyaTn45qQsFcYlzCru9Llqs/q5C+oXCfGOtl4qE
lo2J7xSSeywZBJGkbHTtsbQnJ8AtliwQH1ijxIObC9wiHaDZqYPLLX3bifa49agh
DyWGUM63pH1x6OvHxXrUbAq8FQtjsZkK1Xcp/yT55prxA4SCpLYDLH+UPQI4YqLw
/IRvsx/u+VhpENMc/u+6E7DwqYt/LqrYyM5wtnEBoSmN2tq1Na0VBmtqDbSVauK1
yIOJ0YpEvdERbGBGoCX9Ua3IbS0SxB1q+z8BMumYdqvWQfwfCpQhEI07z9Vechlp
QNLyPNkc0I+pt1VgvZdt1c1YBhjdblNFmFWMmY1PdrzaLTbwJIFNQDwdyjXVjy37
uYACkTj4b/spIV19kXee397KO1Pgdm24Hji7Y49TRIC7UzNdulrge343Z8DtIamC
xa0vjQCLOKImuaS7w9k0c0NE+nEkCaJi2Hfnh3day41cy/aAYw9eovkE3C4TEM50
z6S1DM14iZpHrp/RbgAz4kw+Qxpdv/HScVPJbtuORDPQ3462FPNMxiI9t+526dKs
cxnJ4brCk8BTuEqypl55TudBInSAwshVy67cbFr6uhDByOOgHlCaGmnX+fKzJbNr
ZE3GMHuzFOmgKoxAJwvsDMRAWKPIu8LUovHWoyirF51pAjVv2W6V2i9eNjKZDkS3
9fiCEVP3eHZTNhPcRhq3DAXSWV0Cm5qunj9IKjGSAU28X4QUcr2TuTOAeR+fnBVa
o9ZCpJuI+tF9LVgWhZsmpB0x8DzcXIxqC1pRO3GrfC0jZXMx1c/4mFsHxVijWRZp
hE18a9hM7aIaqUKdJOWNVY2+tddAno0tO3wjEZnafvATNy3hOOmX1OCBTWLYpLfp
ZmgVy2XiwBGG/m1dQicxHoqrjFCcHpqPlkms8FUz4pM3tWeTpZ0Pj/KGGmLGYIWw
ihEQl9kx12DkAG5grYKop+cEVzRbs3cwEpzSQUO+g0zE9B4hwbfpoJ07fSsp8eMq
Kz+DGQtmihfaPMNCWq/WpC9KAQNBW+dW7v9B8zrPCN8KEdR8PFGNR2IMGjI/Rmus
GDxO+hA8Y0/zYQVPNNbxS2SWtC5Ep/W/lEFBiW1oJPBwfcB1qkX2+LJZduXJBlt+
mrjM71SBLxQRzp5W3iRsoJ1kR1T11jMxyq28G4XdcG57tv4vJif07qSFMjwGrQxF
ExBvWGH91O2XpBeB8IyEKZApOPX/J9sOAi809Lq6iecrnOQwH/xxnghumt9ELxtl
exiN/d+LcOGPBzZFckLrA08WFM8I47cuOGP9gCjIZjt677TCt7TSDRGgET+UEztk
+BddAWaWIAIW6lTjadkBN+bb1Lykm9rUTaklVs3qRV3lXDWURSBJ4tbwb2iaq2Gq
vGaeyhflA1SAI0oFiydxUaSZGFhCNUm5Y5tk/AOewtyU7rvDo763+xDYatXcxM/g
r3kggJQoi6rmW3xNJB7Nvn3RiFQcZqct+nAZTb+YPjFgK4b57sE6c/cyIjj2+boS
XaJuJ+I9Ktmlo/64kXrl6lwcs6O67f4ajylO5oCL+8AINDgFMmiBS6GTW/1rBbtq
YmR1kyt+Uhz+Qpq0k4EUim3q3ip3DN4rkUgv32zwejHwLh1lbLdxLtEYZB892BY5
dM+GVExXCo4bUMcr57xXlYGUecgEBG12oRp3dEHW0xJMZQCBvXXDSX6QW/rPC1c7
4H6xWUPJQZq3LNmeeWtuTrHK9VRFOE+LeghOKs3jR50V68n/SFc/rw9nM6vgJKII
iHSt5Y5DmNSnHFpkvag3vHYYpAAkyA/MS2USBsxZZ90JKs2dWxIiIuI1YA1quZIn
KJSD5Q/y8t1M3XyP9sBXBo6szxptaJE7Iz6/KV7xRtY/1XCyMvieCgnba6yOIrl2
xasgm28T3HyTEolgECzsqMH0IHpYgxtlwUY2Tmsp0p9VuxH953fY3NlaWoWlZcCe
ltM0cOpage5cbnXNMzopcDSN/DISLe0hcYNuCztDKgo0QH/NdmkALzc9kYPOlS92
ua9nd+MPS7wfaGnjwtNDA2Iog5/HU4ZkNAlcUpn6DD9bVFwBNT7b5CwmC9Ha74rY
OqVF8hsYQ1qgorA/z/86ktNSLPQ/9/O0KM5GINXzvfoPhmpfpaGMJoWXBBR6dUxx
DlFMNH38jmmZGgtmKSVfQs737mp6UlqhGcVtnlZ9jgJdwwbwEg8goe93idxMTiZy
dz9EmwOrjldhiwC+vjq1sF4fr81h5I+z9lBq9FnSd3QOmIZWnuDuR0SMuJBcSK1W
qnu6zvSvX+1DEp7vAF05qDfLtTRJAePn8SqK06eMeEUpgCM5lJWacMIoxe8cgCl1
Z1o2wDrxBAA48T81+hDd+2uCB6nNnmWx43CoM1RzUnrG4gqW1N5OAjdXP63cMgac
TOTq1W0IUSTQw8BfCUsMpfjZLkOWHgeydYVypfcen0Phw70lLiZEsfkMffhWxCLy
NA9cM1Aj2C2i5mb3grVzhskNtegPInVcLylUR49L+sIUR8hg/AyCpkk2ZOn2pTSC
riFgHEbShwSateMwsdhuXvbQavQ5YMGhdTkDJLD+yg+M0jMjsXUmFxSO7ASFVRMf
7sq4SjqamdeF3M+mwf399NjJ2K1IZ/JkNPRBCYMoz2RPwVKIfjjq08pX8M9qaTtE
qQMD6AvcZzbGXynAqq8fyUHRo0u2z85OBHSMmUju2JKPhadoR3LQzkPO/qi5A1Bc
HUYXcC7je8gmKFAixqxEMBHXRn6IILRqn+nDBO4u+iYoRh8WLZJYMqRo/z8Tkyju
QJGvvWyYL7pZzhdgzzLrHXWXklPsVStuJmnVevEcULJbuSBktE6wHB6ihKZFdSSU
6tSFkRzXLL7x2n1fcQt1IzOWSoluFbwtoh+gHJIa731nXXXZYqKiEixMYXbg3Yvv
x1WAHD+tFyAUAu73X8A9CUMEd+3PiZNbK4f6JeRn0wecgXMF0cAJG9vRuOxYxIEV
6oh4J44QjkynvxbHvSQxv9EzG4BT2O/zk2LwkR39iKtl2iIfICi1TO15xsFdENRA
d7kljAMUKwQqwmjbm5+QBwAXgrQoLf4uHq7Apx3wrsvmIhzAz9bbU1H86iwJRmS7
Kd7ecbxRMx7JpBHHTwKNmigIuW22h/vKBiR+eAn4f3dlmzlE1URRsfsDQp0czl8e
14OZx3a9sE7X4oR57KWURPYsca5G7XDJJa++MVMf0eh2vn1l+UK+/EiUYBT90zIk
Atq3bh0E0OrywyR50D5cbyb3Z7uCrSW2LFDv5VlraAFu7k89H7dFCx7LK+EJoJnM
aW6smu9OuD/0AaCfeVaudaS3qxYWgh0MXEaT0xHA6emn1cslidEqe3TxYNn4/x+5
94ej4gtvbwxpSapqB6Lp+49/Rjlab/o280kXwk1IbhGNTK1aMZaGlEWNyMydULnS
z72yjCzNWqfkBbcW3hTbO339xCiHiYEwX+4JVVPrEK3ov4+q0p1SnSkmHzncjhdW
8vW89a+vY3J7qRkWM/RuUu4wKTNZV85mw/kz4ZO0p6kqFTgK/JbUoHdXz/q7aNni
DWKpF+EoRFBMoTv0GSKu2oTMA7egcQUoLC6Ux4T+d0O5yOQDfo1beSnJZ+nrdvov
3TSa1w418Tp76JHiJJlLHzd1W+vLGjl2/pLjkCWZAfW1ySxgxyl7DRJw01ytMBQd
M22UZyL61+tDJsZqImWsb4ZwQKjt6Zqo9ECuOoxquVI6zjCL4I5hddXWdsVi+Aaj
lqNEo91EvM9UHUTTCavrLBWl4pmYr/IR7nB/iYxSx3nlkS/ZAn7SOiDbVmEwAaPJ
ul8LeSarpuImdrnB9X0iNiFgbn23mOp5VQgrszPtH7Hw4/8/vEzD20Duvx+tmvbb
i0vsE++w3qrdBycU/uy7IhUjNuEXotcv4FJZiW15SW/+lMyDZZ5x+lgTc9pzihJY
c3f2fYrk0iJayBxT98cBU3KVJow/51XzYaChM3KyQUdBa7xcaOnuHfK05Bg6pa1m
blB/g4Qhv4fXZCCDius/nQp1um5tKSzbQjRllVrVK8m63cNEcDl9hf48JxQK0BJU
HkktxdCRYP1cI/N/DUgLwrHELkW+DsVFhC6gXN1jB+ISF5unAIkTK82zX2pZqpia
POx05TgKNROgLZEgqJkiqMU9x+qatUe/1evEgS5nKSsEHciGu4IG+2b81USkWG0P
tF+8h+C/7FXTO4iu2/hhljvrT4Yuz+fZyg8e37rwE1sRs8LhMJFYBC1g1VPvHEfo
yKpdRi8QiLYuQefniY15jpw4W478oKGp2qWQkruB99B/G42yc1C7xPP13IBjsMqE
oFA909i62P9vUkwsK/Ps7CYLWJa9a4lbetBZKnXwhyyhvJZpHpwtQDFyqwXKH/j3
hlcUO0XXKJsPjD9r3HI+jgl/Sn4XBSIb8tRG/CshCED4OWoBz/NLrRA0QvfXe7T8
RcDomLlASpHz+QGwxY4ZX4VdV8KsyBIMy/4AgcuxfQRimMyOXvfyPmvTiL59d+mu
gwYybYZHiAN/T9PlzNplmLxXa74eXdcIz4ka4dnhZkLD4hXEfwjKOx74myLMdMZK
jcynhoQYPUaFKsE4snnd9JvV3aRIk+xfsxzXslnr5vkm8vTLwL79yHUK0BgdtCtP
Mayf1n7bHlqgFlUZ18SyjO2HZ4/14X2Acn8MyKuEFqymcbQ1BMAb9TMcn01tCxED
RXq7EOo8gj1cvyMHDEYv5q91NWG8PXiZnq3x2HpnmgrVcIenPH2NsM5QJZ/gnS2W
QDgneOqlxFltfube4njkWWVxrg8ieV/uW7SCZm4dmnYCA0lpiNGgBuBzU5gMX9Z1
OUswqXJ+hExGpfhd8tlbI4JEjaBfQvA0fNlm6aukvQLkS4NTtUJ9RecmeZMJQ/n6
oB94VfW05HHHk45EdA3XOyRmwFYS7+XY2EAqGG+KdKmkXOgESNArV3INlA2BLLYi
OFSuSmUVnRz1IOolUJuDCG5lv/CfjiKuAxfv+T9M1d3voX+PxMDQMWsG8laWnlew
Y9F3kyIcFJwZmgFDIycxy8oXtsUqvQ5ZDdKLoqC1G6Apc+YkRRBcQGadnckv4dp2
B1rTW47lrR76aG4SXlCbxRjDXUOMAExj1Hb0HQ1zyQpermga1HRjectL16kj0tIy
GBIgxZkqhN9DlR4Pt6R++GsETschcwwL+RL+fC8Kefjn2Sz9E4PcWYtX3VCnEKRN
E1M5n0AZos95cDQ7fOL71aK2nIAt0u7OBJTEpM8PpDqIdrBtYqJxcZ0lNjBTek3Y
3jhgRR5evU7gSnGdPpJFIJSL62sStl0qwqRIVKeJj26G5CvBAGFv+VlEGY4HZuu1
qVy85HVTOOJBdiZDfiuyeodOmjwKyyQIyPXwwVGjfFT+gHfBD3flxV0VK9RxFg9P
dalMX/iRua9RGjcvKKLO5Rk2Uth92/GOVsALYB9w/Hm0npDkSym+0wRyXbD3OzLq
jTDTwzJbY+D4+j942Ekdy16b4u1sJxo4x6Kc6aoKPrztDhk/Tym9OOH4s0hG73A1
NIVLVSPWHbow8s1FYXbYduDAHloCu2PWT4aHAkIWpE0/ZiEqqMhExVqygD7HeFR9
M75XrXf0y/Hj4+knXCFYIY/Sb0O1j2K0zJN/wlryqojMICh8mIceLGU1Ti97iX75
hL4JfsfoEI0iYJ48bFzE4WB2c+IOpI2vX2Sy1W3EDO4PV4Yaxy8bHpRKcC67cgdU
SwWxxVWQy9zaAyDbvwe5DAzrnaeTJ0/C5pgv/xwJLOtgtiniau7wDwzi7Ihc9YGH
Z+dPkBVb2tZ+zTuh/tYeqgkBItg1Ey9CJFRNtE7GuEI0QI2OiiYCvzl27BasfbC9
TqsyyHC5UDOylXWhRj5k6LRve9nHb2f+gwTqBY4W2ROvMQ3dzDdPieDJe3p38PYL
HCaTRnu3nYlSjcv1Ypty8IXisSzbrJ97qGGsXC8gtGruyYbRpLaiKD5Du7aVkEyi
mRyQR/gEwGnmZ7zdrqtmDADBwBJwalFNZQgCXSfcrsxABhWqez3CHoEJDaOaXngp
3jCURutd6W8JSxsp6PRF1kkW0dXRDhvhulk0/YIcp1X0rOl7bwSPwGvYmFBM2nle
YqT+6vOZwwiTpSEeEkjY9Ynfw6Act2QSVyQoW9lTamFDPXEdV7X1s/SMDkWe+5Hs
TIEUMppQWXl6W78sXmfbgf8N6HdlH3wtXDWPgabnWvsqaAYW9qWBMBY6QVEVBW0Q
zxIUlZbGPqYB2sCDWOOsMXhj//pjsRg9cOHz1Ld37Zl7+ziu+ZcvS3RMfNrVUA2A
lUO8LpjeHU0qkAMfR6NH3fqXKCCIfZZ6FGC/l3bUxcQRpHnyp3YdzaH/fHqTOIJd
y4wEx2Tn20RSTKTXHA9CZDt9nTJIsO7vraus1E19VpYy4IZz/clWfYMMHLVOKlZm
hVXbHiQf23iirfz4G04OVod4ai/E9LYMXKcoeBR2z6uHCfCR+e4Dn0Qb0+2lvFdx
9du74RHRbsa2C3gyaq/Mnkwo60AheAqvVr3W5DTCERUoOHbAgQaCrvxNP9n8xhHH
NMqz6VHDEILjh8+K0m9POvOqQc65b6tZNUNyE33ng39OH4anFBmkER9J52DzTa3C
Mkrj8JDAorzWELNDwWlRUL72spzx8SXZxIUzoFbXWMkh5Ea6HGK+hydPjP6XM+Gc
fm5kmLeeKEAvw4+4WruoA6uieWz89CCrz5aPqtsjqVHx9uMmQiQT9sNI/Ga0PxwQ
DesIm1X450y2hG6RY5G/OJkPUgiRp7Wc0VAeCHPLghBQO2LEOKoFfZEdb7RUf6yB
ZEUE0g5OMAdRNmMXofAIU6F6hz4CUvDHxhv+3W5QjV9fTQO0zpkLHFrKZ/ivifcS
TKyCruvNMB9ZyMOHiNHOu7GlVxRNGM5MiJmIK+M/Xsa36cFlOPSvFsIPLMxLRDa2
JF56qLRHEpkk1MVFODLIMgeM9uSV00xpOUPtb7eNi4zBrtqJ3PgVOJtT7+3+DQ8W
3Cnt6RGOp74IfuEhQ656x/1ZPHNSdZarSCGoN0gYTgB7yPzbQwc5XCLbhi9D8MPZ
wh0yX5fehvlhS/6IaMQ0Tf091pXXYOh/PNsWfraiunNka6AKbJWKtPvny+dP7/7P
g2RY61It3iWsgdIP11Qnv9IoQIzM+zYbS5DdY7lViWK9UhRwtgtrmF64FaSzgKvm
ZOAR+aNVEkLAGtkDnBlHOOqMkPsYxF/YroucyiMheIO82AI0CmTYRgxCgzMt93Bs
ad/lRTdY0I5vOfWU38KJoQlrGgMzSjUXTxdHVSMJoyr0qMlw+xhWmQiMO/30jxMC
9zcXMvtcIZIOE4tVlHHbL2z2FpY4RUUa+3VeW/zTEERAxNl4DIURj78o5zwwKQqi
h2+CFuf3qJ+ewwYopy7QN3HB3AwENh8riCU/B0TWfbdH+aV64JplhCBf6t8TXZMS
4n13wNEhaAfqDZsbErQ6qcI91hS1DNjXzFr3xLhRAi9xou2UcfINeof4qDAuupD6
L8U1wlXCrLG2kQWAvrhlFRSLYILsR5xN0gVfBAmAXCqKBxsfLbW0mvkeyzg2Lw+A
rWSLgKP0SlcuEAS2Ups0rC3oWbxJ5TWuF54fdw5E1dCbYeoUBFiM6mfd/Kskch/K
iN9SE3Tn1Bk0fNmw5qZTYhKoLQmHPYb+jBuho80jDA15IyWuyFKI/4z9VUJxmgVR
EZCeq+9qu594toYp+3t0iwOQrqUJ/OGSNR0Ph8UZDEdhspjcmd31IIWtc+iwKdLO
mT8IBtaW7MbvoFkfLjA1Px1TuzxYCRgl8dXNcuC+LZnfegunewXJYL7e/lsUW/p5
dYKPH+eejdS0yHJPND9DWhNfoeQbfeZ6YO9AKoWwDQo8ZdGLPEVnjWDm/txlH1FA
Dyy5BimvrpffQnSfP+WUp1xE4SEOR/Vr442L5Ipe3A/gYiNqqFGFh2iyI8MQX5H5
B3cGOMZsrihosoSPn8ngVd7gLNmE4aASBbq8wspRIJstu5IZrXIFbjIjS5eX08SZ
PXlqTvPPx1mr3viFoNtL+u/BZCkEWYcKpCJYYS1uk8Y3o26zwy6OfvoXqgnslaCZ
GK7JChh4a/HwV8QW9vM20Bj6t6qi4YBHf95zeRwfFPY9M1+4fmkXmCrBnotLZNcw
uaOKJS1AIe1yg+GkZROjEemnqaGez8LF1E+8Xc+gXF3Xa1e7CG6AAIAD20vPkVRa
LXYOOZMKJdXh7vxcpwyLKSgtD93kl/lLDekg6HqBDBVrwWaMETkmTL0gVErRXZex
/uS9iLemE8haO4mEZ6yA4JfGJYv2zJwZ4PmcHCQVqxgS9x0UOSJUTbg8Amwx38br
FSSNJliDDF8HqadYmjtiFNiV6r9Uv3czRH8FK+i6g6WMyjOkVltud3cXYXeOCpwy
fpjkgnTqLDRAMyw2W2TI+eVu5gr3l3UBKeIP3Mlkko6Dkf3QECZRD4l38ZKfYC5Q
vaVvQ6oES9skEG855gmzwApNye860kRvtPWJ1WGQKV4s/29O9BoeBWJLqHKuA4y5
HO8xkQtp/twgoaOVvPeFaMm8eDIyBVTyza2HPbwq1s4J4w5jdE2lJE1HFu2bCamb
OURzv7eEWEKWSQ6EFkYNHNI/WoplvLppHlJ3Yfkl+4xRV54Laa4+otuf77+/GfND
iry0b1YUM7/nz05plLWxC9DcGUjBkPXH7eNCsW6fOKU/ASHOnEGzUv1GaSjwADDx
0NPleBWCsf/BxJHG6h30Fu1Lbw0ZVe4wX8Cw61uDBK4D54PfqBKQgV4EP/DsgOHL
TLS0CHSwZyNDiSzkMz6vWRoqHIXCTL/3Anof/eoiFGbxGWpve8q8yfUlTn1jHz6Y
83PA/HlL+mIX9t8sDgpatReakVhWcd/cuPhbHcRlWi6jxVKGM1+7mS6KFd9RRTKb
1CDj9qwAMh57znPv3BkSl+cQXCv1FMasX1FGluFwuxT85xfquLId64Xi52eBbZlV
GYBnn5jvJ03dWsUBTe/SE1/mCLInz4H88nf04NGHiGs1K8uvgvUbCID0Zzmlyo6p
GFPDFyAZ8yn0S3KWkjF2o6ug/PCsKrK6h9MV2zM+nLmQvighf0PyiZQltqe2Yplj
qUcPT/M5wpK1a2YJYU966tvrBe5pv279+UzgJLtByGAQSxX6R2kSjZ+7RsCHsnfj
M84OeSzlAjXoDhVCmHN+jwz8YO4jzFYtJ7SIz59IbKNFEULAORK6P0Zm6DKR2seV
TyFlqH5Ymal9nLvp0fKUy3xK6nIMBdTiTvc1h0UW3lZ0wLY9dW1rCusiLev77TGn
8TTO1wFk5WWIBZ58arjZe2xYobH575qsvWDn1fgUuXD/bbEM3xWJ+ByyXHnS32H/
MpCQ/ApB+DyzvY4Ul9BCHnHmwFc4P0ZDyAhKFX7djRruA1CsNAl6h0bw9QXYE6Jk
W37+Ud6tt4xXsCYOSZnTuSvMIJst6VHPQQikwL4AdPPJyTuBp8c6tvs6ULcXM2pO
cxYKmMQ1TpgdpY+yDWdrlA59Xk1Y+s9fU4gn5s4PP0jQCLoFJWU2NJC9jxHpRgsu
ZyIOkEp8hpcMynhuKbsr9cUTbLZTa1hPR+Rs5IwnlC8iEeOzLqx3MKSoHwj4M8c3
KsVdunlCmMA5x3HI6WXaps02/PGuqbqCDSLjS+d5Ms1BLeulj+R+r7l8BgBaVicY
sAxwK9uikIjI7Q9ueMU1zBnAm4vqormJ9p25XXTDcjkFb0wVP0OmWf4ww2rWycRv
1lP+4WuO4tXTHIpS+fB6C81jBYd1wvKwC4/ZydNtj1vbIlyia5736KnlLFhUbkiG
xCNTDm/oZH1W90Qx0HdAVqAheHvilSj5PZPy+OjZYObdvnMkCZ/2DnO3425zONyb
AsTHBcJi7Y7Ki+qNZQq3QuuLASZjGoz1aquu/9fOc0tY4DVjuLqHyMf94f+eFUAp
5LOgQJEQPMaFCs1e5gnFvRYJ12KJJiL+tTNJL95YsOv/2aolZYn17gRKE4QNtE5D
hfD56u75LdQZ1eM28YEsGivBzH+2YbOwBlE1UOn4gCtnzCWfX0Dn5dJl6TPaexjw
pLtOBN90Neanl5PhwgILKEyjtx68cSkTvpLon6ipAkyL9Iw3KJkLB3xpcDsdcxUO
ZeOGHng7cmGKpbufPfomQ5aoCS6g53FweYLMDVdv0GfHLVYIdH8JSerbW0PwwZUg
rOfOnIiEgPoNKB3uDPAIhAWsQMNOacCaCvXKqg2Qf4tEpGyub5+S5vtvc7f5EUR/
H3zu/U7jqDfD/47lP2sjy8LHeCkLWUDpquE8gJIdAVUv6zHnoNU+SNV0xRGsn5+b
12I1srDyMRZQyPGOfehUPfGrvRBEHryqiKJurm7P5Sf7zRQP20+EWw47WYvV0NgE
JEato9r3dCVopRl6+XjosgooRFrjC4eyx5erS/CQKI3vtD36CqfJ4lHUU6js2bDX
3M3BFFsugpJJ8dugvK17eQ1jMC4KMj9RUE5kPSOh/sw9Q8pCyVzKk6gdTVWtpQia
ngLwPffuoVwDDDX/YCmTsk2Sy+4IWFeFjEWwxaIxz6dr7gUbT49SKlLiUiUpiQtH
k+75C6lPhjAm5Ipq6weQbmKwIDkhTZE2mpK/pQObI45rtIts/+HfxCqJGlz/Z15z
qHU3GWr4T7y3NXKFIo8o9rEiSpz7b3aLTC2nSKsdXXYDilcqS/BhSNkBuP1aLncI
MNNDu+FBWYVos60F/JxGludctoFrPyLImtedAjg0iXosmGz0BT5YKQ62zL55gmb1
O70TViHifbiM5uxCLGNChOdy566FUQTp30eXnQGvkcka+EE4Uubkf0qFviirF61H
KbORKnbmJzlwQsl0p02EBMNR0Z5UxjKL3nfZ3bzpoEfYEYgCsIC5q83mhrxmzlUX
unswR0F3+TNis92yFb4fUpAK4JjL6yZy0Tmwc00/t2h6pSCyJMPao3JsKpbPqweY
zXOJa55HboUitVL7wWzgrQbMWn+ifJQ8oliaZaejhyTu80ZGZYlNRDkKWps2W+xP
tX0ADjKYAFQLnI3yrAxxAFUQHEIyosRkH3Snwoyl420mfjZUU9HCdwVJCra3quD6
6W2WopMoZbXOFX5CLwvbduMM+xg464yRXvUhFwmjIwBGz0u1QrfTSuIbf9TyfdMx
bkjTvVT/tkvoaf4071dSmtf3Br8ZeNWL7GO6bMHMJPEdfWOOTkcwCfyXpd7NESVO
KIVfOEY3fBKYOu4YGahzsu4JVgzvQfMljwpL0IOitO0HdxxMq1KAuim6SAiqVHb8
32pFOiyQS5vGErhK368KnC319KeM2nhCel1H1O20HTeU0olMc9pGfYJGqRfq4F3a
XKVk9nldEPIB0cBDtxAhH7pstqC34qwbTpn7Q2K8dW6qLGnmI9fsp+6YExc9Wj+X
sMoKktQEbamK7AJk02s7s1NhhLnTqppBqI/oW3uPdbaXS8w8IBVHJ+wLKMBTLkZ/
qPsr9H9/zgnZEkvFax36X8WhqCcwgtKtuC9u4hyNk3jHHCvF9MN0jL9lfNg24MgF
O+b2Bb3Txz8OvK3lImdNgrc3PEurbfpwLIuXcM6WCZiq/wNqAF6urNKtNmfHQzD2
fx20ssAGyE0UTAL8tjv+umLHxPUCujN/b9mYaT3ABjaqdS/EU7EpPiqMhmgkfgWN
5jWMUYeY87LOpyC8IxFF3fvkVIB8BHe68sFcOMFCdS3z42uPh4k43iRia8xqaSHO
8rwK6wlQ5mp3bs7YiskmH8SZoxuq3jDdPyQgwq+OeyFesgVx3MdRpd/pfnzuF03V
izj5rLslBUso4fheO003x4/VFIK+/azUgxIgKT2K5lyDeKvLDhXuyWTIAlYDZT4+
JeLBqpPHTM53MRUHIKe/Mtt1I66Gtfvr7pzpl8/M1pGLtjB678MnMwbS/ftcJ640
vsyhSNRyVC3sZ3cB0ylYuHiBCukecbCT399tMlm/Wiy4DDCMvrk2sMTtgduZYYcn
nZgD9lKWZ3ad7wflTfWHJ8WQxka9VSxhcBTpagxQ/ao58+NYtwwoQWprAm3Hf9Sz
P70wrN4OnHG0GK+onti5ki6Plc5NKNo64fhd+iH+5IKlqx/QB98DxdNjffYWykpQ
MdR9SGbh2wOxH+pPH+xIFBCbWhmRQf0rxjKj8T3G8qQjrP57iDaTUDaplwLnNVVz
9CEt/Bfnw5DWf3qHPwwtoMwrDhyVvvWNpfy6FPo6nRt/TutJ2WfYkCdqMHrQdO/I
+E54tqwtCTk73uqKj1af78gTDtilstJbtU9FnP+RrnxfYg0cxW5Fit5Lm8vnzruV
MBHlYFUvf6I0qlWFZV4E6f4r8+gwK2IaeSMfkql97gkrdk0Bjoo/X7RDGZeeEGBF
v0OgoMWFMyohfej916SkywatKELXWHd+iAZon5Ai39DL4B3o4+oIyC4bubm47DPF
TtqH/BJHpntG+NrxOnQjyDNMLAyiV8XYFa4uOkr9VzDiVWGVSSHzDzEgNfhwLn5G
QCSgTYcXAdptwhBqvnAxJ/p0rSihKaRIQuJoo27vS+XZTVH9Fb1EtWmLBx58oJHE
Gwq8ZXpebLuzTa33yqlCtp09ytS41+I2p/7jIzLzR1MuW4MqcgmEHrZU3C6egWR0
ARNHzsookZ1DMkeg/wOGmCQjqO64qz+BDl+HNJuppR7g72VFYrXFi2esm1DyNRMj
RHv1p566g7a/dbkeituaTe94nuHoENbCKD3TXVssVCU5cWgAmGomacBNggl2oZ0h
ynFRnrKbQTRfD368AQl9Nwpi6MNX7zDvZlL2itz1d0xys5/DqAwczos3kI4vJlyD
c2cbMBLN8wUeVjYWWBGHN1W1YF0xF4kWb+EjY8+aJphNWnRwkm75ZZnbsVNhVwEn
eJ1IZR7ZGhiwbqm1c2KnQ5l9j6/pFdz5e4rcCRnTtUy9i4Q2ZpW22+MbXugTMNrH
kknu6kGquo1pZhL1HPiP4QQ7jhPzOaWcwBZ5qK6izJPGkvM4LwypUgSOkNhqm4KZ
smy07cDweO0tSUZV5wAqffwF8OuwQfbkXYwaC3o5ep2AA+p3Uwnd+HtUtxvp7WWL
Y9K89ylmhmiWLKH5p4zGVPrN3gFQLAE2FbPn2wdmCfKv5tD0t1UEJTSKIqP86v6i
uWbf2dM6/ss4MnPvSTFUgxKf6yLNC3zXE1+S5MWKxWHJ+tYiJEoT+RKNt/itSOMu
aWJWH1AicuGANv0ezG/e6qqbwr92AyGaqWQibzkLOQN1/u5zNbhaeo+B67vgmaky
3HKT7eR8oQTat49JHho4zyP/hFhzC8Gp9qBq4orP/HB63ImfWF7gGUaWWqJnWLu0
XjB5uAQ7oNAWVH/yfdZYlVobaMoVAC1h1pXfTNBFKtCUU1UntqOMz9vtdhDK96L/
neoj6vymzoGeSFMdzZ4XnSGXZfoe8Nqy4m6EpBYGC/XPwa2l8UryoIJeF62xZOt7
K1B8EvwDDgByJVuVdvE+FS0O3jSfSzjCVDrhoG5KCKeWFZXqSiGRTzQNjzAqcONq
15KAcVL1F0axdfAYsqk87zq2ne34/UvKSLGAJsuOM8yFfiJS3nSXQieWMWQtt29k
b3MrjTpwatIMMxAul5cuxIHoa1Ng4nipMtddTP3X9RTTQl1kiww++dWwh1ximhWB
0txP9UbwkH6+LkTX4Lu7I6Pk9YhhOVSim7UVQsQDzomk/5GLB4TJkTBg2dvD8OSE
H7KghUt2EV+Z2s9//7Zk7BE1pWFY+jPjubiwa40OMjLcjY6597Fs1RF+qiU3wkfM
ectNIcOAIE3eZyZBhxjXSmr/NpwFph3GGU8K7iDzCtK50DmtLSx/g2b+5Vuycy4P
OxnmCvFA6z/xcyHQkvdcLGrjr1JQyxWBmSToFqoYH7ETUDNBP9jr4BMwlEpjtk7w
NeE+5TFfe443v6jkcIqOdG6DYPs6oUU4c5YToX+TU4dMJoXmW8u4txWGP388yttA
GiOcsskgCEm6d16ubaCplL/HFQe+Ha88L3IftXc6KDimz2aUYlOexSN+Ow0w5haA
/4H8nOO+objiefvK86ugrDd/1NjW8aU5ZmbGz6SWUNT7187up5mZUfg+YmDf+ISs
Rm6sKimsDWZGMbxmI3k7ALJmVbVbxVLEt4cteHT1TnEiE6+m4tSsWTAFZA8YUE8c
XbBpTioKz3e7POvCqG/zk41eAFBDZEWthnK/KoIB1LFi/cZ94jszdEPIv4tXTGnW
EiUuMH5rAOwCy95LT45SmDp0HKVe2zPACm5EhxwHQy+7wMApTLCN0SeqY4VdoQPw
syVojf223WltvtFWOgbUAdOUhqqnONQLnUk4fsiYlVzaI8uhmTK1kb9nkIvyq1k4
lq0Rme8U62mE7Jh5QMltxTgxJ3be3+YkbxJuf5kiovsJhcLyMTyZQsGpnkgMdpht
vpbexTNjFmZF9lxuSec75dNiZE74s3sqFasGUAVUjZJJ+q0HOBkLoWOpmeaTbLII
8hYbKBZNrk2FG/onjoazS9koegXLhmJdfrQkRzPB/YEbvLlqvKXETm8OfE2B1qWm
zT1jmof/NwVEM5B0wkURTgtSHER2rF5Y0ocrAdODoj+ElPbbjK19FfOAX56/3ylN
9VPc393YTyOS2b96vQiVNAGW15Urpm6EGtkFQMgT09bxDclPDSdTkM30PPaIp2tn
LilmhyS3kVASp4Ws7GZwdCpep4yUkGmjpzwduKwssoQNxhwVL+spwRcbY89oJNDb
m2XFTfCv+5zVFHAOhxWXKCpyDiUOmtTA9jcQL5tkpIulVTfHni+ZCfr7BooSnH0N
XNUal2+0p+tgIofr286fQ8PmdEYkMPdvlHbEhy8PcKY8vhB3AfLAlzM+mSlW8r8q
YTax/oK+HlfWh+7xihZAmBuoiQFdNntWk5G6rjr/3yymlXLlbx7gdVXpWCKiI1a3
MHXhtOI0TgyqXF3Afk+wEmWwV8N+jxTFqakc6NwOMRoH9ldjiOC+mTq76JYBGdec
zO1yfW3kVSEwffl3eXmziLCLKse+tEiGjVyMxkSSC1Td6E+1ion+M93vlzcZHmli
xyD78UEktI/R91R8Gkqs7Lfzi7TeGN4oESVuAgKFmJiXMTi1eieGM/vuyOR5T0hX
Sdb3d18RzMmnfM3sLgVx7UygpB15tZyLdTKyAcV986/s9Vo2hZ8QMa6q3JMUMDIV
r8Lo7JnRFTgQRs8d3S/N7+84HpEQF8pHZRoofOvHnUemJBpR2OFfLo63z2NkSYKy
5sGboEM9237ZWdDwV3G5DMOqvqnQhFMP2X8tspxbE25QdA0MJr9VtoLwF6xFPlnx
JyKKEKDIVAlR4tVhCQNPegXwi9wV1lhbZ/J84PqklPExGrQd96v++0g+Xos6sJO4
nox5DJLc5CfAPca/zhbC8cYCO8kG36m+iKVL4NknA8HRgGf6mM4mNbK7N2KHxILg
9CuqQAU2PSmrhtYglAhbPEa1gkfrPxW+jDsa8TVkooJYFXozQtuRkbrGOGrNd844
+k7im2TT4XfZNh1LuRdevsbjzphkKFfHrMk8lw+4VaST8ne3X1Rrfgz1tyaQSoFx
B2L73rl9tw/8QLZ6J9trE7YvrEI2GvUtzhYJA6CyLce9Su03o4O4/7+cfXZ7ug+x
xq9T9Poi4X97/5vg0q16REoPtog5zyil4OaeKsdocz7Lo4NCjZvy5OwBLcuZAiJY
1xTBDkn1qh8zKivO0FNjBV9Tlu6+pXcWxDZOReriEHXBByY7iPqR3vBuIwMVGti7
nACoHdV9WF9xV3oiOHPNzNsdFhTqLw4tbOxa5Eoz8QEMA9sThlQlih4yiuHyHZ6o
16OTetawgS7iojXn73Lkn+rOhSh6RqwleIT61ueM0fgqzOGmw51p4ojYsL6tg6BK
0dhoajBADSeKZ28uOwFuLKmvzBgBiQiTbrft4mjENrDE7QoWgBq6hNrXwXx6F4+K
rOMhujeOxJ576qL7B62KVnUj6bxq1iHhHzaw/9FMw/FdNG5GQOwJK+GVKOXBa3XI
5AcNUGvzOaaEdfjkE/46Uuqj/3fJDZf6fYPsQWsCLA858thp17CIB8XBUnqgR9uA
PMO9trpLUZo53QvNriGBjUzufsLP5IVPudRtQetZJ3dzk5DeWez0JsNcdFbr5iRt
60vwxubv4gcKH5K+2KbtoobkcF3GFx9CdkI7UpuNcR0eG4tQU+Ff04u6i7bO4G4f
bHTolu268O0fMFlHZDQSDMb8yoVhxxBbePlXN7f7wuQo2Dk3szeSd0L1HQKeXkPK
5mwQrjxBz7bHQCnum0waTVQ5g2uuQWuFa8ST001zNFFanZ77kLzzYDQo0rXE1DFS
/xnv3Wd+mKhghPnkz1T7Tte2hV6jAj1f0+u8y2RI//W4V2V/xAmEUDPnOsiFlWdQ
tmMJwms6pa3dMgkZycuUKF1LChJtDUayVtzlKVySI1ZrgHXPSIN/wDjGYt79vRPO
+SgaYA10qzJ3vp08WQJEXBsxu1mBtJuWrXb6l/BOgdmyJNDlOx8RRRBtril2v4jv
Q450itulEA3HEteSdaO9IcOSNYr6P5Anye1G16Hn8f0KR03TeCBLMro7OAPEXcDA
rB/O4mByjj4DXRepMNOyf30ghCzyq53+lFi32HDcH+JgY9lM+N5wsQOu2g7W3alu
IUBHG/RDXw2prFIKSXzWCF8xddk7D/KFlfjJqeU+s+W6oTGW7iWWh6BD7MXCKvns
9zQs3cx8QiB+bjzsZa+vnXF2I9tEyz1TJiC7icaDC8m+Y6X14VpoPxUW3KVravyh
FxfhlRKmroiH7nGiyxrrk2/XtqZ06jjYojmLypXVG5ABhKPe3qHD5bKhpf5XV0Jz
utI5rpGw6bGpVQvakqgWDzKsEuW5JGz4pgRN+/QjaGuYXofHMYESNMBG8d/JzJJQ
pjRe0TiGEmFGr1Dkz/YFe93UOG6drzWiGF1QL8kWc+f91bFfZmH1fR17T0HDPZhT
cuWubey4Uw+oTLpo0YeKq6GoS028Zo2XLIuA5EZQ/RQUJradR2qatSXPtgvbAUF6
TmgS84o8+lwibZAPNVEeHpiiYaeKctqCHAxxoR606b2JFwM1GQgu/fw5xaGDNOXz
95yLIdgyhv2ledoQKvmCahyF962JT+zRov8bobLaFoVZuKVeFnF+zhoMzOGAfe/5
Ix0gAr4OtSp5P/JiuUvMmQkxBZ36gf4h/GhrtGbA5VQLyJStET9l9sQ/WgBzU8Uu
VYsatIqU7b0vjqCPR9UeIqNeigbK+VPhw3Cjh2Dd4M5MiP/WF3obNMPJr1JUDplM
c9Z/uvniYOEWq9UKdKri2ZwYMS+IYME+U5xkX7REZnaGE7Lqd2j/L9suu3CjeN4L
4hG7YgNSHvxYc6rz3avmgJ6JI2XQI9+FRy3gZ+bD/Zs4xWp0nGPNdv73emaM3opE
7BAy6iNPCsWRWLufrXYddfz8R8McRbFNhosQMb9Hl6OIL544o1vQ1hq7srbxYDin
pBFbat3IHJyLTBIxOq+v1CTp4HPY7bTrbarZe/VGDinDk7K1wUa1y6Hnl8eYNN2M
qN0atn3c7KgPtSItqq1neRv0sltnB2SzhXFL1APzV6aMhzaFbtXvLbZhftEE5hSs
QxvU1N/mdBN02D+gsH+y6L3ke/6DoqkTbgK2DnybnvQr2iLLeKT6xkyuV+CuohpH
Ispkd6mXLrkVwVzZi/SWIfFuaO1n3yP7Ne9AzR49z/KvUuBzXsrBeUSyTWOIDvWG
JLOMZ7Ji8rH/4jqap4iSNFiIFWijA0CKQkwDcWbnczztzxwzhhuFdzWF0Y54Sisy
/uJ3/CrMdmFNeADPNT31qxLiPeCVhxvSBeRnQzcFdufZKPP0QZaMUtpUhJlgksIH
q5KBQbouMK6xXxMFYr8K510Ovhy15BtYOKl6I61gmAjQ2s0okfLCaTQrbtgR9ykX
Smal1gxqKh0ffRQbzI9EBEbwkUEVeuNQc+NFLBSdfEkqUV7ddOyLmrpkHeieR9N3
g27FecyFm0ndL9nlGja/gMeky+6bKoLm2BUpUXN5CrjgsqxgysFtBxh8HGDGd2ao
2aly9EH6Jk8tqrBQ04lVhAHh01ky3bKatcVIIT5mOVUD1R4i/ABK21nf4xH5IHCI
QJoYLqZgOM9YeBIsrU80EUGLAiRU2ycnsUXI2pCV2vwP3zXKbNfwnSntJveWUlVI
HFn0usMw6zBUErsB6CmACzm4tQY5G/iTvvnfTv5m+qHWCjhECBXd0/E7PYmqB0Rq
s++oJhiU6+RP7MEwDfus8gZ1fzJXFLyekr/Mtm6DeqZHWlrLVPZkuKZdqEoeN493
ivJmsm6j1u44Q02E7moqcgrHjVxQ3cIWuZn0I4Oxuwtv90fv7o2ZzpU0qCEozcc8
MiC3y/n6+kp2fH6vVSBjFk9dWT5JT1lj9X1WR5G1pGlD2GVOZJHsmuySB7nfzxLT
QCLOmwDzZlmcuk//avWxVK2pKRGXzysgsk61aSTEeJCUvHLvCe8MU/gx8v4Ld8s+
nykzEMZZy4+MnNMBCkcJzjPILhdy4D0B/vcOtpK0fY3TR//BoaMUqI8TIVd9yvbS
ALQ0gphHnMC0eMQHvNdaSur647IsGCyo/xtVBWXShNkzFYjo8Nzi1sxHG6ccGm+C
eXZSI5PQ7HT0IOUaXM9kOE1vM43+aedCagw7iYaOR4d5pvJgF3sDHPekadhnvZ70
foklj2GLHyOUFqdDQSYX2B9nTyuCCvvyuPg4BgLTbaUB1WtMz5A3jl0l+EaytiIv
K1RIHH071qknvTMgLTQkIi2XU+Pa52hmVkisB5JmvDh/s/o2kAvGuh6YZa8ZATab
CqksuvfBOMG8tCs6f7/avgWrUZNSjFtqMP8xgwiH4bBsDj5tSDZ+YIXsNeyhW0dF
sm/bZRNdWA6gxrWp9Bfl2wHaQrKpJrJCIUPvZqtBM6vRt0ux+yJgwcDVWJZB7k9j
i+BxSM/n5qfAnUEUkDOb78jwdrLBXnsOPuJzd6zrbwrb1+QjIo/bXCmsj5qm1IqZ
in8t3U49Vgp4Ru3SlXOiqwiVRc+JM6Jb3ZH144FFPLl640D4+U4fnxXqOPO5Qsi8
ECKwuYjsgJz/L+NBzDVQTTLgSv3FL+6IxEkLGyqx8QY+Y908/4Pc02X3mH32htUx
LUeLebYLkCePQUH5Pc78meDp6MlycgKIuTqhhclMO9IzsGOGVYbC3dpMf6R4M38d
804FDxjExRHURqjRquq7L8mQyYE+4hX+flnCULOT8W07G4GY0EfYbkWZQv+NK+x6
imI3fcI7+703lHS9ckVmTSaMfcR6Li1DmOxeXN6k/HzbcgvZcVYfKdfC0rS8Nt9c
HluPclsi26dnrhSDkCyr2UWLWELETaU4lngL5ezt/uldBfJkeQiromlfg8PRvcWM
YPMz3CO/prUheBUJf6bTu5SLigACkUPmY4m+17QjHGs1hobS24uMxBAFgfbujSZg
gAUpyPs4rMBud4vFajzBiYmB4aMDuYkECGXtN1FbL5/XTSUKvWBZCZP8EQtgQhgl
SEXpVfTIkvLP8Ka84VqHv5spA4hCX+wXvSsdrWafspn+jO3eGQDoKtWh4nJMuoL/
/X2leoMsze7Hs/heWmv7d/lZ5WCAOODb5FJnQWWNcFoGIbSrqoBSBW3OY6WXkl1N
UB0LwrqVAxGoypdDq/pzwjBu57NS5Offf5i49LI/I4S9U0F/SFf98xxUh94o29AC
5rvv5biem7Sz2e/suzXmfSeUoxPjVGZTpuGPyJ8ukCNvimRXw19u7sX9NEhmAYbg
+Q6DRKN8BF8yYneEIa/Da48PGjy9dnSWsM3FFl/JDWXCURMCHqdqUb/FaYGVVg6s
AaK137Emw5guuzoC43MOuu5+i6Bd5383aNTTQIl8eFXGtgGg3ihfa9t9zbxRodrV
3rf6crs/1PSSBRSofJNaaqX90k7Sw3THZU56cnPAAtXjW9RKYY21KuSeV2j7JmiM
dzQ1GwAktiRBvCxK5dfR4QqwRizBMVxkrja0wpZM76NehS/PwIdIkIn2kDXQ7BvT
A0NsEfstTRrz64yBDu8vghN4zbDUVZcrjbox88SkuaXYfqFemAmQYEyv48L7FbTA
+ZuV+Y1MyQgMg8Xzq/h+ViJvgV/4DcWNmA0Tp5g3O8IhCvkAVrdmitciJRm2Q72b
bPmrQEm+e16fMOwizqNx6rT545m7RoIsM+mfeTeUjhprpM/bIibG6U1vvfuCclW1
6ZrF3GqsawPqYcMkvvRw5qYGOzA/VF/pSiAf5pRwZpAzVksn5yXyb0E9HIOE3t/q
Ito3eFdyKYw+Nx6YWTIoxwb+SLzwIz9TNBO95lwbqC1j6ajun0EtDtFBoDl/MhfO
1C3JYq7bHSpiKoMbNKhA4arkcoFEyTzoyKfizir7zzpHwawcNWzTlWePRtUbLtrV
SGVTuTFq05eI9/G+gYlNb6qPOQ0tcVhUDK+DHKYa04cpCC3gPkNuS++3oWZ+T5rT
Pj8t9uBOo8lb8P/a7dVwu6TEPfr8+xIMAGyjNtjDEPqOQdfRpfo9gawOunVhqOUy
M4mvKWYts2289B2XftJnbiXcfxKeCTf+ZlIFX3YTQ5UyjiZMiqfin2Qh3bTMoANR
kLO+2cOG2m1czgpMzUK2et3wPYjWoR3/LOyoZFgUoM3Ytdp9BbzJdAezIkfieU9k
MUObhFvQWdRrl5sEkWmFt9dL0qAW6pDCbBFkj/x35IbE8qrRF0QdwKGS432jNz3X
Jbfe0ig9YP4ZOaTmaGHEXFj3tm7+YxlTmrdPJk3vKTdNwp0Bj+IT8eDK+iwCWiKw
yZDAFwuG1TOwE0dfq+wOMPoSPKsmCK8Lkv4OT4+jY/pDGMVLJF5ANN5W3dza+AaL
1lJ3PSuZPDmf9rMwMQcjO76CnzoQamv+FfKEWtbecKH6La3jCGhP8jMGtquo2bk4
+BgeMR28HtrLqZUU1LcfwNuM2T5RUUmhjCpinxvbLLM3vAgpW5lDcULKRr9Qk8sj
mvBZEFCBSa9UDn7UOnrg7B4BUYGlwe7BBSiY2tRRg0gqmKdZ8x7XL4vT1BpRHJKL
nC1GvOVb6jv6tFZQQXU/jvXFvrAWTnKFPdQ6k7lLMy17aJ860ibiMmEeACEF9iBn
ENJmyQiUIUUGqbwjWHoRDArUHXK+86m3XHZKiDtaA+aAIQJccEi6p5IIeYRbkaYO
oj8aYxwRzE7s42Em1FribPah70mnKcEaN/u4iOOus5g5lE1pVY7tAXhF+M9oZNtj
TV7eZ1GlU2HBife4VlglV+SjVdVYXuU2OavxyEhwz9BcaUJyH+Y7sAqLiDQqhO48
UPdg9c7b3Kymh1egvjAc7Yk4dCunhQE7YfVGcX3AmgpNtrdiJ3Qkbhz5l/BvuVF8
nvg7ZBBrAOZqdAtHg2/ZXHSofxi+tSKEHIDFnp/T/7giEV42pQ7YRsGZn1O+1m6c
NvinXBMEvpJGzUFswPMIMH6ztE8APZcGkrQ42saktlIqhrcWcrhIHvUX9DGVLzX4
GzkHfF8b1F8Bi1E8dPk9OlzvG5tODBIXZnIKTzMrESXItozAzv3rZrL8sUEr04es
ySV7TzdH2BDxdGBiRcxKANw0ZLD5cFGXmwLYtQGBUi6Cd551OvZB31yrzai3JaE4
87luVbrDyYegjl6rCJBVFvq4cvOtJVImPY8y1AXRUIdKjJrsQvWSeMXMYHnWDvOO
NeNCQDftjuYllo3SJ7D0XGBZ6Rd+bKUUy7k3N2x0RZwGX4MunBIoJEURAbWjzwUq
FeRrtwXKJAFcPXrZSFBeu7H7hv7vv8mFy+iACTXP91vYRQnSc+MyGa+hZ0StR7B9
hN1ACY6d1o9Tz4112hXX13IVPqKfnpid663eJ4vgSWP8JXNc82axr5kkip/zlxXP
f+8PP/jnFbC4OdL8iBSnJTafwu+eyG/Mm8o2OQa6UAUaC+VyGZEExDYWYTx49tDA
e3Q7BRQBx5vRkmzoun9HtXEdQrhGbWUE2mYY7O8YajrOAwMdNfqIwf6Q+ngU9omt
sfYblFRqgsfJmK/1P4c+giaswgV9YCl15DNVtC4acGezkLyJSKZMF5KuesAjgApW
vuIvb+C0+LlGQJHVBkm9JioCXlMYusBZOEOKelroQRhvwUqbXdcYfAF0MMpuFCTz
nPr3uKKD9vh7ja8UXOAF0yyt/40KN974bil0q5tFoSYoXNORJYqrnldr/g8nX2aO
c998ubkB3rzU31lq4w4nWBTUqMoxABBnB19igHa9EhPH1KzdAyCuWBg0wFAf1OM0
xfyGkcmS7rUFv/jpWDyK8RPUOxW/VgPf6NsMZDyFfXSoiTIUMpjcaZf4ugZn4SUN
htc0KrARxoOW5YgwSKabHisGmMSsAxc7Zwn44GwU27IyWfpP4EZE3/st9v90cYPH
mlk7+GpC7H79mIjdEkcw7uXfcN2Jay0ToSv75nF6awhHnFzgcBLMHKcO4I/ftsym
PUUu4/0h7wCf/1vvnLwESEkoNbOWqBM5ZNqr4tdiR8MpSSnlIKd6qBlG4pqvi77Z
/u3zGcjllvmi6WWADHFThqANL4uRyMrVknsegN04SsSgNR7D+wm8pQpINnnd5rQn
QJJKakMLIuwjkj0YOUnasitztlZjrs9TnR8aGms+cAmC8y5seORTqgjrEgYhZ8Pi
YvQqTyJOy+AdHxydUJfRNoFeqa/T5wqwzgewinEbC9nunhq7nWt1wol9RHAIjCSr
f7QdJHHTb+McImrfENLWAEDJD/gP33IxVkFf4jQbc9cheBQd3bRMSdfOTbgX0zVg
BZeV6uSoFpgBlUng+rtlfdFK2yTYcHlY/bEwFUUZ8mCxt+VNyg+LGcR07BKgKGfQ
/w+2Dgaeexnfg1tPtsp6QoYoVOhr8mAXNywNpzo71S06ySj4PNvjuE5r7U8eSdok
Pv/L9+puXgHYwav8GregYmBaBKAGfJ/5vzxiErUcU/M3Qi5osB2qMShC12gAoA2N
jR5jcUWFa2L+/JkWLBctvO4/1zuDNeHxrQMcppQwex2vyl/E0VKXT/sZALCUteLQ
ULuU1IeUWX7I1gmfSz5lI8YKsy/KPDFxykO4+ufHP100FT2zC5pG3qyzP2G57qHl
ZKzOfzDKveH1FkJhsy2qk+jpNhW0dZHuUbzMH8cY3oy4nUz8eM5/mE3aoayM06He
DFXsZ5h3J8V1AkXrNRnJiNK8t75b2bFIATvgBR800uoKfte1boDvRdA2836pkmp3
9k9DDFkeHrQhZ2ikCiBzxYdOdNXsdV857Y/U1lBot11h3Bt9idWuJetKPiHB6w23
f31LKAnEx6QObYyJSiiwGwwrdZu0ga5ciA6wJjf4GcqmzYny+wg81bkT7MYtR773
a0iuOIkJOhIU2SQ/ZpxeraXO5gbcm6z2LieBorXs4xih20n9iQP/2hoEgNnsI88H
/0lIIr5+W6YO9hnARXmTGqiIc9TUlRCJ0p1OHsOyg+duZ3b3ZxBDOY2uTbj1HrRh
/0TT1tqDWGubGPwGpQUIn9O33lEkUZuBK7Nw2fYrhwd1aOhIfjfVtNmHHoD+CgLT
RubMRFA+JDV5F9JH72l0WvOyP2HlIfNSjUN17pcC7nP6xfCrUCMvsVQwTCAMiQTI
mzS4iVgPTllybiOnxSzS8X+qCuIvrD/QLolYubAW0GjIzzORHDEMfHBczjMyUrrT
J/Tev9dtUAnqxjzjShRJ8MjovGWDIIQbUwQgWxRmPrichnTbUEzLn4SQnLtkerCS
S5oaJoM0WDZqUQbEbY03pkCcHrwEgZOB6X010l42YLezb+KK1PyEjCa03obQ6Y1y
KtOMEudSaJ1Lds74MHtIpvl+jEIMUjaTKgnnWbP12VDD7qG4XL/1BVX5ZyUI4EPs
uefHf/LzAW1qsOX1AdJp2H6dBJXigk+05gmgpN/Dpp1wA1qkYTZd7uSRSd4+aTQA
KE5owEu9yoezbEOtiqcMusECERr0VQOZfj1pqGY3zbiSl36ip5mjhrXm8tXlG8gp
d3nF4kjBwNKBpx/cD7tzL5j8DnaHzPoV60gwt/g1hW/iGNbJ/amuCMAJlbizE7Ge
DmZnax1bJxpIVlf+9hA52lSXNIvDWSlKcXV8QViEwB+SGwAaKaqXOWbH73lz+mw2
SwtMsvWMHmB1JNQ3k07zIMVBrY0e008ip2Wr/tAQxQjCz0ADtRa2LItierBe7EOn
RUzCEI21Yunwc0RS4UW8NePnKufSqHDBDrAiqJkedwzoTnHjhsPQ5lC+MOHnG1DS
YXIpK8i+9Dhik9fFIVU0F+T1TwGuSaY2nszkN5dFDjPpY/UBCoEyH9XXi70Mdur9
7G6V5HuBAspICOPP+nB0NZO1CvL9QHYvbjId5HwFzpE7sA/biGJ5T2jGV+kNfbQy
e21XsCNlnbdxTGXJREKozFg6wTEO1VLuerqjFu/TdMyvzf/a/GVeji/F1936zrG3
kR7WinKknasPxvB89OTy6iPQpfCvjBA71a5hGtnp1T4GPEkP7O9YkyAl760muigy
cUlA7mZVx26Kdv6DQF7HvxJdq1zKdiP6R7YLL6yPQvc/KzvxxbEM8Tq88EuyCURQ
9NeaYYk7Bx99DkmINmKd9vn7gInqBWBeaozGf7BmZ94UrgwWxUCLE2Inr0MvIobR
SM0DWBT/ppcFc1F6HYbPvfiTaPzX8ixgcdo3EaeQqbclUIKwnkI53NjouraPZNXK
VEcv9jYI+x+ktYTiI0PLyMM7MUiqNyfHJvPDInFSn0gbkzO5DbhW870pzrzg6/ZH
cgTunkmOpWG0h2Ma6j4+KQjikzqbFPmcEeKz0PoeOeE/ADBV7NhbS2iSa0jLC5/9
7izThABUdJFoQOKP6I9KGwAu8VmFjPjlTyyWXYIVIWIY/EegUXByxQXaqDCLN0B5
GFIcDqh6BmnhWv0HNELEMvFj1Lmi0nOFSNohyc/waJr8GdoZsctCcQstIUjBNIt4
Cj5PX3sySITj05w6uU7w70Q1iZL5e7AwcBqrDwTSGN78/nP8KpOxi9Md0TcmfXz7
GNGvQDahEtAKecV0LhvPv45cfGjgJa587uyiOibpol9A22I/69vSO7M5pZX4sbxG
up/eKCEMTIKU1o8aedIuTpGtQfWhSrziC5T5GO9/5CNF5CKfMHIHKZhwfB7j4SL2
dDCX2Xts5/8TKV4CMqyy6R8YQxCi0qcQ9twaxaoSGuM6WklqVaP18m8yrwKS0h65
6kfTTvOod8RuE6vUwsZNSKDS0vEBG9laGSb0xSR5f/0LEwEFQfsboAMid13msgtN
IB9PJiJIzg76tDPjo7LmTXkWi0+CIbcUaxbIS2bLpfP/zq3E3O8sRD607xpEzsTE
NPyvavDVfjbJZBt/VDHrLikwIMQvL0DboSZKsxG9uXkVi5KfQmrzVzYceGK5TqHu
BnTnpdZupNf3Alsjal9H7MLHCehT68XCPtM4PfSNfg1YBZA+2uELKfbE7+r5tCXZ
RV9Ie7zhOqgbwQe481j6vHxcLa9Aau6YjT1BJTeiRXc6Sul8WLMIRsmTbjr16Vai
UjYzBYASDvPXZf1u/TjToo2ilG0oLEpOJxMqJkxC61CuoNCuxfIm7zI22OuxlA6N
eiylpLQcQDqOEncD6QrD948NUx4CbaqXSCZRAVFEIeiFNF1Zn7ziaU0sN7Ehup7G
SPxt0pi2kQrRVoyi9hRc0oUE0+CK0jW9IX6sK9DVgY3Q5nhnoEMSMIQE0AbVMtlt
AG6zExXU/AVZCyWv18SnWDxXt2qEtfpmIffHHCdIdn4A9qogI+2paXh70Qg395g5
HXhqWzzFkb/6F4xYWCRvoM5iIa/X7Ij5EhjmGdja9jHJUYz9xaWFDOyZlS6hxTIF
sFGaQxONzFkp2HpgFhm2nyrKxrxaKsfZgW1GA5xZUw14Jj4zc4fhFbMl7ZFfEuOs
hTdDTlGRXhNfmx6K98E+ATeqM4HM97K+jHBtnnHXFAK10tLg/AQWnC1rK9mXMXMY
Cuhtji8AJ7hnwTRIWFvX6O+agSWjAoj9zRcMkNnnCB7v4av6vgo1OAmhwqd9F6zk
KhydDG6u25ItKoekyGgDGGFFOgAlo73orwTTGR1FL/LaXWsYhA7ACFCHW8ykr9Ri
90hx1rAE6PMZthLVgcLub05x9vDJZWrQVwKhKAUX2SKsI9f5jFlVEe0WLEQuXv+8
cNfxK6JdGgCXFnp4qUUJmiOCkQFB+gjUVd16uMWWSqkAU0PWZyXyF0S9MPcsRJvP
61UbXsXl2NT97DmXCj+ar0Oipd12Arl2QLuueWAgG+D9O8Nb5ffappsnc7SS1SV8
zavM4fbN1GUrZLLUkUxi8JaC6yAbsTuQJPFRgue5mSO4finazeJUJLyVYwrf48b0
XYtXiDN5w+hq6mQOnhPEDL79UIxQWXD9K9tq9toHaAvvN1DHnyEcDqfaUskS+38w
4dmJifvtZt6q52KBM9WCS0YeAPXfAWwrkpXd+91efmgClG0UffOAb/UPk7VcBPg7
8cZpzhzaadp9QsjQm2qeJ3KhahVJP3ttmzZ1HveSZA7eguLw6vDMTivZhPJTCFpx
pf36eVCJzYm/buo+MV3EZUQNOI85IyojeFMMH0486RlKkcYA6U3EwLNIF+VAiWu/
5Are0wVm1EFurQHSS6HV9eIaGMRrc6Hg+BjNEaC3C8aNAFTiK/1KlzN1mJT4xe+h
qkWcR8zD9KuwZaj9Vhwf78Y2Fn7GgdkJcfxFjEkYQweAP7SnBJA/88wsARfx7JPO
2jNBDJNTMiJxbs5YsCYWp0H8+XWsu6pmp2b30ifNlMjFtBvVIsUvkSDxki1JBMTB
O9AjIzrNiA4gD1zKH9c+lSTzaS3EA8NsU0+i3Duj5EA9HWhbHWG1jT47NKGjzxKB
H4yualbYophqS+Fe/PovZQokT/c5T/KaGQVnOIeGoy0u+ZShczMeXuvcKF7huzi5
/O7LbHFTrEEpQvYRLsDvqSBGognM1ImKTO5u9OK3/OgNiSDvua35vmYkQH+F85MD
Q5cGEw4pr2u9jo/45X7ePDahQiPr35rSyHjJ0dTeNlrUYRd0EKK/3se+EN9sN1n1
Npl0luHXotq7RYyZdf3HYDgA08dmC2zZk8umM1bWfOV3wYbgLjmQtTqWcb79Q9lC
B7hfsRiAAzde+7uMZMJZfuLWE7k4beLLCGXTknVXZvKHVDY1mXKoMnRVP/LPU37A
0Dzw9oUPrN1sUyZzMJJUbLDAYdb09z2+1bz2WFSI69VvZajH+DRslGzuC7ZZG8cV
xBCnJkCSL/cS1ISdBB9lKfVp2GnxldZRww3IImY5BOwyJ1DL4uKx3JOEFHTB+V5B
5AnY/3qxUN+tjlhACggwmRlKxq53qAU6SYqJNdW4k12qW0hsENF9sXbKLf8mFGgR
er7zj0xyGrU0jo1h/o8On2DuVpWNIlmsTuxQ75QM6uBrkzyi5LbsAsZdDhiI7+Sc
FQVG3qR9sMGYvuP+Vdg5mlmkdLs3KfqHRStXXcPHLCOnePinv3a0RKruAC2hUClo
MegM605jlxJI2LJamYQJoivzleam0/I0+agkXHQvFNz9B7A1achp+VQMAHjNz1AL
JdxRpXSOC9fP/HiyvpkngI1qX9F+Cib6ZtY3ZgmSdcF79YanPgCJW1VMNNvaUo+g
PJ5D9ycLtO5ZAmijN/cFY29uPa7AP+2oQkdAjVshaFcxcGralkxP+d7mCF2udLLd
rD6AhG5J5ug9aHIkYUHoFpELVMe7EVDUBKSCVFjWpwrGkfrXkxGr+mcpe/UtTjK5
9GQP3yHbFmj45vuxPoxMbh05sMEAoM0l8Wl5drQ6gKlEZnZ75APNWhLE0z7X1O0C
OgEBt4KRC3+q8XicYAwkAVZdZGcc2cwul767ppMbnpRxd5457CH8nNZLoaEF1/Gb
GhIBhKSoo5U/Kbv5as/YrWQqO3A9OlCLqrHhA7z1wqOUlwsrpPleBRwllsp2O8Cs
YNQy5ADY6M39siC7wBFLiZu98osVOe12daG2n78NLzoJMEtsQ2orEq750Z1zSybm
Ol1r025kyvy03+KyIwG9KhQgVlKfe3IJtelo6C7iStDHuqHQMJ0ay0IhyzlShSX6
m0FH9zHtr6U5dPis/up1+mtBUXuDWdnjWjb+3yTdXOg0N5TylR0ihgubyXhc6ONW
LdF8/Q5RcaikQx6AIOznriQf7lU7eFFtVE/mhqmqGUdOTfWBCO6bynbvFfCStJf2
xYnwW3xTzl7qKj8gYq0C3NiV1NgSynivGbQgsMiGRte4UR0ezcLV61OqPoDVfKMH
DNLRgLgBVki3ikOm8xcmXIKygMxW43Ye/akARfNOEsougFe8c/FCmFSoAhPaTWu7
+KIXrwOlJkacXPbMbSgLDyHKzmC4N8t5pIv/y2BTNaKchcg9YvjI/64ZT5m+TIrZ
7oFoOSeuzgMDtpt+RgmEAZV/hNhHo9dL/6eQLCagTO4LfCjWEVFCcoT7tM806daB
9qNvtUNuZegf/dO2DYMowdkzXfhfsIQW1d35EDi/QecnlnczwUCxmetogexxRTy2
vKVy7/fJ81DCMgO2fXOnf82f+3ee7EFJXHd9NCZmRLULnRwINL1DIg5TxzG5qa8c
moWz3UvKOflYOn66vK/AdlMQwdhgOLE/NIV0fdDVL/xGR9jGTbbVu4Vfi6pgThwN
JVKw1JdVAyj+/Oi1OFwY5z35G1pzp8x9rKH3LIizVZa8VEyo9HkZPjv7aTq6Cjbv
Gq+uhW5NQAB6vOyYocWI7yWFN9K4ubfdVG5G+BxCGW8u84bXcNJCx7BNp3ILFHRt
IFIT15aIin6QYxtV27+YeMvsEyp/JfBskJ+U07vCsZOQp89T46DjhUnClNlBRmsz
d/VouMseMZO0aEGzV7L5mYwgyyJqv/l6HtalMeD/gFx0AS2cTr9AtbrplMewn26h
FuvSj3k5jTOCMYz/IlIEQFj612KhsgkKB2ZCYCiyeM/rZ+XyI7P8U3Ix4/7O5CJU
g6ZEZVfkSBdIrVNbU4UXg69KGOCAv+/I320lgvTlNo9TtGUuokDpVmm20u63zOPc
5nZipFsjojS7frRRGkqCCrMzZllYJB2SsEwpxMc1wGmtsEAGB+Wr3FrtYSqaDCOm
OwnGHq2NRdDGnE23cdXaXdR8wS/v+V1Dj2x3GlKuvD9s3fSpRDNbIVyJWoKyBYLJ
piZtC4m5x0VKGDBUMLnjeuaBSzvoVDSUSqbvzF4hotRGXok3cqN7brz8hzlK3f/L
SRB4ZYdKbHmtAeNqTMl4lrmCxrZrb8oPRJc9OZNiuw6F7R3aOZSlTK33EmXMldaz
TUDutO5CJ3Twj6z42wLxARNyME4hDNAyXrKRS92SVC/MI1OJ8vszProUfFW92m7X
c1DIgsGLeleCx+uTHCaaVRd3zUpR3t2IntgvykWAkA8pQZIbNEqkPeucDUmgqMGU
vtzB1jnl8wF5vmvuy53CPCP2LWC4a9gHkxRdH8VRjhd7shMPtCD1KpipJ8oz8YrF
vPN39yk8OZJ3lV772AHY08L1p1XFUeWJMyqZXRVv4lkmn1xYKqFnIPD+dR5TQOtO
gRbLV2XNZsohzJYfWT1tU8/qxRxNAlYDAGdW2Wq38Uy9OZdFCH/BZpWN8BXU49pr
6vA0FUTDSJzIaQtNT2ec2yD/Aaywe+wIFdlgUnZWqNDBJp5v+i22FXgBxasgol59
92NaD+QhpeQPZQsIQ4ccY4SUf9Tq3876hxEgat9T7JKQ7h/DiJkMb0wK4ojFHz+3
mBoV7ePbHR4hgol9/b3WJSLaWdQ1juKVq5wnIAUBtfMnwgTkY8gKk7HP44u2mtXJ
WGOh7kjDX/j4G09qkNj34VlRtcaxTZCuIP78CPhqyhrxPdcbyb5nAs95c/TAvBmK
2EfpViBkoUTLXDC1eFsaRuQshKhnaSil3POJk08vL54RK1ND0Y47VKYNb/XMrNbL
bt8xb/+l4Z5J4eRN/qo8nvzImxWpmMO59rRatLlEZB2BNsZRSjNM47IA9MFoxwSF
6+swkPnkrUPqgrbKSIKbXAMZODjpeyBa8MBNLDkXRg6R2qg26wVEyAby4vAs3J8O
aZ4wybDQ1Ne6cjYqcCVTSIHzaYWXjWSnob1GwPS1BDewXFRX6+tVuG9wN85Xqeef
ZxfqluEi5iI2QNNRoGPb/grRkBsLKU9/ZuMzB5XCJ+b0iO8AvpFQvU0SwyIGsIaE
2r5emvr9py0gyZGcJ5yzPSjIe9wQeKM/fRYszxcOkuN/izjT4ArxnWE6yEzjDCQv
WVnS+7mMPMvDbFcK51USD+JknpH0HvFHUj/CxXoLEWtr7J5UnMSBK6Y2DQzYEt+S
aVZm0ZdOfdJE+RxUS9KP5fuKAyOb/n/k/rbG2Z2h2uH7+lMnfjwpekxN8xnujTOV
u975TN4+nDDIKQmGUbR5ezEWNNpslAcIES0Pn9ZSYvuh3mRboc9pS1cbe5yKh77O
h4Pi/AJbflKM25dNZ5EQbX2W2O8gDogYv6R0LXFvhUzwVxay7agID6Vt2ECcdUQd
H7mqi+sdU/zlEMC8PCjzx1CAHJ+1f7oL7sFb1OPNMA5TRZg2rmQB3epZxIoumJdD
Zg6/BLhMK7lfRzSBxXw11fbgM3tAMJP9so/6gFLVWVjp3R6QLB83drZrR8606fai
WvsODoazMAyCj3gngGtM5xQL5Ie/2Y62nxeUo0+DC/wh/Im+9wPYeeu5UxcTMYkn
V8RGHNwlFenPsEDE1iKpY6i/2cmaxfRNhxXYaHPCrJQoVfq9OSJEbkyVmjIOoEGq
dFAdgCdjfw6DpxsRV1FYAcSQthkbLQeWOAa53vwwBumFoGs7Hsyvy6xZSTNk1fy0
8zK46U/7qwwQ6i/VNlFPpFjp/kNpCYusLhDD7zf+fW263Oue78UJwXkew0WEO9Uo
izmkfhJshcIN+u/W0XSwMKFoy4R/XaLBZqpQ/7Zd6xd4KjMD/7cY17l8pOflPAIj
3mtvdbKtuqJU64KU/yiuBAhiMgOGyzcjUCVCOG7W9g7uq4Fd0Ow0csjE9iGGbZcA
XXlr312oimzlulibfMOQLQ6FIbe6eNULVfw67hpr+4FgtV2KeZ/9aHUNbhi18iE8
U+epdJZuHOSCPyTA8weQvbv/g9TFSSrOH0z/7lj3w4uYzgDfjk7ULiqhXifePsto
PldRayEZ1mpBKDPjVKXszreFJDkSJYoTQ19ZXLJevkWZqp78USSrOyX9B+yZUpqo
X9Ce3SGGJINxHt/yxsGfUEaMvoLNSIT75kI+EGCqIFty8GuNxtVYcKGAGGwtxsdl
W4I2n1WJ++FnBSZEfjOelzKvu9HQVp42otXVBnU53aO2zPjUHiIMds92GV5n/O8e
6rUETI3BBDUE2dFHTSDQnlNZzZBx3PKTkOdr7+uYMLwn6HyGE3DGzw3Wk9PA+DZw
LwH9n+IG0UITZRC3nHQd+OV4LTGr596kVbVgeipR6bY1oQjgF/Q5mZUewV6NXBtt
evKFkFG8p8CSV5U72PeBU0axrgAZ4Drqz1YCPJDGzalQJ0bWd9gQjiOjCdx81Whm
ITHJggWty1k/lQr0BRxqHTL2Xg6G6SQzMq0rScqg7GjygEDZW5soSNu4NldsunSu
tlRBGbehjPc1gc3V5dHTaniJA7nxqb0bcRYt2dYG3RKqlxJx04icbeEiaNKdysnN
/b+LMk4Og1hyAvo8+hsl0TNd8MYUjMYBnefyetkVQgDPUz2ipHceEN5i2TYOiomn
ZiK68d2rI/VgHu/2pdk0eT9QHbJ7LPe+4RW0eDKNOBui6hB3uRK21QcZVq1T3fy2
xUtLR9MA8S8PANJ+0PmS652G061Ve6H5HjoKLnV+OsRu13FiD4KGajm87eH2+WZ2
LljZjD3X4CcIRg9gYNew2XqH68+OXz0s8OiPp1lb4FkVaAqTJVssEMCIYrDBU1mu
161MyccFNh+xLQOoak1sifJmYzHeqftf2+ZMBi/IocnSbHsg5W2YNnN7r0ZWQhHB
fUPdHoLmoLs4FEnwbaA1JhiWTUoLWsST/+MdzsfwPfnf4+Kn5JTYuGySQpf3pzS8
mdfeSAyc0nqKp9vglpJmzZ2CT/whCHC7TqKdcfq7uphYHbYLiqg2wB0hztaXvHiI
unnphnIqoWJeQYda1uiDyXGyRjC3nYAoHNHotChLl3Dw0HsQ2k7hTSTWXCjrXMAp
9HIQnoFw8Wl5xw80BBVSbImRYL/gbtN9waIeMkbofhQoxOrK/buiPOYVVI6Z/kYp
XHGwG4r26A20Ht7y4UskLObl13CjhZg+Ax4JuMnAHG3gDtyCrZ11jRkHXUpdsWdN
64SLXSXDud+RdwEsGZt/bcaquvief16aKWXKnArFrDOUCiQH1RBYM6bOwTM47D6e
rXyqw3EMUiACJy+N3NDyim32LTqsBjwjvxWxsoXVGBM3ProxP7hQz+CcHpMI5VxD
vgcUa9eBfPukw91SvPqC5Ytt6TODZLk9Glrd9gpaWEdWFC17yQqDV0Z4vidItIMN
L1wz6jotv57/7nHkBQFmSa71UJz61qiJNAnL3XdCH/4fEjbQCOZIoAEyvERs5HVE
rH88B4QHPSSf6qCj+aqG4Y9pmrvOYiAsQq1a0Tm+yygLS7TYT8SnH5+pwGeCBdOi
DGan2i31w04P4J0WlAJ5mmAATNAVaVjKpCh8jzcEXKmp/JSVXTnL6rSRVgwx5LGf
uc5La+A1TConV+2A5a2FkfweHZ9LpkhU1D6IyE8XEmDL9+jpUlJWj+G8p/QW3WP0
ZHAMiOaZrjJCRGVezAJlJHLhKnC+zJcwx76pT8J1xO9HRp8qyw/1lG1COgKUxBK9
PGqyQrZAUMCoXwjGVXKJXLdeJspwCPx+OtmuzsO4Hg4i+8dJTHm25aLWYH6jSV3z
HWq69ySY5LwWpq13rc3DMlRhnqqNP3PRTGDmwvtQBEoTOyXw8qh2pTBS6E1UlN7e
nxoULWAHfgVkcck1V2wWXZfSZjYia8sWPd9bAptWmdpBIIX8YGE6dFxvX31wRF3L
H1F36RqiRIgwtJo0v9PowP0fuKD6hUZYqapJrQxza6+HNuot6XUPttTv+qO1L+le
XNrgBsKYERVDsF6OnWJ+66vHQlBfK89cYP71Jj0xAyWl1qUnWUxC2fJwWPavmi7g
PMjHY8QkND5l7RpK4YncbQ0WKIO/KDI7AIDziN/J3Y3z/8ZR1YUz5x0Sj9ZIuiL/
lJ4zowWOxrgwNYGRAClcZvNnGF64HTGrjTzxDY/tS50yaQ45fU+9dE7FsQg7ugOi
B1IVsAhp6NbPFBeCdCb23A4YSJfvZixBX/HCvqIEtRG/yAZY98cl7oqTqDwRN/7l
hEkQpCyhCVvLC5ecKC3Zf3wXc4aEP+cGG8miuRmfT0VBsNpRQfyx0ThQSH/+gS/T
pRFpRfzk4eT2URwTxdxivZY5LtvLiu/XdlpFaNDnGY2m6GnDOS1lalhssyZY9+rM
5ZcQ7nUNmQq3AWXoRIPZpr68M+K5nwIcVe5f5ysMTqVf0SbejbK94roqeCQyErAg
eyDgUUeQ1k7wrZeZ4Busuls9ndb7HV02TWcptK9rfwLwTPCplM3plJDPWwjqln58
9gjvSlowHSXWj/7kNcLFjBfUNxlWT7/0oaRyJ9KUbemu5uWLYZUt56jZNlNpbiz2
lB1ytXXRP5mzT/Cao/U5NySYxDyi4KarQikOsCXKpVxewWU3M1j26JYpf7iffv+e
RwzwjqhlydQ14hUOufwBGxcrvpTrPpKeBvkOI3mgAfeJhV7khYCMts+7qm3vAuWf
GL7d4rs+UGhQ+VvonLPDHAollSuY9pe0LpHu5bgOXVimmAquxTd+oaYy60cPTBRo
W4udPZMHRPlLVvhGuL+mjrnEjF5YDZ20qv4kw7CBbSEj/LVbgP7mBNQW13PZwIT9
MpnqlRl6JXZ+AU0VdHxKzyRyorH9mhT51nOxJvR0sAE+Gkj2vE4tknlLFSo8Lm0j
WyLjF7ZhbUdGMdgvGzgNxnjVcj90air6B7OKW1MRebvTfi/hHF0EWBokeVTW5AC1
9oAU/creUs3rg1zpZjzookn5yntTW0meMdR8aETkKfEH64Yq2RjmugxQC6m+eczJ
YqU4xzwesaAP87hXizRfUy2pzX9c5v8/Y9iRIrKL3tvPpB7aEDK2/YccGJnuKeOX
IQFStuexPsGXXE/LgvaL4ujAsuoV9LUzRwYfv1u/ryFVQh9jzYgxaPZX5OLsXwmr
1HcrePMw9wqpfSfkuYhM9/8/5VPqJYmdA5yb00kKGau5yvdT7cM/jUkdl5p5Vo3M
awPHYeh1Dlgx+20tnqmdejjmjwrdUniOlyeWsnI+q9AIh3eDHzxliN5/8L+y3BoG
NOBDYEk6ZNr7E6BPb8z3aR8Ng1zwXDHQI8p0VbC8wDE2hb7WT6NmujcvTWQhB8WP
a12scj6v/ikB8xGQ5+haokD+S46ZkW32SwuC4PEbEANqFs+Q5x2sDoJgtH6Ww3yW
iDYu4nDuBMhD6bGtJRJPOmWvjzD2hyfUo/xwl2wPnOSUUpISmyoEMkCnzQMvDKwW
K3OmjPLOZW7MsoYHPzXVWSBqXeeeWjRRN5p6eG0g5/1aR7lNnpMW+NqNw+7/CrMx
m2/eNpPQPDb8X7i0T3glHCz5eYApBKKaS5uJ2YEthKl57NwLgSPRftjlYkxSWtzZ
Jmmaj378Lk5E2Z3PpFf4torPQCVTCrowkx6FZp2UEP1teP77WvfnQ8kAHW4hCrK2
HnWoLIQLMVHJ/8qJAd4krlKXOedAXLdXqXLS1Vrr0+lX4jKsetqhhdvAs9JaM9AI
rPttMFMKCK+NRNsHq/wbJYSWM4GuV9ilO9AJk8Kr+F++5ZMcmn+mv3/p4IVHDp3n
LNKnlgcHFZfbbKQPaBEV/Mt2/pCOJ9W9SAis4i4Jr1HXjLx1kxrOClp/ATz4IV/x
6g8SNA12XQxxm/p9HjChRkwFeoNuQTtXocrYI+YNgTKSv/eQbcxBJyNhYHXdx2Th
QYJz6NLT6kI9b8+HEDbxSNCaEwyQnDqn/DpA8reSKcHp/VJrbhR62Jyyi3Tlntqd
z+ToJd3WVO4Nni+E2xUIQHAWREsk3+HHWtMmiRmrwz06d4AVywTU+llTVNwlsIOf
N8tmP3wRovLHbePzRZ2tnmmQQUx3FQ5yIDG3fu3YLaFPeExPoc7QEmmtyP+gTHgt
uUGhUeLRux1+lGdmkJkfU54neKZAn0Xm9w3pJVBuOOrQulwBa9wc95Zc5tWXLllZ
iFyBxsSD9LJHyFAprKvmHxZ5JKE1QBrOtioxSu0wAjjHngQHw1++mFFI9Z9LDOD3
KW3z9J5Ce8//Jz1M2xcL9p8UkRpn2amYEfnsmfhhyDHoIupS0eUcRkwC5owpFwYD
LLjuNrXRAOwdj+9EN2KvUR/SdvdnLkjiSK3LENLFjlsHHBo1DZzFsNEctunFAsEa
CuYtMm9/WncRaEpJbprr6qyZ0Xmcumn7X1ew1ZXuuH34GkJ747F9DyzNhs3MPAxZ
2W94vR+zcJqk8i2AViS3G5N7C29kU7sY6y8CGCF2zytHcLGLyUlsPM7k7Rm0MlMg
KQCFguQ4LnZM7JWm5FvrUALd8FZiApOkF9c+sNypmawFH2aMGv2lb4Dfrxf10yds
Leh5euBTIX4P+K8FwgXbze86goIsiQtuJvKxHlSwFYbSR5FS5cSxhW83N7fOPF4U
Sv1P3USSeAhNPTcBBWidQJSA/2BLJWgCySfpu44O2vX1jmEGFYorZzPp+Uf9I0w8
/wUcQujvCjloliKCFek/dpRKxCfibra2IA/Wqy6+slQJDpDAuguumypeRI63fgKs
2KsyAnVuUJwGjJKY7DLt6xwsS6S75xX90+KNI5xC4qdy8EOhpaHd0YC4rWDV8D+i
NcrHqBiKLQJ8UtDPbGujrbWQPJWV5wNULuUTwSXihKVv1K4SEVDilrESQJoqVeKJ
k/WQkULHkfQs3t7eyahT8hFjio67oilWL3IWIzMLrWywhU3i4XPPhaMxrq4I0cPw
8fPTCwkhL6CYsoPjAN8gqV1ySqVd0v3ptPgGVUOwNMUCyF8XXNdd5wB1H5t0+ScB
P2KygsxonGeTIJZE3KOTUqM7OsSYvEpi999iyGLALgUx5kEPJuFwmp7NcwMziAwm
A9HUDN/vbVdG9MV1NSjhE9qu+bK9kFqKajytt0O+tsQ/we4rW4X/80aopXbGdPPT
JV/mwAhOM6AlDajWNy9kpj56LIUNs3sdKHWa74nN2BAFybuyK9cU00+7W8+YB+aR
PI6j7KdXr+3bEhRt4j9HzrNKw2Fcb8Ha2T1I6HGsI5zAdbNs3grvP1j/3u4z2pil
xSYynWTUfxcJz3Jd43iyD9gwvjkJCRTMhAn8eFgJtn9cECODpWgxfwM4aeDHaQJY
EJQrkXBzZtkEZrudcDrbPZ4mw5unNf6xZvGiy8d9rkf6XWlP1eIRPaofjZmKXZEC
71FY0Cq7n2hmwLCGQw1e95f8OGd5hSz91/W6aextz+XNgo+ycCPLRb6OYmxwUXlq
3pwV/ukfI+NDZAF799XfX/aEOQ8GMs7ry0vfUOrzBIsv8LPqsZ74uVsjIIMq2YyR
+GP3hE+saar5Ct1rs3J5PLriIP4qM1Qr2jrV7GC8Q9p1IRGoc+JgNgEj9Cp3K4t3
42FBxnqxg4zMaH7tK/ez4KY7XVGfhcJ7U+MRkmRTX7djXqCtyx5zbiQolEoWUZuS
Jw3X/qfQ5k+fQPdExqhSlMEu1J4G+Ms+AFo3vdZhdk5Q7aIjUaTh3td+ieJhEhxR
IUjmv8GAk9Gbu5ejO+TxGMLd+tTEzeiXWdGinSHYOTL78RD6Y2qdsbM6ma46gl/D
2IaC06Rqn6UYICQAL2mSSRSkC2ZyhvtaIBuyHIDN8IWpACHF2cl2JoaSWH7VmdMF
urNbK2zbDyHnqp4QpTtXfJ5a0Z6gGBelkkGeBQQ+nFiQ/7/emtW/mNg3We0BKozD
vmPfrDfbEIb2yj8oCh5vq7ZjiHEXYKFjn+iFU+HqxdFtncKxaqdGKwrnN2nWa5+j
dkq89hGPD8QsLuHF/TayWr0to9NYOBB7LU9WM3buqjD4k6Gd036Cwf6aRJBd9zfA
wBmg5+jD9cmki0Hp8v5c2oyqRTR5SG5DyUKkCpUysfCl76rIOJ4eWCaiU5RN+6MO
NN/gBkg/ka2cTJ0p9fyslNUcrdHxVw6cHdZIFraw/qtsVQQTLzuEYuvHg1zROZf8
v6JbPnlZVSyVFf03FFw7QB0x3wErooyYEq9Q1TYynz2vyeQFZ3eZEVClB8Z9zVhp
PUC9xGKo59z3C3deLMUUC4iPk3dwY19ot19Z99Lo4mzPdV8dJsKfrHrXUURXMW7l
kD2U1iR7UDfd2KcA3W3A/O1ugrOSsVg7eUFLnfmmtgMWBV8yC/55gIe4ZlT0owmf
abnlFV/ggb9/MYxjBFB4WstOZemJTacT/82U+KL+3rknuFj1Vha+Rw/O1HCfM6LF
qSQVsOpAa/7bIZr/9wNB+2VXk00EzYeO75zxHuJynoGHQbaRkx45QLdy/wUuBc3A
vDfcCSvjcIMxsHIay6sAU46G4YbvMYRgFYSAwniTJdtLFWIK689WmHUIilR2+PXb
t91VQQ+r5J6v2Sm5cef+YiffGN+cUPuUVdlVAlN6i39f6ecUuj1piFovkYw3cuuL
zEkEXoPB/Rkgzfk3Iv1crVU3v4NumG6FeTasqCuWkc4FnPuM+CgrBdmIGCeU+Ibf
oMojepiFoVYZX2TushS4+QY6Zac65rZDcPSoj/m7UXN+9fPa5pnCQUeAoxYXWN6p
j/IhwZhT0l1G+H2Udu8o3FF0ncjaHRa9ryPAYxX257uqLY1uIXOZwxSiHuSV0MLZ
Ej/nwHizNOojja3wbJEcWnLVqn2MmwY68PQH7Qk3ijxEhT2YZSTF7BQ3s1Rx/Rhg
5PMpmN7b5j4DmVNRSVEzwPqeNEyDHCLbLToJkc80rgvjPGuTRPhlc5WIR3UhaAna
YArVjrb8knUzXchq+t7f/fhHjlG4nyS8tdDnqwXjcUhYz+8Dzbdbm/dwSiIQo3QG
kZxV/G48PJU5J8YPMdTjT0lf82OJkez2Lz/BZmawv4maOYB5xtCZKHaalbKPCPP7
mrCokNyssE+gHVPSo9/Zo5A2exEdkA92666nfBX6exrWPfySFcSYGMUH5o4f75r2
wNcsWJ+wa2XIjVxcEK9/bavJgnty/qj0YF1PJQHZbQUT8/WtsJ+KQ7wA3fYi0Zif
66RsqdVXyE3pV9Idfi7FdL5Cr5JHFG4vo5i1TV7weO2dyRJ1ZBVEl2WS1K4pN3Nv
KMyM8EU738o30LfpgfnLnAK9kre9B4P+Ha5vyFVbythRJ3YnCg5N0rUWVFLr2oUU
4lNfx+Htsz9AwXxxBmJzbGasK6hBfSUYn2VvMzELvOK2Z0pZr8l234mK7lSeBKAl
l60Jwt6Gf5eGizoJxRJ0lPntxsFXXQaeyxAiu4Aq2Jz5LgXr3cqMz6kAtz+V6fpt
A8A78Rom08JO7ttYADFmLdO7gXeIl1rRExiGOesdTdhRYQGPdfWcNeLdzejzcJSR
ijpw+iodbERUF2VW7sKcZCHdUrH33fHdl0I/tXfy790D2SI90PhzZcN97UyacVXX
TRUkgWsDHIAj67X+pghCV/hE6zk8qKkh6JQGqQ5BBwgd8Bvlz3tyc4q5IeaeJ8PE
BXt7d+s9+ayol8N+X0HkXr6clbbw33qAd/0DrYV2xsG6ehsvOO/9B8HCd6iZrO0a
drm4wsoZyPGBdx4Q1Y9tX9jBJRhuqE8o/lqxI1qQ+u0803/iN0TPMl2nCgP2cr57
PW2juI64TBQ8plbsnp5MAdxIw1fy+bzZaCOvy84CjegPCu+UNOIAKAhGJQj1ocHm
hbx6B/C1pHBPuNkTGUU6H1huYH2NAGxK7ZTSYTjxPn7WblrVgEV2EltxNJXRmhL2
sbStxFthwOp4424hO4Xe4BpkfiEn0fM7u+rZ3yqRIRMPZR79QoZTMebsP8uWnqjz
Flo9XNj21OVvX2qghOuO5EhGEqGv8Kbt9Xh5T08MMC6CD9CyKR0tX3Dd9ho0qJaj
n1L/FYle9h1UdmAOpEJ1+6HApMdkpa/0Hk8LZBLvbs0tM/A+x0dLyS80P2OOzHSj
4VplnCPc92uAY2sHNnkCMugJA4KAikmOZU3VuHIfPHXsDChuSgeblNqe5RHpiHN4
fp4eV6osscIMz2ctebuaq2DhrYVjiDsuqvw6VovU045w7huNcIHMRWvt0EUZzKP5
RBzszOWuE4WKD3cKc5lPRmf2ivAr4PgJL2sBHjVlfscHN/cXLrnG1TNc+bCBplKX
phHk0NqnACMoXLr5jNV8RGtkpiH8lrU8I2kcoz+inRwoSXWqURfarCnzBBHcoKTX
yd0ssC6FIbZnW8wLfO1zAnnQHxYPW6su2fPL/VM5xbSfdLWV+DAnKpCBxMPTvdbr
JrD9K9JUAgxRqVAXdT5yveabDgnWQoaSlF4o1t38vFR2vtACK1PrhNV7e1HhSdUp
Zxgibo912hliY9L3WacqzPu7zCU66oDNB0bZaAWChXIeBRdck2HIst/OE/zbOsP9
SyfI9gu/2TKna+fXdfz8C+jDZSY3rbq3K2Yacgck/wX/YukCumOP+Sm9XNKJzcDZ
kfNE6Ajbb9IyVMS7PRGlKWJXYdB3c3CtjgTZNwfIFfeYyoimbQthPCamNZVlvD95
PonKBRpcn+yiHipdCsv8aXbyLN0y2qXXTbPADbIstiXJywtNFahYEkR92ma4paMQ
IrsDFRaeSwU8LeaaQ0ZDufMoHF8l6YOyFV5A4INaqR2aeLEOepKwQjmfmFkkcpAw
oF/pR4BZkfjtBNt6YeRjCLeeA8eQgPMwGmusq+HFcYJyLO4Xn5OgvvDArrcGQFH0
i1jPnJqyljNaE3tqCbM+rfc19d+BAuWYuXImDvUIPcTxhtMNTYKfppJyek/njFbG
N5I4UiW4DMI+BnoMYxqwoa1SqKQUm48fjdTF3NjYUPQK9c7uok011jEMqtq/H2m5
uLOpz1Kb6a87LscGyXfjDTiD+2XI+cKtd0Tuv4XkAek43+AJKt81RN20x8Pe9v0C
Ys1LyD3hUmtaumtV3DvYDmp46RFBUQZJ4CUcYpCjcSiNT0BBB5KcPbePM5iYgSn0
IKntAdB4F15YMcqS4FQJbJH8RCywZYjtjCPnSr9ZvOg2gbMbcCn1Wpgfxfo119g/
RlJSSg6jSb0HLieDGRZuSMacYDX7p6R3Tq1+xiPcPVIqpVSu6ZAxYZGEqtVkgdeH
mp38qmKiKe+h4aWpVs+AFrTBPOnp83H1UQYv/bm6zpIQBbkgT/0mOz7nAhtPgDQs
SZs5go4YmJTtkn0wDIHnqKcqPImFu4vaYauRnP4Klmf9IRQCvO05I/dm+di7vyxS
TuJI1UnobKi/n+hO5OmeuEZlkC7wtyfvgVICVM0T1acdolZi/BjXSLckb9lXlY0O
uc9Jg4Pge/kcyyizrhTvWfXKNIImg6M1eZira8ydyPS49iiNRdUnymRsR6iEiGxe
kcYtPg76TR/qAGoHppfIGD0xQvdaQbWm2q2H/ef0ZO+QGteltRm2w4yZ1dLh91fV
2Ll4WbajjLxMa8BD3m4sJntin9jBN61JO0BNpBU44UCECQX8BJkz9cwDt/zREgnz
cCLvJlr1+o3bNsw6g43TWyBrszxawyCmZGOriwx+fIqxj6JY6eQH4QvUTqCKcqfm
450q0zR6wHPcK1WI9qr6FGyC81sd67Ya6NStkcLIts3MV0e5xBNb3Znuu/BWAyPv
me0ucEs1QP5C66M7uKvb2QdTLu/ca0l+cNY12DAIOXVuIEzuqEvWWlCXHZYqX0ct
0xfyFb1gHJQLqkWSfADQu/U0AA2qsnT3mYi0zJeGq2N6RlVaB1NQ4y14iaDMRb/y
hR7zxzc9WCv6LaNJwZM6fOS3FLxMeWTUk3mnTK7n4D5GCoiy+eu2Lp1537ItY3uO
gOM+sGOI7EwdJxJcWbiASBo+xQAmSwU8EXeIUGhwQX0IF515EvfgmWi4jVchNcJn
qsk8Ya447lfvpyldmE5156U6GC/RZ47aXIefMeACs/RL07LGhxuLGpsD7oSTJFUk
hT9DiCE3hMEsHe2NbIb71ZZmI6dkSmdsUhNfzHDYLV/VJwkYAlHFQKuKdoR2gty3
OPa/D+btyAdMPCnTZ6cK9ypOxHa2dsTDmUFZeVKsr8qv8WLmyAxbGmkBIdGXdoC6
3ZTWJFb/kx3b0M5LgxRz3J/xDOHBLV76dEXf00uWLr/wFFPgl+mHnvsCHdYHooUp
TvGb5VC4aC/iAgUSpc1yAo45rOOgf/0lCU+l3/uorzGXB5j3VU8VxBKUvdn8bIHx
EMVTacSRrLibZZmxDwFEyqEvxsub022O7Iy90Ow4IvTJ2Xoi+BQWHj+Vv9qebtqf
iMM3qVmZlYuK3S+HE9UUKIyFPGPwOl/vLIE7TFRucfbipWjPwVZdQJkiYy4Ph4pj
Pn22/vEtsmSAhJfT3vT85xzDa8ffhPApBcuWH2xlrQaYGcl74yviMz6qWatsvo3Q
xIsLJFiOXKNG8LW7uC7GKtvub+0HbB4NuOg50UsC55vDRyLJXGEfKrsMyL7J51V2
WKJ1FOhN2iMC1DxIY+zFivBeE7HPKu1B7HhOiGGu/vKWjaVM/h6oR192H98uF9oA
/r15QPI+0qh/TCnIFf3gIUHeOIvWfhRjLxLs+vivAzGxgdOW7d8CyDhcZfLLKFRG
zO3KJwvh/2avN2Yisf9y4MX2Ibgtloir0OGZKGeMN96N1Xg4eg8tQRZc8hXMAp8s
O4gsuMkqxEXmefvsKp6k5V17bs7kG/3iQc2hxTvKx+aGSApA/61MxXhcRMZ3i80p
zUXIHxWsg5OacnmR4C4IErAdJ9i94QOrAKTKxrT4+NRmOwZihDFd9WuVE/LRASdr
tVIaX7BGjY9NDeQ9S/eCfmQeZgo293vq0Y0H+LSlXKoNYXVMdzF0Dkxw5yudibnF
U4MqlOhVnq2VPMPDQqcYF3TZAV5DCVVm5mcY1HUJb52xbloEC71d5MW9CvScvz+S
CHezcJhRmozTQzzn7J3g8CVGv/UMJ4aTBCgyczxCdLn3aXPEcslmDm9n+4P6X3RV
2/W1dsPPV63zI6Jr+O8yjbw7vz0kXGaNXb7WeoKMB53IyYYbEvCGGP3JYfHREK2G
UpUuxWIy0ILVJAalVjbGeniASIlEmSBknsLDlKz/aSy7ouoKt8/6Joh8XzEMQY9V
X6Mlu9GhoKVnlbHW+NHIOQY2uPXrNdGufn/6x2JGgdtyQzcTxzXXoR5n73FCYv+p
/nCWRVZYC7zBjNzDSFBwBbrHzywrGdRf2TqVj1sVr4iB82f47Bj9cEFS2k8Ufaa0
QlRBdRrG4B32GXHni92N4DtqGt/ZukZbV1fXmonYdoVGyzcuavcAc35ed8CwPdLT
R8/xuUCDZCmNDp4gzhUxDMi3Js2AxTNhVkzXgJE07B4ADff4Es4JlXKG8uYnbazj
bSdNP35tLusfvgUfF8l05biAw2zH7DYj2u/WxFYA74zstv9uFCOv/20mq5xT18sE
x6KYgocnzaDD1tS+3JHFSkm1KWHN26QCNj7SPvGC9TqGbBqMVGrnx5C5/Jw5mcC5
1QM2Lbf6PjEdxrSvQd/n9E1Zty8tERw1D1wMQni0r4/r3mImZlgGjybHDCgF+ZXu
p6qfVbHL55Mcd9lKHL4Pf8KaBgA20VO1MZO4wfJFLLUIoU72xthbMBGznowBYtJ6
58dllQU2pZ7Eyhr3ZmGFhrGgBNbEFy+hN8wG8F3Rk4VWjYYts7/Fwqn7pUSlOz6y
W/OmISKQ9j1JqqcihJBHF086NILraHgl8me4nVR192F7SFube/Bc2n7T/YBvjglY
w+K8JIZ+Tj8AnjgaJ2k3Snrf4RhaiV16zQNvWW4CFQSSys7nNo8JVRkYQUFke5ph
lEOZRQBne39PBemurxj7IpvNtBUXTPb2c0l7dCSwBd55TeKWXk/a0Gsfi3/z1SrL
Za7X1Sn+PvYs/s19ZjIVLUifpm/KgZkc6m8XpRtltVP1AqcEM4zydFGdrerhE3Ie
OZIrq2uTb1Ov0tHYgJArLKzpGef4bpo6zO/MnJhAsM69SGhKJJ6xpgvl9WF0hlGf
bcTZsp4t4yb1B0K0vt7aS6htkyMrCQsMadp6kiL2MT6nhkYXTInsmkcNb2C9FNnO
t7d/3d5OPOZIvgQHbYcVc2w+aomfGOGvur8g+swWIn9YZFll9b1FjX/N4gDiJRZK
j0rRv9y7PSHw2sT3yVjuY6eDQC4Q8NAoExpy9PG9oesXmhsWWVhtbSmqavXJx/XO
raLIC0odSP+9jUhG6JgFjVvggZASJuFGnC9EjFREuq526/yjneJpOQtyzuZjLIwh
Gj5K2c2MvjNY1zoJKnkVopG0/8gcSPe7OVle3tpFEQEHcmwdDyctmMaGImL0XCFd
rRRFNQwNHSRogCUmoc4dYGaPolEe02DXvCaNeeoeVDGxlEjYrgqOpSeAJXBU6MZQ
rj9N8+/RvWtVNkORKxQlxvp+A8glO712tkn63+fDXlOGOdSnVNIEwe6I09zQJPhO
kyWtpI6TeW8frCOuGZ7QjoRtwlhYKsGcFDUaGvV9dwKb+uQO5eiLPtsex/2V0+kv
L1ekHv2MF1EfKFHI6C9WAdStcrBw2TppRqmTwqPBmbcfuSkdRVd9l+Ew7UAhDB6Z
v9piiQx+vQcVLcAww4Xjjf62IxPZg458sWhOVjadCopADaQPYsingVQvlIbV7Mmv
MASg3QWedSmotPFX0Ly2bks3rY8ae9v2fm+HxSM4KEsslYDADRmz86rk68QwIV65
na3NX4AedRFWeuDUTx+ULAdjUU7XSYCyr13xAkhSpuz5Xq/yHCv3eszsNesv+KXX
LVXD1wM1TR27TSScXDBLiPEjm0ZlRaYYxh/3UI7OL6OVMeuYRiN/Pc5Pjz0SPBGo
nS2l+5KXAo8q9cEYmMyl9RchKf/JVCzE7mpSS9LbSHVwafanNdyhP5O8KXXZLE6F
PPKurtnUkpBriS07z4uomb3IpXEdmJV5yzu2nQj/ZDJFrN0UZs8PLfO8oyuwCKWp
1330eTm9sbiqofAQ+KzlSFRFyGIlKExkgB81iCGnwBHG7HM+QYL9Vhu/MqkaUOnh
iueAbzX6G0YhJEwmfz5QsUybVgY+fI1xP17EVQUQEQc00rrhsR5mu9QQf/iNm8Q7
YtrkpROxORHl0i11XIiZopNQv7LAqbRBluuLDqTmlnB4yf3aomdP02qfMqFz9OSn
pQLZvQ+Cksvcy/wUTCsl+MFGO2M3XfFuAWNi+QHmq3+EDJzePpuhjfYyVOcJw3Cm
RCX9PtbxtIofs/E6fCqrvI35Tvecah6Yz9KbkJ7tuAlyay+wX0vWimbXbxTEpK/B
7wcFYKwp6OQYDuOp/B/CHZTHhw6Sq5xd5lD38/9o5jr+yzDJuCjAFc2VoBFhb1KL
42in7UvrETtydqZ4KPObWniD3umw2ZJXD1mdHGuNusHkdyiPmxAvUhU9LkEALX0u
8MSoTRP5Dppj8Q49Uf3NWGJ/j8ICuxQU+9rXCn/ONGMiEOQ7HaTJJ6gSsmb64mH2
Jec/mcryHxkqX21WcPgY1LMcGSJm4e7Rg28Lr4VMkxnTUYRThpej64nE8DhiFHb4
vMgTVtP1zkZafrAGyNwrvGLj1uLDVgkUYn7FErj45xmGipUOM141Eb9/9VzJyvlA
7YFuMECfvE5HQzkO2yYhmar26RmyHst9ICJjFanbs8eQP9Ci6tn5bX3WLm4iEUUN
2ijySjCbJ9ra50Zlp0M83tFJjH9T4t4rr9OsfF9BeYz5b8gLq0btVau88aQlB4hM
qJLVkqBP96D44bE0QhJWE3T4x1RwSzrwPkergMNXjDOCIJHrG83KR37uuQ+7U/H2
R931vQwo0ZU4vuLg6cH5iXH+03v547UVDWkM2OCKCOj6asxOgbsg6MhvSme3x8Kj
QBr+wPt+RkjV/nJbTkLSpr4+r/H+UGYXNm8jDq8zN/2AcfFHvxWha4P/yALVSqKa
9xKKXCxus+yKLCy8vxZSiOFT04kolpyQndfaZkIUyj85qRgpRqoZty1htvHWcDXP
piOX8vFVolJ5HqGNGnEruhMB5pIb7YqCNLeScBQHxzRg168YCgt1qAdeQAlq/HL6
5iQ2dycTcQLmGsO0UNuyvGYFdGo3NOuvbBmAnqrDG0buT9YSEdcmZY1e+AyGdvIm
M6wP+w5XmWVMTK+uxzh2fllq6P3POVNMz+MYwOiC0E6VjVX2P0Ig93/x37vHKvjE
5z5Ngtgt42+/GSAAX/n3chnKTXkiqZ3wAQnSOJkrti9i/PBHDaF7ycz7pc3GhhBz
8anfpIl4SXBfSCViCjlJnBFev9UK+d3vlG/+kvpn0BIeuXZju8Od6Lb3MAMo1dbQ
Rft/fn2JdAaEKoO6b4QbLgypSjCZ21oECd2/lTR7dNYg/T+fDlEdAoV1n4WXNZ9n
aLsWC1l/W7dh1CWhxSgIv/H0Vlh00N/vztXWpBdOtrGlyonTogd12JqzvKlFoh/H
6Ntoh7YTz/hRFBOc+i4KZ6DymHxA+i3pp7a5Gf45A/ycqVAN8XSmBYtTLBySXBON
n4BJnXVx2WGj9wuFlBZ+A3jOUFzE6LubK8CANjhz7KVAw9EkVT+p2+wmmjvXrKxG
lQz34S6yZMWQNPi+qpYpxDx2pTbhcuRlypKlGHnzGo+TByvZDC6iMaRimoT8sAJT
yBq4Rg/ndaB283f+kqFq2UyIQEtBEmGINspAUZjGHGr675aiO8Bu+3t0wMGvSSar
/RQBHKDlI8CFZvGjmMKbm1+0GkR85w2lEtC30PIuECXHdeqgSVQLdePPFt7hCLIv
ICE1FZKZsKVuLh9Sgv/bY2GXUcIiFTVT5fuD8GnOLvH4iAXYWxhv25SKCIsD22cF
giMXHh12q/kR3jeweSKh9AVrZz3fPXuZwrWSn67iVMMh9mxAqAe4Y5wbeKFSfkIb
BkxFnzKmqSjCtskfiPmhbmyQcBJ4XEEoPPNOb+JewkSKXlfG4defxRPCsvOmENWL
NfM15kvHwVaA0yLHn+pbb53JUBikXdMFQ3SGdUyLuT/iah8Eqsr5lvbj9i6q2UKA
433TwF9Lh0Jlrj7pRsObaD7nBP/DAI5xi/QKaNkVtrMAwwPL4dZSplK2nZhQzT3A
//wIWAALhSAwG636W2NKg4XGD+nemme6R6RWTll7R40GWgENLGSUeNgqKOWNQfCR
RYNkXRRLaZkX+eMIC5/wWydBBvwU24hV6V2Xv4YcyQ0fvcAZ8m8QXbj99GUUC6dW
z4Bu8sZzxPiaj/TnPHAEfZbFkWYJEnG3tFrDetRRhWBetKfm+9jgWtB2i3J7inH5
lLHQq0Tg9bq9C/4b3OAyAdVpMIE+5501GVKHZ1bqfBSAWs3EaeO8w6obdcAkluf2
H5pn7rLUrEmLFplk0IA9vzNwj8YrL0Jo4QMWZhgCGMxFAUNT30XABbUXzN/w9xn5
DlyNeEMtg7tzvxihtCvUtiYynUO+sYHWTKja9DCTnNkgm1n4DrO5xCpB1FbAzASq
824tVLB1HgFVo++1fT+dcAGHaFNFbpiwKsxTDvN+JuBXVn1gjT3Xa8VXZoYZFKn2
PcXC5GQYvHI3CcDxsvmS/O1iycXzKY19uaXWZKB4+j3syqYfdccWTdouYiwN92x5
Tuf2E9EUHsevnigMnqnPtXz06UWK/4z1hxU0yI6oqKxaBLiQwJ1ewu0y5ZQpkeIU
8a2hIsCIPoyho54wYNeuhU9j7Tnm3Feo62O+JyMQP2CSAqSh4qxi7tteoP8zMBwk
Iabxs8reesrTsnCGic/NiMwvLJ2CBgeZ2TLZADDumrfnltzkH7/R1IYvBdLI8jXW
hGX8k2h1D876vqWP7KuUK1XEWDMUtogeDGO7Ueegg0orK6cjq+55dQQbW9VLJWSP
bSEkHGRa32WsCmZ+QSC2E9Ozf5z2DwuhNlwxO7MyA2leCuBKPM4zPNqcRVnk4ggr
Rw8EQNpw062ieqz72a6JPUOSTLeWs+7uspW5WSQ1/kvW/ikWO/rDPTEZPbERlm3S
hNy20poLUshhs8ISekfhjugsmh3UiJN1l04IDCPowQB8+/yFhAdDCFZZJTozoQhu
JowV9NuXM5lZajjoEeRgoQRNHP2BXWsvzs9cg1qKJSX+kjpJ/B37HvuIAsFiVhVM
U3DW2jy7EaCKYcWczUy/S18cxDr7tJRdX2oWfp4Xg7whssQmBdVqpEhvwq9rjcPG
gO5XlRu17UEBcVolxFbCqy+M2Uip05ERknr0jzMuVqpJgQqHjfDkHMCmHt/XumAS
EjoWRbAjW4AalNu+7o476P8QOcxMvejpWikqrsinwX1spa9izKvJK587SircTqr1
QINfdsvQOyTfN20agbATfcIOVzYM7/o6UFulKvHPU6ukI4eSHQ48uw3Rm0u0kYEg
rxYogtxYqmo9nR/AMWydFMqEasPMzlesRnZqoRqQQBTInDRj6asgn9RioqowWr5t
vKOjR6DlCfPYaUt4ALUggdiHr9NU+MRP6eVUDbleEjzNJrDNclcL3zHJmIkx4c7F
fBEG8hAdN9TT7qXyUMo7dziOS4Ga7B0toyHGKDUdiwxHNkr19iy6S4Wnf7IZdTuh
+z1ebvbt2r90UnxWNyV4nY12zz3uDEHY8IaeUye5dAC/97Zb0B98TopPHiB4skyr
sUzgrMgk6eEPwjBvWWeQBVffXQMcOAFPxnMqeqcxGayIj3i1CTJmKhS+nHbwWB3N
clshrRM6F6wV/ekRzOgAk1nq7M3n6TGdXSAjp9dCmcxaqUA6uRpoAAYvjoRbAcUC
gBW77Cl3kq8wKYVCDMTqY4NDi+UGIpb5X7n9Znxfsu3sboF1qlbf7mMWK6Tccp74
Jgc+t1ja1WnyzB4+OvrBi9ZysltWPEPsIHmlUOajPTFqjMzuHzQNDug3KUzBI3as
5ZgKhPHMTnE4ocsV0ZtXp0mbimN/oCUVgvZioR0J+cvK5TayzNv6niMv8f104fkN
HlVXr5qXfCJVjxL0qthmqUVjnPRBSi6PmHcNa9xNZPnuiNNDOs0CV9khhovPNLSd
as97QaNPOk5Ex54p4J5j8V2YjMYBagu+opv4jW1vvlIg82ueurK7Ft8QaH4Xagh4
tuJq5/ao3gL4qMBr4/5+dlH/j6qXG0mZTD94zdDp3kDop76uKHEiY/UI5wIoTjWl
pba4UVBEdfa5A7ctNI3ztSj+ZVyv0//+N59OPVJnaUVTjiAdK8MeOjhPZvx9aTds
VZpQUpYPXlbYZ0LcA/dAQQKvzhQetXkVscFZXXT+8xcCqxXqtOtM4wWZvcoDgUzn
D71cWNpNOZ+ctEc8b7H9wI3zdvT8FnR1IEZ5TlR5o+Bt4koELFiS0iwRjsF3D3dO
noMjxYl4UCnR0TdWepDeS7DL7n8Uv5QSqFRWNZJWYt4bsls6x2yNPCnOgf8gC8Jv
VXQqbkmSbsPtzID3sdWUhQQ/HHRxyW2C15D2Id7iCtBAfXNueIz344i4LSDvsgEd
hUZTTaEKN/GLHmaxzPfnTfUigKLimuGHksy58hB2l9oLt7vTnZIdjjT4jvV7PXpW
MvXSsp/zcCKKx+zZzbGBdhReqy4P4Jbc9OhcAufzc75UiRVwqoQbgmYqfe68CInb
xNBUgXjKKc5pWRY0CvgxsBhID8xChQlwSHLMklw4UzTst2krAm6NgAlF8eriHCRK
5U1vjULUXGpVe2jTkvC9JBe3Gxt7mMjEsLXb7SvPiaxGw+jNWoGtyACpmWVD1x+Q
puCA6ULRqpxuAv7+743eYQ3UPviLK+4Q7DfJsE6TTo0AsE8/K9ng/lP3oLpDCWoz
q91oOSKAT5495zp2EI56/VgUZxvUbpk6s60prw6PHbg8PXEHa3CzZBF36dqPhLhi
r7opAcMMP0u++OwXKwPhX4OtGPe6iZW4a0LgoZH+46polMxkZGdb8TfKFKXYviBk
siV7+PyWu6ppvITCGxStT/I3wpPskjdaMTz/9hO4mOzAbHkRG1bCmh1zf2ogSc4L
vSnnPuDEOKVEOHrUAHlEcMuhF6g24BVsh4WevemKpEB2NQDIY/Q4RhBjZY4uk2ot
om2Zs7FkFDVI8BlfkmsQRgsAmw7s1otAM4q/c01uyHnUyLuzrAJhRbMEnSu6yqW6
C9qra7YP7tS0cNJQWij7T/x0Sg9Mqxz81cRU4Kw3Cqt+Orr+CW90jpluPWjLgHXG
8kyMS50f0bxyWc9Qof+SkaWaiqLxlLkr4EmjB4HiEklunynXmiBfn/DtK7ALVcyR
tdthe3nfEXa5YJsi/K8iOgUt7OU9xYLl5skWFHNxgP32IiIlsg9tJcMUrYee2ccd
k9lti92oQE/hNdUm7BDu37hYs9zWID8JkC41PHt3BiMy8/b6H7mz5XdD7cBJaSpz
wWaJzYD3IvqWx/tdJd413JEVKSsqMI2OXvqMaBit8Er09KutLIMYdmvll1wf6twJ
RSgkYxlvStOzqjePpDmL3kTurHl7rXxxEgpQWfFUH1DDda7xYbti5oVL6sjxdzuv
eQYEoHqzrjb2lBaRoBxXfqWvbGksifV99rzSi1IyTDc9A5gSSqkSnfO4q/QAo1ag
ET5drytbrcSF1Uv3uxaqULfiuD2LqPOXxPLP0RpT6XR9p3nLySWZ8m5W+pRqRyD5
bC1qcWKtrx6nygcJtpVEqUm3cSJsuvprOQZs5bW0ul0iK1+R+lKaFVUSc3R0+pVP
ef07Kr5JW/3SEQHJIx1rDD1HqKOYUhuDpERgR0ujzI8m9DIlV/Hkslxf5rBMMfg8
GPNBmcwY0j+0HOP+SdyBsZ7rNNRjuG8lH0xU0Y/2E8l4yp80Cp9bpmE/bflGgdaV
VPXiSlh/e5rBHPkOQERMRTsvNeymsD/iaLGyBrc7ObqT0vo6PLAp83aCwZzGaWXu
d4Lyt2hPPP9RtdbHQCE1QJhfPDAKckJIS9nK9g5nAszwLuSIqRiA/9SN2W+YV5Cc
q2LrK/z5p86iw01EEIlTyX7Y9KXV7xcJw5dMhqFZyn9Dwi0IhjV/FjFx2HjE+ZKX
ULWEkGir46GTmcKmIKHa28kMixZwcnidRVV94uIpT1Xq8lm8fxbt/c9ioKGhEAUd
aeTJzwSEmfFI8R0DwZOXP/eVXSqorPIfQ/zsLj9b059wG6loPYtHhh3EUo9ICka0
5sqepY0/amOLIpiHC/xPMlPuWpi5BplChzQLYHYrL8Ir0WuEX/Rw/X9+fO1nhmfX
NM6chec2Ov4N7Izw1G105zKGWnMf/uRbSNV1/dyBiDitiaVjX1eDtIV/LMF+OAN8
SdWH+wiqTSvD0wsDM23dNxeHzyKlRDxzp60KtXDFCrmCu8SGaSgjbAu3L+UOx3v1
bHg8uvS7yRLgWLW6Ks0EtMsfjpxSuvckJCcg3wwYCTEYfB3jhAoI94AGyeRRLOWX
zTgXmlMN7iGwGcJFzu/wN+tngk3+zYuUNNeTVlI3wMcV48CLxY1ohmv1MeugI6ny
pxjo6K/cxmgwKJbPAu8lAafEy0l4L48ftfAaCY6oTevpyVqm1LxNpXVlRtChSVW+
xi96iclwGWlsbvdXgDpANFF4CMxKYIzVAkzgVVxHt2WV+6HMMCG02ryq2UqTEf6Q
xZaZBm4rnQn9jzvtfmrKCNduy7WBJme22jMRDm9DfLRhtNzaPHuQhdAG/bIOCkdP
BPrqtoIKF3/jHk7KnTEOtww7g9u5dCuYuP+1mXQQOiKrM7rhxXN8AZpdtphSEsQg
P2TIh5TaWS4nyn/jnfT0fy/yv4RZ0gM6Lhr/0uoc34TAqXySOWZ8zadrE+0Vufak
sJd2IUGUHJobTuZOg3z5Gqu1hCo5deKiUK45G1KG0yDVj8nhJff+knC91a/a73VY
eMr2EnCJMpxcfZI1wwZRtN/AIKoSIUF8URbiCqjvccHEwt7niBp38g3E6iTF7JER
y33UCLWd9G9IjMA7eMdvHpHEHcl8W8XbQ5AdKbFHvpcLdgTKLBc3ul3UNNrY+Xw6
wplY+85zDLWZvmsn2kuYHqekekphOYRawSmyfZVyJcoInHLlduRSObnRU8xRIIPR
5A/fqaXQ/ekVTbeKQtZlEvQh/MOLlgh7hFhvuVPv2+nriaPr0Z2Z6xP2BnAPLyca
yTHLqsJADPQs4XBuZFEqiI95GprlwtZNwxrJ36XHGmtGmm3t1MRhSz7HT73XzNCL
3/RvER+ZKN09T1croqkd04oMVl6R9aWtSxAEwFbSUyEvbXAg55vewZLcIyxZo6uD
9hDrj6W645rlbnrgO3mAteUFvcL79pfL60RWZ8cc1VY7YJZYv7N1vXn4S06kwW6P
Etq3Tfvo8nfv+BYxmXqOn7CTHqfSBjNtNf36CGlxjlMAnESgLISHK9UVDqeF+F08
y7J1ufz3TqUB7q9X3xtyXIcsY3zSZXPWhdR+eYcRFECaM8GHdcpI72cRLhHTPFOo
ZtkKCbrNnC/NXHWqiqsvyWvmO+jj8gpJ2sLroXEAnxBn5Hst79PvRoU3cG1qOueT
tyJdQnz7AE4r6FkkhnjKZ5XCYr0ZUIOfoD5Kuj1HjQdNB7pF591eqqmLCcUeKNhf
p+LFKVvno7wv6y2iEjOFCEW/HSwoUunkTPXePxqtAvXYUfnjlpWbjdXrp89ea70B
hVGrahPXYgWiv3AdJ9DWZrizYagVH3WoB7VqkFzWQO2qXp9p0wGgnjjE8ucB6CIp
R4GJDOWJKL+XjiiLl1OY/F85NGA16/AbF7SFbtYsJnM8sqs8kKyWesqBC39z1DcI
jYJGXwP3AjjRG3Zn0A70pjiE0wJdxWHwIM52XSVTNzMm6sz7tCo8XJjQOo6UaeJx
ePMsMGrDlm7XAgt4z83DTjz2d4YtIuRgYGW8tnSVdv7ZEB+8XWMTJ8GxKKLwarwD
zgru/U+TQXgkvG23SUNWpVjzE5XKXsyTUTw/sAiZNGcXx0/097vEzYfSnUsHJSgs
G+QIH5BsXkEcB4ubOCVAUV550RSPeI84LSQ9LMG2mq73BqbFobkifPKCozNZiFUc
lZGADFu9LhA+zJRrWL2hTur7IoeNsh5Ie5AXe0WHo5b6hKsbEEtHJC46ITjhNfsv
ItHCBZYYAphjL/wr9sZ3uB5KtS9uAG4axKOJW/nbx2P5lU5s2Ep+I55epmQSR2qa
dscD/VwjYqHJJ7IqnuNj3WXL/1M2szM1m5v/y0pN2EK07mjUsClFAtp/2+2hHUo9
gciB4ZbzjibpnmLHYKCP+kx4H3kJVIo43h8jRdX1DUFjrPW6WXqzuLsULXEI8urn
hJ0bAt9CPYiQ8pR1SInKF9/RvYDc1ptr3sITv8LS76+OqyfsmOMws6X7xUEX105M
BsCdsgg4VSj7FWBcXQgbuB9lCbBZA5g6UkyXDgTsJTY3UxlgCQ/nL8xxbQd+PzUh
WlZh1ynxp3A40rZ0hso2Fr/GXBHKLkO51s5E3XlQN1wLiI3CvtV04MSJkLXv4QZP
Q6INYH5ZRvjzqxME4kCnsaBT7yY/RAadwEuT5lZPM1t7FFeS4I8/cGPMJ59X41LF
GG2FqHzrAWY8h/7bWvV2VEMS1jgfOZqnDYnTuqMWqy/VVoQst1xjmrsRL0TvK0d3
QFKQZcrUf/FSMKRH4sdbtQpUimtstCSh3dYZNx0IEPw0I49du4X161uBRfekDaWL
JNA6zVuekViuA42wlZRFAhcEKQ/SvPZxGdjRO7vQxhbeCADhV4Gg1hqrUJxE4dOL
KHe8ugZjnYb9puYti+iSGMK/nxuIFlCHaxfmKImAnlRuuTTRAuluNYZk9gYMc4g2
OTeEJ0+oK3Y1Qs2Q0MUe23emnq7yTEuNAND6tudO+5lZy2chdLXkx3WUlBhEdhbg
OUaGm+j+D9X8DPLb3e4gHS1BN4gyIjoG9rf/M33qeu+cZrCYShNrEVxYgFepNiyX
n8kRSWq+lPzTA2KUGpqicSXb9Zga+kBPJwzisuf63VPz53B1e+ZFeWrwvVXTHsN9
isEhR4y6LZ1PV172/p1Yn3WzHxfAfAZxYMI4uG0zpUEiFtN4I7ai5ROTqhjUjFmb
oH+PZlxP0IPPwEd8dNchZUVcSUB8oke6GRykGHP+UNUdi9LZeJ+wpDWpyn2PQgZq
C+Fcg31dnECwy0BgbpnULUKpSkJ2FnLkdO4qRM1PABb4q3QR0PSOuVhTW04QWzLL
4jgDRviPv9XjN51Jm0RwEsZu1X++hMuul5CgnrG3pxmUlq6O6HIFanax6//cfZc7
E5hhy6P3wde17dVlsANEIYVgIqXmW1/q0DUNXk5KrvTejq5Ob7r6jv/CFs/I6t1q
KQsSu7H+x5rJCAanGrzUrROLUrIHVu8/+XE7B0SJIQM5RJX5Xc9grG/rQp6+s8JX
k7JgNvUqTtreqE+qTYnTZEXdA8gbscDyo47zUDgvds8hL+K8nRdv3+Xy6W50B4BT
gHgVWBcoUtxXTBmRAQcDQZeYAOfdnQDxE3wsjQqHsvlstWANMD/pwORytGX41mvC
kfFMyY+V21Cn+L62DwumToVWwWWlgQWVt614kvT/bFFqiYr3uz1A/NUFUqwktYvw
cmfez+hzavwz1EXIX7ROoKJhJ6GqOUwRIGgS44EIbwBx4LaLzfK5Tr9NClnPsFwC
aOZE3oUHmou5OnNvD/HAhwMY/JMhzoyOkQfY7HuMAWRgvZNwUif6XlfaDEBHk7yU
yTqKMmpN5x+43GVr579mVWak3XhIjTwhJQm2jETzJnwxyQe5YkPcCtnPnun6DrLV
XCIlCEqhur0ddTXhSjH2mPkGIhN016HImCO/5XmBuf3XP/A7+fYqYheVrQkv7MK/
c4kFmKYKMJkUDt+RsUUqAfHTNPmKjZ83HaOW3dIhZT6jx0zrWfNBNC/7KvQbs6Hu
helE5LYTdzFZJi39xmA+ARHAwrQcBDkB/WK0GiCMJTc1L3+i3VR4MEREZed1cU9j
xylydaVcQoJ8R5TkRa3+vdzysgYh7prDJhohtbU93qBTXDEJtXdpn1Tn/RuNiQFy
C4SfUNo5Vv7AncY3eghaqPkKz9/A5EpakgB5Yq2IWhA200aJd55FjzcfTYmG20FO
4FclgqJGjUbwOKDybNnWF8zSeHvE5Ss8y4wXE3y/5+6ioE8fFhOTAtoogw5SsaaN
asAPu+/eFqXubr/kK68pmMuyc0oCBZ6fmHsAsvMbrAAvmyJd9OtppOa6cg9PZ5D7
+0D+5fAz3nB3ty9KOKfhUh2C0usEbXDaLoEW/TV0fN+5AuxPoEgXrsgibdemfGY2
uZ3WHOGjbCWoNjb4iB3p7CM16tavnokF26A7i5lS0WO5ixMN/MVe/huRFxvDYJbu
nMMmUKkQwjXauyV12UPzmePw8dj5Bdb3CGgYqHAwwx2f7BEqLJ4QEMHxOdU2Dhaj
v/lefFbGKoCzPxKxLVzqhQrKt8DCqUZnlhvFYN4feuVH0Xy79Ao09hX/z3Jk9sIF
jKxgiLH69ujcpxG3VpXAd9s9BNAvfmCeH6KYMXSl3wtXdJ7L+VEmHRPqfwATj34L
T0wURwqJKzQoMdA09OH/wRWdteMu73yjAdn+Am0aSRsHOWb+3yCh/iycZ9p9L9/0
gyKjyjO6ZAjngoCBkxDog3SIlGVBBGEr1WgVCprsXzMQBEs3xR1xj2TkmXWttEn4
MMl4fuspA3i36HWev5RktzPuhOWnWF6mwcCKLGjRroc7tdIm+cUGh5K3aFe1Difc
qIW7mkUazHn4KxCpkecS1hPnZ+cDpRxif+16d2YGqPZaSAVUyjS3w4VbFOb4F5az
USn6g4cxXu4UtujnMUD/y9n813rp5GUjb9QMUWIP4aKuA+4iefbzE3ixb5iioLX4
UNkJV/EqWanR1w9uCrKv0JqtXnWPPyW3s1cTwQHpUisxvPlrPWzt/U2HVtqm9TVn
w4A4sw99fNnfJUKyMHtdSRaggb7c3u8IscFnlspis/j0jdGh5VvQVd6YVliGRmJa
1HeWRqurqYWvaSWA+LaHKurHqzGs6pCv7AIfDE7+1VIajTT9FPo1k8rKSWFXeiSF
s1dIkIsxHiKidLnt1dILEGMp26GHRvnMHgOIT9rZwdP0qlNJHGHvYfu0u0a5t1UK
x2mc+D9wbxHk8wU7uvDj+Q842a4FYt2hEa6fzMLaQSeVkmeGrQcgFEVMkAWAcIIT
4/L1GAJffOED2pRSjwIM9mDz9hf4jpNj48RR8Pkg2eIs4pfCvS/Vd/4/iegNjQu8
LAYFYzV5zrjKJYO49su3EXpcjflNt+hvhLmJe/CCevGiOdILHHaFgHGNCCRERJhM
mXzjZ9F4L10AD8uTMmH5jQo1svlU6A4lnS9W1Cu3AFv/VYuz3xQBQ6mdX8lfig9A
ZPOxAzGiw/PL19e8MZRgg9qyrXH2CNq2ypD3I7fpDqiAL71/wBBxHtjwS0S87d+A
kJ0ZWk1WnYkfDmU1RMxsWAF0GjEH0v14hy/7vPOq8SOciseTLRTHTdNhmXUUsQMY
t1aR/MmldSambdRberVHB/f7uRVOwVfVSvY/RXoyzNdhUxepHOxxYOi3kxNCiVP/
WZTLkhqx+GeBX17m64LxDODuvH7iQn/5zyZwCVnKsr1xZy43fHCHtJTPk4o/GelP
0JNA/q3vQ4RggZW94AUrm8ujQpN9akqKnyKoNHGE0PfeeH6reMNslchNiirkfzSB
bmtSChRLJbG+QPD/Sok1vuqkE6u87VjXXrlKebgmiA/a0xCCIjJwjAr0RTAes9u1
To5No6FMTYS5n+q32XlAmLOzojBhf+UC7GmYHrBYOqOk9uR7X6q3AkEqcRSZHp0U
cbvLeKVoEjw99nMfWqliJnYgu8qNq513c+y0GDft3/l6R0Ia9EIjn/l38+WfZuW/
gcu0U05MujipIVhT5nzx7LFRLsRZ5ZKvKkeEEoVUtqUVBSvWs6TOv6o9oJrPGHER
B5vd97giq+UVgECsAdRsBg7wPJQS5vQ61Dj6rW8Nm/VGWWdjUrk/02oytH7QUyuV
4r6nI6NgTBETgLc9H+bjTjIiYfAHfH6kesVCQAFatRRFc9Ewshr1BqYtlTkOO/TC
nA1P8qhiN7O3OUdelRDn8rqJWY6a9+bGfVDZhDcieZN/DkIQodCk6qTOW1UMp0xt
I02QCXZH5gbFbm7wp8RPDBJpWW5E3ChHosF/EEbL1YwNzJChrdwf9fqM5oGWBn4U
N0HN7O7JNb83cP2G4rPsusrhJXyXu+ZVXZNkFe2G0Vx3PWLWLoTXcqa7b94hRdch
U0yxOoN9+KoYFVC7n6qPEM+IcJefm9ghXqTE+2t42bS57y57DHTHHugx+Y06q7Pe
a8xK4zSa1mZCaRehAduGIWcmBW32kSuIyjFGsHnBSFg+VALxrs3PyBBdVkDjqNu5
FxL+UM9l3B022G8DVWU3wbXvY07At9HimcZ4ysZum35M2IAwxFc0L77hn8Memke4
4Z8FXfopi68y8I4a0mI93V+WZh7dVggdPVugz7sQF8gIO0ojik+xcXK7Z1FWOsOn
xt9fmuof5Tgvu8677UzVybzglEARwOC9c9TTYbqX1Z04v1n4XUWIrNn0xfKgN1nX
6e89fKUCBKN/yYFn/slAyvm83FmqTotBmxtZWok65IIlK0epc8kUY4SCu3/DW06E
TgsbXZlbpBVP73CXDjU7aRkCW4dWzm8OI5qtNYksKNBodaBLvOpwtQbcJEaiKWzo
unWbfZTIEYrahiG5eGY9fW07d7IZH2R7DInERNdaqje1DXmqiLQkaONwGowr1aN3
at0OhJegUPD6yvNVSZnsePsmZy/R5Rkc7Hz0I2Ut2IHIJFORo9ANcC9HgAsb2S8E
AaCSeKd6JRxPgIXUlalR6cFDDCsi8Ts96f0P/u6nzqFFXoR5oAIkt7wuWMO2kFb8
7F5ueF3+qyublY44PlES70zs/JJTaJr8LPhJmLAaQvaFfEErIHzTzpgUA/7f6XnL
rnsVIKKDzUMmmTmJv5AEWGtRIlayrgMPgoKwWfIKbu7JGJGe0RJUyGQMVvGxJrpg
nKRmj9t90P5FF1DCqIbF4yo6dFaLbLuFmvyewOCNYlpx7c9bDgfQdgI7mJXGaPyW
Hw5hxeFDvHDesbHtMi5rNMHAsM7+gQCKIMeGkrndN1tnjG4qViB53Az9yK24aXWB
mBd1Fa3aapcT55WjqPfPPyTbHv4RXTFKb6PhoUo4aHZixBdGAaRX9PQz7Bvezwxd
OcBslZlAvdGFaEYw/AzICDQynDr2O56Mndd1HovpvIhp06/eW9z9RZzT98I/3Aiu
LyOVkUwMHCDBQAPTYpyb1u42ZfXJTBmnUViNPFCIOfHngAh8rLRNsqLx8wzzc7UB
rQDMIIlMXu+J5jAZ6qt+hXh4LtBSZbgQYEGzwdn5dGoIX7w0DZONImcaqNLtdW6L
jOLtSeLCJR54lQdB5OY5/vRvWTXNjykoDGx6+3Fj9gyTFY4j+gmE4UHFRSfufus/
ydNcuiKObe+1RiMyTf7zbrZM04HasGTbm8An523s7TDp6X32KN95sOC8G54xNgEQ
245dulaAQKyekVCiDKRmADhi1E31awTfqOv1SYZQYcWkBd1PRABv0qO8Qe/rRYNA
LCF4s9yn7ShuO5LJ7nJemp+RBMkCoFZzbfCpqaT09MX/g1j5ZcPzxGbLq+JJpVJI
+9H2yqOlpvxqDGXLcaLD/zKpHQ7mlxVIZSvKOEKBX2iuub5koGEWTv4KzsLNt+oq
d+8/UNfVrLultpjRXVR9PcRg2lJcVJRRPkdiJSyW0YViASTgOsltprgiRc7m/jp9
X7GajD5GKJ9iLAHZCMm69OcnE+NvGjKoXswSbS5F0h4jBlQr+25GEq0CuM/DBvRr
bQ/VWwJzfZV7GfqtWtP6R2sEmbNxeec2hCK22ozegyF1G+0I5+Dx3+xJNRqIxPvh
e8sHX54rUQPPFP1eyecktDFdTUNKDbCIiIjeg4byHLYWt6bizbVtf+AzOtmCZbQU
6uiNcNlmkCPmtXN08Nxn2S7b6XbjwE0FYewv5TO60aL4uZWo3s0yzzKT4j4UqyPu
jx+xVZBklw/qq69dkLLvJh+zQSQWSrLeSMf6xChRlr7I3B+utNycrzo42BDheMXI
jQA/BbJZrVeBepQZ+yN4pr6TrrpxaSnKkwnLRYp2YZOqNE4pueXoCgI76KCH/ADL
txSp9DydpREp/rw05lKKb09OuLa1MVALIdpEcCzGWL0dUjGSMbMiun76kfrUzlr9
BcUmJQ8vicbkleMBaXH5cSiAvzwMfv0vnkghkokJjY6fItuqyIkqloIdWscU01uy
SdHynXjwLJru5dcBWVxdNsA739juv9yIcEqDfy34gm7A2PW8itWXa24guJ6O91sj
y+j4z5nWTf64zG3UQ3YpGu2ohE7XCTcZad5qWQf3RcEDd0vUbkGCwecFwGUpj69K
W+d/3QTATm7H0L0YaM8lQHvmzrON/oPGJE/+e7AWa5sM5M9HI1pvOJvfNhn2An/t
Pes7Xg4LJslxXy+mX4IlkoZE22hhLvkghvMrh1JqhmHT4t0HmyNwbB3TPV13EJ2w
Wtmc7Y7TJ6BR2eix6o0GAQl2uZKrZPqhXkK/iSY+e8c9Bano48Nu74xxMarhnqjG
nUUd4ozRH7n0WHfxRfAAxLcQip7jRW4XTWDfxitbPiXDM5IUZI5SjiisnaM9HC5g
WSYVqBg99yP/Go4Pi9whjF/PYEWh4GR8WF1JVLhc5TmpeSMvG8F9dh+uIzyrPzEQ
LmXsw9b/EzFL9B6rlXlso7mcyOrStlVxW57rheqAWgbSvo/x7HVuRx0DlyTo/8Fu
6EiDVTGKSKh9RcseaubZE/GnKBuVko1tkLSUctFIOQmzpDtbdQ4x43+nikc4+98c
rShmUmO4k52YA3Fl+3u+EGFGfgIXJSPsB/FyRuZIRLUQkTvXaT4w+WCScS+03y+N
enCq4Rq40JbsfVsoIySRKvRxaXn4vqF68ZRlQEMoGf2t/1RvrcWctvdXeVa9diau
8UJcIFmbBl7Gbn67r/zkN4i7vpWepHLgSLS7wD1jA11tfH+zW/C3yl/7eeir7iW8
qlpTkcM6dDVt6x9ePeGnDzUjCCQ5NGHXO4VFcK3crRKBqHkTQ96kRXAIZS8P0TNP
n8CBKx8Dxsqan/nrtRD67S4J5B200BAxhHHgzhAE12Z7oCUuzumTq5CxSb5xit4N
y2X4Nt4K771SSHXy5fO58O0A6CtoBdFvUtBhuhupUueZDEp6zkI5Wb3ipWudbZPb
RkXYAi6Qec9VbOPdM2JpkgqHYyPilJ5OQUhfjmvN+XUgwfucw/DCHmdYfFv5vkSI
qMSL9JvbiHXBi4ymJaEuFJsd2RcD0YVJO4GPN/61mIisaFrBK6QYTarDxPrh5+Mn
cDr4/eKxJ1HtLzHAR/6Jhfciy6kNLVsaJXifEfoptTWc5Ap0y0Hbpw247CPF3ugB
BLQZIoMNhCa77qcwuD/9XERHSTkzi+MbBcDcUmZb0CP2EdmYZGpEwoT8ZzYo5V/V
BXp2manyXPfl5w94QhTz5qvACFmrtFi6C5scfjyyFAXnZZPokwDhCpYIpiYRd7wu
HNbgzfdRCdC4IowLXWDXz0CX5mUenq3wmXEWf9xk3CagGZ89QYHJRq06Q4NBkpHL
/6v5dM1DkQlh9l9u756jGaFF4RaNBOfvYJ2W1HXms5f2E+T7VUvNukhtCL8JYmom
FN9ZZ1evUJ7Rizk4LcB4JJiyQfBSYEoJKY2nfkGdoeS8i6cc5Ff809brAT9cd/gw
urgbecSKe6xSt/m+0nm9aqz1cS8+gQWN+MwAQSSYyg9aRuD/Nzdwys+CxlUQSkYv
cRYGhJqHCHTkjWqEbvgUGKtPSf51Xs+vNu52Nd/MZkeli0wokogm8do2DfuKmGLc
bMzGWTEyMrI7xOj9NJqwMviv3IAioDT5nJcJrcitSsWF7izG/VQRRIxcQHvLsKw1
OUGPymGFRgpR9/E35fKvyhEwTuqtvP/CdFq4p8VlWBQRd60hQfbkEx0ByCJvvqNz
sd/79dPU6+4o3ho8a6c0zlAhvsvTGGYVBam1C/Ra5r1eAKiVxFOMG5R/tnv/d+tB
4MNijenUqkJ9uBp7WLDNYtZVpd5zzoO4u0Vp+vZVIImOTjN4iV7I/UdcqU8ZJz9T
kOkFktGlAdglyh0mPLEN7qRAw5vmYGCuRFABIT/2LO7PD4GdKAnK/IJ/5GBLtlq7
sAMTE8/eNvxsPU2r5oEuu3MpYImlRyLFq46Unq/d2+wwqyk3k7FexRQhVnEyRQrv
XTBYDGnu2TUNaiEB6nGJJx4krB6A9/jvkLEu3e+KvqkgQqQlNwOVZnJz7eS3FY3L
cl9LrxtV3fl5IqVz0g/QbbQzm5OBXKNCYUdHax0t2FcjpwrBr5vVw7HE8ek3h3ul
1jsqHgXtS5BIW1f8JhLFriwT4eMHwmcrDVz6vEbPYSYVAtiqGRM3IGrxFcpounLn
/6uDV6igshkh4BJChQGcNoEcgRRDuiyvUFU/nyYXhSDJhd5jQRkRInDhhaoMAuqu
hJb6GLLMjyyXpzLIBkJPsmc5rdkIwV5mDlhHeVrnbmeldirprWRul1rRr6rvVj81
LUDFxHYK5RxQ2A+cSrApKUxzTcO4myacXWwch1kHReERcej+7rOfHh8gVeeWE9NG
hcxUs9rjpEUNvfYsaUZT0kfDrOMhhG+UfTPr/JB0TOtZkNwpf83kvByx2M2dUB2k
HY1IYoGNIiSBJ73GmfAbEnyN4k06DwvlZxSxjKyXnZskhWbosKK0X42x8B3QUqtR
Q6PFF7/p7oDkxO3oQtCTc33+dxZ5FlEOKFUDUy2SSPmmsaSKiUSqqF7w0XLByjEI
K+NNKjcFX2b2q7G9dKyv511slpbI9PTFgwrtfUWIERAqDWG/95pJTXwHwJkGv7q0
DFANd8njBgvXTNdDqbnneIDdpB9qgACxmPTnDid81jrdTu0AGIuJGE/kh+t8rpvX
tq5o4/AC/oIvsZhOt/tTcZ7ar7X2C8PKyTvUEWuxFgsZejwvr1EHp9a/fgklmSsc
kl/+OX0tH61zHdqEHqdWhCzinK15uy9fdfsP+IK+7hrK8G6Y06WdaaQxX6w9TvTC
Xutris/0Quh1U/iY+i+ygMq1UGDtqIyqbRq0tpH9PSru5is7K8VE4OceLl7prtnZ
+TLS0/hr5KJAs4tQzfLJctk5a+mp/9ggox+luaSbtMW/laBzy2oFjbKL/0CVJELT
vPnpMlfqX5JDJ5EHt1LCBrXgUnSBXJdotC57eBu8yyJOUUbtcFw+ni/Y3iK4a00D
CJ6ct/cKhmaZxrmu7Ax2J5MR1B1TLwlfUyshgqrke4Mv+IQyUX5lyjL6FbzG+lKJ
CQHhONwhYn84QVaMhIbD09FdQb6/c5eWogVAYj+KvMhoRc5KdoAcFC3COoJOqK09
aeJwaTRnjP3NpTw4eWKg/cqkotPtXL9/+GICv64PVzrKKpU5e32jT0Hfgbwlz6RN
8iojj+zLVeAcnGT1CNPItWjeiXGo+fr80u8Jhi6lcVAfGVyOKDv0waKwAMlbIu84
cW0fVPdENbgqxY05Y4SnWyPBFpMV9WH5Q2Q1n6zLAojcsqqmEai2I0GpB9PQEdzP
lQFyb89MlnprdYMDGidZGtduT9urD9JxV+NXMxzU8CejWqrGtg/mBmB2RMEQzSGk
esN63q+DVYGS8xUwZqwAYoZFW3+l7tPQfOLbdTgXWQfof1IicjWAKF5hnQqnXn8A
Hu6McLQBAeEINZOgP1H/V7jOsGUo3Phi8LhSoBUFyKjekj1OAbjR2SW+QrQC3FLG
nY08iv1JhAwKcAaq7lF79bl1zFLtHTpapu1tDux35q/iIUlxHtz+0Y/Z+q/9ztv7
4HbGd4AXfP6er1PIaUj06Gy32W6vAM9MmRffplPa+rMPbey3XH4Xm3k3U+s+BxwD
rmv+iF3m4w7x7H2sIeiMvcw1xb1Tcsw/vHREJRUF+h+JkxfE1s0OYz+yL1YwiW1i
3mjw5uIJ8VvRYlDIk3EviwyPG4UYQGA5JZThuIOs+mSw5XsKdbHdRZfGUHsHyjp3
GrzNaDt3UiU9k+nRMNCPl1HIAie92B0ABt0CQbKs+CaB2T3tCk8eyzzgnTLvc824
JmlhS4/DeJAyq7MJnrn9RP4mogwX55cbxeaOd1QRu0y4B2lOnRNTG+weRaL3ky5l
uoIYFCd2lj2MiaCAai1SVFoITl045OKbUIU5YpwhltcLJRld+Ys62GTMR7nacJ+B
DKRQNFodGBsC63X6Kraih0WCVNz5GRBNk8WHG9vCaeZk5A/IKzsvAO8EzugH2pmP
yfbxOxIk3Vfv0ka0Kl0uWIuqCmJ3zypRgy5zjHoEUmiqtPlYURlsVbMQ7xba9glP
awH5r5o52phyVw5IHMs9HL8Yr0Xmh+nFbB+02ZVRYSyMTU7Pmiqmn40a/403S4EK
iPsoej4R3hcyA+fvUTwI7YLjXH/PHsHQeMAItjng/zS6eOSUyiHFZ2jBWAMb3VIw
3BQhReGRChwQAW2CdqHRO6CzQ3tSBzTA8sGwNcOfs9D42b8/bmzRBFX86pEtDJ+p
PQgSrdOFTyXLmrA+cIa7IvKa65ev0moFyYViFh2fMoFlobiVimdtvyYOfxRENrSH
/vQ8apnPLGnji8iYHpI75S34yNem253tA1SAdIT2rkLQmUMIFZeu/wyH7Qn5yr4v
gs0T8+GHkienNLcpLX0B/vWgE+o1G/JVCIcezNTOL5h868rWCWdPvRD4R00hu5tE
pA5P9x69/JOopjaiK+o0YHjOFsEQgt0XPSSt1i9+67S8TJY+VqCXHj0+rTGLT6Ut
wQrUO9xjSx+Bq6HsNRMP5M/P4lbX8jBulF+afAFvBH3N6sVFrKm11Otn9dI9zG18
+6UhI0ay2ISIx0xahoFelHXg7hoNixw852fj7+CKN8M0OrLME4SlX2pppGX16nU6
VR5qN4Ms6P9AKZG8v310LhNDmjFR6raEy3XfiQAKRprVNzCqtKeR8EZyRR0mfb/q
lfx/UDCZ+AN1GNgMGf/HV6WZ8OwqQsx1MRY6EDAj1G8w9hGYvDF1qygusQXDXIZH
rz/LpPNw4pM6IyZFqXHFWaiznaEOLkfIsL/WmIPEeDRbSI0yWgJ7jhvQwouwJHiL
Ur/f/wAxdiGU/sfgn5ji93vvWSzmC3lGpRcKK5gY1nPi9yTEpDSSuYXq7QFegrMO
lt2ZZneIVCJ88mhXBVcS37akzbZrK8LFa5ZsIgGRW4Hw4e4noRj1V1V/+qSfixge
tu79PKIOViId+k+iWC4X5uAVbmp0kzOQSsLjZy+AGEcMNbdBECi8SiUacggut0XI
X3s+Ka9H8pDf0QhGMWBx862j1v5Q11wkbl2iYMnKCmzB2Bj2ToT9FGcODbKBVKJ/
5/OVYowEu3LYpMOMgUxfTIg844rjOY5AD58dT7eXzMADgBF5U7GkqCeebcIukHDb
m3QH9MGj1qbSI0eDZMeXxS/MwnZarT4Hpiz1HkVSrFY5hn8vkIfM1AzCHwXromWj
6ajKZWJCOeSDiqKQOWWJ7nrO7M4BJyrx9Rz1zZmR4IbsAJ/t+fQIDo7KybHZ1vVT
5BuhrU78211/1Dceqha2AGaBE1BApwQQaD+8B+WYeRGGBmdgOLXuLD3MTDZmG37M
w6VA2mN9mThsGfyHnjh5wVsXH31xOXNXaeSY6C57wX52gdB1MohnvkUcjPdOTE55
R3U+bUP9Zt5Hv0pFAZb1C5r0A7Z8TSj73ioYzYesx8TDRNsJooSWCAc4/8gB2r+/
msMlUEOcnN4K1xNAE8H6z/SCcpSJiZoF1pHTrmNg7bIDPddJ23yMPAaZmI4Klvjw
/FgX2/53ScUgoAxvzfonVA2vkaBimu8gyHZG53a9c2eSOCv4KBcvh/AtPP1+hfYd
8aaokuodkJczmJmsTiInWiHvW7pvv0Ho5Gq3gvsaVkMU0kkCuHZt+/443f6s2MJy
sUMXl2G/myPbWmuZHwVd/mLzVL94gF5xbdsu0AoI5qCNyWUvnGAqiBL9Cfu24Rm5
6qjPrTfSsM5OS9i3zS6el7zUaGdFvHqOX1EsTulXPizRfXOGpeFi/jeSmt7D77Xn
gc6UFd5G8DweMqNLCJeNQxQK8zZVdWzwDxlg23eVF5ip0hlUxjWnjS+s5PK7cC4R
Ld/bFW6LsjEVgxgb82GjNwvAtD6H1fyL8LjmghTMk9zQCd1O9HM6BXkOOVGlZxR1
rlVPe/xo6bqTSwxswjKGkal5Zf8zQ0SfvCvca3US68K6rt8oU5Fn1IG/aJbOOmzA
lkTg5gZMKvz9aHiTy8qp/+5XR7Gb1jHK8HjrBEqvn/ivqI7MMzNQ1ZH6xMKUMVhS
wE5JHBZnnADUsVbTuB+g88Hu1Vt+ez/7sn9Im7ES8YLsaHZ7TT8X0waO+aRCtqBT
C9f0xv/DWMdexHnStyzyhTM/NyYJ8IFlpPuKcgi3EtYWOzfEqwnyl4Zb64w4ypj3
UP12ZUKjWuWt917TvxPqJhALTT6v96upt73AFbzfQCYSFyU3XCOADHvq9eP6zA9w
qLk36SwpIIBvP99kX4yTKQO/41DZ8pHL0Aybi9KQNYI3OrldgElEClz5E1PPUKYR
3v3N/rvPwvdak1hfpMp6y0vo9tFTKBl2xKPJCBpteO0E172+yjMOL5uUFuad5yXF
t/nxpcl2SnUlmkldeB6oE/9+ZxvJw0K89de8eqiv6SxZU6gR+TA8zgCmtf4/JKfH
I43C+zBLraDJX4YirolO+bYHfsCAsxADIRFnphq75yDxnfTGMscphnFCPEA5copc
zWvvvpx5P43/3RwwuhSM93Qu33GcLOCkEmDk98OBKtPkzFeI8CLclhKQLAoAwLih
9hBvCqtzqIDiqvJaC5WsqeEkBwYJy5N1a/emFUm3BYx9bzswWh6g9Tpp/XZ5bj1S
guypTFjP8g3bt2gW12lxaJt15c3oUmH6JSAxXpFuitYXPuqEOtN6RpipcnQ+lkQF
/J36+8/gWFTN94RE/Ca5uDZFQdQyAVfqrAdTRw4Mp3rIn4Z5uo8ucr+Z7V7pXXPS
7ds8cZ1lnHrrHD5Bz8IycZrDff8uk3/engo5hApFzyWuBUoD/8wi1IrMENzNj+uD
XxgEhZeRtfnxGQhuzE1WlhuI1I7KQF+RQcL44JLuNq8XYHdW+uklvnZM6TwJH3wR
BZhiN9L74kmCi+b/4ukRxbFp7f2eeKn8AIpOCO+NXTtM4M9/nOM83kLP0SKO2u3G
/f2HJ3xHTrNEGTrlHwnwWfbAKhjBuWZBYVTlLpBOfzE5S1/XyAQ6uSPEAeiZz/XL
DiU2mE+zQIc7xsVjT4P5xvn+NuQa7OU4KSpvNpuVaqsGHabp/0EOtfHlRCA9fWSg
+Fhs/p6zvBB3P/CaM4rZi2r16qVlkGj4InknSEhlvXZGimvHA216aYneeKei4xG1
syAZsKt84tQZvtJO6UFGlFx+TtHk4fNR2rGXJhkiqIFOct+6ki6n+LbmcjrLbcQz
z60743Ge0DKdOA1jwjzmsv7gYEtj4QR5bxLsoVdLIAVJfZ99Nz1GcqplwNPQM5nC
2u8xadZJ7rUnPyNljZGUXymnIxx3gQtwqmf5gVS6KzaJBhwtyoePGbFwKSCW+XtG
Ul8XmRjnzB8MUpke3MvL7c77ERdCA8CcwJ+L0vw3O3QW7IRspTwy1OnesyJ8a7T0
5oPDctHg6ZG29dB6oElO22b3gfl4arPss03mWBU0SqHfWPzZlY35um8igwZ2/Qh2
hbEFlliysSCDr+rdw+/Ts1Cr/ee2xCwiJtHx1rmZ6f//J4lLSb9wwf/iL5H5Q7C5
GysRLmKAr836hMykwaCnNRtEvl2fx3hzkLI5CCGmeC86A/fitTrx7WM9wY7yTV6O
ZwX2CR6qDbqLs5RWQj+QckB82IDNvSlxBihYk41WwihmD81DMZjZKDjQBZD1rgaE
V6VFgHS1nB9XZI34Zajtc+AtYACDtnhaZXkWmPoz/KtPyiBRhiNXNQS9fHRkXj3/
eeGySbgqL8ofRC8YlX8tRW3CgbGZYIEAW4/90Ly1t971EgT/neTyFyY820pmsp4i
U1Bn15X0nXOVcUeEaUO5UIsBLP/yPyprJ8E6JnPfCW3vwJ/I7vV+Du/a861Lq1yO
IyjwndF5/y3rSmXC5UychzRnZYCqrHSnqMQW69C4yt7TT1Gchv0ApaPSYkliTgty
JF5TgyFR+yDc23oEf6gPsXI+Nj+EmNqKtWGJzZA5f1bnHYO0p5QBxoGYXFac9ETK
GP4EVbwg225KyX7A2EKHMBJHdLsqkhSBawJz+DrHFrCdQfq8aZLaECWD/iuHez3g
aSA4RDH95dGdXTnnkSRgT8YQ3rmmJnGo0Ef/e75SQoJmuiEYDc3Z65QbgB83CnEA
ogPWSSDhBS830gsQLojAeGSEfBkzPWBn/Ex3GY3PjWaiOO+1W4uQ30knyfV34fY8
0YqAoZ6pzcb9q7b0D7CR+Q4B22UHu9ZDIkTW4cVM3ppfVvexELN4lEKsR3qWiANN
qmSlahVsuUXek4hKgl/jpYVahPkRa84/K4sScEUi8/wpYUKmA+J4+ZzOYauYNJhq
UTmg47levcDufk5cl9u1kjKq4ZRXDZMBldOJ3BZNAz4sB73rinTvbgAsSAV4Xkp2
BCI80Ls2XBmgvv9UkgWRco1j9b6o3p/ttA+vW0i9NqU0doNSvnavRPcou9TaCn8L
E46hS4NR6OGJu2k+YFFi/dGT7k2tvIOuJSiMqVS8za2IdgCgOwOuOUMdx7n6KGd6
U+CFeJdV8YToaHbNLYxjQI6XHb1C3ZezibprlZU0OPGzs5bgXk1DucNzB/d3kXlq
xmPiDvnhACGdPrWL+pXRnMsWNs6LWw/rQSXOkp00i2TJt2LH3m4WrFHl23kGNwIA
iZnSspPW3fit8NTsAJF7aScmhigJeCVBm8ZbMWJkZlmMkz4xpICQdsXfeE3zn0nL
B2y7dKtt52nvagGMuOjSW/fEH2OeLi0EcszOd1pu8ei0dlWbLOc13zdyXzIc3LFy
8HXQOdC84STUbCh9cHyNA57IvZ/YCy+J3fSEPgYlK32isWPi4N/NUY0fZeJfktWF
iik+in/E+Vei8fetY1EAOgASIBXNbxE07U+9I12knDSzUZ7mOCzn03hhrk+fyn5N
GebbgcJovoBydjPk9whWimvgZgo73SfXE00YFV80Jbs8qSLR9M921CzHpF/Cu/uq
6deG3JJ54AXJjuaO6DfivJW8fXe7R+DpjLLfnw4dKFE42X8ciGHHcc1kieW1+LF/
sEN20WwkPGtxM05dSj6Favd/A1iYCghDSqTUab+YI+YEdePYOq0cbrmfCMB9Nfu+
CHvyG5OjKc8GiA/XRO5ihb+cKDex90xi5KJEKCihZZD/+RCdTt2xD+K6w2MjZQv6
1nRP905oxPm3xBk16NdiY40E2QOV4Vrgqb+t9E48OxzNQSXW8fc5ft/W8ZaqxcQL
qQs8ZX3gwxo+dLtC2oPunNJu5sROCZwM4UaTxr7tYTg2NMBMlho4HNyhifH0xpap
tj22u/8JJt7xwdZArlqLbJEmFhl6hAwKK+en2MLp2WQ3yAifBHYpZqNHW8XxFCtU
4GXXUXWtiL+VSArX8uSt0/GggdJEBBF/K30zANxEv5CZF8GPx43qRfsf8Koeu5iN
weIItqE1eozmpBjPqiZao3nrx0YSZIRgi/aq3VGrTqY6FG4jqSy/o/Y+AtVKhIiT
rFnkqgq+grmqb9FMOIV+kY4qRjhUOGawrNtnHCA0chW20Mq+vOTiF8Qfpidzwddt
D6VOr7kB/cdSycftagCVdSPt0P91MJF2hIYmsDz12iMleao6MvbMBNiQp45nAhYe
C3v8+FdR/KEqpQI6KxzJf/eV1v7ETSLSx/3THpdCT9dhxN8mvLNODBx+Rt/rM27B
1xe0E+0VDbBDCep1uAeDbONlG7YT8TO4XbOpIqE4oVqodCiA+yr5wVCUFFRbsyQZ
uHf24JH0FZqA8exWlNLJvzztxrjxsKNTLbB5AQ8JhzNQn5bc0W2V9qrPDmmLMYmU
lCzNFy/sAjcg6yI1ACx9Ll1aaybOBSb3/hkKWYJVDtPWzbLOEgyuYksUNqzBVcjw
vXhashLuIxqLoqkiDYd5lMGPk24ZfbE9SGUu/nf7p0aFFj9T7W409wPDW9GjOoMV
lm5CbAiOWT5JKa7iftAT4Sb9HVmWSXru8seM4c+XjRE3rTQXZNiVHy5y5nRG+Bcq
ltiiIG5oReB22sFk8NcinGfEJvyZrN53r/+a4TbLIri454r/IVFkJRUuC7RohAAq
gdtS4ygkpsvZ0wGL3o9fl6N1ffMXBAhM0Uu1D39uNmNu0xb3ItKI+wFKHq46AqWS
7eZEEEFX7/O6HLGGWIfPt88WHljlq8T/iGHUPMqI6YgzL4/4O4BQG06/GnGv5NcQ
qE4liCx+4fnLlyE64SX9TfIDsre9xc4eI+GkmwdGfXDfqKUWxScILNfN/WKBPcRh
NyLnLaF6zY4qi8/tUnHxTCwjRtgucRKebSx+LMrOSCFzz9UCPP/tnBa1t4mfzrwm
Nvgqr6m0GikYxXbI7FGV9TpdWc9huP+gOCDyRW7SqjTzWic3HgB1cvhMENVwVVil
xPxJZBOKV1NrArWKY3gjhpbpZPofEmT4Kn91soejVc0Jf0RnCr9MNxjx89QKRvRm
ZAfKymdAY8P3aTQanWWECHfx+2Sky3DF4fpJZLusLm34Tj5qi9pzzy/NCJc9H7uw
HXCvPP9pf3Z6RoqrE3bmdfIPmMm9i9e8ypgL8+cJcRQFoy3343M6/ZCmVxMVMUTq
U07Nz5eiFaslPJfbnLhPmVoDNPEr67JYf6I0mEkQVl8dN+DKGuT9hDxKEvLpje2s
bPveVuYAO1Z6cDhozXj3bK71IApqVhhvBIFjFMO7/loe5C18YGWS0rcteYu5O3cN
CyWTP5FEvTA6a91tAs22rqmssGIK5LP2o9V2UDjOet4CFmXH+UMNCVMjZ+zZhi81
o4Cs1nwGcN9sStJ4Zlxlp/IUtuBm1+nPaU5xbcwT6VUKqtBaYDcROBCR53Bf7/SB
TZctfh+9TY+WfKyjuKZ1+FlP2yRO7B7ttYAOBswd77KzvPSTXy6d2NoVYKMcBnEn
/5gmu8/Zk6dHSvoLMNT1i5NO1GWCL8juJKcyIj4Uljaxt7ckCa1zbNx3TNn7gzML
Xs3DQ/jWYUge+Ji25aiCWRXwivd0XmAg+RMRtxlHRnYjCjGFBaZqCriWsTYjWYG4
IaNxzQbkDZramee4qXxYL7mhq1TNoqPs80vj6LtS6g/sHGdVgleZzRZvjk9/ruUV
aEL+rJgetsLH78//n7R2+9WJaenYsJC7LZDaWJ+JPRdmbuLOwKGap1/IQhDFB7qu
CXkrLHZr63tJ98Ujm1R1XR8QmN/J/RAymZPUNd+ofoaNStAPruh/uwof1lz4J3OF
bGImQIgvwVlaixp2+WyEgaes8v0KOONT7ELQqznqap8pFRBglzpEv01vAYuJdozw
sENqHYvC4KpVA7MLk8fWR4FQNBEw6fBG7VMgjatsbMH9vHSe3Gn4jKiUcL1sMnje
V6yFV93zYsdboiWE6OQADd+PA0PJNI1C+bzwAnbpqD7JKGUMd/4DfR/YIiy44yuA
9T7kdwi4YIOeWwAhlmcZJyAo7/tXI0RqUoPkMszQgq7bX5OTZMWEj9d9n/Xp6M1g
Xn/btbiseRMCqjEGVGDrvWsUW1H3SsnVE545ldRPIsjwqwvQkT0ZPWYjfdg1e6wA
USBWsiD8LS7cePt9wE3gq2kOtE0ca5TMb4tnNgpFU/h+tH7uR/ef7F0Hcjjp9cvk
VRltwe8/O5u9FtRFJbw0M6UtORA3cTDHud36CAWymavyuzi42vRLLaIKqhxW26Lo
e4lW1i+Dt2t6vFQECa4FpwVHK8wRW7EWTy42T0MOYCpIVX8svnbfYoLN9nq/iLIY
Fp0rIdjBQe4/wkNnB5xq/vN1fy+3wgzbGlkP0mtsSf1T7m6QSq0z805T17C8ePs/
FgadkC9YGvh9nv1LWjdWszV16RqTWxIa909M5SGOKpPI+0JsYQHN2EvWugf2LhBX
pT7YQvCVX6uR9i4bUE2oUhuLlvxpSW41GmNr6SyU+4rl3oLnc2XFb6qT4jQpRE34
Gql1MRoSbT38TVoyGp5xJFdeG7f8T63lIAB4MZBB6qldwELHmPF3Zp7jdEbTEsGe
PMmjgJVnG2D70boC3XP7DH3DNtVHMoJA1oz3guyw9ZN3b2oSpWrTtVdYe3BRNlmW
lwn1jt7FeaoVeTtaRWPTY5R3D5Y+yBeYlBYX5Iip9VblzjP6FGhvOX6p/Avbqls7
yRk2ylAk/0PcB8B/R98E+OwtNizmZGQiRZYhEWQ7/tCdhsRL9+TpQgKLxKNVH81H
OUxannf/tfft1RIFAgLf+eTpOtnH/XUwyCaiWz5zb0DaZZFF5LEdjirkDRqNIwkB
zxqfzUAr7day21nZ+sOlOYCveXHDU32At2B0eKuqAUBGAckKYc3D3C9vgCwThnpl
ZnkHq+VLP2WJ0J+w6NQLRy3mSSjor+HbholYEG+FW0rEgB6NiqicGPrt0HaxO2WV
s40RDJDgQPATtcgS8X1p3wUZeEeBXIzMIwENn78fb3YOlEus5pQKdE2pbkkRPto6
2gmgeUiN7pdU9sEtp6b92artTkSiuILMWqQindgc4z/tmYXc7Rml5gVxfw3Zqii4
4DxF8N5ADdMKMLXc1Q1CXvAao36xpSVlGw3EGNq605SKEuPhomD0ipJ6+OfZ0MkC
I9T2Othl5RnkCkaAiGL2ILR37Mfjt6uiWRk4WARb/8q6P8xZ8GMbVKF0KYhFyn5G
25/I7+k4jVw7eMP7WbHC5CEuS+p3383og5CkwJzmUV5SFUQkcFIENJr69K8CHQJC
WQGhKyyOj2nm24pUge3HmA1b5Nzf7+T2wGhwsJdrF1DKa9RmqujHR4DaZojP/0aH
/BFEiOlMh1aZncNrPBlWresBO95HzzfbU2KnlxzKZPlxl8dgiYrb8gdD6p0d9rLk
7HlyAfjIxUbSu0KX1zy2vwdqdJyIZQgfU/+J4iJgV8cOKAL5xrRE+rU8fs27R+XS
CPIrtS2UqxOQ874wX9HSekaaX/zLf+jlFB79dIe8UyDJ+8HOIRy5zxHRETlHxWFp
aSEipjjFGJ+h2rItO+p4aiqf8z+D852WuYq1XM9ueNhlAvg2ZYekKdE1cNk53T3Y
R0B3b1mDYswNXLgYGhzwWTJAKsBVdVOEOBsSYRXjMVD1nw1Xa/4NLOVEkMP8P8WV
fIQaHK04j3PORfrKhoize0glfV2GSPKPAu4GDf5F4npKrdvaa5I2/cn9WeDtJ897
rDHx1hnU6AQRnw5pyXnlvgfpMcfPnpelbl933DKLd+M/QXQ+qFb7IQhD5QEkKOu5
N/aIul8mUDaXoYUbfMzjaV0PIBM7BsBgktRPJd5I2XrrLxwU2jxK9HU60OK0XV47
DAz2nseMaNxqlenqYodQrwdBrqDX/Em6Fy9HNBwJTHUjgixOZDjEHxKfmf3SGTr4
huHGB4cA3llg7+JidGLjSi1pkZ75eBqd64W7oHErglAAcVqHynb0P+BfjO5uSXsb
7rbLfV0lHOCE2Dhisx7Ros6msB3y0r0VAIHj65Xf+CSSsafcbVkTn4lvk2HhgpPK
egtg9HWUsTymV2wIa97Pg4Qctn730sxXpU/snO8FBjKFp4LBHe6b6fhr2LTrzldS
RrtgInSEMX6MbMM90CJrCgaVt4EmwLPImaXSs6l1WflZYzvOjjH9rQbmKoBUtsza
7qimvqp1JLrrubRxwu3Xv4Ifs1CYG83nKCIJhQCe1GYcPAGqFs3XqTVtgISNqJQG
Df9lekU49Fa48KE+4KrR7DieYHWc5IefcgTiaYfIA9RTfYEkd/+qzMOC1Zl4EXLE
LbjHKf7ysrb3pn2SVpIhP6Q2cDaZ9/mdLPNiUvHzgV9e0sgHajnAHlU/Yc0wukKj
Tj5uxelCH3oU0w2pI8wMmYMYt44V7XOau5fZmLTNEkPX6iBzF3EChFvR5uMcsG97
SWj6xaBps5eztuBYN4ot0nH2JX5v8s9u7STSUoABV1SrXiPzkcmdbjOWxpe6EU7a
nVnIEmci3Ya1Tx3hOQ4iLHdaczy+Y6xhnNAepA4z5nFd/0I8qZU28qpSbb7DG3zc
SSSkcsaeKny6KWsaWpH0xkmAFoeqlcJwWsYrSFDvnicjolV12f5M6v/Zmt3a1k0q
1gSMAVxM5q1o0QN4IqIg/aicrBl+z3nJV7PIBGaDrlpDS7Uj8n6uH+rQmWq+NjMe
af56n2VF2uBaGkOtTx6mag4ikmyQPlJCOIchG4XCxkAQqAsNH7YsJRVb9nvyll9i
0WIzwPBpMp50lWieDyXk7oBipqdFzXp5JL6sqQJJITv2uudYaP++KQJOIenDxhTA
xGwTAp+nOpBaMDXv6n8GV+z+ueo3jQ27dV41TrCSbQBcC7vByaD31I+cTwXH48hH
quoDbN9PjRq/PWo1cQ6ixr3Gjii7Mh4lB5ELdf2p22jyg9sAQY3/KbrqxmTs2NjN
l2Uv90USbDihubv53/BAeVZUPWip4Fu3QjtcO4cR+Mm92ivekfC3MRjFHvPKTFhG
RV6yYrFJN4cf/jVOVNKQufDnusG5zascPi4B+jylSZoFle2Xa2hfjEFgE2jeRSlK
Hd7e+APtwUxMODDF+rd478IJsUb0TINIuG6HiPRScKM/f7LvhkoKJOomRPkx60rW
pPsLhUCd3LIInnoMJahxnwrvMgoKyghwWwOcE384w+u6bqS5GFM8lZoC6jbU4CTS
9eGhCdqLa22ZKLeZHzzoSToSlJxNmSChXBDowgbi8uI9pGLIluLjsmBqZd5TjDJf
lQiVTt+vfh/JKRRHKzPsuldsDeb0IGvG8pnqPaRs8ZINfZiuhkUg/HZHv6NKzVyl
czlHSSgJ+3CAfFl0MxB1hYjNZ/GZBsqvqTJh5UpGZB9eZHr91F3RmVLJQZlX8Zlv
0spunivUnABDFnI6ED+pXkSBjR9z1ssXRMTXUtJdgj/fQlE+qtGyjIjc2dWYQXhR
qQwWYdJjJNxfsuxMJy2N9+puScJamI51+2709Wt6gSvCSpdqLSrUKlntvRwN4whG
ka6LTztJt7RiofJSbED7hSbj9GPythb/UGKt5In0XA0HGYc5BDZtiEHlR8AWq/47
tksKdEG+R5BHe70Ww3kd0GVEOvD6kk9gEi8EUocR9QXCMzN7aQwOSYJWrDk1ilcx
9WPD+T6etSTuLU9R6g8p3xYAdxlmAnjGES7+7XmUGOHJkwI2nezZ/hBPdqaQcxG0
elThIHYT0COcAjyeYolBwuWfsiRKq7b800ZLHH3UJKl2/j3KdowjOmnxyT6C6pHH
8ao+WdEXjFcVYsdORe7V2jrZWc1biEp6dOAk/9CYAv0bGc0wmvTBjurDPpq5qmOV
a+LZauvD2qXTYBCzSl05NkwifjCsBfv6rKd/dkdzifru03FoYRf2Ge2VGFimeRuD
vTIrxA5EUERnZKmX/oTuNvF6vSSbY8mb8BH2hli78iOW/gYebhAtH3oyiTqBZ14X
VWBnO04isXNYEhdOwbaORc0jPXTD2tn29h3QF30KxIdkhGg9oaPm4i2zDgSaLzXf
yghQmA19XDsrDdxQqiij1z40I7yJJ14FpnZ1w119dEGd0rNCRbz0g6HemKqUgEpC
3BOIqIbd+DCKoSK8Xjr3MaKJWi0UtDqXcLxXtPwKNtxCU1/ip1m0QGiluU54f1CV
m0pfJ6MGODc5L5i8aCBxV8mSY+K8bWRgPhTVxMlTj1eFUIboWpLQDMQCm6ZhTZl+
UU4p9mnZ65yxD9hUZcE0gG0ree2l2D0Brwd5qIGuafFOPHSdO2a4P8QPNKXxb+Kc
k0cQg7n5ctCoWagzJKXxhiFNWqUhq0Xjjz/aKQ9vTOC1cA456hPPQWWJAWwxdLhT
PxeGLqUU2r8TV/DlPknRWKf7ahV0OuPu94zljQEhfkiFAfvEgMRJuHjsFxYhjbiI
f0mE4klfphGggjtkqQ2AiFz9XoeSxx7qeqO/UZWK/YUPbl6JeBofsITSKSiSwvuy
62YAeIAUVG8R8GbfQYoDJLdj6qcEzod7xsCuAFo9nEWEdGL2DC4pt/epd4ScDK7f
OJOj0qY+AmyhV+zclmo+M6TOakYEU7bcUAW6TV7ZoNSPwiM5Go2vcThWKc4vjR/Q
inuthRgZJ9GAMCF4wz1dGWahybX796tjKRK4rJv9yjZENJ14w0yinbBGKBtAivPL
CXfBKAW28fLBqs1MnI8k2gt21+4YooPSzpwLKERKQu1XpSNoSXTy+3PhBuT5B+lG
5oCFmj1c1vE/VI6rVyduBNvGD9fP0KXdiuEe3GP7AYveDAOe8Gak1M95FSuEwRi4
ffWqkoZgygJ+YnMGUKVNQVX1Qi21pl1wzphKz8NYHi2wvB4Cy8pFqTwa0nb/Cl8h
NlF2dJ0sNZ9xW8KAVc9GUsjE3TpCZAnmACwyCKQfiDJXNifQkQ3oYNdpF+H0ba1Q
8bbPcqx5FA9kW+rr++tWMTqLH1bn0Wh5NWIZaYK76/WHesooAbV7Y11x8iGvbh8s
AyybCTRWbcbtvVNfcJijqKXpJ7RTCmRfsp23Vbyyhm/6J9XQqyBtE7hiEfFm1Mrp
oY0DQCaCHuzMfrVlRIAqU3tULQJybe543K7wpYBrlgPehaVyl0cF/3Kg9iv3Se+R
X85S6hb/VML6ClpJTv/+XWnqt/Ul8qC/DmDOjplfasy25XIXnWCsgwSIM9R/HMIx
u96WxY/C8z4PRdYvzY3FHaqi6Vv46XyRXC2nP7vHIQ4XhjB00fvveCzygymQ5z+8
0H7N8sGSnpQAUA8lVi9LVcQdxH0LERl1iH87Vmy9iWbv2lbcOh11LD6yzqmU+Swi
YccENj7Nv/x7yQ/XukI9kqiNxt00Bm4fpuUdwCDTgjeVxjKiH2NM+sLaEgYRovRY
f9C6yPmqH5J4ajgxygnrDVV6PuM6lSRXZJ+xAcaak/tvKiJlTxQdK+Hc+WOxZrBW
srvoyBzfswvG1GF8RJExMv5LwJqQrmbxMZv1Q0sxlg6f+1+VIP8IQFiD3x6wUBZL
2AiDI9cBRQitgQaBngByQ7MPx3zw88KbDJz3n3PbsMUVfmTZnpjhtgMLD/8zKNNx
6DnHTMG1ZaJhBJX3p4/eGlRdFljZGWQW8ZbUQ438/s4AflktVput/GfnHjfd8GlN
YnEkXRKj2XLG1p2r3KKE2wpmZ7QpW2AQy8REQ54RHB2BpFRGTxTwS5v55mqopUYq
XCfNhqNxCbtuaaoyYTUhbOv/KsHcojlwXUIQQPWffRlxQqZsrZEmN1BtuyXWJvbE
cqOKI01/Z4h1CEgYHnLLnC145kGtGjgaz1yNPO17eiir65YYJRFlWjnkPSnZBWSr
k/cjOIz8j8aBHXg/V7NZrtrd+24FylZYtumoLxrwf15h7MzDTu11U+aByrkSPLYg
26O7QqUoHxX0TNY1nEdFTdiWgmzfknXVB5ZOACFF1NQJuY9LAErCm0pb5RwiBj9w
KZ2s1rmBp8Q1gMpgZmTX1qgWyAJkzGLMMfy7sM3OXFQRwESDBuwP0KwpDQ0bfLLp
+b15/P8YiWdRg5I3Gz2jJTOJYRAeqKT8Ncyb891cHuVCCEUnGOr1Xt+ZHKb/rRWk
FPMvREu+nl19S793Ev+ZSqeb3OLRAntJuIUW/p2gvf811iAeO4UNA/G76X7R2Kqt
UN+UPH7VOm0tEkhfYZ0UvZ5OGFboH9GgxRS0eEzh//w2VhxjXgRlggZ7o2J9IW8G
Eu+DTP7J3mvNqlPIRbp31qt3vBdBn5I19I5oQy6Uq4Ca/1EFszj0JLtg/szGRInk
tW2WGJoB/g/sBjcSQD5A4hYA9M8vz30oQHg2Dec3ZTQYoq2G8fHL18JiDIK5k1sq
fKUbQousHVk8qNwJUfxrlHFcDS49iOxCOrSAHJK5EIVHjJVtNvwP6aEcrV2DQvwX
0k4tquUZlRAweax8TBvDYq9S1s2wPFCWe5l4vEH3lAOZKcAXoDtycTHJG53oBZJY
SurJhPfFUjHrZip8isV8Rvr91sK//ZHOJppmGyX/MtGsqZNjB8HCpeFT1q0+zrpy
k5E7qOQzPIU0w/oNZLqRkfHgorL2TsirFWOs/svZd44EHRPkft6Dp3WQahcCEsdL
iA83yBBr9z+sSUV5UwBYaTUeU2V4RkRLEODQPaJOTeQxbB12XX1nXWErhGHg+jK+
spAM0KHFTf+Sz7zoE2yyqU10ZxYcRM+yLi20xz/Ejc2u14BEd6dMD7OoYIwq541D
jDQCdbg6bvJFwo+PqKt6Gt2oNp/qHBhlHDA5hheUvrGNintnx3Nca+a0Km6W7vSA
q0R+I9RN9jTybJeGjVzU4vnAEDS3DO7skibMsKdY8Br/Uh/Lt534bVShyia6q7Rm
zEa14WVD6qcqCFIdxUNlVdi86fefM66OOGjUDYaAnVSVkXJLHhpw2iOiZVAgp6P5
wyi43xV1FqgRQwhxZh6ZYcPV33RV1kESGYYUTdD2d71MNazB7NWkQbIoce7idH6q
ZkBz8UfEm7hJ9OT3S91rYzH11vXDYTSjyTKUjdR0enFuoLfFhOGUS4sIy4DePHIK
hddZUWxD08fA998TYQrAXqIeago4V9F+ST+2lrF6BG4pfRIjW5oO0EidA8nSX+XT
TR9+nvPGBuX0omA2PwHqdBnFqmlke3cPIx/knFic2TU6tktCzeDMxWHTE93zo7CV
EDBtSLz7zhZQQ5B6ifgceaqoMdhAchAX9tQwN/Qlkc9PlKT4oY+lS+qVfUOKKxCT
XYD6IzU2hW1jFLDSSoz+rGU+sUuY/1Y0QLd+vKOi6P9bCSyP4zT0qyJJhpoRqkXh
/2NNircQIZ6sdMP272vPzf6zLFRALDXOiEhXbYUZ2nIDcF/i8a51oYo1v0G0gcpn
x05/sTj9HcA7g7mU1XEVfqifwnIp7CBK6Ea7AXap/oIBOw6d0VBp0oofY1GG8EIi
3vwjUBbcF2XKfpU74NKt1DdD7reOqQONJKKEpESj8xop0fTbpUSXGtDBMtfKFn90
IeJCxiKBLO10kC88TIC/K23XBHpgn3v7HV0EFtUxKm/3rAznRRnSMVlQyzthBxMZ
gGuz2/eChfeFiAqZgjoxNid0Rb44HmElxURJZEbs8JEElkpjF9VQNQppB0J1y6ln
hxN0v/mWlI19NU1c3KmQ5T9KOBW4SzWw6FZoFKIw6kl+iCU9PwVWF8MpPG8x2MlK
8hdOI15AJenqkrIXVbvATPb2JlngJr/DeHYo5ku61wooJPn63+4WS6cY1ckN4Cm+
PBPfhLlGjr3lXyowtwsOIiuzkbX5ILeDE/lT7mWs/wqEHecItAqAt/0WQ/xnbE7q
6ksCaXBrfIQZPrG+YAns2QIWJyilXwaDJkfegSxEZ66e4Y3PBATg812AbZ+p7a4f
E3EEzr1giR9DvWlgFRPdTjtPWd60ZBMOSkTkWTF45u3NI7yRwiS0FGugOK05mdKd
FPa+a9OFmseg7Jy20tCKeI/BjI48DM+uKtXMD8yNPd+IpT9Q/o5F4SMv4H5Dv8gc
+PdjVd/uJFovD/n4az2eOyOAX4O+In58S6ags+PZuFE831T/GJGcQSGzfAb2JIzt
/Ygw07esnpqN21x0SuuDBfi3cRxDJ4+Z5dPfhpmCfcFmgoePiqgf5QIH2x6TCA4W
SO+tdUX1rPxF9mbb3ej3SkyprjAa5kfwIG9XyMa8pbOGyWsWum+EbkU/Izs9c1h5
PLPVe0B0fzJdh6taXdRTZFYxxqwf6LVvpdXiCbUjD40+e2/Gaa5tLYkqiwQc7yuA
TuXLLI+6MR1i/WCB+RVT1DNJGF/JWtA19jt/J0Iym6QfaA5tODTYM315/nRJKow9
ogbklViTA4ySXYHSyz65ZlARfvjh6lJh+A0aT+vMJOfmJYvICGWCmOoclxj8ceON
w35pgQbDHp017h2HofNihSOfCsCUJMY1BeXUnjRergXGaVhVZ4HdT+ViZm5BJO56
qwkke+uAHk8ql6WzkPOig+PVEb2wdZJjOjJ6CnvAUXVL34gO24KKGifAm8EmLRXi
jyq25/Qpe0tzxhiXzxIXH294c2SFefZTCpCkJpPbM5nub7tgnxwnaMcj+lTPs0Bm
dUI8ftEudO6OeEhScvTYmoDb2N0kCTDnCSWvWNfycYvEcupCJof8r5hliJj2NDaT
RzkWuvph4OVEjaoLlbbQfphdQ4MQ3FhSqVIOhpry915eZPZTpM+dvqjxQb97cm6V
HQtzklJitcXkhpKR5SOWtFdVb2N/qWFIisKXHS5BK0nH8Vihaqeifn+t9eqKNKWa
a0JtcLeWYm8jvWRsD3otOHNf2euovEQ7rD/fg2BzF7HESwITqytGLT1Bg58goQBY
oyjdv3nhGTgL2sEbxkWz7r1vVIKUHPFIdryUMJceFywOpHP6mw9CL8q5StcQosEq
hwmsJJfJbSIZEUYuqA+2j0G1Z8y7841TmAUl66BzD6X7uz2K5uznK8zYtlRejGJj
Bgc/TfvqtBdXeCN3X26zs8o8wq0O4QPIAS/yLzbxmlSbVZakwMrwAwajZfl+46VC
uQrwnMlf8qLnp/6XliSesrIGccALb2Pd37pNQJOmx0k8JZRsPCdyYn4iE8lsHkeG
/IP0GGTMYJCL39GkjPdzvYli3asqvbctCXg39dX7UY+INLinybk497PJmHRtyti7
I7Pi8fPTXPZRhevWjPy7Bl7N9bf0sA65x5Ghl614jrEn3v/QNZzWYwQzp+1AXfQW
jU5bQBHYS38NezM980r896GndAKl7TMSEfebLe5OsP/DFzWELQTIfSvu7edaKxUc
V2/jEk0Pnda8Iz5VXA/BB0HMtzv5sA4cMbvJjfgwhsRtipW2c1OwMJ6ojP3PIemf
qVuG0s1B12iMumWeBr5rokgt4Z9XXftI+J0QFOzBDMdHCZFQSkO9O/aoD4k/W7ch
fQwqJ4rrcYigUdd3iT1mHq3F0jjJRESqGO4z4ASn/+rUpU1t660TSubhix0rgKV5
8CufnzlmAlzIJO8CIYTX0rxXRtwX17XCVpG1FIrt1GEpfSIIeqp3Tq+9kxGbz2FJ
aUR/zfm/PmXYTg//MyyfdkBsJ2SYWn4MxgUZ6zBYXJyGRNOa+C/KPWi02fxPT0WA
Cm76/iutUmpuusrYs+co3qwimGt+euynRWPaXK6yaPZ//zcda3RF3571Ki1QQBRv
tp+j+mDP5NMhyAmkJ+rgK1mELiFbLpKV/pYmnXRBu8LNV+t9LcaIAbyNzxv0Xx96
zwqjghN4n5PZZJzswl7qdId+b4nUYcBprE7cP/dNZqbYSwWxBC9LhSjk4c9CpC/u
5THIDV64X9AuHCpiOfQvR4bOex00Pk82uyAYFD54vr3iqyhQHEhLhhEJDAio5yrR
OWxS3fFskNcCY8cCqLrvddk7q82yEVe7hTdhwVhS0ypX1+6QAD3/AqJ4HsYCWZC9
oMSeCiQbMl88/AyIxw+owgJMIVw/Zb+OaiKYioCD5o6Lw6FrIiBsetQoCanKuAKs
QjTrnovHbW6iLEtkWuiDlcn9v9wC0gRBSaPcnzwo55xkht+JeKEIfvfscH3Fq+kw
Gqo6CP+OFpusJmyy0oVY2egBVJiqzolVUhK1ykWLssRdnNweGrH/GT4sIV1o6jAB
Ng/n5/vxMeicfUf0d0Ecji64WOZEScVZ4MwPXGc+fz/461xUQkpiBKBpLdSEpoax
NrW6oIaxVwsgHcNUQY4ZAsWZiZ6HN+V66e+Jfxw1b6Dehv1wzqAPwOXb2IT4bWwe
Q/Uq6ImOnR9yYYaFt/Ld2JMYqaJfsGWruA/TJZ1u4XI2D10vdvIuDGzy8Bwjabs8
oAzjjH2JfmU1pNBlPIzQfk0D3y3f3ZK6Xa0H6Pb+hFXqfb3Cnu3cPB6PurYBGtgu
w51Zf8T54je2WHJo16/84B07H8yUeWeLMKwqRZN5BDZa5LA0FNrWtnOmufcXymrR
zP84cPgkibhpf5PKc+eIeEEZ2PI+A4Xn9NG/imOFJkxhZrLy9SuOdsU8HdyzzpMG
IiAeMLppPedw34AHi1xNQW8OobMIMXJr4uIboqSkZn+UpJ/I9cFCms38qw9MRnIY
FgTFU1YUZl1Xnmfl7vSNtXLfz6totaiB4eemVn9qDGwvbq3NFG34PikrK2I7e2wD
cvaeyZhZN84Uu6Et4NorAZlx5IzlPVNKtry+/Sq5GWP4hB2sIjGHXAkO8zzaK/Ht
dbjNhX8oqleBzaE+DL8CHfE0SP7OARf3gGYSGjB2m/pudQ5NNDnEKTkkeLDXEXPV
HlYRUuW72O5ChKy0VkRy+cyw2XRTkvdO0DYVG8dHNH4nc84/IK02cXeoJPyeUAFI
FLprtygJiyxOBVLh1QJ3CwXzmlKf8yj4xWXzgtMyWYjtZ7owkXEj1D5LzlbFfyMC
lStG7BCzGfoLtXWDw1DF9j2BqGOxDeOCLBJ2gujamx6IqGvqZTqL5Wtt0NzdbwUB
yYLD87WcAV8yCleMSCKUNveg8JuhZKQ0T9X1SFLtq7MLY/0PuN3EQAzDZixF9wG8
pviUoVvaS02il3wB2OMyQG32xzONhsdskJK4vm/8oD4blBIsLYSg50JjSu1qLonb
90ROmrjnqDgSJBsflQD05bXq6qKd9cxoDPr0RcZOIlpAEjUp1B7meOiESuPKgm3p
whY3oldw42BCZlVTi6ALboXoJtVx+E0/+umwOgLE3Q22RX69yQK2xXFoC3r7dEgr
Wuo5YcYuwRo4DRVGbKMFvVRQ42qX4yeKblr1maoo5U2qIf8YpGgn+bhbClH42GF9
foVbqkF4IJs4BZLcs9H8DrXVDp1uCHxJof/JUGNz6B4l88syCXxz4te180KMk9Bc
V3sCakeUy27J+GJNkwdMWSLYmzkZII1tOvbamnYErGiNPBH4LLF71Yg7ljaCryYX
0PKLewLnzFV8d33yq6ee0qErqlcpEJoIJjYjYlRim7nP7gPqryT0cp9k+uQcL2HB
RHeemKOKI8H/iJ3H7U+tWAzPvSEp0Vi1zffYnAGjI8LOGrQ88xJunmCLmY1qo0WF
5IpsFC1HeivPZi8G6Je2LnvxLvlAyUrh3uC6BSb3cqXtzNaV+F8IWipMMt+Qxddx
yVzblPOVsRbexEHhcd1X3kwMjw3KaoNGmHIz+OtxNsAFLvnnWYEg33unrMwHK7E+
+5moCtHhYk3+Ief5+kqTLgSu18WCENTlhfdqwDYI74rTJuR0CUZVP0u/JrlqFRFT
aiFxo8236hF5LUj+MKqQBCmrsgku53m53P8ZYr8j61WSpd2d2eoLfaGI8VoSSjuf
AVyCVSwNe5jJH/khplYm4zsk/rdIahCNKs6ryyr4oOCzzCpz4n0/mJ1DcTkz1Agg
i9dyFvZBSnXubTP35LzwXtWjL7/JNXtKwHEp7yf2TEstwHVShBASeZPJl4VOgSbn
tShMpyH6mtvkf4WaUcheG9UhO4AfhxYhivFdTm1dvghfBJyxbgTobDnsCk1omzXH
ZRDQL0Fslje0iRgljFV/g4AxFiYsk5pv6lzDFlP5KRJEpXlegXDicMBIpjvM7EmK
kiBv33aph1seoIRYegwSMypr+8NGTFuvZlkGOyb6uQo34ewNkOTTKI7C1T0MnzLq
R23ocI2EOs+fvv8oCe1Oj3IQSJHUgHJuzx0Ud6YIPSLQTHretyS78ZUXZhgPcesW
8mnn4mJnzUvnRxmscEvVNx841I/UnOfqFF2o9vWFFztIvbK37LuK1WfOpTILxNgi
IdyQeZ4aG2kJnGcOkXYnRiM3myX56r+PD43K3/U8Ok+E4eQfFiNZt/WFLeSeJEIz
FyXUEFyczq0GVZk2clF3RkRqyfvAEvCTtw8SySniyCGo3iVf2FINWy4M3FrjSt+l
n/WClNYvjXR8oQi4rs4Lvs+zmDXmKDdtd6x+GwkJyDOodv+ctJSjygj/Y+YcYCK1
TfuMxZgyuNOPnMM6KX/Onu/bBdCCJ9LpSB6ojUx5y809XRFPJKsSqQE7M9NIxBgG
18NU8+Bj+bmqAAKbwHXu1YCD54bdo5fI9vlEI4PTO4qTfwMNlFEgXzmKXBkf6qgc
GhXvoDlnnLxMNxi1D6+yb4A5LJuiGK3X+eMfXSKX9BEUk0xof6iuolYmxR6ZljZ1
oLrtgktvnMETYUqYHKR0+k+6dVqMnrG8tzN57OrXEe6PnE8TnrXY39NgRqb05tAs
RukkJ0gybZMy98NAdvaov6eWNSy/UIYserbnBsmJPgObRQQ7OFfCCVN+iozs9lDI
4ZSv9pfpQFHySRcNGMUQZLhF8Zrm5UxFHUf2c7TQwJCux7ZrPEdHtU1AgXwPiER6
ruqMCeGpx3W3oGp9C3VfFnhERTO7lLfAw4qGSfWpv7BCJarkzjZ6Jj3Wpuo7wDWl
TLbaMAXBLyYXIyq3pzQBngiVk1wbqDN0lfwQEL/INYPbv/puSPYnnaZYoD7dZnEZ
xk5oevvyaxGrSIKc+bnvhNN43y113i/+bVtY3wg/qEDIst5is0yOsjYp2xB/ftsh
Lc8Wy3lALZyXvyyWb37W9vdps5DmixmPdco8ri/j/+49iMcVpE6Y9OmqqMd++j5s
UrzzbtMoWor+9qOkXw7LcHj8il02j2wSs+efqa47dgMGD4KaILAJDuB7KHU89lOd
Q36XYmb2WwYJJnlGl3OecmUJoxezIeDZePVWxssChMwdgZRO2Kz2o/Awt9Uy6Pkr
Ga95e3RYjYhDaU6Fd/tbHEASMvXdlWsg0naZ+Ev2jF/Txyg1KmLyGPKRkGrgppu7
q8IR56o+XBKU/4J4XK1FGVtQYdJXX4/4VtQSbr27Q9DpSYB6PDBQIuM3R7/LA23u
43KmZD7goZUYrmNqFEpKgZ+SefNYKkk1oqCs86Y4h80nvoXydwCSPxZhZA4VIHrM
6lawf3xp6c5PYiRuGCX7MEMa6Eo9DF5rD75Qk5vnxNtjtlpqKMiSk43AcqHOBmJ0
VUfoAECyOa43pRW4mD0fcy2rSlVohUE1+a95fMGjgD0zJ6xn5T/p7jwE+1hq1MzX
caV8tLcaLWh1ILmCm35IDpR7wAPOnzv/bgz2j8jGJqWoTy08BUL/+1FkWN5VM0Lu
bXLXv2TIFu4qwXA3MexeI99iXTHMB5k4koV8/uYYxlrVPhEJdqsXUOsqKMxZ0+xQ
gkWn3Jqak+BghHMg4DBhUu1YzOqlLKyP4O/TqUILDI+zLCrdgejud64K0qI2t+xU
jusUy0vKDEO+upLJEHXaODjvpH8wYr4XI4JGp3VUevoGXTQu+byyGzWuA5C4yewS
6maSD9fgCjaMQasJDf4DGSAZD7z0MQqK3ZqDGwX1QjwnysM2m3QAwOLMj1G6Of7H
8w4hVuXFGQDLBOtJTG4f47wxR3OT14oA32OVcWAqJ7dD5QdDURBeTZihmb9hbQow
ne8+uJFbAlwXErH2p+o3KyzXDR1mNYaFBjlhPjOGJQ9ArLkxa25Cjh+PtrhgCWOR
cbIeA8OUW/eHgw4R0Hl6GeOkYO6M0Cb1a/P2uOIjujc9Uc26xm30hLKlsPK4y7Vy
MHtfgX/D4GjEU/PiXmy6C6hlajCXlSRdv68k2/vuqIMIYZ9j0zjTTdcltdYzj4ZO
kyF8GnGEqY6Ei1mp2sIqfJ27g3MIAEKZ6QJjzAN4m7knu3lQHaptLH4494VrYSxV
A2MHrrK7al0A0n0TU8/WDWXJzIv1M4hMjawk6+Ic9Vgzzs9yIGsv0k4I2UHDYpIH
1yCp4dHaooamwS1fRbyYCezogm+2+CDE1tnbzmJ691Y9xpVxOpJ/7Ogt2aMs1KK2
Wci3AghLtdFkt9VgQLWgsITSLjFrsMklq6yfgboa4rHnNgDdgUqtjeAPHN12FB5u
xfq+dclNmvZ9sdnGpeY+4TdgAmHZ9hJj6Zx5hAt4TM5di+ICO0vQ+PsHDG0V7qVd
8ILew0572JChvwL+e15i5pWczVYFfP3hDeZObnlmh1T+UQ+sJeXdEtw2XgijFu6G
qaZsHBE4tkSIU9VL3TTN6bK4sZLgcEs2Kk2FkzOJZ1Vve/K6bRRtgVoeShJMja8u
Am9Rrx4PUXWZf4B7VG6UGJeYtrocBVJck/8TR5mNiKNVD2gmPeACCPgtNjQTC3ow
4xncYY5krEwqtCXcLkuIBtE1Mcg9gahQKVm/FfgKIoxB+SvNhHbLjm8O4RP4LLB9
Er7Xs6UBsFaB7qtvyAJROO8TlbYx8Qy8CxaACCmlc0hPRkIy/xXfn3fgXskyFTiw
q+amIrOo7zZU3eoPxC3EEvQFB0rBna24pTAYGLZ42F0a0DkILLucv9qi/qPDWMuj
7E3WVmSO2OczPw4li19IBQNV1lUQkWH0s1xf2c2YRJf/kDT936d4EBh73bbLy400
PTxk6CpRrSGeTPhnj/VBDdRUgQWTU/WmCJL32CPCzXL4J6+KLvciyyo3y+dSg98f
gEEjOcvyqaNatoKThMuGhHnQS8VlUyY2O6injYOOnpcx3oRxi+M6cb8OyqZNZi5g
AUQnZIpFOCGZYZXhDGqKCj8EJReIhTeQXf46DI3CgKPX+fzW0iFFdLATR2E8NOuH
KqdMfBToCkBAK/i1nrDSVmhbDL6XbJtq+AMDow/0+mEp+eC/9HtgdJNOj59BCTz2
l3/ineziThPmNh21BpTlIXASegoinMjcx7hu1HNG4hwcmqTosacGs5im6YR2YrTB
xYNH8PJ4RbhaiBSktbchEMN9+zEa5/Y4Lo/60N5z2GowBKTLUY3fnuKHo4IPD0zf
+OazKtjG8RX3WMbHY4gDJE7hbNrcHTS6GtVoyD1pozrUnfkmAhMk54fQR8sou5pL
Vh/Fnj8r+nqxUsumt7QwSaGtKOwLnnA2LvntssH12LZYDkolH4f/u+X2Zg1M0nLT
/O2kZwHkqTNq37bIqiA5kjVat/qL3LivXbAzByv7o86NBJPwb7J4jcVJl8/Gr6PH
y6JsswA/aqgylNQCStX4j/Qp/KMzOWlhYNJudNN7mY+7SNVWSRprNfI87o7Qzlba
zbw5sSKHVSteh39UYgO/NxIoAa8tBZ0EPhyHKo69ip0wo8hd7e2tupHhDmp/TfS9
PxJ23AMuih94+fLeVeJct1bh38WrPpJ+2QG7iTfbIrnhno+WZYafXHfkvLrxxnpQ
LLwQ6LpfUIF1s/KcaS81+W4g2v0eiUozGaJDWLIGieMH9GwiVO38zicXbLyvfMlz
t/VrLCt9S19UgwbXmzSnmIPM+CUHtSoXO08U2JSWcvnuB749BStd48mISDsO9ECN
OS2ZV6kR/HdtEtWUh1taxeYzOaCfD9jJ+dHWKcPDgGlZDcTExd7YFkjVe/7xxTjA
nuDC52v20JS0YZ083RIKDVBXPr4BqKKYChaaWRgMNeszNQiud0lvY/0pyoQpTtMP
34T/UmVdN9BP8aPYwlSCIbGkmpmz31rZujfXQ+SYVcntIIzrRkRD9aGbWFLb6TCo
EWBFcWcHZNXFYRuze3inBo8ltqe8nHvShxS9Gybe6wYX/LFOIzfNZ1uBCTbOR8B5
rNxT9SzFKjOccPcG0+p0Dm1rjbZuxFL0pxYd57w6ozzKUdnYzopR4jtF35xDhcMF
XjJNQ0btVDgjuA8r9cw94jwmN7XkSRTHx3DTTlXfn4wNjBFkdn/CCPZxUxypuoil
NzpWQWjuALXrjItlPnRuE5WL9wSZg10g3AO/I6lRcztMH23/b3L2tpDBXMMdcPyJ
HIwme9damttKl1zpd7geFVkkyTJ6AIs0NJO12PugHyHwk/jRnhxkED9uyIKLXAaE
ICuMHd+0mBSJ2Ac7759sfTgGmpu7O6AlOxVvUPOBOntt6xpx86dv17OCLXATmfsC
e/ONJr05h+T3FgnUvFUdGN1mQE+54OvWCIW5Djwo39M8t6jaVgP+1eV0L2aZyA/Y
sy1QBQX0Q/LUwdNJxIdId09iQKRbOjGJNnxzm7qCU+eBcWmN+rGG+i/yocJ7sf06
HcGu28O48tlpzvBnEsvNQifvc8ifu8Xkc7lOxOIKTOfRTLZ9gWXWV1Tb4RmQz1VE
ZuBWt1LhZrZRT7nnWuUMo2DSvlGrm5HGMkM04VIMLguM1hCTjCc41axTr3G5a7WB
LAfWrTAsURH8sX5yEz4OSs+9u3zUjM3JSStAGFlT3y6pA0R3LyUnuTFnyWpHMn1B
P3xMlKzG0qU/wMrRHSjwHGVO5cvc6HME9fnPWpnAmCvoU+91RuizQO/IbmBSJlpx
+4mNXMfryuKLY02fIh5jIeP+tfeDtpadmfWeEIaGBxTkXSyjuDzF+VEUSeQxfZv7
a/7cOe/PB5nmSXMEwwYp2I6J1J6+gpFVIOkboVDCws02fX7V1erCPu57L0+Svdra
x63XVWB/sT+5BBgl4Us83rx/ma+ElaWH+bBmR+LDyzQvBTtuskJmOkHAYg2eCpGI
yZCYtjgMQhxk1scpa+l5raaVpok1ejYKBxE8B+0fjd/rtyPtKVJgUiZb+wuzM5zk
2VJHkizw7m8PcBTjKQrmO3VJqfnWsPXnFQEeD9CQcwBn6shinv1s2RtyTEMDWGQi
JLUUIXjgFIQEy+T+lrQc+ny+jPoPHSStV5fj2NwTDY4/Wt4+u5yxtwkKD+EERbCo
V0ij3KCJJaMfyKEX5XJwq0r5p6KNy5U6XHm5JY20V2tjF+Ez3A1urBhHxuCK79QS
uYEv0g9zWsucqLjUOtOkg6+eq4caA5ri7rAoNTVGBEX1naG/+Ltl/jJaGEMrxRCy
0LFuSdk1GA/hhji6CTlE4z9WhbFBX3GdU4nxUNy1RxsB3KUUKqX3vEmY9mUwkNcv
e39xPXUiYDmHAf1amRG7BPf+NLJ+VznFa6TREMiK/SkK2k2vlTp8RplUDsaMXPkB
rNDypsHG5MWoi4A500lT/MENadnnarFNkKfgVhE5MULzHbwpYy84T7l6qiH+wae8
co/DGVRViXmmvb6qbd/aG3Q8724tbJdmp5VN5Cn97FWlUnjsL3HS7oce8k2jyZCX
zoMNhm4o6E4IclJuEOz+1HkOBRQq5Z6VLeRoe4go9wzH9ebCKnmfQzRjtRzS2RI1
SjmezpDEFAKKypeM5FLrXAe5v1WeHjvSI8MX+gwWXXkP5ZGQ7OghobQKZtdeFIZR
IhxCwkDwMm6mQpW0gpwqYsQOJhGldnt0ueSsoKMwIeJTvY2g0CM79iNlJGcfTkSB
rifcjRsM6kHUbc3aqTl7Sj9fBkHt3m3BMCcoxyKDOic1HVf0HIU+rnrrtpEcSVpH
NpdG8TBlRvyP83PPKHPxPg1OZPG/NtSdW7aPlNbJF5gB8k4tMs9QjEeQWLkJgHCh
55NtsPzK/txWEFDlfVbPlvLTgJZ4e89dg8LY0yoKwbLfpqwwPCbFpPS4Wr3wtwi5
aYBLY1kM8CZcDNhVs+aaSPldhDR6vmmqqGrlnz1DgodALvJjmRTsbW4t2l7n3Ur3
SFd3nj/A8C+lRuXUuxSE22d99uqj6g/S0H0iUe5rQGG+mjIhsgfyPOkN45clYr5c
nLmKY1LtsHkIfO4eK65VZjZK8oYoMwBw7PvZmQvsI4tro9HSTzlobVHXlxaQF9Oy
OQ7RwJw5lE/DG9v/sMHJull4BWkK7S93xA9sa47UnXiJzAJjy+nvu5lyFvEQcw2P
+UkS7qJfbcAcpH9ud1iLhszK3IrH7uYQ+OxCcNY9RKUy4/97ElSoF35BZpZ/LVOB
CziMsUU4TgJNJyuBySDNJqqUbpuULvIatrwDQ9AG6caODEyrCczZk2KV8SHp2BAp
MnWAG/4kpLUlfYqR0eSAHshb0v3RLYKy1N1NpoPkrSNUrL7NMs4M8T/YtgJ79Y59
YJ45CFb+tC+xPI/JqY0l82Z2QMf246CMwf/rlvbvT+weupuhkvHs8/Jfaj7XReLw
QLU35xJmL4PSCpVMub/RHXMMkewayhvqHNPJOx6CO2yhndZy+QUB1NLL6c873pV0
dQLuuid9djwFJ/jUwdUvR6LlxKLiZuWdHfNPJFDki6s1lJA7Fh9JGty4tTw//GQ9
5Ma4oN4pJ8VL5jUeLtsv9BzI3hWYMSrWodfmwamdMeavKXY1KqhdPQVVJfWmyJuz
p78Duhb/MIrHSkCy4tT+uxkuIk3gfWEf+bCid6Bcft7w3D0/OfdPtrIuBO+UW7aD
lZiGM0TPrAmsmKx4RVjvT3SBAXkH99LlNe3WPolgmDXdoRg4y2kjAtFBqDg42pfL
x0bF+6dsT1OgcBhYo+UvjgYPgQt/i/8cfzbXxF51udlP1PF0PiN3VOnJyB1Hr9Af
hsPdlTM941dODs2MwZXasr9qvu56OSOaK8EqnmqI5sFqnTpdY50dSRJb141c+r66
mkI3tVfcQUkPWuxjrZK3WzpdZbWa53QmMHjgEas1vw2s9z35W7Rvdih9BLeBwZUv
8uDwuLqDpO3iqCidxVUEoqVGHBr2W79jFtHlEi1Q6DQRhalDYYJezsYrPopPxjWo
8jjF6sl/vdkYcdmk44pdf1PKfCWjbkgtgi71P1yAeyGjP9TRPsqTtBPH3CQPmnQm
EGLJevWJ3Tp/nslR5Ymx0WlbJFy8IpIc3bEiYBO+0EqtJN7ouBEm/g+6OQKUBWE6
j0RfRD4Ka7v0NigvTASguLo4gc1Bga5ClMp5HXMG5WyhqTEGia8GAhz2Iu9kMMGV
sNHxbUbZtKv+GcnV5KgQ/o24WnyJU6lUNWwj2IiWlhXKeCSV8Ppw2swX0WKR+65U
xOiaLcYADzVNvE42Cja7l2n+jlMc97Kv+NbifBRRkWGmdfOONHGkoc7jj2gn6/bp
GPp/sdTo714k2zgN/571Vpyt3Lm9QSIFDNXfFJx9wWpf5V3S5f9Mn4aQW3mbEF7o
2mTgo5H5asP6LsV3FKhJxD77vimLImfiphcaqv+Tl5uznoMWuuYiwjLyoS03X30T
g+qsAAgjAjalHa10l3WDb2LrVCoHwB4qAcmGACtKpZpBlrI9SFV3hLD2vfUNIaZ5
Lg3z/BA+UfboExZSe64pdUr37DZivv+AbqPR3OeHuj/yVv0P2rfZAZZ0cRCRUWp6
OyhMVykByn61X+IypI9t1wFdLWxKt9LAAsT1F9DRw8YlPFYVDSQOZ+ReL1V/d8eQ
lJekD6gd04xXzjeLIVmermKTD7YxME6QeiEOwDMA8xfEPFYeh1lfzvFuGTX5vQiP
jAramCKIcNg4UtIlNTpxJtF6m8LAmQVwbS0MRJTiuHUGWXo+mIyJusvsajBIk0GN
y1DYIBT8dBOGht6VswUyGRD9wSPwOBd7zzBS6J8FLqN7m9GqP8XADTPCq60MJwGG
ccUhSLshXGYor6qKd9hLAElHNkuxVygOmZ7b7wXq5pxjCPJ8zRN2vPl4axy4NI0q
CRIf/bnBmBDpCBsZqaFHqa1z8K5UD3gqbGQL0rUQYF5i2CMGjaWobuOslV0Bjxew
tnvB1OqHVLZDMdWqtG6eSjdQSrIv3MyyosnZ+Ly/26JUAFvyxzyCIOv9RclcjOOn
uO349zazr8IlWk7r3okROr+0tZZcwQTrcCrntbpYE84QMCByG6jmDEIYTBvWRIVG
AKUFxhQQVn25rKJt9CMRWn3IMrKicrWAE9gsBSyDGpPKVV6Jbl4d/d3j3RI/yPnY
7ykDJKBUic0gbYHUYQwZZP5tnfSvgakm8prymvIGXzmk2mrh5duRVaW2+RIsilUZ
MK3DgAkHiTqBfDghM6S9/h2ejtlR5s2YKPbDkZKF7m2X6qJh1sGhuMLtx8vfrQaQ
CJdgJ/ON9FOJCk5Tr0cxDpMh0ufi22nIKxiMAxpdz/D2FNTnLeKutGKZ3dkVRGPr
pfJ0SaSPW0lAkywKksiwQ4LIjWTaC4Wcx4MTJabbLVH5Euec3fcyzsCVd94R1cpg
E22/ABl81B4Ks4Hvl04zp9jcPUItvwHCEu/joRm61V6s4LGGLrnj7biSmgb2llbx
A3B3f5+eYXKsFI9T23Nk/wN07I5QGXnT+muotESF9Gi40Dyhwh5NVBikjCW0MYFk
2GjDPGGIHb5FFWuBQxIdtw7Og0pLbDNS0cx/Z+pbot+gYypEXdz//vjGj9Z6spz9
pGf1L+dqR6/zrnPPkpaMnz93dSJ8Tt5htA/56qN7k4GDxK8/rnkjvt/CNwOc7kwx
lON+39GQtkvzfXmVrbT0C5HWtoH8JoOAXThxj60JkiIpo0Se/PBnNU0ktTWGm0OL
QaxrIF0h7jG8ZNK0dIQMGFy24rWHPuIPOUgTXkDdny9WyUUfYQzk3k9ZNxuzMpSM
/FBj05q1U9YUn26BqNT3CoHTRhrCZ8XWQNGo/lSaljTjctQIHJJQNV4GZS7Y05f5
GkzgEGtLbg/ddDzgu71avXjfciWp8S29unYHCB8my1ig7EJYp5twCzfaoKUAjFI/
yuty81EC7/mlhdyW3BcW3jJABMyMzK96nnAWBH14IsttlImIQUcrdemqTdzgkWVn
AUY21UQEvhoWyKpcBQT6tw3jgMDQCZppvlsOxCiFXJ4VKDWkNR31dMVQCdrgE4kS
5406R7kXK6ukRWqpldzOCsCv1FRqkxZvJ3zRiA5CnLabltJ1EycoFFTTlyntJRXg
zTlgQttnLEpPRr0m6XuT315+rCgy4Xfl4k/DSunLqjTP3kWgwsI7iFY4JlLSjQtm
cyH8Ky5djV4WWYuaB43C9SUnVx+F6LAey+A5FD8RSThd+FO3nBAZ6O3QA+zyc24N
ERRzFV9fYsTsR+9EH4lyimc/dvYhURKtknb+BFsYdM+1Wigm2ccZAh23KMJSEXqa
SymQpI4KjOLADM2lM8hlfNoVMbJnH2mAxRrzlgA/ZEnchFjOqZG8EyIs+x/FWvqs
/tkAUcnq7kwy1XJ5Ee2ZZBItDwKJSiSbOvvVCpO9q8a9Xp8wBn3rRHRbq+cJnXFt
mj3OUNbcIEIcK1Agq+Z1ShTTVqWvsG9Uop+6ZabtleGfzot7xg2FgO2lmqAo2tij
TdKDpibOnRLEMrfjdRkG/EYZazM5iX1fI5ah/jt60ZwkGPlrSppOcEMxPoT2eysk
daUN3CzvOQUurEb+Cne403ykehB/HABp/yFXdP9btsgZ7nwrxyZY8PtJDFs6PTSS
09ZOo54LmsKkJICaCMd4DFt9lQQCblF4/Qk4HbSJL8hOz/AwqjdfK1rWtEUvCYMu
hevO/CGJqOSoD3oKc7Rkm44eGTnXNTDKpgccRTA+K29eaboTE3e90o967ZSo2bUh
n7BEndumephCSkKyLRTvOz6Ut/A0AhyvA0T5kllW/3NDFA5u52ofGvMcfUuSoclT
d6VmdKnTosnajxxUyrTyf3wvM0JgpvAbBMBuQSqWHUKNMeJDSVjUHfDz6ROPhPl4
ZKUNSvDtTieklg4sCJDuc27VuhH3EAmQuLn3Y3ykroe3caO0oO1bUEzix4W7KYT5
PRZCypgvXGdB+mNbx0jpKNSlBlLgIbJfjXonVQTTaC9dguCpESI9vyuQ51+NYQqU
bfJtMettfUKIUqIsSQU4e+jfSoI2oX9jki0N86Xfu/BgF77dlRSbAy8p034QXJgh
nVxzywpjSphof00ainyME0RKdy7UM6DSXjAHqb7PbbC33/Iub7U24IRzBQyuNhUd
EM5eDE8u9fmI/OoAZMWB/lj1Wpgz7AKCkz9sf1H8Jy6ku75I5f9lROLG559Php/w
WKHadBEND9hEJ36izXj4nION1Ex48EtVW/s7BseVUa+K8lP0ZHulR3ZI/YCsaAvJ
GNN6B50bWJx6r/B5comoJzFcUt+b9HIBkZVVETOxi9RXigaiQCflt/zUWqw8Y4pQ
34nGmyf6EaAaweCTuf2gZmS3tV6KGS32M9K19Wb9H1+NJw3kC0cVjeIZD2hQ62sG
gdwXtKxW/YtYaAlOhM/SLkaqhY5Sc/kPJHO0jsYddnqsYej4DyCTC+KJ4Fs7l9MF
xBwwtL/wLOEGxW0tH/E9OtzqF/IkxJ7e96/KTCZqXyvvwMuNTujxArepAIP84BXn
/8ceVoSZ1xwJaXSIC4qkTBSYgH5Y1ikxv8I1ru8QSstBNxv1VA3XVXz0l05GoeYX
IEmqJsdfag6zFWfzliIlP7rA/MkI290A3bbmZiblXRk/iQFr6inSpDfE+Jg9554e
GAd1UGYBeIEWR8OBrNeU5awsHvnlsnLNXe8YFNfUNFcKrM3CjcYiph40T5f3TUah
BtZdTlZkMdEPBeFT7se9Duld6ZjRkmYvcnQWKJtelY4iZlf5jnuV5fFgbbBEVKZT
BqQ6kCuH6xlgps3VyDULC3VWxp3hXAsrPdjEckIwMKSIUok5JeP7PtI9/ecXLNL3
KAs0WMFWlFTxZr9M9iEJaev0nWHZgRS3tbZsfDqJ8oqqaJj7D9Pv5q6xi/Q8V19F
8IKRBkc+BWQ13PIX3+ETPrnrn90sws2rPeBDddf3zDNd29UTgYThqLJ7aLfHrCiK
CeYaoABN1KgmaozwOG5QLaYTjn0CfsTRfsmw5dWEmXQ6eRekuek03rrU50jTLZgd
UkmJV2EoBXY7DD9iTY4tnlI0m+aZAfTw2JLh6UzS/LszbUyKyj0f8eSMTfYQlwy8
hAekogJnn2ayJ31OxNCd5k0QGBcYhyPwYeUpEulmugXZC/tAJRLO4ineEjy9F28p
+y/Qj0PWIsifTqaUvsTq6x8CgW56+g42ij1L0AWC3pVSvI5GXxolxMiMnSpdsVbm
+fZoDvZLsHgifVewi3CMtRKh3JXHL4vUf32Odmz0egglJHId/IUUURG5GAT+Cir1
hSj8xTqMvUW4RGGj0LBRBD0zP0a0XL8AKwXv8atp5scXHDx3uLiY6u+TCGq5/vPX
3zKzpGNGU3I8GYwFeOaq1B6FBCL4B+/cNRZLRWLfUap8G7ArjB+gRA8VqZG8QhEp
wBOqmYAfe5ycPSsd6i17fe8zvScZHJf3QJ+GVsBWAdMtnQMF848RX3ZUvHX0yD8Y
CSVljQD+KeeDNhL6Qb2btx/Qe+TYlQYZ/ivcZvLcFA3k6X7u4/ZB9fyOkrC9/kAR
oer6vf2wKr0lt5SoivXGfOpVPi2QqR1L64tWng8Rv0qVmadZQZJ+TLUT8nm8dDNC
n+BYynhDRIFY5uhlaC6iBB9a8N8LHZl/CINtbqXdsOxHEQOegxLX7yQtUHfxlD3e
cZ+SnMC80G1XRDk7J8Kwx49IQm9BXbmnoBA23Hqe4Xf/XTStM4yQfMc69qJlWE+L
QnfN4VneXH+ollzitegtRcZixPV5i0zYgpnIolVPuqV+SP6BEb4Z02o6O+V2bAZB
Zd1o6aUPe4TIH86vlxcrRL4eyZeW6nK2Dsv+L9YFCitD1EtPUUbSEKDj/sWUXTLO
yxWzSLuVN4PFle06A3YkE+qpkzH+jdKvv9AzHBdDpl3jIlmsLTGkzHR/Gv+1k5Wa
cykU7cUs44/hxfPUjV4GsD2KbXCUrxYzClWLRLE3YtdxOunfbZW0xZnDOvNkO2Xu
KJT+XTZce2TiUegPvAJ2IFmfw0QW8pXw3DczCGB9DFC9j+KznGWvZVSBXNWuBc0V
FeU3AqRa3gsboKV8kgKsmLrWCGqS8vx/oJd1uMfp4OtiB1SSX6MAjV666ovMPhgP
cjxoW/7xrW20gL/MGt8NIiFOL2zFWj4o5xe+SlgG3PZV4XYi8Qs7+ay8GE9mtN3b
gl0S9tPyyEBzbqifd1SEzGzYUZTOCvdYjnhsbkkdzoa9nDj2k11wGAWKS6m0cX9Q
wOrIbJH2GTvmh7HN2F9k4Qs/h+uh2LCzU6caOgDQSDybpvgbZ5pCkW7+4lY6Z/qw
NoxqoUl9NN6sGDwHiYMLsmVXPjtwG+cuEALXhUN0a+7T203wHRUO3T0aKRP/wkYf
Xr0LwEefnwOXJLExMprKc5i3xWH+wD/OdfG0820VjvjHnmnEGoiVBjFdHJ3+0EbB
wgf3Oc6ZTgfzkiC2SMy2ONwkRZ4rYikcRpj1+ONf9Ls7/F6Hf1DokFF+xgCLj2G4
kkwKq8AxZUAtlVeeQA+WU5lz9LkYhgzM+rg1wkt5GsKuBXxijpV0LlwFBt8R9sTu
2KawKAla70EGPy2wxvGY1/MgmRH/XyY2n828WcK9PCZ4SBKYH0SUpj/F4/q/Ge4r
8HB/MlRyvxiqMcpVlV16D3QJd1pgC5BfdVMXBTg2jp/61kwEPFelcsjXDPypFUt5
SGzL4VTqQDEgMYg3zAwT7wOtFdjcT2bqwYGRRTC2PR7BFNx18J5kms8IeF9iK5bb
un8ec1b1T/J6hN0hMOCzpgMu2k5v/ev2raQ+uYqrrtYjZcnxccJXFSXQI59TsNxG
WK3f5VrBJCKnMR/3TqOJizCvPVsy9PopF2dgNxFLDCqPG4TVkSkBmnO46yHi/3GT
wZb1gma92gDP+ndkAUl2qIVB/fvHv+w5/O0qsTcQCf21mxLNOuJ82hwTsr/DLBVV
/sCZJFYGoWFRmk5/2xCi7cB2UJPQ1dseP4ykvV7fTyCmA2/d4CFnJSMm3bH0CTk/
0FAJcHaIp7ypFBVELCI9NBontHXOPgcSy4YIcNgWGg0FRAXAyPQUxE1evfmK/lAG
UwpaVDEGMtRxKnYzpk73PpUujOF/qYbtm5/1ue9bwU3cn3Bh3GViP6iB/KqSB5Pr
bMkTFP7OJLgXHUh0ZV0MKwvroEJ0hyRDNvrwEV5N0TjJFA1if9RJgn9oE/dVbAR5
HEeip0TipjXblKDxrkb03FX/6ywVkm5xNzI7DXScWa1R2xGs100R1On4LJp3uYt/
0YWQpGpAz9473lIQNhe4UVHcKdFOiJZRTLc+B0zVcwBKtN8ZrGd2PbmOk9bD3n64
V+H1ZUsMFGXQPlbHCR8x/s7HMs14QyWCB4eXsdIoqxIiUm0wGZWjTIpmPja8mhJl
vMu0E5LgnlndUFeSYYKNnuTnTTpu/5VzVHywcS0RfWELgGjnnDwFM14czF0lubda
FkLSlH98FgdUGhKaZy5YuJpnkvLHbon9Q8fYPU9JLgUhSZOFMOa8OOeIeWZixScn
fHZ1ZYPOrFwV7hxs+Qiecv92qraTRQcXwrKPbj+z2kVsDOuVBdFQJ7jj1Bh1Nyc4
P6lrrwkXcWFIBc28smwfIdcPwBsHql2X5w+KmfkyuZ5Nfntx8U/MQlmp/SNDsQ10
5iMxhewjB3oS2A2ylMK/XXCDZ48EWZTCwefDFDOddUK+FVEcWttM+cGtN2PTmg7Q
5Ot8FHyl59BEeB1L/kHuTB0xxFHbEB3kgWqaPoMJ2WhY+Fs5SU/86ASSMmni4W1J
2LDfEWQULyKS72NIQ7U59eOBCv1m6ijJZHZ1Ys9dkeFNoIfOJa4p855NAe+//J0a
b3FCNVPzmawLlqT2LalMPSAy5RB/8Dzne4/QiBjtCa6ybQvyjP8Eh8hQ1gVYtzJE
B66lBTZeUD1gKZbj8A+Ule/Q4IpgqZK2a6C9PwQnJ4zdwqNySUVhN3f4j4f1LYXq
exxx3/lLtqEWDFJ7cfUW649FBQWJKcpBDd57wk5seIRMRyzcUKeSqyVZBkRqOl2l
TPKeOM8twDJgTwGUUSbiLbs6F071fPT6Ulk69E8oQA6RIO+4EizC+9LSNowJwnoB
MnbiEmaFgmHsfRw/nyhKw7skn6d1AZqc3H2EfBh2MvgUeLhW4sJof5e3bwShha0p
Jk6CjTwxkoRZlDDNiWpLeulaRljgCAiIjUiAuxc1MJHns/jQ5w/V+ZU/hQ5znPyW
iMIRYbNSt05Cc1ggxaSjNQUAGfwTZo16C/1lz673XI7yFo4JmEC1QmIG7l47B6wp
YKy12n3K6Jvs0Oiyd3M0aDfQfFGhGWuPPaye/F9E0xnta89qnMNKW9+OpEFpKYUL
9Tk5/JyuFfQktDLmuv6fc/aT2bQwx4iX1APAfgheIHwdCjDx3ZCHGOth5y5KZv1q
/Y5MN7rbl/4WXXEFZklVVTFJ8oplO44rdhmwHW/HOQKe1MGph2DRGGXo7iL37kAW
m+5tUu/lD24ocjA4Bz+c0ULII282p9GdPFnJuoo7Sw+5hXJ8BcvErEuIdHrkoh8Y
+WAM3quOwovCYzoeNSWEANGn1ijQzlsRWRIHxx544PJ1oDvHeMII4wKo/plYlkfz
lOKRrEzqRYbCBLQv8f6mlV0UfB7YJz0EVWHrA8pgbxh8/AGpRvcf/EgaGCxb1Bjm
MMOWmnePZAq81hr9+Yxb3axF8s9IJah3oPgOT1cJ1LBMV0otBIlIXQlV9avoO9jD
VwVSLqpACWj7sbyEGJCBEVg+bhbttN9ZtddEPF7LDkZVNFLIgg9UHm0XheDw/OYa
E1pL+HSwW5V6RlEUJeHrFPawhWe41P6XH8xoBR4IbWiPqXI+y8LVJa1aF8lgCDd3
ZpZIWhXGcbad2cCS0ce9hKGX2un+mV6FH7s8HV9WHGlXQIUgtdFVWFmNGl3x2bGU
ubo5BePhZz3UFASJgAfjapIbKQRFuDApyFp/xP/9bNxOAd2IEcCYCFUqSPYQ1fQi
PwLBKWKR/prmXZ/4nt6V0NAL9XTKMrn2lM5OwebSBZsEljmc20e0pxZpncrVMSZX
gwZNjzA3k2Hq4QfLk4q+nSTfjf7TjsEQKBMyCSNQE2popPOgEgApg1kXju6GxZ+q
AuowHjCYHbjj6bcy2uKNSvB7rzfwAEeR/x1erzSQxhrB0q0rdTvKDuRchomH902v
ARESc9/PigIurLsUwdPN8qL57yUFk7x1/4wjskGx/8FnhD3jwBgwY/naCM1djdha
QHoUGneryaskzrsX886Ij03TRNyZpNHD2Q4tHwzq3MfTzw2E1VLocjzYpP9d4iJV
9Om7pLp6lmGAhygODhU0EAa033ifsNb1AjdJ9EkCdHt0EsGIOU20KrBUMQDacjVZ
KyMiS7256FxgPiRao4fEiLxvUvIVfVBWbuomOsk/jdmEQD2iR8tg8KIWtkfSGxba
7t3ngFCriv+WXLf27C8iCZ1KeyvqSgrTYbMZW4zTD40dlQ3Y4UUB2CkMJj5+vetp
07TzslXv9b2CPIhF+TpN56oWlbCzkQd/jrn4oQym3AAszJCuSksQdiZHPBWdV49c
7rf9jxX/O6mPNB1j7vBqySzy8M6KX3g12HZIDYxmEbSqUu52PahKU7w+YyQBApyN
fibn61tHQb4dyvt2i+ezIQDXqejptF7YyYePprue9KrHx2hyIL85ys7jnw6CYLL5
n+wScSIFf9vZfIIaAGnt8otJKa1RN54iLHneVuLuGYJigwhIUiW9PA/RgvI7vY7w
lXkC+WN+4+lEy0MCKju5Bo6pt9Sr16d2MfcTSZ9FGhI7DpFrNaZhM2UPH2RtAf4M
78zvW4hc1nQxgF5Rip5XQqMTMFxAFuLCsjmJyaeHa4ZwT6xf2oLWvdpiKomOVl1s
4zr/vJJkpSP00xlqlxhhkb3kcjHh/Jr3BwX+Dlkh+kWVkPbn6u5bq7uAkJutlPvt
u84TNF/LDzra094bDfd39WzyTQkOZKk78yux+d6XS1iWTtepTcqHbvnSMer6MzM4
pj5c2Wslx6TvfgZPeNp0wwwLgwNsfnG5H+zk1+PZ7ff3pY2ypVSQ5nXqcFith+eB
qW/FW5XbOwGSkk5WOanPVfS2pc94RnJbQsr38X1YNx1g8UsOcvjnNLiVnCv/xA6f
8GmfTjtLRKYX6sKVm2NYFNjoB3rBGijYB+W7XHvW+IydRe7Td+aDsaUXFOwJjcJ1
gHfC3AZiP+zp87iBcGOaRR9yTp52fn4fLoWtLTW//7NbqEBUEplrrcdPt/gxC/GJ
02ONC6wZahaQedBufx96lM7LpGzYsBH9UNAMXxSrsTjhP5CiKiVKKc/9lhHwj57P
qJHcUuqCiCdh/iLseioYf395YsAOQ3jNCLVDFqqJHwBX3wBpowU7aAL3iFNfTH5B
o1kIy2WPdTjn6+hu2LqldnQyFi0E1gwPC2gcDCu53N4Wylp76f8/O8LaWeCCJW1G
aNLo5SHA73DyOacy3+AEAm/xgsHB2gqBrGTzaJnU/U/misGpR21ScKJBGDVcOSrm
ZPzXYr2wlx3sQXTqX/ZhRYNAjjyicY0jXeLtovAVfKMAuA/5Gm7h7wSw3/5iNubw
uXiYIkt0NJeN5IubHf4qN3dK9otxuyInrurmqYKs/bTMXIbHrPuN1PQ4sKWPEYu3
bi+vqMK/s9EC2gsuHaqW7gTaRSLqfqYunh8OZaFlQWXAnhiG6BDKO7JOVK+3KgPL
SSXiR5o2QGqASuqyjgyfuP5JpDx3aDPAyWhKENmYGIlg5FP25wxon42HAjofbSPt
qVdpsH3rLb4zeZTAM84Jtg5MYXKOKY2VLiCCxsJDo3xAww7ovzKhoLmMjMBKexyF
FACHWFvAeJXeyvvsKisvce+oC+99NtzXWqQ6M42PYqztMoSG6iOLd1VtrVB/VRCT
KK/JWBHg1lCqWtoT/+5yJwX8OwE31Q35yRWL8Hsj5z6S2MhSsHXYfyrgZ32mpCvZ
PzoWkfne+K6Yje6I/kaRcYoZWOT7eDn0JbsbaJnJIcICPeDEMYIo/FTyI822RuBE
ppMi63nJFAJj8d+PgXvRD38h3OWkWKWlXLPBpeiGTkbGmaIG7mowOuE7Heo/qw1A
pp0vK+FkXbG8yBl+69XwkrPMV5qZiVRKxC+SrACR+sJbCOiv6g5GfYGDKz7ORld4
Gs8+SuUwD77UEy49xXOK3xPp/VJhGq3BOmhw5tzF81ImtvNgld5W6bZoocBmu0d9
J+7DRqpcCmRwC0Kjb/IvpW1jYF2wupFSTcEEf+h/Q2Og2Dv/sRRrvLeYyh+jE+QP
YOFO75WnGh5maSi2CBRG9QUApRGv0D2YxQfSs1nXSQ+vlOfKiigQ2acfhSshgbND
fA1pULu1AuZGEDzeUF9qOrNZSmlq/Us6jCjnLCPjhouS6kluL2fzBSPIxqZsZf5b
ffnxWRJOrW7l4fqYYSGEdpkj5YGjSehN0HHBQgrXslG5drZGt7QNybv9fIrXGDfj
4ds0FjXsAgCpCtGVDCiAnW7xayyxJcX52T/HR95YT04YTi8R19CC96G4r1c5Fg3t
QRfbJYdZPpwCBBEPN6Ez0dO7d5L9lp2sSSc/9p0aX4WVHTDoT3ee+y923gARtfeV
9YAmvY/lExAll8qGmU/3rnIUuS2Fnphabqh2kzW/kIfW0xSTwTbImp+xiAB8jSn6
nUMIJcE//yIIkfNswxzhFBlIg1refCYe8hlNKfLl5RVoGZoAk3Itbi9zY6yy6/Lw
FUyzF8JR9pyecH3gWhI16vGUcQh4zu6CSR4HNWsbNEeTRpOAyY7NhOFIyR9VAgGM
7NcqN9fNmxcwgzhyTQseLE6P82ucCO7VubAA7ZqB/jC3UvE2f8sJOhG0nrg2dIul
lPc+fsaXwQOJPmaZT0mSRdMtfsHMcIWU+ztQeiNmZ7yysAD+K2r+tmsLzXFgMnJ8
wNlgxtF5waIAfdqQVizSNzzqIToSDzAcsHoADZ0geZsFo8owV0V+Q8ZgmqYl75Dz
ABq7g2AW3DnbGK21PmyNBppXSN2mR5758n5pOVnr+3cb6JbDy44fh4w/PrZdAESk
ejGax/iwPQW/SRZypCvDS/maAPtjsdA4PlfMQ1UOcJhvuPK5Z38zkVemS1KUXhho
iOr+uT20PumpB1Kgg+5jH6tsUGRY4JMvNZHDLJXfhNMuOIt1nGKysakWr1UvxM37
ByOzRdQunfee6+nVPWBfVY8+M/xpPrrtOeSUnez6Uw7AKCNX2Qq7mvov0IgfDwpx
p/VpbaZudUmxA+RY8WCWusTpHYeCHx8elnoWa1L+Jjcvvgd3jOIvcDqyuq6YRwrU
olq2i5QTtQeKzi9uvtLyH88kvDFV+ucLq6wLYyxuepy1Leitja6VLk8xHTvjFz/T
Elxty/xleERxeYN6DINbdeueaHhpjrCuKOOBdmAkOyHu5QfTFzusJPiMTijfdjA4
FTyYLuYV4y4pU4JzeGFwXkTaVf2mnzUNy/d9FHDMzqW6tO2ByHVIIb9xFtNG+4Yf
e6ub0Mj5UlORWhlToXT9tJYb528osQvzhnYLtinxSxPiureqc6zj0xbchw3lfqq1
H9tSEMfhU+/c8IkIMbj0Zt48STeVaIEx4AuAfO6IyG4dM39iJ4qj5koYRPylvgDK
nLFp0dMBY9DidDNWj8yi3wScZhg31HjHmfCVSFOkmYRkyh6M2lQPeRg7E6jaNA7L
50Ps9GQ+mOCSvEKkHkJ8+JILsl5/04H/nyFvoaUNPwDcKXgEli1FOxwhk7EFlp+k
6h4XlToLp9ixFdy6guQ6+Y7Wx6QLy6dFdmwPp4VXasOS7yrAmo78JtXOop2EncLp
mq1yOs7QBOeIcTv/PcQtE5FQMSEcQ98pZQt23c6qydhWjTwQJJKQgn8jZnGsx7Fi
CifBcgkoBAAjAZ8uQgRvS5UY+10f2XzjDaFITI/AtamrNAjCJo8GeWYtHmWRMEbY
wxpsSxFrlI1Ms6+Bi44Z+dZ/LEeE/1xm2jEsfQ9JtfmE6/aGl7q38e4EFrV0YCz1
MfQLCTTLPJWUCrA7zskulx7VLH9Sh3iojn0Y8Q5oxV/vFs7+m7UhEDNyWzMm1g+5
+hUH4/5td2N1WoOJcNFlYTo0NGUf5ZjrlWAxjYTlCRZX6O1oeHL9smWumLKp2s18
pWMxkKiTPhn8/DrQskcqFEV7Mkj9UNCcauSxHiD3wnevu5+ox3HnkEQjvz1J0roR
BtEvgUQ2ZxUUSjm6OGZ4QkPpOGWUC/3lPHQxF1FiOTZbIMOODbkbkcQlqM6yUWvF
tqOOEhYyvepMWPQo/enr1qNTwCRBOqwyoRSKudHYEnu3bVSHPML81Rmrnp4BSv7e
09YEX8RKpt5weFiN6Awlcy7BhjPmw8OD2nCyg84wP/wcn/so7K6ykI/knNim9fq/
Zli3R4AZNHFynuN725S4nP308rz/uhdx4C8kZE0sB3C7lL1CSGOrDpb9ooFlJ+JD
lPutfTOAF9GMPpYpKHaFSthcibhjYoNP0afkPhn8rzSYV5DknDCelzESfZ6wczA+
XqnIzvKhqGKpC8N5xiuOPlsyRQGtbDdO92XmFP1kjj2pcy5aN4QJHNWHdwTWRslx
haxdZWEJExXegPtyG4m0lSA2Gocz7rog//xUZT66yRjItQ+NHCbMnxls2M7n7w7P
YojBs512lvG5DTAd3jLmUh9CZVHWGjj5jZNBVU4w3d74GWl8FNuhEB50Y0nxZqpK
u9de3msXuqBe4/aVWK9p2lpYN7nehgW1Gwqadda+1cy/rah5jGaS6fRhQhh/WR+z
+WXmRAMMmLR+USxXvkvuiUGRxan/yCKHpDwyBtgyXFA02pqvaYG3Hg9uIZhla0er
6F3JkQ3VIhydwTf5+16aakzUMPBnjhFrh/cfAjYhUPYtDGu+ixpmYh+264bIkdkY
pmKO5ij8699aKleK/oZVM+bnwqTtThSl728Uce6ThhV5XKAqJETu99PQrMtE0IlU
6reXnlLiRdko71ne7TmzPQlKX7ObbSAwrggCRfh2/VV3K278wg+b2bQ9W58+Nzxt
3H8+Do49T6G5eoFsKqM2s4YU1QEqmCi4wZtbXKboPZwGFcob7IEtSFF6m3vDPgvE
0xEVryLw72Xb7/6zl90DkWmAHCqUDbT3z3vgvGblhF9UjEeEx7wPIAOhR6dTkMR8
h9YWSqZbww/2T6W9dniYM+1HSoBbMz2tAyzUcGDHB1tIU5gbPwkXjVOJmdGZMohR
X53jafAFy92JBRAWb5soo1UhNC6YMmmUhNTgITGLmQlCYASHaqItWF4hTh7eyZJj
C3aFxFIsAyV6Fk8teTI9FEOkZUexJA+QJiro5n2q3ZZv7bNCfIIxdV9nTXrBAtZN
F/0W0HQEqIS19FUf+IfE8bYFZ//48qYPvtCQrduj3iITFc7FTMV2Mwdb0XrBZYiM
mJkazWji9WHXGg0nZSjFNrs6QywAiYDeZ4YFFCHYRYikWUj6IsqNaoFfrTXKZwp3
wsOYZGUOtJthBLkjUS9ZQgj0rOrilKZJ6nxoT6HfCjDoecTdTCITQuVv6WA3VURW
G9Xs2BReoNqqq48vJK9VTm32R7PL1BgzecKXLsSTWootGTioIRVGh7RRWtaBk0zI
txaaJvh7BwzMVK68uMNMVJ/P79b5x1fVX2v5QzFqT5UewG5RSHumQr7Ahc1UCdMj
WVPz+KzePxFMi7Jmx6rpGqN9PdNKPpAv7+LnKoDBF4ZvofgEkSFPwmbBJ3ZlO6AW
DyJbWqqigfQRCK0vjICY4VNdOJzd9JaN/XipAPCtSgxCNl+/E3o9zcqoUPrGSJYe
agEZdfRCeSyeUNLNsyy8M3jzjHNsUTp7Oy0Mn7+RQk6WNUbWzA82Ze1Zy+efj3bg
Xkf1GIPDWAI5oppkXodHrus7J1zoaHyzqj5HiyIC2UlupKVgffUKDzvw0Dnmeo2k
Z46U4NdUv8o3dSoMbE7IWVhcSuCebOOD3M+R+x+8WdeVw336q58sqHbhUiCT2EG+
KOdQIEXdFwEZPpF29E0/IxszAb224vAtjcisbxqjXAIKHWF1SUPLbqFTXTCWrqMH
rAP/XnYKGd1x8aKwY8SPIGuAJToR2cBNEcOdjMBnctn+1ZcanY6fH5GfNFtdoCfz
MxOODPEtBtNCf0tEvwzA3uye5xjnlCRtE+jYk9IgVOGevxiwK0ukW0UzSKk+vdCz
PpwdodP+8RkJfyHBcYEgt+r3/hOw/qnEdz5Zy32kP3oB4KGLpuR0N0f+lhmrvL4E
pCxOJAPVndh+GTwLnzE1WLZf0A63ObMHmQX6iqRr34TxAE6oWRn5aztRA3N4Qcj4
g+iDFChYnjQBBZmTqaJPAsmZHyOWGNYphTlQGdD/nRGZU+WUHGa7KIhLmG/AhQeK
TdMBJI2EzpXGrmjZign79PHc3o6oS4h8VBmsNtWy8KUWeyG8F5Rbbp3/eJXjZFRn
4qtVKgPa2xSvB9C4FPEC2fFiVUWQWonGRmMy1Bb7kGCOVgs30Dchr+7EC4tFhRFh
vgfFOSQniOREGgOvbPIyqsBS/mmWXtNqxhfBb2TSjOUeBgNtyuRI26dlIxN70Dai
+xVFVEZ6DTrSGDySJ8nFXMxCO6SSk6KDMo7M5sJDR9aRPH4dHqmOShvJF6z6/vFz
odt7Q5zSHeWy6D2ok+X2+B2XC5SGisVmAe5mnZa6KnWaLJC6mo/RzfEGX0uhJbuV
kT/dHIqTEN/zK8sNRzgrovMx4VK3JtnFkMgiiDxAM5XX4RN3HmkuGgQ+YAJ3W4Is
thN4feIpAfsgC+wNj+61T4aV0CSR9bUuKcr9hiJlZ4Su5n9HPZax3egMrKGQTGHa
pGVdjkzUyveaaX69a/B5mo0cyU+PCXcE9/EdCGx8bWYyECqFV0xUpg2LwT7NHvww
BgyOBI4Yx3kdu4mldGIVCQAB/L5ZSkUovCpLHX1b2qpR7YTeTypfHW7+zPwOIube
zo7aqPgwiw2gnCjxcQTuy8AxWrnwheaiKTi5pCSmr2RIA2GSYryoR5FgwNOMjdwc
z0sytY52W+XRp7WzKF/67G9FLfaHBR2ktTK7wrCUYy4APVRLkuwOvJLh4gzRVmxh
+fIoo1VfddMeTKxwfn6uXkYxbmRkZdTEpfBFmwnOCxohgzhur5IXGY+R14DgKbVN
9PI3/YJ3lJWL8mZNSAXQyRWICDxsCoRylfXnfkmxS9hImiEqHkZtFSwpTXTUjZiB
zmjkOvoVflu3tPwqSnBqFNfUb2CiMPc2XCV3irrsTv+STZgwAc8WGDEFAU8+tBcI
tikJJ5kFctNmWHE/Uo/37DAK+AfB4cTzHeJ2ZKfXldERMLisPtvnf5Re5TAiYJYA
Rglw0WmS8IU/qUF9kVpjdoi8PAJEH+rIM8Y35OYtR7Puxj97JsFl9dfUSZoITuzd
WZ9CJ269G1sewctgu6yIdD9fk/9dbgRZutdvDMsq7wmA5IENlczVCE8K5kBhCEwY
05xJOKmTXCYTzMBYrTucYLEA5zpQ+KexTFcKBH10DzN7IHs+4P/zG5aGU6+g6bT3
IsRcao+tAhexQ48B8noo9MSsCJhIQII5uRsfAQKTtHff5CcTZuK7t8DMXfZcO36v
r/gR2jCtsfPouvPfg9oV8f7Qr0mp5epWqWFgXZqHvjAo7BXFxQ2GZwdPVfA9lany
ITESSDng1zs9fMLM4y5iy5myO/ztQx2qCJtjZh8e5gUQFX2hLzmFFxP60aoNCxZJ
Y9b49a9uAqDSA93alfDQgOIv68tdb0P+kgBuMK2XgmI33OJdWuT/BggfMr3hRmCN
9Qk2LQpgR3tVlb5SJIkEhquWzSXtpLq0K7y2TnKpLA0Tvd51ZGeisoa5QSH5FPdj
8vfc5ZuAVnWhiZPVjD4WIyEEtQNYikUo14xrb8XHIyNx9Zr36+n5U2dbtvnK6X95
su4zo+tWQGBx2iEDDJOdW0zgxF1+iy8CnzCxhdc2wHo3jP4MABEhRlGCeorb7u1T
p3uz65+n3zN4XyAVXMqSjYdZ/yJ6cFXM88raWou0BHpzWk4m7HMEtP71gVcJ3LYF
ny6aRmzbg38MphwuwAeLmRoFT1SkplygNXR01SQBj+0sDU229ZQ7E6aOd750aE/C
h7xJX84kOntcD9d/sVWEsAq1+1kCqJagg54MVUqsbQ26BhMzjwWPE9yMu9Y7m9HH
lUAsgk66VsJLXq40KGYXRxs0HpkFx0ptLeLF+cXuE1yPi7wyIpk0AHhhUxqpdAQZ
Qs+J4cPR4kzbZ+85Q7k14Of/qcOX9bcWnXtrzH4lBbfUXeLXsFRmEvR6NFAuh/3D
cZFKgoZtgjYVH0Oq5wRUfXPRg012oHsI8SgmE3WWDJ0O4aA7P7NThzY5gdgfeFIg
vDOkN2u/pILXjaepIxY0KdQwqOqD6B6n6/kyW9KeRjwYqOT0XCyz70fLM3SgdfQY
FZHeLvggjUr9ddWlevTQe225c5R15vsNJL7x8fD0eWLro4Z/BQ/uB3JGGEmwNxIH
7CPyiMpfjAyzhAg6n4ZgH9HmCtlfyJ7LLs+Zn+IXXeY/c4SkCCiekyyMqoabmIky
cu4Z8LfIJ6NVOuzfX2ZmpxL9tTL9P0IE2HMIOH/gxH8KIabTUuSV/yv86p+65khb
z34+u0raDgMXGAz/5WQdqxwS5w1+/iFKjYHiZbP+iVSNrxMuVFOBFNUhr+A2lbwp
9nXojckbKen37JpHfkdk38dZXTBkw6fX/KLFm9yI3oV6iWfLidB5pv2jMBwC79Ai
8AR5dyUXSV8qM1Psmz1HyYJgT2S7qdAsVp2nBrjsg32ONLd2lO3+oTLzgK4xmXGi
Cjb/io96CxKBJXmcxpS0dTbpkGqx4GapxUHnzwTwzgLu3Dsvknu/DKTApZ5OM5Sa
LYn52/sM9iOcsAbREjOzpBZdMmbLc2k3BSoZ685kmXvaHomZgm3MvKFaCxXj20Hh
6XFwKad58BmGOv2RTD6YMYmKrwolSyVp1JiEHufnMy77tjwuu4lRam/p5NCxIjei
CGlSAHY8AI9JshyNiMljpRufDL3gJQZhZHvqGsR6crZs+QMgcoh/n29kHvFvZJWB
WTHTVZHDu8pk03ra/uLGSRA+YEliIJhvBBpIS0sNfGkGbJGA2H7oLTIru4MFj1fd
49qrGKTO+cwdUWXJDHUJXCnY+Z665ONrqJR/DvPtFJtVCgjJ3737Rbgn7VxdMY0g
OKDJfHjzoyoZJd30HbVp17JYnWibhUFLiRTzRKv+zzh+jdU5KRrhgEOuQlo3s7oM
cWlMc610j9hVyTRnPWGBpErzdCJoSLKSaMHwYfoB/wAZlV0och1KsmCZsQ7d/bpp
GQZxoKUUeG5N24qKG5gA+1GnlGWrUfWucHi+uA33izbne4Ceq1xvDGO6qTVx6Lx6
/0hWI79AKTjM8Kp2+U9QRVwo/p01zwDzQh44ypvFy8IOF2d2nNd0WbGbz+XKw8X5
NbADgyyGZM8cX0QePHa+s/afGkFuRC7rmSAAX8Gwj01ngTZsl17pK7GEMNmR9Rxk
wqWs7ksncYWFRfZYK+JLpgjVRNYAQZgLviQRBKSlbbgDbK7ssNHo6qblCsn77t1q
hfecEYcB7wuM9eY1ANRfrP33yreCFubsXjv8fiEctxgb/rCZtK6s+7t+YNSkunKu
Sy2LZzOd/GEVOCX7osLLzS0V/6v8sCIfCPAy0OCi7Rd/BSP44DSO0BfCN3WcOE/8
VVgm9GeqP/JJE06slQLe6+Mv/FfJ7+3FwyPUXuBY6H0fQhBKd7lMZwDI0ZsRRcIV
AJ9rhDkrvJvt0tzP3nakeMcq9iVlZyghOi/cQX/Oc/f1ZOB3XVyljAj85NYGn3wA
itpUdgd0Mpi5j/nHwuegQiPOU7lkxF4jPYE61bQ5hYrfAL+Shfz7FTQaj4IGM7Ah
CoOOZm6iI1UE6UIGNKqZioGxHvVCImznuiP3a0vEwdnICge2d/61eM3TO2CBv8xL
Few336I50p9ghO6DCJA7TiIEox3P6QmRpOm/5YanQMjbTlGHciZ6fOIiYAkcuJua
cFjPIwPJMqoeX3VaZN9kc+NnLLrlVHsUNA7I3WSIPwBXIn1Tu6QwBzhbgfSI4S/W
2ZWIxc8XHsKasCbbSZ4ljCOTnQ3IUCrsI5BEdhQx1FVjXRhtrFl6PMD6w8SN3VW+
VIzwUAuNuLjMN7imUaiz6zSQblfnSxuNto5YHwDauIhJxFACnDURAioJe+H1+R+u
5EZXh8SwvF12stV3yaFWzdwAn49VhRV3GiG+QQQ4CCTInTACbL9NHZQBfFtBNi0w
WDQ9tN0ynMJ2xunXEhaYnnEzP1D/FoQ1F3Fo8pgvHE9R+fiSJDgCwifzwDHOoEur
VY9nQ9q2nIH1+WEoVIQ6mY1Ri9zFkYWT9oWEpI/ARwMSpJQmi83Lmf/TkOqrKKE2
Y+8ZLVQPwbtGP+Ltc7LGFfdi4zPbB52aikTsh74CEwEWu60Cpl30M1BwM6/E52D5
+R1i9UmF0ZOJzgaK0nWzrrSTH1eJ7vteBahr8fpjLtLbB/9Mqd/niBLv9Dt60Qnq
8e6B1y3AqA+gVnJDD0cxaY0FNNRiaQk2JX9feSr6tMvjdBjPWyPSCsJLFeibH1h4
rAvBnTc/cR1eCVlLjAaMVkCY7iU19PASpWCtdNHrabYutQqHwVwZQ6fmRDB2PQ1d
GONsRv57ZoS2IQpHDPcZBJlcsqRpHuJZZDjGhMKe4K1JniPaZZT/6Id4Or/9btCt
yHDmm/AXX9PyvZLUxFBEujUur9+8KuU1Gf0F9G0SbTjIrd5ELgNlrEgBWsCDhRYn
hTEPp6E39a323UjUcts9tc7NDKcgajGvj6P2KZ4FjSmlq9wpudPgAbabhzx1ud8R
ZrWCrdJdy5a+lMDWKaYyzVKdpqDa9/HsUAU8ylG/kYm/XO7ovQ67rMD3dkwdVzEP
4Nak6aWq9Q62n0uYa1zEMnls+a//IdjMsWa2Kxt1j1kNNTAazyC5n+dkE2FkpYI1
co8/DMrbBOL5oFq+ZsnctCLKxiQqseUhuYde9z2GmEVsQj/pFxfSDd7doxpbE90g
YnusakKDHrE/AaQFIdhUqTLZLvdtmPAJArAzS4/4puz5wWvkbd4ytKvnz2XWb/az
uDTj6Kws8bV3H6Zt6sFF801eVOAe0PqL2YEhezvMfDrGnIRa0NTBybpzUhNlWIsQ
XLNNPbtT1gwtYxGRh5G4eOsr8m9pA/ra5XbixP2DBCgXvAp37WQX0Ono+Gpmvc5Y
V7CUw7L+gil/YEbUwZNIWKeD6BjIZWwqgIcMcWMeb8R19zSDlhih6ZCTkcAbO0jq
JQsBuoTYoiMIDS3wKcbFZBAtw1k7l9KKvzZRYbh11ishoSqR0m2v0erVjlgNPh3O
SGq1rTtGizjQ3J5xzegveQpN8XiKpMVBMqAvLPWA6Gye9L5eXoW+dP3XLTSxbfgZ
YtjnUTDnimrsiafFOw/oVbAC7g7gMd392kJz2Z6vJsVWLchNCUsAEkDlZBQpgEEc
+XAstt9+VyT2UdiXO3+gcu+Tc/UIfkJ4dLPuGUa9tfgA9oWfMO/UMkoLjVcET/DE
rRYqrguiUGG92cjg/y+MVYooJnXBuf2jkM1AAPZkGtXXLFXj5CEdWwjJ7O4qte0w
E3eXs3n3FclEEA/qoWbdaub3Kc/1M765NXw3W24wQZoqHf+7b8DfZzOnBeeDGSAh
tcALPtxRV5ABb/40qT6KVC3V6fXt7W+NEDS/sesb2JKj6tS1GRjtx6dBH6JT3eVW
n/vcpc8Pm6bl9x+GVawKJZLc4ahKT67K0kEE+g6wqfzW01tuSiuKDZnBljS8DK/G
2jfU6NuJJvuiHWvdu6vBlEU21xBaiepbhBcSH7KLH3TguFnd9hm6eTfL0bRSg+RG
6rI6G2xE0TIUXjGsEARwFgTw7jSSR1VG12/P7egwqzuRn3sFcvy4hGDHiCaSXHxO
/pDVOTLT1U1YEs4SoSPUile+7KcwmBY0ml3c2kozOQiXuhZh/zlHmEMRt7XMmdGM
9ZpL2ou3Kik8Am8XJZuCEJ6OTDFje9UmTrYQH0pM/2Y6EId405Hd58FlxiMGv86P
bcLTEPy0siQfy1OmsP4yWJBPIiPuHXRw/DBBXH1vKfjHqcdf4+UshSD4YmiV5Ngr
7QTcgYOUATLHIJSLqwKLqG6UabtzCRNdF5CkFpTDomTW7GeV/Ca0xAgflpidPcXn
XsY/BSpH+Qg39vlbhSz+7+xoVjz0lOIJJNmFXOOV3v9Zd77Xy4rTjECHfiORBnZq
CUQ5lVFLvtzMlvR30Bj0OklSIib7XtEwrEl65U7axqtyjz27KNXW75rZwrcISjdD
0FEfGA9qhwDHrP0G96HG6kYP66v4F8tRUlNPZzfKtcSjGAaFPreKPQgVHRdfKYmT
jrKsUnFUBo9Xnipdw9zguOC2DgpC7WtuQzv/x3fC2pTNcx0ulVIo2hrdbHV1ZsmA
MZRMZzSIrsi68xprAQfxFETjBcfDslAraccjcXGEMeh0wUMCG4+9xLHsL9UZ3Qpi
f/loL6NSuxkTm7DwOavfzI1tucyffs4ko84xSBO1swHHTe2wAmj1W9L8VP90ioUm
89qGtDRaOMlqcudUPmROYiRpbQqVjEeRvS6+q3YwdMOLJxgh+6KXJmhZWud7k7Yp
yC4qdoFFnn/7JMWaKIMDYedP5uJJfx+lCbL1/RPN5RvZxbmBVsHBZHnxKPIcYc3p
TFsVZR0MWx9jh5QhMWF/VdCl5SjP9yd/L3KlJrqf5SIFEPmmwNpwtUd38hj4fnw9
FZABq3VKwJNdl2wxTs2CwwO2ZgGqc3XXKEagHa257aMhnPfezNp08gldmlqOOJox
yCM5c7uvMpL7ZG/bMlZL4T+9JquUCqFASxlWuNgbEyrLMVU98vjONCXBfx+H2JX+
noG6dorf7NOcEoLd4ijK8tzS7tbu+urag/ZegSEncnwIDaCuvP+VL4F6B85kAf7x
2C4up/x8FGWo3zMUzY3yIEoG+o/Qdyi3hJ7QxpYKK0RWWrOFKUX5NLA1jTKYg8Lb
+UQdgIklMZYehIs17WruOCq4QyJgWGAcG5jtHhBI94KHhkNuBsDUIN2noMJwfJSe
g+Bw7jkTs/BckV1JzkIB/dzF67pLgftZ2uS3DSs+Tb5hkxb2cU4c7/NV3hKe3U4D
eXqk5HuD3SM2nIpS9ZECMJio4jy5MzhRnx9a6mnXVFXEzC4ry1z12w7q0ySqp2Ey
fofpB72wafw3A/Xloj91iOMcAnq+Sh3Asp0c2YBXpWb7ovJnggM/RIs+vHDCec1k
5lBS99TPN2Phw8+KX3SX8lUC3J16LSISlFDFDzfNz/GU2cOaF3xRYCAZgg7fgStO
aGUjqZPzYabOzOIXP1AaBXolVpPd5Oe7N9pQzz0PR0EwL5pMjpE/fMHtDKx8vYnU
DXFcarFWFT54z6HZ3hWASaxVGd33G7yULs6dntsLqdmW0FUkh3o2+v9i0NySet8T
08bAZyjskf4FYbdZ1suqu+JLzDR29QUjwFX3AAN/tJotfz4m8Nx0jlLQxU7lPxd9
mjiAPBC+xarGgF3SOzdK/96faYLeOjG6wXePXILqzylIFuiwu8JrZBxipuGwFj/k
GoRCM3n+cU9tbvz3OwmQVwF35R8Is9Uos7O/VSi5HV5tl8NKx8fWrSARS1j2dcg6
C2TOzYwE3hqn1GJbKh1CxlrdexN0/b+nbd+HppEnlzIcn0/P+AvpWwBPWI9sEBXo
5vB8gLUDy8NPrcG75daA910kWIRDMwqxOA734aFQ98416l81D0X0D0UXES4WrZLn
0+urSD9Rq1No5o45JrHF7fShxqz5mr0hzoowmv1h+bMwrE6Joww2I/OhDtz/8MTR
H1ywqU77ubS+ZrgbZDpSlg3p7K3yc40w5SYSH8zqbkxM61pam6MctsDJCKV1B8MX
YzqL4qQPlb2Iv1lWANRpz7fMUSgRcgTHAMcmuSpGp3zPSWQj35QlylqxaygYC3jo
MNDs3bj31TbhGjNcNWi1gOoSjw+iVlDbZUQgAiSrhhFX7+lOaKNzVAvm6rQvaU48
KcpBzHsMfhoHBWWqsfZ0nTfNLHx5oM22ZsmXRjydUt2UCdmpgCPBALVkhn5k1GIj
fWdOskue4o8PoALI5YoVN41NAY19K9CiIs1yxT5SmVrQCWhg2ffyG0dniz0PrnxC
2CGvoisG66bkTY1z261ytUJ7SPbxMPh7xuauE6jqaSCPMDDFLKu+AHc86ES+/v/e
pRbHTaNz4oPUPlxxnO2YDJX+hwr9J15ao+ouRyO5fVrIfK4qQr3Ihu0IT9APIJ8r
6bixWCi9Y1mHJs/G++hypiAiB5sPQagnNixaNEEqDPJplWM8DUczilR/NmBXlpay
fBFv4rSWLY/aIysMQeWSJKFN98BiGonWceV1A8rFkYila+C5zNPCmbAlMCKuQrq1
6ypXrnQZQHjpsfBrbBcvPD9YAwmIYq88yUemBBHaEYawJu9sBeJTATHPz3uZt1iJ
Jbzd5LVJSNxVNh3DLsndSo+SVdpiPPmm4Zvr2/kIP12c5wSLcwS59MqOL+wClKBY
KL1jSVtD7EMoFul8m+8DNEKQ4KsA6s/U+d8h95imWxnvuIaVowe7JGfmn+dq/qT1
OUgIaGA9FEVHsP9KsqyaZkAm/FdPbI3f4F+w/rU0HrCRYEFgEIWBAFaBMlVdl+a+
zEo5MQ3c4kLVlhENUTHF53uwcqGjCuee4RdJd/dhv0huxmu758Fm/RS4axP4JK77
Uudy1zO9rw5sp1Hr8TtLHzG2eV8uhqtT6mw/lIwEs4P3NXSNkKW+IPVmwZJIDz8F
tX01wz65dMFhjJAqJZu1bDp2KbVYd2ZElQ52Yo8aRJS08hpdBvzcdwDHDovwKV67
c6UDJ0Ti4Hh3T5NOOoBjmZZKA70GArWG/zTeX/VzaE7ERQnIL/V1oYqdIRoU6T+f
AUqi8njiVG/AunLMN3Auj8rbYK3zrU4Kdo0xlW5nCN5M1UBSB75B5HXVf9P7GOZa
yeHCLBM4VPx2fCoKWwfulboqYs5BjBBWg9mxwO3Vfwz1DokFWo7/0llkPEycmt3g
iq2sVRR99cpsXczA19dBS2kTonXqMxdx3wg52j9zXPtOSAQFULcUhYKtZcwwuZuL
0C5Mls8G1vQUNMCjptQJV09NqwDpRJx8sXD/FrZPELMUMKTYksjTeLUbAg++Qzbh
tyUjhN5Zpn31EWniVT4i+RfM+bK7mQJndnCUhhZQXOU5uOxftwHuJlmy2HRnsSat
um7dPmIHfuFOith5QZeWfD1DmhEnWID25+uIYlqEbjmRdEk8FccM1xyVxD7AKkZm
JLdCz9aMYDKw/YyvhpxVU+Gg32hOdTzYolN264fmXng90YPQvf0E8PDm/EJyXWSx
BFFpYeGQE8cRF/UmeHQ6DEpNYdSoVVKkRdDoCxFzQYFY/UtsbxwPAPUW8wmijWb6
2vhCiUt66Fz9Y0oUzTr2Pt18qM+RVD0NzGFgaCO/g4/uI2rXnnj8YXNYLCMk/YpV
Oh1PzdM36wTtWyZwGKUn0PFiw9VLPOMpWXNpotUm380ZyEnznnjjSrqFa68nv4rV
QlPjsI2emhmcr3vd8joGByU0Gn1C7nsX5UXuqAIJMs9KBC5cJeWOme+r1UJJRi5a
R8HmmhS7FG1uyavGxKHcPODqAhqQWEz+GgwKOOVTi2q3WLVjDQyfvNQLHxPQtv45
5lqp0nXeAM1dUMoEtLBCbSXH3iuBNOuZd5iK3dEzZvaFBHBeLPWbr6KjZ0M44t36
/MqW4l152mgmvZ4ESD0nh0EtOAqta+0wwhGeRpzn4K2aAYOpNJ9bmeXwZtHI2BtK
84EpDyyqrvtrnATrc8jxk5ZiOA0LCN/52nIJRM7ZDZW7smYj1bUE+5OHAaEMyHYF
VElkknHAbJ6smQsg0zvfqYKkaMbH0jJDDWsnNVmy5HAPNQLV3FxmWtZXzf0kTEgC
oEH8tfRlE2h7MX5Mze62Fmqoei/Nhdu4r+bNaRRlobr/MwFidUgOjOuZvw5GMifr
xX0JXL2YccHqeH664OH5veI23+oe9kHwmibc+H5CEQC2vbkKAHhi7Z7tM5UV/tyL
bmsz1GJxqIAmFxgfr6HMA5dz422xUkmkHOGDML2zPLiPLEKVDtqTo+yRJ65psWL/
G9dYw5B9OZE9RNkE19G8up6VuVw/rRGTW9TRwXjSq5IXJv6QTdZ16krn9x7OP/QE
5ADXaor9DG62Uaz3Iak30CtCjQkNHNJbvaVG5HXI7sd7Uk5PyLJbj24FIVLf+Jes
fAU67q/uLC2hSlowLrzYAnKZOEq2UZwngIi0zLPVWhr98Lpv8uztniPOQZOa65nQ
26o5EwXliEbhVgFFuO0DcBcLHmgvNpW3ho8NUUtV8LEsyEQB6wcxKYUUQ0JDoly6
5FqPjYsA2zzfehFtL9hWIJEBF/GPFaO3tg4FmGBmlSRszvnZRdMqEVKlUGfOOBbF
yx9B2weuNBwa45bqvUOJQaiZX22UbjYWC7oqItULJgLl2XYrEK3qr+bV9ri2A9gu
NBQ29BnL/Uc9Fnv6OqktwcjPiOYE1ysOMLvfe+Y2ojbFPTgmp6NRQoDcYspnHBEx
ZvmhX60YGCaQdSTBCK3NONawEaofQZ35OHdTafpVu0Gi0cz38zjBciPvvDHKbFIQ
F6Ycwka+cl0MqguSofoztBdUdtEYtx8sVOhOvXSvHbMOZFXE6yPk/7m7GYVG0YB4
RyHHfe79EBUXYeeL1casAraH6xXTpGu28SJDR/rp26yxvRd9ZXKiBKZotFD3/B8X
iDh3T265cHygKFW9fPWybnBRR6r4mY2mzZSBfX+I/It0gUKaCHZwrNd6JC4bdkDo
Quf2yJc+gtIld1ouaiDdXi4Y8AWo7gIyOGdTNCUHNir3K2LxNyGrnsyMgzNGXNFi
unf0eQE2I68W+/cDLHiBN4M//fpXdmAWAsY+2njFjKmr4cPm6muC7AeTXzKpt7bX
cF0NL4fFddWtJeZv5tVZxU4tZY6zxVShW8wjbheuup7a/82O4RQqNea2k4Bonyu2
y4Yl93CmsW+2lViAcJXG1qY3onSoP/MAfK008ecMARnGaoiwQfS3mfRD0K5bDCPa
ZP3AraycTHdqQ8vxtnG49zghx+JpAawEbAY/eYOLHGGS/bHXa0vQQLJzjzYZyAjw
soIbd7jdmQNohSh1VeM/l/FI/vJu+WzZiPUrcSj9xy1XUkJItG+6LPVYLlUuvbjD
VNEjJ2ZGNQZ0bQdnHiDZz5iFLKmnAQeLqAoSXdu60lWtwjSfzDZsTCVeuxdDbtNZ
RsCBMzj1IwbIyWpiQWNLGLEiWniNjNUm2FTbmYH2Jq36ARbF3cJOPDL6OpEhsqiv
5ghrL7gpUCZqyGAc2qwfT2EwItxEciH5IULwvxp/epWto+UgjTWZBQvBuZOAdmYb
VQi1wKbnldyyeBAVTqLGL5iStIkyYMUW/IXDdgUjAT36SZPUXyEmzGpQG+nGwuxa
TPGISQCVKMgijgPkP3j3CKC1bW2fRkj8drJKnpXuge8m4bhR6FZMdXXqe0hIw0ER
M/4SCfInJxHFinIVqgQWLFtziwOlrV1Ro9V4x6sYauoN71LUHUCc+l6GhH3/lKts
cmolDsqImHPnbdGSP3FJOUr/53MbvpjIYLUP7jyKbD032C4phfg3HKUFbHMPx9P3
zCoiT9Sm2YyTOeyZtmwp4q0AtbfROHGCq9aO08U6JHlV7z7pQsr427j/PFncMGeY
0M5M5v+r9bU/9mR5ffvPY7eu4D4mGJ/qtFa9gi+jdMgq+F8hJAAPE333b12Xpv2m
4jm3TRSqrrejBbFjAqLlSs9MX/uYg74M8g0GI5iMNt902FQ9NPPdvCnEgQdwxZqx
b3oUXdDnKXE6Rb5PZafezlxGmH4L8VGwmTzSvToihvrRIRnR6MJOe1Y7vLKbdSdE
3Umnh0qcoFjHVkZ3EXR37JJAhXZsvwh2Wq8XqboKlEejqxrDNUwEN/XlRCv26xzz
Nyzb+6sE6FyfMRMAtZ7e1HloJGHOKTI9AJmkDEVPYefzcdIow2kck7/AJ24ZSkLD
6T4x3n8Q8lWOfLndBX4bva2k+x0XBP8mVnvmEedtUtwWLaUQiNB4PEEJ+yZPvR0D
rGeyEsTeW4Z5Tn2PAkyy6aFl/wgCWM5aVCRGHK4WLffTWIHiNlD6M0pW4vs9BTTi
wAig/7nI34uiQYizUb7RGFcAU0a105QwuZr7D9SAwd2enkcvf188+ut0R5Ww4/d9
0l9jDF/Yq6Hawc0U++yp9Ck22SWZaMo867nxKptW0P8wUl/MQ8VeM61CkREEkaUM
sqY4LJ0bd13Ee+sorNs2mUw8Dok8FXl3tqClq1edGsNgvakgsJQxXjmdJlU9xuVd
yBrTxNX+jGgy9DTViaR0OF6zMN6I/p/0JBvOU8M8AqS8g0/SFM7anyYeE53HdPvw
z70I8W1oA5NndqwhjbV+XUWvA1Mpskb5DMMintvd8ZghNyBp+02cG+ScgWJAcQWs
PUUn+wHbQc6D2U0F3p8CAmdtf7yGBjemwM3jtO7nwcsZOSG+MurOjtEJdQJySq7O
kt4wqxlZaMUow71tZ5H6IwQjUZXSCQYWmHylz/2AlzkOglePLMOs3y9uG5bw/2EF
f/mlP3fOk181bu0qbP2qRNEQMVUoMgbgGThyCROo8N85Cr16cN4VxA5MgEfWJQVX
MxLqPpLJmLhuiOghOsSA64XHDMWtYXwf3lb+lu7lrkp5mLPB7xt0zNppWAr9zYyO
zMu+GRJ5wHqIZAcaXgWlFFzX19YnwLj+W6rN2aHu5EYmxBM16mbLAT1MkbvHqYx+
a4AF3V49TUDxzzxBPBz6azUnwgD/7phi+0H4q/vLfFOjBZvXxWvkqWZeaXAKIVtD
xgNCn+QUP7tysRuFCzJgrvF+GXyG92CIMTbO88t7z5tZKqZQQc6fFPl8C+UTBhTi
QsmuE5yg9hZUI2dJa+bI28RBm5sCOQYOevsa+mItrdNG5zVp0fqu54kVHyKb5Exb
nr/fDb0WmmxH6VhCHkyvAhYESx8KtOTOPBWo3fgwzw4ORaCiNSTnUejIo0waYEqd
SEZ0ay+J9fYsJj5felEQA71jpskkCxbdDbx0Y+Nbwvd7QHmQd/Pr96RhsScsRL4N
OAyUF5RHdC2B1LvT4TXgzYaKMJYQG3pz15AH0dmjWosanf2M32LeuVqZO3dsTyFA
TOmBxB2CEQWjerxWtlAY5j+H7arbA0A/EV+tzZFqVFZ4Xxggi9lej5Z0CPKd3Zqf
mKyeAJ0Zo4KXLEFSlB8mo3pSpeZhJoc4nlkJE9CrJORusruDutSgEY692hPOO5VQ
JfeUrxnOj+ZOtKYPGarun1Gg5bMpEla6mWeEPho1tM4FIByTRQEDWxH1A+4e24Ic
3WFF2HBVeI7oU5V9ZJ74yesGA3fbnhmfbupCn1hnemmiJof7xbgefp1/bDnLLnUs
ZalYTa1tZ1We4g9+FEdTr9N9FglyMXRN1qQEtEQMDjpiQle6NGaVbvE/3JmfyLp7
9ilXt4tRiFyI5bQnT7HIppPm3v9lYrWrMTfeSgUyorB7KPWIj2hnkxhtcykx8Znf
LtWIy01z56K7nzZ2q295XINprCpdBWKGSa/NMamly1y4M1+1l6BnAMr+7El0Vz3N
XZJWHXNXNhxetOWKk5EeUUa1B0pCx6HFtRZ+FlDdwGEwYJk2UzWoJ0goVi+PDuYH
6tD/hFALjjwfnZP3Bdl+cCrSXsKcjl1sPv5YyWM40xIiizRS/rZd823au6ShGpqG
wS4MyqX4eksgFJEIckiNzUUBGFXFjbDY2Ga9aKsfaJ0N7w8SHd0wVyoPn2Mz/aPi
QxvtZVf8py95/EDd0grr1kquDErV3hxurZf5k3U5nJGE+f0IjAXvdLhN8ejvVKZT
zJcUQoIzB0SW3gegpqeQiJnWnv3a9Rg3smSfkh4vvJHc5s1acPpBZdzKyiWOxC0k
pYs2rUZ+gAVAwKL397K14FXNoSqU3jUzQhe4sPsZYBsQOKpxEvDtGirwS9iPktfo
uhU57oTlPwx8055tHPmj73l3pcBiNi9CYvv77mMH4K3ccsMc86hhjD3HRpO9b1Ok
hbkGkN21fHKNbtEGl5rdGnYMPLRF8yVSivkSWlicxPuBL8CAym4MC7ljlbZUHSEA
P1Vfq+1V62XKQWXj98/z90tZsEd1Z9kf00WzTRvUu1dVzHTgTMVkYdBiixj5whG3
rYxeNvdWlUDGlVy3gPpVS4xNtqgHBM3804dSY0HFZdSh1csmhvaVmhRzxjTeMJS3
ABUvwR8WHbK1LnYyQiEuYpJ/X2RHipylsiDAlBNmehWqlXDiRnK6BU9zn+aytBZw
KcpvkP0n7vEtG2oHCu4U88md0y4iQClLHjWQDOWSwZeiN05N9DwknO38v0PmyI/P
VzITUb6aIeSiI7nUz2stHhS/bkpT8blwM901NL57SxoHvqtf2H9bG2BItGNl9FRs
EjCM02PsfzmxGSupzVxR5OHieA1aJq8aevtrCHNV9OJllqHk0EW0FJW5v28Q6DLV
6nG5y4ZhahgTc+O1XC5WpsT4cR9TYxe35gpmjwsZRU6a+rH1JxChi4b3KYpJ5ITb
5gv9BDAnQvNQHYbEIrkGulasmRj+2YNrPELuEq6pLGQ+tsqpILSDQEQXQSs+A2Oc
VfFbwdevB6opJsqJa+ea7B6XlqZmUK3+eupVLLjBkiv0/ASwxJFibH7q6P6HtZze
laHT/OOFhMU1kWepPMvv+cN3ak5fuXBbH0+AeWNNsX6Qhst6PY3R+J7hd5N1jlOO
+qvv1LivloUIt18zWyQdomklKQd6myp+Kz12Jc/bru5HPuzWGBhLcH6xSQYUyLca
PHBCSyYvYWvgkk7SISVmsFt1j8qR2PD4ujWHweiCAdR48MIZTX1E4PeAFB1ycE20
mbZvLIkIxJXrwS8t/E3DQx1SxmBZZQXpC8dY8w5Y7NNTLIMM50itEiIR7P6EFRt0
vzYa/t2t67mhTYcyqf9KHRrpAEnVtbYyDKRLU7q7LCyp1uE7O5dnxQ/CdEOSGNry
E4pjoENr842Mdyg0FDU4Z39hPXYKkK8J5lxZGGJ8vSFZJsyws4/qgExYiOunOPAn
tmmePAR4qf2xTDDp2JghwkbEjSKTE8DaP4ewDWjRmBsBTM0Ba890R3XALled1n9d
Ze0NIECZW8Uf8y0ihYuFnkTTIuKTen7IRyrcknIw0DKvPtx5Oi/dLOtk9S6tycLs
773NoxIpdyXXU05AjZhnGln+amvMAfZFkmt51GOQRqNqRx2OZvT2GrnM7f+h9wOL
29Ktv+nb6Q05/KzfhOZhO/iOO+iWTrXmmn23eJ05SfK0TYycAvxO1fhEVxVIAlAX
rr0GFSdSOYmwkZ0UA1PXIXfkCg/5nBSucZccgsgoZSTuzfiejTSrU91D+d6rU4A3
sHl3jXFfPaDEyf9mlIGRDuzBL6YTGj3oz9lgVMHO3mTUy1ZTMaDbsl9iuqHkXnLN
kQpQHMLbw/S4r1x9VUG5XgleH4uL+2abfyG/8/UYTq16QgVEXq1IXD/jgxvWecYO
atKDQ9kKfZ713Iw9W24tGRFtX9B38PBVvQ0o+xSpn7WDP0fmnrc2YYCSHo3XRG/J
EUUeC+u9IrKiwCXNmIRzWbErUEctYYYdFGjH68/sC4HqVExFlL5279nX0kgrH7PU
2bjWcLUcgSGt+XM4DgmKItWS/eMJJl2hCP/BXrsr2iFIlBps+MiGy+eMxMnMzq3u
2cNPRW//cjurL0H6fgfWcSakqXAY0lsV1hnnSmIesL43L3T3o38lcM//lGnWgiTR
zbI0ilUhmOY9E6jG3ROectDSdzyLBOQAujCRUWddIfi+O6QlbASCErd3bvW67hVt
Lilq/kYPWEZO8aLqUcGlEdaru8/H76VhxVNYFrcHRBcNGKkOYxqyZYBkkbZjUq2h
7PLKLsHBwdZ0IM3Dgcoog8lqAzjsZqx7TZK+RGvENaU1sO7YJmKnJ3OmdlDLOSaM
Tnr32DlybbphTq2Rxdk1tnCu/DqkRF41p9jmpgWoxG3HSy1X7sINDgJx7x+fHtX8
JeRxa3qnBIqCB/4bI6bN+sIrVPxdzGXwuUDVOUCxcKxK5c1tJLpeqWEf8QwEdI5y
oPWgaK8bCi+0DGlL2o2fjNveqvJuX9Ay1pv4wKc0UkkSrj4zq3hSaq5VwOL4+eVc
xCZX4RMcINqot2pNtvhtPvdaXEz0EKPcGfAGaSEDrdIXvAmsYOGvVjpzZSqwMON3
ndPowr9mxjPel7DfyjqkU15u/X/EixweWni2SzTb4bjTIlBMA8fFLJ3hAt3pKGNJ
DrZeOGWb4TEneuere8+RTLZrsRBpuA+t1ExHUvpsQTx/odFCpOB8G/WzKKk3IsL6
6PApr9bA8JqeLRrQMhz6JxT055NbCI85kDpnBZxX8gl06LDOzXMKi1x2mmQ/yfns
C+RC2grV9wpPcmTF4R+uEK4aca6PIosiDU5FMebCZL3OSG/a4cmRBu/tnVOBD0YK
WeChWeTAINczD2BioMRwShx59d4WCiNeum728sZ5FCZfBZDrxjQmPpTzhDNxAirQ
ugwjXPfqftUIcCTwx6IkEdNJH0LyfLbtAv78fxtzH6Dnmci7hk9mrdog2WMeNT/a
CdXfFpswkxnzBctolCT4mOWREZVwChUYY/guvqyY+aTG0pqJWxEi/tJIvVez9bkh
noyTrH1csgfM6PHLrdr9OZL+Czbbz+GvFH1Tt7VjOiUyVkvoy2UYJviBpGyHyNKY
PN/ARaJLAjYI3zU7BI5RqJSL1k+R6e6ZRrnrdlQTs51BGSJS/mUtmm/aVE6vURKC
R1xZXgyOoAQ44AhYJKRCMtjs8g+TlNI8Lcan8RzEQXCL8/78qcH8xztMF6A5UPFK
2TcTgp1949lfxafMmjNC1RXRBYELQV7KbqJ1oBcZc7/GGXD1au/sCQvhvH3qq9cD
jCyIikmuob8zkKzjpggCsfUjmFtNzHewHrUxrZTIVWMjjz+SCL44MAf9wuKFYYL3
HRSI8u00l6DZYT52vwPrg/OreW99B0R0EYjssXKzqmSx2ZNVmo115K0HHFxm1+rs
1EdRq5oX8QD6vHlwGzHSIRZwo/P5a1/9SAOWCR/qqsBrVIGJUEpHtnXogluh/Ihh
LTmDZeBVxaN/4t1S/ym9xz6/+O2jeerOsY2fcZ0P9w08Z937PwUBUym5joV1jOJG
iQr6fhLKh8jlk4yBVC6ZMdYLcAQO5FW4EtggeiQhRuoso6U9Hltzr+rHyx18PmqJ
FeReBb1RlhR1rpjQX4TW8FUw+PTSZ38RfsBgLwnavuKz88nbJpKR6e8bkKwVbs6X
fWJ6+X08Id9Akd+LoOnCfSkyoi5Tmr5WSkNAPWZ56R1GgweLTlnWFVDaRizDB3JT
mrulJTf5SfTdRafQJz5Zwwwmcebb4r8uy8ZVjCupb8k+gWQxrYhu3lMGHCPXuv5a
TPTZqT1r+Wu32u0RpTwZyq6C/uwM4ocKMkKRVWqTW6AMwpfH/unzmfZ1OzUM8dKe
b13HkVrn03rA/D5XVyKlnyN0KLCbBlfiohBzflV0XHZBLBjAaletnDJarmuzZCL5
9STCFKXRBlnQV9ltRtIei15HP7UHO0oPbgCuOPuaUx+UPwNpNmCVa7DbHLyVptjD
bqgjYT24zblKLoreUVCX8vyICjOJTf1+3b6Z9yfRQ/IppOfN4MPHMR7fxu1TMcGQ
y0jIRSWPWiiX1e7HJQx7ooOzimnkcbKFwQz51HA0ghRRBa4eA5w5jU3keBGcrbU4
UhlVF5SM2+PUpX8/Q19h79zdPfdf/Rn1mX23GtoFyHiJix4+ahu6mmDP69S3MUNX
3t1Sq0woyU/dJEN5bBMQu9ys8oa+MX2W94oWeoSRGLOHIDP4v4T+bJs3P7Oy7clm
2UMsq7FG1IwElBHtSa8wKxyDmxsjmAouSvqm32Ew0Z1ghFoRHRZiRH6M7Ajvramp
ptCOFP87uCSUxmp1GjIWUTRPtvQupS7EKU0tkfXtflCuSyfBcljusNlcekXsiJfs
seJqfINYutJOlmoXtHjejZo5gJg6dDzb7pMLHzm5vb9zXQuVYFYpB9srB4pIXC0s
4Y2BKtp0eF3GuytMfWrS65mTwyD8q5hjpf44brloN1FYMRBV1LmyR1w7VA9OuDBb
VPeRDMeS50eeArwcIY4fcS5qkZZnzhWTLiSKoeT4AXrAOkwZe+RrW+20JS4bhkQU
zvbTX1telO+rTxxskMz+WS4FNU8PdT86/3rwLjWVvPd3DEzCU4W4Lqv90cTgjpzI
UDSzOO3DIV1Lx81msMKF9+C9l9XbL3zv58u7Ps+cZG/cShGajRdZmwwgxHvDAVFQ
95viWPFNuOhzgC3VbsWWgt6Z2klYqz11cdTLi1FYXf89Qjya4OGHGWUq3EZavWjp
Zl6w8fVFx8j4+WSw+1AV2gcBG1X5REzjMrUDcT8xRITbgVnuv5/aYElGlVT7qQMH
Bef5PxIB3qDMbgjkYIEG+o6APgGaQOVjpXUYCaEtNYLDZ95L79eihvFcSdGFmS84
OfJ9VyMMWH7IR290jWGgq9ZaEUTaulpGH7KIjrd8faEx48BPQzRnYG12MDp9S3je
gkxV6Gh1f6pHye2qMT5/9IiMzkfWNHrL7lRbloGcplfFaZcs0Ytm/5SPNn89NZWt
T6UFG8rXMBYYVMVc0Ci2HLnW9nMEytWamsC1RPZ4vf9/Y7zLgYgQmt6928EB81Dd
t6q12tnWDQt1i22wAVrKxJPaNIkLlU+PprlSm2WAF0vQEOjHabSbc8zCZ6DzOTdR
Mqi9R9zcPBSlqfmIGX1c2F5Rc0Z+otPyjYXBhG4v51GsOHhUf/OzTDNXk6NtQd+Q
B4VIVvyqfaAn0Ou9/rdwAWnx4z74qmrLzJ/EReGBiX0JzIz4CRWuiBpC0i8SqDb5
NPCqeLlAa1JP14ce5H4oDs4iEgWhGkHKcTza+VwsZQ+tqEAqxkKVL3fWKXv6IJOp
J6wD9vhLwkTmEApXbTbzmLF2UmYYQNNMCjwtZRbwK+jeFsu7sOLwwt0YzJO9fz5f
xo9mwuxSpyo9Dv3t9MqoC+g0iU3HIEUzUvq1k8VfUD5zrLCqaRjjozgH9Kg8YPIS
Xz8hqQ5GydNTBlZp2k1/W+1lNlc0/phghe5zTyhtntpxP2yDo7sd91AetI5k7Xe2
oZChbTdgXyt0DSGoTb4qweWvaCIMzbeYka0A25awo1mJZh7DWcB/+76G592N4910
SpID1wXNUkw5DZy17zwZmi54AcTfAhh0fifViW7cpaSy1MzLgzFO0Xqh7+0taIkX
LghlNTkHtVHA7kKnObPnH6lRTyzN4ofzgEyrrOHC3gRmXIsNocnmUG/TLF61biNw
hhqPuGqkqxYlZAoqPS9zhu6KSlcRnYsTCmZHdnFTFWEgpCoUybzSa6Ex4JSMeGwW
B1Qj0bvSxxcd0kLjQRHjFrghTMi6Hrz8NAEetCdwMaocBxiqWHm5PcEeE4wAwZuK
/VGKKGO9kV2V+FnWfRvAhEcpYhwRxwmFURMAvIZlkYO82JHC1tBV4prjkSxk33ga
qBepK8oczVVCyNCNQ9sqeZlI+VDAJLiH0yhiXNsjkdErM6oy4OXJU4bw4QdYhaqn
9ErRosm/0R561UkWSaFYhyg2XfK2+N4PWOxLwJgxKynEd2aVO64ZEFfyBB/owJEB
vbccXUVW/qQfIoxRZoxG+m9jSg0rlZ32HIeLkyzPeGlzLw0Prf8lyAkrSBI/Pt7E
U/VCOIVlhZSbIBW5kYGFEJLiR7L1OjnbeL/lPLBSdrNi0rnB7w3Rtb0GezvOwP5c
VqVOu7o5zp6ggACHse964NInv78QIGUNN0kphVBkGCfivIq9Zl69eUqXmjtbOcCl
KFf7GtQ5rb/+TIQumHFOd5c/I6eGTaYiDQvdbrYonR3gpFrTHZiiPDC5VZUx73sd
SG7j9BC7a0QqzCQCQKmbZB3o4FiBRBDO1iSTzHsjlfloYF8mcd3WOSB8jWCWIlsJ
RehO6fw5dhpnlvWRz/pzOfGMx5SAiAuP8R6kOqHSZsE/dSMFfhPkwxaQ0i2rJGd5
wLyDqauQLh7lOtQBHYaSnZ34e4DeoqnazeCHNH2GC6dr7mHqaEfvRMMLgJz+stD5
phN2nTk4b3a696gVsqwScW2fVVRJCE/KHhG+gSshYsFtJcqpBPbz9WsPlnspE2r7
bjTTsuroLqMfa0Ofpi+p5vKmF7z3K7Whe8CSAXXnNtGB76mDe3mlOA6Y1Lqh6jgd
o9X/Cru9kvNg5GllKHDgwCQVCwYYQnM6SBC1WgWu7tG0eC41h7ImLep3pa1IrTNH
Ie/XsyNh9iyqslh9o3qgB8IV/xw+lzjg57eaQR5Nt3vzg26/bLv91ZUuH2fDmR26
dadB3C9z6O+HCR3MvVnSfCEIaFu6uxL0UPJnk4PenTtaTiuboDCF1tmrOX+INj75
jgdJzA+w94KmVEoXSXCdY5Y8OhIDd1jCM7fRyEJ7ij2rrhXDeYwBUKDadR+v6S9i
jwre4KNu3Fkk6vKmTdz81URysn3AuPM9uG9WYTFoOG50Z+sok7WQsUA6BkKH1xSk
8CMrjMmUT/75E8I5M9xxOAvP+RPdbNpkSuP3gQ3DnpSQ7qF7eXwVN/bkeWu7ibOG
WpGyI0hKFF0TXGb5f7bmjK9bNAMqLJlb6XUU8mHVX82BRF4o/UQE+z6/sZQIfScB
caAX+tl5jAkAsYrSbgO58tcWXHwKWs09cn8DHRA1HF9hW0tkdmj4hDgIn/RKCmeB
PgYT0UfSB3V58d0ASy/sGpPkTNKDezE02a1Wo7hMfFR7AlAs78Lx1VoLP3vX+qiq
s3hcUBzwP2HJGGcgwD1ct4AgA3kjPcD7EQJqtSzmBKQfkbMXXkVm7AisGV1wQS3y
TLen0CXFnQAqdQz11gaNdxT3Ml7ol83TPfu68PGwe1wWsggKfSXr/Z3vNUZShDzB
AvouZVfZgMPo9fHPIMfgMhFh0yCUkyortghPE8lFuHog2B1++ZZm+emyocYr46XB
I71z1KBzRh6hWj1/2iog43dSF0rL/4xkcRg0NbHLor7RO8RCAt283x6p2BopI4lu
OKkwr61jpcT+4I+RfOdZGOunE1Tgh96SjK0H8yFEPlCY3DPtTwtFfMvOtIXUHYqo
pe10KvOuzPQVIohflu/SU25J8bX33eOVGyrVg9gkR+1qffAj8INcckc1zcoPqWIx
Ix62dcB6F03HLYmYg8Cglz4yi+Ih3yiytzumJz0NRb6z1h9UQdP2mrAYEn+LztKD
J0jE5Ip+BMOq0cr/tXyAiZXWTJlrK8R6wtwUL9mL754KlDHV91JN1Tb8L0sEaDlH
CjGU86aCsCWBl2cD643TyZvVMt2u7JJr26TPyXd5Di+dMnR9TRhp2VNsXSGGxGtC
WALS1noWe+J9AVi9aMzbDHb0G3XQtpFZ2lhWUuWsuTJ406XhodaieSqT99uuQdtu
m+Fw/uY4OtjfNj4UHvM0ZQPkvrNf4kqFI4zR7K1FETSkhGycEBdGb3qeqbgiTOsF
GGPiS6USzzTBoYfAr92Rho2IVJSCswIahsvLaNBfZHcoF0NuAWQFhvTOx8qd5ynE
LHFtcLg1NRJ5nxJnSoEqSxWVwzUumgsvFXUCFrGBHtaPm6fe9CkvdOzsBcHxLkV+
2PDwUvbKZL2+aegNpKA8PMJiDAfWO09gwMVjutbVx5LwpNofjhDDt7/IeEoK6TqW
WvZjJc7sd/34jX8dOUGhAKFGTN/n9EtAq2g4SFS5qWbkyhzDISNgMzrejjw/8OAG
H1GYY4cTIOmcNAwU7Qb6+gMuT27db25reA8yybSUjdqvUZHUeY2AqFs+95u4OEp/
Lfz3+FRqVqAVvuOsAhCSVdGzYkJpk/X6mHYJFxXKHEeHnq7on84Kvwaq2Oh4+u+/
opiq449uzdBM35AGasqwWxMTNHuW+aBje9x35DDDTLe7DwMxuV9JWU56VI3vYNN0
jXJ6Ujfxftx1v5sfiAGBsrjhl199O61x984o19Xe2NrLJZZ/mg0RkDHqZZU+cV4U
gbFeFqaTi7eqnkVIP5Acz9b1Qi6Ru179OrxyxUyarD8P0VreeHEasW54f9mZPf8m
X0lP2TaTsbT+hryagtP+/vVCDA5HtxzaPNaCgA0SRyeey9skMFgiETYNAbFoJTDJ
j1mnTf1U0VfPj3s2PrZzPS+o59PE9yiORRzao6AfpsjNHcPPSIQs8c1sZFU1TOcP
t7kBc6dy2+bMyiy12tGZcmRlUsSa7xjVsXqFRqAWvAMZplmbmZ7qANSNPtRqsW1R
ETp8Y9niRkRZDiZ5pHAEnvw+CQCeRXADmTdJxCx1gkht50dsIQ1VyG0nSnUeFx81
Za23TZSDC6VvwTjEmQtTBE8DvBY1NuWZlKG90ri5w8jrCRVqE/Qwq/4yJh853lu3
2H3kAikY/rGucs1M1Jeki4k62R9h4wJw4XEpmmNGO1syMbnzZsvgaAEyoQHDmN9k
BoFw8bdNDi7Lg40ZsDmhuXJ8TIh0nQEOTHB0ui+gKTPGAmtSxYMtfyvsaBfzuF65
LjS6/koT2eCwn/pX0SD82cXxfWaCWizUeYScFOlFcXjCRrGCKHD6dUJrGcqqcRBw
HQ5Q5EWDVXgoPjpEwm1GRRkqnMIOzA9CVoVtbzXivDUmIdEWRGzhklZhkjCmQ2zr
7nZ/szmREqVONa93WJ8/vYO8OmUJO9AKzyPUWKnEThrZI9C5Ft33QGfiwiZVHsAV
+/91SH1DHpf4r9nzlG14wfWxWNjKPrE+W7hXWHeRMvEeLh/4xveigvHj72AjG82h
7HZkPkxecRn6FCDAQWTrUIdiFlm2sd1REmHnPRxoFVFMiib4d/r26ey8md+jUSBe
95La7PlddsNthQ2+8Fn4GwRAHVbb5orfEEtCpJ8ozz1P9GePJRmwozoYOyr1+RLj
xRUPVUPl7sVp+r8dM9581nGaTxTcde/LEtn7vNwXkN2Br9clFBe2goTxPu0r9liC
L1wYV8y7NoN6pCA3WNiUzfT12EiDHLU+CbBN3DrP2dWYk4l4rWYiWQPmXlUTw0yl
e9l2b1fS2t8iU/9C8qb3H+PByiUFcuGK0ypEy/7nOaToI3Unio/EbAG7j8+5KKV1
Q5vDjQqcDsquYt+oRZAAu1r1MACx/Q7iAimj2zQ7EDBXefOQy1HJI+bWWNTDbmfy
J3+zMoVRspRiU+6vgcdsmo89Pf5TRJPMBD4Cr1pMllZzHr18wM3ZVTwVd3k7JMgq
/27iYH50WeXCHpeYtLWFeDmQJ/Wd2/tKbD6FauuIRCq4Ptr7dCdiNhl3ENyUT9Hq
5hP9+fwMwkF6A4f1FofCLGCGrRN6kfi5tXjhiotJ8ETm8inO+I95RQGGs4QN557r
USb7TCh2GoGnM7M7rwXW3YmOa+P9hWgm780ZOlhYHxYRPtpD5j+NYHAflfGCHWYs
57veWyw/Lm6DQEmYPowLvJtfAMtmiS08/I7Ekm/KFVolTd2vEitercg5cCtfz/Fx
jT6Hr6goOpn7PhxpDvfAfl3/essSxV3SKOFS7f6ne1BXPKmMpAxDuOVLY6GHn4GT
gvcNREbpPotLudWDGJ8ER/YTCeZZtsDs+GZnq3z2rG1WvCAzT83T92ruFd9ZTzNM
mBXhy8ubs9UKStqYZHW/L1Ea8Y6xMfxJ3Z74I1hTe0NVtXQrD71qU2Y0nDkV0LJI
LF0MfmjSVhSbbmtGPtg+RTbQzWIbJvUyHrf26sW8PMhpHuvRy88CbkPRdh10Eagj
bMsUZbLjYtAs+32S1zX4SG7sxO1BCxX34FDrmY+9kodjO7TYKQsy0L+NyJJqhueO
jjvReLZwjpH07gqxZ7uDzXJlGSUODAElfN5Vq+W3ur2tf+m/J9iVriuC2kbC6j1T
ODJsE0ArSXSBPsenEzdhKeIChBW2XEIbj+p3w3l2XDy2nxVaqadAf21vdml75PVb
/m0xTYjl9sTTGW4SdSgy76r3+cteGJsdwvg1xxEyKarGzSAZf4zXPVHqqir1v56O
us7ht7fsnd7rtl5qR3Vyr866chDc6GlYQYZBbgVJXe+qA7RlJvI9lNF79NkgMXub
un7kr1lAuuDM/ZshX11RXm6bJsh8llZaD6bBUNUYc8r0BnQ5dh8cnwrv1/ONtkem
DZckmu3UARcioOwthj1TyhFVovu/Lh+GufN9zRkMYQKFBgLI4BCXCFkgp7OYOrbE
0mQ2LB/wxQZRP8EcOi7Nc7vDm/BbJW9MXl0SL3bvQLUqFJNGPuTT67hy8emQQRZ1
Usm4O4dTXhmNckvllOm0iRpkuUJBPxiwu3l3z2JPTLLeyv5qwY3GkwZyzmONZUZ2
5I9t44PmljRNM1jhaa0/hLoWmMNlJvEj2EXrUEWRR7S2fx37Gc3I4eXIitPKdjpr
HhOl0z4fgeV5hsINrgLRbhQ1dUh9JSYtHmw+tVmmdNBuK/OEN9nWiSmJjOdkwsJL
d2gyOsySmmJlJ1pgJiepbXRJdIYU0UBoAuHPaNqcTL3g12ae6L0KRPOwkB41/xv6
nIabZ0ijl1Pza9kCh7QPcSOb0npbuZ3AyAf+mVRo/sTeiguxZHtVmnmNyZemHgMY
O9MET1Wl4ClHlVWdYVGtvrcW/+RNyYF95ysXqjSHzSDJLHkxul1G9Yy/6WhxBEsw
zKIm/P3J42l/vnM4ln1Z97uQO18ZTvxIDqDZ6WtjO1SddDPqlygzkvcZ7xJs+uTa
5f5tDDOAyFBiCzeU3YcXzuU/r/LFRkx1+UPLHz9dGr83QyP28/qW8zzGhKGUd16R
9zLbPtrH1H1pNVoqIfcQthC5z6RLAFaNVu9RGVGuMTkfwaWLtIzKoAS4gGWnJhdx
sX81Fa5fisCL3XIKakP1JIvj0ov+VISlo36WFGh7Yr++65OgOFGXbsfUst+eycXx
uguad679wO5rCWdKV86hS6dvdvsr5Yp/57nph7SL4mthUTyKTUjMQRSPnvQgve6H
hgvuU7RWr8tnEGz79VMtBO8K9tl+Ogq+YQbORjPf+uCn8Gi8dWKAdkh6cu6mUzix
wO9pHzt1fRLEZ3cjpw6hGNT60QDFFhJDHZKhjS1+E5JntbVDmogrdF1nKnkLd06p
nxdXw4rSs3gtRgT5qTKJXEe+EImEO48mD5mj1f5rOxFqilJVwtQbPNNSAw09hS6C
ulaTTjNEJW3drWex6DaEhLodctrn2Tl1Ja8Ld5vKxh25ushElWtsYnigVlMPwOqW
iAdfX7Z5wMyF///lQzTQ5dcVo08YbGAJEB7opASJICgzRzY+feWnEZbTHECoCrth
wXlX0Q7ly2hPzsE0OwTcC1dn1cy84ka92kOmv6lHQ7nSc80kELlS3taBvdKywX/D
ynyyWElv0V3LY/O+2F0GRldm9vAsPACEpS7o24+KH+qb4hyCSe6SycOOxpnxLaYw
CcxuV9tvmvAHeqN16YsX+AzzLe3GibklLzFEYyF0tCodb97uqFPBC81zd6Uzj+pp
cfjk+EHz/N3bN/oHq0iiUnUIsCXJdcSqlAHdMKt921P/JReGwz3wcxnpIvIkES4u
KFlJ0nXeLu3afWL+exrponRGTiJbf1oDXfKOfKwWJyKjb/YXoV3VnTruzeKeMC2z
kjU0GMrr1PKQsid8mFkkOC6sRuQ8i2dX56z0NPyL73Rp7TSg+DjaXxb+mT3MlosN
aijja3B6nQngVHqwhjikRdkSuHTGbsy3TH3qQ3yYFjdjM2jii5tU/qG/NaAbteJj
iR82owC0r2nF/JbTynnzfxQZE+3QKg6gXNj2WL9L0vxeLIm0SEeTj85JXcjZnha3
LEiW41+icJackCxZRLlKgMDklgWQVLgBRl6I4Cn8f/6pjGLCmlvUtpwVCwHyHICi
T1+D6ZLM0/R8VFXkTL6gVMie+XRzfjT0pNTxxfzah6kDtqLVOof7FGh6nNMqOBHo
jM/kedOz8iES83Awa+UEfzYVxgQLdD3wlfMaX8sqf55OCloGiGO3/3FmLnz9GSw6
UoqY5sDr1TRiDfo+Q9W+KRBYW6NX4DmqVVF0LFpuhxagj6diZIn54md3hxgmv7Gw
F1Low0pA6SB9HIkjbL/LvzQIUoh492N7uPoZFlB1YMXJUDQCO9MUHBH09AJxI7Ed
jMhRK6pN76iX0hJD4t7gtg1kNoBl/bt8X+jR1wVx5AcTcgnCxCqdTWGoAOj8ZHJ1
ruhyzvHSxqUh4q57Ez9aFKEpnd0IayYMtSaHpRuKDU/VzHcYeyKmeVHvgVBJQ5fc
/yOQrOmuzxaSTTwPVHbwjGB2x/IYmYhCQTNY6EY71UgaotDSlZwgMPn+niGP9jNU
sZkW+Nc3iwodaYgM2VY1jyQh9Kiksfx/0WyjwvItMhxRECBcJWN7l92CYxOzuLBs
UTbKXSGk1cxk/2Vdv4Q9YjsyRhss9e5T4XdqpfLQGQFO1IaburbaWkVG2WZeKmeZ
5Y6atfi8iBSBksATDO8mmTdErQXZ7BhTjfSE8+1RweyZhseXZkH/WKGm8G+DPIF5
CNeVdqi7JNMpzw6HIpBXPky5EPVlNMKdr79i/b2aXd8BVe2RsVSNfYJ+l7nfPcMd
1bf9E8VDfsIo1hzeouP8djXcUc+dknygqF7l8+ET0X+1tqUAn5p7+HzTueGx/wP8
TdGOBNJxH46jWZlH6yOOMKeBXPeFSteh9m7Yf2J2KniVD+W5+5abnkdBvw0sOZHC
kuRYLTlplR51YyL/KK+lA1zO1AkpPeuLL1y5EjFLlkGgSEQSQgyUf0lyy74w0aXI
39nGvb9GuyXSq0VDIfekvb1H92O1Cke617ax9i9UGQdOhqF0aHeqsFcY2bzpCEzn
TAW3MDUx91XnYLMXdrvEEWaDA/g6nMCGOKaDu+dLbXv/LXA0Qprx2iZNQ58prfSP
AI+ps70ckkZ+pJ1IJXTa3mik+N98wRx9i/ZjYrOF+pRmW7PSJTvfLeeNSNocWdb7
gRuphFu+iOlqpk70BnTqUVnMteWBpAFKj4ifmfLGfknWRqwjh3FWQ+pfHGpHoVmX
5uYNetXmPquUECpDWtM+N5rwJTdgpUsVvYR9Odzk4StzbOAXODjKTOghad+frGqE
MV5wvL2TU7Aa0VilnsP7gnVqYEqd8gpzUW+pwdKULtMuoo4NiXPLrIje1suDhHVl
aow+ISkSRABdbyPfTVSnOnz+5997nTE5e1aSeLzMzw05iuct2sBmAOa6gfCvcu0+
N3KD+zZlJORtTQL637sp+fODyH16+ymaCjqqcDArNspr8PqVKk5lNODV80XfQInF
rpANJT49t9br/CudVqJPIFqFH1RXSCdhddYl4t16d1V176n10XziZTg15mdpahQL
/wXAOIrM5fH5sk5PJtN3PRfjeHTDXu7L0XU0Ho2WXxuXt847KlOyQXyEd2vABseQ
Jvaisa0PdpKSYM4GHIFciuqAKUHry+4gCEurAFpCQp6JgLQAg/M1ol+gtUYDJQV2
YJ+4/60yQkCOgz79hflwmRemHbotzEpPnQZG/8wF3lC1EnjQft9Nj/voxZCyNfqW
HPU80aUVHHwzHQuTGwmwMFQa7k8aHvzgXRwlADEWDm9ItTHL4oxXJhsk7ZcDv9sL
1SIcHW41JXTh93nhoUqc4cE/YLtCRLD9Kq7POdkVGI5ABpK8fOw9K+M7kQXa9p47
UzkU8Angyxr6Fo0wxeH9AkM6dDa5GkjZK9ECMjSnGCjzjsBsMEsiCnVn7IRsdtJV
zAvbLyNuzwz7uejkhXZ7SWMb3sisGeywYJbYHZBU0MAdcFAdV2inffNFAVMtOKtY
w5ygsrjGW6wwWsKR3XVilPw09ndmijN/vxVIvYsmtVV//ZL38fq1B0aH4sZMTHKj
b2PGpD/A4PxOGIGH4xKlw7RL2Yb/yyltZAkWL6WEC1OfCuaWK64d+AcxUtKnGh08
JmizN8hb/7HSKPkGmGnzAAjZcDh0m1tgNwXouA82tUrRo/d8kEnNKwz4epLnIO2V
VFs2n+3QHrxUpJJoVI8dNP2wpXhLWe9pKh8OPA4kTVIZBl7bOWOtKYJ9sr+efdRh
QEq4GKXcW4hTDSdJQ6O387Hp9zdcm55B1/172a388MgoiVxFwFRHjF/8pD2nwvRQ
cGCuJhCPI28lfv06POAiLuRWBts8KfIXZmkQGHVZP7LbF8FDlRtkb3k7rO1CsJoR
jUei7nUaTJdzQmbmBxNRRKax7PIB/2stNy295ZgslR7tnbJWSgecsoRqlrZK7vC2
b+s9gfbIWsANBG5dIzUDxQTdnaSB/W8xy5nxjP9YgEXzqspD9O0rEmFq3Ib0Idwh
HJ/dkPm58qYhKoeXqWEL3sNeztdhVH02NwubDQFDg+BdMFFWGz/GsrF0rKDkKkab
KuAAxe5hzA4dMqhU3RzW1kIRhZwd8uPBlICltIYgMCcp7vkEocPZgOHkzhzvpIXY
eWTnQTceznrBq+mi6KiTA5qYzuOMoCRXYe+7SdNin7bgpOI3huHGn2z/APmP3S1m
GeR+XF5Dg72YDaWPleXQYLqmre18SiHNFP6rufYhR9Ayv2eQSQIh9RtWvi4wAK0C
4Delkh7gSDtgZMpSnwqmCbR9s2PyjWrVaWdPZl2TEEU6zTQojFbpiXVZ44tXqKgk
HMfhNOZSWTjh0330R2FjA66Ak47slF/minn7BMkOGinCju15xdtOOfBgX5ZQYRgN
DIEeOXgBBxxgKcmJ/RaGBLqvt9jYM9auHw2KQa+QuNIpIiKFcaTPfyLt4qY4ei/q
YUJqoA1SAvQiOLnmgSo3tMwWedr/O+pVV/EGrRU/Ztnjc77q3rSV0cMLzAni0Byc
CvT3sipY5fcKoWLP9gV2ICTN71Xtn3vdiZnM6l3raTkWtc2JS7z6HcxVgg2U5xJV
vv6Rf28uD2aLh5yD6VcNSIUbBu46tCqQER8f6nuiigYj9mea97vTcW+JnjOKSyJG
dIsoBqhHCFIoSCo0wOTy1f3gj3ZF43E3GQmEv2/3o4aASAVG/Z2VOLSRi083Ay0i
mOBARqxjAP0p8ZcpZLz2F2vGTPkjbxkBc3ZFDxDskL/sdfYErF0eNFi8DkEvSEum
mjT32VjZP+2sWutmAWO6LsYKNO9LcHd+YOxerGDU5m19wubbjHAL01LoWU9aLX/o
KKE24P/8HSI9A+LMViWsUfh4yswaV/LMiaoSrU2qiuO42Ew7AR1b60TkfDlCmO1R
MZN6RfN0ep1ne2I3KzwYD3fzRiYr8pvQ3ORJ6vfjR8+BrSX7oUsL1khjBfP7+Az5
e8GfcoT5BMPv6Dzdlf3GxggfPqCsCuuceECZiot2+m/oZo1i6ac5u2Drieyqc6WO
05jCVVoHXk/nW8VYAFGuEXa5pFI+zlocZLYjVfaqes+vwDHnSWVnhAMn4KVp1VNo
4ReYIhAdGNngO5ZH0wtbeTpC7hLWiFDiHEubBA1QeP/tZ4xvKXtX/Z5PuaDjOWv+
7X0Xa14ADq1qMcxctA5v2gCvJliFtoR6+kErNeYoy06qKzM65/Gft/tU96Rs5JAZ
8xBZ82aI/1nW/Q/sPfZwerIf+pND15MB5kA9aQ3ty+S5wILNJ3vDIi+0uvA9nl+l
YFdiZz4Y3K7Od3/NclD7f9pmDOL14nPmFrRJAVKUfacHcqq+zpexcMNyAtuBqf3U
toLAtxsBPLdOtNOelMnpoRgtHL68vyoIaVHDk/ZcbsCHIsMHoXVkNT8Gu3N2FOGy
yIgc2R2s2YZxEpYIr7h+s/dCohATGV7YEbtPTBesPgzAnlpo5LgNh0bGeW/00MLI
g46A/PqnnA+k99tCQk89Wn+18cLPyASsV12h721FlZInq+TSnFuHa0k82E/N8m94
eS3rMPZ4tTCgWI6X56hZFelJlbSu+2kbmbM9lmtmwbJIVKAmdT8xp9xeEV69Fj3K
6Q3rQmKD2ZQt+M3A08YsTWqCfDY6IfoqSS9YPoDU+KBn+GIl0l83mBw1b5nNjPQu
yh23YQUAhWzelt74bc8OLbXS3gGWGu95a1FfzGAviBWsSkdDFVE9udk7KL/Rw0rZ
ko+JODNnb+56/DDVOpICYm+1l4PGRI3O1B86oFBgR1wznqOdo1ot03AT8VdOdgna
jQG+EGdHnBaLibZs/yoQylQEapJZnmehLPRXKWG0v3/1YcWTUorG72/UH8Q/CI5N
++tcyVq3AJ38222873Kb3rl5zaEtk68vpc1jZllFuTFX6YiLSYsXZmOT5uiaCYVM
V9Zbi486cqog05+CVj3dXT3COS/kjD+T0MIsPmZIGOXrsueD5Sd1tSjI0/wRYGKg
4nd24kLXeyC/gr8N3wQMBTrpwmLLtPU1Ac7ymDlbIed70qReOW/XG1isNVB7gzf5
Pz+fx0yToUIATuLZtZ4LWXJVFJCK0ghNryKJ5X67Ey9mZmMYxufiJm23JFJzdoyd
fwzY6BSavUgYRxHMFSpvjbSePr1eTBFAGYXrA/aHhWCStDNim4ndFs13P/UJggoE
uaYZSchIDlvgkh44gijY1zBHJoC4VcyXBMsjcScwMX9nvczQuH6DizWRkRfkluts
eWA+DwVxAIl+zdofEO3J7mAnIy/kqFwAbPadCjGm5yAJsMuIclTfLHIQYKv05b0a
ptJ/ka/GrZUqUjiESyZ92urvKeN0tE1CmCKkEyllK2/ilLAU597lTza7AUv75uBD
LdSRLnC8nLD9//DacXKQx9aQTfguQmEFSUF70o9YT9YShae6fdXZk7hSm+zI7fi2
37vDYMl04i4OQIWCLYGf4r4GTCd3PQY45NI+vgBO/HLzPPFNzrX5yBFHHlMDBrKu
TfAB0WjDZLVmjLys62m2E1iRdZb3/BzE9EPOpWx881aWRsyiDZ3qrO81CcU2gcqE
lyv/Yy/n3jH4SZ2rocXlu0CXFNTMlLSo5Vpjw/o0yYGaJRQ0kvxK7sLA9003kv0n
HnZ2+JEifD9OEKCqRVeGbvgqcL3M5AxE+mcZcbBIPwARgvUNQkQ7vGByTmizYvMJ
sxBHVYK2Lf9t2lLvTbkUtUKbHofrWCnNUVAsgm1vSnOO95N23GOsy+ipkcr9gCzD
QufutkjHlwuOuC7T/AUVy8KUpf09j8BBVeVNE/E23R0gkESJYcW/6Od/0BPfdBmX
CGv/D7xcO0tiXpf6fXD2ebpn4PbvpoSWij+BMA5KFZzwF3JOc6E4HgjTBzcEjmzi
JIehtKyp2cgx/FTX7O04124a0IjGYbQZ7TCmJUxN9TL5wxitXNZi5fxCIdoCupWG
tUd6Bm58Ivua+DTpTdlhCz/ziPMI0WlpRuCu/qVSWSHsvViC+XeQ2G7YDRCzSiGi
9/8MfkBHxS2Gbbxj+M5CAOuLLYiLZJbikKjrm2vsmtpCs1mSDVgY1ZTkdHwpAanC
LwAuuQ7BlBWcTXiWk72tCmMJUenepe33bougVjgH8ukJvi6klHrcQhk+fZWMACYp
Z+QAkhEWYdLAwj4xDGU48qR34NoJuDm818lcUkewGiWW8O3srAMjVt6fBBmAimRL
27rtUmFwZ28DSZwJzXLlAFxcMuIkJr1oZ2YjxY+g0gsxzYYAjrJGqNYLDRHILw6T
rXd38fwY1nK2KKMY7DkLakPnoFzdlrz8qRg9b5A/TKi3aaBRyx6wEnrFkVfArRzx
GQ97UzNFRjI7gBdh8Xl8K8tC71Qh2VZw5gb4rLZElGbJepJoNOU7suQwNgzwxZAR
pTsfjNHkeHVfabZZZDO/as3DDZJOMQSUMZJLpxwzKPcvVQqksLGk+pVJcwKF3/7D
xE4CViF/Z0HT+WjcgxoGU6vr1MJyAWFue91rlAz4Cx+fWa0PQ4fvUSatfngAbSJp
+WNcoL3/loI/rVR7pIDlZ3Uqe73WSShJxFFcjqPpYFzWbW6DWqARAJLdCmlNgUNG
phGUN3V8SMW650TgPFZfBMDbq01Qipf6zciAxuC72JijI02HVco+k1kG4ny2z7/k
K6WfvYhw+vBqcN2hRmk48xmc3j3au1pYRy1XChL9GjMdbPp+Dqr0nbc9Lp1ftIgp
elJ29BIL7UUjx5nrPvC3V4p7Xp4iOzYdqSYVv8dX1cEgFTRSxBy2zb/mW2QHgISe
RfdZqgJ/KappdkOwCvKh4Ba8vbMiizqvgWfdXH5Nnnjg94w9peZ20QGqxNfdNDxJ
oLKAy/sS0Xti6Kq4joqEF/ci6Ft2TPmLQ8MQnzU48Es2IAOekyaO5SigKDXHFjru
xA1rumRLKofLvTTJbDvYFMSZyH4aEBfRU3dHKTna7FOqP5q4YrCgwbLC++T/Y/KW
qevmNGNg7pQLLowwNxbu9lsaJdBDdC4dLc7T/jXieBAOEMUDdD81ju2doZBepxih
d2fXSfAVCKWYILVnkwcR9RT47m7Sivs5uW6NPtXSW1gCYd9ejhJsQOhpdXpKBlaL
4Wzc+wwebBz10VG1gjmEHiQHIW9H8Yj2eJy8+DfbGQJwnZWDmD9IPq9MD2zfaGsZ
tzuvCfTLU6poU0EJmyi/laqrvuWsjr4VD8pc74Zg8TAEVrB0fuHxKp3dA43rHDpu
vpG4G1D0L/4v6JOPNxzIxiWciliz4qhmkn/FGe9Yp7wqLwzr70HtgpVrN6dojejT
LuQXirWai43KcibzBLrNEhatvk4l8/q2e0o41Xnvbhbz5cebGsPQ2KQtUQNJTjM8
W6KhNG2qcUpBz8IV3TY/LDs8JaFtpBEJwlFAB7vR1viyqtu+R/DufbnllGfPtW8Y
6iCSJ8IZgY6uC8l4nQJGTtyFVmCWNcOs3fwBxcTis/z/GHsN0Fatj27NS0matU3d
GMvWRzEEDvVKW2Ds0iCwJ1fCx9igL+Cbn0owZzqJR9+DFpb7bsiMhMyclLJJzt/b
MrCtUpvdZF8bRcJYP3YNUYSMJm7P7VTEaOdzL0A7Q0kLc/VgHUPtQvE2k47/o3gV
2D/dD5yr5jkcyieRm5RGK0HIzJzdPrB93tcN0BSEgiL7Bs1ZxvYyTCo6hKyFgGoD
ELOfp+fOdTEF+3su5hYlL/I9H4pGUhpd6vs8vTsJJSXgECkThpGzbcs72je2Frf2
MeeWG6MdOxFX0dyvQnkNSWqZDgioy/iQ55E8MrwQnqAG1YRz2goc/Algv3chlf4E
+p0Lg4kYeXY5qj3Tbm7XDzwnAOW9sTzQj8VBUOIC/GI0Ry/y3Bn8dxMWFEouryIg
2oFonWgduZRAVaNa6//HMUHUn2bKvEfeN0HNKJtqluROoCc4aURmOgkVCMrUSzd+
lgv50Skv7LQ95IZzevc+2NRkwc5i6S1qjT3/vF1I8hyLHSD3dE9tlZQiDe8DMv7K
CNtPvtF/zdmCUbWYZbKJb8Jmomq56WPuPOSsMC+N+c27AFvUbH7fdVRduVUACM7N
qw/o+pCfoHTVlIkYvoK/BftQRwB7h4OLyTPqqBfh4mwHiVQfnEOR6mgjonIfJQVQ
Ey+8iA3p9jywWf5o8kvps47vwqyYGNh3DdiUMq9vz6Q56o8XHNTmfNabl4Z06yKz
IIhn4zf6ZZcuoxKdOaUQpBXM5+mm1Qb60hAg0f8D77xqStXr/HqCTht/EeG+0Q/0
mypjPi1xzOjGhMU4o4WxDTfRJl6jDjp/ExUc3kFriO7GqreTtE7WP6ihNMB5UElJ
z/BFFE0gyLOpzmBCNXFZpWR48Q8k+FhGsZoTyumm7gN6Z9oHFvjpyiJfngziPPcj
MYuAIM8ArWTOpeUN/z542awI5VUJp1vtu+tY3gHylh1k+aNJ3sEX5JsSv7L2THUv
tBCW6L3nHwstg2lyFI7ZoL3GfVrk5rQjX4A8Swc2X9lb4Sp9iKhH2fTQNYq6vKY3
SRBxQcOjcj9d946pVw/Y2YLs6cvWuQCO4jT/xxzYPJZ9EvSB9ylldfbfekBfL7rV
mvMZeXG+uQf6fyAQ6FTFUo+l7zyweqPWOpknzLEIk3BDQQrjtfA08RlOfTNW9oBq
hyOY7aSdOvajMYW8PgLJd6A7xOSdiutqV2nMQDjWsindDOV3ek4gxoicDd39naac
Hw3u0/oFfgCSI/KADKsCR9aqUuB0ERrplGY2Abv3MpA0B0NgDKC9hDzJfipWUiZR
CnUKm/wylIs4HBlkXYrJsXJWHsrcuebF8gJJpQDGOf9AUv7e0/S7BnjS6hE4+k2R
HxXxVUw9qR98r/8XEc/hw7MQq6FYPQjP+nOiaOwIGFzWci6XK+NkRkpGRmP5UQS0
2RTS7nLtzv9yYmdy0otp/jKQAYKF5/dhE5PjfFu2AWxo4ZjbvESMc4xZ+vPgu8lJ
7H/aJBvGfYV/Nld+lZ1GnPpZNjhKkppzPL2lH4GzL+aIrS95z+7s/MqNVkWLLz6A
IohuDUpWhxC4x529yPCpxz8vE21Jp5MAyV88Ku4yND5Dqw8UoLUBOnx9Kfhd0Y7q
R6yORlrpwBIN+kkIApQc0VzpdM43cHLHtBltHuB1NOR8HdVnehZKZRgjQF+ijvD2
UMjvFxHbyTAVUSRvjlf3cz0msLmeEtSrsZoqpcUQ2aHXKEd1DeQ3R6IpJNC/uxES
v99rW+gx7noAoC45w7vN6/Yb7dEIrp7jnbVe1Pa0ON+i+Tc3qWyMbNUBrg/S09Oh
MuQLrOdoKSPTph/E12zd91uvpZe20fVLRws/lEo3TFDwhP0k2o8Qrh4uTgiZ6VBv
ozvF0Sz8j8rWFcSnt8wlKzh5PqQ9J6YQl2V7XezSdQT5qajkAt7AJS+6HHF1AZc3
iWlnpvFjYdos3nRhPbMvfshewvkg/yRB53WeoDtdCh6hkkagUJHqOxUeAbsmXvjh
4XB1YwJQX1H8VKZJhig1IeXM3wS7DsjgE4qzdeDieKN1gN8bISnGUSPc3ovEJzhQ
GzKGO4sKLMmkWqgZOI6OP6suTdGJxc9VcSbhdU7ys127yWSoWaINEG3Yr5fRbJAg
CvofZAxlj3PJtFE/bgOyDzwd8E08uafgB1Ob61T2/GKaNVI1El/kLUVHk7v9fWpT
oIC120rHMU0sC2QWT8Eh/rNgWV7MBF4+5mKmagvYtTwMV4Oaer3iIZackYodfQRF
Ow/Z1CIt8WFHRMUy0qnQ1qaYQ6b6/ykQD+PoSgfYUcTG+VvDIDbe1jwqNWpKf0YV
LKLSw/eWyeOc7RGleFal6XUXiPG09hY6a3fg0uATidp/T3zYj9HXa+xbJDewOKh9
GYCC28dJy9n/zI/V8l3HQDVZ22SjKgqjTsmnFTXdlFRC/+NPv7Q9q1gCM5XKUVrR
n3uUgfdrx3XSfzyIe3mGkU9MYJ7Z3k6sG7PXKLfHTmbpia7AfqebtDntGd9Fgevb
U9A7GTMdIb0fxvykS7rwqjjIA5DK6siMdKOUJlf+aqyF98pIDFKwbGY5fj5HSbhM
SpkdSOrMnX6s/FbP4NffCTKkya57ipE5oqyWA1hLXBzIsujHhDNXz7okmmgv/2RS
lUwkDNyQ7yHEm0+saRbl9p8bTy2UXC1DbXv30oG+xWATliDy+rgFNDG97gwDin7R
wm5zz7rRpIjutxQusfkkdd+uj9H6D2IrdVmx+nfAFK/cAE+l1GVjyRoB4ZF2Mfmg
SQZz5WuOzy7uqIAdglAMOHF43tQ1AZpp3p6pmzJyha2oj4qWw48WNemKK3rvqqsH
JbroYVHaiNV/QhaPGA3SEDSjmmh/FZNrFOk8sKN6GMkS7w1AqkTCkxdMvypEab4T
l2upInztbR0ldWl9w7UcjhXHDjJ23+tvdatg+N10I7j4vCuuqgBtE5a/QrUIcBlD
eLWbKKkBrBT2dIMkwMhJpHeqhFra4OacXS2Rakmo5dUcEG4+i61BRCC8A6sD0ngo
x+2tH037rr9AMpTgOBo22gQdtmIdyU+K1JP5IGLkBII2nyv3jBkVRU8FVbzRTyIv
Na7yapRmyXmdqlgJrEtjy5fJO1wnW6u0NYGjANfhkhJc0vm9UYWKkzQn7It/GlQr
oOWH3ASn8txM9NesmDJkTYH0/aW9zbnbEGlalqhhk/GvnLvxl2asiKV3kBD+JtPt
sI5Le7I3jNgV/PuxMmPTjiYcRdUd4iRP0TlSAbz16bZ9FQ/Wa5pRVaFo3w4Db7O6
jnLoUqgavzjOqVlf9D6wkpUh4pm7Pq6DPDLiT0VqZRsdffxMo6S4qPywfOk0A3/r
Oh/NN5ICd/hjokh4vuvJWXPDc2UkGrrS+PJR9wmR+kmLetCMp3FiAnRg4WFpDzWX
Oc4bmlV1prNkSPihNIcUKWlQTEHnxc9Bv9zOQ9S9OCFYYy/ORl8/q2mvN/xgJRfu
pg4cYTqvsuCWAJAlKLTSE/3LYnC/ZFhNNZmkGR9S1Zo7VKjXuPQjxHEUEahiUC6g
E7P14fdHJNv/lDqFtAR6Bn7zZkSYS7H6rs+LEpIRGExvdLZZgPEBqdUudm+KwECH
efFC83l+ggSN/PUeFvIDiYkIoOHUsFuQnn1Go5ebYmYmWlLF3C6jSn6ChzMa7+kM
u9FmhOHJb7tuGD7iPDN+H3YRV40S6beLYx8XsQ34lxrvMsN8SIJoBdhATPUEUVgk
GEzK8s9t87fQDfO7gNnYUjvaFRHyROdFilAsL1gTWsKfRqPwIFDtttxdYSKFpsMv
4HVCpppTEzferKMN7nsge0qq87p/w44csu6+7y3ynM7botPFMXT9Rf+3fu82p86n
zoxQORsRGGWEdnhP/xsxOXPZ0u/OKvimFP841x2kLGGgEjUgF62yWY2a6br5uvrk
imXUqDetQHP8QvMyEUDe4r2gcRdZfNxtTZfjEpaLMVUhIpEtOHujo0O6OXmTHYUP
njx+wiAHBw8VKm5AgkLSiMcCtTJsl2vNQ4ceHgDxs1EpwChrI0bxtoSqaDgMpgif
GIUuISmi9rhqlVvz2ZYCQh4iypTp62VkFGCJcn9MklCrjDt6BHdj+Y0oUvJKnu8T
niN7CSdLuxyEcd9uQaGlePXBR39WkuANNZxdSeMr1RjSMDjQ1rtzpDFW/JHVWo2J
/tgAvwpc5U2QGb8czrqNJshNfzVZ7T9lLIhulBi+cRzjDuYLzMox1LdKWP50wemT
63zyZBH3NElzrhM2/1t+UgWXfn+rZcXwAEuzxUE9JnyFBli/Q+UyAmnkUPcSEy5h
Uj2/G8SVMp7QPWqZ8OgndVq9rNPyf6pmEsTu8qDyO5G3NKxQz7AaPfVvFXaDog4b
0qi+ub1gt2njZYn5i2ha6xXXBdOq0hpPkYxYYg3DHHRkClh+k6fmU77YUeVvgRbF
oPQO6ohUxrDe5vO4lf5ppNZyc/RTFhcQI7AvpxnGkVrzVaW+Kf9GKOZOcMAMVrp1
mmwM6N2JRzDUiP5Gm4rGXM5gnObzyhXDnEef+lUsHoem+4MA7DhLHjAaiq9H5Qa3
vKQX7P+HP1FahpZUiyhI0vsC6SQaGjjSOLrf5luwj8GB5pQzz1JHmG9QEjI8/Rnw
g1lLFnIB3NZGSlw/GAT+N2ns7pyxgps/9Ut9BK97yMRzCXH/+tW++SmkCdO6gc9d
wj9zPpOB/pxzhwjr9aLokeALQ2Nl2utgRC//TolJ+bCPv9gJ61VPwFmPuSLjB1Yl
bNXwVukVun85Dh/pqEbHYEGrSp5BEpW+mN9YqzqQLS+NU/Df72y949VCLNTWpQlD
eaFHjThoak3rhX6raIeCMWunL83J5w29WBJzi0eRq/qJLeYv2xVgnrv5L04h7EyD
8pn0hB5DcNWekAPUIqNaYd2qXB+VrYgI9qzRcb6wlM+ut4DevIOhotmBZ8Bjsoj5
8lYYbKTHWqG/pk/eh7Qzh9kiaSaxQe1pnrnIaRGz/biSlF9DSAWzP3YTy6pVM5qe
WwEIjTeUOZoEMb2ru3NXBdLxmaSgn4IxNQNCRTMWZ6hHFwQrOM7w8s4Yx8prWGeO
hyqt+xZc6aKrH2Nj83LLbtgeRhYMtZfmrZpC4ZfkaMR/PgcdCZg5HIOrLsXXtnYx
P4uPxA8XRselvGujuLz9NbkQuW0hy4s/Hhp2S8AvPddQ5F1MNsvYbWoZmA0qc0gB
wZTKrDs0FdVkN8691mLPUdkPFlOCdKNRH+HItunwWqRNM8bj0S+OCmGqJroxmUSh
GVAi5bmV7nuPT8+iKxjL0LHvCuvKXjD4ZLbxL4U0l4L/QtAe6BZIB/5B2ICy0I0X
1JcBRPVhsnMLzxlERb/G0Ukuo+T6OPkFONyoKsE8sxuTYESC+/m+WGP2jZbNnWL2
mSRyOpi65FyDozixOHN8blyZGKOg6TV0C8dLlA44jh+zu8Z3He9RGRCI2xG066PH
zZgcmtBcDM4Pf88A/bF/mDWSmEzybTqC7IcapMKQo4XFbuVycJCRsaGznY0tu++Q
QHsp03/9KhnLYLyO/DCSmY04zn+TrgjVmc/QAsuP5dSQx6iNYCUKe4kdODYsfqOY
iS0oZSK+E1RS3tgfrLJOICxoBcLp1eFBcHid38RbVK4A8zD78F6bhNnXvqSvQzIY
2b1ZX9VPLJLIkgA8bB9nZTIMfDKdgRVdBwXCYrY/QYOBSEGzpW2FTlfpDOcxZP/A
rokJ1wXWfB7r5dqWf+s/NiiN5jTumvrkldnPg2XLYF3FuJPKEVln76TKAA76s8eV
R6PpxBvc0rgL/pxPJItjrpih9/p6bR2FN+v/ehUCJB8lj1soGD6lYr13CKZtLv7J
alJcTiUwq6oKjfRJ2qMARNbdYwxrrocv3pcYe8Z6o1pRii1OnbO1BfpN6gbcpvbm
uUwVS8LpE89K3FZ2lbSgAgB3if6uyaakXWG2trlkp5Kdgmxdu3LZdYMdBJciEvRD
X+cwIdxBoHRYGjbolYs/dExPJT6r6F1LJrnNkt40rOZa9+yJeR2+87S/xrk761Ls
qJbQN4axxG6Kn0MElufT45VPrQZmlEpDTdE08xq43AiU9unn6EIcrRZ0y/dt7tPs
40I1zqCuOJ9MTm0Rq62a2QL0s4qXWekgaeYNOiKZka50v+Gx+WXyHfDlmMWP6UK6
6LKrxGyifSQ1mI6m0R7VdYZ/L6NpVtzIKLMaS6V/jyXG1qVsvGvuhmfxmZMfALju
rB6UJuZyg39EFaRTGWf0S5KD/LZNlD33Etqr8CAuLIR2LyV4ytTmxDms95mx7asL
EYWI3ch2IoEH1r1XB9IR2p54p0i/U/GxPE+xk96lRXIo5y1W9xdqfCWe3nzmgmD3
zniO5Y8t8iPX6FuSbnuvnQBDLCW1F1hqty7UdRvPaZ+9mdpX3gCqYcqDTQl7JKl8
4arKReUmCePxWFWi58R9wBLuWhuwktmF2NTp0Vyz3X523n3UZwfnFVT7mL8LK1Rt
fDCx68et+sPwQaFi65rpy+8S6G9vTIoNpCj5ngN5RcnSHRMwuMznddjrkXWfWY2T
t/Y0rn2WI8WIiM55Y1GCMGKrKpn2UXmcisU4DB6oHinvkKbrWBK5yX/bHwN6s8Sb
sHkIS1zTP0g06d621rBw7XzySuKwBwebHUK8gZntEaZ0kbzHALVGjf65+XIN8OES
LM3pTSxJDw4eL5d3/arFVtfIapqNjXwfj1+GCNiqpwWyTHZJxl6RTLZfc+1Pdf7I
WbzgF+dgTkYdKel8ZLpnDEPSisKmOuM3BB6NOtKaPjlChh8doX+O7U5B9jU725Wd
5S+E25W4Piuy+2dfo7M3YBARfMqnI6F/dVaFmjOFyyUFPeLtdD8k0t0xoNfNr6jx
tu+XfIdxQoI6Bxbr6Ydx4OKiY8beg8hckXqoT1D/HOuj4TICRddijRAeOl6WWpXZ
wuyDCKbnnHTxtaY0ULrmE5wo+ekOpHaHut0egHNXPGY2rlj9CW2sETtw/OYzRQPc
D69s40PUGrkl3bKJAeBkJg0KasHIdhG4A2TyqHcyqQmRdiypV4U5cXg3N5IfPnUi
L1LcmTjHDWuJdb1evF0vmq9Xy01jZ2t+8f5p5DDduP5vDOpSpAAshhDc7/SeBi1q
Ln/T7uyKTzAl8ISK5UoLUg4dUwtRMBpa42RFbG8VsjTBaedGiMEkmUt9H7K21iH6
qKNJdR429dFi/KWAsIqByEaJMpvgYBIlvpcldR4TS3am/mbnOb0pOKhZhY1wXnTW
NHlXv3Ifph+lnua/Wphfbx1CCXOGqlzWTVKy0UVFDov9n+5h6bS1aQSzY4kSQZYd
OBNyN4gV9ZsIcZuQzls+4kgDvL6FNhLjKPtEmHVH3sYEwEeJdID1oxDAaidt9tc4
De3CqkXf1cBOk/pIOwejil78dNbjlKWMI9hniFgNPzf2TWu5WtYZ4HM+ddgapsJk
4NmxMsbt7CBZG3T+eIXZjeMGKSp68qk9gPtAgV7ZRXVLo7zPmoQghaNbMa2PrI5R
cxqM3KSIdKcRsgrt60337+pFvRrEyu6FTOLHCamS4zAJOibc6UPMFoN4oTHcvsVF
GjtV8iCBZzbRFhfR3JwA4ffEdaeik2CPhfiMG6dPy23WO15WzaZVerDpS2qm0GE9
SmHM4S1AG6wXdK3NMYtY2ToKRR7mpdljOsav+DeG1Tn7f6jT6USpHJO2XvUs3Wpv
oRb+twDpYhiNHuuUoEppkv+6kCMzL3f06CMqdFQa16+DIYECNQZaH3JGdirheqh4
a4AG0FMzJGDXiPH2bWUaOXQXQYjJ8EUaNBg1zv19rPznMHiq0ZN5BOSryt1WcwXZ
/5M6sqh+lTvdjSCKr7iYoTsikg5U+nVTbg8+B7AqDx5yPJSUblRLmlGNL3zfWVbx
CX2NlYU2sgZwGQ8/ETmJDHoI5t28YGXjatG97PQmctWlJegXu+gToS2FSv64dl0D
USBGT1049/6LnmGWXr5kHO7GB3xrbXZ+qC1TxJbBY+mlOYF195O4NqZgQQDBNWv2
tw/zir9jho4fWEBqKwZXXWnfS9M7pldm4wyOWs+wQwSohHdG9I4xDHqW1KM7fUoM
lKl3A9Z+rVOMydud1GNqd+KPzgYwpH8DwU1mjrU4kOv/QXFv9JdWPgUnGpsFCoMb
Z9xZVONLEuhp1QmK16eZeors/BjPAnj04A7zhyBcKPIv7CKjD3EPBVX5/Bd8+3Yk
auWViueFwqcvo0fOStxmy59+CGSsmnaQDnhjnXKOamKOHp0tO/shp7JCi8XRPt/w
hfLZJz6TKSnhyhvv3njxOggGUWN5W2CcvPzFgZseBxMJ3IQDYH7B7DCfubKI4Ss5
4h21jiCuWqE6e5MhUCVd9rzYtqnnwkIEftqI3R1sWzvLG/kOi+xOMpXmREFC2GS/
Tg4fG7gkfm1I6GMHgQVzmRFUnXcRJzYa63tR+SmswxfMiTIx+BOEOE9tZdUEEVD1
KLzpClPWEsjblWVFhbAa4VliWAAct2kOKGaOiFx/RKas2DblZHRljmJGt7lAllcJ
g5FRlVS2+yIJxeT477twTAl62bEtygi3Jzk3FgUfm2HbqdAy75stLWjNVa8p/mGZ
/wZZ4kuMTqZUX4hZ8mJKkUQgM9O0EYO7tUgPO53Mili8viyoXlTARXbwlscmTvK/
ApALkl/L47P/bSLdsqfy6O4ONlMpbFJVH99oHOFnB8w3aZhbKmyr3toY3Jt8tpz1
RysYEYGzRz46P1UyskYp5MimV3EERTXY2liXBrncc647Yaf3Bn4UUYHOhXmSOUOX
r05dQIkYYzkGv7kXrgWAdj4e3PB06XN9AB9mghUNn6E+zsEpKq1WQ0NR2TLyNoAw
wdteJ65NgwcgSSb/M1mkCXCke1d/ztBQwMo3cKHjwHxfbd1tECFPkWElvX0inKZr
ZzwnVpHnMsTavXHGfpvd0wBmQU7P8188r5oAIe7V7FeNldbL4O1t3riSPJ1HfODB
u99pNdnoGh96iiESFUEPT4HVQpZQ1Cj9JEIlbpCCIcxI1qr9MF8+Qhqgz9Rn8VT3
U71nYdCto9kEVFPQ53+10vaCZajS1gcpQqlqv5Qm7qs6MX/CuXWih3Shy/9pE51F
tGSMciZ2T72FNW5s1K/OnyYrSrCcnfKOItKxiCE7arHR79GJJJGmZifPLuFI82P3
EId29BR+G+BPZGMsHcy5W5epRpzxS8JPhI3Hvx0o9WBiLmy5MmuwkXr2C7bR9i3B
JpeaeY0deexqGa9HQOcoeNICBxQmgO/W42b5Qqlz7UgnA1TGcjS3C3daQ2qlf6k3
zoIW2gn1nfwl7O31aVmW4WECRBmxKZefxR5Jd1H2FX9X4MjJDc+ELRYmdB3nRjbe
ZWr/Z/ow0CWHdihquumpCnNOXortQM3c4xLYHofTwNaSC9kKktk7L5s6pDLMnT51
n0JGeMkcFYJzgsCogshw752Jk2KFTURO/CJmMuMgzxwbGQ9ML/FUvSKe30kmQDIZ
sBo1LPVJ4JQXzStOFYO138Yo1s1CRMw72vmmrEF+HtxnYkoNlDLivg74WYRthPmI
NoDk59Nns++5eYyKHH6fAotck6L3pwlB8hRWLcUUG0bg16oQKhq+LCrEiPM9O81n
qsdVus3f/3CH/BUOBXZiuDUTmiFal3GZ2SYVDmLKwSCLBHYWsoDNdw3+YW+23jBL
Xn+os7m0vtM1hiTWJeYxnI7ospr0nMp+Ey5DMO21Z8WVpjpuIzxJGqCYQ/yHGjJa
azQ5xqOwGWZg70O2x5hKkTK6PeMkmbpu1S4OfhMN4+yUn1RAxoPUetL3tqYKBEOE
uxhn/nLesIS95RDKlrLdr+czCpWNeXb0MdRxm4PY2BrsdHszBKXFUogxZXKVFOK/
LuxUveaChKuXBeOxRwpGO9VL8X0G7etMMifkPRQM94smfOQ/rrUXeUEXpNRx1Dzh
XJd6Jcut3HlmoKpr0U+yBvZF+O4yPrqWxG/YljAa14tslzSdiuwdk9Crdwx95I2t
GZmI3zLy2D2jh/LgqROqZfCMcQ1Bwbz15niuZeuWxK0wNb64sAIDXVcFi6NM0xzW
FlOXd19psAHjsV+6M3ovCjsQy8JDGRBpyXGWl9PCPl6fx7CKVQKKzbNdkZ1m0VYR
JUOCrK6eMM7Mn4LlLeOS1TP2xwX+9pazmvhteS0MuHfJ45T6XQOBESsQRgIY0fP5
/P89dy+E+Y9aI+h/rd/WjosbQM/7LU1f0EdUx9E8VgxDF8p1iXLuqBdslPwIjJFh
wgp7K4/lrrdpN/gVZrY/sl+kChbBkvlZx5AeVH3S9CLnqZecyNcOK3VUNQN3kSNS
2/gXcddbu+WZGRTHKX4imRxq+vVLfSGTG1fv23qbZAFLVqM1AZ09btdkJnrgXmZ2
HxT6LACD41LGPSGxuOI592UyaYL5NJV6cOEb9CKvzYWFmUf1QASOSieOoTVUhkjh
Op71IaojZP6uuPJtMkTRhG/B9NVZvYFmO0ICHjUhsAW9M//JhWxsjBCYUxZ/G7JW
0F/eY6q92sxyYjbmfwQ+6Q7BIXtLcv0wyr3wkw8SPCLzxLnkkvvalQVQkn5qWPNK
6hpicUIMaghwiRgKaTCp0DZwcuBhpQLpS/xZAGwXZ/4XHSR01DvfTWbFr+n183dj
U+URF+giTfE75rLC6kOIsvy5NVstA5g+8c2iyllPcPtUM+aM0Fdb3JUOkZpXPmJF
jZC7YnZsCCIAiGg/Ls3zuYOvvjcA6aZogVZf/k1vWUrW/qDLl0UACEj26bKXRo1t
Ne+sUUwsr4rJhk+xs4DBCtMMiowrU2arvMgE083nHJhPkchORvgq5/pNAUQ617eA
pdskp2MsoE77N5pph+W/aHfOkkXwdJkK7ys5Qm6p+vOza5l/3nS5qgTLn3bC9FvO
Mf0pqxzBG1Q6ExL1dRKhrywH+uLNcqEixcUEcGp9x6noOpgHkrKD4uGKTJYza2OU
CemJHv184oC7EH80wUuURd5Fyag+K3moHIwi2qB/hrvyliuV/Rx0gMCselZxqX48
rT17MIhw1fCY494fcoqNXNnNDpiZcEE5o+An3tFQGo24RdyfUy5NiTSiCGrBZUuc
4XjYc9s4PfrbLQU5jKB7KXG8X379yxuEmhCgti2F8ucLULNcbxjw/v3KmWvmainS
JOiyF17oKynd/FFbGU5ybzOfVBlu0l2njcAi8kpDu47WD5hhmB/6ipgnTSecfSG7
+o6AkIAcQS6q5vyIwL6JHoFMS/yJa681l9seisY9tbldAbgO8kjiBBxebAcogn8y
XeUzJZJXWW2eC1ZFoq02xAnApsWDc/GIrtlNlCh1EdF2oblao5+wPFXyWP0urEr+
CVBgs49Gdiin9/2lJbZCHdiF+4cQOhSan22I9JGzmsECHgWckhis9zP6dc1U076L
RzX2uBO0/tzoylglhlhFN8FSnYcTDabsbKOTox7KogHVbbSsnqVXCkETZaeu7Tc3
fCTdPl/v/TaQbD8uGW7ZbOCiZb8Ch0OOysqoLF074rjuqKgSE0etaBeBTFKSxQjL
A2OvdJvgWQZi58ZXHSe7kfUcW6jiRxGitZ9T7BLuheSIiYxdtGtM31n4Rn7ooXwu
hR5R2DVrKQrGvYg8bSPkRZcuORk6/+dY2G3fJlfbuIxAExaCNJ/iMXfZpf5k05nN
jnLQLmi4//8jHx5FaFrydstMTQUd0DudrYSYckmYXW5WphmHsvfHoAk5wZAiEn8q
wvcIuAJ43OlkG1TU0HNzxmUuPvlK+1vcTUr+ChZ5nbZcCXc6HXpZf6qWmjD7xr2B
BbI8frQYsUUV5WxhOPO0rXsoet0lZJdXaMj+L6JP+49+Wr9Iu408KPEVmMJVru15
W8VzjB7ftufILjSa8RaXTs42gJFJXXTfW/+lQy4o8xw4oJ5SomcCvM+V8RSjoKva
bAMI/eajawBYA6WWcJxTWua6sQLu7Nz2AsM3+zoc7ptMhUrbDHOFl7Q2IK3J1H9r
erINIkbM8re3UHjvNKCcW7Ue8EjPB6rDqcS0b3vliV9XYcYPS69Km38eLVdsoYp2
DoVfIIHwU3o76V1bPyJDdQQlnt8ulFYBbIkFMzg3+RmCSxqQmCpLsj07wR8Tt+8C
dPuAoqqs1p4Fff0srFjg2gKswTCl9Zklhqz2TbWsl2GwQC6bqZZiPItNcvdVIAGJ
3QwGsZ77zmBLRd+/vBTPOtIYizFUt5LmN5mOm1xv6WOvANoq+hSdNSpMkzhL+0Bg
P1OZ+oTEZ98e7tfn2c9FWHSfebntcKB1MV3ntRYC7uM5G1mRUx7ou/E0poneZnn5
8AV854buNDXjYaqKNW8AeFnd/5NOY3ggsk7uRpviqlfyzeoPelc8uby/hCMZcFKQ
89b27GL4T1zSCqGInrI4941Lgi8QL7/eas9ddWule3ZSbgcsdWVYh4EreEv+5fzU
oMtE/Kpeam4ABJkO1ztmknXrncPIv1Hg7HTCojt6Mp/eQYA7WFuA2JIi9/LUJ3cx
VhG2dByw102uyHqTypZNdVxo5TqHQrFITTR8N8UKIS5GywWJhEjsz2edc/GkNmW0
ZsqVHvJ8xceOzz+PpiRf12mx8paeRv/bMmWx7kPlGHTVDvNlgcb3eTVHYvM9bQQW
xiF3vnLi6PPXmvf7rRrgTCA8zvFvF7hVSglF5FGLe2jTYcoDII2dGAx8ZAokOBBl
0ugEYs9fQ9UfBt4ePwVvm+xZpDISlP79kHiw/JJ4mIEd/5giCMo2ZUMGjm8nFqFw
ePfSgIY3xaWR/s/M7bn3Ol23ARMggzdmAVENocV3k1lP/Gz+Fea1+nW2zycCI66L
vwGvo0Id8ai8XAA0frbWkAMsegssGkizb9DRfGKDpnl1g51i7zg6kGi/BwaTVS1/
VpElHMcVX20T/jeG/Uk47QYGtT5UMACtp543sJpOTUznJK+LMFX1/QhLwknK6RQo
0GUXXgB5oeaLO3Msqj66TmciYRSBSIVf9amk//tBQpMoJH1tJkjqecU5NHFXDn+B
cYp5cDbqV2PDLYN0sGMOdtZP9nYiPOiYGMZWUWfPby1TmooS/3F8cjK1pHZ79HYC
dec9ejRSPamMeoVGgIuVnNNTQ00Mx+PrZD7qJohJWBLoLjgb1i2jXhncPDBRKFuz
J6znktZdPHQzQbz95Xvj6rftiujJ+KOaVS/pywr/FqL8qpyDH+miT44tQOGrLym9
FvDGSFnrYA5pBgGw50fMRaNQMTZ4isaWfVOeMM6Z3VG2F2/f325ZTMRXSsy9FgZB
f4Zq+I4/ve8MI02v2qS34LqMSFA0BAyqd7353RsSe5RcTOqrgnkygXg7ryeKKBYQ
NbICStpR5ht8iEA0z1VTWfhxs0E8EOLeAb5yeCqV/8idrUNzDl2X/lY9KjLgmZ3o
ZxGCs8hkW8JWdYmwLEDVskWGKvhOCCDUTFCMDj5MZrLeMZ6+welcoEhrDlwXYN3t
FJwHdKdOLLm2/XGw0/l9O6ylvRzSUeVGMl/xRe8rc00BDIaEJ28KxYybUsTjvtJU
KY+NAiGeFl3PC+uaIbTUyJIvd3Vx9aQkFdz1Lkg1j4OsDS+3V/ZvotAjT0asfkkG
Hi/PFYk0VcfQCHQRP34+QjnTN48yt0/e1JTZiiSXaoHYPzIG1gYijWCR/7lnl+FH
tm0c2LAwJ21bDwSisZSWoYSeadW/RyPb3em/yeV2Nk6D6OLLpibdaiR1oFPf2fd8
kBVpDmbVABqZMcRYe4VoL0QAwcjkrPzXQvLcbP5/2u9+yaq5IdIA7/LIKUzlAwKX
+tx6GWIJUdpfDkoxyCv1wz/BlVDKnei67wA+HwlhqWMCnavk7r+7DDKqXUlnwbHh
cZQhsHX7FTTqxTEaA3V1rJhi8d/KHqaEkX41m9XseDu8xoeS3mygPlI/kQ0olqJT
35dneLGVCwJvhnuDygThxnQ5/PleMLlWlTpsqAQh3lkoziuD5Zw38rxRY04mHAzU
32uWmE1N/AfiFnG/2NDvR+fjsmEbrF9d+W2yFJ078x5dM3C20kvMHjbi5O4mkF0f
PP8MWA06UogIc/kN3O/ZPDpIzNoIZ9f2I7IFyoo6cyQJjI7UlPKHJRKyljPgy3C1
SAUHi+9b9ztrLDGS0S7GyVqYb6LTHYeBqsNGV6lqg6WyE0uIGeiVBYiNPCtPXYy8
kef0RJLno8MIJ8gh8NMakSONU2rkZAvLfx4T1lQB6utRV3ZkfTUUYojuVC2ta1Cx
h/3iN1BMh9f7R1e4npGa0J+Uz6zh2mpxdvzuMfuEoALzg7WfncV7VDZPLpW19RPg
eXOmaWzP4DQ2XNaQtB4qDgsZvCd4k3OSjQ65HI+wNybAc4SVtk5M8D7P1kNuDs16
ikcmDPksrjZXg6kcfPKbo6C9mfUCvbDC8wDuYOGVMlMLCloawLR7javJ21CLrxB2
2W9ffOYwl48Gr9Z4PBh/O1eCnB54FLs6wUO8HTOG6rE+MqVvpS4wIRMRFKkX8iiH
G4S8kfl8hb5Q7dHu00r8R9270xsOyteoOKJ7AV5j6wykZf+vxtaAkaPkhHQ4ncuT
eTAbQm9TQHdrZNu/Zr7vEdn0Xs4eihplbqg3/UrlNnxU/y+cFWSTTnCoypIm5lBK
1uizlesTsgKgREREZNIZEKF/JvH0ObwZvpWdbD/KQVCII5K/3t9fWhfFCZavzaOn
ROew3Ac6fBJGbzaxxsUgFUZKS/m1emyGDjvW8kkPxj55c87uvV1iCtygyFYgJcAV
QY79aVpLwtnHwjaHm+YQeNXh3a6k1i4WGkreJ0UDd/Hoqoex7AQEgHf7dVI8xJXf
6fDg1EwnoqE714+95/6vyI9Y1j+CtpN6Xy0s2SmPuNzbav3OGX8u1K92z+7PAuss
HIeL2BqBYqsqTNDusJwkjgVlW8ICUfkVC0O8ekaAM9wIsp8G/Tj8xbdOrJirG3OD
UfxxjhoG4Fej8/1sU/zBNr9qrk86/h/ytBHWV431g+ayY27Q4yeR2wDl1N8pds4i
0ySsm2MwHoGXJ2PTHheuiVinho6VyEYRcRGvo9KI+iXBU1Bgnt4R5xd/LGRDjzni
gWdkw6FMJ8pkNOgF/sBmvt/VAPqGxxwlCJTEacdOd5n5ehxrflaUXtaZS23Bv99C
RIFHIbqLNvKGUP64pnWLfb9xzeBCIa76ajy2NCNaNrNrlRIdyO8IKwMUp66FLYCi
0YH8JVmrUD3+R6EWr7VY1GSBJKhUudxx6VQ3FSYEhy4BXCRKrsxwO5uIQeDGZwc9
pTp1Np3JmEb1Yi/sq8GnHlo/evF6S/xXOhLBgIqkSVgf+GP/h8kIhwzDmUTQ6nbc
MUlJFz4QskvJYQc8Oviur3wHIoK3fZZA21DKvsLrfeAWUcVYRuksD4qNn5vQxhkz
z5efhbgtWdivbEh5+xMUva2g5JqXjZATqNKF8HcHiF7n9usDkr2r9IlBpREEvEJi
xHCg5WyKdayokkTfllFSIOT8L6sBpGD6tmbLqFv37J8PxpBqEuTYSEQ4HzhRzyQt
+Pqx7rV+5HWzGynEOckYV/A/AsQEnisSFd9Y655QLM6LZy69yoYOWqgUtjXmIscX
kW3QwYbPuGbAFpx+KKCeyzGC5SSOMH7wLCehu8BcAC5BzbJIdugm35b+HtI1jSJk
G7qy6k8leT9cfxidg+IvAjojYauEbNzRX+R22t4CfpTy6Cg2OHYrqspaeetfcAwy
CFlaGi1LNr6iiC9FwBzlWb+ygY3A1vUyFQm7S4mf31Ya3AT9hJXw5lEUZTv8t8M+
bFAU8T4Vi/Ez4WWeRyfko1uvenUFjDom6xyymh/77u5V75OUIHuBY1DC0ZDrD89d
KXd03Q0VJwxagzQBTzsTNm6hS4jVqv3DmHwhgT6ZAsePGiMN7rXnp8oMxjkiaOt8
3OzV0BJABIlrLc+qvRLa9SCk9g1GLqOaqPeRJ6VtFkYd+ikZKU9ckf6UytdeZXj3
hJ0KV/qTL8mcHwsuzV6uR2+mQDqtmuNyUN4d+Fx3HWCAG6i2JUHerhsVd/uCtiTz
p6cnbP/0dC3/P2E5fb+B2axNWNQEN7z6IOEUjde22vdzxcogorEttHuXSiDqw73m
y+Ia5rhrpGVq4xGY7ZjRFMUfyfsNsa3nOkde4FG/cWdxxvmzDLHS5MHhRKC0bm4o
WhbypMMXGdfuEGFyf7//64hoby8gP/A+AF49Cdo1hV9b+w+ivxWFBiJW1P6c04aH
rbQqNXHS8Yt2wRoGpvKD4bbsajJJBbxE8THGi9z5n74kZv4OHYxEGFgmUhCWoz7i
GaGfVX4RHfShvoNKI9OtwcCIP6PclnY5Q3nDwKMOCOejY56lfb8Lqe0djgroihX7
DmHjkUOUVjKGW3V+26moTwym/oloDwKb2GsTsAqXwA3l5/Wrt0FOOaNSRMk3YJFW
J15STD2A69B4iE0odIsYkndLvE0ZmyzPCzvj6uz3SrR7fcXMT57vxcg3SGQ4flBO
kFQlIFqoxVoVf92gTmfaSHmB7p75K/gJKxJujOBHAgcqfbk7r8p89yK8Sm0VVh/N
1aY0p6r8htd6WVgZsc2jz7M4LyB54dt1pgWK5YsOlhYcmxYxH97h6mI9dN/pfTTd
zBMDsgApRbxVW5JhtTou20GrWzQU4jT+rutQrgTL4HLkkKNm7ECkmmqhQu9gLFWt
qn/XWWkMxvLRbGD5Qd2oDGbHNCqJusX4SgqDrpUE6TBEYKlUm6qCs59Vj5MwaRdm
ubPLXZRlpcXRAnWuxUZXxg8mD5jsAC8A2IHMknImqO0K2GOLPot6zyOATsTb2kxx
G6rU8JFN9XltMAHpvs3XVxZ90ouVx3ue9Kz3C3OLsuMMBZq41JN8OahXrFX50Vgz
1z1Ieqh0XSdvDA19kuCIOiWWJbyOoehdhdmVch6x8qjkAwxF+zXZhkcmHjEqeSko
PgRmi1VjOe5iESIJVs9o0SApKcVL/w3wzJrd1GQ6dGaX8HZxhX6umCeDo+B/PBQC
xoGSc/rDAMn5jhEY6S2EAh+xv7vgOkIQm8OTBuPtptD2BO47MJwzb0ejq5BxG2KA
dLVP8/o4smh3+0aq6qWlLqiqL/MAtrsr3fNm24NG/8tWRmf8KWG3OepwL1qeuppH
9avDg/rJ/U3rRJxsC28gO4zC291/BS838KJ68MoHQilEiMj3WXengpjFUOSQeoKt
CbEFRYEmoXHQe2hOEG82RGqmTT4fmVWdJwQ5v9UCbX2YD9I6EIQbmbrbOC+k92IW
F9SPKbzirgl00CqpvCmPxUsJCbjyClbKT8IDkXa849GV7sd4lda57gP1/rl3C7Pm
K5COSrLwmM7tlOpsMD4rOkLmE5IiUhY4YmOuGERevzEUwztmMOEi3VyZfTcJQIH+
ExvmpBn6SgTefas6PrKCCVs6cLqRLBJ5DUmuYBzBUblknsYJLjojyknuoM4W3m8I
3x69Wh0oM5HsfmbtrDEkAykCtT583/b0Ji5aOF4Fm9B6UB0QDak3c2TDM+CHODvf
vvJCkfF51i2S1c1ACe6BJk/hC3JAw+XBQQDJXUJ6cniCyPXL4f+Xpaso8ApPionh
vyHQtyF+X0AjIe0pVXnHgospziyVFiteFwtWUt7ZNl5v1XPgWZ2rjrFwhwoBKIla
IgdDl5pXL9TvFCqcf0MGT1mbvMYRm0dQykTZ/KuUsz+FBfAVaNYLaEa4nIVPZ7df
szhlnTL6LY0diRTz86ZKaW+gT4WD3TlXtl//mhGLSmH9orLZWFLpHgyyfZJAjC0a
52BxkGRaB/ecMEDzjUyNEXkGvPhs3AoDtMrW+ECmfyRf0Q92Q9pUD7mrqzUTDBv3
w3A5Qs3i+TiFQ+LQMN7/mOjegxs4WmwIr4K79FMmPeX3MHGwT9sE29dNuma6X9ee
CaWBwPcNh2myIZnsbkEqvHibUcxtXZu4Ym6HzmgcRJbVWO34eFwC19FJS57OhsPO
M4Fhxt0hlaGJDqPHZo7CovA5ygjsezZK/BuNPaMN6AgOSM4pe33Mv/W+fPTsmZD0
egFrgz/8G+iIvVW3No8PBdCPhccwteoOr9nm8mE0W5+7n5J13InAxgFNlq0JNag1
sqKyKkvzcHDk1X68pTZ77KNk2GZW0TliPh2+qjjqCWyx9BEzvzs0Ogq6PCz6I+Q4
J97VvDg89T2WX7cOCdxR0Atf1XQEjpImDW8FX9/ZjIXd7yZRdvDPNLFORytbN6lr
i3cgiMYeO6a7gan+Q00a7j+J+8hA6GpVqNRf8TNUxOcJR/f00zzmLDTLBj1CrbcH
dKjXckkJDlv5+gEVumaz2gZI8cPzvnEpeF2oGTJwgVq1d5ing6RFQTRRXFCUaZVP
yRm87sdTGTdfHW8syu12Q8Y68C+xZZa1dhGV1+2vpFDO1dWjzdM9JE95lupRnSMG
Vu4Qcdt2Rlo6W+pPc8Jfe8g2PeRLa/V6fJ6RyDAVdUWMlBFjSd8mHMRqd0d9rO5L
mqvGbqNfUzzsT2C/aqbtVhOf/RLjq1BZNwNDjcPmsUq8yImiWguioRD3/uSu3xaq
CO6M5Bc3pJ4v2njmpjK3pK7xJw8XBypApScfAPtKjbjOYeoejPKtOfulDsflLXwI
GvcmJfJbVroRM8Q9+tFEC5fH+N42NFIenmJ0c+HAH4WHyzMKVe38HAoL/iir0J0W
Teb7s6OGFATiRr+Yzka069gObpB9RiCU++sG213t4bBco2gaUty4KI60CVaetggL
tqDiwyHjMWq8gv0BP9lREtBmq5pya1qSMQGEaVYFMr8KLsJSuZWpcflUZPFzYxv7
Px1stRDMRCcVtX1+dtr693oMEHuPX3rbHAUoc+kKbPXu+ztwJ/zAcgCduDhe6/+p
t+sHR0yBhmvRvYrbSJC166Why14PcgKDw4ajGxHo8E5hl09SPWnyP7w6IDYAooVT
7SdDvLVuRyFjunxIXZbbtxkrNF8OMWuggAijHR0FkbeTzqwxYcvV71smpAMJfRkB
j8+cv1SCKiTFugmKVT9WPgtZY7pRvOJ2jJLzo0R4NUULHlxEuMp2MgnNSz56sXzY
lA5B0SBBNyZjAf8pmNCuTO/GxFLDP6ZB9n5yI0/sD7AN7hH8gu7yb/16SsUMPoV+
LK6gs+f55eo3jBiec0MJtfIQg51SLnR7r8FqNI0j41R4cubzqVnBTa7OHrScyQav
P6I65KJhmEZ6JEJU+7Au+5lvvYGccUfnkIciA5sI2XQowvIl+w44GQH9Pg+8zi7d
Z5z0a5Rsad3dDuuFhFYu1ByV4Why9gwLhUhE0NSPOQLEbaNPMXxPLqVflFPh0ynU
yEJguUxsBAbw9VNqt2YSk8YGYyU1mZ+ia8K5+48hCaVR8RyGZ4HA2ZSjug7LAnuS
K7EHoD1hjeEoC+lCIK/6i0c+JaNNc578fX3SJwbfkpYvPtbYSn0G0Hzws2UbT05Y
HNTWmx83SCcQWn8DXyXmLyTGMaRa6izdN/JszfZYm9nkhy8/h2IuOP2taAkSVdB/
vC7vgQenaIVtf5uTJMeSZ3XBPF0MNMnDzV4nRvOH7brXgBWMUSqgYDa65iQEEypI
agIVisvnY/mjNC/uns22uhDDcrF6n/8U9vpJuwVNSZi3HtTKTwLHwl62wVdZE9/S
qyLmvEWDp4j9mGyOj5c2zKDW+Olzrmz4hEanyHwyWRsSEI20Ijc/kJhjvrXXzkA7
KvLoEF5GhbzimHj6E8Gr+chCP7uCMm3IlZvNDeRwJRwJw1oGUF8hhg8SbFL1sQv/
hnlKsmVj+4oVs2ydXa+eFCvDRHK3xV2drMTGN0SA+6QgUS/IlvfaAS6pBXmuKjIo
uTomvWQ7nKwFtEtequ4BGqn/ZWF2OQ11Ej4/Kpq6CzAizpv9ISWi6AINQvhB5+k0
kTI0c9G08RFi4j1bhaXPQauf+7rqf+YsZbMQwir0rWZ4qsuRlvToYroRLEW1NJpb
2/k8QZnS72luelGCeFjXcXjiAQXN+5AYRn9/HyGDs3NLnyIqep/1luL4bnEXs5XN
MMk6ZzEmrg5xB4Q22o4l3Z+rSsCIqFuRLedma66kyF7WdzVlM4i4klxwmX/TX6KS
Nc5RihAr2jJmiWhugQ6JnRfF7aaKGQ/jcO2pRD6AfpCqWLlCgCB0HUSAcKpK50mL
yaKCElJ2+JKygmsVi5jL5iOvLofliAj2uCQFG0ej0H2uOsOlQMONxIkKz53Ne1HQ
oNlW30Xxlkgx9RVaibEBK4fCK11ZLokoFuaVYaQydXZsOOKoKDsf+YTA1mdp4J5+
Sj7hWDYcqCuksIs7jSt41BG1O5Z0NtNJt6jL0snOozWuvAPVU1y78Xe1kH+CA2Be
5h7zIZQcWORPFwvagYMAiI80b0+ahTFVqe0x+DUIMCzQ8KzfskFgnn8tbMW8KJ9q
Tua7OgatiZYjOu8GmQQrIalh8ZgL2RTuhE4nZj3ABTE3ZGkQv9FMHt0oRw0AyOzg
sg7LP58PLw7j5r39z5Mn0NII/8Jz4p5dRJXf6Ht3SmgHoJon9p80GIr1oSzlvZln
frtFc8Qof73gXd/aEt78vnYO/I83BMWa9aPH/YZePYwHqD+QEt5pQVF+IhoVt7NX
70QrZ0R4FmLWIA0l25ifnxeLCpQkiK7Y07RHkTp7bBdKxGYUYcQe0PrCQecMnmwz
DJ7XtbsE25Kqnya1zf1mlCJxuPy2Ic4JV+8g3GIN2dTjFUdbZ5vyMsooJFfa2zTk
jacsO7iCG4s8KV0eMVQbaeCyWG0EbAu9YYq+qqfY54BOzitCl95y35OZIvDRw3cX
xmmUBOQyfxvmuRYnOpdumi9jMGKkKwtGsl9PyzfWkvXFxaXZ3t5OpV/ws5jbzw1H
Uu/IjweX7xJByh4r3Ln2JQghN1pPal0pxNeiWN9Glh3Va5sLSwTF9wz6/OnCOth5
Ij3V9997c9eWg+Xv8kPvRhjqoYmSecEWv91M2E/0ouq/WWcGQOL6B7S28jcJdXLt
fyugpo/kcylT7HwOTSrX1clqeQogkYSDflj9B9hqF3399lz5drm/KBsa32ImpaFZ
oiSc67BiNUihyYW0ecHwn46GSzu1FyPTrkePIAo6mhNhlaw3tfTjA5PlXC0ouVl4
v9fisPIN0y16OqIu0nVSWiluUufmH+cqJpQQfWi9zQZVylddBRKM+JR8/pvM+9B2
hacPnE/hbvHRTuVN/5Y1gAXZXfUvJktApUBqGSfAFcF6Qpnkg0WW7YBoWRosijDf
Itv97v7x6dcUZHTJdM7q0ySrPqa7yBjsFtD5NcazP8306HeGL6EVR8y9cnxavDh3
lF7YV/yXKo22wdtdpDzVcdYoY9PXvf5GuPF1rjYQPTR9T++AhltbDbkuPZw6yZze
ZXZfLEXLi4IkqMKF6vNjLuzcyIcnypdox2iJ0Vzo7vsn4ZBEEI9CIGI04yoKcT5I
J786IYUhYDEEFJwF1Knqc1P+Zodh37KhXcqygoVa7/sCKswDi77zXt7IuwHFxstI
TgJ+10g3SHVe5ONvRPN9KcHQOXDv1uMGhcYMH31lJvbSpQBbu0OZdXlW4OAbmo5F
+mm/WUWihk+pDEOx9xp5UVIfPPB7dZ1hQoktYNx3o+D3V+BWyBbV3mRSTPNjLDaa
2dmCPbe35dGZ2LfXPCGa2XthlHQ4H+Q7jGEHrnwbTBc/RSwuq/oQxDknpvO2oczV
Obml7LGOfWEfRU3IocS9M1hQdyDKK+iEYFKNzJkl9m9WLaFEdD1jfGvYH9hSXTXz
pNEb4DHFsDwrrRm3JNUHuVOA2wpGGmT993dfXRsmRDsRVHvjePMarene3gqWs8Nd
ivDT0uf0g8IBFGyz8Ktr8Q12Z6IqyY5wStaC24Ke6yOkPHvcb2MG8qpPjHyebZhb
1PDCyXgau6mMCZcCAhm6SHoNRmPkz5Ss+uD0azOmCD66kp+lJi0pGCQM+kqe7ang
kdUvCnbHpAI5phcTHGNtpMHLx9RbWeSPmROHyClLNi8EmrTkjxRo/C2GTKU1fsOw
vIlYsKk6OsrdXUwXaHI6+lBKmJSl6nOVXnbdLDn6vOqabadcu0pZ0k0BPWg6hNgV
/OpTYWRYooyWCNMY+lkLK1Kt0nBuwjdCeV8blgKUWrn1NElggrnqi7nC7d2sVIK5
tXnhu9WUYvBFm9Kl2n86JaDR6pz6nKxTSXwCQE+v8HFzVVOsYsqBzNVVueCDCP7x
n4JVBcg8jNM2XmA0U4m7PLOueam8C0t5YWe9po+H+NV5DDkJO0YqPZirm4CvuLcI
y3j2L7Z6rAbQt2aj/eKkhvbRAo0O3N5gvZKQPagn47x4wcUcFOFv+JiV8bcM366+
UfPWAI2XsNAEw4udxlTOYNNsV8h1RrCd25+2+EUeO5rOhxbed9tHPmT8uCg03S22
yNkvG2wHJbmrRrfynKMuHyV897juU8Rv/kyZbNt8U6rBBXUlSSG7gOVmu9KyEwQS
e33SPCqiV+PmnhkBTqtfD9UFNfMLNUAswAvLOtthFYP4dgxmpIRjU43PP9qIPisQ
Xi392ulKIM+ighupddhLknXydhNddmwX+Ff87G+lPqj2pPcIOUDh0TzNNsLs+gVn
+bYX/63kYhXhQxzVh6JP8Y5/DTbmvY+gdOHxK1X3sSwneLvBWRwNxV8M5sE9K6cX
9r/Ufu+Kv+UVt5TTiT1I82tIXC5EGVUzPrVjojQMvtyz7UHLCFfvIctotmXf2xYR
z7wowbZC5G8RbrQz1uAv5OwBaBuGoXrgR78Dp6P8tCLJDajcQYGjOWGl2FDpB6Kn
9D2kb1IzWKKThVjytV3VUcnuxuUbUTUv4dSyLBQWhudR2IQl/NVzb1Dd/0Tfc0ss
DeFlL5e5lnLdFevJnaZCDpSYbpyM4PN80IZN/7liMBRZ4xhj2K3asIrIy1V3Zj9C
UeBMCH7zVHIb+jvm0yx3qDiQkKEoRNCm8dfM0gM+qNcDYUQdn7Z6NE5UNECyZHqe
npb94pRER+ZDxqr1DQIvNbSPbv5Mgi2QAKZ5DeO/Y5mwrTKB59QNRQcIsVKDLVpo
NBUqrfpBlFIYU9y2uAehG8BoFmVI5wYx3N76vaY8dHY8OPjhESn9O1qmCb67nnQj
AfSD8aMmM5ZNoQxvWPG/KaE4ujXYsg0qTF0/zXRIgM7t4eBpASnmVBijT/MxVu19
qB5ZBUUy8TfiB+K6/D0zGfg/kLehVBatTVWrgyyzPB6L7ia9ncVyhPme55GnwAo/
lwghl+CSguTQtutIKgb8E8bQeFRcWPJ95fJsIcBuNRsUtcDcVJRjrHG0HJxlVB6K
4fwl+z8hS509g6q6Uxvd0irlNeM0QMaQ/MRJuVm++d9H9koiLYdLKdKxDXHzRlsi
vnUx2WZ+fgzZ6M4hBNCTa4ZTD3HNp/rDTL2aRNNpbCI+5E0RiNeK04eWY1YAar7M
GUSk/wpIxyhoV5Oe+1i5XmjPVM3rmHUPZw3s0VL44fOKLSphI0jGpJ9oIGp2k9r7
ZKnm31azdFyfzXgnYFzYsVg6Wrswev6s+n+1brnc5T1YszBwlBBU96vRw7PDqDkB
tjC+xNsvSO0LzE4mki7Wqm0ZwlmLjJ83hIgEPjXZsLjRsOb6uh9zWQiVjri3zCr8
sHdsHXqfRCNxd+T6W5RGwAjaVZjB7KAa8of4ZuVIYauJ/nZEF3iRWNXuzziQuR2T
RduD1ZtUvPV/Ey1nmBZCw2ZBEXfCaiKU86R9k2qxcARKv937RPsBVnr4KHenghMn
LNc0n67ZPRvxHdHLYW6ihq1fCPxkmWVfFYdFpkAvytZrS2xP1Cgg0UvJUN0CCjHA
+YPPLQ+e5wVEu0uoqzCwcuqXgH59OEVz3YGf/0Bx4xtiajkjIt1YkL614Rde8MJj
xkUlaXn4Xy9bzWfqZuoHCZK/BPr4WY7J2bl/YX4M/vI3fQLRx9FpSXebLg8VVVba
WNJZ8zx23tf+Vc7+JHFl92FshS98yI7X4FTMXg6NuY69lX0P1qq78iU9KZNcd06Q
D6xtf9vqPF/qMr7DxNCR5Hs6DwYcW27A0nNikjMiqzDCCgrVJkTyDUEDc+uymNOL
fzrcC5ZI3APYP9DPRRDvMit1T0DmS8SSsSn+lSZKnhUqHe5EOm0W9w+3jauf0skA
nnZCh5cbXyjkTGPGKMuh4Cul7RkiaTj7m7JtnQg3eeZDAJRqV9C2xMEBg3JFPv1p
ECvRf6mgvxYS7jNqwRWyneEIxpo/SpraM2R8HXZbc/eEIT+AAWG1jpQD5EJh2e4u
m8BXp564fFoWmZ9e9S12pfqoBH79VskZ4J6FHtK20DcDQf1mUEE53qHF1m+5Zo3l
F87G+Ry2Ooa3LK1J4Lf1v2eEEhDN47dzi7Yxxt4SVe2wfHrx5KRVzRDNs5kXX67M
B+LKodh5GJKZzRU5SOb2bD6CYILRqoh8/eIeMMN135RGQE0JbdQaFuooPa/WTfWR
kwAv06v829BTy4LR6klwf+78tE8mXQO73CBKd6K9pGDpPoNlh8m4rFGDx2SOf1pQ
quSJcw9l4WohAE/C4gcDDxZRECFw/HoxLsj5FIOdBsNfitQrMGK1+2if+Hl7Py6G
UepLE9DOjWf4QUSY8YbSMEuMrqvFbb5z83jGGx3h4kc9u9ThAO+tnkJUcvF2a0s2
Mc5pTX8q4YT8pPlb9P9kzUBJe1y3isMBJnD8YZuRixFyYJDNcEzl4/yQl3HZ2Coa
ojA3L4lbA/PSadjYkBO+Et0BvfFY9IC104lilYlL8iYS0tNkOZ5s5HvyyLheEmFN
WkqVczcIoP/HbWcd313XOU9b7O7SQqgu75vNM9Z5IzClpJWqFktfGFOppkWsLl90
XPpuDZjBAQ7ibT1VUdRlVeV4v+ZKrpxx1fTpjfeGQN7LvjYD15KcoJO51IVSqoSe
rsVDgHxfHo/yfbc23AlR82C50/b0jHLLqYo6F2IPIuhnobVERGPEkQuKJu0xWkU/
50kYLtOAQiWPKPA6A9tTIBsSnciB3oh8lUy2d/lLhQlW1mKQkh8972M0KhndHR85
gzu/VNBf49gcSl7OIRwp4nBltjbwygZkJLykT2FIdBJnBwNIcKvwBgZRGPbdGEEn
kFcE31EZc8cCS2q+fC0tDld0c6Ke4xkIsJ8qb6qsDcKDLlGna0r5fnJfkWIvPFKb
TYWmU0VQhNhnszgs6zdt8IXi+Ud3Ybm8TeS0XT++6XNlab4Vbbc+JGGPFmLxQZHa
JxX2tJvkMCjsjj4EoI9jsmPFVoUQp+Srv3q/8lNlUcakjAM1Q7HbOIOxIw1xOONA
niYO2SR+AwPD5eEgVAiouHykGRb8IzW2ioYi2KDGNlV9qu8doJQpsypeY5r5uC92
vYr/fC8FeHFscg/PvaW+6CfJRoFBBcdpQKXANx+iUC3S8lxN5FkhRdwYG/DPDoug
shTmcRK1HecEgAWSvDheinBAVSy4LIiPkim08l8zXy/nktsBj+inZ8UCTGejFmWN
lPrwysFyuKT1dvpwl3jaSKFrs9FHvxO7VRWuMM3yVHoX5wocaK3xw7gEMFgvCbwa
iAXueym2WZlb26jEXxZWnl/CAItAwQmXtEL1Q9BhnVyrtte17JU7Nj58tY8PEGoi
8W0+i/BiSbitrGlqxn451hjHF2Bsmjc6vevPMXrs8VkWxhiOgB6kiH4fvhabOz7W
V4ImJG97MyNgx+n0fNfn5+msoZCvouiPGM/E+cxaO/ESHWqMdEo8RuAzvVQfpTjx
6gnpAwvlOUQYf6hJZQ9DxqgyfHw5oE6MmCojpPVCBallaGo7iMJDDKfEdDhvHnHX
9KLY540XMZWo6hWG3zafGQ+Ba/6D5y2tWy66ABAaIwhN+VBU3ZT4dSZMNTldUXyM
MNJ7FnJSI+xnGJAbKnTukJ/aqbnIpOHrtlDkdppE8PWOd+/kvIlf8kbJ2A6YDVYa
o/0XT3n6IXy44Nsq6VsZT7/ilCKaNV8DQnxehCgF4613c+KbIWyAv73afcFeu5qU
A/T/NZCGtdeUwqhlUmHi3TYEwlsk1WjOblrBlDg73ddS3m0hv0w11WLbdl1p6Ce5
AgeUDrZzynC93mBJBexLxVdrUdLUeYgXDK7Ri5zr2dQE0NkMfbIIbV8plNbv3FwU
+L3zLG8uhyLES3CkkKx2pQ/Ex0xnotodZrZFIN7Ztrtud7+ojwfxjB1CIYV3gqNV
/V7zJQTx5rBC1rJNSPOF6Rh2s5N16QYfWyQ+JAzQ+1QZK5RgG58SEj7tXNujfB14
yDVwnwYlES9lL/UX2rXNquaQlu3zOE5p8sV5imfOA1cNaG5XmEVSgQXdfpHuZoBw
WymOEUN+3xxNfdpEsDoYY1HnyP5okOfjzgMooJVpJkn2+Cguza5vdxGXZ7kld6rR
3UyeRUw7CvPxSV64dujV7uBocApkgd7yhTV6r2XnoTE/BlbLkXX6HA6rZg2JkMLA
xJ5PSWEPiGAUj6VtEMTFsvpYSz7rZK0cSDD8iSqpmTVXGAp2cmVjI8H9abVvOCen
6Aln4sXzvuETPopzlxZKLUdl+x02AUwtmoPv7EYyNi8ASsgD1p+TfPWttwPLfwDR
6xeSaN67hyKAXKAn3UowKKZRUczrhGYM89rnxscdnizrejdC3moHum6Q+8kPTsAm
9foYfyUSaAzROkm2ZjPDCokdvwb4uKRR8poreO972Uh5z17Rh28dnVpHZJ7fPhX9
/XLuRYtXms6k6hNnDSkh/nwvr3U6slunkBBKLqLRhgnKFdZwg7iSvrgzlmluURYs
z/tV4Vgb8BDyJ80zFi0qizPilISQ/UYU0CvIbtuVNPbMMsJQ/2xtEAnCLVfRMRrw
yKraUR9vDAUSwdcXzI02gD10Tp7QNvLw4x5LBw31DMogN2KA5A1lxXyBb7D2lLUA
+aJ5SIFvSfJw53mIFC2IOiIPDGJ7UfPvUkHSdLp0TS4EW8hxMaw8DzSgDBMAi1Nb
Pq+oKwl3p+OYzKowwymmFvZwc2z8HFq9MR8PngQkPk/T/iKnMMrt3XV8coBvDPi8
TyeCB40SmxQDgRHfZ5II1RXOf4Difvj4L5AUfjC61NcVu6k09XagXpIapA2g1P1X
XCLkOYUdX1FvjjfuK4vmHmfVySsuhBMkiPN9z2o2FVE7mditTYQBpRhnfScksGkd
g0gWCLPPMIRpdn2HIbTlemI34KrBsRFdijTXUB/yIrezBAt5Lz82hgovdYe/3gc7
7CV5eVmeHHymcK9lI4cuzhOSnIcQhTly3CWkgtbkfni+dpEeS6r22XGGiJQAllWr
GP/NyXqsW7jGuUmEI1+rCd3JgyOHqbgt6CbQuqFdUyeP1Z5JJwLd50h/YnGEWYJk
PSmLuhXZhw/e56ZYSOwAaj/Rp5s4cGu9LJPd8xdCtXUifT6GjOvAv0AgBJ64J+Rb
KWReqDsACRZlXj31il+8r61OIU3eV2Blpx/t851lKCPNNaRamxi7rfR3HzskTL7d
N8rHsh9rxoM9M7xirToGlDmDZR9U8yGnLUFnT7ld40GYN0kfku0Tdk1U4STx16fk
iXkZZXcVDGFRwTxDavgX6YPpcI8tNkHL6U7k0yqjhdOiVuaYSEdcJvnoHDqPTcqi
y810FxL0dRq9kFgDMNGqZVy7QKqHjDOTvE+jfyFZLhtJooKc+0wkXw/3Jj+t6KbV
JcBLJPEKww6Wh2eWGpKqNKMAIa0My20yGtJJYCQv6MUsY+kPHurOkQIoDRMpygrM
yhE91aMyxNSSLEwOpgUU92ykFmyxuWdjWtw6fSmJUarZwU9qxWuaS6Dc7DGwxz/m
UhT796f/zgXiHoadMUFyy4ucQ8HhwMyKSg5s8Rn/vL7wXhHQCYXwDo1JOU9CXW6z
RYRRP5SWUCqndPONqmkb/ImiOBRfVhVFzXbsup3ILf5NeuExF5GffHtbqsdV8Xxs
9cRpM7gI12IrSY6vIVqjNDgArGhidI19VRyCyplRxJ/9O75mgNeLYZlLFvc+9D3v
lIS5XukUBzcJQeyoBo1rzlzV9NdjGRAINJS9WyBlCXb+BGY0Xo9hJwXr1DK2Tngw
yNxbmX4EXdpzrBHmffZw9Lj3u7WvArLlCRXtCvF5rTCWvtdE/Ql9cwIvU4aGIsj9
3tiCUp7a3A7hmj4xmrlRhlXFlAoH03NFaxpCC+z8hzSI+SntRuZ4SBmXn8LpbqTz
yI64gO8Pk2CR1b46VXpSU8jT9EBgjiyu43XTcyw241G9zvOanyb3TxDuUHAO5MhX
n6SK5P0yqQH408jnawv14rdFUlBAaJKgHnwMcqPKw0E/caLnomml8WMzCbVIYG9P
yXZzqHKCftJHi3A3stBSvbKUH+9+7pWX9veyWan90JI169MSSBHYqgU0yS2eDVib
91ZyLlGEAtQwGvqzgMGh+krt7lkwV0UBnlPaFvMXidnVYkMjr45aFrNfOY5RD2WQ
E3BjMcoSo08+HDQDpfWaZ//bnaFdPq480z8qEoQb5qF/ZKe8IzcpC15SNxoMg1Cc
dYSLlfF/w1OwGw37c4jA0Tx7foZ4b8h56vU3pr+RLrywom+AzMy6wKtdVSLGXEqK
kt4RbH7a28pThQd07CFSDfFSxQ1vPxxYaDZL3z11PTmmo6VRbEeNZSVy4ePiDKfL
1agdS0idpP/Fl3QiRHqouKw3HALjn5VnLX7qfwB9OH7LBfN0I6EVhgAZJVTCq3qY
NMNSJlswyjKOgYsSXi8p1ijmgt+PZnqMfxrzSr0wWXEY2p/g7mo8S7UAhUqVl/96
6fKjIVMqaM2HPbIKyu4T3qHxG1ijXpMS4bQ0MqixMB65QtgzT6zn9Am8SouqG8fq
r2JZAJiQMtxel26RUnhV1gtw4kxgHLXfcsECfsfjBdXIwtoKXHfC4bkpgXxvbHUU
NHkoRUKyADQ91vcRfX6ycq37JfMTXQ9x5J6SRQ6PmAYI8qJPFxd//6A+nD8Aw2gc
lAyrsN8sh9tnUC9I/1SczyfGOGIHoHauYGWDselUgLU8vC2qrt+1Y8WKRDuNuNxA
/pT2cW5itkWzVHN13NPpAX+66dHpq04QQbZUlinQA2FUgYfruKE1rhvULddZEcmT
TlSHe2U1+b2fTInXvokyboJz8t46ZNn5rLwAxv2LiXmjhccfcDUv8BZWzA5sYn6c
F+PRO1i9kWQzVXA4Z+C8DFZJTxSGNVVkcuCdk8HjS4F5T5V9O+gxODD/++F+v70a
bEV+HOmbeNAmxHnMypXjqJKYUFoEmahcHpS/iNeBwMnDOzo87AN3CPLfydHCslQD
SENNjUiZprSAPcTROA+GZP4JyQObxrKsnyjDGpAK8d0MFIItTQdHLXhthffPUlFF
lYoi57MSv6hW5c24AjemmECQr2uOeh+y4Dx3XbX080/HVEYmaLwTF+lAv/vXoZdk
8EG2vzTBfStuOL0TvZ6TXB28uP+mLABoGC1A2908c1b16lFIbjngb2xlngOvbcUj
dU1yI+NX+/fsckTunoZGapABRt/eablSf/Qpv37Y3CDhDXp57U7FB81t7otzOBNx
zEu/fvjECVEI7vmlTa/IJUK/wuCWnEvYSBTrme2RZYObLED5KCjfMJJS/ChsfsfQ
iMYlxLuswNIG7JFxLPl0wxE/U4k6G5OJOFC/FBLw+s3BoqELaDcao311Gf5Qe63+
jBbEYh1vKhpKCk7rHjvS/xWdBbi0oKh8XkhbOicTJlPwqyZtRE1oictI5Mkt3Xsh
K5aykWy9K8ss0quPXoVhDiRhmujkAjaALzrpG18JmPrHvjJuWJCsqHx84Cg/09fW
tBb3UtiIzUiJs8uHPL/1/PZ1z3ao2/hhJuP62KpEy7Rlxwk0XQnapNi8/lqLOUAJ
C9wN9qjYEy0dzAl53njU6IzVc93ErBRCC29ai0Lhh+HDx5h3TAtMGcjoSQzNnVIE
psY984fXK9q3R5G2ENsddvg5uP1oaZ/gPa2gp74jRQ2OR4jRJEShogCQyZPi80yc
YF8WZz04Y9u0uzAG7MBiTrZAqhR9iTxRQJ4wAaP1Dd5/agh4HMWflILfZz60GhUY
KtzY5v9zYVvOKQ1+w8DwjM9xpG4D2CtyaMVTZa25z44sPC2Xca9z4j1ohLE+7bIB
7PpSpLPuUklQZUlEa3bNx1fpqNvyxxDQIO/3BDrWufegiIhfZ5e/pQGK7sDiqVgM
o/8qDQHQLKE0vtIAwR0wdIFmdyhkxEWsr+dnbCg7urgbb2E0yguzQJLOqupERU4m
WCn8HRLIZYj1yN9uWwQ8WdasbpF03JofJNzQSLXtfO67+VE+36fdXKkP6+CbapJu
f9YjcMC+gHaUNM07fIqlNda5QPvjK6Knx8IXpPTLUWsx17GF6tRCvIAv4nFFNXZd
oQiL0PKI6w4ymdHled6GIYnNRA5O4L002ByLD2KZh3D1SCkaS9cd4piN6TqzH4KU
UZb3IpHHInq16vSnDf0gJ5Lt60vjFg7BywD4JXsZ02uMIEQ3aUgUuqZwHtVTZ9pk
KzmPR9izydp2YaKXyZvH3E0Nd13UjFjLsN3WC5yd0eKZbQcJVr+Xngv7gSHKMZJL
X/n0uhqHJdmx4NN6tagWiqS04GLnB4bvc6HcBufnxBWS0UyBpaiOQ4R3nNf1l0Sw
3TG3HpNlEYz6HTQNUoOfmCrnq9EWpRjRjZnblhn0CiRWfhCac5le+Dymxj9DSzYG
iOUZNRnqrfWkXs9GJPR1XVFpdZlW+IvRY4D/sYSGQeaOWUtmVOam0ovxD0XRGFEG
DoRM/GBkG+4EZu52JJviaJEqsfzRMZhn/+LX3oqDHcrptkIBk0z1Q2IodBumgFu+
KMMIiqiD5PgkJaO5wkBARIogGF3cpl5h9yVe42VwDZbHA3DktnbqOvC9rMAbJCrt
wrI07JgtYjzRC63mEZ/uf5SYIIHYU7xr/e1LwdolMvzHHySAF9PrlWHfjtM6u8ax
JcWnKeAEqO7JebLP+rh3bBB/AIxuuSRjO8HqVyaQ45LGbYRWH7Y0HolKDcvZMIMV
+EuEyPBqFhkn7CE4CR8Hz7pmpKuFkLNEUWVc4Xa2nakkQFPuGfonOHd8emsR9mF8
BxoOP27CZqnGRc3vGbD4Z/rKYJqRWcJYNXfX2aSyVgVqtYsPW4KrOm77jWZlMllr
c4s1SnAtkmOq/6BKFI4RHsppHCU/ap6Hikl33PwURKwVriP1GZO4RoO/fbrhLtKI
9m34gRRvCkk7G17WcTDGXct7bli0HgdCLGln+E6CyMjuOD81lsxfcGuXKobFZgXL
pv/RAz9Q/3qQFgM6SJ4iSst+r0uZm9Qq20+M5e8KT811CQJZFL6BD/c8XyNKZ2JF
nJULQn9LQZ0bg8ZS7MKoABkISdOzpfNd8LMbzL78TveW034LMUWWV4fLoL5lnH+d
q1uCNlbWYlw0tVlHf5sIwXPQ+MUUH+Y8U0u+H87l4eU+05ADu+GVUORMEVbV5gbc
+WSNmwV5hSC9fseB5qKUwLwpU3BBcZJqwAPacf9/2DMfRNElN9VxULk+BC98HlNX
WS8A+k6oSSj6bskADx2vH6T5xXR8moQI9T8h7Lieycon76laRmQQNfnkA8QPf86V
6EOFpV+3xKc+DS+2tyUEYSUN1qLLclV+VC2onC09kdcfdaKLl+UdxOf317Dyw4lN
DUVKMOgmuqC4GcCikPMM+aCXJFXs/i9k9ClvxNGxrBeIu2UVJDMoo/LaSHGZoxGP
0hnOb/UZR1xW2cI44QIOUM+Us/J8UEnAadLaTVDqHBaouc3M30vGlsXyMeNVoCLa
w2+R2nnkryIojmYlY9cRDU4LbNT8h2O8RlCkzSdncYsVAZ6VdcbrBg0PDAn8b6dC
aAU2WsvueuFF4aO2Q7GqsWLqQvYAptEIzmAXOq7+hS+axpGp1naQ+BjnSagTPF1s
vpgsqiBDSk2U/fwtmoVjCMeDx62F7h1J+3y5gP1ITafySJvcVU3phfDjaS2nhbBR
9VIIufZGg0YVcqqF4KAdskWr3hpXZDojnhYENRFag03YGfOSJxw3IbrMnWV0b1tl
BlDe7+l2CD33RRkWDeXHrf5y7sDcwwskA25NUQOsF9i8zU0cVV8hqRAUnxQTrRgO
mUYA+gwx1Zdv2KPfbAxq4BhuNAxmfpSyDnDeDAYG47c/xYbYzDE3EHkriEB/a+sQ
RY/BqgLUUheigAvs5j6ekomOWAENrpJctZXK4KvCHdPAA7hF77gj4T0Gh7V/aTlr
h/BVOM9pAyCc1eNmG18qitI+tlgFggnivwm/gnIaz+9RwdpqeiUkjiHGAA/yZsOx
vhN2M10HGtieayYaZdqNSPt8d7NxoKGuBvN/uFkOta8IBaBDEtm9evrsJOMWagVE
cBm3hOzBOBwA2rdrPgwwE9AwLy7enEFc0F/Uh9rTMHRS20OEFiEKwPNCSuO3ghRd
9FaXQzFOEczob/AqDWnFYVm96Xseh0pdEnPFxoQWK8q9eTLe+pL74GqTy8iiH1H9
KUPMctqZ4b4hlrFw5My6Eo0nS3n4TmH9dsyypIFuYeKPNs/TulZEdGWCgXGLL9Xi
A8I0aioLxk3pYQloirPmTdPVh8sZui2S8T+Ze77YztXq9LvoxNYs0zCIR+H0/Krj
NJVSeK3PGJMQtToGsvPbahttHNU6v6OrKMCBBbBwJE6A1r+smvQ0RsFYG0OXOE7Q
X7d6hc41VPY3sbEJSM+n+Ci9sp58tFlmVhvTY5dyg0L3FtUgzI53xlThF9v8fTTB
S58wjoaOfJ2BijebcwuqH6leAiRzrshKzaUkRhOU8X/vcfDusoEaEbAbaEpLSvBT
fuBVgX9bcY846haJZOeroJsmcJuq+ieLcgeHSeYzdS42jP01Esxc5oLPzE7tw/q5
+g9Gs1zC5vtMFkwEmG2vvx6XPIcBCDAXjCrU7OM1r9vBtFmAe4RvqUdgRSKCKgI9
YLa3g4MZtYTls4N1Uvt+Usue8oAxnQWj69gri09tRSo0oVrU0gFmYc4yoINI2Mb6
yLRNRyI/YEM8eAdFr9j6wMjS5fJxVCOH3fKfbvT4qadVuvEoDjPSbpXOexKR/ooR
KHzxe5n7/p5f5hO0+kx5kCm+RosXfmEHpwSw5NZNS/a6gzoBkY0UgaD+uwDmYMmy
j9io8MQFyKmF8k292FkLTq4X6yY4P3yv6+aVW463m+LnRF/Lo4bycga8HtHEENuB
fUFLLURcfIDa8gZRD4tn3BRgbbzOaFKk9WvRDSSRYaLFp4yNLdK8llSX7G2izXp3
BU79++E5K4b63KgsGuqk/sZP+c/iURwcEUzSwYBwF1TFatXtMCzMuQ9IorUDsLLV
M32NXC51MhynSCMjA0rsxULLyiZ/iSu3C2xqs0Q8LFX9Iz22/Eagw+IiTPExlSfg
3vtL3P0Uu/L6lceZWYnI7D/txTnvbelzLnhYDEuTFaHkrPtR9pL2oCIxH+zHkjo3
xLAYb6zmg82vL0lcaT58ycRmoULr3BDBQ5DZsrfl5rgJqU+3LgfH1LsGokPJf+ma
59A3RkdhlMGvpk0/ezJk1wHUoGv/M6ddmce0LCxeDEoZxUJMuBhGMXklvdvzcSXl
T9XbeSXsO/VEKPFyZZg2uxn2e7+HmYF/8SBvZjdQDu0FT1GGv8mnVJYmuDHdymWq
8C9uczxDGwisZBQlA/eydmcV3P7khFjmDGQM8BYL/nrvLwzUYQGjRcs5SMSU8nMM
NosVL/Fe0EDEJYyfbC/XXjV+7CqYE86vqk+9AyCpKX1ehPrGUw84dLV1yPZH0/Dm
R/MnNxTxrCRMld5XRCdDkcRaAnRsF2P2GZ5R4gtRaQXs6i5jtVx5mp+3n/k8JfRV
PO6QOBCP/nd9nzegfNXkGmSiYQfpUZ9//s2WRmvwo6aHziPwh3IPUo5dJY2a9s8h
EEoI/zCZpxcdYjLnsk9DzubGXlBvrRfgxV4MjvG5rUrOwMBxdZmIpxZDVHxK8uBF
fhzUkMZR9tu3Hr289MBYSxVe7Zwo8afpoqVBuxUj0UC/xRLpEqd1YF2nOZcVjZmc
0xtBXLhBKr9e/6Rl/8dj8xla0ptwlSPeI3zuNY/6I9NYyOFK7PItRm3fQlOHVmkv
T3IxABZr2LQMRk4tieq8R6kBYXdWVL/GmQFAUPn72TfXQ0j1rQzsUQdxbebC2fB0
nBmHTE4KF9X9biLdy92I1vWlJZmUGVK/Twi9Kb0Z2WIGVwZicWlNyEANEw1C+NhK
w9ydNGcM9SQtfpApEaOigSFUw5r5paoNXiBo4W+SLWd0PzdCYhtXwwoWBin35Mtf
EAONhTvkUTwF1nyAA98Tj0ClAn9sdihDdBhkqm4eRRcCVjUBxa64XgB67/4qeCqK
D4WQegQ73QMOR6Sngb5sMCVy7OoXvXdJJGjokR//H/zvTwCg0khKTYFtgwg1Mvy1
O2lNgwh/9LBM06C8anmIXNFQmW2bwMC5DiEvYDAjkggLowbOwgaYOAQJoSctK2rQ
rbEpQEmzEc+BZ6AUJpFqQxBR95yT3y0jCjmH2cVjPT92Kr9mgkFK7FIHXvtSBrs4
bZDimxcgWYYECABzdKET4JzHIvXoUXmvi9c9WUiMnJgOp3EFx2pjF4Ipb3Bb25TQ
8euzqcHg8otmsGDXRXKj7SiHbZ4rjeHHKuYPO6tqmZ2samQa2eGfDo9bdMd6rNOH
QQdl/vyvrUwcNJMklHIeXVjycw948kGGHGEQ0gHLJxtPyZH9GmiWEGTFUy0CDnSD
drkize1ud8WKTp4dr0n3whTJjc0mwhVXWzC1X5HgP8TaZkntRNDe20fVx2KNHiU1
7bFE7t02WRDVpPs65yIooIYr/72GVQyABuHMc+koQUhIwI8jnKy15D/X6dn9lCuk
wNAnTJXvmc1UQeQKo3qiWYyZvWEBKAEmlCMX0iM1/4ztAh9D753YZF8bej2zzKGM
ZIFMLRedf3erx4EueHvC4romh0wOf6NaIPTF88zFWhynJvQw2QaqFZ3opCdCVuYk
YQxL1hIdbVmBkXlpfirifqiGhWPZztfVHkApDfvEcWXczBnI1L46x44C1lHm36mY
SE0t7RzlOMuJVhuP+tM7RMDVp4z0RYSQjOiwwXM1R6p5P/Jr0Tme1ePM8NXy8gkv
f9Yuhf589DHIGD6x3RaotxIALrAgzFyKf/qcEPSJ6GMdYKaL5qey9gyjut4Yr8eX
UfaWgv5OJLP6Dq0QNdxBmWR8+pvi8qgjz7C7FPodyWufkTT1pGN83BN/nFTURhf0
23rYj9mRE5sCt7BSp0PP9v9cI5ij3gZOpxZY+dYhzb5eHQ6SBp0OBvqPtaQEtTaJ
hkBjgo4/K+CLSrgprIbrEKe8FyNt6RtB86a0O3Wm7yuLmwsypy6z8PlQ40sYsL6h
LMPS7IS+8VMuydquCOoAoSSNdFYkb5z1+gRxceiKb9FTl0QOai+mQn1hJiBb96M8
TU5ww8QZDc97+NyXRB0ic/0I9Q4wVMTQQNRaNIE4Rnufb7VMPTebeaVnP0SNLhb4
JKQ8cgXaFl94SZLjXZQ5a5TduqONymbX8aYrtsEFYwmE3jMGGWR5iEjHTajT87aM
ILVPNEopNpl8kRZlMg/jUFYXpJSPZT0utnCSUTJ2Cui6nFPJNCzZ6+X3qCm9ldiO
2ToekidUsljLZG1tDcWAx2aPHnT3yl8HZ4Fc263b6hvYsLmgKJJYAljXVqmCUlEp
8qHG/ZoBzMwWzUn8D86q8ifIbat+lpIsY0MqfOe646GqZ8oIzIcTLZA34Fx5beSP
Yfi4Guqh1ywiqNrheEx2ptcjmapnI48WLD6OjtdfuSYf/w4diK2g6rBjOWOvO3re
cL0ZimNkwXpnajYF5lwWbpUd4bQMqcbjtUoI/LZpe9DxIiB9XfT+Ps6zpmOW1lWN
IjRfVSgRPBXwb+UySJbhHzqm3WoUy5WwkTIZHISwth8isUyVtR0N+dJxV3eBYBxh
D787Qxiv0z7LATOqIehqAOyGpm+P3tuMywCrxXVmMXpoX+/eMXJRBbjUf30Vctvk
T1nr2GWJxp76Sd6keq34BtTB38Rti73BouxjL42V8NkpDx45gN4K+d9ehEnGyivx
K09VptPv+fuO2Jc6hc6Pk4xuVQBSKsBvvrE/wsv3yfljgE8b8M/LlW4/kjWRU0SY
msqb75HDdJkP1CUzAapUp2eetuPyYcPzq2Nj8xHSly+jwZO0ZGKmY/04OrZ/Nz6I
QguT+tr/oX1HnuTrVxXYoeZB9L7qcgdeoTEcz6pKsqD4+YWTaclHwhd3kQmkh8/g
g4UQ5Dz29JEAkTnKyjewATBOsVttb3oKmckEtwoeRa1Qisv1RrNJ0K8Z5QKsCTDs
pkeMV/omZAyoQ2f9mCFHkXH4SOXZIkN9lV52mKDDZmUzIXKj7eurv3fuMcT3YA6D
C0oUHXpEJSJosbpyRT9pwIwjZIaYlMXi+vRvstFBoWVGEvUpgPh15fWNsvda8BPY
yvpU8mO/m5ZyLvfa/20mg9JShFO8/ogKHCHI0XOCGosTNzsrIT8VytytNLMA0WMu
HZCWIyiYkOgKHV10yvpoA3vqYi/vtOFeiT8IiKSZ1sfFB3XR07C8q7fkARBWkRG7
nmvaICyAAHv/AIbXyDbdqIizWZ+t9tnRC52UIfpVM84/0jN0iys1Ztcf/42FsSlG
Wh1NmxmvPNiwjYin3Jja7Or6xPTWFh4gM6LGCx7y6HT9elxVhQ+D5jNfbxanaPpK
6z+6Tr52MZoCXzrttdMT16SFi49ent8xUJZjlxcHML6+KA1MQhQOgXkinmS+TgMF
rhTjeFDPYxC+CVOhw1QEmw+MrqWsQ9KDuaccMGDhhWkUV9LWtLbl3ULEm+Ga2ybV
Y/zAI2+bO0vu+iQ1WlhbqZ6aNGr7GlUx0dRnOzlilVArAaNGT1KKJbwA3YYTag4N
RuQyixBAOFTlnqHF7KFbURL8QV0ModCGXlNzRTiqxQCbFzIB+OhDVn6YWggvyP8V
xikJ0JiSbF927ywD+yfuCINdzOiF4ouc8fP05yemVvJ3xJN88GdBDG6nAlnZMXYz
N9uep1rzXB+a/gJDlFMbJ1Go23TlbqolZKw5vzX2ATlSu6HtuDD/KkA8BdL73Fjb
OqjRh7UZn5/JW3FW5t6DtwjYynEgKwoFL2XkWj5pbgExSkoLQxFUPvA2ftl1rYMv
HrOQRX1JwXY487f0QoNON8A7S81qHGw0XDZnLXssSG5eF5irq6+iDWdSOK9CttFU
Ww3XP1Kvb6n2Ll6NjRKkCJEnXsLDTMu4rX5asIgl+Gf/mTG/isgCH6Un4ToNoDUC
tE8jP+0qzboo6GS7GjnUVC1emEuiBKm33NlwotvWdSDFmHIEIRo+L2oqSvTRWL4U
pFSP8Leqx9XKGEvNm/heC0LUBHzBKMtmfJTcqD7sENgsfoaoOzVOo0PPQBhgIjSe
wtMW33ccjiJQvLC7RxQPOHC5oa7tFfbPJRw9dIqGFiTq0wCh+Lcvqk7DL/0g7TSA
dPO9v5LA6Ge8HgcE6HN6mk32r4QzOZTkABrGAlGl6EE80IpqY0ONRajDu0ryCLJS
3B5SHmHHs9+T83J6glA4IdhdVfHfV5J1ngzCoLt0UfEhKYatyCePr05/yNatwpYp
5zXuKe02pKjmZMSVw9sMp1sVeTHwHpP2GvFQifyusTC3sIjlxcSaMt2BuUxA/er/
ERZzAjLBp56ea068tsjwaPNo7ijg/ej8Sf/ZorAOuu4TsbcoP3pVk6Q6q75C5b27
sO6FAolfV/vebY4ah3QmBWexOhIn9Z1SnabTGa9oP778YxHQLN96eJPXHh07J2ao
4OOPNEN2sup22rdcYplxdRqzRJ7vAjplOcKFoCjfhUpKRYCa8W5N7+Dy3gESngDg
HqrEWtKT+/EmBZP0HJxtE+2EcLMIhI0uC3/slWUcrU8s7dXokoEiFltjae1vqT5l
5defkgqyKjE0k+q5kKLwtqqXy7HYPrUVU80lOMcAIBE+KeZL1wYGqucitSM8zkrL
C7HUFa5S6HV/BV983H9617f5K4rcxasayWoJvs4QEwx7br3Ne+niFFhOYQFU+1vv
PUgEU/hhAt94jXvStzYjchA6hX15vII0hlF95IWnKqk8qnAJiOjKHJQhSeHCilM7
tZNByMK+VkwMsgDehlL+Y9beLKWDaIKuXbIgYOzW9Nu1hbqyl7rO43uaTQnLJu3q
rhx0txGLod9VBbB1xSBtyHN1ANXyt9QgGFFI/mj+Hjp0fw5xXA+OI0gQwFKzQUnJ
eWtz+l7bhZ+K6YWb48PWNM2yTpTNfM5dExhzDD/rb7Mt00Dpea06vAKzFMIMnnNA
VhJE7UBoRgtZLWbg+gHkXklo6O90XFk42YvCFxAXxZRoALkK1uZkdHO3/qup2NWH
HC6bc02LZQqD0UKvXqXsM51032i8twuqZb641WvxpvoTzYtTk/XukLIdOZkGOmDb
G5pjThbsofou9+uEmZSc7+rqEkosq9sG3xkw+uZ604s2cXDSigRY8hynlFGV7rYX
T/ZdfSscoHbTFdhK/2spc/xAq1cCx/0Wui607yWfBLsX5Uj3LxecQZOfvOU2DHe+
f3+lYK2xRYcaT2j5Bf1BC+Do0jALc9IshSpCU17uOtjRR6gCMrbC13VdUxaIcNhA
w86KNelzjXRzTK0eYR9yfQ25OWFsNGcbupiWOMdpjwOj23WzPebdNAd2BQNg6bke
bf/TSmCivSFe3QW+a7nzSohCfWjf/SqcUVK2oQwwdHmmVBa88BhSu3oTbGCWCx8E
UHuUew6CW7YlUvxdkBgpO/XVjB7DRHKcHkY6sSqm5rgQTCzc5UpVd3jnHcWQAJGv
JA9ZTqx1cbbPjoS4B6fKh3D0ynQlYAxLF8zKpOSllLWX6+coyDsFoTMd5xg5uKKu
yUnWpBgKP7dH2gGUj2TtkyPO0mxvsYye6s3cnkLQjLpOpwNl0m7Ujsn4sA9WCFEt
OmFxcciH2isBS8AzH8T140sVQoWJSjeWj96WaKGbNnVC5rCOtSP3slvGqfnNr6NA
vYiihSRIS0KnGZyUnBk/F5YUFDDPzJM/ZlpK2w9c8BZCPVC0377le3E1NgYLqA5N
qwGknQzz4zlKee+jDZdMz7OVFbK902FQZFp22ShdlJf7fmGmsVcGbCIfLyxfrIU+
pWGvq5xIz9D8O18A3TMZJ+rNZQ5OVK3jUg2KepjSb1bqZ6g+gIvbMLm2FeHAph+b
HQZvWZauyz3PxqNKMq3ciQD2o6j4pj4C2ikDWkns/rBdUQquW4nKINBr4XnQWzBB
tHm+j7tUyF+Uz8kp748u5K+fPIlXOZ1aciq1oJQ+GtC5IjM5Mkw3IpYAoa8xg/e7
yz2Sv57P6puCtLa9VP4z5L9IQh4NR6VGl1qpEa+WiVhjgr9Nwf1YDTmY/KNGEbdy
Tfww4yzQBGYvkoIODM9BkTVE0EsoyzwpfWRmCf2BW2L/WoQQ78fTIJl5bdSREZ1w
P47X1e18gWMJUj5sWCUonQgw+/5yoboKQ3jpV2NfKNjFGmguvdO3comaxmYBJNr6
amygbTJU/7MLSEm0sn6Nq1kGEpK1IULNBzi37LVFZukGuV7Zw1yKNzgMxRkRjY5/
Y8GQ2aP4spSgW4nEvctSifho2uNB+375kPk1FXZb/4/HOZWshDeW2VFO+3Hm1h+R
AxY9m2hSXmXy3mlabvLjAo1H+c8Iu6tbwlZmxAlV+KBC41Wo4jU3S51rBfo9HsKw
hft8MoNa7GjX5pX0h6qx9FggMtz4iQcy19J8j6DxchvJCgdye/tBa/uQR+4Ud0L4
yPacD74BGtGY7G2GlegO+LxC3fQdTNXEDZ/eAsOOOk8JIoWRZx/9z0F8e1r2/Ekp
Pc+j+rc+HXQXICuqPMk62E0B3+gBCDCyMB9/QT7hwlIGDM/hsGI9E6ZjbMV0N2Ew
sMNCs3a0swWbZGzDLdtj1MqKcP6f51x+iDODeSI+R34xX27vcTNL1rXXlCrkRYW8
aogpwisROd2+Cq0wo46SzEiaRyviy7sk5avKdkRMXefpnBlSD5MlcuGGckUuYaPr
UTsU4SvPxkqX9nsvDr+m/q+SMal5FLpyY4HiK1dnOlpTq0dNKVNu+id2NAI9TPGZ
zQfuAhUtcjE+UIRmsXoAgyLr9xcUN07gMa/piTi9OB/SDgacecxZaAnwR6U2OYO0
RLwAeoOLcOtOPilUe7vJzZqbGmZehUPdCNHkCVkIx3CSKnZLBLYW2JAXGJnYdIJq
j9muM7aBfr6EwGFbj/M/9l9i9SQsj8EwA9dcpqv98Suf2h2G1I6LXDrNPFOlARQN
9J+ni71NN1SIqWKIOrqCGsao8LdgvwcyDw0/FQ9xXTAc8VVN+4oSbqYpnx+LF3Zc
jBelCzDwhu/hlfxk1/OJv5zMa72Rtp/ycvGJmgVt1MG7AlAd2dB8avr8CsZiubsl
1EYEzceB2Fqnuzk+jyUwF94nYIZ+7e1ut89FOzvbrlAXwAbU3RieqmS3+m5a0Wn8
RzYLRtYcQMugD5YHEdS88ZhHIWwQQlg4Y0Tr7m4OMSyuAlMRX07SSB7KSFpIuU8O
PLOCOqmAc7I8l84JNMXLh00fJkf3zsQs1eGsBrpYmWc3hBu6KYFbiY0ktB9eam35
GSZi+Fj2LJnbTtWuVp8gKfdQgnX1wJNhF4eBRwUAKOv7sGVPSKc0gABjI1Cwh5N7
QPdtX95bOjyiWwlVxm57QifOKK0WI/zkwvfukPkGsPbbLHps5ffpobBPFipd2EXf
OjGYboorMyPiM6zPiHfm1t8aaUz7s2LfURNBlBNL8fPVMlb0MiueBAwprL3Mb9Ar
0TiKVBjcxXsjPG8ArZFI5yJgTrAGL/oLRgmwr/1KfSyyXe/4fZoIqw/LjZhZC7G5
dh/mWnomDWn+SQ1UcK3n1ufKtJ646eyOsdQs5js6bv/tu2YNJxeIwj7h1U0kP2NZ
SqG0O1Lh/0moKWkKbV4cNEAwHwkruz9se8SFMpdKNibvBw6HjprbOqpJgXvgFqri
W70TR9N+tkLSBGUUoyW09jb1HI81b1Wc91aT9vkTv4cG5ZW5We9SbNUAf+b/VyNW
fHtiA2gLsEFKzPYpzGGQVe3NaCDrpcQQ14hN64HesjlUtq4Dby+61hfHq32MHdTw
kv7TneL5z1eieZhbXBGo/OnPstvkhnjMf++iXg+p447rtuoqcl5fD8KAmwlvoqW1
EeVoOqel5AAGHsNhDgIbWL3KSt+gfNwfmeKjaTnV771dacNiySMikg1y4fdWi9DC
9oDnNmgCpLNJP2hBZkYCUoK21ZzG+plVjp6whH4JclVlkzjIffjdbu4tegOUnFwq
53IccEkmtbYK1Zdu4W3NsHqqJMT72sHVhlcOQKU6/4/280OCxyTIKdDKGteVcEdF
XZAN9z4X/yPI7vWZkclQRlVOMHqXyBflz1qhCwSw5mwXwnwzt5QBkHPAuP3v9NcW
cU+nibf6Jw16BqBo2lxYjh+EiKYBtYEaXL6cmCte6eI2/F8j0zo7YVEGD7Y/l/Qb
OcJ1fWvWlpekVAr4825gVFcjhccvxD16HFx9LauafmiNjwlPPzOj1guSl8uKHDyb
gbQb6bd8LCYWRkJqtgz/f4HcCg3LPH3lm42rBMwlG7p62gtcJle+LXt0GKLbOJGz
2Im5vNpx1DaoqQTsAFPDN75YXgLJokBNoQSo+mRuUVaYeI/UMPMpjDKCOYe83gA8
r32S51YFMrYg2fXAfJ++Swg53cAX+PjNU/bw9pNRhOPEYT6HJvp7mcbyUJSBG7xj
1+YNMZ65XZaTdigaNRlAM1+fD4u1/DXZe/2LlfiVzZYd02xyjstL7cSpHsJupERA
F4oUbtFS6D2Jo1oCQ6xbyLOEvwZmqbT6IimNxIu6VLL9b8QsP+FDns5EHttCRGxC
2iv2J9IzE+EyQBGb4L7JTBuoTm22iwSZGl7hb/JctAsKfxyFlQnaSD2L6fLDHKZb
W1c/rzQrDQ3NxhrAo4s0VTWWk8AbjFl1xp3YCGIEfxpdpZ3pKfUKEHFssHwKUgSc
DyP8TfU2m0BFh7TA1UlOO2BT1DpYQZlRp+WXTz+iwJ/eflIOv+g2/qGgQGA8FPZ4
+7swByAAxTQ78y1jSG6jfM+4D1LKi5G7JGEdIQ45RUZFrTNUYw8j9LWaCCqNTwXA
88X/COr8sscjgjP2I2CHFMiVl8/erxmxyHye0MKw9tmRnnoWr0wcUy08qADyjWqV
dnCUmrMLwQCSqodqUXBP7IqMvk+CLqrfKspuXjrM1yX62KJne5P4gr6Tr/47LcQ9
4SL/5ffTwyEgl2bXg+8rNhgr+olclms/Hc8c1uPUF5yE370aVTx/yjp5J4QUzW6x
CHNOTEmSIm5vPbygRYw+Qj96ID9VzbRrW8AcYu/6of0G4KwGJq+IIE5NMbHmMSr3
3KdCgfXGXr1sI6KMVFkn7d/YonIosXiIODTXC0uYOZH//kPvIsByl5MwGJnOIy+U
nhJc56T2SQzcKg31Q4SAgnny9GytLV0qkcl21I2iiTODdN8qJtSkEmlD3IpAPmvG
i2Nol9cEVP9q91l/9V/PNAAPVETJ9TDzLU9b45wKUib1fs/1BAJ0znUa5zyrcpA6
QQnRDviDiPQMZYHqOXHN44pv76n1C/3sZLwkRAG+ihdsZlIp4cWQoIxn5ILcgHos
X1RdTe89lIPxsuj2cfc9/FgvT/qOjGPeHGjbdLg9gcjssZQP6jdleyU+YNoplZD5
box3YlSO3d9eMpnv4fQPHI+Odc9nj5ba1HrDtZuc/TINs34m3pjcPKqShAAipG7R
EFRKMB+LgimHLMdlO9HgRABO9S4nsTe8tKh962ehr+LrTmNYGsGSKKBp8A5v/qs7
HWe/axX5UZOAO4EsCLlK/YKWhbR2D9Drp9Uw89rtNn3oZ2H3mkk4lELsLxG/g2p6
rVO3FNABHZBDbjITS0wJqgtIfjRx7L4er9i9NuzSxgQe7E34laJ1IQmV+A+SOlZA
pQ07HcQEOSUhzMNBcsRa1JkAOkxlLTFDaMdHRfVUmMVEqLpUUjjgRy1BfHXt0v/p
hQ51qtFgephpmCEWzPZHyLHNztjiU5uP/clFCYQZ3BNSas8YA9GpcmHuFFfOfllr
5Jx1FAEjn490Q5G6Vv0giSLo9W/oHcj8H5D7XVx+X+d2SBDlsaN7av7shuogDOI8
uDJHCB/kufT6jw8eD/AwQciQaS+KF+/pDS3GBqU9xz96tv/u0M21WRAfDdmqo/ej
CMhrKXIUbnkRMgyNDhqvZmy2OEVI4RabRLh0WrnqUmh966nAmypV/FscjT16JStf
qxSM/0jtTVrmKzdt0Q0ouM4tJFevbVhLWiy4Xs2d6i6OGUAZ1FrQoJyc32GKNQKG
Y1kKRvThj40/2xeSKn/XCs9fDnPEMCBmS37m4nSGnb2ALsdu/bDpm1nbjr64UpeU
Huw7JTt7zkvdBv6y/BDU9cQZ+voHZqR7Q+v3I3+qr+2p79QzdBBDO7/DB+8V+9ka
jXXrQ/LiRljdmvwxS60hx+jScfzb2ySQO5YEd+I4KxUcZnUS8DvVv7JP1mp8ql3l
BpUhE+l7v6/YiZEVtVplDD8kpeNiNOT8otEoOm4PI+ckKge/rDUZCU2XIP3h9kFy
Iw55p65UffBGgqMxGc/NsUTiYug1AoUyUgorP3XVsX8F7D8bKTNPZENmm5gp0hGc
g06wnwV9wGAstCvJ/s0QQVm/BFV+yPnF5Ap1FQBlRAZ4OW9VM9ax0RxVrmeKvT7i
mvguaNeCOfkqQ2H6CScZyuUVMxlxq1Dup8cNx1gkKgWh0d0ULuwiQta+1gt05hTI
33thrgKtN+x6BW7YkrttE0DvijwqTHLyi+OiR7hpc/Ml141U1WnCxKDs5UYQa+1w
uXViRm8+YD3US0jcEFur1iQ6rul1NtG0Yrm10GM1I/jdQH+79SZvtSFvwb5R55/C
ShoN0fMQMHbxGtBdjv2Wdw1lkXuXD/8qLsnQgq+M3EChC7GXK/jCFzz8xxVsritJ
pTM8fBLbGEORmP3b5sXeJPuEEtT/aBAIruhKKTZOidLnT0ojZnxZpxA972yR5tUc
6Ouj1SPDoyR17i1NfTaFqvG0mBUbt2cgT7oKwGL5UYcuJJrLf6V7r7yKbBPdB1fW
0JvMth/jsjBvb5phmlt3MgnZYWDHM+GNTlOcIZvZk+GF/cahwNDHoBdtmAgWFmuJ
bJsLTEflb1Ya6KhYcNCxYk9AvIDFBzWq2l3+YTXv5ZUfFgHGK3bxPv4aYCt3SOqr
YPYSc4aQGBTWWEUzdlX47XXHdov/EtRCMY/JYboXKuQtNPbGQ/sSDPfpT0L8JrEC
cIEIIfA/MZtoc+HB8EVLU7B2W8AYP1QTqnnXxHj0LKQEHvMVw2xP1KT5VjpUqFxt
77rNlHmnps35lAB3xtElthbxu+/9oZIDW0OCXFWQe9QYLOPg3ScQ28Q/2intJDk6
8CUHwO1tiYHmyH0BQ6WBcHOq6BQJCmZA79QHNkQimHCHNe4GV4g/L+JksiNmt6pe
0jZ/Bb2h7uVBGgooKvEXTbPhdz1oEKXJR/pSkTK1vQDvP//lVtpyQ0gI9p82Cufg
nkhKTc/czRSQN6b9edWJdtTZV5QZzlClpy1VJ0fH9rN+P1FJdSCAsaTlgY7hbdvn
nztPJdGrv1ROevXRzNpG4dXzt0jYrZh8ycgq5dIYvlDyz+DzF6KvIagWTrKyJWuB
YRdt7IhNTU9hQbHkXV6Nufp/gDbBaXjPyQqkPcxLB+rO0++v3B3yIf5+L/lPVAnd
zIR/hVrrQ5yOUdN+8LPDt6gMjVLo5ggr190wi7fiSqr2sbudCB0LQ9FXgriw6Gzk
Oc0iXiW8/MzUG1AgZXQxrXKvUm7G/pb85a23D9lBp1piOa2iEU3W63bOvg+3rHC/
7HTrcWQmOhm0UhIQ9FAqTD/kX38hwIGEVY/UJCcD+x95kuWX9n+E0LfzcdA1RC6P
UI+LLaUPupdLZ+M5Fy0TZWc/KwHV1lxSSyLug6JseCPaES12z4MW8r88UVXog0Qz
BnTKXFCGAWP8gCG8Y/LVlzi0HMcIEz8RNakzpV4BW31Ji0Fi6a1CjS4BRI4kI/br
m+GdMP4AcS7rVTDI4ai6G7L/k51FAGAFnvqFCgd4AsJNyHetzt9tXwF5kjBKn3ff
+l1XuaVed224Cbc4UE1xwgw1wYz5AFITMwKa4Aq5Z6r7+chKD3MLeuRLfenbAcpz
cvSGZA7QLLsZk+/rETKngGbH8eKbqWMW4Eg8hXqP8iphIo9O48l1SN/nYW24UjdQ
ht2DxizMUauvWF/WCdfVMD8jT3B5IkuHgz7ytLhvnnwPsz69Wcdigh5HEmK0LBwH
085b/2SNeqexoIa4roblVjU0S/LTYfGS+3eQYVII0OkOrx0RVovGNYZOZRO0mfYh
EMDLFC4vGqvWuEgbohv7jNF3Juf2mNFZfd6vamPXk+HpAJuRaEFZaEz5YNn+e2bZ
pPuJRs6Tg5fPJ3K3ujOnEUAfy1E2siaw0Pp71dpMd1khd78hr4Is8uWm2c+4+xy/
K/Lr2lpzh6MgLbjymoU4FAkaLA4XzAP6UQnKPGfg5d9n4asN/yfuYO1sfNIMfx/M
J0HQxqUgwSU3di15nj4X6gvDA6kxv7QFQCYSl2fziJINybdwPTkL7MsIuoX3PWZx
jgtRDE0moQsfR3IXj7FAnT8fOa9hS2F7Ten44FAlGi39U2+HV/qoA6vdW44eBvpA
i4wJJb7WiIYGZnY7NP5SOFmM5al2pK2uHrcEMiHlxBxNhrNubMZ51acM6rWbyr3d
Rm4lyIpcUUgiWzvhx1F4J1iRa6K9HDLnwUdCe916E1utIkbueDC3ZP3wO7hRBCPE
yqO2pVcBOgGEzPvG4oC37GYSJ/0+u7Fy7y0PRpQ71tgWP4vrmX0Frco4Y3Thbx8e
/AGo0ahN7DSmUv+B3z/uNIavYVny3yTykesD5uU25+Wof8NNEeGl65/qaP4r5Mo9
RMEXQVyJJrah9ZitnJ9JMf2j9vWBeDRKHT49tGgvHUsNsjPyED8eO6z09cTAly+M
LA/PgBvA0Qs49KZMnvlQS06W2iFGSu1j9O4VD6QZnW/7D1JcyjUtYgmLPMqaIVtV
lQF2zS2BLcyY4PMS9EV868QKKFh7XTpfj0eHSWm5aEFHiBMoe/uLf1qpQDNQjTT9
84SGfOvGKiKpAjNKBuOFODQUGpv8Kb/QkLY0MbfUcNDArrb7WNciZnanpClWu5ku
O7+qbgfidv2Ui1VOcOSfxwmloImkILK3L65dSa7dvfvg34QSkuOyFvgvTdjgbhin
XqsFxXSsFwkNKFq8jXLMUIBWZZGtioV1WOmsLzqKj7Jbb1u5d4LPF9pVXnWXPPKJ
LmatE2FHh4SwZuYiBOJ0MmIrvmVniQpeqgHta5LHSRcTPSEGoby/uOW25H4cBjym
Duxz7VUJD8p+RULPpua05u7OdEsjxa3Qc6GNp0wBeGQG07pzg/YPZDouu4GDKUJG
OvYcTJo4O7ZKQryaCaQagwZ863Kdx+xGCoP5CP4SqnGk40ejdmgg2pXx/8vYpf+9
pUla9lby07qAir52u2lkIMdaC8yo8TySsHXRyabHYxeDXpt5ExQQKH40X6+uInwJ
BZ9nk4fPW56uSxMaK4x8kqGrTxOy9jzS9Xpj0DTs5f/eovkmvocfxZKiGYIu7Z/p
BR7D1Aye3fADBb3CDkA3uNktLh9y+VkuE5oK5u70gNMpW1BjIGxENoiaOl6KYYwL
80b7xAZiMOOX/MWoIvjHxwOrXAsMLEjmWZ2s2CRXcQ+KBssO6F+EQ9FdnoV8ogQI
GxVcYT4ShjOzz7aYAw/g0xkHQlSWuvOgwk29wOeCBlgWLbby+akQlSKjR9aA5vTB
khThoYEPa4UFf0UwK8Dke3w8VDgpufXU/JGgsIda1QBR67rasWSUFz6SdiMo4ThM
WKK8nzaPwuVEFRQNLSgqgISkITi32i62MlgRuF6Mkj6GJpjpzcX0D8zK3zZ6xPOa
YcvKuUxGexfYh1oTX3bAf0LUoiD9R2RadBqJ+0KAc1dqRxQ3DLpPFhj/nolpE4br
Zxdz8H+IzwOY/FMHYrolbwn6BBaA/tgCnzMdWHxAJK9FywQHG4l+eh+hAUEEnvDb
tlwcDzgfs/0nbnc6PSJrdgNWRdCUVDOEy14D3Ix4chnIcQLmlrkweR4t947mUNE+
xNay6QuDAF2SwdxolmhxUFgfyfRa6aAqg0bHnh69rLnrG4U8DLH+q9qsf79Pgz07
t80ALv1Gsq1AdQtERyHPK5aFvzrDksbF2zQcqYe2bU9siEVa/ryJD0BRdH6GkcGJ
cmBhR3XTMBIjWhsPbmYaKj6oYA4oVhmg/k7UaUXK+/1xTMd1yEiC5frjUb3fQew/
LwPeploATBvHzQf/53EygR46OBHU8JR2avgURJY6ahqlw0lXfrIGeB9FGLemk1to
K5Hlwrhebe4HRRrGc5f6yy86mcDmZ1PBpUriQX8Mi7qe17Pw4yEVvn18z81tFKI1
MAOjo36xa4WBXdLP89EXpO7KpHXfG+kNgJ2AY74JqvS3LTaE5vNCN/c4PYw58pow
jIBPlOQ5EvEWKQatEd90+1gwPEx3ZK7TB+AZiPc6cMs/ZTWfkLRGwkZEggDFOy9B
od9tKevuPTQy87dEPVB4EYCpqmJhrycr8i8D+2sLRunza7CiMGttBh1Dy9HQxTAv
3WwPZuCUB/VQHzMB1xmGcl8skz7k8qom6pqgimzzh7PS/czJ/l5uiAg4i2B10D6z
6vn5w1/JZq9PaoDg09Up7bVRTiMPBfe5b8QhJxOscraaXXyosbv4pljwDLyucAaz
aQ+iQ+CYCEbGE69NQFr7UrjibMuiMun3QG35n07XUHnYGrl27tTKv15qzfSAMxzh
y8MpNmSBRVFY9cDjPPgpw6HC83QYYqqgr38Xnw+NPg8dNuH2kRFv3FVgncE9UqT8
Nh1gMAi8jg/qxJwv25aaYhuECNzJYZciIHuet5YoP5HzjLE5NVwo4XzE22biRaDT
gURGfVnmZDipcltON+Gp4TLS7naNfOZ0CtW9pte0g54/SnyHm2yIW6dmLWfT9mCd
rUN4AxlEaSq5U9/Gn7/5NwyYBSZTz1hc3F2PNkzCI98GAoOFJMtLLHXfxuqcM1AS
E61/85QO+tr0NwKDjJS1sh2qUnhiBnnOSGnfpXuWbV6iqBgscnjinPniH3VzTdi2
oq9Rseg4aThwN3RvnrSggt/UpyOUMGA8BDgSPD9xOO6r5wbltGiJsjwMRGmzJE+g
3SrtEwMcw5qr8Fdyo/hsh7Rxptv1k15TP7mENxAvGhJFm9nRY//lDBGc6cUnGDMv
hCH/FdlNx54aBBm650MdG98UrptVibCV14jtzmCPigghf0CW2X6dpf0ire3UOX6U
yc6mVxBWWZ1V9fN7rVL99FGWpfZ0l4BiAL2NtMD0gz/jxtOZhcRNUVqr7OhsVygh
p6qfl+2nyY/Qq1QYOkUHuzudZGBPd8Djpf/eUkNSnaOXAByJ65fkNTz75km7DmpD
ZIhGhUbb9WR4VXrcpa6fBWYhkzmAsVrC0fsjaYDhVwW05iGiwnyr9i2o/GsIJj32
eHCOwe1SCySyulS0j0KrgIMEyv1uip1r1acYXgLx7X0qyvLdqctnvJuEZ6KZGPxN
Fx09Ab74gkB402UWyyEEKT+7DccgAnOVHd4ezdAjVmwdkT6iwBkGhzSavqadd69B
kxcbs6zwfve2En/6kSrJrnYgrN4jvqVcDLixWoaIBDsvNVosZc6fMQUZALLgFENP
pkglplMu9XCdT+aCRgSyf4eOISh05GrTRDPhiwjOEto/JNCZ2po76oa6PktYQkce
tgffL11gd6+afwr8R1RDPD64YMNOSNsGN78BfqlgFDZ6SPLM1HmOSZHYwyXONoap
ukNpaNh6u5WNwTzN4xnGrf/9qeWc8KKhLe/F6zLApFMYcspv56YHRo0TliKl3xD+
m1WYeberajDD3l1M6YfcrGOscaHRk4aVt1aLd6sXhsJmpZnNJs1Rhs6Q+yaMj1Fs
oR96bLSgH/5jDPJFa6JQxaCYoxYpsLdOOzbl/NQP8QSpIE7ajwgPfEYlWEgcjnc6
JZ7lmxrhNLU4UTam2N1jy3FuVMxRQpk0+zJn++oYHQAA5Zqig+6Ddfv9T6ndu45j
xCr44f8soaRBsSrEHqh4mdMglRMG/Z42Q+zJzU72DnC2yH8HdpjfJDl8/qfLFWs6
HbYTWusFZ1K5XHW+6eh1jtPY+5hWDTwdT/8qCcBMIsjTpaizK/6CQeDavAXfUMt0
YR24UmubUCCRL5ythp4v6gU1mDLbQGgjaMZMmXtKOqlYeEVLv+jzxljYVW0y8vwS
8gHfNY0F3z+JgdxzewskXYZ1weh19nP3Ed1amWZWSM0DGw1SDoG8WiDHuO3hdbSl
s8FVh0iC8nWh32mbnt+iUeESDXw9H1XrO2XWIUjMz/7sMH+2VGWl4M4NWraDMwrE
KhjQrL30Wc7ladEIX317+uydLQhLieO0ssL/l0lQuwrbm0yDKBKXlruruhdNRYsE
te5VmOpfuH1ycwmwuiX6+U3ZQCl3q7+xMySPiPX3m/D0mmkH6sTSFwwIz/Ya6XAn
R58qTasW2Jhe89JZQY9Y5tbjwHLhMezKYTKlimAtn8I2Wx1EdGIybDgh37GiNzYE
TnKbmldTYZh+MCScYpryE8K4Of7DrLEzi7yC5hn+vL0WqayAGxn2ZWzJZNcjLC0w
iMrb0y36XQO3bZ0qbdVRCfzAF9o5CKT6iNvNS1pfTndIjVHNNgl59ECCY4m71H0E
r4Is4qlb0vFsWtWo8gg9daf8z0WNMqyt5lnjQ3xdGx69gKU1RQGQp/WyR+P4Bx0U
RN+DpkHgm4UYbDYoGHX4NTyKU5xDGG5tIVjcwQ2WJVtdkB091EQTUJAtbtWs84J8
blKiiTm2SQotdu0w4AyljYutq77lJWjGpUZOgwBLzPpDryLXarHwEyxeMZSwSQ7T
SLd6Lc9AG7Wrq4H3SACG3g8aeLmkPNry0CKX2nZzbOHsYDaeFAO7tH6zknxm7+KF
P1RglpsN6el//MO+OLlvCqEu06hQzwa3EHiMw6TUkPA2C7VLKAy40+BrEIFEfr19
DDr3ms2H1CvPdLwxfiOMeYULS22BodlqnRj8TrqkGHgyjAHrEUUB8qI56fanHPpJ
zfUqJ9gMt/OSdeHK/80H4KNCNRTpwbW0Gn7Nb1TLxCnYbFxbBYufk8MGw0erV2Nx
AN9BMq/wAlhlMGiGEqdF6CVyS7K441GAvAb3RMN25ToXxTooGr9yBEg6D+S7KKxN
A18DyEngS9dES2rnNpIsxzrU74xzCoZeOC0hAQmHChgArB9IotcdDvX1E8z9NAx7
2AtNVY2wo/nOKo1Y1BaSNmK2vbuO/8uoTcC4pwzq+/G62738sP8isIBUbheLze1+
btmPwq12TkHZr61syulb4Ph1mQscjf9s7OzzcJonYRsgEzOvwpxp4tv78qPaWpZq
ls3AM9lJ9cjYocwap1ngZa2LqtBN6hLGuAjLm5rl6o89Ja+YnePdbuKCZ+zQPv4r
WKPGbhkSoPeF6aUL/HzPU0WfJ+6Z5/qohETwI4f1FehvJuHb0WIAJqp8xQzcPzK7
PR5R7A8tySIEpYmZlg2JlTZ9Ig4Eeo9KHMcfawyDqP435WXL6hO/QKKfStw7zx4x
wpPSx6Oilo2e19GIOq7yFqmZaKj9A4ADtulwm0HIdBvrTDQfCB5ON2gtFw6FMdXi
MSFK5YKOy92/VShDrvIxN6az/qrLdiedwEsczJ2KyjSBy0vtrE/9nIUdGZlJSonf
O6RhY1qbwUlsb3BwT5sqsog5H8tkDiaQwZUQZSO5yN8Sdc7A4m+QfOWAsEDZX2PL
216zSDnzu6iqDxQH2C0elQ+5ExYHoRV/r4a9Kfij/IBZ/xSl4zfHM3ZAknKUaOCv
taW5Z1xIrwMhgLRo2yDpirhX2lM76xa6BT6UfC7daeURs8bSpchLihDyxn7wzB5T
YasmkCL2WYWfGWrvrcmTN8ovAfYIn1/gT3PJbooyqwomLFhvfEteGEYteEpXbi1G
JlHEOSwWIyJV/gTDlqOwfFJjmAMq5l0DV9AwYGTjx7TaArlO9MlMaDzyIeKz9nyh
TfJ+HDZXQBZnbnuIeXtIOlcGMHxhsrDZN6kybtUA+b+H2/Ya2uEIPDgRkmYAp2H2
ETmmMbcEIOg/EoeT/4JUxm1DPCIPNCvxzNdVZbIwYZe080azUTnWMhsSDAoLckwE
5uaSVYeg5v1AEJ/7XgJ+5Bfnlfj96fDPPaD3lDQyFs6C5ZiOIMLejrCoywlfORdj
EsCnGBuV8PfUF/96NJ4qEXwkulfeibS+JEXy4ANQEJ9SsUbluCsU6x2VSEiozDEi
+J7VB6Qbr5Qt5WT+zvGAnD4dqOw2I0oROACBJ5rhpWgbthUR1JjItM76RzvaIVmZ
QnbP4ccbDEzicdVTEM1RwLsCOZFe8wnIOIxAXpcMaL04HSNI2fSzULHPC/gCS9IH
TQ4cH/vYHC9cSu/xcRs2E9h9Lw9GLMiOwSQSMXJzic8HDeNIL6s2PIMp491chiCE
QAeb+lTARadjOUGsJ7IUipggFEpIrVEXONs/hcq27mvT05AABYQ7fsyqLI77aJas
qusYgnz+BF0weDegoJZDcAagIgr2djDwUHQXtNY1Df5ZhmrYj3xb89MzFooj0QTP
XtsmE5UidniomjmVfemg/fHrM7kmb8QSe8I+wgrCjvqG3LdxXYMIeAvVjdS5ZW9o
6ug5rlS1QcJ5IbNhq5MSRfM6Laaum0jQz9KS1FxPDoiKGG8a4byPfgO6OoNLvnyq
DMuvQqSnfr0tjc8rQDb4SzTkntdYgc0pb3QHCIcEbeiEkehcaL9J/rSHLKAjYHr+
kgZq7wFaUx+8HVWgJAxYjFWtfTXuffo6Pdt39Mraj3+Tg9v2u4De+xGCAsvIn/f0
TVAmToZoaQdpC9irhIxUTxsmXH/MsvNlUHA8noc+qn1F4fIbmR2n3M7oPYt1VfXj
oW8skRjCv9j/Ws1N2QdL6sgqsYh4HScSbIJsK7BUc2XuxHMxfvjNGA7rbwd5hF1I
agmMnd4ycQi0Xa4U+LGzJqNyUcCyOt+JAJ0H9VDbZeyUwXmwo9ye+cS6YTKH2msH
VH1CfsA8BylUL9mFsghrMXLdkA3KzrIl7NGWm/uCT82C+CNTYoyEQ+P51wey0J2J
ZT5gMbv/lykqonhqIaeISdB5TVfnM/PAoBRQunhK7BJO9ubzUzSRfrCLdX1X+OlS
GBN4SyPcA6FECHUg2/Yk/JyvaGG8F9x6bxUyW8cQKCE92NgsyVOlm7/LFa+qQZjp
/1xjqt3V/eIldYvrZYmfzwxsIxdOpru5ItIEvbuADLA1uo9DxtD6GYrYBcGubkbj
1k0galxqUscXcJRWOqmV+ShnrRj1JEhUe6KuTbKYP+GmwTiXk3y+aGLq8G7rvEeC
sA4k4GuABzjvGSePvUmnbj2QwJjtka65q0T0DPNJWG4sUiu5U0wsJbYi3/ctA2Gs
6mAZnB+PMVxpd8rgot5pMSumaI23h9Aa9BjupJtf2vixyF1URjJq2t5LCMMVuXv3
p4usviJLVTClGemVBMq4XziPz0ef4zIdQu+VauzBEPCyeb+IIRZwgNpm/0LytNSE
4pN67mx+9fyFCuWqzSPR9WNQlK4o8+0Yk+vsSu/0dkIoclALIzOraXYqAt7QHjWo
jIeN0p6VvraY+htQ7sFx8PTzYE8Jsug40fupSRQyw9AnICvx2ALi0K09BoJ6bUYM
884CZbyaNbtc2dv8IoYgzZvaMQ5WuVY9imkanzmVjcfAMsV8rdbiUbxhp9jZysAQ
2qx2xcwJEVn7HkpgfEqmhxzorh6DSPqmVHmjr3ywd+oiJ7FpcH7sAZQ3VDMhxCRQ
MYAYcq+T0EP/2ALajpiXLt4YdhBV72rxxIkpJv0s+s8rEbYaNn34RI02re9zdbxb
NGtifZPDOLBz/9/COjtDeyS6QNXJH6iqvpjnx1z1gsLj601TB++2PC2SG47nk6pI
KWhJksxlUA8MV3nm7IP8/K6dTiZ7HEaZ0yqa4oylyKJPjyhXRYENXEMxjqhikXcZ
QSz/08n7+itHf/HGKcVg9jvNaTYMPD6yjPYVYBeLxae3/cKoQAWwal6B8ZKs+cIq
jI2Y45YDKT891H+zXXhY3R5P8nmwZHRnNks7A+25Pmsefpn5T8KFxRyLyymP2oks
G1bULF6dWQIcc37BYXTGSKcjZQi3we54eeA6EPFcP0UjsMqBvx5Svda+345P4EJi
j8FsqDI9XGWEXiIgFsuyaCcm4Njuq4o+JPoceoOKH5LYZFEePMw/YHydIRgFOJIH
twRvJ2fvQhl8iw97LZONpUJCTjkVty0xZdBHz7KhgD/0fB8Vij3xyOT9qee+vpbT
qb8HwL5pxygSSWeUMsdMkV1zM3O5o7MhqlRL65PUfEPIP8s35PrRhIB7TNF3ErUs
incKu49egkOWj6urgLJ4AlM9Jr1diKFLYWfqBE81SsQB/J6IURyhdJUArImMjOCq
Upr8Q/Cbp/651GcE21t/pqXyhdxTKMPb8Cr9OmxF8mPxsEQM2m4VL4ZCFQD4qBEh
sNOoysFAN5vFqU/spCpiuxFpHRPtpqsn5OMdhlTnMYFN/ZJy/NjroQQruul15HlW
XjBbI+86mCKNMkqCFBr8SHPOHjHJmyqpntg9VmUZGQzQHv8wrRON3SgFnZ305tF8
5b+vHjM15zefrlWVWEBnuMYsxt6CruQ3I2vZQI4H7uorXcSFwdcjKzVI/ETv37jh
M45rp+YIX3OWydrDpwH0EnAMHaE2KuV8HUgk8p7VWupcBkg8t5QnAT8910VcWIuA
p0xHGcnCcppIaxP/Yf4tGPwJH8s/EeJoUe1JtEUsD78hBOFDqUHRdyS6NGNW+izM
FgJ//k83kjG6ugMbtdqzKc6F0q2AflDnBbZLglNFp5Eo8JnX5CMtbGX9LbdOKY+1
s79Wxd5uHtLZKX9mFKEU3YjfUsqy2lRlmo15DK5+sQ4aUq8yqrrIaBdXuVpM4GXx
XWi6x6LbKcg9V+Aby2ajbnvlGcZ+nalRyGMqa20bQx2zr9UvWgtiUelkQbDa6N2Q
cTPSkQXqqt6LHtHpSCrSRpKvXSL7kgr52u2iD6FY+6bFGoBlR22WqgbYipjg/rn1
uHYjcin4/WMTLV4F1AYB4eOmzbMJFUITWeZbuul4vp26DW5c5dEvY7+8BkNVLNCB
8fbwC+GZtYCNae71T3WCeSkkT6a4AItKiTBaGnXHsy8FZUUR/cHM5tUv3VcXOTTZ
zuaubm4111MtUQF/H5khr0sAMtct1qlmeIRHXks8PgAIeVrYxb8gWtNvjLpDGxpC
wxlMPRsuemoRHwEb85gzIQPfOToaodBjZGjPLQEsy333eP2phEBkd4oIYIyj2O2n
4XTTG+AU5HLEOsrYsqNjYYDCj7ctoqMxAR330w1DGHtPmIijfcvBvvIC9DIAxf39
CFVUE5lvTznsD51dd7N8N670xbg3Im6qB+DhYKzTvaVE48SRFbtpKpPzKVsrqmFq
2Oz8NNnFB1oPTp8y602ELrwERkaGwhvph+mboY93+ljCt+8Fv5qmmVvsz8IDPrSn
GEWCDHi4Eht6o0zI8cAaSjoTvNdiLyojNBJBTih19PAhj3BUp7pyKWxitwuDJPk/
NQbSQwKJMUQyw965H4TBi2i0EHNfv4AFhtQ431GiFvPf4vgNY7uGMxK3k8Oe7AJt
Vb800hg87G3NXPuWGHwCylprlJNjpm75od7mYl5J0N/Z3iOHLeaVC4zvfMPiJlt3
dc3DHI0MH/J00OcH4LPGz5bsa3kBD1f3fFymkM1nDszXgLIkOqmI/mmfJEB4rMHn
N8u1TqAMfr8Fj49wiEnxuqTbtXTBsz+WDsVa/cqijf93anWdOKiqm33e/ni+xdSh
hhEOM6zlbIvNT/kPIDZqhqMqC2C7xen5nCfmCWwTeQh7lQg37H8M38/9wLD3RBQ2
Thhkbtvrk6oxVBhIKKKRI3J5ZXRRdLoisfSfhn+Ck4FgxZ+0NY5dPUpgbKn6T3f8
GhJyXpwCIDvscCz137lilV6IQsWQ2qFefpY39yzEdfhYtIxC67hypgJFOmD6lbaW
kwxgAJJt4388vrCeeAtw9iw4+rszMc7w/1gNNjdgoav8/vNxHJG0D8A1FlS971EC
pabRCPFlszOf7fV6ZzateaZP8TT2OttN3OIyFs1YzdEjgBC8Sl4zXRRZ03Y+G1te
VRqa/IuusLPXTIgrcZ/TJrnDCAYrB849jjCUDpOI1xuFDDh4tJq6REymmADshWHT
879tv8S+zNxmNm4DlNkG4l2Ew3asj3qG4RhhB6Opw5w5LlvQCX1JtLJdjRgN8nr+
RiyhCgib+DhuPixvFSm6wpJNKZH2vHeY+CpOJV3lXHpp4sqUGs3FetCyz9n63fIc
SNdNeHHiPvVQSJJHgN08qskKlH6s5Y4Vc0jNI1HZAKFHsUU9NPz4D3ZeAa3hS79V
6feGXF/33yIcP4g+DO5gOftrqVG3zEDhZb9l1y4MAtaWaHM1hYczZpa7JM7p1D/d
auJCcqhVWBIFPOCdvNJJWzmPnhClRNIhiSxJc502DG1g4tkSrzR6A+Tq0Zxjkb3o
ZwhYR8alFUxXHGpap/lseuuMUHiekJLgE6ZDJ6keDPLp0v9SyRyisG3RBmTb8BNS
FaTeIda0pdMhVerieP1JS5DZP6zsjaPPidVifw4y1qaI68Dy0QMsGnFM4kiIkvdp
sQVbVD8Zv+yA2q1Qvp+ISjkhp5aHr81OorvVAQX0i0/2mXZ1ijaB6b2i9pgWg+9v
VTsyczb1jYOtvaRsZUmI80kszajsbFmXSONPYEd10CAjwaFv+b57AmkCTnd2L1sb
f1EL/xRGl6TZlCrGZ0g7uwGrTs1moxkEDN5kbWXsZhfmIss3/DcOJfQ+aOlXEmWD
hZGQFBBlv7Y6BmjsCZiKFSDWY548Zn+0sETE2igh2FgTB6ClHPfPrh28KOrC0j9z
6WmUs+bCXuzFhcpPdy5jmK14HEXr+PUFj7xuqm1/32uyJuRO0OR5kY9lbRbuQ9VL
aO870+Ao8GoQYfP1aYuGK29z3cVErbU+iH43azTzvGkLMnG9GeQtUOkwSAoxSOlC
5WGkGZFA6ACURlXr+ZcR4dGVP9i4g1f74rtno6BNkW4YGRBO3B3fzJ5j5VDps7bE
7osUjsGNTu0K9c1FRcg+TOsg5+nzyzpU9S/KlttzKkE7K1bhqz7kuxBgc0nluBrL
JtYJ12C3YKqBFa4IwcMyHZSW+V23q9mbySWzh3hp7y8h2DplKCv/Wwq/fXiT2LvM
FqK+ASuerNUq9Qj6ZdexFurVBt/fhPIeW+bmR4YXPMcwBIJgmEBht7Co9q7MR073
QVQHAOR2v63jvxvfJ6gcd0KQsxOUpdFZsapSurTG2L4Ye5dIsgOOi7Xhugwtzsi6
0c2VlGRK/cZoWTORdvZrgN5FhJ0y3r+daZdL661dGFLuq6cFMaqeEX3wO4YrHVbG
RzNTeo0YZn9bNrwqzi+pMqiDodw0RXeb4vg4Hvv1xEL6C6vb0kbiAd9Hz7gs0Iy6
c432deHshxV/vTb7xZL9DjWmKbNYEsqx3JWrBTNT+iw57dSqcXrzPkHNKgDk/yNV
HlKTaf20zv6EmEP2Sype7tb6wWszPsI/wylssvF2boIK5wtvn/cDI7CuNpKHHwtK
FH/Ojw/eKvMMgYXAAAYfmDvDI0Fk/d19SPalwS4Tkdp3wLyUah56etxkuoJmAunE
u+2q3Y8fX7toiAaYUWlmuji96oameWjaWvLMYRl3GkiVAKLzjwM3zPME/hlFbRvo
4XUderAWwWCSWprgjImGymzDxLtI/6hBXhX0u2zcjME3i5gANy+SSRvBp8DwkgbB
3D2pji0EJwLVpmqFgcal9b0fytOvpBj6b6vDQRY8jrpcxiZRcBAj6EIVUOcpvRnG
EIoCuJ5moyJI3yZOSc9LaMVZMRmNFD1DjgvJV88gm7kczoznROsnnjl10BadFPVv
mQHghOmz3Gz2/m7fLAEDohH2xC5tSFBSMMiSNTzkTNPJ+l4wd2PDNipu8v+NFDLt
U2E4VN6kk+irF7AtZ2tSZr0M1QSvJ6HZWCq4jqxg3zQUkvDvHXO6Mbh4cvom6CBt
zVLYTA+suBsX6N8TRFxfFA15hL7lrXG/+pKXjHPav5Eqk2HdlEzxs80MKwO45Adw
1+uQuGG6WQo7cRBQpTzXYHMk8ZBpIiYJpPTfhXkoBB7q0dro+nkMpdp8uvsUYWNp
Jh5ni88Q0HWOgViW34bzkdWbxe+aun2gHC03PSogAupKIwibSqf1l+uCi7Thlw9M
VoRu7ZXlzQTB7cKx2ICExcX8Ur/d7lGPvjQuZabDRrB26vbIh+nbipoXcTbC255Y
NJRC8WMB3a73ss/Wx7Upcr+K58PL5Mio9qr4AU+dYP9/c/zfw84ff+E1by4cV74e
ee83T0laXwJooYFf/SCXoFSGSxu1S/y3JcDEgX84eu7ojIcGZxvX0KDhrb2jp1Wp
ZbeJuuSu4UkWdzCzJK3NQEUNv+VpmABN/b9SbeRm+StpFnopYcmrxN7oVGDi1B02
9T6rLIqqNGYj5wdmxLNYGj+/yShHjuNJhrKQ6mai0ekKCFHOJC3pZgiOWl8bzjhc
MANMu+FEj7H4eEMCkegh+yG6zvcWXo6DC584o+DvFm5D80Q4yYMcU0VXWdUvLXOm
ueV/MZHhLJyjXpSHFswdLJoW+WjjuFUeIVgAnFXDWYkkW44mIx/sMzYqmiq+T8h7
g9HqZtuimWp6daUkU4dXrnIri0MHhUEJsfKkVxtjk8KhavN5PR4cxHRzX8ICaw0K
P1oFJDIy2pbJVeQ+vDv7AzMPIgTAa4RQhnfYNpgekgWxRBDhm9qBF9bJc03N7KnE
q3gt7g8MgPmDDXeb+W6mnQCGEIxgg5Ay4RBhiG6S8cUHQHFEj9pC7QEG+aiJWSAu
YteNeLTpOrD13RsUchPU6MfXdtFOFMNbyMJ/UT+JAuZaPMHUWO9mCGPtSEw421Z2
MPAOfKKQHZ4btvWuTElKS4hetzFxESlsSfsgyDsh1JCOeXyO7ZkHxE8ThcyMSzEj
55RSQ6d1XjoUXJ+gHSOL3xoOTCoKWEUYU67W5medAidrOXDDi16a7trSy1LVQeAR
MratwR5qdFT905+5XuHCybh+299xQoHYXY6RMJ9pykOG3WiyJkko0fof9E9ClRQi
3tX2qDRKy+bwnThEjNIqTTohyjHOtM4aslFQAUuUzqSFiKUfulBd5lXLYbjTxbpS
HmMjcYqtR5VcPRK5NcgFMCGzYX3p+z/5KAirG8NWDJAkdLq2cO5QTTJl1+zGIZtr
29MiTKpG9FHFVgxmdR22JqE/UPbchIU3Y4V04rgaX0GyQbchBSkZ8ZCG5d+1GSi4
/IbfcP55imG4tYB56tUm6N8xTU4yFEYCnKniBGCuq6s/CHonTVLJbNIqcs+aVlgO
QpCY34x1fu6DdPD7xRHDxgAZ68E1psJS8Q8bOscMIZXzE9U6k9FocIv1lrLp2O5B
1epWmtNlJ8qjgqTWD3yNFj48tfNa6/nKQNC4YbPLqQ3YJ7dM8BurlUosmEt28k23
8wwd6FNfGVJ6NzdF/FVoXOBxmHFH3EV9SiuVaxYI0/X9F3oF2lENQ5u+tPdEH++A
4D6OJxDcfasFYuSmbcc9FP/GJbZ8cp2xbXkQTXln4Eq1ZhPMGmenK0FJPKptYs9/
9Qum4iWh3uk3dKdNySUpcGWQxt/qO0wV2iZDA0Rn2SxDgJ/Rw440B4SkUqclYMzk
mPLoUSxvXfUtt6NRq74yU9jBMwbgpENNjjdIgdBsRzjav9s8/byWidutPrpkZUlU
iA6PweorMANUMos9wzdPJ5s/mrHAFz/zKpntwNEQasmk0wfUmXoqEWR+QfgVn1qf
rwNUUulk94XhnqYdrKbYO1fld+L1TnnEmpHJ/pG4mD1qp1nUF5FWprc8DxAg4GdM
+XGZhvC3CLLM2+xRtdsFuLYthxkiITRaOGKnqOhYsxB+nUaY1/QwD3onhkJ74dxQ
08ajgQzqVwdYX0urTwnArZ2h1WdIZJ/defT6a8QazYen5Jcy2fAx0TOlIL8mSNBC
iJ83qQ4rIsZwTV5eEcvLE+2pQ7C0+6X48UJskH1fwv3R4CdNNdtNioGH2GaJsk6R
uIE5fln7JPBqRDEKUw71+5QLx7tNEFj7COcw9VZwNvRQsZ99B4R6Gl4nsA+AC1MO
Nn2JWodLt5bM9AcaimDiObVpsQgyMQQvjsHNdTHh3B9WkfVJb/X4eYqGn/Xs1s5d
Lfl9OwIQNu+in+SiC3jz9jlyRdfhXNnvoTe8BHl+d1wsl32EsMp2dvUItleD4j+I
YhpfHd1XsTGgfEFk3UYKgNQmdPMxCM6Juvd0gpOjlfb74DQJu4qqojxkFzkQM0Vp
XwTQT7KkPdUbFGCsR1unZI/j5nYerDp73g9ym2kk46ybA+BIMgPZpXsnkuywK49L
XRErCKS8jrNBYA/lMg2KzbsUGRh1fpsSGU9NYlOA+Oqq1MkWudbG3nyPGfy42li6
gQVNpUZ0jeZQG1sAIdjtm0QZy9dPgWlCEXmu/SfpKQuEY1E1VxJMruqS2jDC/hDP
75AYCu1r+HkxrBMi2c2Qlkd8tGvhymxGgkd3jHZc1nCLKUNXCTjBWBASESv4ecjj
ymkDPdUvgaOJOUT1JlYU547ZOrrcjzfwGbkZuh9k3dhgy3FOn1UrJETvIuo+E89i
5olY0FxfX6HG3AKM5o5sHS+mxE0MMI5BdvvzR2GBtrDXp7u3MTeTKoGzI0j77sYW
tzNTIjhpPovD0L0NauaBKu2hjzgiCkTByKqF9MfNRhRDr7SeLV4+GvCs3YfPmi3X
26japYDd7xWfUqz4onMXXfuIUD9VspPf+sc2kOtzQTU7q/bAgn2Iq9RHMOU30Oob
Vl7h2tRlvj+kBhKvZ6d2myppWCw4FdSbdbQBWPfSQh37mcn+ZIfnE3zKl63YcFiU
yBG4eFCJJCXh0kFPF9cHhPKTzSU3VBi3oCm1pBA4xJSSfKsBz99Vqa/azGfk6LG7
jZIUOXy3MxytxzxpbMpL/hlgS9T6C95SRQiobEmMuFNX7hjWOmXLggf+APeG/G1t
FuNt3efM+zJuJ5T0E9Joes2s2phE3w1JNTzphoCQ7YfTqXdQBs4NA78RWTkZmvKq
gJZBcS7RD2qC3wuuvTD8LEUFRiNV+8TebotXN4iNBShXz/9flgmxoyAoYXBL3n2w
XmAhsAIWcuFyGMmpeaURxizP3VhWVw+XL+MeScltv96rpRC/lmxTagfR/tg+p/6+
7Kfaz2RggVHmmlACZwW+AEDqj2Kp0owFBuVNZVoDpByaflGgQq4V/TaQMMHHmlWZ
/wfmszcgFgvOSKF+KnBgtw+pSK04RDOQiYMZG0EY31+roZWREsoaIE0t9gl8vxlN
iZ1NxSlWJrG4wOyYtDCYHB67CqOBHJ6WG6/FVH9K9DtiLt0pNyhS9Uw06hGNEYeA
QGOLoyJJ90nPmN0k7avKym/Pdsl88n8PwCAfMY6CBPTiEmBMD4eq3Yw/8B4Kx8l5
lIEJhPC8v1A/6/837WlzdsAxcCYQBOSqmMtgEmJArTGmXuDSYuuUfgxd1DLl3sG9
UTfagRH8HiuVlAha+wSG8gFLo1BoEDZFcS32dXtihWMtPdozlyXWLv7AOZTix3Fp
sRFMltd5SsemK2/QesLruuMNkGUZq0Zu8X5E7BlMqqlrv41ohhjRajqKEVCbdVOz
BoxTfa2ONVvTy4m1FfWjJdVcn8fF6G5RbWvffibSoPe1Zqin26j6KcpA8q2EpV+6
MNyioAmEhnouPHkNbAai3olC5rV5KJ2Tn3NfpeZvF8oF7tQxDwuxAQAonDTIcnJ3
/ZkJW4E2kd0nza60JN5YTQ6G9YLMynBIVQot18FUxYqzQgL6zWkavFhEf207HRWU
8BuoR4fmHpkgS2KBu0vQtrCneatIf8AfCVJvGU8FKdDtaji0E4MqcKAFusN3Vyor
TbXLag64HtHghr/7L5fUajKEGhmZawu5/Hf89A8iCECCoFloM21B/Qf6Jc34tET6
KCjhmbzeJt/TMIQsdWWKK0HtyR1WzMTil6XwwGmdBmkvC8llAhI2dhLAgeosZ3fz
Hier6IIJkWt5ZkT7VtxG1i+QCsun72/PXtfjEUBkZZQsA9tbgn2x3zq8bvrDKqIK
EcWlp4mDGvObhYv140yEtM3gAk7YnC9gAeN6alEiHfEYewud8m9tyzoWeq4q/KBZ
qY9ss7srEN+Jz3jLydOjiKfRI+BRDrtJppy1RalRSZAuXsBFhTtTFDHPaliEQdJ1
H43m4Txp2QpZkc9JBm+HiJ5rVZsneMeCDCAmcdZXVC1QDrzSJ/KWt4hY4Ra9wQcg
0Ieei3JBrjhiW3D8bTeEEnmnGgA4PPgT8Kh0++lkDYSd2iXUFTyn5R++uvstizUu
MRV+sxcpRSnPlWTlAq3dNJvhMwb2lf86EQNizT6KVZENlt9f6w99IUpWduQDzpKW
CkYo7YIs5lD1Gtqt8kk/I1WDF2tvgjbLRYGElurwAbKvQ7wyYweZHDhz2KrrZX9g
uQPdk61EvsaCONZ4UuryU6KvDHk6444hkLM30Z/hZerm9ghjoeRsO3w8XhdpGJF9
UDJ9ShKhXOxFcFvOwOlPzIxl9ikHCANOhpbkK3MiechQOZcM2/yJAEOW0IriI3p+
28IagV01sWcT9LBhPp4uS+XskggeAL9ryq25alEGltVJ+voFWjIFYiTfc07q7xaJ
9eeZSNvlikERg5l+UJxrh+SOlUwi+yqfjJoVaDkiD3E64BVnPH2p1Y10Ox6VyntC
Wzxx7TDBWseNhu3n4hT1PquVdWlz7jOtyvo1+PqiQ7o3oD4oE2BPAIHZb8XB8/89
Zr4rypFbE7YuTGI25fo/aGnJH5/WXoPHjCHoYE7pgyvME/cl0wj/65x98OCSLIQx
lIdCokkQRkg1yvAFrjCuSHC6k1Zs6QJZwdgqBt6+gbO+vqL+kejo38YICEQqRjQv
L+kUvFUVkPDuNdaClIt0VayCYVlItxoS3bjjyNiTqcihhad5gOPPJhGz1orap9hI
mn//bF3N5h9LhOGollptZCP0yubnG2Y64eh4R+b2AyxrELWSPmIILVhnMfpNOkUx
BWbQHVzW3semI3yuB3mBA/HCsYBbFFdrLfLvYqqanoOrBWElDLZblHfZbproM1CO
wIxhxTaUF6TRWg3d0aUBZe7shCqOQ7E6P8uI5Gc3vIUbAi2tHrPsUV0RMM8ZQBwz
7KsQm3SNZRQzCvrB0yVoRfEmEpIWCGtKvdz7kym23RMvtyz0hm2AlySd0JaH4+7/
lUX+s8SZWPLH12LrSEcj7zCNb9uFaCvzkJsF9kS/7NkOi4JUpVswsCP5E/TRdCKR
VD2ms02mjkWriH6+efI1iysu4VgTTUktycMMZmiwAPQ8YL2hMtp+2+WZY0COc0v5
ZYSaquIu+ILUzRNj3c1YFSSqs2iiTBm9orYwnqBkIRlX7uSU74DnmR1tiGx57D4B
mTlQN9AVzy8fH+jfxHzClb2eIWOXMSscM1OMwFAcqUPWdKoj7VEN+drvf8UCQrBC
7xreBFrnakj7TmXy2S+te1bx2YdUp1U0gD2knmUoXe977wopeqmrhVu4QiUD2RCg
quNCg+9NxvPcbSto7kSicjoUf0RpJpdxkEzuj0IUv43LtZqKVELiTapv9F2hF74s
dWGiVyTR+voxHYfvycPtUBCn929c6yWsJ3zEULBJTz7K2WanELjKvx0B7SUtlYdO
u/9cjxkQxWV2d5uPB2G3WUAr5wrDmiVsGm+Qty0Sa2mVyqcWF8EHrpIX58gue19X
GnQiZwWexjCRExs7ygiLv9lsQ4o4uZ86ayPIRCyuhcwviTqVuhcJ4S3VlnpttQCf
NZk0piSacjCCtK3EzDBG4Qd4obf6n2Pv68w6wJfkkpCWenH5vL65gFHnw78xCg4G
/iyczMNNzyySn+xNpJKiKpAUlF0x957lHAulthQqB4INTG4S7vMkHrb6heihvKCW
z6yI0xkjhor92EKyDhdRTFySK02sUNlRChN4eBCYuu+LJ9szukdZxXRGzuEHeL8+
d4WaTOZn4dPK5PMkShgwFNZz3SZiwMv95OjvRfvUZnrz+81KUfhcKXkqzf8dWUr6
l8FM+kKY7Q5SiHgb5RmpxMR2awuXuw9nfxh/ZzgP47BU4IFCTxOEdlrnu1ciiRAH
05BcG845+o9Cl+zSITOI/OuvHOSzZnEiHlYpT5UUc8Sd8NZEKrI1dJorBvqaNfLq
RyacZy4SCTfUXo4GB6iozgxKWXQS+reBj2gm1KsFIh1nN6eLihPdnr/OrhLYa8Iq
NntnuKqxxFf3Llmyr1HEZ3dXBEldyKUYY9hYik03OlA0je8GIZ37YH2sHsiV9jtB
fjOtFekoWspksSkIG3piD4dL5T6p6GCL7QUijH6MpRFFtULTK0yERJBlsfuO67lR
VA8+oOhywLpkwIaWDe/fonrZbCDyGDdH8vo7DcBlJ6ypSPsDm6tqHZkPfr3eORg/
0SsKJqle5ckTXLgq5GxL+8ZvXvh4VTLrzcBih3KDz7hMqtEmgPIfGIA1tSje/f41
nqnrI9/i5R4xZwDN6IuQHjYN4QFyzCfzELvxQHB9TzxZ+ItNrZJb4MHWWko1mHFV
295hp1YNr4lo/k93sKkVa3Q5J4fhFnki4ZZA2ZKnslb1Ft4iHTykImW30fdfGPSO
TWXVd88B9fdnTHr5vuOAwU0uu4VoQ2dwVOMCo+fabFIQbkCyIAziMgNkQe8+k9J5
P3LFZ857lbv1qzQsy55iAAWLlx6v5hElEspHbYZXg0A9LqTs0TMn+ceIIo+YYyqy
500TuD9yTuOSqxHIhu4ewx8VbkYll21ncp7dPOnltittNq3OkH74s4tSMFN8uazw
l2UZfluLcW7ljZ7C0e/ZpYv7bjVFiIf6za8PlAsddzxRqusehqn9LhARtaw8rFwp
G7IrWpNcQnty1lgNIGOnoBSZ9BggSVzYCRBTcwe+nb6026mWzdIUlPoqtvsQTgMw
G/zAUdSFkwRv+/HHDx+X9OuTS4Q9DUb+eUmzMC6uhteBzw/hnaRNLyAy69PTIzh5
Lnp2MYHFb1+oDKWTBR21ooEHUDieUIA/BN1njzIwYKYYfFPeTI675jEP3hiCsTkc
oLrNp4aw8kitwF/ZM/6xT2hQI11RWf8i/4hMGXCi6nv0J5Ud2WNbyTgiKuGmIBwu
UwlwCwon3a3tIgTWIX0+rj0sOX9G8Zum6hoUZzyCL/1Y4XhRuc2EI2nW+5RkBvDu
s4saCHnRvF0QbwumlTH8/UcTlw2e4zPWLYP+N1bcGAGhJTC9KmlRKbWIhAzDI9CA
ag48qsRTTtIvWuQH4X4F/sPCikCwZ9x2CHETZkTzqBmxVC8PUXDdXcQM7cEkoRXF
CWYlhtxx9mjcY4EdVA5P+Maa1QoR5VdzKUnxzJRnr1jBZX6ONhh7VMFK+7gXx4nS
9Sv4n1kvy4PxDkDPTqi0GZ5I2e+bdXeqjyjLqJt/lWXy5EJ2fU+IvocA4YR1oxqA
J4aRApAw/xyvnJHcSBJUofkSf8lKoWO2bNmcKq2hfq2RKdWerCKq0MLASGqeR6cl
ZCp18Ha65/VmHFxWN5gf/nE56UOEGIb4jVrX/ZCTEragY9hGCXGH0/EJB4u5AJeS
YsljcXFTWpxO3Jw0w7MbA7A/PBznUJWFSCIeBnaOZ3RM4kpWyKt9S3rVRs2IeDfC
DPlW981d9h0I3HmjO3ER0f0jIfUo6TAvXJspQBkrYGnHM6b76iSemH7kH4KKR/yL
/KQH1vOeBhMb51htXtTl4AMwYCGeRDt1e/OjP8o55L5ZgDHPPPzDxYLsjB+LXgjY
wlT3WEe7JKW8Kx+0voYpDBKR++iJEK9buQSLMf0/6EufhJLXACdUpEg6RwrMIWcI
T7s5UuvJZd6M7+TiViFEnN4tMhmYzVxSY+6NJU5EDDDIflXD9RZQINuAJ9quc/pz
S1VMNGZ4IBdQqMQpqGTSKqL2EDXX++M78K4PDBvUZpQqAsJ7nzeieHwu0h+BiwWk
D4eQg7lTtNX9GiKUhLXedhfVkH430/8FpUIk0Y+J8dyCoC0xKSSku4LM33ecPJ7J
yI30W8/hmp4A6PvSm6jL+zdwODKP1uMZ1JPgcayCUsWgNoYgWS2svE3rEqjoYKq/
21y5vMdyXoL8axWTLvtj9y8aGGbLLxqMXBXfVdmk5j10mVXWyJ6Z9uRcI+soT14D
DO3XkFnrNhyaMU/IMWOoGOdbKsOrZIzuHB/jk67T7MBftbHEXvnxEQg+T2VtPVUi
TyPue7Mljb8IS7CB2xAxJSc3c8RKi2cXIabMcIZ2Ub0R4eX4gHMlX/Lfmi3NzWxL
w2NixDQ2y4JfUAXj/0SoCCC9qFXRjFQ1deGaZ+CgFDZSTkky9Hv0bj8plA5iniKy
S1Vvd3bi4tfPck67xN8kS+PQ1Uq7n8hRRdjh3arhr1IVBVRpeH1EnrqT/XlF6Utf
xUiYlPsdDglGcI78DKDaSpPkDMfAGiU6ZJUoKELNrBc1ubRZwy49rA7/IflUo0UN
fQYJO4KX/31gfoORj0S0PLWYCe5hOM7OzsI3bEU1px2DlTOUi7L2J5h8p/HIUwvV
HemO3//rfDrCtjjxLeQKEtViv4wUXWaS2HCg6jWWSkMRBNzTZr5/SeHKNNR281dI
MX0PlbthTGTgU1IyhWMayQTBDqJrH6I3A+iQ27C5jKsxmGHOu2ZgrW5PpwUJ1lmB
PorYzwWd3pf71qSPF+0yr4s0zlJFsT8Zp5H9t5Y+JAh29QpWE/90e1j4+Hyuz4yr
L3+udne6imGrzwyJdJkzJCBKZlg8HG2CQt/sY0FPic0KpwedhefIjs+/AXm6AL41
/gHdbOHz8dYZ2Zec8sVJoRWpojWIgjCF0KBXlr3bmTyBe1H5ASsRrEA6VJsX6HPt
ro+vTnUcEaSni2sNz+rBYSdx7CSG0MDIGpckgDXnvLzwn30TWpoxhRe+7QkJPsnA
t5UtEyCMlVu+gax/iwDMj9uNio0dmVYvVbx37FGhZyoshbfPazqTjannkJQ5LhLm
XB8ObUZMmODVaIoJvtVJLFUDggwDyfVPN9k0nBhBkOLu2zOPOXg3c/2Ac9b5Qmow
13lznqqxvlxMo0kBegKukiyhLiP9azJHhT1169KWTnGnQXM+F87ZSWxNJ0Bgw1xK
gkqxaNbfkpPivL+LVmYQhSOk8cMHIvzeR+XYbQxhYOIL+78ZMTsqxWBBeH3b4Jfl
GH5ncQL8TAy9ldkXdSaKPEkA/rSih8DAU+M0FvU7rOUy6fqiKtQPTvtyxlOZpsaY
EMnb16RPAjQpdRH+4eai0K4IaKdM8+3iNT+kAG41ypbWLWyQy7bjs1Pb7teqLZiw
nMCU4XCV/104TPcmCUIMyd6zm9mX4L6c52FEnoi/6UtrG4TSmh18w9tqQPNhSulJ
D30yfoNMXK+/EXYrMJVpFYtaEJz99qCJcagRE4NfK4HqGplwkY847KvcG52QXmYx
HK26dm9wbDT8anB0i/PjlmDAzm3e7jO58gK59mGNrGPIOIL1SMpMrFkKkOHeiwfi
syRdp63MLrup7X/ETEusJMswelo0g8bJv6nBNNtMZz3TLqAiZbNnWpP4SBhbtw6Q
ygNQ2Blu0cMr6whJmfT3HHgMgqPGfqwNB0lqj7jDG+PtlkcbVEcLMs5ZH7/Zu6Rt
LqjB0YkGJJqRtCvrvSLGBLCkookLSdtVnXDuLg+puZxVmlkjzmy5PgRp6pJbRmw0
0cBG/d4cwTpjMqQXtS7Vgj6IxZnjAesUU7MLF+ahFhEkO7OiuA+YlPd+vsayqFOf
dZBPAxT3giwkJ5oz8MyrUFSFhWd2XevQT1BpXXnfiMQpIikhD9tbPr0E66Gi+Uti
SzrfVqeUqDfp6313FE1K80uinbK2IqKTpWgOcLadD8nnQux2mWGq+CY0OJFhXGOc
qi9L/yaZcBle8ldwhb6Go8dynTuLHrNiGweltM4OuuCm+U54z0ShI6i8gbwpeqE2
u6f2fEnvbBq+o0IzfyJvTJ5bVnT6g94XWV3fB3mGoyz2SXoboI2dtUOBEEpVUiZS
w9F5vBByfJYItFDCDot9ZeFKLbNcV86Bh/yL9ogc5RKoSt4p4KJFaHEhnfSlUobG
P2c/gnu6ixerkE0qpWOkTdM+zzcZjx6OgT/L2r05TMeI6YlngoWVEpbWAOcT8nTk
+3M6mTV+6ow54xXdIBSSSq2sHLbB2zItp78LEV9F8E50G7v9Av9/kHI5yllj05GU
9ixTQHXSBCiCWsi05DayqXwDjziFURwg3xzmjt4uKey8YcP9jor6/3mZaLUo/YB2
rDocf/8DfQRW+SumwdGhYl6BmyGH3kpSTdwzPG5ZbLPS0wBc35hekh96IAVo/2hX
emKFXUBs9jrho56oKFqnEOlCFpuS2Htp2f2nybr7QoileskRmjGIKK7GrO2Yvpb3
cABT6Iwd1jD+NoOgA390zoQyWsOkY4pFbH6Y6IYyTkTJNIAIin5qONx3jZLVaHyw
C6lW94Dxyx0/N6Lb6PJqRNZrKJDvN7wihS/2IuSLuxUmgJ86CxOHrVwyViCFBe5X
f8MNeMtgtttLN/S4LUf7tw51HlPbw8uqYplVi/mdC1vKhh/inLo3ZUXskb1aMP+1
9DDPjIgN+5MRc0vSxtJe8R/xxYgHGrkcswIwvfqsdb0sq2PrCRct6t08btHWnmdA
a4R9xWyryVwfRSclUvDboEKjax66cAp5E6/E5snKt6tvxTy0dhl9iUUvgpqDazdh
nypst8qVCPbobrG4GP4YUZI0mKa0de8/MtepLTxZuok1S5d5uRrX3xD90RdHyMzG
rcqSL1fkZq4owBFn5nuCNkVzOsPmp8I7lzGc9WSHg70N2yyLZHovPrf9dCwC5vEr
j8A8kHiGrALjQLYgBUfauD44oLTaiiSJmiNAWTxftWOXHlH53S9whNQHMj1sxI7q
XXN/MOx4hsMbC9smlTGOWbfVlDB6KMGpt+plf6Ts3CqL0rRRNnVyBrPwCFSo/3Zi
z1IQVxvLittsgrZxqU55/LkK0wPucsn3uYno2EB4ZfVtCJR/IYw+qaPA88tQXJey
1Pyg4b7ASRCNX1Z6NM4LIwYD0aW2nlYUasMZ2CLPUKukngc2tbn4kYnO+P2HAljM
uzVL96iDxRPugIFHQeWhwvaoZKVykAmaLKMtrUZsGSCtcULpY7Y1bgOlRR4a5IHf
OaQswmfe9yIsgHtwVOpxPdT3DrVcsJmN2fCvCVox4Jiaw09ilbqEOC0tcjrRSQ4a
ux1NpicELfi9t+ln4Df//ovuBgAotyEMrdzTdvAfe2wGEP+g8h0c4PpwAan68UhE
6PrBtZCIXdbX5JCN1JntiQP63YRVqKQF+un+0328CCGwU1SPfEjTamY2m7PDpLNq
Kp6OfxALr+VSYBWv/LL9YA8v0Od0cA0iKtzP7eTcdVXJrUAdJXb9NuzMP6dwZbHc
4cfvaynswlDWfc8XLtViwe/V9Vn1+G0v2j8GduonNMMM5xUuw5KUxEt1Ov2+Yd+g
eecRsRCMJZ3Qt7GrVkDvO3wSrgqn1et3DMCGd0vAaby69KJCLKQPWBfJUZADSpu9
5jXxzQA+t4Qgd7kTAHfCu/6hB8DHqB5rmxoX4ReV/KdF+USfr1HeEHGJxqCCVj2y
6rUe8bwMQb/TlpsVyX+g+RJ3E5SEbHdwNl5WG0xl31JOMj9DNF2/30VWPzyT7sGY
FKfzc+dWMSE0oc8en0WYzEIQTOwQaVdpZNzUG1Nd0EhiZoXH2wUTl9s32NGqyw8l
B7HSpAJSpVYW4q2UvKMTF3GHBRHWvgbE0a+WfPs/Fq0cSglls/K0nZBJ5XHFkxKP
wNwIon7cfktbjczGPp49LP2rkWdqyv0915puQuUIB3NDcJ3tlwC0z7zA013GpNZp
pkkPAdpUY7n9DgJIRCEQ3S6MrpqDvqbIO9GVIu8e1STVHab/WqjSfwr92nO0/VT0
H1CwbZMOoY1sqAvocyAy43vuQvfbwOIEOZ5wPCR7BtcAZTV3OQHmUAl3TtX05XWx
dRDO2paUHNlc64yhtW2Xj2bRhncLMsoOCxePrXtGk4V6YLcciETna539w6x1H6av
P/yyBRqsI4FLuzejZdOtb/ggMIzxTURXAVjwT9pEB58D0qFAsj8Vo8tqOwve6Der
isKhliHiV/at3W8TEJ+cF7lm4C7Q6FF3Yz6vfCOmvs2V99IYgaZ7cGNTHvAaJFhi
Zl4UCwJCj9h4TlJ3RaVwjUqAvGIU3pxwW8jY0y7djHDp1pkMQvq7kpkOfxat3n5D
FXb+a6ZYrk21A0SG1Tpw34Fm8maunLkdJoWwbG9iM416E8w0dNEUDntX7wh2kvE3
1O15Eg8/z6Md7/D7KGEJVQEHLwr4ewC5qrYDTtcYsyAldYwX9KptULkdC/T42s7v
KllSRgwydKI24i1jOpcuogtALEgc5BWpfhk24gB8wl9EKC2UrVqkElTrstmRmiyB
JMBBpdtsYyfkme7kgMLc4R1aUggsJFhGcXTjCz9vcfHdv8ZQr11Nd6nRAhuPY8oA
Owg6Nxt5ma7JovHBYNVAqK5VYZNH0+PBfMEHgsybuvLH0gslZf4QY7hnYsrS1Cju
6OPAoRhmsARhP9OEc4a5EyJ+ZJ9tR8DzORhFD+7OE3CUn1KaYM2MbgHeOf0FLkQD
mRrqg5KrOXvg47SiY84eKnfwjGTnidbWFgS3fmZKhtuvZp22AI4O4x5rrKZBMIAz
aVkeurNncEK1KLF0TjUu6pmlivf3pXIBcWxNjA6nBARrLC7Tb6VbXPmiSCHZbE2Z
KBQvgkKr1qGcuronxmqSOTQJc5U5pGsG+d9M3z29bG5GxIJ/eUocYmmY/X65Ithm
t+mCTQcZcjCJxOKFt/NlLLB36pj6Rm3uul68VJMGulPCZKsIoedsbKjNfKBkQaXQ
efpiBTOFMeS2vHjivYHeiPmXmqNX4mGsdjdbmol9V6OZTDPWvDN6IrxqfjUcxYLl
nhtx3DCV1IwCC0zZ+bALCF6IzEg1WKAp0Gaejc8SRkleGTKnEHIfv9tNcfvKmmad
GmVFbrMRTbnVVtUjqvep4NMEe18oQO+Y1VI4s53A3+ew+D54aBLzvFWDZXVEFkO7
T/LTq/Ua4KALgpMMFXxn3rqfr5s5xEATWFHa+f6Ia91f2p5qmKjgf6EdgPP+pXg+
RLlZwXiUw8vtfHPNLRdRvqcpAzBP5P2Ui3UEjyVSd5DPA2ZHxxn6hEPrdnCi1jdE
kp7beUbVzCyv4BkstSbTDMPXv6Ob13ImkGfbaZgXt7zRT1sSs6nV2VlljoCIhE6e
JQNod7Umlz+pTM41ELM2uAJxiaH6Od18019yrodfvC4/cVc9mgrliDaxgZHIaLAH
nXKyyQhGkiuXYwyBwn8qjdubR6GxoAPhtmnlJUdsjzH3PN7a9qTM+gc12/EYoBQu
cwHO4TA4GYnro/7yOQSjLvVjb1vReHqs0eAoriDf+M22WbN/+O9m3+7Z92mYRwih
lk1wwCtkG5WinfpEob3lyWq/7OiSUHKZlUkjAAKiBESheFGc+n+xOvsrszxh93ec
1QtazlLxwb1+bvle14oBpjNd4Ur5g3/KsoHvOE1GGfbqNaRlGq+yWXCVW7aSYf5F
bSSJNhCRkli2ASWj6Rqyb9X8cpgNuE6ixrdfkGKLHRydiVQ16CuvVk/iZdm7IIiI
QsYNInN7SFIDRGWRgzr0G20Q3Wn49m1nZ+wyZwstbGta1enwhsqTD2HbTe4S4GsB
YmYSySd6DGtwjfCL/AayapVEJloVYdQPmMHGC+3HWZpXLnPbj2bY8bi9jfKI4lRt
+Sa/Y2C93U2KeJK9H4ICYvvUhdj21gSEpM7MM/OwTZXiXaD6Riiu7yjOWgvxXzVk
l7VIr3vg2wIUgsMQeoGR+kinFkP6c4WQsT9ELf9K/qBsvgVfhGYsC349nIAd9X+1
ZpggPpW4ezSTUQesx5aGsF1yEpdDuagtBHCjiN/MgQIAaYenmc5wuIKasEtDQNxF
o/Q9RgiGAGFSiNWtEuG9pXKeobatQ9sig2Ii06IeS/4lC5s8SwPWR/pJoL/abQug
dy+A8+umeI9KQ+TqmbKpp2GTcdB3pV7LNp+EB10yadSrXgCx2Zw1mEOlRAupYm5+
wvSFAeDyePhzi76OYBFbgPnVJOPihGxAccXuUoWjpLrgXJuqXDOnNpI0sWTqYvVD
AkV1imjAGE8U/kHrxStvvUaH+GwwljrzU4CIZVfQtW0EXXJ9Snf4afTmqvobLed+
9hNRQTXr+YahbJt5pppJfvHLGLKndVQR4n06m9SzLdiqtpFISO+8ITL9RJGu3TY2
WyWkdoBQijuAHjFcDed13BQmFssgETv/rVx2Tz8VolhkA/7ph1A0+EVBUKWdf6B5
2ZFRhXdqR33C4IXKGp3VwmX4pJ8DdwSGwLkrsMJYrH8fKn1hU1ZiqP2LEIWgw0Fc
pXc3/Dj7NR5WWfUxmaU44szuXloTR9kKi8WQM4qfjqp3gn4QhB6rhQjSSjhfs1qw
fA3ia2LwIlaBkxJdZcg1epSL+QcHD39D5dbo9owq8yuUr6lfF0Lt9QjyAM+0Ceyu
xpV+LzRIt5MA5xaBd+NjeKn57tiRpQngwnqPLTmTGMgWSX4tjRJIjgGDONOxSQ42
e9P6zCmcB31jEklGZpQRadD5wx7YrUBxM4usEIIm4W04T3Iju+q0qC3neHB6JuXL
0qcpcQTwDLnNRA21oHtp/008Az7U4ilgCRDt16zvOwdT//aiQSj+uQfnvE5PGyFj
MtcNWfzUjT9eAg6M0ETrYx02cX6Dek00c/CLECTVE5YNW2oJzDkNVC1AGYcpGKKX
ZXwfaon8nlkwG63rFmftkjVz/Vo00A++0u9xfyr69hpJX1IVRTizG00Ebg9jh2Qy
rhc/BpOGrLfl1+IlR4QG80Z9z0kySw0q/9gWKPo270F/xcDrvyxgo5c/9tk/Km5G
JyI4qjFyOOJKr97wHDucT4MDD2ZIhrI+YnyeVwZC4VL55d0mWNGg2/nouu4vuAmM
w2f2pZHj7zzf2IFs/iFvnzx5e0LAMya3gnga6Qo4zlB+DaxL+Us14o2Z/8rFdVyY
mVdb+cgvhUYuV6odyQJgM8EinGqv0uerZdtTA5dYM4Oq7ppDiB9SuiE1WP/WOl7k
BI24lELV8raJyiIUg7i/d+sNtH78SWA0gTbOqkbuc2IV0OKFiANCkj86JxvVdazk
d/BRWUoa6cFHf01lXY+x4GhHQpt8wWR2/SJC+fPQiUJt2sCOCEZ48rpSypfxQ3I3
Ro+s3tUQmoKmbAvkHg+ykyHDzgMfDTT7zYTMlN19+owpX9erv2C2WfZV4NY2ohDf
a2o7tJ4+JYfFzRoTzCcl78g5yquD7fPdYlv3fhbuAD4SBfp9arSsJQhoghMvUwPm
DwccyYyNIvTlosZm0CxENwpAHGs4VHTMOKoYcBOyaCYL/q5QXHWhresxt3hIseoI
JBOJdEs36KLbjeXSTiPt76BkA7S4yp8qjNDm4Ie088pyqEKiM2LfVh5m1Y4/9AC1
YBXyBSs0p/w33CaR7YO/fCLnv2At0ufuDW0Zb3a3gySxRW5BjQiepHIkDde+HzOx
A2RFvk9QFSwoe8dOs/z2MQnXbPbM2AfERcFAOlUjaNJpmn/lCOMgHjGui3Y8ghzF
u3eMnFGNARI8UEQE4XNE7e4O4na1/8RVwlJgngTS9WCyVsGmlWRmuwKSDeLFZkSk
fT1jTnE1Dh8FZKSxwiYqisMzzHbPUtjvPXJBnsa8w7Ez7ba3M4Crv34hncHDkQ63
Xs7ZwpWUkPdSEsnhvcRkWrKfRkWV5rM6FvnajrW9K9Pre7CIVuwsBlPgmzUAQrDi
wsPn+r6v4oHbzRNZPfBHt+ckw7g/vkupvOUWB4PXD0IcFZSvSEQTNsi3iwsdldkt
nJqsUXFEAgNzs7ogctNi3RX5OBS45tw59WPFk+8/lTa6taxrdY+dSyk6V/H4ISsU
lssv/Dbv8YF/cF7X2S90aTwGJ6+24YdlBPoXPZJdp2Spu7kq6HhF2ZCUECF+MuFD
ZhkO7LOq37VixWWo2aZmOraSSCX1VPefn/l1JVJPAxx5bYBe6ncOwLbkTMRh2MHR
KukuvuIUhBrOantKtj1R/HEmRIHO092Lns1lA6iebjcH62gIJIV9U4LamFXEASn5
jQIcAKI07FrjfQwM9o93QHWLegeY5njwYaSeqWmco43Eq0Bpi7TAJPxiPw4M4GTJ
fUxkmIqSCvrW9bT+hT+mpzRHHSRYjyRGGqDekSd0cIMsUnk4KZ7YPp5jmSavxkea
WFqeNSXHo47SYbhbXxg8NnhJuuKF9INRERQlovVzBBHQz7kGaPOFfje2D/jE6RQp
hCXHkAEW00H/I0AgfkvaVrWpHwF8gccGYkA7Cq2EsCM1jBoh7Y06wo9+D46eLsUm
rrqVf9zx21cIJ84PEm3yz3jqYOJuAs4gAp01o7YWQwYnELmnQpLuG5IpHnrC2I0K
C4UnygAMlrlpqLXmwf3vCyaaNiAhedjGjR+VylHyr/xJSSC8QGWfgTuvCm4qTWff
2FMOD+HSoLfP61MZswa/Uu4wnqE6uz8MgzR0MG28IY91opIV5R7LZEGk+/Jv4t5v
TXWY+Z2eRehfcGiXqbXL37XPJoDpRdV1hpsFzhFqN7YFuESqfhh2i1d3LA3ybJdv
KpboOh8ocupVgV0nv1XKlwB7syq39xj0CpJsp3UbrgYLeFpmUs4G3Lzbt+AQYl1+
ROzdDG2vzL6EoiE8NMXALsgt/kaaR/9SwBEaLrzWuroJy4/K9dwAO+kLjbYE1Bn3
oPqWn6iPpU+t5GfNhZMgqtK2Cqo0SNSqAwfcuwQMzz9oH2pAo61T1wP7Blgla1Wa
6cGxkm0HSnl6DKJhERJtS22+kHIYJd4lilo6y5DkFYtDgX39157yyoVD5g4GG6/g
WQcapx+ua2EFuqGUVQoltYvOyQ1bvMbwlgtjUr3XOah9Dahr17b37Nf9n7aOnsah
VOjWVpy8qVCTZSeEPpOp6siOHyq1Dvfej3OItwp82WhG7GKQuaL1DG2C0FEfsCa4
Jfn6njJQvhvlAxkH5MmbA4f9GFqC5WBMigylMezYlTY6EddfFGZ/ZaHFlbwOBUpi
5+uHMS82HJVESYRbYn/hP+7FUFyyv8XHXTn3cc0IAD+R72rVhiNx8E5Fx0X9I/N2
5OOFGGXTSg2F9nq4CKhU5sIvhXkSC2T0uXvEwldVIb5uqAO6NUjldHGc/7JYHVdz
aVSs17OBHHRlZQASjtnqA+zX0pQT80iFqAY9G6+eU9gpubDpFJhwcduYPkGRN27h
fRVw0R48nH+ujgxy0F+VLXwsZfvKel2Yk2+qLiqp9eXaUZNFzyhd1No2oht+s2FT
OCJQivjRnuHLIaYMcXzlkDCCf1sQyTtUHWiTZnjH3OqV/ilBN/yEPV7pwsLBtE8T
62IZzxgwYLM8OpEyyO+dQqcdo8nE7F3L5T9u7F69lNqOao7BPl+DR2MqcsB6QUK/
ojD0L2FDwMGc/vZJxpIAlqT88MuFfeiLdYehfYzI6+ujScbJHcFgrNwcDBE0qfYZ
GERzGjK/9dt+N41SFmrzJ2+XzWEKFdlM6FoS7CK8C0InJ0hb9fWbZb6lLxKCdkWF
f+ji6B7aB5sOsk43g3hyUAsfiKKZ3dKtgFkzMaL8vr1sqkeobQ9QHoZAdoECCjh7
ncf0AKybX/E6dwjdOoUsLTqtk1w+4wkk4JDycdyBhR+WFWyl/TnsEuQ/wjeoGNh4
rjYreyKObZ40/R9WSAASntc5rKsYGA84QK1ig8TkMHAZhh/63lPuaXTUruZiQ4no
eyu9Xj5pB3Rhyi6C7I+ygFIjbFnmz8nknv+Uo1sB3uO532qmEY1izoRzJ6rXOl3M
VvyukRZsbRzRusGde2dDkXKaIr+ZeK79JxDuhXHuv98kKH+nGe06hHr0zrhOHztt
bBBlQ/lXA1MqkFwDN6P3YdO2ZLkYQr0XHnh6s+Ja0EvVl0HeF+7RgJJSj1apKm0g
UPSS7Xv7IV50T/XrasQ40gzeORd18bNlYIiQaZNOojwRJqWW+u1pbAd26fqv4sjG
MXWRziKaWPnx+y/yq9M4aRo45IDfJ8SAaxoZU6OVliyJ/jZOh+9ZLHoj9ASPYQM7
G20NGHBXq+Z5Yla5anZ7PikP9knywJV8PBepCH1daO6GNgeVaoCuc0TYgAHCuqKJ
EcwdW/nTUy4auboeAGF5xk6eQf9kXLWxVTRd/Uhd81poESN7pGftKarRe0hvjD8C
INA1tmlqWLSPUv3BW0L1+qeOa1r4+XxBL7mTRtJInhYr8hnLl4dTz5EfTaSLaXWV
5Z9kZ3m+JCEiqlSYYzbqQ7rSwnNKD6mJIPXtncEior7L1Q4SR08cwqjmpWZYj2iq
i2v1Eby8hy0hE0CQR8/By/Xav/kVsl+K7llPplPigz9nsybrz47h0xgHN7VsWSkT
FB2+uHEBPWZHp36LAIbRpWhZiwZ5kKCh17uikakIWeS5kNkhzObUgzLIQvAjc9c+
tNu86yHeMRtCAERkTzDrAYHWMYo4MQgNwMzb1f6kJ49JPUMtrH1kKvwnPZNoSkae
dUDKL2qTkncQUG4TzyNRZ12rl3VthoY4sZwq95tA7YQnjHrQaV+ajLFteyOHfQ3/
GSO4Qbo5aFEwNZe7YSq2KLPJ9lYpGvMyB7tgjjFryNm+Y3XqDjMGUKpSVEikghhm
8wmOT+3zm8bLg+skrEgpOfENS4A+XGc+KSgQc2B4OXeQu96LNj+F7z8kko56Zya9
1HQk0+mc5PSINK0fqaTiwPRRXQ21LHrctlLgbOCefvGWLq3ke50iEnA+TQqsXaQ1
WdJZrNVndiEakSCeKdZjqGsaAtqBN6Rl0t9f3+UT8ELrSb2jUa1HoSYgFkNnLuyr
vx3QV6I5Fwwo3Xdx4DGdVgBZyF7ZzV5aq5NKpoIm2EFyqEIgiIzWg9IJ8ukIXn3B
yPBgwSYGnvLCJ9Xs+1xIeHv4oD4r/KKwikKTGjHbjK+fhAXLMnFYC4AyJi2gQzcS
Defkmfm54vrdw8z4WJw0XS62qa/eIRi4GbYqQxh3/WS0Kpj/OsAfrZyZyPwIZ8qH
JK5OSA7mojujaQqJfXOIVkhtkEM9luURBN2740JRSiUCQhn0CZ38Lm1WXhgW6eZu
ZzGEbi/AQS8Lqz+9THJAG1TQ74zDu0IP9i/y+JCh3Wl3AwVYxJQSYCHMXn0kjAlq
K3noGr076i0WOWCgsC/LNz6T4aSsfjnZPMjoCn7DQD/z1GW0ehqltBcFDXlihCBD
ozKqhsNlB+Qj5uNA4erjCMClCnA5071GFmmSxLomOcVoN1nBRUWRG3IeLYJlBp6J
q/lG77PzGFBGaH/fVw46uYhGDkGGMYVsVF2bZ2F7YQLegFwDn1FzMTAqj4m/uZyt
Lf2WgCKOc7ARO4MPk7yVIxTTsVAsHwYDmQUm4vU5LgSYx3aratazRhi/zEbkfWr7
RJsRhUwelxzn/1zZsDQjG5emAr0j3bH8l6k4Hf2opzdZfhyZcrxscfe+M6uzf03U
OEL3V6l9YTxb8uGJfR5I5B9q2nvWtY327pytUe/5bG1NRwHq35rNUvyAlscbMzsA
/WXXLk5S4PZKnRu4Ul5vs5i1MI0z4iLuK+sTDUqezk+dZqP30Wc68tGIqkQiIXK5
dbNf7JJrFABVp93xU7tfAVDdClNfj1NuWOnmrbESUJruZVcDmCGyJF8RzN+oAp78
uEA5gZ/F55k7ibRW9L2pnfg3ydZmJl7cmR2ETXat/7LUQ6blc1ZjfP2NsH4eANSn
z1H/II7UxR/6Q2q5LEomlvYL8IjdzchvFyRxbljNk9Fsui+eB9Jw1cQEmOyiV3DF
TJh1Vel/U4DPpcbPcIqCv/7OwsGLpDGmq0FeRQr3bh1rPwczWS3jq5mqs/IQrJ3F
VidvISyu/H5XDk7Rh3tLdFX4NUxTbaRg4w0nxXV+f+Xy2syu0LUdFtrhwCyaNIxw
x0GG+Fo0TOl+oi2I5JGslwYbAxsbpe/Ljq5Tsfxgs+ErThUECxMeJF3HL+mIQCbN
3l9LzVP4C6PaMRdrcMubAYSTw+ftRBsQZkTvc+TNe7wFvcLB3Lo2CnvWb0jB9/m6
RZANac2jIxiRgOdcvo8qjOhcxnDco2saVSmbOicr+TWqKp0DHvxkNf4HhaL7s/sv
M9Vhn/4GU8sPTiK2rBSZkrYW7pF29Y+P9xlpH8SbKBA3/cbFsF2ssizM1Pdn6ccP
6WiXdVhrdP+R0sEQG2wv5wFIAR07X3oivtfE/eNK6DO+xnGZMLBrjj35Fy+fS+w0
kMJvCS85ErWgFvPcC1dERBgwxTKfjLKWqEedPR9wkfMeAUbs1oGv3yZeP7XPUtbO
/CSl/fTserDOQlaEfYxDMtfpG8bmqN7U48y0K1D98vNs05AzG+VtCKMbwgOP/gz9
HBM0dCxq0tAyoshIC0qCYImvEUwv2qr+YSRg2OcpQ1D2IW82NFtNGvBsXoWlLnMs
apmlBa2Hp0syglleEmD221uD7+sIrvilHZO2ZOtaZeMUX1gIHktgwfnMS/8cxT1m
o+c5Z//KLIqaclkVRVZq+aDkQ1X8u7VigFJs/0gJERfoo39ltcvkHVdbvmKlag1I
3cWLGdeFqbZLoK58mLyXFq5sJnLcVmv4OmgxAI/h0WIWn8Y3KQxKxV1k4Gs8plQH
KZq0/JeD9vndFk9Yf1v8Ueojx3vEeWfaJQvy+dBzjbYCLtQ2hbDnjFKcyBaF+C1V
dOey3Xp6WAhjP9T6NET0c7g2W+CP04CoXn6cVl5ek0sK9Xo6nAbqSEScXbAYQyOn
nsHvM5U6uVvUk8o3IlJbFnEHQ1w+XVasjJtH0boSoALNw10uPP7bP4brUkBrQubd
EoZS4eYPd5CTPdPEydgqi/11ZbDr0fHc6nC7k8aVlNiOltdP6ObVYi6SFKei1wgo
HdNIoxgjyKo81BpPwty1VMIPpH9K9CL/OsidvYbfX86K+MUSjL0vX8C8AFGTwlah
wv4AiL7YmkWoEBk+GtdoSln6cqy78mbPpeS8AnjPONFwSL9mhe8Wpl9l5ph7PMOw
upQhjFT5U+Vh7cE1disw3ILrnkdQ+gQRAt23gNeai8cSIutI/CrNU8dhKicTvCQV
OzuM2m2dlPL/8fQvzvsaJRINVyalVVSEYqU5FlMwm8+VOLDbgv7mR35dvYoNBs1Z
yA+6YjZzth2rFLGk0U1qY1ZlgJnZAxPxlASSg7vNC5O9yZ91zPt/lYiDBNTrpM7k
J7t9NZGHX/HYk/xY0uIQAb2B3uwZYzC1rHeizWVhYDyxwN/WbvAyA34KP1I2xdVO
XnZ0rCdyC2Jov/cnbg+N9l7K/4DIFb4ga7TLp38EZTjRC38FVRbAlA/t//ODKVbd
bPUoq0DHRTppnMcUcPoIG9hu0rGs2RX30Mdbg6uEKfkmgbYfgfRa1J9wVbiU/Mjy
EWCNOYkbyeydm40HEchz2dBAtEIDGBnZXvV1TVW7dNAh6KQOQwaTG1EojCtzD4uF
1iXRgiZaEtlAqL2pZqiYD/H0Q0RMVdRlrYJBNdkCiYKByv1nNmPgQsHAJLMNO6RB
gmrYUgwRnx3XSAGnvUU9lwh/1IEyTUL5qPhlCuGcTvFPspZ7q4xnBeP4gJhNqFe6
RkGNfPfCI95bQX2ZnA+rbFlH+5KvcmpuPuMQ7rMEDnecmablQsREAXqcuRlXaBsz
zMAIBzE9f56pmdnNRuQ+DqLSC2P4cGeLoeEcYNKqc2CiFtyLhp86ooScvBMYTXKU
F56/ShoFixzzfg6E26j5IJbvSLT1CNUkY45JwO7Oep6dkEa8FiuNj80zh6afNP0o
vSgAORCdu0OUzDGAIW/7KYFAXcoRNSFOSopQOQiqPEKXjShuReZPiWWJIEsOSdzj
WA5ognhFFX8ACgu0BQnh8tN8PzBMNehRRvvjW3RTVJubJcFUChmJc/yiBWrq/smd
IocWm2NDYbezR9poE5/5ajAB+G1QIilsqyQ9izKvDkDMbns22+cXDkh1/R1hv4nb
vvzPQEm/ndzl5dTVaf2Js/q8W1anp6Yj18OswO8m+nbF+dZx2tD0vI4Pr03kl1C2
5BYN3RQ4otPLeFAZDGOH+W3HjT9a7heJZp97lc4PAWyIu/4BW4aW4z7JqTrOLaWC
NVBLPUs71X4QVo6Q/JDQj/tRG8MY24NfbUaFg9oIe36BmiCa5ZB4QawDEyGKxgE3
ASVS/90ZKb+7kODcpkzcr3dx1U71FDyCBVB8+PizUUB4gX0kTIXY4JrTdOtamVo6
8MPcDf7yFBvln9PmFGD1YEkueI6l+4YsEdG4z991E17b1ol2BL7AmpWyIOw3I9My
MvqiE1uBQ9tqKzr9feAg4xE/rZ4HDxSt9GIqqlSMl9t029i7X6yi51r1Q/9BXymP
1Nj9sTVLuUG4jLVkl5agEc2ul09ook9WhtDCsQ0VlAmyw7g6aimA8j0gDon6w/Xd
E0WoY8266G6Dylw5GoPFPYLyGSFWMjI2RhfQnejyx3X7VTEDEDGO2yXyTgf4paBL
X332hyjfoKAAXzaDkT2HxUejXzE3Ki4gtzi8Mx2bjsE1fHeWqn1NDBTqGVrrBg9M
Fv6hWgdwUuL/IboKbKfIVhGKZV1mt1NB46vZPRN0jq7JzrtnVgPiTLeoW0lzunJh
8yps8v+UQL1kcZQGMqADD/lVy8/EP9B+VQTB9NuvE589POmHuSOTiHCKdTjJjUXJ
2ye7Kmf9nOV2Sb6KjTCk7sKFLWtXiSCT9i7KleS3vuwHw5hsi3m/ftFSnhJtcqYh
0kAVLsBhr6elhqonmhs4sRbULnwrnXsMGBKAbINfBEX6WHyG40A0MYPkBhX4+JAY
SHgDu8MvykHVqld0uy1JRJ/0TFYJETbDjTg1vBMp1ytxcIuRGr75qUvWdfuRRcn0
yNY4L8gnpXep0toAeJo/ojxd0kZFXGQYxlwutLwf4xux//wSqtd0TLuGc4w+61eT
6tUoT5ARkBNEiElzPklZ+ga0lEwXmmbBq5aWCFCIES4EUoAhwdSzubUy0t8WrWCz
EUSgyk5XrtFwVID/hlDqrEBG3l5hDdVAC+XJiv+GoGV77jTw7KbIgDXuMGhOGV9U
Kk7JI7GfdUFjNLnGvOZlCmNIj8PXk03YI33TpJLhz90hPL38FpnDezzCFD1Q31UK
v0jcA8lya3f54fncc1/iK+xvVjRVbtkGVSRiOqvnDTQg4KJ5SjpW0krd6HX5iWPT
8TLIbrvxd5CduiN1DBoGkkWbuIjS8pcDbXDzPrxNc8V9RV3/8B3XNtapNTZgFl+U
e1jNT0U3spm0gEO5gez6PAVeDS8kkcfzkqpOpgVmboIL0aOxy307CyEE6iQycjMH
Bfy21IAJ3NSD/5BGlRCX89QI+0oIFLvV0O3De9d2It9UxRPywcEBuVs4b6SCXPfj
UMpdGziLWGzfc9bz0iWfeUAup1F+VzANAQuptbqr/vay3NtVVhIPZ/dlmArV4sKq
Qx/FR0AJ2BFyVVJacLcIPh2YukbGLhUbvOT5Ry6CQL2C8WvcYdR7snS3yBvqT8F3
vnpTpsKfRj49CQ3+XZipoMRUF510TU4B0WMh1lAv/9fKNsy/TnI/Bn3rgNyhBVpH
EndEaPn8NKDQBiRQ1veSz4wGpdYnGWTEL+efJbewOBFhE0MzEFHuPccRsIEc5Zuo
UDMPB+/GH9q7PDjNXenAoYuwTsF5ZF+kpe1v2cZy82p94zW1AijRNmZOskOrReAT
OzsVXfDGdC0iLLzQjG0QCx3FvkXOv37zs485aNV8MTAYh1xF9xM/Yl7YtPrMpile
QUM961v0AzhST0BV8EccZkShcdggfQCBUT8Ca2BmBe2NXLbWTMk3rTGrx1gPp2bX
/l4rv5V/UhQZ8mCsvkKZFGl2UvVus4YeQ4GUtci1tzxjbuilquDZezzxJA0mpP5c
HzFY4nNcfnfby4552S1GurumziOWS5itWTen2mGrzd0Kw9yHd6opeFTvIigSAEk8
81jDJgVj0EX0WIe4zUrpEfw1jIfYnyZ7xDFwHIdMGqgALp8NKaJrQ5ND0AtxRiDY
z7/g+wRj8pSTdVQmlwM5tM/rDRwVghPyS0eOMCQ7GBS8nRbdCfQDYHiKGtzi5pXx
Nh81HFqUU0EOF1vuT6V3miWGikmrkCyc0RhviAxRs9vffMav8uQzK+ctOASFeK8l
QZ95k74/dRRxV9k8Ujl8P5b85heiwGHSA/pjk8TqY5DFSFhqVYFH5OoErR7h5Ts3
0WCLS+Ia8K0Pryf/QRIhRYb43nxki7FAJ8ewvNLYVehifx8CSoBcZ+D4AQYt1gax
WV7XLR1eX+KJNZpcp437fOnVWBABLhwExgTZV0YVK5VIfczGXi+shEdjFSdT5TTG
4Ivkvgj8IaLdryr54yBJPHZzmkjGamXaKvYextBkzsRVwQs+HJuW4KRRQEwhpanD
fOnJj7Ql505HU6IIftvekxj0gKcYFv7JX6Xy6t8UrjJcjS7V+kOAfb2/ivnRKkfw
m/xXUaB8VQe3REX0jj+OyK0n0zbZFnqCFO4P2/cujTWM8Wl4ArvwSq5I+DL3xru/
w+t+5VR8fYC7rgH4GuMcFAdoVfGSF4oFhal80AASrbLD9gjfSXtf53yS/fBDQhlP
y9rG1UNqeG0aULitGbNmhGYl6GZUiJVJWIvroVpxkGFa5T06AUxOz9MRlKlPiBnD
nL47X0KZh3vMroZ60+YpGHWGG672Ieaj6PisEofl5zE564O3R3Z/UeBGdoI40un1
jkmZym25rlCbY/Db5qGQOqQAPNuvWih+1TGrQFVbk6JRcY5qUNT8Fr7m6RUkx1F6
1EuwAQd/OL8o8UPz5xku8rJ6EA08O7qFcc3ih9GZyZgPQcllefajd2M5bgS3paxU
WMsuf209umUWcu2sN3N/iE++QEB2hRGwLO8Nhy/oW7JGgzot2TSrNrbvT2Imo0/p
txGivbl3PPrX+Ktq9ZyL/u64XhvjHKnYqYofP/qx4nskj0/wuMuQs4Hl3F02zy30
MGQf6hCJb0G4SNGIEcMx+buxtiJqFXcy8kgVfYiYJ3SBORQNKojhFyYGMmu4n1Bv
T6jMRwG0ZSzS4H8RfoYYjDz1xuzRc5grLDlcYYO98I6zBjXY0riGXM0r6z2Q6yt7
ejW6CDpltgp4huFYOeRaCf63CzPFIVLJCw98mqsSMMoECdSlzeTyh6lVI4frmUgW
sM7YRN+ZPWCTH9mMwN8pCLwNcnH47VDj2v6CJSyFkyValU/NR4l+2wsoBqVbAYc6
Zx/0wG4vF9i81vjRTS1AGMckGZXwp2F++5CtzrUECJS2T2zypNB4sMQw7GPSaiIq
NGgwe2pThOxzJIcmnND9ICWfW6wXL38F3dEp//ND3JsGKow3T6Q+8MnYmm86uJ/d
bGeBz982R4QhvFJVPVKpTKI6VoEVAZjfAOwkc1Q8B+hIwEygYnAQb6eq9sRgiMMY
d4s5LFxS+66oikcQ9+dk/+yt6c2i9cKJYOE+j3ErNlDtWU9nTZeUqeI8u4XwlkWN
8+OKC2vyqQX0Yb14WejwqM9kb+WOWc7mER+/czgFEtXTMPfxIOgNgFl76zCSq6g8
TsUBKGE8eiTNv6s/V5xnycDqkk89haWwDpooUeAKNBx29pUc0hVhvy1Fies0ojhy
qEzdTIIReBDgKkMhiXrniemMD3weqLOt/p6B61cUbq20UAqRUtKhNnpc40VkUHFX
qlJwCPS2/w8S7e4HOCIWRKdTeYZRHXAsVrjtIqxrrsnhAQrPnad2BaDaH8dq8NlC
rv7ruyyLRPiBVHmErWVcfzbBcbBUO3aFlC6vtsdi0kp8pRNJsFOOBzhxQ2rRs4T6
EOb5HSI3VxzGPr4n885VSp07NNSjBrgeuTGcSTRzhwRcJAn+8c5+6n0FzSU9p4fM
2I+PkgM2kgog6N36cfRBIRmfuXKRwQ8x1Nayhw58YXr7oWmkLtbo0mXhPBsebuG4
rgbC7yeoYT5PbR7bSInEuB2ghQcjpsNQy92+s1HHreCrAFBCoghKSi0OSdQ0ZAe0
OyfOYncQoA4PIJVxKb/LW0aK+lrn0UHLFOUlDUjk6PesbW7HNz4I4AOaCPIlxChd
oOXx6GbMhiPHpVRoIsQ6IW5qmTW+YPjyokixIhHhUvu+Vr95yVTBDPqO1gSc2F45
X8FB5X5hc7XuvtZIWz4c28iMrhVDlcqUY5iEDpabql2ruiiiN7wyAEQRBWGxsOn5
l1sWaAkD/hEHxZyA6ek7Lax2e/x3Ky8H30m85GhcvcYtVCQZDkbwMdfazlsJr6l0
vs/3sIxD4SnpfXElwgR//s1ADk+7r9d2AtCG55L7xsCYTiKkcxhiLpVewzVzWAoz
IFeMyyCHq6tslET/LmPJbwhE/2m+H4djW+kyDA1gOFPWruxrPLgNaERLF0Y+govD
rOtn3dKobVlQjmP8sH7y2T/mCQ3m9hR0mWI3Z6UUbcPTW/ryW2kmTvrslx9tXySR
WzatCzHSl7VrKq+Pnm+sfIbt518+YEG300GSxiSqyRALF4dwxg40ARKylOFGFWmm
X9qK8CHbJXJ55wKTFY2+3bEHdR8k0EEZOM8PpIArPXLLPNlOUwCP4c2C49A0hqtn
7G7Ajz591hWbzT8NFfVPuqcVvqSwEJTyVvCB+iqy8a4Ikl30KogWQ/0gBfI4ZSqh
LMYsF/dSoEOKzWRtry/xv4BVIm8G/DFhXq+rMuFdPkzJHvXZnIOxLZOzjqED6tt1
M1Go7+5JX5WfvW0UC4E3Qfyo+UZd1H0IIwh0PUik2xg0c9Eg0SAAG84sAiA0hqKT
MzBxbNV4noP+Bb4zrezKmfleV/ox2PyXqYiGJiEeh6JUW0hNqrR+0Wglrrm1VOQ5
jzxA/5Z1B2IeDJI1pazCsAkcVwDG/F4xThQ67quTqjQ9U0/IH35F6xeeVZpuaMdY
i8YN6LzEEghv1koP7yuAOSMje1RKROulMDO+3iasSlFkcWy6R+1PBWrO6Z4m1L0T
m+v2rag56bnUZpY8tunHNlgdRCs/1Wm3IgekSb59Q5CrL4OlkdSR+HnSZvbCB4gz
yQPt/V6+gLpNmyjdqWo9p6/bn+vRHRpE5B4NzYNMPMdaVfhZ6wo4dWmMjqFDYN+/
VY/a0i4XkPmyGUUoOM5ZRYM46YJSZav/MAY8r6fuITCUVEWJoIWMQkLKdwsKdw+7
SS95edjSApezSdsL39QAT6EAPiWrNi6HGtWf6+58QNWYDNHAOC8AeRxVatmbElRe
6OTseAeLKQJIp3HJWke0WFscicearhD1t822cLR6NKn/KkxZm7lJJXo6vnxLqpMo
9c9dth+fSlTKUwPWeac6TU7IcEz7ax1pMERmrR0s7j5rsl2oe5iUwctSlZBk+ZH1
FoRJZspTbeJPjHIdzK8tYnJoC6X1qsIgrZZjr3b/JeUhJZ05/vBQYuSgCbU27RpB
hDciFf57MITlbKtRcjshNlh+ctG303QKmZZaiiTA/qvF+1Ys4EBBDSPsoa0gPH1g
udBAPHC1FbKvyh2qqaKb2lcA7xm/8I6ITuArtnBGTauPAcY7seE4+EjOlgJupf15
trVy9buzIc8R83El4AYPxxUK88HpFk1mOXHnJhl8yL5uwDvykV+vPMoqrjDCqY9k
CZeBIz0JJsvGFMP/oqtoWlZ9yEMolWv89bhecA9mFKSrjdsSNVf4xACYM26Zw+LK
Y15Zwr1EStDU7KiDb1pe/ckipqrRyWX7l511O3VYL7KZi21W0xUm/D0kHLbuuLVR
6ts4KA4znaisupDRYQaH4lmZRcGLFOwjl+SsKVj1udZDwhLbknd/JjmvL+8n6Sj7
HN8ia9Dh51VpWakZUrvEGvQICdLuoJ2zjzQQI5K/eX5JGLpBF4xMgDZ+ic8zwKdv
mP9noG8TXBWSaBMazkmKiDINS7Ro7KJEbOzZfrFpCzUSebsfBJen0IbgJ3XPCLzE
F+cEJoZ3oUYkYeSCBMnTekf/kPYmWNyb6Cc9/M34m59v1lmOrqY5IvWBsywxEmEv
7eZ4X+kpl7Yp3KKuK4uTcKOteJF9DX4QYLtnMVnoPyOv11E9huSeBbt457yzgUyH
D307ClNz4Isd/UCkTVFgWkYByn7BX818hcCOSZGpx80lkzCdbXfqKula5hUnMQSA
q+9ezpmh//x/isu5vuakelnT6t2wXrKsRS7VNApDRnwDzcajhgh/vWVA9aAwJH4C
p6NR02GgVCXL5/1xCk//MY/VLTiELlTRG9o0+1DL11K/N+oKyqBdEe/OwWa3AAHX
01FGuzm1o2nHW1gu4h6eww37Z7UYmboEaMyyUnrbaxmbW4+R6yjYZ3jEB0kQoCtN
uHltxtZeS2Ygy+2LTTTtzvx5I6/DcFsq/JQtu5/zy2cp5RjhQhMqiWXNxUL69VZo
yro5sJLc63ImShbCqpCF+06qqMNoJNa8oSLMU+VXg027TimaUiUIhxkMZUOLARPF
UhBLe1twjqO3GYIvcuL6jldkYqpgazbIdHhzM2qSdsZUm5eCGL5AaNn1vjyA52wG
u8WWjePi7nnQuSALT5JvkubFz260yAGF+3FvK4ddcUHNrlMN00IKRBGYL1BgA0Fh
VgP2AkVtc2sHCXvKXbkHqTjsxbsSdHxkP88rpVmGTzj4yRnSLiCgnI2SmlK2FZUY
Ns2+KSOwFU+rQVpIFXajgU+RSC8VOGJ5RreabmmsRG6aiYHzFBuiolXH+99nphdZ
gGuqmfoO9ZI5SnWQYsFD8Adohzu7Hx52Bsd/7fLn7L4aYs7yHvCpXaIgavNr2Vwf
kn3Fa4idvXSMI5Eb22NUJBnZuggkssLCt5d6T0J4on5uS5ABq6P8MNxjzeXnwUZv
zY0nSlajQg8mlSZzH184zA5q0F1Ms5QLblEsmOc0NGOG6hKbiYFQuf6evVVz3yJh
Rq5l6CYCCWMa+Dn7yw2UiCeJwN4747/zcWsmgMSmUIkpdC0y6G4UjkRHvv7ueDUz
7eNwtoFR7YmMm8FhwAekH3jWYdlkwjjbX+Czg1f4251iZ2cbjGBpQJR4kcI5AeQh
EIZ77uw8q3qL+QOEXNwTtFy/KjxD0nyCTiJp5Rbe8b6NtUOfgrALY3aesG6Li6kI
/0oEZ1Fb/5h+pzR8UR/b6/pYVtNYz7sigJdz/jBoCAA4dLWakDNtm518RZ/SZibo
ORPBj1aJ9ho4dvm+k44JRRaHc3b1Zluo8m6oN1aYZbsKSGSkHUVfUfLsXhtcgtEe
CimbP9nJQDdzEqw2SVIvLlcwuL4aY24k1g/lvbU/JYWw343Flu73MX8tV8nOHZXk
zPev0cm07JldWmmRw8F70TMuJapZSuXvUZ0j4JjEqfDUttjrsFkaa0JdczUFbtUl
L72Iy9B7g+VJQs1aGAIbYMBPTU/dt+73OvE4ZocbaXjUEztIutZ2v2r+NQYiPEIR
6PCrzOnG9a3xXqAvnVDPGMz8hqhlPeeAWtKEaLR2cGQSaKFylDWdHpxNw7LlTMFj
bxykF2ncKDS0KsTORvI4fs/zxIluyQYjGGlsFCHcuCu2xm6gThhngyTkShvilykZ
/LeDP9FW5AFM8tyf6bvS9NlzvxOvIdQcEMH8LYEKGcG87yFWHz3B/XYCTyqgQX2n
Iv//zOgt/+FKMtzbHoreX59ohKpwC1khY4vRR4gPr/zlCMnvXdn+U/G4raYVfzaU
Z7zBlKM7tVgJEGiSC8AORW4yHPd5s2xxNei7oJaztzeQHod6qx5VG2cfarZPCozH
Jrr9K08ehWqo5V7FRX/uaB9hAivnQdphVfp5ImEKgqsG059kbUKtLF2WYVRficqc
cOLTbUpUIZbnNakKj1+5uezBKv/JAGZZr3arIZgj962yFCGy6BaGqEkyAlqsT9Wh
CvMsAAven7pswolGVU4d7PT9zRLNzuG/lKqerDSCzcVZoLXbqtKzu2iKPA4ss9is
2DbfXNL/mnaVnsbbSTY+CgCDZgJDPlfvWW0VLxAi1p0dbRhTCT8noB82zzlg3A04
nDJk5Hh/1v7vejKBRcEOW3wRJXJTBrHdET1rGAY0eMRA8kW10/0C/5N59YCqaTUQ
eBEDrcNtPgzJY+i/TWyWknwZiPeN/gMF+pzmUDWTrSvZuZplcHLeBSfv0Agmq8vq
2GjGyXZbJBrzMMsjuCHy6cT1hAVOyz9zxe2bvNqJnyiy492TwFoEEy9pk5B9C2nb
yjC/OVcjZj1zUCrXhHXNJ0TcdAhx6cB7uRfmCI4kLImxfzf/HCBVA1BViDJYgAuL
EU1RPeIf4g3c2t6HdM5PuyvMOQqsyZxx0qCzzaFb79PLjc616fuqYER/eGzAd9WB
+4LHd/o+3ZRNx42AN+UlFltkQNAiJCkX/Qdu/YVQfg0EGGZeyzy6APZ49BNkQ9ns
k5hBi+4fKcsp0u0PYpVCeJjFkqdAy8RwF6HmRQifIhy9o9d78ztZNA0mqN8kmNtx
KX+wopP/mD4UVeml4QjuexONgUyF8X8E3cFH8MnRxohA+lJqNfifGdvZLy55YgjZ
TPz2X5ZHbK/s6hX65wjcGNx0NYn7eyHuwne055aKUxJAFTPktjVBLuc5fwvrPoNe
vQyfQKWjKBSt/5vA5zbR2m6e7+eAaFcpwYF2yBSzLiwUgKCbfbuFbbX3dh3TNrGq
VmgkjJ03O6dIkJf3kh1F+ESaiZqvpmnVnaMe6i3v0Oo31sNnDnrqUf/x3D36Y67t
20bFU+7rCR5jZfAbjDUhC0ABCBl14DhYThn9f3aephpqNP0HrOk6TEZD4HKF3pDL
m4KtwUeOA8t5bvJwIdo5ZXoMCU3WN3VHTmSwA5kXXBuhmRJKuXflzVr8FDx9SDSp
AhxbKEKxSAO2q1i2gah8W0Yo+C8cCd6CAUZKBeRHwj2N18Mxv+VafV68tnR9Ewcs
xbnzX0YNhTdyGRnvhNjY6fCIXO0xZwCb8nL6P7/AX3bsECPQBjegA/SICTJAU/8k
Bb2cHGfAH584um9tqYQ6cA0XBm0x/mAQIK3RcUAgz8T5u/BVBEFs8NBZcewl7rxx
IgJFYdbb45rVCNx8Du+fszavJvp0v+xz4zWCied9QfIeGiyN2pR2l0DRiE2J7qgs
SKL8iG/JKXlWhq/6FS15RllCS8JDaqMG/rkW1YFOM8j0rb5LfqVt4AzQ41su8cgj
QuzqgcAuO344jwVTsTOpPcXG7yXKa/FEDBmJM52feloOfKFqWqaAEJ1kM/IIgAQJ
aZUcG6OgtqLzRXu53WiwKViIEWXqiHmDV00itq855y/Wb+zzdmjYZneD2m+No4FL
3Mqvlh5AuAJSUiE+Cv/ajr1WTKcPxbBExWLPRyQ9ASqMRs8XuFThz8uxF2NbHmJu
pM4N1RhP3I+nZhv31Ya/RI829qC/3V4Rhvsfxuu7Z4VOUwdopgchb23IsqaAPPDH
PejzomeYSgj508U1eyYah2Zm8Nwmkugfmd2AttZT7V3dH02fLskrknBr4ojDMUq4
9bOmYuqsoazkJRJtjII9IcDsOGWRFyAZjgQA38+EL4BXMTuK7bYS0SLd9BtEJs7u
fSve4bEMp0/rMrG934kTxUf+GPhmS71r3vSoN9s3wMKLQ3qDrQCUcAHtnEHgXrah
ow3cexer2qiJYcLS/9ZBeCV7dzsHCamf7NKlPYPvBiU8C3EaMG8xF9oM4+xH6tPs
WmDx5Etth9haPQ2R0TfUZCUYfvMNewJQK3PQ2/bxNqooYvmli7nYoKadzQPN80Nt
b8PfemN2ZbiXcU3+l3wx+qKlCUslKrq0kpEQvElRRYHmlpM3eD/0ldNDbtHWSGn2
/BkuEpQ99K2iwtZd3B39zHdqK7n/HBewLymIyYS79+HtZ24nkusktPUUd3kSLX2H
qzCy2kSqh1Hd8B4fX/nUAbVnTY+Qa9+QwoE9a6mwg8piS8kdW0n73awAeEqiRNOc
XLX0m+2kftOqrURb3MJiA4pf+n96mDpHOqeuKwrymRtHT36Z5Rdy10M40gG/yCXJ
sJUoz4mOJVXviJf0dh5yQhEKQg9ySbJ7P6hpflk2SiM/T+9V19iectoxQhTrZhwD
zkgnzgOEmiyeebs8JLEAdMsxI3ACAYC1fYRzmJP9dhKCd2M9hJhHI4PNbAIlK8W2
G92ned0xCIB8RT9ZizonIX5yS72Wt3/fbxgYYL77UKzIPghANesIuy77zhxYLk+t
Gdt08ljEmkD2xt4RH95DiL5kEo9fWUb59w9zzcxMKr3TfyGHmc0A9CVuaWgi9ZFU
mv5ZuFfiPdH3633GMbOWd2yjZlAj7Ra3wNQ0CkTGYRIzt94zhvGlfXrBcRhpxlLU
ZIJZSXUcG9KeCLzM0+sSABuu4qlbslgVIs6cN6qFw4uuQOn6vWLHWx03aJN/F+wz
fCKJncIoEHG76HuF8MPcTd2qzKfqc/GtdLrpSoS05MK3qLM++ZP2SM3APrIS9e/2
eir9fVGTZymfAYaylZO2kENsSeNoDCEwcS6rUhAMZ7jfhwMEqKZ5CmWTwyoLk1rV
vAaMkrpXcR7l6/lAb5MyGJTJF8IOGqRQE8sdBXhEp6mmxjie5o91TixdzDkSdea6
YXea2GNFk4ODTcse8Sdt5Y/Xpn6jXvCxBL4zpTtBEFv+0I8sWyrVkMqau8Gxoi4G
BbdoO7iZALKfgST4Yn7XkYUajBeCrmIyupsv7lkaN2mnryuhpUNzcILqKBicqQxT
SVpNT1dAqIOO9GQadIzNV9TiXIY7tj1031n2unQXkvJlBiiNCFGK5DZVPR+WHz4r
k/mY7on12jEgPO7bALk8FGmTFe1xiLnJ+ojEA+eTXA0B/pzqkK88hxhrI4NpaG0M
XvGwMoUE/liDrUPZnthvvm3/OttxSFmMj/UBf2+cLVA6yLUUv/tiuX8h97o78Q7q
A1CzPElYAyifvlPv5byCfAx1nBaFP800HHwz6P62uA780fsFyck41I4mcPnET2U/
XEcDs7hzeygMXst3s6PwlsUa/u4FymPaMyZaPlmsjJK5tD9iio9XIqMk+zZvJmQr
weIOTDE1PDMS09MYAjLAF6YYnIADWdeMijpV4c0ONoAmTJF+X+ypXRVIgYTWnk8N
zuSINwkrmTnTCLt0CfxRNeWyAbIOuL/UH1ieoZY6XhjgKsO4SOIFfgcHpw1aqA7j
Uj2w1Ihk+L7YKj48eW1UxBIr+0f0sSDtUiAr+stcrW4mrpxc+F3zMzFRN3qyj1ws
rZPykwBDoV1hZVv+w5YS3+PcCYgo8EAQwt7YzyE3Hymg5sSnQcCvO3VE/BY86aAF
Brnk4XMZ9Pjw3JLqdMnXB6//5G3bqNEopybJwAKALdhevq7lv6a3pUFAlaS/D0bQ
g90NNtfO6mlQcPRUhgNnOaVg0WKECes79FjMw2j1SzsfpSqN9em1JGcNBU+CUBUD
jNqwK0qSPz7OeaScw8qneheWxAT6ku1DoiI892z+OD0XzRTfOOJsbtkm07togPuo
u2haU6Fpe5fXTcWoghmD0g1fX5lK6P19eDO8+ZPwkENlZD8gh8nBEEDF4w+Vc4pH
IqsFRx3w78nv4jo4k6yA0YKfUqwpYoMOOfgimtd5BlwckCHONLJQZxMKqBXqZzqf
hlQRyGjXAqx+0IXHKymf51ughr0KdAs//jJWhCwGzBM7R5ofjldbmM+cLefocElN
3631so0yP7kqYFSEva+mV35BA0Cdn5gBM/WDglKhhSB7MepLz6yinlMFjhkofmVK
z+nTp8/eXRYcwS6htUqAY/BF8hI3gjKfSav6x3HDNkVvvf75v163A+fDVUCHhtXO
sNvhdEsA/ezb6Htkyv/9/R4hQ3aAwr9sBPQQ+a1Ldh/47njXCPWFAKc1POIT8o7O
fGpVm+A1b6NKMOH5NZGsFHPrs3rp2jf3LGIu165sKcd2xs90AWo2Ec4s64potx9m
fVenRBF22SwSipP6LUKrcEX8p3Tpznp0fatZ05+84zQqYpUPpj15cvwcMmjuZw7o
pq+1WE26TCxiIpXHIiO7+C92wMY4Dj7OR+dv2UpTIRnpXDpIXq0AYdvNhA5Cmnvn
5zhB4gSWGKRqqYcXFmpRynXDTDucrxye8FnkaNAjg8ttvLuQG2ndzNZH9zxyuzSd
M8ky489QU+9c+7HhfeqwrxhD4Szq9KM6atvzM6diVxThnQHBFyAzCgwJtlAm/luq
r/wJ165Ae0B3oAWyLD08jhu9jlY81m4taaQ4A4crPnoyvSUdbKqygRUWcDPHLrDR
LGmw46zcYIKoRles4RFXGk97t+Pk19YxtERA8GFE2mosfOU/ivhhGvqwOZ+rvvQR
c7toYl/6bWmxDUtrNeA5P6ERJDCh9woDs5FuKp4TY9vgf0sOhWKs2uklLkSiLKLA
OQbbPxj41EQshxHRKWNDW8d1Bg+D6JS5vWhgpfbALfkGJSwLmvu2mVCWkzjZEzJG
MWzKtDR+2NnAjKJd/gZ3VOPGhu57fELmadyjYePLuJa2J4pIw3mm0mqxCed1nUI4
h1yLZtLxO24MtcIVqIyu4v5CHNqgtfBaIODKe8H+lLQ7kr23alXSPbHymsX+T5/K
sZjkOO+TTX7RhmV+ds2bDBMp8fNousQKn7hobTCHxGOObjs8/x+55FKcqcfjk6cI
ISRiKviFWdNne1JRmHxZJRfUJWOtnOTpgN3MmgBIjbsTlmhWj9XQnk/artALWDH7
cXoAwCmqtMnjF00Nm8YLlZNYPOd0zIbn5JVIFCGAV1j2Sl8d5m2R8FEWE9v+vh3M
aTAmjlcxbCKs5aKy7x1RONtLwzK1FwFELvYgeUQory2hBHf/kTOZHwszELaI1FqC
iDuLAN18tQ3e/2f68yiTZfBX3hCnGsYV8NgO1P7yLiPfJlzPGrzjbTelXEJorO28
k3s3gXSM5pKG7NJUJMmCL32CIWiMUvaZpgQeO9PK4yw+42O/EpaMzduFvptjohj8
VisGiel1SQNmxyZZk1SmH1biX/rJ2OphP/yyx4GebZkPgrm1clisATbdx/Pf2i/j
Bn4jMppIkZdj10wQqz3rLZ1fKGYKgoxQ1+IRqefkP/4aBTfZjsFq0b5F3as/7DSC
qJdqsHgWI0MZIfZOpMcrjPFXfa9cGRb1CKFY53wlL99BK/QhpTY2zBXx/uIUoxBM
CqZNf1SW3Ix+E8vII/REU2L8cd2kRa99Mip/WKCT2WYM9iAG/wfublafkv2TeVa7
EO3wwlT0pdsT44pA2dgMUaJwwZn/vd3p/+5F0wo2KWBqKBdbb/GXKK/OfiQxbu6C
4NAYk32iFuGKvClCfcIIoDOY0bVgfFI3BBPlayt9JuNQgOl3Qim+gyrYoGRZRw5s
da+cVxBqIvtj7XAxDlbOBDQomggyTYxgvyvEWBTbITdlLdxufzOmKEhVyronSbRk
ePZ088tpYKgX54CAsmt5cycsYCbdvssEP1r1cjt0GEvFa56apxjYJBU6Nrs+cgIP
HXPuO7DRfHWkkfLcd+fC/Zj/okiylmWmrQ1B6Bw+RpNOSSF9LUICFjn0kOYmDbAP
fibJnaOBKNPpolH4ylelwYM93aaxQ4TAuwYKUTE9hYyS5ZoOI6pSGIcQMt/thmXK
iG1EnIxQprrqtdssDs031G/6LtDm62D99LnQshADvE1qH4en3NMBl95hsT2+NRWH
ykfYXuZpqIWZCK4ZWjor6NIrwgDWaN5aWfSoOTR7e6t/0XeaOvJV5NVY8MOkDGiu
z1oix21HyTtILjSpbEGhnloOKso/Z7I1q2SpCG7Wzg0Iz2GNySY/cZAcNiL7V2Nv
EpQaEh41m5SDGxjLeuKQnpHOx2UalerLzbTgVbmUdMzoLpKBXz/vaNAVxALJGfAP
beCJxPBWj55N2Qfw4bueBHZySV/rRhEaOwuoXcCmRLhdqxty8c9CI/b/hDqeTNIt
X3RlIl0TXh7tSqRSfinh6mmJpt5rHO4HOCoVlorOzO3/7WzbkJo6+1o1zeSOnPv2
5x2i7b/5+1Y8XVMk7tsvuNqcXNVxHD/TJ0LP8b868T6i1IvqGp1tfem5whEvCWPj
+CcuLUce6kyjt2GSdJKsfDpVQjobZxpV+EqlE8Oi9cPp4gM9X52kef4/DhZyZlcE
FTBisoUV0esf8MCUFTJVZboibG4wqQGs67Ib68qzs/M9/p8xxAYKt+6hDvd4iB4m
jvN0NIlRLT/lLoHXMMO6tacqtnwjWq98n/b64pUBtknNAHCGWqHE4lYwHmJcJAPQ
TIwS1YS706qxwj9WdZI4mWHBETZTxOjGzmy37c4gKSZb37JTYRRDLagB+LpFMPp/
8M8sAHeUC5E7jsxHPmy18GSudb7hZK7+WGFkGLtkCaeBcVey8KS87xpG2KG/HHLf
mvOdRbEGsho7XYvFwaj0C2NOJTamjBDnBcR1ZYXrRJp9uz3xNCz4O29hKiUIUrnc
nfoPAP9jtX9q7kzzAoYV9OKeT49Mu/IUFXcN/Ryi6srytJuP3CmNQ1eizK2AK6z8
L80HcFGhR1S5I5CwUducqPTkuzP3DX6kb0pZVbQ6vdNbGAdFG+tHbmzAPNPYAI6J
5MHqu2MNgS2dqW8nsJK+4iCdgzchxPJNONR4035UWKgI5nu+2tG2NkKo6OUjMgy9
W5sShrz+S+UXXn5MGGFq1KstztXLhXPsRGUjrzbG+yntJ27w9+JDaWUCsi8zTQzb
y6Vm/FRciAag6/51eb5eZDOwMbTUacKdVOJL2A/ycADHD9uotIXVBRfkEkl/KqbF
87p+4cHQUeh5PaTzbgADWckNSuBl1z1Sf1GWtHe8jzIvI+23STZ/LHf8PISTR4rp
1ANxsTX7aMpyMZmPw7hRmazGtWFF9adqTZSifSGJsSHfHY3fDom4huQa8l0XGEaH
sEBSZFlEKUkRxm1j6gIBDTG9ESDi+h/b4B9zxajC9k7ZLu6IrvdWzqZhOtIq7lSY
HScn48kBIpQUPTosqd7bF/I5gH44/pkQ/O6pzPS5n4E/pzqvclIy6DaikBOPfuQj
ML49Smxi2aowtquWCWm4urXDgL2iORGmXzbJrvwwJzqvC/ooKtE3f0IqW08+Av5g
pqEBvTsd3ukrASoRVsj/D5Z41T0UwA5mKY4sidu30b7GznGDugg8CiHwi6kUAqQp
pZokYIdX3wXuLt+SBeDJt58RrDc4WyvfXix7YTwmvgwakNCZSm5lSVL2n3Bu0GfB
FH9F8XPmHwJkcT1la/TX1RNbsJwUOGFyKWid0d/kEQAO/b9eUgRSe82SWREpsHaX
2jXJr8YEYESP7dZLy5KNvjJvp81J4wP8n8IWs4B9tuonX6b3V4bDuxcq6CpwpxeI
J9X3fSacQuUz0Uga3qTxmo2/WcENzNyB8CRVziNtPXjJ5trY+1R40WkPs5skJ3ZM
+XF6eIC4tC6OCYNC//6uBtHMZCy/T6Xvhm/QqNMdKrEmlPDqnYHAAovaxCl1gWhg
RcKdZi6KU+0A1ez0LJwqA+gPCQYv8sFubHrotmgRLjVA6fl8R0ta+Xbu9csN7V8s
FC0ecBgJ3OYjhvOXeQ9Y40ran+Fi29KQ9LVRxSWo7EzD/EZA0XipzOlHo413bbCH
zl0601L1ly1Rmf5VyUO/jZpWM6k55d/8pPHpFYmcKJ5H+1655/0xm2rNKj+2tJAk
7jhAbGF7vx5cKPl/53y5SygSEzyLcdCcKmSG+Qbkk5Qq3pgQCym9F+xB9hPbIRKP
1WRuJycHNQQoNQWG/pWukB8lXMDykgesn90ogvYQyretB/bkRSNougdXePaqld8V
JDLKVsjnFy6BJeQnuenzYP3OBsrk7H6bgxajLJztBOqj/hyIAEyONKy1v+PUrzmA
deAAtlSOOJ/8jNniHTg8ojo9E1Hych6GL3O+jt7CBzVtfrMInRZJLQbWLpCCu72M
J35yd4TWL4vup3FFdNopeIsGvaOS6s70ICaOKPE1z3SJ9CX2bJV17xHwtxU0LE65
KrMNa6CVZGA6pB5N/1q8F/UHpqfQcznCngzegT+DctH5kiF5/7YWIccTrRLE96zn
Ex458//EkWwe0VHI4w5eWqee3RqtmBrPO65Z0667SnU43WIInlPQE9lI7ZWWWpPt
XwU0MEEXZ4zVR6Z3vmc8/IGQRkJmjLcebCn4l7F2O6m1kougs4agKabd3ARqrGd1
vQpKwILHDRHOr/UgDyKH2iTWcaeTCsK8bt4XfxEf1yOPG0A0xYknYigoeuSo96wa
erlxoB+RVlhtuUmoSO+wfluTjs8Six2v/z6lBASpeNjn+SxldQOQtZPKjjCvWiFS
Ovu941pp6BhRHNivngHd7Yc4nXEO5MU9pZkigKEsCZbx23JVnXUhhOrDkgeLR6kt
q07KIid+8+Z18qdjNKH2Pe6MVxgrV1u0rOenJNoja6ccEN4YSVPFJzp7a+rUKaEB
LnV51YaJcgQ0oXubnl4yP1/x9Ms0CIlmbLH/ahQyGzWUbP7vQlxJLzt9t02ioGIn
CGPYqh6vSJcRFnY/06KOe12ITUyvkYoVBsnnSN2Rm2iIWyZpLFf5dQvdHsnLjcU2
UX2loetUE8QG1P46IB/mG10DigiNmeXdS0eyx7B/XULeRKxD760i0SeupHL3OgJa
4kmPvt6Kov7K8zGiCc8viZ+gZH2kUAQIM+hKQCIMTIFOmm7lV3a8fqYMRJoaeIs3
0fuR1t6MVUnRJOP4dq5cj1x6eiqNqRfbrIvorlT0G1SZ1lylAjJWB9t3AH288ml9
8tJ9pmVleDYR+PikWUPT7GD+41zjfuZX1/bKGV3enyb359HtVyYR67lcZXZ5wCHu
Om5q1DapPX09MIoflsmnvIx8RwnM6KBjIzuwwCacuBrCyr1rhfjHF1txr+LlK3Sy
zxwITD3wOVUwlnlabWP96nc9MkhBPuJrOr0/JcdIPXYPXWL3h2Xyh1TwFtCNjY+2
2XJlOVdMRxc2vZo6BipXvAxVz/zAKnXewNtliC5ZBenIUn3CJytyzVaBhU7ObeHx
PBYdgj3MKP0EbDP9afgo18aSyzdsc8LsbDTz2vFO5RiIbwsENIt4rdSeIUUmuqkU
XMxTC29OLw53S6oyZaSlqpq3xgzoPRQK1ODlPRlvmefl8AgAyUZe7TiL58np3xrR
KXMqoBKf28KXzVbaEdbTD/NAkVXSVHgHT58r6u3iDaoIVCqUlHrUTKyl4TYQgsrM
40Nsqe4uq3HnmQT7zSOUfBCswKbCfWeIfH3htNTITPcK0YFCFWkbmVoa00/k/4gG
AKzndDGDerR+joGp2Kk3v3RWcm0OQNIdbz+QyznZc/TgQ6M0vhysNWJvHpD6nNqX
E34M9RzCO79IQZIjFMgYvbO3uOiSxbycZ7S0UN8w+PUQ0lud+tdumcK66y+CSI+9
mB4Ev7hdoDN3LTmzrXF8prQcd+hIkIbZvwUpIn+8gMjwQykfFM9qdG8RkWJnZGWS
sgSfUWDSitF9Y69f8wHW4lmFpIFSAD7wAhhueFqjDjXg4p//V5KTYPbLC+lkb1es
jGP7yVF4PpnPZ5jtdCkRgd0PXQiCjBpmk88K6YVrts64S/2qO5hTnaHupJfeEcK2
77azm2P1MsXsDZ+6sXhDxo5YM/JH6o1/0R5yiFM+F+yTIx78fS1MN+CbtWKxK6Y2
W7IsGTykmTg4ysRp2V0bsHsNR7CT2XDjbd1mKMPRdB7sXmTIb2KVsrt1p16p55YY
XpNLbYebDmrVo7gAWdte2Ve/SsY/6sy0af8eSXqSnODY7ju6sXMILoU8hYZF2Da8
GJ/9xYYlSwbfmRNf5Pzk8GBkALQgCxTzkPDpmza4igc8kyzNMKcLVKmmwR/6skRh
KKnGQmZi0Z5UkDE+cd9onK1DKpaAKCR5xPH0PjQiTvZJkm5FnyuCHKzDsHXyIkAi
YIOxnnxRbFqhfyC+3gRK/lDpYO4GSJiGBtrcwF5VfVBxH/79CbN7m6/X2A7GUHv7
ccgGYhpwQjGlzpYc/4BQtAmSoMWHJ1ZRAOVCJJ2y95HJ0i3hSEQ8q+CQ7Klt3Ovr
0xjwz2cYUwXdDkUPaNV2g4Nj+DFZytVecLp8+vcY3Vj0+5xA8+cl3CMkMX4V/Eic
G2FhlI5H/ODaa6eiZG8ZRgAp5Z4G9kZiuoD+Nbvfgpu/NbMfLo3aENICrAnHDpev
rfw0XXUpaf02qcsWrfqVKU+CKMUvwDo2hpsVn9GQ520X5/f5SbBfNaN1pzbFPCBk
TBWFo3T4CTzUD4qeP32swIk4Mih5UIp5KwPrzboSVMJb5DYb1kyLrHWvNVbRMRtj
RL5wWoBfRavnllEEmlj25WgihFK+38jtuZ+DsKTqBzXuGmf9SScLdMi1vULIAPip
eIIschrVEWmJFfnji5SJJissKB8mQBrdS/xBM0t8kygu26ND33icOJDdse2N+gaB
erqKeGOnZrxs+dk/7hHw8ceq38n29a0zTt/0j0r0FTpzgeZUjb805F0sBuo74so2
0qR2A/3dfGkYUXcJmFVqz4bvgILuWM4lRYbYSj1Qtd6BSpIyJIIGC1952PgcS2zK
VvBhGgmAxJIb/tMEr6T5roTfPV1ZhQA+4SfIq4T3fbYXBfLuYeBpiCRd+y10Qhg+
ITYvSeytOzsSWwnwCABXC+4Jg1x3Jp2N8mFbznzrCt4gr32YWnr3E+a7ytHj1kzh
P05xPS+DEwkUet+vokmor0BPTy29C00Rt6YRTlYSkxB9zyJY27Mx2NL/aYz/Bx97
kLcUlhvuqKbb+bkxpn8CdU0N6D7yrhacPD0Y+WZpOZ6h08jkVSdqxGLDUS2K3E45
GFZXtB0iIHzWebCkxDI+i1ctT8QWBbizDtNaxjtrzRXqCzmVfsjCCBPa9lcMG5Ww
8TiHtPB79rk/O0CobT5PZTjJJJW7uTdmlbCedHnTLKSYgu1hNjW5FbKbQrxCzbFc
SnDUiXOR2pbimWqRrbhbIYHhdRK+VVlHoLKBbcRx2vJKdcY3a7JmtAY2dxyIACLX
EmZCvFhhG4aYy5QBV/+gq4QyZ6UdnBbfbrlDzJMtbwvFlGoQyqN1jM9xnFA8qP0t
s4W8CjDj0auR7wEccqIqaEFw6B4+j6JfGnhui+n9UdHOVChaG6qBxN2YrTTJVehQ
tNEQo0gkyGV1gR8ZNbYraRcaB3aZtvseIA2MS/4r4F6InhPmmZiDT3dZL5/CP9rN
47N2DrZr5GY71seGeVkGg8uy1KvLbmJ2ovEZ+ANO6Zz+scrH6H7VnPN5Tbfw0Fx6
MUyvymLwy/ta3VXzg6+muUQFuT9Y84cK+Qf4YuHwjMv3VMSdIU+U4kDWJhoPlRha
xZTkJDOC1BUFpbnJNQpL9Nj7CxcumaPJN0k5DyYYLvvyt/VMpxzhXjzf02rWNAvJ
/6gyWZ1tn1GkIogaqnsPBnlGQf1URZxkZKU0nA7gHSVWtyovS1Nv1L6jBUhIyBO1
XBJs4MyyPHz/SgrtvZn3z7WGZquVudB0bu8DabscYxe9QCePx53/JR80whIWogZg
cAREr5JlQPe6lMGOQLwnX/w+zR1/jj78eyY9CCGVQadOO53wAVoMwVVCLOqcxPeL
x/RZtk6G6wq+q9ms7mtEC3URIRquzXRaWtQj94luDzWi2QHH1PSUHWrsSCjFSbTr
SLkEUT5GDvD04q+hCMBuME9stMJXOD4PzbZBLJx5wTzZXZ6BjwdfHTNJTzMqMx88
DTTzxweMcpxaxsAD/zLSYG/UMvGvsRm1je3jZxLY71x1vv6eS/XARv4CcYbiV7Ab
WZK+z2wBM/0R5Q364dlk/urfGE0/QRq4iv+U7BipouTaX+BsorDZnSHZpFebp1s3
d6Xu7Q+4G+zfyuC4bv4+5xkjEKIurKUPdkSrHwjZu6VlJYvqgE/6LZHE+IByo7jj
85aHj6ad0MsM6Gt0cgCclZHtA5UzbGJH8YFrZiyp3t7ybWsIc/IkiznJqGYjfFjW
P6dwEYlGvUknJz2VmZgKeweNz6wh2NX+ms4zWJWGhTr2R9XLe0B1TxgZ3OgAVXPO
8d317MWNgTGmq938Q7yJv/spx3YKd62v5g4xUAnh/jn7rW6aewSO9RaZcrKaCLgu
DU632QB/ElsKvivpQyBv2jqyRQPjyg1RGgpBV+rIJ4ssJjIkXmzwc4xSAbNxkuRx
KVeLTLgB8OqqMYgUvcGgkkbB1Ba9aJlqoT16cnWTOo0okDj9+vNf22I/yZGK2mvg
caHFzXRpJtuqdqJYjFc0ZoJDb8F+91mSA8u4SH+Ab9TX/81uyIvK9QticLuwm3S9
mev+rBg6mas3GvX8bqOlGqBcnv+QqhNArR58FPveREKRcXG2AArl7NNlkZPcM7JZ
wc/FX994soTIvdiM9EVWuvo4yU2+qnWnWs/prq5kq72YDf8Rofmmr/2HE+KVvylA
tQ6RcRJE0YWl5cfJ2hQ4p+YINl+/tDRIKKweyWJIti6NicaC7Dqso3a9RAkrngCs
GE8pSV4v9ASsJjulFWSwj9z9AXoTNial5yFiIrbE9LbjejxRQ7Cey4r6deNNeO9Q
Gjd78y/Ujw7c0bhsl7XBgJrF2HWPzxMmIfRt/yOXasWxerK7DzPakSUySKY/oybv
zNGQyJBSXCQ1TJRFx06vJh4xoD0sFMsbaHVAfsuIXHAv/L2bwKrG03V2REYLm7Be
CvQeM4B0m/l6O41xR4YPpY9kRMQTtE5wh9DdW3L54sBdE1GgKz0T4lBuJO4dllEK
ffG6SWBmGv33JKfm96QhMouIIkEal0Y7aBYzKRs8PFlJn9IlARiPdZThOj+07Qbo
87h8CGApvn1XXjNK3KL+bdRS+lZc/BwuiP6EyXiyQn63YAXnOjW/ozGHEvfr0r3M
MmkbxHYLuf5IlpkL5bI0reFrpBPWyKfq7nCYbLMc5zHhPWm3Bn3jrVyGiQpBeHII
IxyTfQpKMVtfci4RfjMG+nAaykhpQeW5P/a7B+ogMQ9mDH3tvD2uf+svSh47Kjpv
gtgJ0FyCOEc0hBSDcyNthI/JdMvNeItFvMz9UtMvL2EesHryBZ7GEOvPmSf17RAU
5yPfC8BT7BB6FLiW8OJxD+/0KTrjwLpUvTZsOERuuRuNuL0q80CO+QymEI4hFcDq
R7gRO+6JUgBOThSMyZKrCwo9wAWVL4Qnpz7EUq/kpr9j6iWjDPOgV8pTs65NeEik
WIspZPJPOd6FV9+6y0rRaO2UIK4SRsCxeomeZuONDAREYMGw9B3OH1gYdATVkDJE
m35I1LSGvZg1n7R2Hro2RyxKS/RM4qlLaM9/ANYFzaeWdYfgMILDMhZZiSBhpO2Y
qInzPIXP78e1/RjINSG2HzLiGlKkJEQh4xXdz2ETtY3xUQs5y68ptyA6JO7NgA9k
03YSvQhk9e7ATgQ9SkEl10aW7bu6TzBW1cG8urOvHiGC2z/RH/UMd+6BTKkafS3z
AemZbca4vCuI7PF9OUYP0KjtX0sNVQIyPLOGmdq/x1ycajCfxuZ0M0+Gk8WBq/bF
2xlz8ET60OXKbsNL0gjaFBWoKBq8cvb5g1Xh/nvHvdElNuyjVwDYKwCkdOm9jqvg
ywbUH2S2qbsFOeWiSmurbi99XR623u0jg2vWQ5lKNu3kSwqVbS8xgUuSERCvggIy
IV7HIMFXqayVVjnZESlWsIjs0f9pcSB0csS+f1xD9KPfbvNwPOFf7HKSBcWW7YYB
H/ZMXEx9rwBhlf0V9tPyo/vGr5Yip1a7ILNGuo0LNWAe8rOBtANInJjBSmSp9bAs
i3T1Smkv/a81y4PceJ8NtZK6Mqg2SAlwJ+WhwdLUX8uhGIk+nd9Qm0259dD9CE5G
ilr8k3H+8mK40dqcUDHdBmlgZtQr0UfNgZXIz86z/vHspmeGzNVFTo+ouqI69SSQ
iv0ezbksaq9k7l4hL2LFjv585BwprFxyHcBsS1NU0Fw9QvyBtdtTwEyx9UiR4PF2
VDwEo+ee+DFJWJJDxM1D5gVZ6O9LjJcUs89ryn11+72T5plSrSEoFDmCCVFoCIlq
VRyiKDq8f0BvlpwkISjGVNu/IRdY7Yi6LwjD+MuiqNSfdbz0Tfm7rNlbAzHjODU3
sKSAcptHRaFbdAm0D30toDnvSlt86I8fTsMWFbCeXkbMbCVQH17rr2L2WEeWGYxZ
FGswaPxCEliCtlZT9o8NMSQIa88f6cNh4V1S6vgWcFYLpJTHuD9xyHsCLefABtqy
WDiUIZB99UjiJslyijabXvgLD994f4UwxL47wDuyy9MJEnoSAg0N26T1MiInkist
D2A5hbRSTX8uRxsvPghtkR4xDrpS4hbaLvx2FF0mo/GHrKeRruniiVWVTfFVxFaG
0CCdWqnIQzcx7PUDGOkhAGjnZ9UbWpWp6LJ3ZwKSVhol0mbosqh+aU58sSv8bzNx
GQAUmrlu7C5b8Blk4rIl+BPeylu7MeGKzpnXlbBD2ICVxwCWs14HbZddSKU6s5al
rKxKaU+GxipayQvyJybFBAT/nl5/+0FRTLibSSukntmROIYFIBQ1OddTzQEYekPp
K9Q+W9ygLF6RuWd3J1Mp73/w8Avn6PAkWuAnbsnptTJeeWAMR7ej0kz6xZCpiKEe
V6//SrTNXtYCMuRQXmPvBd9W1NA9ge7Y9NiQ2Ak6fG2RK/XhUuL+T26GsJS/goYh
5vHEZ88Zs0zNVeAMlKx1Y+S5rU7g8dDE3sFNVmKqipM3bLShxf/FxfH2UepvJKEg
wJMjf7CjTpXCWek+yevxRcOm2Ko/o+9w/PI95Ch1H1/VQSEXGpDbswvSVSWKk+ZX
aQlj4JUGwryn0DYFzotZ6SJ0Wt99o8wZS0z/qwlmP6D/ISZxE4HpxMCNoKwfCQ2W
Q43pLLJYqMWFPNmiT+74Wq4XNv8rH5vjvpLFCdsBxtbQNRXNBJZfQ/pKhr9h5KZx
WIFJYENa+7Yj6dMpjpnXgqliLda18kqcpDLA36lM3htWFSo1Z6U9f8zFbe1hUKRL
wRQegz/IwQ4PcxROny4if4bCPrwH5mDwFGTQed8SniJ6/imydGHgzQr0vdddYHjc
901vERBziFeNZ/PkDxkB5mVaTidpvmmeYcJCfVK/631uHZ89mGSbXuS3zB3xLI9v
CyWXUJdWY69pMcb0zLshOmk/VSo9Qeiw6kCS/voCjRn9o2yzdngPaeN5QQvY3GCR
qExU0Tb3efsx8QljtvmEnzsOdxb0rsb/RMQytPTDfR+bF8pwedidnmUdry/iPNe7
Vi1erJaiAVmZ4Ue6YgyFqm2tpka0Hjy3bEBatRjkMADnuQ5ZnvmKvzbmkHK8/LsW
mGcuKhMIpEL1dPMcbDGfgS+nbMGedL8aJ82rc4yzs8Zo8P0XoF4f0zemJgvX4Duz
q1j95jetaLIcGbIXbKeuQxrX02LcDiTr6wEX+Ige8XXlkJenhstCV93tbhEoena/
FMT+H5S6j2hipi8P+zD51l6a1a1JiRFYxpq4PCnMf8N6E+6np/rSK3VuYF0ZPPfi
IOSvxmt8ud0L58hadODjCD4qitfsCAqcD6RE2U+MW7pa2fLZhuhvdKKTxNVutEMp
ZCORAk0O9jKlu0KEkqIcbOPTiHfYim5k3rf+0P3h0Sco5ERvCPnXMI4rXCCx9Vg6
8EvGCdvERfkzGBoTXGwPHsnmssCv1hWqoWRvP3vfDX8vIWVmzpLJEzQjRP4zQeX8
S+K5p68t+fv6+CNxbtjMFjxlYUjZCwsjTW3i9Jl+hkObstWj5qWxpD++7VQIIMCz
g6Y9oGasrI1dH22Dy5VU6e/38/0PaMn3INYbEXR6ud3DCUex3OFl7i0TGyIkF2lq
qFmFOisUQZRrjzT75HrdjQb37wGXVqsho4nlGeSX5z/rGoZcDXIFgL8RIolWXVAO
RsC9hHEmiU/JfE4yP13eWWmq8KpqeeUCPjEunqAzw8aAdOFOL/xaM1inNbALPux4
oSkoJ2Bjxkx8gxbNNmJMsRErJqQchsaXXqiOgIWEITlgwBBaPafSYZyMVQnCIMtg
SBrGnndXjU6abCKjD7A1RjfZT6rUmFQyDJ2Scx28HUw7zZ9mE1gEemhopbMZ2yqz
BrCwf/ezq537rEcbmczhhvmlcRrN7zq9RgRzbOcncTbNqUNnKr8m6PmDqJ0KTfWl
HTzcZtZqAaQA2+qeE6YADqLfAQBVFj6AFBO13fpOe3mzJecQy0hdxCAee3+o14M8
OYNnLxKBayJaRjsIfNoV18nX2oEp56/nqwhHKpMtd4WV2gpFDFy9YnkM+5Mz3q86
Pi726z91U/V7DD79lWPdYJRAsjaCOw6PRcxLchO5B+ye3ueLrVXfIIsIHKKhCgaY
FP3/8PlxRbxuVH0ClsEAiJ9A0PIAyH/H1qYIouSOe+IWIdfjbivPyJLLGM4uccmy
C4yt1UwAhsp2gHaeAOmFq04Ui2wYbcoGT5yLdz6IxqNEJt/Mi775QzspZVmWtyoS
OkKpV21dqWzZqRdt44EIYmm8oxg9aYVpq3uia4y31pqFlZCAd4DU12CVW33KCDhB
2C9bBh8vnR9vPJPahtV0mGy+AqVwJNyP1gQaQ+O69bDrqcZTManfQVaBEs599kOM
1RO/rUQxMB1FJ3axKggqWPDqOCUvptBPAlDyc6eLIv0OnZtF7bBxqdGeLu7XIA2n
zLtIt3eoyFZ0DbzMLVTIq0iNSNp0mK3rgeivKNYZIbCD55AOsFcPrFWiROtHIQlw
36nsjJQ+B6ZQZWvU6xDJPBRZ8HpDmsZXINru6fnlNMZxEbrTggPgCgrY/v42954y
xijrN9KzsEfDVVDKNTSCiLGNj7idfnh4zOUSKW5SOkogZSTkS4L5lR9RFKLb4foC
qStUHf27Jwi0VYf7+4mM4exIIbIJv/CUKRp6KiTjikZz+S8n3SzVw8izL8A7YpNN
d3zIx/3CkwLn7Vu1G79ChCEuqkTHmgRl74NdBuIfvNT2lWP5JpMQUkSl/ZvtmxBu
ER5Reai0EvgtahW+MmWOsNlbaGJs7cSEoaLedNe/XNlKBOzlqB9LAV/eYXoPco+s
U3ysj1sXydDsdaJvLp3X1ZdKrfmXUnA7VVnvLT2PBm2urvTBMADQu2gd8Y5kDHE/
trurG3FtW/uPC9+gip4QMNGpR1rY28iD0o8T+UhnWrDjx90s+yJaMR8hU0n5Dys+
48JG3OPozrUQ7EsUS7pvXvGCy0c6XHDrUPgRjEMNO8usPiaszoxbnfpZjyamx0cP
56lJkVV5ZmbEmcyZLQI9gpe+YyxTL0Ch4hLrkAvA2YJeyuT2tp/AN4vVkgO/A1X2
fZ9xwqcciVE2NT5+5tQCT5S5wrC+Bo28fkGGcr2DbfG5B/epL+OD/VznYe7efQGr
ubBf6bqPRwgYUsJx5QhsuWBStdeOVJ/5g1/YfqD/aO6wtgc3N6L9Rc5Ouk5iNepg
2reMEk+09dQvKv6sUcp7Wc+IJ182pSSQdOeCdF1SARVI37O7bFEOoA64ZQ5vyJip
7CUX364WEHwnWiRSF2ciIMnR9XaVn2CfCRP1cvMNKkgPbW35WZOeWcNDLN5qNvJ4
FQ7O6MUR46ArQdvo88l3Xq8hzNt3JoVQ3EEEX+539Vliwjr5O4JaStNB9mUZpYnA
FPZORkM0gS/VYCTIxEcSr8ulUxaxMom4A6iOl8/4riaFcvZVW7HR6NjI8bWWcpmk
+pKUd/VhgEZSKrLnSLrd0IHH+uBIitfje0sP8KQdU8sMEXdDyQGBD5xEk8pBgmgm
aCEqzw2b2uUjg7wTiBTyoWTUwgeQ/QqBYWVYJjVmHxmCKuYPuxuuAuFWrNl01h/h
gvd6MeAUDBLAz2je8Nubpref9B8VODa3HUVwjKm3Lp5LUGnQuPYuXJJs7vITmf0c
jVO7+99UI32tFjaubzwGXpJ5Vnkh1DWONeg0VNqm0C10HAyq7/SEFLikcaHfv/7z
XcYjV5iyE4n+/fH5NMnauPs9zJUNBDvsDM2gvLL7gAWBvbQf3IrqStUWgwZHR0J1
rHvq8jf6DvRwW823dyPw7iYLnZivkCH2F3KRiOBJulsvNx21YlXikgOcXRIOS0mT
qHbthKT7M5uMfpvYMUgF3FyoonSSxTgkwlDQOeoyoU1r2rVQthru3yY/ZcreIsK/
khur61+H+vecb8CpxMEMOAqp7RgV/GRmrmlp3fm4sOGnsAjVBpxx7Zavp5Pn7N63
gVrpXCvKIQaA88T4NiOCfZqMysEswETtDZL1iUCdhxqjej3lcQWOQyaCp/d6leEh
CHnmPFU+c8zbfL0EGyLWtAPW6YEsVHKWt8AhfacmLDHVoKggFFJjDpALBKtLk0HP
qZl7hMk6eT+nP0+mu5NRR16mR33haYLyWTfuPRi0fHF2bqjSybOzqmVEz1/yyjfK
OCzq3/98VfDEnM12pNGona96ycrxKeMHmfCDxqMFdXrjVlw7KKz0Bn3KoF8ILHVZ
fsBUSCPR33JX/j+7KmKSgNjQkP/WbouhdPJbrXBaFxNkqM6X7R6hGADWjtRW8YFM
XsjGIjc0CAQ5k4HxtuBCpj2ZxTHKLRia6AFW8GtMYvoXTBzJNHruwi8LokbBs99r
fPi1RJ9WlVAXMEFTl2y+OycSzGEtedAAdwUsAVT7bERO4rZeNOSJmLWAd0OgZlxP
0ecuMtCnOGWgiLKEiA95NvFbXRNoBh5lT22bLOAX9pffiEm1HIXhtdQxteDs/mB9
gVuAwddc4k6OnndQhwBJFSpRpNxhpdxlbk0fIM4ooOeq1kGGokzxjUo+7LurhI4v
OT7LXwbjlinAKNzQkajy2IjZmJmhWHAp9V1Saci2o82qxidrkJDg2dXVun6Lm9oH
7RpGNIKiKTGi2+Tlurapuj43HYVWCMLC4tWXxXyIsFGFuFbi31JP8ACe5sT8t5wN
MHTFBZeXXgy8p58d6qEPsaY2uY2LEO3rFe/QV5fuhK0A+LoyCBOao9vzDg5qfEvE
IKlqaC/v5CPyj1pTxsuJx3lweJSq451jmMitjay7ecB0S5fHPtwV6AyM/InALNn1
MiI/5dTS6UHpWodjCAgPqARC1leOlZaPUracRnSCB9XiK4CD+KMW5tBUJPY0TdZr
Xbp1xxlogzi0x6wqxu77Xto25ADuSQTYnFCMvdMn0Ya06yBcNY3shfYlVNQidGhC
hQalVfDfkQEb8icT3adQ1t+Jg/NtJePLK7WsIxQwh5LtKSdIGk8GNOI4z86mLOLK
ozcc2O1HJB/eNDHApOdOWIB4NUSReb5wkknXU/9Agqaj4qQ2tJ4dOuCgD0S4ycGY
nAFuRLhx/4vznyNdOtF8cqlLatKPX3wHJ57hXOHupW8noLchrvpffcrkOesraSgI
DB+KwJxPS6c3PvmRO+FFLEUvorpCL7KX/p/FMxWo5F7S3/pJ/2UuaGbj6y2TaTZT
hRqtbPc78nnIKkF1J1NjEfcIaru04RipiJMPmWAqhWVot509Q0SONHU7PX4Zgbgz
BNnEVe5iJJbonez/6Himiqrc6km5aow8GkgowM02vID/BG+gsVXEsDX6Ru53smzv
1r5IHLaO8584aI4fpkaneUA/0huYInlL9WXGm53TyPGdgQgy/xcaJhUiPvqZ19uZ
XhANto2csTwgWhrLwYwAmapmgSlxkqRF5q3TnQFD/eH+W8nv6I0nu5mourXJsSq3
jSuEUqP3VCymktYy88asb2n+nU9+bZhWAJs/LP9aRFiCX82TE+KjeFgBeXfQ7zkb
4Rk7IwAskoYzeiQ8gD3os508h2LzjN/mVfcYZydxm9KkX6dUr/OuQ3IX0AwpwzcU
clBNfV4bh7gGS1x8+tWKhrj9YEmpbTXy2Rg77SIHOKq5E/gbUr83NdvJwPAwbHyC
uriyJTWFAL6ehIpTe53jh3yjai5f0/2UFbfDzliP1n3YMN3ntYXETFsNv0ZZm2Ub
Q9IstIXlR0ggM/R4a4Nh8aER/Bzgi+4SfXaROXDQx4qaUxKTG0xhCSO8B6Vrsykk
wwlBVjUPQBdHXbHIDuxjoeBJhyl9+8AGAy2B+vn1FZKNzxmcYeMnPQw8TegovQXN
RsVj9rtxSnBC91IY05Cp0UuW6G67QJx+0Ht8YVtBtwG78b+kpct3qdg7QXZq5z+2
aF5dUWjzXeR4i9b4lcUSQZqwCA1tyl0n7+Evbgk/+1aTXcz4ZFQgOnAcHK0DyEJ8
+kTQcj0eq5S8co/Z+C80tUCjzaJsIxI12ZPyef7UkiGrewsAoWgjs54nZpKpyFDV
JyCjItxZPHv4w4rawKXZEOJjLL/vsKRt+bGrngiJsCw31sAP6PWD5GkK7QRQ7Fuo
QJGsSxiPTukJ8J2qUvTf0/+nvPQ+4T+fa6Ia3EP0uTzTG4ACYhui8XmHD7GT1FJn
p2DCGNGR57ZLBlHzGPLY/HJFi5RCPz2S8nkbHpzur1Q5yjJyM0O89gJCpn8dQieU
86YmD6tWEY6aJE4sGXkDyJv5pJ+XXysV4vhKfyd7YQc/J321kC+VGi8k+mrCRYsk
orvsybYlIsM5snO8F4Jn9VfhgtGunX3S9LTvyGM9MkjrSsM5cpz1Ay/4VwqyxhkN
XjapbKCV9qXE6BuuJpjXgvXlUkGLXNU0aKqsI87njUhT/AphyRvxMptE1XMls7/u
u0cUGZ2mkBCWCjlnHjfLFDMh8jFHjIJiSLHlx7m0XOuhdZ8pxxF7jo8Cdf4qchuQ
2iUOhk5YlsvPumUa/OwtTFsLaxLlepGHawNH4xrI3VKrasx/yelcnRj4IpH8AbD6
vjqp3x1JQBxBoMxlakf8/ACBXI+pkHkJF4/lfdnQcqi4had4fSRYZYthnUgT6jfn
vj0t/25xil3VcUOqSN9me4nPoc5YLImqwL67jRDftyjqeZjNr3+4LKwWcSQWLtKf
rLW9vHyIgcoMNTMxj1jsWIwbBJAX3VH5RsrFMPaUuz88t+GGYEZRpmOjK16y8NrI
yONxOHptcaGD8A5mVRSxZN02eI3iDBtvXkpJjSRXr6W0n5vWgJ6jofc31F3OCE9s
P57m5+evExNZZnVgPe1VuQi5GvVQQ9Wh/b8Z6AzP4aSzzPOHiD5nBFJZqtCYNhMi
chpg6ypzX0JuTIXd5O2BtUqRbaj8yHkEPpFamLlGEcAWIYnSKDj/AsFLfcdJwOQO
8Lu5c8ifVdLFaGN1Z3K2FyvPwEKQlHSih3CTAjtsPhvN+5sEVmV8bqOr+Sct7BhU
0un3GchsiwCyUNsWwViTk8EBSqkwMIq6g1rVH0WHC7RFTpUa1c7q93eSW+FWWgfK
un0rYCWQJFE3I/AgABOAnZLyBmuzRaf2iSqjAnNqFspQ9JRDuJCCKvZw8AADCzXs
cbehl+gq910dYMCWFlXQDu+czMsAobRfgmFw9YVFE4hNtlXvxoBa15DFAqGC8Xtj
GPHy0DOUthfV+lSib+leRO2b8P3HzRSwhQ3ewIIU3M/Q6QH1ngJPMm8HVuLOGhAX
KgaNVd+kLQEt0n+M5KEiJ4U4S6U2mNK+BfNl5uKC+ZQYDIHHQQBX6wuMdheqlPaq
Aq1obhiq7XX5+llpxfckX81poLQcjN3fDwvwqDb0luvGZTvxGtjgQreSr2M8R9t1
6yvlFj9PUwInyV8mhyThftyfdtIXOnOaunRnuFjk/mIjglmzJOJfrCoPOq9JPdGN
Mt6S9EXp6nkrYmWw1nfFwtqoawvy02ZDEu1HgmWGxrQPTE5BAGvrktBseVhQ0Ru+
hgFe5ENOT9ImMmr/iu8JY14Hk+GHTmDwD77D3Tw5BoJzAgCHnlfTgx0RbuiEKJpz
Y5HKlBQzR8QG0ZRJu1KWA0nzT0WE0rPIy6vmTYJZsYOSLEQARjyFpeqnaGolKWnm
QZhDLKF14nUUGjKELGGCLFiMFQfWJul1op94iY2AVtiW8EdrOVmZEYJmeXVqpr8Y
6LQrE9uLd/JdNEdNhSafGxJ2zkjaaOmlCLkOkE6ny09YaiI8DkJT/P5ip7062mSf
i8WVyI6gLBJGfwwSG28YvQTiCDKTQcEqGQLvz+L+gS+aBfAH0Aa2QrFk8yNb+5M3
fbmwksc0zFd6wETsKcRSl+uAaCM+8Qx5TOgVYq7HZzLLZZQxWFU00HLzLFM24p65
yI9oMdzbEQD+4lnRBsq2y85z3+RMkmnyDxxM7tlRG5HYJYqy27EYt2o8IOBIKdny
33l+Im1YQ39urygcNRrmw+V48CH585MwksvaaTujHFKiePSJ1RsQwnMi9YYtGrSw
R1SUkuq9vj5tHty23CcQwfcj24O3w10JHxBHWkvkHU719I169ei4RRDgz/bZpPoZ
aDA/xA8NtqSOu9grUoQTVSfp3ofNajPRPKnBqN3qQf01kyP4io0leyQN3itHcAqD
zjFwiAUFfWAWZc4lIa3Jd6CH0nWxc5i5su4nnbPgz1jWIUftrDAm3pOzyrjDZ2e+
HwdSBU/5XeBqHmu3pFid/juU1jOHSEcmnsoU1mCK/sM+/qVq0dVWjq0TWvsksRz5
yuwTYiIKmKeYVu9kIOpLCzeswQUM4rGcef8+QRLFtf3MjVNtyFJ5m0EzQF0mT8dl
5oZegmZoPT+Om0DiB7KG2IECrTK6A2+kaxeGaHVDWILPiMlqocWWr/TFAhqUVMOJ
v4audsbswQnVfCvk9Jx/PS+ULCDu7oLwd7hIl5RYLK9biDobuRZd8sQyHXGVWYzr
TbM7GJm/k2Oih+DBGg2poy7ZmD2joEmUbzR+pN+p9d9Dfop1pPFszN8g2U8ZKPYG
l6RXa5ocmA/XtLLYM1KlbLgF+JxAnVQp23ysXLhAslzT1a8mKDU5UzuJL2RlTw8l
xAAriia+nJ1/YaDn3JU2kuLweKV3JYV1mn13saQWhdbQOkBSbXFhZZN5EQ7H3f60
bdrr3wjsUPFsvjRiBlUNMBWwQPtpsHr3s/i/Eyx0nnkHKaIYJWv/qIf5cIJvNPdS
eLtZ7/1rL5HAuUMbVl1qHWa0jI+3m+mzTJ/yNLkVLniaje8Vr98zrg0FIPQWhmTQ
BN3t5B9PmbG288RuPP2SZhAwoxCaHkcAwq2onZwkgzGwUTD6oToZvrlpxrVHFVOq
XFiEZwV2ELMiWATMbNyBND7CsAlTSC9mn8aceNWDLOW0Fkz383uO4BxW6BDRnDDK
ahPrHmtbDm54AIfkZxPYyLQyXVxooD3DDGGwPU0HMIZCRAF66Q3RCkQMCJzVZlzP
fbKxpTzWSCipsHyn6g/vmQrSleEBPjhTmom1XI/y7eztC6Zy61+htmZpWfpfC//y
E4Imkq+dyRccodHBcs1xyPXTTvOIT9bEd0Ch8wx0HOim3A9+RN/DxWtY2keDzzZl
Dyg0wQvYzjoSyT609z088mvk3wM6Zpr8UgQiOCP0nyjUT4em42ZRUgQ18trQPlBd
BMfwJSHz+OWlsQyoiwNDi4vJVVqQCULw6AGwt4vKVYtTFnLQQFtAFKCaSh9Gsl+U
wFsDSmUItzCMsvom8gzX0LeB1ezkV/rufArbTRlnvlbx5zI+dzKEk60XqUwA61Yd
E7MFOWJw1C3egX7UT+mLsEyznP/zJXQOoY1r+4Ao8O7vmO5V7enHDGyYRRbNjcPg
2F/sEF4aAWAjRGPlSBFaOk0gU+WnHBbd1m9eAPf2nIkCN3LAVRjpVTxuTLC+KU3S
/YoD14S08t/AyPFygOyybepDUX9fd/QleVtfyQTQOuJC9aRcRF8/hJhg+mMxOrRh
+062IPF/ztuB0iUxCFWwMkik/c03eTNwmSXOeIGj7Fu+apzss8OtOOEVRIozMNiB
kP7dTJDlkkafgI8fV4wGpD+HvPu2lodqN6H8u24a8nbqM+XSTh0seFYEoPTah7/u
owNXUv0t2Z0JZjtfkpqGYO7VE9FZCaSZZt4qAeJVsTASqRhUogkOOOJBM2pPdRcL
Zm+QOQJHakEAu1ns4nENh7MlhHWI8Xd1BhtVH0b7Ytw09MVQ62SrAdow40gElslJ
PrPpCFT20FxKXBzxPfNLGugcCXNJGV3gZljTVJPXUC5PZzLsxLRmA+3ax/UgRjjU
VaXwztt5sEGn8pdRElNbrcE8OPyiEJEmy4De48W4m2jn87YQI5dxdjwYzqMSThSe
g3amV6LnYKJzYmoSPq2SFeTERX71Uu2s4P0M4GEomjPr2Bs3qvKmhO2AHtdjP2iy
1Vl4ZTMr3TFjV+BZ7uHwlHCZ3rMB2UcznsGuCyJz2+RM2i6kOGLTYPUkAMSSWiqE
8NJbYqWJPYZExXHhik4plWDjyQ7TZyqDeN/jO6E51kzr/t7a0Bq2t8e1AL+o/pst
y1BeOrfDXSpp7+vKlEPisg9kFch26R7qNtjC6yrv7w7c8XqmzEjNNY49I8709IQh
HZyuqCp+ejcyjnSk7/vGDx8OmPCG2OiPA94YL92G5ilYB/TViOvOCeo6OSpvvvU4
WsJUQwAsDRgOFJIpTwDann686fZayo+Jv5LFfsYatLQDaUk8hf+4l91iklcLXrhZ
PDt14wOoC2LwQcqZwHWuAer6t04XdesqDdcpjBlycXgbrWYES4EnR6kBAojToCzO
gTd2PnCmO1DwRNdhkXjdY8mNuWbxy6wiBKm0KQDRxRhLjXpfr62X2XxwkXxzqfPR
aesKLvObH3MsqprnpTo3h+Dr3QUg2gXDvfsy5u514dZTWqxD1bkXy9HJEbZ8XNlX
KiNt4Vsdo2GOu5wedfql1PJKK8Sqr/gr0++kS/SlqS1gz8WRmIie/z5IOB0criy0
O+iGS2mYK3Rql43slUZLt4uC9HSHh30ijNJ6LnXS8UJCQn3MGsP5ySnsZbckcUJC
bFem/+CHcNL1L9ESTwfZY2PZRS1aIUHQbZ1jQST5IPqCLVTQ1oOhhNH7Cny07oFI
ttNK85dC3kFtRL3a1XNxmLuBLmWz88PjT2R4wSa59grR1UshyW5xJBBG7N0XraG+
/JUv9bL0PR3UMZQVIsMlM3/6GuQPhKnLOLSfBHTagQQ0bXgIHDVyoSNQStYlduOm
rnRuv07FAK1BLXX6ES/kvF32xh9D1fOx89bayn/FmSmrudy1VO8JP/GjOmvFnDfR
OLL96SryO+4a1aTVAFh+0fH0Q4ttIf72PjFYSdabotdrFYnR5UuzuFfxup3Hh+LF
OCIzX7ZQ6gNrULH/auQCabNbUuvM3fI+d9vwsUOGK4Xdj0ClVMMIWdvys3uKn4+y
BOXufpsx48JH05ZvDvJxgvZG7la4XkbYV3gp5T8QkEP1wV7SRd00a/uFGoXCAbyM
AmFklRROhHEBewHe/bOZeUoly43mgubWYYzoMWZpsXYYYm4jGK1ehr6LazHj2yGV
I1rb13sPa8+suIm/TtiWDphDZbwQYI+/7SlE/xmx+nlTw2v8V2+fIbZLa++OjbsW
5W7D5uAx+6Hbsh4RzLGrrH0yejTwQvfSdaN/4HqTaBEA/TdUELys4IQW6bXdCwWj
uutxYLMGx/bUZM/cxguWf3i7Ztjc+6pMWYcYojgAP8rFLep4IseTMqV2tP/zes7M
YWLW0mi2CITluFKJLuaeiFIoUIVRl4MiXaEgmugUA9D6ZyMGkpEYAXo32CRNQn9+
EiOz88UislgfOEzgAoi77DK0y9VTYvcukerkk56rflX8kT5DZzqVOWyywcd4OoVj
2anm0+6PG/CUMyEC6X38Y26AYfh3nvEPgseGlZvSOQmDUz3m0fU2c/vLCDjU71Cb
RuGM4bGNCLGTI4lvTzQOD7IDs6fu4w2fiGlYe9eKkj6/aqnTI8+LQZuVz74d2nCX
9y9qGOanPLnJGPuF0HRusFpukTDVfK2KIr9uGVpDGnLBqB5jnLm+gPpRtWqD+06t
TCTy3mfM8x+Dp87HHZ/d3xG7hqiVLRyQXXE6T60Z5DZ+RmxK9IRsqbc0zNaNXVGw
ruyfZrQmgYRa9Ta15QVMNBTE2gBI/IqkN1wyZqYIqLNTDX8UDSugV7aLhYwErBoU
aM772CmLt12WoV8VXLNChL0FeR30uztAszNgR47oldelXuEW1SZ4mh3L3twOsGOC
X3gw5v+ybSI9fZUfyt1VR0KQHJX957iKrU71kV+Eih318tb3/Qx92BBWoC4J3j2Q
UrVr41m1G+Xr+lXT4Ed/dLXXMOy1TtjEpe6hUqEPBvb2eUdLctRIxMpU817ivlIL
/WNYGys+yvaITofS1GHyupdzEIA4uSLJOAySvgCsG3/qCT67AGNUDwOuSHVhGGQf
YbsdQZyRUZ2MvfWbjkGt63x8M10asZAiC1oGKmvKEpncxTEDD6ZTuLABP/5mU2sf
NJPXHXOwiyscr7xWWSx670vmJiIJzBeYvuX2J+pNBpkge+LyXRi2uYPcmGp5nOJf
p8HobZT0f5wPLOdGhl5fGGNLvpJZhHavU3m9UBhCbIKko0ivjIb2ZWgDHvzggvF0
Y/EEtmmaQ32xNin1JtZbL2MCH9T8/zgt99/fK3onO2DQa9Msdx49aBSkfeb7GfBl
Ezte6RE8eSbCgNscy5G8Z844Vm7f4b+rXkWUF6YnUQPChi0TpeRUIII2TwP5QCdC
7Fdl4CaPlqFcSBn5UX2R/eY4lD2s0zobxAOVyqgc/J0gij6cNopLq6WpihOcmLmK
Q3dfSjMUyIVRN/NAjYedAKciKre5Luai7mNl30+m0rwwadpzmS2clgY8VOYuTSpz
QxrQ9govwMLrE2jwHNknzyhpahJIv2ZeEdzNoSeSnhXvk3DhLpv9fHYQElijZ1xB
VR7be4lApZLQysSrC/InvgzzbqvBrA9AfyrQYIhSefeSO5fdomV64ceY0FL0Afga
veax7guDwu0E0TEAmDN4f136rtV/pYb6XIFT4+J5U4vlvAIY5uHo05AxwkdAXE6d
DHIHsrPTJwLiPv7mr5sWgLMhZM72SO0ih5DZ/RJU+BIJ5I3ROqDcPTO9RnuVT46Z
mShZVpjalK//SmHdmiP6EknNa6ETyHLGEuuesKCKT2Kqdkxw+6KDTfZQfAam1TQD
3PaXcMyZhhRoED3OVp07JeSPHs5eAWt4gFfYdMrWloy25cwDCEavDSRFwnscMs3v
YnLyqsTf468GJCgLBt/Fm96bCODfG8RMOyeBgXKaByocCsa1Z2j3YQrNVvbzsa/E
GM6jB89QPMoIREsrN0IKXaWVDhKImW9xGm3lMAiKlP+k9tWVOtmSMqm5B7AV1RkF
2cgvdvzvVubPjvuk4Zy/iNWuhWkyZDxss4GTq/8GDcMb1d9pzog3rXskwM6zZLjZ
zucmuG60tFeRGxi8CFSXS34FWgAur0T0FiEocfyOO9h31GKTytzr5ZYuq0gDXbBQ
9YC1mKzsqNdzseULm1mAGfCdZ2Cww7ng7wzjTz3vAxrSkZ2mJpHcqi7oXdm7nZ6B
sYstyL0pzw1zrdHY3G3ZavMmY6Jm00jDFyXC1UszBGkoxSYrZ18JJGDofSoqCvPf
g9KLGZLrDaqyy+Kd6WPTLGTsvYIGD3X9f9JeMbyatTD+A8q4FXNLbJeUYHI1DDU2
gdvIlSjjBJz58NYB2+EmKqsh33OjHi+wmP20dYkTqnl6DkTbdZGmRp/ocxoXcaFT
98iDgc5VzTbiotPfLbBgVcLkXWFcmyH8JoLzGMC2C/rQiyacSXsJHNCrtBAVYn4E
qHn00PcDCigAxcm0UfQhyeUo3Ytf0IlSef2uaqxP65e9qzFE2BsvJxgPbpNk/Vlv
/zNW7d6DJC0pSLI2pNHv8TbkGLlKmfgzc9/OlA976n3raWuhnjG+ep6ttSISsapO
nAmbDWFe9z/EdmND8GLJZ9u9epFTWOiwa0ZkYJ8UuWpr5ZZyCTa3L1FdoCWzSdI9
xoT04ffI69L7MBUWWlgteehnKrGgYZ2d2PRkIu16nisrFqJuxADsDUsKt0yOCoM4
ELVDIgRVjBUwCQtUV10Y8l6KE68aW5gMwe7pCzVdYFmGbBG14cSSnHzAiQMXuUUO
EMH2GPvTceKs1HUNMkbGFljTNwItvAf25lwD7wRwRgdH05YhGNQrXQOvN0OUKfde
qMy7ays8EpZCdmNiwKcol7gbWPu6Kk82PIFUKC9XZeaM7Cp5DAF9PQ1nxij9t6Wk
4zlLFU2l0Z07XSKgaHyVjXifADGuAPUCp/faG7FtpoNTrY/torpZ3RcHcEoxpZmP
FIsXFUNukNiS5Duj2in8WE3BC5wHp3Af7vAOXM0Os8ReVmhSmrUNC5Jxza6DThud
0IR3Ues9/7M6vk8Bc9P13wtSF3KwyKBl7/U1yCSH9VHF4qn7C2zGwHru+FSHOfFM
trZoTzeIZQGoYjdW4jGxhxgRqHgTj2/WYknCVtvG4YHsCfHM/Zg2oqnxKVPCT1FN
T8zZghFHEsdg5nno1TGslgLot59NSgsKfi57IFtju8OSrRC2paHcHVhIIzV00gWc
tdr000WO4+k006GxALg6csGN/xleD5shRRi8AvPGBATgrZLDjKLocx1hgGrYJjRm
fdiTKYc2xb/k0oenV6XQPD70pvQg6XZAYml+3MU5BMrPHsAmXP8HQc2Ag0nr1cR0
49WsBYYzlYGfxAxDE+z3OrsGh7emRI9biZKh8ZG/xEJvaC0ox0vb2BWIGY7zOKwt
TlAsn7ODi7TG7a6tOyCbjw+VUSoWwxpyi0hPKDQM1AP071qTDkutVVs+wiPGSXd/
DLo96/wXuFsKwhEvql7uelc5rFhz9bjjU/vHTrIN64Endqk8ScwXaRzhx/vFBVPJ
hRgAeZ+LiJcq7SLpk2gTJpKxZBQIW0oUp31Fr4hYGvAj9wgg0ZFqy6L7T98Mm7SL
zs1cJHESC3Kgy+ydrKGGfOfiIQ0Kl6NBMhs1emj6jgoB9v2UY4x6Yu6rPtHiR5/j
RlhVL4B80uF4M8BEDhgj1A4MCOzMtJm1RwUV/qNnbvky1Eym3/Rn74HKHdi250xc
pYgH0g1wlkDI5dRl3Low5jlHEvnPlK4NJr2B0Ksdbmm4MMBf23zoS9RUf/JBo4K8
zhIhPRb0dDJJjj6wAD4Um0zVr5zs2aS/S8PGT8nimoh1FSZbZVn+Gsdli1K3MI59
wl1vJ9Y3UqK4wsAq+vY6pCugeI4gNNE+RqlJnpAMf3yImTLnOrJkGLo0kBW3Eb0I
f/QAXoio/Def1O1HV3SDwPVPhRkhybLwLsrT9IwbCNbJmrvilOms242spE7QLsem
cQolhWJocpY2AfTAEyz9hddeFRVOIkd7RsWJphn0dBtK6aVDcUkaQnMnExcco0dp
H5H6WNcgdX1N9ukam1sgAvd+rdWCbNJsRLpUt+mxL2o/K9Act4fYGf8sR5X8wpzv
8SOz9iR1cf9TQsmotJmmOC04oSBIUMfhVDWiCYp6SirxCrYdUeK54Wlax3/zNEHO
3+eorf6IqezqbBiYV8bUv4kYwNn7dWmzQOiTObadnmSNtwZaeyHkv6Pzt0xrGOO1
uLV0XIg3wnAL/C3y8rCA7BlEgmVFeGnPfkbmbJ7Ri3xm0F5LfIEckTqfp2x9wLyY
A3+WFn0zt9gwN8zr6cpVvdh7pXYYnA8qjtmO8DqFYINcve9XdzM7pu5ptc+b6wfv
5bDn7KpnPVPOihddkfNFg3dOthZ6ewSN1fV0s7pPTwX5aHai9V64r3hNJTT1qleA
2VjyYIyTPhh/ZhOt5wUy5zuB9khU22pB6fWNKlAG8LuOEL+/IpkJ+WefYY8BgWpe
cPD1dfKZo+bdf2oCiKtbcwUHJvR5gOxmvkAFYllgusqZpNGtGBa+jW4h4a9uWqo3
EoEYwzzYLINaGnQJeffEGhC/V1FTgqePpRE4oaKcX510oTnSj9C0TQ1yEroXa0NF
33cSFxy+7iuMd1xK0dw05+tFbLHNQwPwPr2qkpzwrqH7NICPe1DvQes3dE9iOmEK
A4urVVeHu+9ij7PA7bZTMBiwi/4U8Id1g0moA6J1bKyh2MtMBEJvuIaTiz/fkpmQ
TwkfXe0RRskK0HOWYe7YZzIfZ3N0CkPAl9XXTfKPdNpXUrKd2ZmFkB0BXCTB/hhL
3VxF8SImAAdZkaUQubBiB1UA02SjxiAowlr5IvGktc3JC+afcQRTcWrnM8uW4LZ4
e/CBd17uNwLzZc3gNMri8zWji45jVDwLBR2zPLBvCgk5arwuR668shd7jj/2pA1Z
OB9wBcrNDrRkwQOaC1tVwI607vRL8qhNzXZPI3skEaH5AetlyrZi93R1SmcTtyVS
2MLO+vm8sLCEZm9Fs8pfdWTRFWaeXugpxQTJk16I1K+/L7c14dFPR2pI4q3C/s0O
jOagzZOIufjdLtmBotxWctiQaY1L/Boo6E/nJGJIi+f2rXTXpuBIP8XgA5kfJ7qZ
ljHUMPLj5LXbH5sh1DmqXYYMK+V5s2OpBkelNzKMziu57JJYvWB0GGiTS9yCvgDf
gK/jNZs9S9o/7j81Dzj0K9pejKDnDVWpTYZBTtk3/uXwnATnqPTQ8LzA7uY1KudA
bw5fazDLooA3afJClxGnP7Nwkra5Uk3AbhxXUg+2asGEguHGQ17aDl5JSPtAMVab
uSGU4ck7VRj4GdNFMsHpLvsTzQGZp+L6zEkb0shmFevtKyRaEH3Zsl7u6LUHQ3em
pJ8bvdbl0WdOlR3oZvaKVIuy1RfxyYJk0ktBMm+Zv9tRjd9wrWyr4yfWwV2E45Dh
fPwQO7sCD04jIW1xKx0pfFrmXAWZtgM9X7u+aG02MAqtMwJXTfbF15PpHcOdmY+t
hQ99ezSkGxrB5WIvjU/QItZlVu6o7NmHQFEFksBPgUfuO3SKHM/YnBZQSCu1rq1+
em3V1VMdz8kKUUlCsPIWQfGps0+DQJJd6+RZq1iSwRt3eojfsodz+olbpshANG0A
WmeucrVKmD3QQzvIwMZkqWQjMu9kABxYKWvH6uVwIdYOIRUT+eIBimAnWPRXNB2I
pvmKS3Wx57QP7s4Cq5P2yGNVN+N+IWk4Vpk7NwG05ozoANGwqj5jCwGHnnWoMWHY
hk/LJWjW/QC2zDHCOfpuAIPuus5XL+nJ5QOOmgNe0nMkEDabDc1Wv6yLDbTp7qxn
zZKwm2iEWpiUSYwnq7k2BPhGH9pNTta8gDEj/WeRmasK3z3OxwdCh9GdnSahwVCa
jXd5v7O8vKpm/2A1iYXr+HQ+DjKetdwWpVm7+boi0PLirujwgt4Sz+eC+AY3j9RR
QJCzm+5KG+Mxc7/6kPvDwBUARn/Wr4AGdHWYO7rXi65zhbGPrIw1znufyNlMk6yP
17n3cMSJF2aE2NOAmzkdWMGRDyYtceObc20Dy8v/gc/prH8DoBA5o6tzqNZZ15Yo
6qoCSJsFWIBIgd4RnM6Br6GGLR9jaooaH3tgLpbbH1ADH+5oUfIlyOaMZ8Txxji1
SlPq6AXgG+VPMPG12Rx1xg3ZnlPZUtQGgYHcqpxyifsPgUl0Af87o7sMEgCiK/bU
6Jy/RPixFkTb9aEthnKBTZ/kSHJQBQ36E3dQbSimaRj1GfnFkUdNSbYWU3cznxxk
Q1gPYtiXeu0POZYBmEBGOCLM0+rTLySsZgMDAGsUPxI4m74tFb4aOelfezJvJX+K
g13CDj4M0vOynZg+kINJN2L3h64LmDPA+aP4rTwr0ilqVe9OsEO9JnAypipSOwrW
LN8ZXiQvhNz8pp4sqD3SnOFQcVK89M9bSu3otxqHlUr4PSsSjVcnpOsFcuaza8zw
WTz9m40ioJ3kRumj/8BDOoGm+YfEJ0oQPjlIaPYarScK1IzoAck7sHjwXOiO7ZiG
LrAKrogFtrzKN9eJqNVOxaQP2C7PL2Djqjw1Dj5LYj+q1mGs4jL2DoziXxNXe8vY
BwokVh4k2yDy1w7bqtU6q5hab6C99FEezPocyX/vthwKZuCoc+wnVOxyCPf47l3E
M8ZLTG1KNWl3Yye5M6nJvPT7muoGVh0MseSpBKw/u0IXBwf1ym9s6guiHpUN4L3n
fLAmgxmYqPWKVWOS/7mFCByPUA9/MjD4BYiHAh8E+uNFWsdrI2Wivvv/lbGO9FWI
WtKiVPf4MA8WGDj9c2fWHf4Rh8/FahHFzoiRSUxVw5bqNxzOW1swQJUMwP6k+Jmv
RZqA8B6yCCKW4NJZ54T5GotfL+AaaWIk/lepbx3EHdgC5OeaFMPNCTfTr3C7z8Wc
z+7unUzkY26BkuL9icvFx4FW8hcXdrLzASe7x36+6aN4KSPOyH8qcbYJgDIxzjUZ
gY1ghdsxrfFsxb0QDLYkWYJFtMUW2B20QmECTYNkzC6S5v+XxUuYzCzqU+TYcQij
JKii7EBCG99Ee8ZHtjfidiMNQxa85gQwfgeAqy1qe8c8NkCHAEaz3S0tdZrpPSf8
LR+E6muojqmnl2ISrOQL9W+orMISiBmV8EmH6O7OX0RupOiJ8i7PbUvgg8V35QWA
uZTt5o+foxMWEyCyrE/IZeJKHzPg1QWJmLl77I2M9z9SD7r3VuQSfcGSGpSidWJN
ah9YOz5+Qp10rDSGgRilZxQ9eesC9LYkJ5440kb2GUd56nMC0/KW0HrCJMiD599f
1KYLz6U2md42aXuRFBF2VBRC4+/u0CQ/hdgY+CmFh3qQyeY7Rxl51CuQaQwskkjv
bVNLDaX30YJ6pPXX4xaO4NIn6gKlTQkWgt7JrzM5ct69rjSeHObPDMG2sDFl6s1y
5C9TUu8JW1cmmk+ur1HxJe5izw0YzXK1EISN1/5vhLfDSv+QmAPJb2VeB97Enb29
myLu2GS78QT7wxuGqHa8Ud21ebAO2QrG84b8uHlIQWzpmMwApNRWjvrEXrvuxNuP
LFLIENz+YDydkkzom0YJkxxU+8yxm8t91EFqxri7jvNkJOlKmYVpFqTyv9GGeCzV
OpCO1qso0mVuZfuCF19uKsb/WDKbhYvbCktDBVi9SswbPnvZJNhkRV7nj7hzKoYW
WZa76+8m6I3/jOnCMbt7luIn57NUWTelyEjf3L1Ib95wfhb9onxtKwKcwW3NLhgf
FLI9xkUej03mLzhxZ9zAgOFfLFcPOX8wfIqeEXATTWTQ6vQORuVHI2KVzHp0qBwj
6/SAi/kVI4uegvaMeu3edKR7yBq2Cw6ZtFm9UKapUQnlvgL01caHtFcRjvFl4pCz
t7C3Vz2hFC9nWLE2n/dKhpqHybY07UX81zG7BMJkVom4POcs1VVvBFKrrcXUOPBZ
lc8suzoNuI7YlRWzsy4MjFWDwslVOg2CaJ/3+V69Kg0h+QVZoLJhJRc73VNnLlCK
T3eAhYR7ecHC4sYtEcqtfudPhdB6d3vw/wcLTe1kmlyC4GwlMAdR1YsUqzVupwo+
Gl2rQsiSqJMrW4zM57c6tE6Rlb5GbG+zHn3kDH+keC8HqCDhNLQxUmP3+GqYD/Bp
Y6PdmOZRtisxXe0lHXgjyXeKy2SitNqAz4dAwcFuQS+UWneaTXBzbf4WKvCugaM1
Tw97n7lEentEQFpTYO32V7qaWjwsYP/tcvQfLZ6P/cOEM3dUQXjFq0+Mwol0tS8p
WbQJN5zqP6tmraheuqT64B8ZTpcmyIhoxg6dYTf1O2g2Gby25/+bwoeOt+iKzJCR
L31stcP7N6YEE33GuY+aJdvfPQlWSjUF0RX/AHi8DHmj26cv6j6G0txBNXPuMdqZ
sbStzUNNArmJBwjyVpdUF9vRxI1v9VYKejQIjoaUHtL83okRrHCdojMmliRdh4bB
ILXqwRJJO2PjyCATVdc5PFrmZoQHpS0DUlaaqmV53lqrhwkE9z5j3CJFewQkE6ro
4pdwl8auMqYtxUW6UfUcTkN7WF6/npWJHLUPtjDR3eEYxbI8WkUcmxT3wEYpv1wp
c0WRigg9vhfY+e0AmEsVOQdULrOjt+kCdFTOXjbDU8QyALD1ZdWI7NgoPI6jbalN
xhYcpKNj84i76+W4/kVeS0mcyGcXGCdzfllJTjpnOlYlTNMQiSjA/AkJXVBlrg6H
hRxRv5CrFfBp6eMy8dH5TQ/g4qLg6QX/sZU6S2MTjRyc8xHcNu9Y97H7rfDhI6JM
z/rnT5xLpe1powO2iA3+lwCek6ksEla3uWJlnN+tNdjVFdZjP/jzD5Gsw5D1io0A
CKm9ANZH98GjKK4wXLCUiYHsTzGTkZmfgnxy+RBrmmmGaaNgllk6QUlKIOmuJl1T
D5TGRFIp/kKaRTZPC6bNbSKZY3SrP2+HlWDbO5IP5mGBfOriX3zeZrmh2PYiSZvz
eYfqII0pvGZ8hwbkEvpowW7JlCnjs7RfuZ5PW/IRzVIF6KLzI6L1Q7tuiHOrm13F
DOoM7Z/RZASQC3u+eR6KdSRpYGzYOO0uNW3j5CdFAzwfs0j8Z3uAYyllmOOBcz6t
H103B4JqrIxF/mex37o8KNPKOhjci0b2NRTG7wz1pnzUDsEhgX4ZqQ1bebQSuJRL
ApV0uPccajE8UU9L7kfMhWSvqt8fd+iPDTpfA+EeoN6ecRm1h7T8Q8F9Lp4vQPNo
Hi4AB+PrAdpP+uaVlwPjz/Lga2mAFfJPkS3sNiPv0LQx8SxMIEklIKaUD67UoIPG
wSkUDWZvZIw6EJCOrEA3l6TT2Xi5GywYn+CknR4aZrc9EQmq924Tp7yDok+3Oe3B
QHUpgKvZLHeuS8SzdjfRu6WRmp6RNipkPpaVUNKMtS5OC2L79fMTnMwMS+AcQDZV
RFP+5ZeFc2zAAZxuhM5Zxfd8j8Glt6yj1/QsySzwKOBKGWryqhWuT7WNQpHDVSh4
vpmF3f4Oi48l/zo9iyAzyFJ+GUqWjcCSWbaCDyb/luTA2EYC8w3Aqi0iY6g24P8S
+XMeJoWwuIiA2t1VV6qGU2GWzVR5Dosqixfc84BfEGMxDM3e6Ieq7VvAVJIIg6s6
z00sc2QRgonTQczczsjg873FlDkhKj6bNfD+iUi3HatTez9JmCYpAaolcl6fepx9
YY4rFArT4pHXG+nvu2BZUwYy18YTzIlrRzt/lpIMMzBeY7VHzujITwAbX9elsfh/
cvCE/dQwVadCswsZ1Yoa927/rC2irYpBi9ytxjm4Bk8RRrue2YnyKSAITxVrjzux
6DdPCZI6Zbezj+3oi4EUmgM3PVhG8YXQdOJS1lwUmHOi6rDc3m9z7YV/VS0icyMS
81/7beYSs//xhwKpaBRWCzEni7BPeBSVa4NsiAcV6LvosD+uiPs9eWFSIeJOdBXx
jv17+5O0vcAleJz0r+hOg3DCGjn4tlwKTnapqltk13lHxkVq50BwX2OisWTfgoHg
VPvaZHizpfRoa6i427LEJorzdb6u2VB1ZJ9NdJRzSBeMLCiCc3cs82eiMZBm3fcn
eYviBs06zHpdjl1kt1/+O3FYxLjltlSZKDqJ3jWDTapohyoIPBtAZnCRRQ1p1qcm
vVk17Paz9fiZUyakBia3VP57FXSD9AC2Pqq1vtYgDWoCZE1QHh269uQ8zDmzXhcK
PD4kCY40YY9gwIbCGsALmsQmSKP+6pJEZYriolyw7cIoAHV+7ZXxLIIjnQAvb/yH
5zuWEUSMEZAkw+IEtbQkAMFONl8ZtOc92T+8+IiaRq/KM0KXC0JeWtpPXwPW6B5D
EvRhYJ23MX6cFAfQb8CmhnE8uOOkyozWqQHrnqDY2q3//kAQ9hXpWfjWLE5vRbCH
xiFOuI+T46TBcvqI8WqecWPS96xfny+hzwFDpvSl/M7pU8P+ZsGAwnw33kqICbno
oyDJIyCEMD94Sb9+IpbJV3hwcqX1Z4PfDLMGYWriXn2xPigse0r3qbBvSCxq291D
qCmEWENLtkVyxZt/mCCBtc+/dPNHb1rtsklwfcsbqkHSNYidc7KxAIzTrdEAuMOL
1iVdnptmffN/mFLgOK4/Pxx/UBMDl+LMIaYo1KIG4CS/3vCR9PJAQ9uHFcV+9EoL
D0J7aCK00mPkLS9oHCKW4LFM/E/oqeRZWpPW6lxd3yUMOSa43w7rUTkx3L8XHg3L
X2ipARRgxHYSPtE/Qn3Zv02RHO2dEM2UxnqbPYAJGdTyVu6Gz+HBd8C7QlpuTt50
cpCY9PZErfEgmeu2XRRexfLy9zgfNEWa4dYXnZxSHT0qNXETsO6NxTl6KuuWl7cU
DP/xT1cSn0mm4sKbLLJnIqJ4drWkvIMKSaoyMyX0HbYXP4LN5Fb5r/y5aq/mG0r6
ivi8K16MsBh5XjYbqH+JLFYb/cqI3ANmohHKxCHlf10aIla5nWEzzvKCXlO/Hguk
c4jg52VEZ0HB9jIOaijby6YWrNy4zyqjqk4kQJCC0C24LCvx+Z1PJQeVhbV7dII9
IaiTKWv9KCiaWKBK1bvUPXiWGlY4ijvhh+gff0mkdiwQgyANXOD7xkQf+OZO8DbP
BflP0EYf+iRrSNH8blR8CSi/8TOLOehIUK4jd3ZY2j5MHVvgQ5HweahMkV/50oKz
6NNYHcXT5JvfHak6kKIt8MKTJ7uOjeZ255THvpKePZzOoZxVCu8T968AdaRlOL0q
4erMEfuLXCwp5GkbY/SgrwnzRx841xHAvUT1n+gnnLoIIMf5H2iV2bg6aE9iKwkf
0Fg7NavG1btuaTE39M+cNqI9k2uElRQyefEVtiKdDzRRZFW9nA2Q6mXgojddqIux
nSxR2RWSi6fED9GPb4bYbbFEyCbHAyJTd79aUXEi5QiU8K0GnbXaSI4WjsxyLA87
tP7Q5OZKUJejE14TuH8aB8VGgBs+mCh87l0zSwyzxRc5b6/mUmoCzey6uSW2veGG
+TgNYBju0M6+MqXA0npcHyHWY0NXEXDGawHWLIYfylXvdCD+z0AVMmJ5NUQHfxpN
n1xHQYrOfxffR6cwGCvcNK/OJF3fnV2z6II84GXK/R5pIdr5epAGKpbTpDhzlpJw
JJFtTd0K757M6UQwWXpkhqTtDgR3zLa4tzdQD54Qpr0Cq6uT1eAafgKa7+JiLRRQ
JPS92hmkGp4E9NyaNhYB9ENDObENUVAoIX49FulNlVY8sCFJYViHpekARphKZlgS
klezhHbYGBldoPXI/wOYR0ZQ0Ig1YYx0K9F7ji96PwtzvU2QXN77c/ZhBbVyg60I
BfKmB6RTOHSrgHr9GMpAZyV1YDnmgJrpsj4CRqmXwMrs4rCOIGqAZnOHEF5Mzr2g
iuRQN0jZea1LXOw6j1GfLZQZhpE7RocTwIJSONYL5f41swapzogqKGCUHVSbZg/8
J2ABOLosHtf7bWgt0ErTimJSdFQb6QILvQiGLTxMTZbLk8US8xfTmvrTDTFN9WpZ
nNEyPQiTjvjY1Rti8dcegIYS9QpHGbSSZF2omYhCApvkEVT/2K+N8ZkB5RDWCZTW
XKXlC1KgS39FszIfU5h5m4Ha37sr+hb064BTTrBmn+oIDiYvsIVlyk4EE18xmsZB
5JgF1zXAC3DhLRLvl7JTgoCEMKsaBgjZjX0k13W4HwVRH52fnMEUnM60N2XzTH+C
ItVELtccjgR2y+4zBDDnTawE79p4x/GjYdeC0x66bS4IUuOzUt658W0UEKnDzl8P
G6q6zlG9TqAh9q2pQEDBsXHtAqVnyqog8coNJME4GXEaf9pb8EyNcuUQjF4gKaFP
9jETVR5iSqatXWruvUHvkUI3S0U9oLPQDEw3REwrQajyCULosNMa0ifcWZjj2Nmh
eHfnTpML9rr3MTCKcIWFrVfTBQrB7VGK2ZyLACBxtv7ajvbvJDi4e2fSQVxma5fu
hGwBVzF2XNz4u+3RpwuQMhCNIRvGGFppdctbzAfGGIzAJi5QvRXFzcBEq4w/wYe1
fjelj8JpbYpcrXitAyxmeXQi1g039TLMNIdKw+IfqJUbk7oOdBHJogB9zVqayadT
NuuirD4RquqWJaHJIcUunJ+PkO+ZeYfyJaARz2b3WZVlanXhoqTGVswjX/dNeeAj
FAWtRmSGUyJS4ACA+oYEtIovzLGYlGwttKX3DzKwxr0h/gUjlSVqwqKoU9yU8m2T
ntOCI1Fcv4QxahL63fm2DrrPgL264DDopH88Fd+LNDgOAWX6+oWQp+WFr+/rKiP8
9xg/SAEAen5xjzpgEa2HT7FhOk/V9UPMdKvqtdQbRedVg0cGuhWBMepUkPOjy5BZ
orWw4wDoi1Kb7fWuJg8ueaUZuuiEpSPyiX5m8vQl2rcQvZSZ72KbWFwx83RISddp
MEpAEAdBzKxFdp0uTSeFnc6m7+AROizBrQC4DxBYwcEwIYAaV8w0K8SFGVvga76Z
WWpRw4NnLl840UGA54T25Tce6yHslpzlDVfy9XsgRqHVM9GqFm7Q0qkndW95eyJB
JG8+QSceC6sHNXGpnWUMAVkdw/x+i4g753ACeuJGK+HvpMAaWDmsTZ1j0PiYFo+X
YWZ53dfI4PnHz3aZWAllWmBE4JFImPwPHIDQAZ5QQxndtk1OLqrTJ2ao2CseStMm
wLR58JFgkHxOLOf25+c8dPlBS9+dwX0MCnEmw3m+SXNMbwZ89saxsThtyUyzEdwF
n8Iy5pC/rIje4y+0YguvdITEnv7vNr8Zn3r/tQS5T7MrTw0DP4OemURDR2Aw3jYL
hr0BoLAZkSVVpIfe9ZMlipydeFWWoW1K7tw+2TeS6IHkOcU4wzAVOKFtoS9ISQQp
41CTgFNC6cfCxErjSWsgihL5fbYBACBDCprijtmsS2MPlLzWC9JaunHPU3PW/vgM
MffpN07uGzfbtD3+9UYt9seRtQoUd7UYoavkDnSAueNhKdfDZ51oeHtIpkGk0DJs
Wr5/dqssmC/gicBb6qY1TfWvTbjsT7+eMq/MRdSkbqffVXE7jsw9VtCt3HYz6kLH
tzsJhTtk+qUZPwlrKlt6sXeMx1lT0bEpa7aJBOtt4pzNCHkmB/2EFatSdMSKsofN
QmyBzsLppeTL6JMkypVlIoNYb77LC1CLwX+A7wiQdq+MxsBWPfPotSOvkqFPyPkF
46f8e+B7UTacIfUf5c09wdjf4U7AozPJJz67zWhreeZd5ty8Tgw1DZDdaPEDhu0U
BU2qm4EFKpO8O47QTO1blzReZap1sZ/6GK7CI9HwcuWpU27ecOSDmDPW0nq20c6M
cEK/0S9pWTCcXDNfhFZOHKm/Rk54PYO8p7ZH0KbmstdGuwNGMlZA6+G/ja9EKZE9
P/QjHco7Q67xNoeLY+JL/PKsNBBGQE2noDusRknh3CaHOAG+N1+wKoWZdt6IcHmX
c0fPngZj0mhYquhu1f+xc5onu40Kjdsg8OeM2oAuv+ROAOVqrJeeirDQjxnUxm6+
psqXSgONwsT0AZx9T2VQRbuYNvLFf/vGypzJO7QzzeMzDHkLB57llo5LMhO79JeN
jsNwn5wgA96ihzgZlMdQaG0uOb4qEpSA2qnm9ED2A4NSRj/Pp9IKR5t4dcS9qdA1
Yy4WAEJce8cXHNuaj52Zq9UCfY197bCTdPu0rjV3g+AcLbzhUx9W8u0BvpMbPTr0
T8Q2Aj2mI+51W68J5Tmhpo3rh6ckO9Y+BFlbO+C3zO/+QFvNOCMTP+XIlRdHRc4u
i4yFuXMY7fuCrdFejdYIbwSDYvAPU2T5ckrp4KclkIIQkTKlTxRvSQ2T8wUebmD3
rrPhhEi7ygmvsjSEFOTA7cjTzNMDm0f4KmJBdzwe2z2oHHBdug1LSQXJItGEGoh7
2FI/5QO6CtXSP/0EXDYjXexqPwzeHrFvecy/Af0fdyGwWRmvKxzEudzYJdm7XBzT
R84uih8b1DwloTlCYdXpq/e8NwhcDqRkBdPgzSiIMqejV6/kpjL/zL5lhB/vYF21
6aFEHx2DeGPJyuT2OxnEefnaxTR+JynAwYYGDfnT3EiORmmy29M86Ni9aMVKJ12a
af3BDx6FkLbIDvmp15yxY6JirwFW58nF2E/G6nXcklZ4p5/vBLZqplVYHaeFu6bH
hQXId/hD8zdYUp38bn47pbtLi/0J88BDCA9W+LC+J90ERZSXA2su4oiJ+WUrWUvK
l9AnwRd6V3Asg+9YndO96ZhB+e1hLJBy55h3qvpf9Tbkpse2BT3mSMAxGlbRuhVL
j+6q3tNvyM1pSNHrjienrkJHax+BwFc0ZUQF381W9uLgPSciVs/k6DdWEq89fNIS
WLm0Z2J2p4aFitCPJc79Gx0NJjEOQXwd0wX1w1tKCuxyY3W3n+4ErNlVAikbxGxT
NxuVgRNv3Wj/2riEPUxsFuGpfR2NpnRr2ZOAQ1RTNJexLKbQ5T7sbqFXfFbdK1vE
O8Bcy8CjqVOB2tq50SgDWOfIxralic3BQvs0xFv/c3nNQgzuLg8wXzyXucnq1yih
v9am3EcgpjzLzMBBUuSXdQpEInXxHQJ82r0fzl0754gJAfRvt0Cu3HNsk60zaiMX
rP29Yem6mY+ioqJYyX5MsQietGtS3FHOE2LsKaOXIh62gay3l8szDP43LWiDaHgb
Z82XfkKI70f8DC763XzMq7Liuz1zVwIN8D0uF08MjAwc/kA+dmLq/JSxyLjQIr2j
7cmgT64obQPH70hHF8XFFHh1PFIn93lA/rlKoAWN8QM70+INJLSkPo6g2Ar15CIw
OcMAWRpyUeuYINpi1pHbFVt/oD0PZUT3SmD1rKmC0KGA14tx7ji8Q2uLKbj2vPF5
WJ2AioXc4W8Z0UouY3aoGe2Ac2vBQ4Qwd3+nv8R28UVhg5npLzRN+WOXKSSR/Y73
mhe3yWjJzFUdb0GLaxJf7MKerSYISKvti1l037Lwi/2wfb7v0mvE6dAzOLlZwcMa
WcX555N9EhL3CVVaAVm8e7+4mkoXmDJFkD+Q7IbTZRpUWQEXxEBiQQf23Z1kUnUm
AerY83+gV3ETTSVXzdtxAuaYOsFVZZtatuAG91fhLgMWjQVqD0cbAWdRpHJW2V6H
3t0+rqoqK/3z02MYZiMi+OIvNRvO6jooszECA3tQUVj6sZfS9GrOLIpcXlDos2ig
cxBL+nWv8XZgbum6y8vXt1DNfyVUVrI0IvS22zJnyP3k+M+0sOJ0VzvdYUg2YpCX
Zu6nPbMFQ2iFGR3lI3anYjxka+Iw5V68hY67iRAZdtY+xU1eBrFnBoe3W6FstFWj
SkiwfHzMYzifUd2CovVOg6Oj4u8woXzvBECpANDJY6Kkdq8i7qVVf3ETeChJewzj
SypyschPZ1eQzSt5GMmWZ3f1q2rdFlhkhfKCk1iFhIc4F0VCVsGl9yInZLwHPoyU
Z3538QCCCUm0iyg3lgMaawVN9trD2hpsUK1hlwRG+ujDEodaaRQQEgC8B79BeJmk
S0WqhBu6nBId3J149eAtkPT3g2sgQ+BQI7TNwciHZtME0+Cuodpgzc8ALabrlF2s
GyPxI6lQEnwKSY1cE/OfxCwukmMLxN+9xgyjyOWrr4eVdAT0w4gt0IBaMC8Bmya8
V26OvGnAaOPLeyGb6D6cusZaJm2iJcdAEcSSZD4haZsT4TxAp52dlnYOh6E8q4Zu
gVpHWZbkabQPprw2yC1WcgZmBYeH72c3qSnoWGm8SY/AL7PwuIefDXyVzMYRJbMx
v4v0HsfKUeDBEcPpa+vVwChqkfKz8PFqy/PvQC/Or1tI9zuMbFvjbrOjWC2pD/z6
wfXJDCrDGqfkWvARqLZWjQZvmWiA+Lep1UWL7EwwlPYGYy4RgH74ZxA9qfP8XgUf
XPnubhAvm2r3qUj7GYW3Pq2LYlEgO5IkW5yhTLzks9fpVlYtPpqcnt3/WEP0pTjv
VMIedkh92VEz8QHbDOCdlGzifoXmVclRln4OkSOjRU5ArbwJsjymmTvus/AaOI7q
OGE5qoT+NG8eWNcQnOdm+FHsz8rndj3QmaQ28AdkIEzpI5r5E/2Vn2RSt+wAIU5j
XNcCjI4kcqyJ7g+OCfkch2lwdP+LKEjVVZsBdqYpHDriZ2xAVHnHEZtsoO9qI9hL
xydbAh1qBaJyUarA2nS1Aqy1lAXgVRD1ZJtXUN0727+2bTVoWQUUtvOok8+asgnd
wl/Wii4cjSat+Mjhd+/AqtW14JzOO7xvUwpYMpIZ9nz9RYH5z8feuJMN/ClxwKpL
Onz2YrbZe4I7aDw2LgDx0CWMLZvoULE+OTJoql01SKtK4zpgWfK7+5bNsJqI4qod
PT/009aMoWzkHLMwRIT0QLZaCXjtVEP76kpYCBMbzrS91jw0uKjiu73sks87gBKz
qIv3tbVvtLazEDPo9xh/vgWiQcetNiyIAEQXpdbqlWx++e0TuLo5CuqHO/dph95t
zYzdRmBoWDSMdxr6udP6dfkxRTcgQr84WoD1a4/tyIR0qVAT+TXtfJLt/9543G9Y
0VASoPu/0iVViTQK4Me4HpQQ1N6tAXHoGzXpLeZmK5qCFnKUsjvM3DEy8OeXcJmh
8bJPCbu2UBASWP2bdHInmJNZxfvTQjOTgICHfpW/3+Wb7LEgQ1CGQJyMRRgXbZ9w
EGRx3UO+3+P1RcF9VGtRKIGRVSuh6H6XPGwjpVhGlbn/6NqzUqn+jDoN3KmO2AQO
5k/22eiLebm/LStk13jzvuxUxt+MHthCuChz3l7daKGCSpqFl4yRwGZRMGS3mfRR
F12OI4viEs+byUUjhKUch7Jv2XuJrU7AGfxcplqrEkbtRgjY6mr5n0Ym+iG0wccw
1DBC8XqzRIz+rB+LEyCAEPOaABJmLJN0inSLxMf0nHHfu+cx3J7+1bwVLyzG7T7U
CiTpg3LIYltwqGun2JjPZTzHURRTvEB+n2zmNHryuP5EUOsDBDBIeS/2wFGATHrm
b3P9rICeeX2sXo6IyuIxPsgiTtl0a2IKN3l6hRCV/Hv9Y6Z/cyarwf90xfcit+Mh
LCY5fzl887m+fO4jKhhOf7wtvcb2A7O6YHoVcOrAwKxz4t8lvfYUm1J87Mg7Vxa/
hRFhVYOTfSTZJ9smIR4LspUAWct/oiYbzM4s5WroQ64T4Vz0ItwMszFXwuNPKSUn
o9vi/hhGWChrcBuCavKmNyHXXWPnxT4HJ/l4c+7jL8ivGeQ2C6cvTzS2mF5XOHvA
IqT7CYqp/XR0Fi9AEWtTy1PznkQ+GPxs/LUdfJEQs2tGzsx3nzLH7rA7Ru0Da6eD
0oYJMhPuUHDtOVs8sWu8TAjhEFjHa7qplac/QVPXHgyzm+Y8xclkVuiH7S3GxMji
4Du6egxmEiEX0Bqct+MFuA11XiQu0ik+a9/AhTHRlcOg3Hn1dGF8J0NxzIOakTiN
wHQqy9HipoCRKH5/ZUE4ccdVbEZ1Z0hW8t7oXM0/xI2FMPgScnXmU6Zr0JFOgWv/
seAIPT8Ou/ZUu19DDoKb+/nBzpASRYNN9Ktc5TdIrANlVFxHr/lo/T+Vx2szsfR4
r2K0W2h0DZEfFSpF8S3vwOWsjcv83gVa8XnN0CN768doWnRHKxaihO+/6U1VUxBO
N5KvasnfKmTdrpSW8smp7PjOBUPHUGLI3DkBzxvwh708s+I6StEDrbr+RtUBD+R8
zUQADd3bfV1a7+lTM+DyXx2K1z5Ou+VSHNIKp8vYAoYT8WFAB/A3/PZ9ScQt6H8H
AX3I54q+oykV6+Oxt6Ay0BFSi+oaLKR08SH1iFKTSTPTaaed3OlHIqF51a/VAUiZ
zZ/Xz84VmbOLysMCgi/c6aR82k3Gcta0ZUy/5xnUINjGiueZKzEvo7nqInhj3IqX
KeTY08gjj1cZ5c/KTTWtmoqQyL21NMY8QthWQKv+Gj0lcQ/z0JE4FdzJsFRF2T0i
wGKW5/KV5Xd/PFUbC5/Tqqw3nYms3Kz5aBUPZRJa7gg/9n2v8vQLNI0hYYIFex2O
aNtb5PaPJ565/aD5zsP9Tp7LgA94D8+o8CkxpwTPlLjzgrdE7bRoyVymC2fpKJJ4
ARjlqLb8IZPt34SDvpXSMY3qyIEyd+yEzcOpDyz4KVSCiYaJ0cshxAvPGxBkrAjl
My11NxO58xXhjBh814c3tmeJAkovfZpVJO800rwKHIkRLg2CtxILvh/VWtdyYcNQ
XAxz/azxxl34P+zjJC8Pc8TSUEoIBw1Qg0bzkWSSUt3YfkfINXKfV8VgRYuREvRk
AXX4ccGIS89hiDuQDGacUlTVYXPMVtGyN9A8ZyUnWWMcceQW8mo/udZnqN5Zj9fu
m3k8umoGY0NZV0+oYZwZAKZ+3fksDNbK2PXl8CRKoRJgtihgimC6Lal2Et8kbwHW
1QoNbhPl0VvoNyT07E/UrjCHhH+hbmyMed7HEbdbj0XCGcHHfmW2n1f57jHUmRMg
yLb/a9jqWVAfjHkTKwA/5NFgcITQSNzz66om6h3e0Lu1GNdE6S8dTCgVGna6iCuE
CSED4Hwz8MkGNi6+if7LHzcbxDr6R5hA+1bdMBGLUuntDDtJ97Bo+V33k/nrArsR
hUUX4ui/Wf0y4dh9QbF/3SkUnU9ugy17UtlFEVEbrMT0JE2cpAapDDH8k+l6NNjP
zRbGkyxqCf/xOW4tkuo7m1XXByYBA+L9pLx28lWnVEKhVxUtOAzK5GppI0yG7wo+
0dZHlICNUdMx9dvYuiZaczLXKfKIhjfH9O9vomZ8zCV5/SSlAqoUb9LIkG5RGOS1
Q5ncJj10WKvRQmRfkmO7OmV1jHqx6Zyu8KtZSurzWyRyecMMsVvqPTjne/CW4luY
L5eYvkQk/1QvmMcWqHlm5G2v28zed6DYZ+DMBDyjBUzh5bm8tvhqFUu4uZuZFTJE
Wh//zPYrwRroKDNZhFIlQHokt7fQn5JOJfG9kMMRirCtuQXX7QdMZIhHjoj1vXfP
SxUEfV49eoM5hxZmlGv+m7ZEdeH2MMfZWt/T4Xqr4xSCxqGpy/6nOhXo6p58+aEH
wsLhBAqa4+H+8CnI5Vc0MWrGdIPByGQcXD1tZZ/W1T+ZU/9n+wMYoHT1FwdKZlEZ
vLZ5vQfpQzIN/UYPeq17kbzhAn90GQK14qoat5qfiXTcyW28YhQ0OpLuakKG7dlE
G/tyuvMO+pH75Yr7eonlkFND5i797yfXTP52aRTgb6wPQKd27rmRg/wXXZMkkPmV
coDDYQoMmeFd3U3JhuSZr/7umq2RxYCWZIqgK9TIEhiYHyAG9idDLTfZjl1tRli8
H5LZmZiuXSrwJIwp4jJnyoPEtWnJfyX+JoGV3AoKO4Qy3JbODMnLEHcz/jkWhh9x
ORPmynoBrZsDj4LHBMF0AVWA0ZaHe9Zj7CqTs4ENmFtwvckQEsaY59iwwbHqd5ZG
t1IiUGdVSdvjFradygv0cR9sX+Xy1KhLVXcbkYkHH00KN8ADf8f1WddO/8PU6tN9
y+rtlVMAtO66r+NOBCrxYQrylaqUaxvDNz6G4rZq3rjuhtrkYYjtu9cGQ4BSs1xl
7NXPwhApXzQyYvr6vgy+Dn0bI7Y6yJzhyzbXCPy38626WXvv7KRDx0Ue+neMZ968
N+cZSc5i9MBeuZGwJZj1iMSAcoVmFU6/9Xv01r0lkY4whjuu15W1uME4NpfXNHWh
buqhCjNKFjG40BATNwXhBi/KVZwf8Spjq6BwbBXN5Un6UF0zgAuLAAayPQ3JHKRs
X3gKM37W3oHKEGIFgVk5Rb55FSKIYhBHGP/xpwLoIFzjQF3R1M2wwS3UVt/QQEFI
ASmUKbrdGwVwBc+4aVOlEBQPBpnQqhQQiX19r/sPAqna0wfRt0URPrLMjb5Lifoo
we7qsQEDoGbrN7n2AyaErHsq6Y6uiBTM04mcNQ7WQzdkjAmgMG1h4NLDVEESSszn
hrq+uEZA6/O6KOW5+hLryz+uT/ZpiZsK6b4hDXFgTcl1ogm+oX00hrPlAtNosNZJ
QzTGJ5nfVDXcHxJiOssQ5dohu0DKyae03L/fx8XrpE/NSYTSZMJLQQnUvUOXdFE3
P1Ju1lVNp4gVhUOWJMhQq4en7CEfVH5yGKRQekcBMRf/tWZnlMRsf/cjGz3LgyP/
E1az8grCM1uAwY3qCrkPmmCRjXlfZD2nKt8uPoJBT/+fMgcvU60LU3K/tIqqHLHQ
pdiUPITGZmLgAqPpfGoU1CclOXLDLj+ftaGfe5uWpyfTg6cmiq+QQLVrJRx86AGm
2UPaaevRJoQViworgYnmG2aT5R0CD1ESyCRUBsDANbPPCXZWZ4M+wQbCH13AmlcX
hrRLWYmMAU3Ml6ICOfcu16kX/nfDYMg3+rjVXi36YtpBwtF0+O0Xi0Axt/p1qWx0
PNqpzTDGpxO/CCnr7nV7inuVzQtCgaqKHfScfXHts45RKC5hlkcA5I4Cbyf3VEOW
CeaDaJbm2p4O9shcMoAXwjPqyESElziDgY8769g8aAWMd4hiWlBpvWUhKT0CYxGl
Yaq6ztMl5kZhhBYndWzTlmaR6sj3HdrUK16eRycx4n/21zwRdYJou083cY24DfCD
I25P8f56DFEf6Zzjc8zO+Fq8KULTpHbAP4Ct54lB6DHUO6FBmBgYrMwX5wiWc5Ef
r4WwMvjh/hJ8/r1DYFO9NC+a822HCMldw5q2zwxR9AHemeg4KWXxmQ5JVIv0ceeW
ZGgIExym17uo/EpRL8KryNkdvws0qZ5CqhGfNy5NPLYgf427LUd8QP9sibYV2kIi
+ujRDCrrBtAc1Ym78GKHqoFBQHmvTGn0aJt/+ndR+AYi3MDXlXaHnydvoMcuTere
xPCm47kUIe6QSGmFdvVcaWJGT6oNHSRyga2sua0DMxQs2l0xXx/OEqwbHHQAQuJP
P/7QvnBDlLyn/6h2g1X1QnHZGkpPunLFgeWgK5vnI2ENMiCGdFbZki4eY6ctmrgC
3sZKKI8oojiZhGytex/++Q27a03PDpWbbqFEx6j2jadC8Rm8ngk8eVvCfIhwaaFp
uyL/93KLwuBI8dn1DybaIC67mj/vyh/2CL1gWVo+rpviAOuPVDANRmb8EN8mQcBQ
0Jsz58fSg5sHANVhI4zqUuiCA/qHwM7hWWZBCWnzD5kZr4tOtWwuIaEDQWEgSukU
5uQJYIJBSIapMOoTsbIXHNP+ms7/KY/X9AZlYJkGtzd8liQbmZ9KIZI/5KUvDknn
jjqsmaKyX26473lXTMPixhL19LP0e7NpVsYfd/jlVCTAxnCNlPreMp/eLgncBSXW
B0Qe/wUKxJdG0QaZyFCbPs3w6h4YCeLSTEWMnoLsFIPU2AC/FsslPDOCyOWxvhRb
AS9ij3NOiXtAqj6hr3RsNHOQ4g8iCYLE99rawKu9PZ66kV36agbyUJdvfngMntnB
hzTLHHSF76kzHboaItI8rod/YZ8J6rcRs+W6xEEamLn/nwcd4b4OfkH6WwvkryiD
esCyDW81BX7jvRLC1tJCigfnPCmJ9XYDg3BMGNYT/dR4adP9QP1azcW9dPIOnOWq
NouQwHAodSdbehph+Dn+u2ecDStqCgg76IhSvzY9IHspYLWXT9lPgksglgjBUxSF
gj6F7y/DjEcVgoWB1SBNsVS4Mg28rMVifPRu1LrTfndJoAKJeTAjsDFQMBrY1BdX
ly27QI39737FCntorvwqEDuO0V7gtuubs3n4Z6sf0qNBvRy5SggvfuM4lg9ek3uR
ksp/kg9fH1u8Xxphv09wo65AbPPd66Xrp1u09ptyel339DghhfDwOA5htJJq3nfk
SUC1JtaqHaDp+l3SLJ9mIvD1+LA6rwK90h9LkVFixmNzscXxeT9ymvgEBB1akOYG
V0rNvUxX2kXmzG81/w/VMewEyT6YHaNvl2isewM9DOvGzUmmMQ9jIHj3H//icJ3L
ibnbnN7ov6BtXkRm2dq8UzSImBtGxgg5uAi19AFPoHSHeOUlbFeqYtSOeijmJOGw
ix619QiWRw1r3+cLOSGWiphRH9q63dlcKU9VP90aruki0GoKLU8KA63igd8Qi44p
VEemuurW2b/4fyEvaVlu3H3JKe41d0xjubIU3E3zbQEjbvGIf9IMCP4rYxIRQuuj
TLdjq3UZrt41fhwXqxSilB3gF7y7NihWJnj2E224BUXfdeeP5Xh+RzLM9f0k2bki
FIIhHPPUvlj8gJHwQ8u3qJApbl4RLvBEG/UyHgNXg5pbq4EFm+Phajapenbfmcgq
JCBjtR2VXAfScZVbA+PbP6S9nkZHL5V/zb+cQukqqWZtYCHO+YeKXCp1YPbwTSOc
QBuAQsMGFv8wZFYbcd1jIYoRRAQmQpaPF6YDEhBusfiLUbuWBtwfIwVwLBWiiM6V
Auakup9l+ahslypgEITqkVw+fbsdpMrvwasXrAJdGcTMFE1k03AfDzSLqNhvqLJq
j1haUmASGV1R0umSJ18R5fKM+JMoqXXex+eA1XBCC0hjXVtsrLUK/hKOHezkFxBv
JWz9VEaJye7spwg7EsV4KOxQ6qTBhF1HMXHLv5WY/qK9aoc5nfXlLrBBPE+jnXRo
aoLCVZ/yi9RkkPCg8aRFybleas5rWBI8ea+IzniTGDev+Fa72hYdZC53VXK2deVv
LT+SfVzdYi47xXVRyI5WNKQfe/uXaZ8jy1qhDjwmYrawj5DNUgXjEb1KAGkk8W/O
xg9Qs8ixMqM3jnpgkkUeMH0bvA2JbWOa3ykIaQaFeNe4BzoBgWKPu0R+TyPxyjuQ
OXgcEXNJnf28v/qnU0jW53gIJGH5YmImVnA8O02XGwK4CWrYyPMtdlBah1WylyGe
5Y2U3Y2co3dndbZXX7+/xDdAmbKxVkVIkd9aPhMgjwsybA1YsUGwcvbg8hORw6UO
HRN4GlFsopkRwOlIZF8vhwRIrEWMx1mT9j6b/qAOiPyB+vQmS++SvBmu19fN9DYu
ldHEZsPwEEizvOy0qwfV5NA63M7qeNe9pFD5aHtjYUr50InimOIfaas5c/NBh4Ak
fG/juSvGo8LFbuy+2u5o/nAAaeuq/LfnfCP1lzIdHqK6ZheXFRks7c5642YPJzTy
QYR7ubJNvmEC1oa7PMd5bZ+JoeetAo38mwzRoJ4I87BKNKcaVd0BiB1gl950h1o3
b18MiQamSbEuhJa575mw5HMk7GKue9hZXAlk3vECarGTXD6HkQMhQIAQQLeJ6s9a
t2I+kD3xZlnZtN4VuSKbCt1i6sjXcfLjZGGTUncf/n6h7ailCYWfKqGJ4aHg3mSw
u4PuYG8sio7b6tLVMCzMFfWKQdj1glj5TOKKbf541xkcgFEZ5UQYTMNdjp1fbOfW
wTE31BTBETHEEfgwecBdS4pRG6e8uWvg1tepn2UtuY3YIUb/ZN20dEhTLkrWvWBk
GKLMpAX7nMrIi7SBdG4HeaZdU8F56I8X0D3f0CbPq+EBOTH0UZHJUrXOXN/iUZWU
vk9qpXNIeMA4o3MSDeAfMzqz9jFW3lokBVILa5buEswR/8ZyvYP+tmNyszaTYxEA
/5IQAdTsSgft23U4ZSO/r7jV0QRMkte45jMhrp7G6D73F8CLfpfNdlx9ercfBQNR
52HyIg6h2YzhSzPCBrcqjthunFbfT/QEwMH3XFYIqNJf7hA76emVdjqPBiCHrcfN
b1JGonFxAZ7+bAu9GlUbvm4TsOJqwKr64qzDtxnFuwIwCkygyso0wT3L9K8tbJMm
99hffZ5rsC8f1A6FMK6My5EmDihE9QPBpGseasVFbzL5ul7SqfYvFHpSEYd42+rp
HKJTkUCEhn39fclvbl1gG4QwSfG6zjjlF56fNI6j2MW9UHpg4pICB3CZKyBn/UhD
qZks0haclqEFnrmRGA6Xw4BdiCQl/UmdbB9ltAwuZzc/33kT78iQEyIgGOk0sL3h
Rn/Apo4bhpvY3G39tjht7C2MvtEXiSjozUM0uDiFfMRWs3qCkZK8KOuxFyOEe+TS
yMoqrgFxeTQFT7CveSUrMEcw0lnzBujKtzUEQQ2cKIzp/0YE6hKEP1WzjF1JRy8G
RSqiHBasRnrUlcvw41khaqAFJGStBGZHHUb79r2Fj9jupZXEExjw5t1sl3vQmEqB
dkjgGtnIBYNye9Z6qYJgaScRWWgiMyUCPGJ6RmU+3QhGSZ1RYutOjiPMqf7qyCZR
FYAdE5VpAmcaYfGbQnm9skw8Dqu27TlfRLpfKi70gyzrLQ1VutriZb0fB+zvZhiY
5bkVFxqse4MJ/05LvdjcHOlBndm7d4Tq3ACZfj1VwgaEZzhNzSVgj423F/WcrRnb
bVM8jGYxO9EUGC/ghNP3z2GgNdDlnIJ1InD/aVIKjlACx/C7E55YFitjyLVV0Vg6
3z9TUFJntGqih69Diisoa9rt6LF1rQOPfkekU0U3CPeJUpXX03Sf3Nn6FhDbk7Qc
oAPgRElT2BMIsEwrPjJHsizraPjmV/ygT2IDTUOJ5sltUwcslAVwTU+ui8VXnhVB
r+P7T7H+cCmweq9PkS6Lk3WqHGoZWufceakKjKsWNSeIaRB/fTEZmQ8y/S6IYkqV
LAcGjL11XybJLKmMQOCEsEQriGzzTHowWZCv060b+XYUDaC6YbrngyqaCJxXwI4c
BF48gTgBIXNQSj+zZcnIKyXM8Gp27ko2u+mi83LSXPnmRMm2HE+cSJwf0yoLu2iZ
pVPBWFGyjv7vmH5UMvx7yUahZ6jw1m2PAH6TjOOHd64TGtzhWECm6bwT+3pqfbI5
wdM9PDebwyQW42cQh4kaKBNjtPiqHamoxpF2kxAsqyzUnkpiWoEpN1GqPpgW11BW
TSIeKM0Kv6cnJ8aNkt3NQRw2ZNqm34ae2Gf3JQfpiFHr5tD44djmPVw/iCpcDkGF
9Fw7srMwoIKk7rXjsrOWkLrk1tmr+2Pjrl/7ymzLEj/hv6sWAQ0lvGgp3F0WL+cj
COVZGTUD8Tprwxa5+51jXO9HxUBhkLqc9EHbbvc85I1v8XPvjrkIWGwXmLajtjsv
siV9VIEoa1SahD+vfs6k3fRsGa6T4Ma3AxiYpEyTfpSSNcef6qsxxDHiAY1ZE93w
5hkumqla82vLagE2eFOTyU0JJi3DqNM8raJxA3FoE7O8nlTCYLOMJxkh8jt/zDZI
C/TjeHCS4ldcem5A+S/CK/7JPastcJ++oaMepuv3quCs/dla/K/zWHGbyBvY+jBb
tegwZKnfDVekt+8OEMjavH2TtWJqJNsex8louLTov+IE8+sDjmBJIRLEhNcbIdM4
CuKkBs9+HtybWP0Kf7ZWIjyCC6XHHTvhRcxxBM5GBv4tnlL1J9nM1zYS/7tudqj8
LM+OKcuZwLVtK496B0I+9unlwmwyd1Q7bLuVRQn7UDpbyquQfvT6CzfnketJUj8q
dLMbe4amrxDhEbioxf+PTb+MNpVrfUrdX8kxAcvt79S+VdXw3m2wd+goDUzjq9bi
F9YWgXtcYPaHL6aREV62XUHWDM2XtUurVAFGsBRz4EwyMhsud1iak8U/d4uWwHi8
tUacXuky0Uoe6JiR7orkUr6U1PBG0JCxC10FmgiKJNyQdOHHsm1+OZ4OAxAC/Vtb
W+GZS5VsBLTr2J3KhzY8bk8Y1csyP9Eyf6Xng+s021n8j+7+rj0DcE+iftPhYsLB
fSf3TKmQ/GsJ/0bjwBl+80xLIS/2EMxNtfsJpoJHelZwfz6NiL86m/G/Hd1GswWp
RYiBeAnPmhu3kdDe6mj2q3QLtg+TwuzG7PrMRGhhe1FYrbqKAx8D+8Hu5sEXeaHU
PBkpj8zbLrj/hnQBnQcw+mQDYT2huj2jGR0YPkFnnGhKXyFhmL6E0IWw7oGmIOjP
NgNG+6oYWIw6r63QBBYnXZ65C/sA8S5S/z26JrMVnH75sf4LSauiSF+gI6gnEVzr
dniwGEolqT+Ha/N+73yoSYft3QFzEl3dFXfJF5zBY9BlREzGps76UagTGTP/MgJz
RVH06bJLMlvscnYeK0PxGexUgxh6TZ3R4L8aTb7Vcf/kfE19qcpfW27u18Tuw7dU
L/ktFEjVf/kz+NySgBEYQcT5mEXdw2mDtd1ZQk+RylewCT9ZPx1lMzkfe5C+tGA9
g7Jeh62z2pAd0fN+6gFHtD7ZwYCnf4tGbYOWh+bx6V1rasxWcm18o+sdTiMlXtA8
vTfeCVBCOdj2512IwT74OdYc/BKxG7uEAABj8sPVM9qKQSpZjZFhabVcz3WIqtE1
KIePUkhGRFtA1TFu9qbO5Bgy9ePonSAu2gvvzpAD0DTP1t+JnbUdx+CsMRvxxnEs
ULx98aIw175cw10y8yVLraBB4XXlRqvQ62JY9o+AWkXGp91w1STtH8kQowDwSn1J
9VhWO9OM4KsGwdihPOlc9+djEGyaI4bsIv2qWUHgVs+5xeZl0/k5Rn4cTOtbgP2S
It04SrgHlh10jddAEQO5Gwi06pSEcMorrfIUSAqPqA0BWfFobnCUicX6v0H6imV4
SeHZ9KEW0Q5z44j8L7IKfKu8/uAHuA2JDI8jiyTtAoeMTN+Hhp+lImwAtE+0wbUE
QnaYAHcH8UZShiLfnOw/VP7mfaxEobv8yJTRSOZrnWSmzI4vtKrxhSOK6IgFjZh2
K2052jiSRUylkC66p+RfMb32+ZXiUYwvxnRYQO4qqrdgV4L3+cke19osY2VfWH0b
l+rDXtuMV0CFybuwMRZWXoiPfJwCzLvFrDWPF+JvJF9BPh7YoAfhgkIjVaAlb8ne
W4TsEQbfJQ2cExK3AfO978PvcNb0wNWVy3MOQCCriVeqveaf/il3cFokeukmEOiB
sZ82VX0foSC7Qps4QqyG7eoUPkZVBTELcGHDtxxRXlWjPqzRviGWXDxRmaCgIR6B
ZKLYDN/HPouxfg0110rPLEGYCNo91IT8sqqVbkUqw+nwXGLzfk7OO0ehsOcfsYZz
QYzA/zxsLC6F2Z7O6coCOi2yRF+GhFRiRy/xTDytbowFPCte4hiE++Z5nkOFFyFe
boLJdA7IBi0OzbCXIA4vHyyYgdJAJ2dO857RCam//KY1bgsB+ZEzhftPAE6k4DPN
hCbmeWGKuxAjcuT+P15r7RWBDoQ2NBYtu0L41ZXC9sBmrI6MGjsD/tOmqwld1xyF
PsbIeK1sPwimyof/1irBCowqrGTUsxKLguQWnq4KlGfu/5y2J+z9tl3vR4rQmM3Q
YIVCxNcXe4oao5rzDbOd1G9lZd34mYQ2gvtMrNXykuHRVGllI9DlMjNWoPjfsOt0
SMUvjKXpZlEqlKnzRhuwdFYpfu5NrZs7+oH3did8+p/Dm3/qdQcXmi9zRAfP0azw
MxpVmw4wR+2pACqTHfLsliosLI8uzTR1kXQpUbj75bgVu9Xae48mzmtoBRHpZ4Bs
CVLCPqt+KXXm6JDSopdsiLF97UiLg8u6WOVMNIaPD+KeGaKkCywNzacM3jx9hUa9
jFc6rLpt8/A1WM3tXmIWsPXBgdP1gxE2vu57oXHJopabqV3ae0Ii7FFwm2R4mXJ2
U5rJp2TovFGWpR0bs2j7guP4yK68n7TjHx+rULtp0dWYcXO/t2/qPNQ4LblKogvR
q2LcKMzuFpJ5ViGR6vRFv+iUDgKfL78XIsICk71ZhpnR5e8Ib/uJXKPcMggDjKLv
ZQUXnjx58DVuXR1yUVYGhuRUJBjthxDU9/FtsWH6fqsHWFMQPEqaWO7aZVIsC/T1
NPutYB0fPtzjkEEg4ocBqS3fCd7X9bYS2MIOs7U6Tx6pNg65nVWhw+EVM7hFBdUD
li3bkm4TGBbmHkzFqCHnzHSwDKsSf1jLKpeUr9TnB9ZiH7KEUGv6hv7Z7PTlzbbA
BSj/UNrJCgvFN1czAf+T8ELi13ujvf3g0Mbu4JJUhxmMoVLd365wW1XMhvN/CPbq
AcQB/9YIjhwn1S0aMh+iTK1jRM+GkzuH/8GNxt3Y3abVBxJSEt4IR7Ny1UPcoLt3
FXp6EQnt5WlCknw+s7ponXSJN8ffZHHkTtkQmrno9GswTVn5ryVKD8WVSIypPfNN
QduawxBe4eclitfmUl14XBwU9U/JIQ88w/Zbh7zMau+JDpOjRGWSzG9rJFPW/vXL
yoCFoDWFsQrEF84R6DuFUUa55DUSkjXN3XGGIWzlXxXERwkQmZsQ9+luWIKwYlNy
OOMr3yUFuCR7ojK+zN334ndQjDJPhGYlHfbRKbxsFSjOF6KwGWvp9GCPPgoUv9s1
EBabeKsJ3iHZWsfGkhx7xyDT9NXcLusMtVUmbI7iuMl7AHZaSd/wqiXQsJ87Igfj
WbvmcVwXtKmKkraoK6exx2LyYo6HuxNSzSu/jKdxPK4suzuOJ76hJZQetsD9JSZg
pqKJ3/zPNt9XgnKZWIs2vJG9xk/Fs2PWdgQyBlUvDKQUxLScpAi0+lWVNWbvPOji
OUtQtd01HMTHF2+JiNQ3oQtrg8gu5/HsHmObMqT1SBk+u+VPT6zCj5rrEu0lCQ0b
bE5sQEp6eXi0wWOb+apkq67fx71oIvA0Zm9qsIkSfyd2S6oraeZP2uUfnNurC5sm
E8w5Caky5y+/cI/CrtADxT9ZOC+ar6P89QCmcyjl2xoYSfA2fa1dOklNjJdj9BtT
KESzl/p1lwJlZvnZOQ4bL8o8XFVpWxrjmpnpHC6s478lPn78qjP3m2FAQCEqo18+
eQokB6H/WWP48JZOQNRUv7cPgdLBhpN+hGB2He0JnsDSjXrgAZqfUa3hHm+FMPqw
BjhNd5ItzksSkAHaH4VB/LZy7Ju0hKJUDNvT6ZwHVDXA0yaiJ23wwAKhw7SU4k39
qBmfmcASfJOwjAmJWQ1HfVQzY8VhVqwOqFzX4lYeYsQfQGV2GuTe0RO6AjGKYNI+
HW5Z7Ego5h7rOOkbGDPv9NRVaJEyUppESUrSio3oi0Fq2wLFQr0LhVKvai0/XCfD
fVK9woYDGruszoRYNqCKg2NKRIQSNZrPPVJMIpyGWiMO6eVgT0FD6ZLt2heZ43aU
tkrg/UkfUU8Dz2pHaObwVthPlpCZpaVyQ6bDh7HIl+qnsOcixdyLWZjaOqt1s0m4
8ZAUTXtLxugGaLLyYB7Lzaal5cBdJeS21HUe1e2zq4z6qCBpEgCcJEHsUbWvJetR
gTsSBAsJu9YwEsvopPz2c6+iAj9xS+LX4qoSmAWbFjForMsHnYq6UG+h5zHTZZ+I
/rNFvcAdf+azVI8UZQaRwypwLDZprE4z3RAP6HkNd+2ahKjYS4RVSgS13FKFOuPL
nWxcIBe7uKTbAfoHIzPBf1n5EtYpGlx/39neIZvVx74O6XR61E+Yj7agz7YE1CdG
5mLzdwZzl84L+mGlM3wDQpARZ6CiNijt/DlU3BptvwbWieqZSZLAu8yFDGqg0yVU
VAvmejFq7rTVnpluZmt0k5UdRFjMzWlYy5tkDHz0eEcxoIqm1dIHLAilza5Ixy81
e006MnRa5IcBKkV4ZYn130sQzmWUHkzXhzZSxwmvXccbJCQsDYiNJY+YO/7AaOyA
YqP0Nls2qAThlv1UFcsNaDoXANUZN+KL17YyF2koNAfLoXn/3UHyWVOCPTuDvIVV
slf1V///plthlTKAx5TSwnacagSk6sIXlC+/mJskGoaCcL9wo4Rrg3i7VRQem3L3
2Rp00UoH+9o5ZneGPaxILU9oxJSmZr83F/X/6Y0Vc16KfOP1k7FMEYG7yBSdD1c3
BPWwmS3l7zh0p11GXz6dN68wjfHaw/gyqS0JPpYvJEG762jKwb7NQfYUq8sWP8UR
sR5fviTHq9xf/tRnzA648RBGgTClr5H6am8aOU+cLZNNF3kuYzLo9KrxFIuWOD9e
zuy4Wlm9TFiW5VMjyuPwBEn2PVKRMIPIuqMDbuU7d6ISKSfQDs3ngHt0kIz2Lvq0
Q+iiQJBSubAtZf9S9OmnEKqVf8+9+rhkwTGJ1un3l48XOcnECtIM9Qw0J+UWYZuK
sOwDKxzIIACy5sxLtmGvIrCuRSXw7D1kZUdNTV4n+m4WLV59Cg5O7o2P9buRkqfT
DM6ELjzY3P7+OeQH7KNnrjWbUDRCHLhkBX/sUSMN2Gzd6ZpOpiRiGsUu3xGOKe0i
LW/XMi/sOkeOetsHbaFGlfsthTiyNJNXhQyVd7Nm0cVEbvoTUT/15fmFezrBpe4I
4uNr5dGLD/QSQn1qAiAZQ4KfP+/YBa+suz7D37rayXF25THkMlWESi+5g5MctjZv
c6EG1iCrcSnP3lyT/rhkAlo9AW6QSRHL2Y0gNE/uTw+7z02K2sF/zcqBnF5co6Hh
BgYcK1FKVkMUKxezVvrS7DV+w3tgpZNcq7samhETshVXjvTuwMJ1T69nqUslaCVu
umsn9eZfbHSU6LXt+o79z51Y4cOmf79uIxNSjtsekpelqJBwCIg8yiOFTxm6r3K1
1VM6tzqJvE66oBq/HXpTKuJT759f+4oI/UqwUkzNMaTBGt5Xb70oJiB+Oo4r6KQp
M4xpYnGwARcpS2IztoVWAAhwHchnJe59eJu91P9bCsj9/VIqTpguCzO3mITAnURg
kVO2Gx0+LsdbhOptklR8FpLx8TFfZ4eNYmki6JNdHBT8Rrs1zNL5YzDiCZX1cmzV
Xx204hHY3Grx5VuUXHZB/W6rMniKRULT6v86wTrhK/EG9yEgGvYVfHU5L52U1s9I
X5ik1XwHlCDk8hqDRuOUbdF5VbAPB2kMJnuxzQgFNlzyo56YAsbCOA7asSM1GWTg
0bD3cHHjEw385GbHoTcdaIlaQ4tW+VE1AbBsnbsV9GnXEqFlfZidLr7wFpjBbtmN
hXSP1Hjs6J0WNuMa8WVOcvdhbom952ZPO1w0ZiPANFi852XyBmZalefoh0Bjw7wZ
GXb6BVm7J1dA+EgIWqMiQ4i0dXoMAuO/vg6Ei0ZCAIzO1VvUEI9G/+pF6OIv84p8
EIJvpzJhAmNK0XSPzrA9F1AtxFzIeCAYqzb9u7D0eqlMmf21nhP/hhzdsuq5pJ/6
q6ZnYttixX01kczld+k79NTsZ+i8Vc/yR3oofquFpUOGB7tSjilVQtA3y1CZb5lh
2P6cczfwjZQSKHqmGTp2LMFNI6cuMDMU/aQE9eE3DAKW4nMAbZ+r14lGd/dRyHGt
/Zn+7BsXLUDqy2DYqIbtJt3APBkbRWUMx1AiVvKD8MCZapu3DZuA1wgFeQr4EiMG
ecHNKrii7z3GZifzJ9TqEHtKGCWIWZG9wwIgnlPje5fpNll7qe8q0qqX/j3KyBCB
WdzQWQhqqu4qDkDQPWSZOYnIQ7bMNBsupBjd/IvfW4v427GL5v1fMVUjzyCo9IZf
uxQ9Tznakf2Z4Xe21RiZ3Q0r2IG/r9HZZCIdCDV1dw5nr7KxUKsXdNSiAyvIkNCk
ZfNkUP2YwVN5HgOGAt29ly/PTN5gd29O35iMN26XLLTK73zfC+MdoLPcTOey6/rR
aFRZXSeEVJME88Noiun2I46iB7Tyief6YVH/qYcsfi4Jcx+FXYmUmW06Ojap09JJ
YZIfWrSm1oZabFpRYUUEzYsg6UWjaisizs/AHF2R6CbkT3VlxEF0p2XcHgWMZ7ib
HDE91nlDsnDwVlpztAqaNp3T1wxXHxGtrsQFsCtikc9qBWualpWDoYIF/jd/8pD1
4Wjj2UqZYOING3w+TJAI1ubqoGwi2WdWUedXwCgD3g0kloEr2f61n+osfcKPR5Xd
5asIGxN6SM+r+2IXnEXX8VkOFCDDQRTobfKTchY9PA3UJg+ObO+NFUVj7T1Y8j5u
xLpfj8yAaUoNDifyilT9FZ3xbCJt2qU63lhs7ypngY6ZcZu6AopYu8PAzLiTG3Cm
+beoIDIF9jXruziijxEEj8UZI5kwEDfMLofKXOUaap3uDpGz9cpCm25qahpNWRm/
uZemNawjEcnBQVuZMuTEkGubEuHoeHRGgQmqOEdJdAB7RLI6puQvceBODFvzZ8O3
kF4WnOgOspGW7FT1tBOvJCPvkP39O9tmbRUDjv4Bft9GB5csInc6p1UeAIYx2l1m
9G3OQzZs4KAEeYTP2tK+qKpWrrr6MW0JCRIWjkKE84x6qo1VXtzWDfiVEj+0I9yL
HS9D98nI9AWcyIsnF8qukwg8L7OFQ1Ej2245erx8EEQ9TQPsZ8kPJel1/WZhgw1z
2a0d0xncuXodnqzSqjCgI8f/jvSnG07e0kBr9wX1eheB+EJ1gX636buHnIKjMj9b
sLMuHhRB+QWlT5k9yK7P3c1KCu4GSCJ16Y27QJT4uUyFnWvB9JtBExVW6W5eVK19
akmxqPfgVciJ/COru/GP5HCaRtGo9LcycLkelbaUxqlWVPZu23i7Lw/cJK8C713J
s3+UJrVz0wlxvC2TOzlC0QDxsvoCzR5wxri7X8mDtV+qFydZLAwcyzhyr04UyWaW
Y08ZsriuxBwfYCHs/bisDALDKD7WcqLbBGg/D1dWjGqJsCnitfY8ZtHXHVSdw3J3
sxeceef5Cr23gb9D2IyMyT931vaHeII8o2Xy5+zpnathVQwvwJkexpRHG9QmPQDM
5gkczWVAKZBFInvorkbOI+vlpTnCt5cqa+C0XDweO8wxrSs/3CsjYwy8KUDwpKPB
MCOg7x36SMpoEK1kxSwCEbcBkLUXL9yWHFWRt+OphcLd4opFNX/cv2TDLCgseN8i
+uftBDdlGIkaMPabsZdJjrrUoCp7ZN8iz0Z1GY8AspWPm+3Fm86TypvmtnY8qJQ1
zNldOEZT97Fq/Gu48YcpBLwUAixHOPIxHXBorlJ1lyA2IpWhM1DSlaOgElenNeeT
xjSCbDMbleGIjWhimklQmXIg8kDMw74ZrkN4TCHCUrGbz89vUveIiWiAVfz67QgK
fEYSZSm1+1VeSTF1Pvw4g9jk3I+pRu7udptTaoKl2dUrm5PVT+EgcerCmsuaCYOc
As3oku5WH+f13iTDmXyh203BErNG+lLsKIwhet6bcB7OmSQo37ZUMaL6Jz3PlzEK
l4ea4d0KH0anqREnGjczcBv1+Hyh4AB5T8Mk805kwBKO4abjbSnxYf3AE+cNhPSZ
2cfoomEa40w6KByaLHxppr1BFWU+59QRh4ka8q3PMRbVQd+CacNSTMSJJTJs/RAv
DiAI8JFoH083ufSkjzRmx68Ptkaf2O6KTd4GINfcGWJTbyA1yVoF2CS31eklCafJ
MDpMx0q0qSzsu+sN0YCIWoxno3mrD8S6N+2bPO1/BpdRYdrgy3efUOFcQ0FH1rYI
9Ade77D0nNtT2xyzDYtaiSwb5/fD3MUP9XfMNuoaDmZNIKGbNfdV4HnzAmUGxV2/
q0HzGLemTuul+e6CqfSZHBLqHtpWKzQYeO2TuPo17VqDLFV/VOvnhrF9jINeA9F4
y8aLSD3363G3fzL5NM73E9R8SlUGloMy0nimryWQBqi8ZSqo/H3AFMKpx9taGr+K
nIz5HlrPrNJZ9+qA0eM0ecF/1G3+ZXW2ixe+OqXKuAsyc6+jjFfCCiAsfN+rlBQN
6EzCtlAJri79cAf+snNC1RDKnx8aXokSQq6jTC/+iwfITX3MVPMJBgh/o1w0bP6v
cpem8p5X2sV6/Hn5i/huYz03NzvkUqjxede6Yb4Q/EZcnlT+IVEJUeEUxabRRhhr
UASyCowKtl1snK2YePivx9TBmgPAD2ePkmgC+Phnn7aUIQtwZ9P2W46E7IAe8eHo
cU3DfXdxCxIeWIaaL2vc1xYuZrtVjz8Dw0HL8oTTSQbI8VTV0ii+Caa2hDp2xcGe
gHanXQJ9Vz3uC7ve1A3pwcmedVf2XaYSaLBZ66MJpnwzb8c7yDUWFcgwj0xhvQEZ
SUvgJ1JBUXFL8Dw31PkoTgq8DBK3bmeRR2V6e++qQszBC3pYk9bkqan01nUH1hyG
Rj8ZbgV/i+t/vAll3iXnQzBCvVD/uZZ/R9SoGOKB9kiGhxnG2Rzy4+tQA2RM7ZGa
cp0EzsogPEa+jX6u2oO/wifrjj+CKHB/NN2BMmFXXBT/SWsQPbhjgaj9cUS1gw/D
ZlPGsL6cuHhj6+gIbDM15NAfnqD6IlhYnONtXuMvXp4+BqKH35s7LwK4XjqAooZI
Lw76GCBRa6r72OUg1QmGGpstz9N0lvxt4nNQVfTpTWvUEVJBA+04c4ns4yv/Adef
1JQd4Oz3UQTJhzBIcGfFryU5OcqLsIKN3G8h0uA4cQtKs/Uz4KIZPh9PgAbs5SaH
7YolD1dwPqaKT0vXUm86m6+HSPip/5LJv11zk7DuORp7/46RFYIVHpR8nee/F3TZ
Mrtu2OqPVOBEZgP8gAYtK2xXWuBgFgXwc/YXoqvKHY/AHG8qaK1AEyt8OLplPau8
JylOhj+KCQ+oDElaG/BQUuGUhmzTI+UyWzwpF65QfDc14C8IcfeNF29NU+sVwnaO
6d4DIwkgRSzPVxCzWLq3zK+PQC57QDa+VlEZx2O7Z6ILB/XPqOv8f4+W5rw9jD2A
BDSK4v1pf6jnpGT5VIiDhSYl9emtThAjuh+HPwbWQsNaT22gVGuMhHB5SHyEpgTl
GQbp9qNAQalx48NZBssekkOW2tYuyiNxW13mzbgjBHS98MS0dEKYH5oH7P/PSMSF
3nV4p26ju3yAQSy6defNUZM6JCF5WoJrk5NUdvyUJ9N6qlZzbb9P/bDNX4tS87Pe
BTfSnNA3D+EB27AHek5FeOxsy0nSQ6YkdEhf7wOEOlCmQ1SO252pXF4fL8kiiMT3
uUtjig6gg1leS3hn4PeDWGxZKHybFvvZzRSZgQMb1OSWEbKrmfFKMlUcdLyEObt/
N+FpiELTAiuske3mtT9vxyPnU4GfbziojuZc/ckBC5TAu9vjfUJWCsFyW/9ePNMd
8fLCfPWNTZMTvppyOITMYmkdFJ8M+GNm6j2eK+a0/cdtkgqh/L+Q2FLEVKPwrHOw
6ZvwSAUG46KlPbk1djaY+ixIvsZPwRMgbCkUuAvHVvF6O2ACLr1r6MmFhXt1dAC5
h+KlaHJkU44DNHogqo5Pp5LY5CbAkbgUVQv5WE26SvPyemHB+BnVIxaIQChqxwlv
V9u8JV2M3EP5a5aRp6oESuHx3oM/RnQBvbltPL//5VGOIrhjT0sW+SUqSjKsB9JY
CzdT80nin/ThprnPXHplgv0SzssfTCbolwj6lAgvWUkbDZe1fts9EKO5s4m4USYT
JN8uecJLsmCH70XrNqEZiweB/PVltGZuk8Dzl40NcgqWapjsxn+mt9Ikwhgn5WD6
rwypa+7mMxZOsG+RCVXwPIqTh6xF8bNG6s+34PUA8KIcBnMMbLY42ja2PsKXlBnV
Z03ncG4MHa4Q8BDuD0ZuLmtpUvCMOSwcQi9LMeJ3Ap38oknjIbHzh2zYhpM29EtK
iS5ymQ8Lq3ZmShFcqpDvYLCr5psraY+aDY4ISGKsZsFNNY0kXU7gXi6ZNh2/TnJ/
weN/MwC/NwjmY8Qlru9wc67hR+2Gy77b+WjpkVF7LuBxph6UmqLORnpXg1JZH57V
5FFN5NVFyj4By5gPJwbyEXY7RBcDJjShPHCIuS4BO2NHj+59xUILVNSnQbsUA5Ad
s9RoPAbcp0VnqfzKRFBxgTThIcUFseb9IRT4NI8lccIXDSAjhmR9TKoPcnLShWJy
eK/EUIkZwh1uQTtmJkf7X8rAu5aS/98Pgryea6XMl0Cb4T7NyOBGbODeDIuxbsYP
mXq93PdMWFiS12FyBN3FBuaJC/LfvA3NKOvVtLJwHQEf1420mYJ2iO4kRwtgcbsk
d8yVW7r+tEanFjkoDEXtVqCJAaNl09hNlTu6BkA8jUW9cmEzazVMGbBfZN70yytY
9tzY8MlR5/yxmd5u4hyogVRQmovgcnEUka5ZmXNUIBmbSXQaNfBYufPb+BmL3PNV
ors7J7v9u36oF3frKv/YYC3Ken3N7uj5BxPYlAit6Mu5hB3McrkKskSx7BMDucpi
Ts5NmJrM4PkM6T6wYT1IabyqYdEhDhVO/DUaYtxgRaQp+l6Si7Dbwtp1TDQBFuvX
sHJvWEFQ7WhDL0gRlwORZSh8uHn5Ty3PhSe4YCfEvvhLl+j1s8/QRZvxzaLg5wmE
MaegccRyQNTcOvgFGTobaz05QFZ3fNGxjgZCtYFLDsuRbWr50d3E8MVpvan+fJIP
ayEJLFmnuvkS5fvGuOHcZoI8GaQLKZO6qB2r1LQt50cixAhMyEhfX6Z0HNlKvamK
x/JLutGNITlYWCwRx8ztdemhM4nHyTJnRyR/Q+m8Mn/soVHZQwMGkHAe6CJI+5gW
Q3DSmajdEOhqGV6Xb1kTywsb4CQifpzJ1a8ZR82GCjFYD3HSZ243i69T7fbH4Hw5
phupzAbzeJYpVNWv+GLlQ/msQ5xuem6liqCKwsxEUeIH7fHinI4QTK8Eixa+k7Gb
KzqRr4+Vto2apbdKiEqmkDG/ziFZNc87zPWEbLXuZFn1V7TBJyUYc11xxeF6jlWl
oJ7MYKNCv4GfyXVDcp7FU3N/QZ3umUgH1JlmjcxFAUHuzqzYWoMis69QEV6NL165
kjrTadXhT9XEhuFS+hv2sr1kjqFFXQGipo7JRmt5xQRpLjdmS26V0DK/pGx73hUP
swUHXyccNhYIbRewnrcsCLKN88ehX1vX04z3uZcAXGehZjWrh7l+s4Hil/Z+cVwA
xy7CrPn4UH240nj4iDbxYBgm/FnaPHqk/yb8JO79SmSy0nDnVSIl/MFu+s9ZYtgn
FoGRxREfg4bGbtokwsvLV8L0kUyWEyVrfPr8cYrG7K2stP5X0TvozxmYjlcPgSRx
y02oMd3X27vCfapWCxm0dprVxJjdfzH254+YwXsqpgzElv9aXHByJoesosstrEPP
bTVJxEtnKmxZ6DOOzgtN6IQN16JJqbfy0xGx9pideDo3seAneKGowZWqs9WZqq3f
/9qdSzSmq5ootn46ZouypkHAJacxtAgd7Sv6AIneUTJTAuNSmML/PEzNaQJuLaY1
tr3W/HIG/uVetdPPTtz7POdTR8h8i/n8Ih/4TMWxZ2UVzxcZvW/P54QKqvF6uQ9d
2pxObP9/P8aeOnyCdhMZZ2cr9V7d2YRMjnr77+Zf8e8AG44fea+UjcCMLsV/62SO
Rr41QFM7ORale/d+WlEFFcUFwiY2XWxSitE0YWlYFDdoyWIuOc166RNYlhAxqNIO
k52Qz9I3Rm1/UBC/7zNo+Tm6Az5HtYh+yWbW7PMYO77MoM1jmfXsiZLkmsGtQXJ+
oVx4dqo+t+hKZAb1A7lk7IWJPdj2ff0V7glH2KnbUqeM2QDWLlBM3wYNMgnVYUc/
jBXuDd+yQdZSYhhsPMxirNSRJgIR8g2k4xiyMbTXpaQnXhkvoRtuOmTa26oOOJ9B
co9dERtuw0HFHqNsvaaBczXweTtEC9YbXzVKGKkSyHqCHhEeQ5fp8pwjJgg+tg1Y
lJf4nap4+lQl8CXu+bAu9rH2fre3zcwRvkb/5DrWsS7zfeO4x+iMEVkz11lK+kZ+
Xf23Be6PBHqNW+41L1j8ZUo1HC9nDRccUTOPB7YSbHTtr/xkgqvuHkVoJ8F7UNZf
Z4Nrr2JTwQXfOAjgblBL7/JClzfUFYy5+CYtVlHfroYf8oof3NPyYOmOxMrMstWM
hek6cDUMmSJir0OgD/WtY9QdVpyQqGVT+sWsV1TBPocQVeFHhhT4UYsxqOLvzcLu
dVrHtzl8/AlXbdKcHMN8IdkkTgVZZFVFNGOjOcy1iz1DhY+nhVzHXQBw9GwXpkkq
hWpAp+n+eA8/DkX9uY/f1L1apHwqhiHZg8T9XHcEYg2BWlPsEWDGXMCY3EB2XlQa
e5W9rDkBAUjfcVKAJvOaEP3lQhY9XvnmcIQC1CdcF7ZcCdSuA5VdtP6JCSxPaAGz
h5svvQ9kTJ0zyTW2Zo8nxIJm92LqsgLzzmG79s2V16UpCsf3AeuKl9KcIGfoNFSe
4NqkdewpdYpuv1Wwnbm5E9xEjAU+JbTYsIjj+dez2MRoIxAfC0UmagGaAcBdAqk9
jqREdbUYSZ15Ioes6HAunjpVg4UyAcc2i2UMeDbl7tOgUFh7HX8O8dhueK3M+f3J
XZUzcOcdGsPIF9+j9nXf+ptOJ10WTIiWEmppJColWq3MUYN55q/4W/rYfc3V/HBT
OwVMs5x2Xue9IWDOmYvbaG9f+phd3x3tcHwqUATEInXKoxuOtNRm4jJoLh2+p6Ct
JLsuJ1md3TTv8gx1iVgkfFMO38kievO20o4q7DuHVkJVIq8NZ/o6pXzL2FJwOsEG
k33fv2jimQcUnzgnWg6SFrqUxZM5RBVePCcryURKZLpssbxi+DwoXF3rUP9uHk6t
pQVwyWuT/nkxVLt1ynn/5PIgSkqKe+BoXOMJqMQKVE8qNQeYx0Gs5McRf+gZhkAA
Zq4CNHOTzLlIxuttf+8PQaVtu3WvroaWnzwa4fYLlPaLzhpK/jP8B2ucNLv+SAsV
bC9KOX37DWjyWMY3GCMMwbJD75W5gFAogNM5NP2ubiTdcfKxAKUnbZ9dKMPW7Nya
fDgvcJEo6AjG2tm5xtUXpGATnh2qarAHtp5JJj3Obn5ZUur6iDjiy8yk/fuVahH/
Pmtk9koczQqonh/2S0WZvGIo21lVmC3aMWmIi8Vs02l7g1psFj8IkRt8txsEPBW2
Gtg+w4Ou9npBH4B6CppngEISa1LykDvVMdngcjbSRGbVBZVmI/eO86DsbOSRkwaO
/wQwlNxf+ZEkfZbk2PkHA5IStvDYNFIGe6J/62M2ngxXiXeWcu7KuoeQX9A4JEz2
1Wtw3Stn5w8tklZgLiwyTGPlPaGiipV0oN8lRDfdyKpk9rjXgyFaROCCMfmxljtC
p0wpv+WC6RSSorh6SpKH9iBE7OyV2t8yOc12w7yF6EyqJq6f/SXtVClO7H3qCsCN
hHmrkjNiMjdGP99CYVfPtHADVL+bBUSAMvDFZcCf8zNGeOLm46d9JKpcDMddavBc
KVoVNWyZz5UPk4XDFSBS43uP5IrWZ27aR8GjERn7XzLPOAHuUQxX6kr2xAhdU+C/
4Bo4XbnlDKSB11jyuSqLLX5uzjn5Z4ds2nNbb3HBABA7ZCarGHVcc6Jz+KYQvzF0
ENZMarHP5bn+/FsGVWg572bZcy0+2n8CcmDPfgox5oI8ILJw4ku43WeLChf+2DV5
xkCU4epTnR71b3rR385OXfzMOJMKZry+pJy0EcvFGE11xoDImigm5xV6WO07Q1L2
2pl1gnsfBavj9QTgrv5piti+KB95XcBmOwC5S1OC3sEQWBvLOk0ng/9M9WtcTXfT
ZpDIu21x/0K3OHNsclXM6Xl9+/Il2gPGUGSQBXItlr8fSHqUCeFRhbzAB1D9ID/D
GZMvWtkcQdSbSdheknrRuA3AzHEdSwer0fKqteTseAJuPMOZsMnSvW8/B19OGBt6
J02m5BEkBjSnpZeyIt/WEZBJCvx4Wlb3nnlsbtI8MUjvUGOX8LYmycznuGuQyPEJ
UN0TbcR1lTZrS0fC/lnXz4zDwK6oipdoe4xaS1BBP9Fn/yeDHoI7vFAcU0JLoGcq
x6vwlGqyqMTkaDyyGE1MCXRchirIbzcZbRkG4qeWlTymFx2E/ui5Pu/UmilVdRlM
5VXVmQ4Mxyi+Kr2cvMKaftdPs9Jk61f+ZFRv2kN/riYx8qv4FIe7Xwcs8SehojaR
WCUUFukXYckFEqwrtbcuzFftYR2zA3iEhmVo57mvMje8ZoIk9OaLfSe9fbqlpDiD
B4M8Lc5ZNtmhoryubYwyarZDDardKPH2R5hbSh9UJc6qNCbg7dm8QoJmyevk241o
vmruQx9LFOIXy12J+5invyJvkQToQS83/N/Yn7rB1oybAgbeMby560ten7/I3P1L
s8qWowb1I0YE890Y9UyKwkWfL+FzXTiK4s1C6CDahpC728a9LPBpwImvcYQDLILF
nMpi0p2Pg4bGNtKogqvJeNFOY/iKY8FhIDh8zZqAFi/XtpB9f6WS1hW6rB4wbs4Y
dyi9qC5QZjOTMZksUmiiGfyqpm8FhdKFQLU65Z7eojD9hEMvnw4Fr3/BaxOvutqT
sufMj3cm8jOIFrZqpgPHphtyk+irJGZqxysb7CFicBtSmMfscxqUAdsUcmuwA/GR
KKzVDCX/hwzB1vWtiazZ7X0Eco6RxiEn4zwMBPz0C7FzuJrGgdK7ZuaTiadXEV6O
38GOxmPLcmPgtCizNZ2hdgXtOMlV9rnxHlxtxao46JWrAXZ+k/zeAndc7G/wBAfg
QGyQ/4doUSZYhnpvU2gpvFbQtQFqXS8XIxasPH5YpvR7jXXhQENBXO4TaTVh9Fwc
BYq5OYZJuySD8zf/+MJByfuv8dSyAQC8vxFrbh0yypoNXLOkw+/cBm55oLBSL55s
zSlVIoKA5a7UffxawT9is+J53W1wSVslrYOtWZeaC7Tc3ZZ139qo1LKd/evwyatH
yc5NvpvNCr92kaZiMB0td+N2AUFwRcuOgroMBgxT4tFckcKMgQ4NykvZTDMLrQTD
rChNaWasFaF6D1QJI4QTE0x8GD4bNXVP6Pq5IaFgtIsbv7Cpuxo9WMgTDaq0s1Vi
LxiwVG+LBFzk/VTPCOvBV01dZVyOF8CO7g6NG4xt9zPi4Wjf6LXX1Pm0yjxjNlx0
snGK0n9CUm/ftOO6E2ETKH5UuHvXl4AmIruXey8mlqvkL9oB9wl/dZrYcWQc264I
Zl7HLEXOZiusQZ/b1+BVp2GIQ6yvSzMTz4pFR8xpZqECiRhc4yUpTFWcb00kmGQ9
CS5u77dnIwOD36VNItQWgAjXmtsu+/4/unCs5xrROxzBG3E/HblrTOhj/xyXLLvO
xOjZRJROqo3ceGFpuki1u5tB49JZg+Fl9kOVnyZFdJ0KtMdRyeASTE1h9Gf7lUKe
TRjhv05VOWh8IcS/liwcvf/RxY/cXKxQganUdMY8dRCAyGUNwdgQ2JeJHkdPIdtM
vTasTYBYWNKN4q8pMI328oXk6Cih46PF2gd0ykMmCY8oZz1mqBN1jqx7FlkWngpf
kC0w0FiFoHMgA7/dbNJY+xKmIxGLv788/G1VULWaCjzPRfv8Tq7hHog7KGqivnsE
VGNKboDZ/x5r4MOqUr9MMHkIX/V1R3PzXRsspqWY0Cg/sa++ch9AEMa3yZ1dfeL5
LF7oMqk1QqbXgSm0gVfqqTAzHUTFwO+QfAPyiyKlFCCcf1E+Knh+oqQZzAHiKKP2
+JlukRRfkx3B5rmpx+Rh+T2Ut2KkZ3SIIOMOOSbrmvUf/qF+FO22QBDl8/fj19I0
vbM57DnbVNpBJFTFa0HgmrnlOQvwL97bLWzwBxpJmrOZlToRsbChrqdJQ7H4ldGA
MsVShWwEb7ZspEVBf81GQI+rDeJZE8rZXP8YzGeN7qwOVbwdcMIgeKct4vHCQWnk
iCIHzXopGIjO4TSh4jbpjLr4VT8/3sSavkc7UsmriHUiXsuyAPq2rTK8c3Ecz+tR
Q/+M5YqCzasNTlj2uRekNmdFx4OETPt8isqIhAJPmHhjaKqTdx3ap7BTiXebLtaW
gNF5c4m6quCHztQP5h5183FMnI0yu5fSMB5OFIsDKj21p5RW3DM6rLUK7ScsgarI
hZUGh+vjiWwnizEbylpOKL2Mrs/ifj9hS9b7AWjEbUg2a7kUOTuM/UBJdzMvEoDG
TXoAUEngzrPn2hSKCuMVbQ+hJtquwYT/e3br2X+nVk3ki5dZNXJM6ougmIVnvUSy
VU8snOC27j9rDweUacOe1fQgVnK+PsznXJlm+/9WIMGeF5BQum1AoMqWOr5lSFFd
H3Zq4uYLOyxcm0Kb4kWJ+YLvX5mrcxTTcw/IgCoAqB9syebM9tII99T4oQKD5d3d
vSe7zYyUh4QbBHrduW2x52xRFydKXMhz6BLRIddfBzDWXAdD2RSXj2AEdvN7pTqU
ICd5WCQBBhjBtaHZYEkxAuTo5pfxWC4cpleepQPw5z1LMS1qeVG/yp5KzKF+NC9g
OzKiYeN2WS5xDESG9ymYn/echaX8vRaRAd7SbE0cpj1apdQwu+jBosqq30F78G9n
7ZnhedlRA1Epk2P6MSTOs6Glfo2RScF8nzTXCJ0DABvP6FcspC1ZzhK327MkgyhY
sJbpl6NX+pevld+thGJXdfxuJ52lPR5xZBqg+Qc5icipqdBQRvEFu/dcUlLaRcBc
ck4AkyZk2DGInJt3tqdFeYqQ7ioydmYyL7awwUHMwzSqcUo0NfXChMOdKNrG9nBO
01Onh95yQ0vmsWPcqJor8lZQfGPTqJ1v/1PAdnpFBUcrQ6PoHe83EqBW+sUs/hPX
ar0xCevKw6kRCjcHQ/mBBM5cl8zdNUtq80JlxYiONMfKb9IJxWzIF7+C32kItsPT
VzXenqVbATOyNlCTsFs+ayq+YOBrSueMT+559fWsX9fZClezVZBdbYvLz9TPqt7g
rwV+e/dmQ0tm/v9CjceHMr8keJz9LVu9QFScbCyUwxdDy+jdk0yMzrOwhu7VufjM
cMVdv5re+aZqfKwgpPCumRSOBNjC9hfK7SuMg20KV7MpNwHd+d9bOAB6zCAFJHuy
00O+nLEOHDeeURYP44RPSpu8XaihiEG/68PadkoOzOrXHgySGEm+CJcnj8rqr9lD
4yBpWWcqoR7xvXkVXO1/xfx8CUSPb4i2w1GpdKpqmkZoEScBPnGkgzCyjg2Pa12R
5OM83vZ2mn3YtwpQmy6Uo3h+zQ2ggXUDyeREYnSGklBeJWQz9qPZJxien0DbVt6U
5Psoz6vr1qlTEYoMDJdrAqnT7wNflTBXkXZoF4UZp86/IKflgSkJZ7/JhaJErCUk
y/s3h2YuuGOFoZaK+al61Cw373Ak8lIBMavzDovrIMwblvXqzeqbXsrSkrtNdZU8
MfRfNP9qbAuxDnEzCwNJ6luQzYYe4FGd1DVg+juvez58VcSe3rI/HyS1JPnWzIlA
IZ5gpdXKDlH1+VDz9/0JE+SLSrhusuDOzc5n962kG4Qv0xrazKyp6T+bMt/vpILY
KSYKZ87im/89fSvl6roTlwQH8XyMNaiJkBwJUPMByEbDJBmZbA6SwRuyCCHOF6Xd
Lz8qbjbfpmdlc24q8Zi6A51GrQPN/cyB4wAgg9WfdmH7IVg+6bT9QZZGhnfWijWu
H06VfxhFy0hQ5iMGO3W/W37zGR0NaMiS4TDVjSVMOVsAKnDJyQtFoncn8LV2ErXU
D7KL6png4XfGrsboeP6wcbASuwQaSXjZzFQgmznL50L+mz7NpqCBkcHd+T6hqU7o
Als4galzt49IaQZC7RQa2EYP+SSfDQldYo5MNmFVrDrTF4rawErCSW8m7WBL+2+f
AfngNQMu4KMN8xQCGwoqxRBxJAYV7boAFBrVzzSS5ism/PC1z1X3en7QMz6JyFI5
TGrHbvadCilNxUNkM3gR0ogGnOk03URSaXOM5qwMtZvimLavox4zLWMByVFzpDjf
kyb4PFMqYQDuRZ7BVAjfLCA5eB5Kv8xfXUhl9EoNceAZNl4bt9TCZQD/f7gDzkRV
Ewgn4DsLWNwrei6X4y99JeAwVmhKNBwX1iZnG9OgQNw680+LGL9OycuhGPkcC9CO
/zYHxrzdfBTWBItjXNaOi4+xo9CBjDfJVQf8c/DgCetZG9AXtR9kRUVNVC3h4CeA
1iglQylGLW4u2U7ujtG2XAbT7CAsWbdEvRyRZ3eYWjjkQrjKvcN0BTnmmP3BEgPx
mFeKPq4SsmyFShiD70SDOAfbTzWw/zZ8YlgG8HYMnHhGzpXz2NUvK8RMDoRMPi5d
iUPj2hZulf4stVGBZJb0Vjs9XTPPQm+x+M+VfNSXl0o1JZcLK69vqB1zyk55c06T
UE0xEVLDbNPXSGgTdHOWsMVmxrNMW9HFvOg5mHuLiDzM4l9RgaKMFfXvG9J3zWvK
a55hBVoIVGUGIgK+oFprWAuJMpaqHdVzwqn6aNgu/MHzp+NyKGM0H1liNKmo1uy1
OZUjZQNJC1Ru5gCAWiNjCuPOiZ08IRJLhG3kARRYN4HeMfUbhg9qcXPeSaqEo7uP
7o7rQL77BjTGBp1hg9oXYCav2YLL/Wg3V0J6k/+8cwjalgOVVYN4wa6oULMLsGxo
SkXvI4lF0076Qxwy6NQwvZAy2jua0rm7hp6LZV3dvedj/o2y5Qnadxizauo8o5Nj
s9KY443bfUxwq20BmRPQIRfEEqPlL2gaQNk4rCcuVQIEomWR1/22ib76rh6/oYOi
A/NauxZ2cNW/Cky3Y0Z0OsnM8PjP4HFaGFe5UccfpRQLTpKmC8RCzob0yWrINogi
9S+cb0I72XyC3Nv5nsWJ0ad8B+IC5Qnk3IzOY3xt2zBtwHzl1DfwjVFb5moqq3TM
fzbpS24azfzNIal82vfl6Fiu/CwoQj09UY2hUR2LnW3tPL+wA6Wyl2OzTaKeqdnv
Nmr+GErF4uHEx8tshTR0K8V/e4eXBUQOhCWw6Bcmt6TJp2+SXzw7zvienuSFDtvB
aN+PH8Ick6j1xKdNT/qnHmRG32qCqFM9Tl9Oqdbl1f/8NkaHXzXwHpax+iRBaBs/
FAfwqnRI6TreJZSKGdF1N3h4KQKvWjy5lxYx9EkAbP/UJzk0TegJ3jYH2ifYGKPk
d4anfmYE0G89b6G7INAQYo4mPvLABl4OIEDhpdPsvkC0jmKjgCEOYoWpaC7J6hB9
RKtnuvKqDi6WXCcjz3v6KN7ZUOu1NZ1KLO7hTuIR/HU79c82yeZS+9FJE//BOIFX
f/PPuCzKGBhe9/erArbfE1VhWRP+DJ46cn4GK3b2hPbcKMcr8tNDzXw9BhBohREF
HXPNbwfVfcMkhS3URytdTkoLwZErYaryL/1LGeQ9FQBgpxpGuhcxvifVW3emXXMe
1nTumix2j8lAJiVH003emKBb1CDwiv1FvWsPlxYIyxxDJ4/ncAJXWrHPUAve4KyY
RwJbRh4jVdm9BVeD8KInc40Uc8hc7sM6DNOl6Q6uye/J3b6xqejo2xUBOiBrf7W2
D80viIXrZjB6oSt1zN7Aciz8EklOKReIXCW4z0uEBUlR3svpq47ydzVafSlF/4n2
inc/NJte0gSoMyq1r9UJv+Ou/FSkXaMFuqAC4prmnqjsmGVG7LGp5uZnVCkgXDFF
t3L56sDtzQrs7XnXquC1ihpnZonTNn0rBKvMXL+A9g3t/Ojyki/k1E9lM5WMDk1d
9zDb6RJdQ2FjhTw9Rl86hhIlDmu3klJwPOMSSeAk82oUqZBhg1WEKmKhhf+2/sfm
B/5nUFnB1gK/9aTz1MqmM87EuRyiUFFz+rwZRZtuxRwH8xqob8hbHF2V5wvtRc24
D5zyCFjN6GWkYaHiN31uH8zG7ZhA6puoo6bmjDFvlvWuWBVmcJAngyPLQHNAQ4kH
1EVkiPtU5DK3+497tv/LbCj98kbp3iAmdYlWxLsTrLyiMaKdqPVW/7tkUPPDJ93A
uJsVboEDFCsE+rNHFxu0Koa8Ax7jQFDgAp+uHjCcwwGjZXPbEC79G8Pipa3ayZxY
08u5/BgR/sOYCrqmipPc1heVlcbOkrKEP7Z+ojZU/Xl90tAn6u/MJr9mg9ULNnID
tYK92gbay9PxpAYdjV1JN/gnYjLAmzMVtkHjYS+hus6f+dtyV4L2vTq/IgTQqMSJ
iWmhJ4cUVvTfkIWbV9oVACRA9BKpou1QDFQjgQNlfFZhBIUrsrHGosZJI6mM9hLp
wK5Jt/9othqW0CWsAlLXziToCy4bSo3dj1gJG81iI/+qjFco35zwG/ZSGxJwko7w
c3Fp143zBMoZf+3ubtO/4rSZVUEVC63xXn+0KeDneKtHxkNe9m1LOAgUJjMP+1WV
u03c/q2LIXvlJuK/dOQq4qWYjW6VnnUtki2NkROGxGe84ucjCjRL8F3Bw07z8Ni4
zPnWgQPXyOUev+Hv3BmPABvSZo2WbIq9TG4cnhIhxXmkUERxQFmMaJPT8q0dJJYX
9MOoWaaHqDvwmHrYLyMP+t4OWprxDNOUMtiy21SpLm4P0/yYkq/rAt0qt5l6rKY6
hO9kE1HTPSYZ6yvZh+YjnSnEdADqJHoNVBn5DBnma6MkxCuq3Cu2t4xnODPkuqMS
Np3+OU3RYJLh+XdQiclCsCvNyLp/kOUcjHGxeLDsjCywCVNURlQemhTwsdpwFlyJ
sdoZkcI9gimzOtbvYhR8D2ddCuzA1+zdYmsWOrxhxYYXP5t6IKzN4gQGZvg1erc1
xTJd8/RxwR0f3fvoCSsOE1Hj6+ZA1eeD9EASirE0CzS2+xPunC9eLJXnlVpnIXVG
M5ffDZ9nwPaCnCr5EkG+zGOSiT0KlZsJYZ/HtqOoNAvtq4g7PS/+2BEv5GjUM+Wa
ggRv9ZU5bphSoUwsGPzx3BbGYUmMqtEyC6JHnNcRIvDn2Pn26TxhCZE1S+wshKG6
+QSgscU1m6ofTt+K68NUw2uNDLpujwqaSRvKlDBwlXKrljfC2J6PJEn7J91nyxtQ
TCZ91DP/eL3oZ+ZW+W0qISuOzVlu8FbQReBp1gPzcC5km4DMp9CjiKTnEcEjc/+9
rJb4hb5jD3mJx9k1XeQFK+W8DoSkGTYklW5CMMIyXCLM+U9jD0eiTKzz/V3DA9Gs
F3j2XfDOKO8gArT/jMXPvWzVI3LQcMUXAdi9raXGpWB8NX66SNAWNYNPg9ISgsQ7
vOduNOsgGiwzW7VbAQIPaMAMl5eGAPjkH4sQjUQJiMTenXrSmTCKAn786Vz4nldQ
2iPjYgLbnmC7wc96GRnptSmfsngeXfEtDgxQxLUur660maBvyeX/yt0f5CHt67UT
bQzQGgjPC9Toxu0xVdkxPlBeF3tu4CRLDvuxHdD9tKgmAK1GYqLdoyyfBu6iFvOl
TOWWCFfk4rmBBhn3x7wNLjmQwiFK1CysxQODNn377QTe5BAWARK3B2cOsEHOv26s
gzGfz1SaWK+4acKpAAJb8oa5otBwRdM8Yfex0WOG23vDUOQYkXCFxOi4Mi1AK3uv
23/mPS72pMN81tXBDp5rveJO610iv77N2hAYYo98GSvzvkXqQ0O3eawzm6k7/qOl
r/IT6DScAQpL5fxZk9kB+fimDq+X//hCy4WVpTantI6AEsqxSYdA9JQxMndG/vSZ
5Sbpkj5qzPRFq3gkk0dx4+VD+cVpEwYKzCNGX/CN5YPNQORQYHFv7bLf3MceCwST
5L2gXv61oNMfCI/711DoC5vCPvkTwrqXlPrODisjC1yzxgyeyVJJWJto9fLkmvvj
UGWWqdSLPF8GG3Yp7jickmWwb0xO1QkSZeRTJtgCW11EQhRyLeIFEIgSNlbjpUsB
FntCvBo5ztuOEJn5FRoBbwDjzY8znpZTmlJambsiqfkgJvpsyieADsl/NXSfiqwp
uY1SfHGi1StSAhd25vbytVRK5Mirld2+VVTap0pAz1yOJoZpMjbHlTIxt8Xse5N6
UWjxGN/rXBDu7z9JeheGn3T0XjQ4F5UlttbF1Ba0S3lwi0hfwrjP33tA0ZykUM8G
dzWwLVlozCM64LDP8owwqE4MzYRZ2h8C7KgsRXYi07FaYB5p5dhLkHeI+7Doo5UJ
gjZjATiVL2i38sjIMp9/0SuXhPad12OGyocIy7qL48qIDglZEv62aR5MFKvfKdfe
T7Xqykq2jMsLigKjM8b9gvRD/Xz6/dbhlDcCJKeI73uIari0E4jFnlEgQLMf8vO2
BuCnGx34VyFnawBwRs20xv/qRLdqG7PpwXL7ICFPqQvUHJ0d65hTH1dBH6Ow9FUC
s3x00LE/wdVSKPTzf6F8ipqwOeftUcN25U1JkA4rBvyOfh4a/p1R6pVZNbC+O0qo
GUU49WyhDzIDv+kA5D99BYNkpbt+dKxn7k8v5+KZgXyZcTsgz5RR6o1ibVnZ6qTg
yZ5e7HC19MowBFMUQnhAvnSE1QOrbY8fNAOZA7kn/7MLIrBKH2HJJUGHxf0h2usm
d0ihKZG9lDMyUI9scl+csdyXlm1gZAoAwJ/E67oAKbFibdesQds/ke1mJArYP1np
lRFXLU2ASajSle5RfQ43X9fR3ns+iVDkH6ncoeRV0MQ6vw3ZCaEff2GwBRwZD0BO
j36bup/mEXdGCuk/vm6Mwt3e0bRXQeShI0/qHR+s1DTeRmm2xNAW4Q9zrgPINFC7
FBGUuIsS5aT2W/TfFHKHB4T97qCVT4vEMzflBPdhiH1UGFpMCyF4n/d/RAKu2Bll
An6HHEZqh7Jwpg5RqXEuDxtKPS+TWXmp5PyZC0gSWznK0X4ptjrtRk2wL2OnQmjx
11D4DpF8zgprga4GqkalludywAFwyVkHFYUX8MxpLuATkayV4L5B7gL0+J6Ilcn8
tf9P5qShyPzLzOyVLRnPtB+/rjPuGrqIYzg7Lf+9FxxqWtZHNF6/G3M5lCD/5Sl0
nyb0MXEP7xJ1bKxYn+CVdI/60aaVtCn3743WB/s6QssJrZFKOd0xcdaQuP/4OEC6
OMsy/fu8BlLplA35Ifu62+hExi4sbyA8wLzbBXkIVbro2ebZ2O6TvyDCo7gRm7CU
Aa69M8p3b8w0rxnrn/hUxTYeM4TcSkz+nwSxKF7VHZ6VRsSseXSPrlTD/yOFkb6F
0ugwIk04VVoaBblfu72kf8EfGCQWpVxfwJR5NCqnhmqY6WZ+8t8i5eIUQrfptgK6
4JvisEwIukthTLCumakO6xv/U34QTEuCOMOVAbG/6VDD/h0qYtDGjR/sHBvt+Y7v
buaTAvROiN2bjB3sek/klj8ToyvjREk3U+8xbc/bA87oYQBn0tsOft5wg70Lf+mc
1LrOnj+SdTrD1OLQ2Bmz4yehbb6gpR5mQrgyys5KjpAs/wWeAtm5APY2QdOCSXK3
xj2LKfjvKGTqhhdvfpu7k9t+f0kQHwDoSFJd73yTZYjXt5KvBcNyKKfNU5Zs/llD
7GZsQq9OFHuwCsBPIWB0bGJe1fX93b4Ll3G30/uBhX+kg5fjUwd5GyYl2CcphVND
tFDPiiYVjxzPpEV8u0C8gOHbQlY1E2GHIJVbydNCIvxr523/sNMlYk3fL0+48Njw
yT0BUCkTcj8u6k9/OveN6Xv6rDcZP2tYO82tAsofHBsp5gSyjT8sbATJ4DeFNWzg
qmJ9wy05W8jfkLFHqqakVaQg+fEDEBW+OdXIQhyxMlVlmD5Of3GRuOS3xpglQpJk
9M35v9CcD7nskh1WdvRRO1o49XGDJA6i09oXVoOFvMSk6DlqpQ3dVYA+/dr8Xaqh
Jh6XhAYh2UoprSd5uN1u4QO1lDqZDEwBLGRyZUyTE1euQsIPR/sC+EoFN3dv5leG
U132BwCCAiwAfysdaBULCSYY7vuuWPG3DMygNF7Glqfr36VklnoQsXX/p1vRBEH0
trk+ZV3VjSGnGyftorpVqzxtXoENheGYn6ijroA9Kh+vd8rJYLkKOXpKQEfbYImB
/cavZIzcg0YqWy8rew5DDkRWBtQA3ncxn76SU+tdJqaLbgqh4XClSP7aBUHVpcw5
72wrkmx9aTOSl7DyR/Gk8BsB+w3zAjCd113O9qvHofhAjxsJbaEt6pnkeNX+JdUV
QnTjuIJemclGwndSwHF9vqK6hxKjewJ6BPY6Lg3tCgT03TbKr1S44QLmQoswXpv2
QRogsuLU00cSkTg610W7LOiGHmIdZbO52f/ADJ+yU1wjIy6MhVOXQRbaQYnWdPn/
BE0JYjGn8YwG5NUTo3HBcbqGG/thpd6t7bKaeYKDHRXqPafqqIh/FAL3EyIocq+N
jFw8z0QnemmWFU2Kd8VFo+y2sK0+mCTXB/SnAmy/vXYhWFviFjTAuuwFXLtyZMOl
/Hi+QdQ24l8u/MmSctx1Mib2ug6DTkcLNo4WWePFS2w93hzox3DjrqUzhGkHk3MN
vpqgxhB1vx1xYcJ2XPOc15YZGdoyNG21G6nNom+dG9ufxaMfnU+qHHdeIUdE8eVf
o8HM6HYwKltrWxLP3t9ShsvYKk8kbDrscFK8L0hHkk8R9gBMXeVK79uxV9hM0Z4N
3TLPadSP0KVAVGJ/nmj4mPTYJIqkqpVw3CkFASfR+nhWewBiodX3j6JsWTUEqrYm
72lHpbAnjwe0PJOFEs36pZoG3dsosqTlIVr9dgeBITBXlXApFTabKgHtjwa6nH5I
vqBMyAJLlvBqJ31HfsOikZ7QL2NZX5qAXbcTF0zeLHK5Df7BbyM3IS6CnOId+bt9
pDi0cfNfULN07M0MSpwO+RcosNNSEuxh6MmVWIzy+DHX5K84uLdjxflV7xDc5vCt
+i9ve/lKv5Fxdx0ceTBkv/JGTCTdZJUM+TqMtcHERgqeICayqT9KD9apVXZ8TSWQ
OeratNcQIEFrZXPOlVzCFjDKqAdRhkdyWzpqaD5kcbYX+GwgCtrLITSql4xpjG5T
hWPlyw0z86M0WfUb8QI00L3f/OSe2nFvbHG80BnF9arQ6RCwyTlfPQ0wj8/0zF3k
dZ0YhCZxVTY8+3XWiJmOblcsTLirVjwHN+NJLT0okbGSyuCj6dGIEe7HQkT6woBK
xPEtsJJ31Q2IzvDQokpt6F6eWIENEMX6YcvmYL0oxJkojWETlkZAPpPMBfc2kxXT
mss6ovAFob9Ql6rrlbS3QL8bf0tQlxYo7xTmurbhPI+/FWJ49JqKr0duZgdxjh8Y
4ADnT+r1hPTg0nuaczh0Qt6y5QA7Ar7h001EgglC1Bgjc4GDBydBjk4gScPWzCTu
HI73Zww7eO5TI1fPDvvIKpvvjHPcWXCPQsu69gGiP9fyrwMA7cFfPlWzRpDbKzOX
5diSQIG55Oi99eCmb7Liw6V94B0dKeOEq5cVhClFzmdEoAK3BUgtXMhLC4lgq1PS
SPH5mJhXcuZdtY7Kg6a9W/YkD18Ptc62tT6C0Z6W/1jViAyQjNQILor/9cXHrcSU
fa07tAOMTLTaiGJrSyYMP1I8H/U/pv3lK775noq9kkc1HIx1izU4IKtJdTGN8PtL
TYf3igJTY4iIctpWzqPN4PmZSsMlIJMSgSXyy13GtWczDqCLFkXtHQvW0royFAKZ
mD80Dwc0EWeAKICM0PZqod7t0pEay8Gmb7/xJpLcmCnIU63jmdiC8/2oXGcnjBfB
9m7rvLY0h9lyQt5E15WvJy+6RfPN0lBLfBGaipeHi4fM92NLYJbK83iXynuRv2F8
/4G3au37Z/X6ugxVu5CMEfRS/Y9pICegFAbdfI8wKrEd7Msy/GY5K25GnBySFXB+
8vm7a/uYC3b2jbYaE5u+tDCnHDolGPJLWsUBgYXHGZAsQSQ/YQiLo9mYFe/bFHfr
Xb5yslH5BqdQx489ZhwJCjvK9TOQRmWHn1rQRnzQ457FOyBcSWapkBEPyIT+A1Tl
d2UE2IYDaOdXg7EjlN31HMHevB0EzL64+H8q+xRXanch7ZhegPo9xn+BZsJsrrXp
Sz3buQVxsyaFsbheIfVM3mcNey7EHyRbKxxp6m5oltlkxWyutN0oLAxyX4TmtI0v
fo4uPBVvFsH+to8qtCBc8lp9jgC71ltTSvi87+zcIcanwhW56Pyb5CaCnC6WC0mh
ahIOxPZape054pKPOYoUAjaP19Z2vz8F65WEAUbGUQxXrz8Z0tr+8qwlb8Auyizi
on+LQdwoKPj7ekD3hMYKA6uJRoGswErYolqNAh+UDxX9rB8x/W0CGz7N6w/aOCeZ
+1FGFL1TyDK/NIG7pVLrjYSWwlA1cqxnxkZ8MZ1pRIqVAvcRtRn2u/PlAGwU0FEI
5Tn1ANiS53K1EcXp0Cx3ZYSGBGXCwlIWj3fI6NyG40KWz7ZhYV1G+q/oDd0+ucf2
ylYqM5wKDtuSAIptjt8qYY0S7d8qMV6kIFzrOizyjVK9dJoogZ4deKcL9fgjngk+
6TC9ptyTtm8OKk03ILDWtTYelhKxFSR7wtXXzspz5ciZ7NNVZ6uSX0Y3mu5ExUuh
SECMtnNJcviVpsQRi7OrJOFTttcPecaRBizWwP9WbhmtWC2OKmFFv51cYSWy86u7
yyUSEtdbryJUf+ofm4ZPAd7NYJ8UxLT0/CHxE2VEo0ALn6unTqM/DVTumbPNQniU
ySSqZ4xGNiXM3UusXoSzLRdotGj2FO2mHyvYhff31sWsFLWsyd6iMbhNEoASu7RU
T+lqyNK+QdOXvJTdGVPOQNCyf868MnwdaWR8nZ/p1CKL3H5UwJzUNfCxR323O3G7
HcgBJ+0LDPduZWoUixImV0x/7VyBnAQum7+kwi7RKrpJtsgikch8O4TOI9sA4hKO
XAEX4wtF5bt0Xigb9xdUJSR14yakTmxU1Apcg4lUMjVNKVcs8F3rw4vgcI+zbBC/
3Et5ABf0ovAEAG4IOuHQXpv94HoBwnEoajNRgwcmrRjynwZBzj/uQC4aHsI1LNdI
TWyqgwMlXORIVHE0yfCsHaDuxS36Fdb7fbmRwjZgT5G2c5wdcM5q14E/xxrE5C28
0muYKqcNYQ65d9XGZrMRSMgTbmbvjxT8hoXmMNaYpztZot4yAaU4wuacx6kSAjl5
N2bfemn2RN/SRMDtoUxLPNKlQJdIEBtwKsMgQG4q3rjpUkhsF38JECyDovxSKRtM
ERb/84x2+oqcPUSS0PZNNCiNCBGGyVxlM9qTZFc389lHoSfTO3hvehvkZBbXP0OR
L4zAdOQ/sTjrWEpImzU3rJRxd82rUS5qCySdO+gWl/z5nH9eLYbZ0Ci45Le2vmLB
VaDP/BUd2q/t7c5yQv9f5XiPFX5OU7eMXWc7FH9WrHZJ+qQRop5ESdTNc6EQVyAo
zU7w6jHqqSrnb6y02lcsGfDxxjuaGE/6qyYZgDmS3+R2kSO74r7B5gaiRiEYrRhz
KWpN+9QFPjd2ioxZC+xIGl/I5VcN8BIrkzUPvHjBC/v6OqBTv0ynBwE0mPc+cwy/
w9lVoP0eWrJO9+ll9EYe5ePc7QqbuoXwlN26eJPJALoM3RO+nGwZmSvYeJIB9H/O
ePWWdN0HUWPtit8wJzInFyJxh9h18/Y/aT+rUXmVzapmTQoosx/AKM29jquDSpF/
Kb5twJe5FFJ/0rHBZr/dISqMRUAlsjATY2yRmJz1ym61sy1mFGUJmFv9yLkJl22p
5s9iFwbkcj6kTI00tB0z9Oe2CZ7PszPgWIB5SWwWjWTka1Gp2+5Xhgynmvw57U3+
5pszapRV4tPEAiq/RW16pXVkXeNl2qPGePIk/kCztaBXZty+IADJOB+RiR96auG/
cSu1gwvgxS30QQVa1d40j2iMw7t3JofLgtdgT+AyDDS6tix4pRRnHGUGQQEJTFKy
h56m1jvBELZtpEaP2znrmbYfiJmn9PsHJMBTKDCS+BZhIbQzmAC8CSy47vzw47h3
QoLqZ9qeg2pul/2TanCJKfGOoVuw2mRWCxCVpwynsWnA+8IQqU1I+x8bgdlaCTTH
f3HJDIqZv/5Z6MFA/8VxDKDF7Sbigqznu5L2b0Vxz4lK26H6JlWsAf+bB7agoXNR
6G9hMexrAqr3K3vpL5oXTwzD6xQeajBXbgtPMqvf3BSHbsq1/623/AqcVVtRDKeg
Sllyk/QurTMBexqNWeLArPdi4IBNPoOcv9CA+GNoS4cHMa/K03Ghyj/GLRSbQ41b
NGdd8YJ1KffCXpeSNpjAPku+blQEOqewDn26wD1f8ivK3Sgg5xKuMrYk25CnSFzu
TSRkkL2q4isjrW+SvX6/XE/SQZLcVijOR1Dki/MrtXrk7tpQfMmOrW4BcIGtcWlZ
sa9/7gKILfoDCm54TsNZhXnxE56IDwoSjiKZH2aDMlTUtH1MBWOvAgqb1YvzPYbX
MuqEyql6ptvcpknCQnTIpS8mZTiE4GCGGpcyt1GgmmX7Al5S0zHT0wBX4XYwv3Uq
2FR2WrXN+/m4XUhqMXbHQuEbv7YqZDurYT02KE5O4xfxQQrzF0K442OtffMFe8nA
xQZH5NfifAl5L2GQin8SuP9EuO+/ozAn/cPKg83b/1JtKx4vxGq4oSIDu5LfiDgR
AGNSxzdIS6FAybRBzqv6rDV398OttPk5l/K7zdz2ckvh/0bRLK9XxINteRYdcq2v
0KyIFNj1+H6gY4HXfh75i2ySsXuaiG2v2B83dWlejJc6DIVkp1pO1G1N+FEVyEuO
IFMzwWi/Ax1tH5yn1JD2PrTc9TlS0oCZ6jrBI7fOIGZ6OxHS23+eZBFoGjbDtCNJ
fnR3qw4Ve13s9T9ari+dRyvclCOQqXJ5O0yDI1QwhfcpO2KW4J+hRZ+x/KtSs25h
vUjO3teXOzCw9l36i4OiTZWRdy4mXRrY/pPn6L4kWj7PtBoUv4HENG2v+QPlgK5a
8BwPNv/DQkDZfxz1TgHJ67e2gLJWC59fIBxekQ697aMXwA+F8gBHSPvtuaqmRA53
QwBhLBLVNPcXDFzHmJtX+IVHpGtToLtU5yQRzFUwfWEGm9qG3n5W7r1zqlg8ifI+
cPgshbKShvW5YJL77+inpRthq5VEf1NBlrVu+A/4OYZvWHGWDPl9JHzEaL2N1/Xr
tLhLNZ+HpJ/3GwKK6MM5lAKBtTZH2pqLuxsvVed4SiUUn69oTPjI0wPz8XSIWKsq
HVjLBKBIPuQsYZ7U6UUHjb22X1azOgdjQj2qzkoKf/WBDR97AUnI0VAOLkk0t9KV
IzptuMKKNynGpAxBSzoKxAngCxRDnhMaUofQKDbKzDZgrLcyNQfJYPNShJx0YLtC
XNJtRC5N1hvQKBYi1vuHBEixq1KgQC1tqQKB9LLy3YxdaFbfb54sz6mwEYFLf78I
neGEVUze8hmO4rQlpBRijTsLY5vciwVENXBsPFb1rrSTDno5e77Ii0yax1141N2b
Q9RXoXKlqwnSAgkRafxkfC/A9ULgcp4Q2u0tp+/VRrpTYXIonDhM7h7tv2DgCohs
1KYiA/XsapUoOn5aQ89e35yFz6eipWBugyvnuoQW7s1rBiZwHb5MB/LlIWgQX8yZ
iqr2v21M5QJJYAYBFroPzR2wxY+SsMzTgTvXfengtDMk9jeslMkTpBlhrkc2kIXq
zajjUALotcL0OCkOxTMNu7UXmk6zsw9JzgStB34PjK/S28WenZZPFzoVn4l6lF0F
EyDUSoEaaCpNoFDKe6OK8b9okleG1ahBEokAAbUjsXz3gv2QUYt4RELq8mxPPszQ
xnloIdIWclrBsA8gnC/t4w80933N8RXkrp/kwdrm5Ah6PYpk5ITOsze7dWZuLssn
bPXSfHc/MPydvwer25G+jgncRJAFHey7SNdNOhKq88ZIYLBqZtRLe+UEG+Uj7rIB
i02osMpYKw8D2nbEnVRI8FOax4XI98NQ8sQALr6CU449IlLgaF4WVrUty+NQbBVq
ItOljFDdCsq/mWMrXMpC2wAaZaQ8PO2Z4PB+V0Z1KwachQ2kxvoaqEbJsXC7BVL3
sQwyX7Ni717N2w0JkegmPFuOKs0IVmAQsQXjhd+M38v/bFHxAbKCB9Z+3UVm0LxM
n/bdWH2edeqNXr5xBfIAj1WK1VurSSirNQIb0/kefYOiQAqW4Fz7e7hnSmIACR4y
8ohosXktCHVzpvu0UuJgUO+uNbiEPf8u1MkOZ4dg9fkmQkp2nYTVgHjb1FzSSG4t
+zxBwlSWHGjW9RMcre9jDBmSD7RsionFDkGf+2ZLUNMiOpNSeI5lQ8YjTBv6brwp
7411KoohWE7ruZdnhcVsbhFQ4va8a+D3FqaQaZDL0xqq3TlZa9f34Id3+j5h7ZkN
827Ire9+TYSwgQUA6ip5Ywseb2hguqkLgVWpXY7N7o671bNssNHo06AdaDvxBjTx
sIlGnL+rxJ6mWISREF3iJdOlQcvLVxG0KVHFKIkeYnc1DbFQJZCyMAHpH6NR9+Dw
1MitEb5klGUH4UXHCssDiJv2R8CiSeXdQioWi77pfjbRMxmrQjrk7bjSJd/z8rOw
SV9tZ6Jtm9KYlQOdVjDJ3gKNZcu0Gd/Vf85P4qsvoSOIqt5NTmeIIWo4Xj4iIXil
7HThKlSjyjz8XpdqaAEBQlWLyDBClq4viqNlwKU+k8Pah28oYOGOwWMXmUOLadO3
orQeIZB7Kq02tbtbtKlrRJnzKqQe7g80LqNJc8LnSwpuAxqvMMxzjrLVPaji+CEp
GBx7ULAwnaA0FHZCTmrexcxk/USnfpuAk0aL+39ytNdzDXj+BBuv9H8LTN/pLOMC
NoTMm3OVu8M2X+Z2driHOWiA1rsylMqQDh9gzjLoqhQuN5FIONKtLM5Zfo5XHH11
zMERtlktFRjzIPNLnxIWHLybjdigKFt2MsnA7V/y9+Skr5l7iT6U1YPLts9qvRDE
B5tq84VtRLFsXB81pzJsH0445Ndq8uzJiABU+SN5jPYq1yTejQMb8+wcStQIWiAf
k5y+aWoi5lqetq8x9jUZK6yYokBBezuFXi/uzzbq4ymMua5Alu79yqEWE54K2r9S
WEosH+Z3kx/yg6PfVz0rTbBz0nnvI6QAWQ+idgUVKdSZheFbI0J3EtJ9dmOVMUHz
jAFHbz2tQq7ChtRvdBOlhA0QYcEC+eDAUErylhfFfpJkrf6nYc7GKmbL+nD4ud5T
SN0w73AyTZ/ccLtyGCiNMoEya2tx6F8OKQd1dqAcs0NtNzF6TtjMWsk75Wd3356f
SiTeKh3FZVGgDMnGzwg4oXKuK2IQVp6zfa1V0WHhGJXDcHPYGzt2RoPRUXuKQDGj
FHiqUtJmpqIF/ikYAEuSPEZPqZxUh+D/+5zvYJMFPNxyc1enJ+rvc9JtO8NV5o1x
U1sVvpmhOOyjbglNh65xJGuPNheCMK0Q8awRbQhxLXeJbEKTgJh5aSccdxKhfeqL
NHCqsiEHNGe++KSTNrgTUDYq0tB1BT+bVjXQgB0xRunkIhNNe5db0zWAd48VTdaX
Da+UBxAPltwzBGxFChSNcu0L6CC9Xby19ZGbqxeqwXGVGeiLK40iCySt9+wShPJ4
d2YA6ur7GHeNh7NDIMvwveLBplDUj5tDVPKOCrG8fjGOT2QuJ/AZo28OomsP9w94
HHSuK+5Yo1BhBf6KwGLZ2tDofqckaOi9yFotag2V94vk+kc0oF/9DbL/SxuhuSDm
SIVeve4LJ7VgfQOdLqtgXTuXNXcnh+oVRVDhNuh5AmTfhmLR5hGqhH0V6n1sOd4i
FiqKoTBVVhEBWYfBqJ1mv2kGXsvVoLuVgj6q2yy3R38LqO63lSmbPgY7haLp3FM6
zYi+7aUcpaQ4q1wkybCNtDgL+Cdejy4+bg/VqkhC/jkXvCOfP9R5LOQJzYTJGxa/
sH/5SRlqSxrqZy+yqK53P+pJj37CBo4E/PNCA9qwK1uoY9dOXQnzxuEfVPWd2zK2
538Lg+DvAAw7DUCGw+A18ook5XOL71JBvjldzK9io64/nkEI+m9xB2PQ6OXfIott
xLLoBkuz2Zi9A2/zvZ+7SktQdt+eTudrvan+ei7RfrXBdriVKGNYodVE2iyIkW1H
l4E3lNnjMIk98gf/DOXcKFa5GC7jeMmaFwR717CtACofQZ2TBl/fCh5w32duC57j
nF9rCr5hZlPV5tHs8+GgxZiAHS40szGUhx/rCQVzWoBj2bGf0G4zDGMSduzV1j7V
t5xpw2lwE8IqWITP5YdGJrh5Z7S36iBXiZFPRu9z0eYNJvcvecg1I4P9vwK2IjMv
PlGMFqaWxuoOcZz4P7YLud/U0bGJWS5y/B65xKmvdafP8+IaAiCBJ9rwKsOkllX5
BaYT2gbmNe8hhzxRfRmxjcMh9eTF3FQIOmPeZYyejAUAAX0ngHl6g6GHsbLKcUuT
y1L24QeUJlZ8ZANNV0W0qDf1DCGavS+gxlj6XBlCAjjxNWhdPP081DxxYdQGtSFn
UwZ8xX8z6Hi4g1xk5yIlyUH18QgS4sxNv13ghBei1R61mO2Yb/0tIzZOWPmvzZKq
CmcHnPCOG7Pmx8+/epgxPHTLSaNGHtxiI8gr1tfEiNTwzR1qgtjKdT9DgmeEnShx
Un78QV7GJkxOV0OPf/IFPwj0y+f7hCsroDOaT6ZPU+6m880st4qMxSXCne0LEksd
Arma4a1rqdjy4/lR25twm/0SSihuWzqC1/WpptsyFAWKeJ3JUbN64SSgCYJy4fPT
V1yDBDv+Mj5HkXXXeHDo7g3LYJ19+ro46j1AlM2EBQAGbqCkJP96oPWgXcwOEAOq
YBW5PD2nGN9chp79DlHvaadQpztAlIqZmCiFSSF74fogAhpPbwAU5UBYoZ9Yza63
+ueVHbPHb1j86yQFkrrelGrLFTjFSrboyXTOxGJCgpaLcPZoviODtj4JMUb+xqRP
ZYKBkvaXoHRPVSTJ5rLInynPJhqDmrKTK2Hf5n0JFbm9KOhEB6cghpfk7zCJHL+J
YP9hP0apQqRRMIzIMIijnoT+JZQo9NfR5+MlrSVIQIso55r2WSXG5xj7UrzQmZIA
AROXIVsux90CatLyJC1DGmdZTVKuHWaVatpPocTjQUxkGzwzYGJWc0myAKT44eJA
bf0QNavR7Ag/xONrfECkR+opNLGtLg70ez+ERn910+p1t9BqkcUqEYs1Rv05ohrm
wGz3wzPdMenNYdijIdzVmboFVqW/FgNw2F24agOQSG5uLzSdWZzPp5lWmgUr4oPe
naMpUbMiN9CnGsxfg2W0sz/87uCiytcn2QHj5frz/xurmwp0vkIwl5QaMB3XKkj5
gHfffVJex4vyDZPM56VtGU23S2hDNqobXoLvZ8QZNi1Rs3N2CS/pMwaxZFomeZEJ
lOjFIZteG+YpEcWpdcrefFgkdvGsA072wo12J9cVhBMvUumA+xijIIvhJQdFM1N4
fNo+HJ44TpwpLTdJa2LOJdPqqMlZ+xdYrRLGU1eLZ2IfWQExz5wdAhPoZln7AbNW
A+95rZPCLeAti9AQrJww2mAmlwUj3JdumwE/hPg6r6L11/uA8YRsZdrgKTYZDeNv
GVc4E7zvhoXUKr4rPZiAeFZ/c0LALivpA3MAdV5Sb2QMlhwlVlh/MksK7OCi4Q3e
cUTFPrusHoGJKl5NKaIBrtikTUbftCxZ33NVaaOvXIPO+EzAf4q5psWy9RAqFwe6
B5n0KX1l+B34X4oT17rYPQBc8R45RK3Yl3toEgmLQCb7kiALmJkLml4Y9RKeBZa+
8ZXhHo9j1Q5AP/pKdQhWWrWDewddelvzxYIl/agIRmhNQsdqW+odD2lAeuXDkk5o
tDh3k4SO/vnQpbD7L+fxgM5wlwnpynzNl77fpusbcyfFGy/TAhO2Hiy9XpuvUx2d
ui3YGv1G3USBhQQwjHiJ+z7vklqI5dzCz4mrv+Uw9lmkYRzL7DSZsO1wOC8ktXzp
Lge3ZiCneV8u6uOttbsqTWuZrRaBLn4EcT2Is8NlJXiDqysALY4rz7cW9Ykmp16q
o3wcpRR3hAvtZJFUKwIcMwLfU7cYldAvs5aPhJ7NogXOt4TGVNxaOem7ubHx/bVm
7RYjjpGRpCt9mDrZnxVkcBS2q9UhWMrQ9KNIY5sNoAPiO+mS3QBk9VPCkLS+vpS+
xqsYTT2aIP2XvuVQU4ZfRJbpQtbn+q/wvbKvTaCkil05uO3UxiATx6PGA4F6smw7
TeIaNhAbPUCpuyUjvac7sKe+JoeBCEgS6yKnVXcMEK4AX1QS/WBd0QELAqNv7ujf
ILhnLNtrc0RUrIhy9/dfcTCNIeZX6Q5Q7wH6z+zURPyjXY+pKQuvCWZ12AtghwvR
YERf1Lio4oX31Ns7ZV8HF282BnnabsRzExXxAPSfQ/Im+64oOjoUFa3UHevjShFP
zKJ6e0ClOuflQTVYmeV7z9EjPj/xOYA9KbqJ3sNBhMoKt3t29Sl7jdLL56GIqXH9
zoCLKf84lFKBjsG2+b8uejGsEyb6eac40OnpiciPLElUwJ2OH6RyZsXSpYFXLsX0
eqmLGDGdhgBVcThsy/NxpWQua8etQO0R15xU2ZwqH3NZ6M6lOuD1xR1wnJw4O9SX
+7svno7RDfAsvp1NR0N0S+xkmv9SM0r3YpjPu0cz5w8ZF5NcY7hKXLx4qUx2zAp4
Qa8S6nvYfX4tW5qaWFspyjSeOhw+6PGvfbsS9BFciKTsuNUsK9XS0gdA9zgSF8AA
eGPjQXvBm4i1pcU1fRhPHXvU7y+ayHBvn3qsOiDS3n4SRzVXd7kRJC4yonxgGJga
rJQeUAaEocKqwN17xR1CLEt/Ldj5amVcJHOQH29myvLW+I8X4foLEqAP8WDMHnc8
SLtKhIIATPhGE6iOCl8SF2x3sFTrlYTNTf+qTtIdxM84xGvnkQILYY2qXRKApUeM
wkYzqophQQmP/udEfPZKSGUqAxr8EqYgqN3Xk08cNLi4+LOGRj1aD0nUwiaZoMLr
OgqBbtpGOk7g8QNr4DAL/FYyXaKQ9n+E1MwWURz/uF/9zS0rv4oZlsjQnWnTLV66
bG2Vo/XABNIk5LQPFEXm4aUfBsZydYSGG2KZlv9eefVQvWxotO36IRkMO8MAfST3
/CwkkLDZmyChfribuw10DfffOW7lIDI+/qj0UaIEOImHDxTEilhcI9ZWTUSx3ccJ
GFDEWzcflzFdxV84p4o4VmXB7xJ1JUW2CpeLtzB3OyLcU16RkNY82SY9PokUrx/j
hRn54li+9TKnETSV3D6gqojbjtqTjpLOQS+lFOOluN7cPy4PrNoYEnqMxBD2nVRN
mKiVwXV41Ol88tV0FLF/pg+jsM82uENoUkuO19Srtf2WPGYyM5rzRZMhIMqwxVF9
+DrF4hnUU4qybY/+kgmfP0N6wcLepnpA7IP6NBqTWkL7r8h0eCyRjwhVzheKSF+w
asgl0RKOruBstmMkNpTsXOG7e4OyNa6GK3P1BYr6fft45LCwYXOEOVuvGEG4+8G3
jdTfCbndPhvaGoAsPI8QJQ0lAOqRMp67AbgLFdmjGoKf9otjaAZ5TebqOSXsJMxx
TyicaBJRUERja1i4/KZssvkJqzcBsgJ/U6HxeQRmF8E0armMCqb5ndhf8Gaf23iA
uIiHCqjypCq2UY6Vuq43ClOiPIwAcYiTcWhPKs7XM5t0oZbFFowKybpYjNUOBZBl
gC8EpSC5UNCgAyRnNMwBjcOewPyUkCQ/VIJgqUPV1BR+A+mov3LkWgBhPF6jgRNE
O2MtglkL+krd/SjHMEHrzME5YtEYvVhwcU4bEI8bWyy4sAwnsA52HgD8FDeeKG5/
hkLXu9uvzJ5Vc/rszxF6NPfcrTibVoNL4u4AinKcQjO3DIthulmin2gtHEWBSgzH
0kFGiXqrAPtSWNNs+KNGGXkFc6rzScIp2RjsXjAZDIAjvH7PcCAS7a/o8Wwcl5tu
qcMrLWcl+6TFitz4fMOIRdC3zlrR2eQ1mMpSklk4lcDCJk0zmLnmG+yDFRDEalZd
wPDBRF0yLJrigfmjV2BSv+ynPcAHL2xRB08ELC8uk+vB+DiIFz+K6wHkiJ9suxy8
IThNJAXjJzzbwr5EQnnGVefzH6EDEjI6Wih20usKz3hLtLq4DmRJBz6YSCKyrp3x
A+ZbDLteya4j7hmz+VW9hgptvKSBj3uVXvNwAbo6yPAatcwohgManCnWezAUHbmv
wGTJwOCLgQJCj7aiPFD3g060EXQDMi01N6Dtjw6Cs6pSXbukxELix+8T0IftQ/Ej
MqaOVoP6RYrkjodp6PnhBJeBiG7WAxs3H+3Ijj7800DIjC8q2HshJnFGJv5h9T5R
j7gkO+ueEf3K2d6wIQQImqidU0fEpAdVh/wsBk3rRsUYvIlzDbWrgzfUCc6rmWy3
cnwHedY4urE+yOIjUXuzDode86eZmTZuMkflAG/z4+8a4VLlvc7iAI10ThATYCSf
fm/9NZXNl5H3P+cn5bLSHxZIN7iKd0wUsj5pzwy1AobW/cDWyduZAxFw07pqn6Mg
D+G4OjBzNWKyOxzfUXdSH8OOA6F71xeAPTAkwegcXN41lytpM4MMkAbZeMIt16wE
ZxgnUocmMgdKAU7J+4+Zfn5xwOeAO5cQlMUb1bPJ1fzNGvq/z8Wl498vVtIUd9yv
zITtkIY+QhUDdGKy30+IlQ5Cq1HDAjBNvxF0XY3g7VvXKvGE7adF/iH8sSqYRohA
GBQEOyvtshvBgW5iWO3bxoRSyhV1LN+WNHs92PEktjTq5jed+JYHQxUEb9zMMnPs
6S1prTt8CJMNVLhq4Hz3nWYC5GJ18Yt+DQBcBO07caaNegrCoHuiTP9+NIKY5d/F
SZmp3DGOnl3ILra38FU6u3lLrLsTQ74y0T4Xa7vhnNfzwf3UCzHKi79/cu2jOtTu
8cWyEhCea3ILkBNDdhnwNmBs4eAvV1ZoK8swdlJz+zemS3EKVSvGWwF0jiMc5TbG
fdXXAUB2RCTfbkuN7v/HJKM8gxBD0NoBJuUXquBQYhBKikaxih+lNfQfbLhUmYFF
ADkSjuBw7iMA4Tfqn6KpRH9X0eun2NRr7F0Uq/AfgucYOy9GxPVJP1GjAvuGKUqg
lZXKy4E50gxMWaNH7g1YIWEHz1GQyaujEX4pU7xYQy5YG4jFmc/+qPHP0NeTmJmT
HWXz+8WSbOetjd1y2Tvn9ObXp6D8Uy+ky0Absk6sMINZXns917AaPs4TZQg9DfeP
CNReiXF69nE/aDQFX1PsZ3za8XJL5am/U3FyCjuT8JZu4i4mBDbO+6n4NYJClF5V
wVmF2eCeK7EIZowcoDeqEQoSou5E6FR9hzmNGooGUD6e3jeZLnqK/79rhbhSqBUq
gv6bngcAQkORyeZz3mMeZBsOYRHtPj/K6n7q2tr6GpkbmvK4ncxhdYLAEyefndwG
JgfbIC8FrHSkS6veUWt0eqlVdsZPTZCE7ZKSkQG8jgyJ33xZ7dKrYPdfaBYjlMNe
sY7gU8g0E0m1wLMPWFBlrUDeBGvYMxKyU0aylUClanuInRBW8NpW3yBxrrEe1lf/
cmGahnQuEOgE/kvmZtq8IDhoZJp1aC4q8lrbxzW8VNlJbNGt6WYr/giGhaU+xwhs
f/0Xk1nFS54LBeH5J5aStDdhMWg9HeiHo+Fgn5rwy1QQ/tl8ubeKV8MMEIRa79Wd
/ALeDjcJ1Engtirt+ibIqrj9MJdlXe/7n03LhfhEGCqBQd8Qxjmt+Pv9iDrS3g2B
ehVGa7/rlUXv1ad5oX8Yk9C4F0RdOTlb3OEryTZfue7JLslY+AzXdqxAucwH8uOd
Nm61E5CsxOYUwXpmzE+LIxZ/oyArUT+5Pv8Cua7PM911K5kGMNSe7Jeg9QwWuKQ+
y5mSSXnHSVvckM5JOjHpQc2pr2ZlfH5g1N4r8Fw98EZdFP0l/UDJpLwX4uOT1x3j
S4XnbfqTNcHAPhbxLd89glwqWqgefO6HHFLsm7rsxSXWdSNgvSosSMnVbn50dz9g
Lz8CAEjem9MhDd0CrQfjNAdbxcCvJCqrWhEW1/QZSpBKFeKfNMVwbSbKYzHmeoIJ
6TMjMYaRXV2+1S5xCDDcreSmuqnCfKvXWF4GPvaTMr3ofJhP9CzIYI5ZiDcHXgzM
63DJHjzcqLUQ9BDMmV/Pb4Wh29jnR956iwpTaKNra3dXHAr6NhTVcNXaFNJvJy+8
6qTez4QxCzOrI/XN68jshF0Ws3DnNZjW75aRwpcxz0F8UcPbJiIe36BgedU3RwIo
DjEsqx8Jetj2TjGDym1z5q4px4yQjuOHDsJzg0H3rC6qUqYb1EZlK7is4Xe1KXkY
hKoTPO+m4kziQmjXP9YBRXY0IAx3N5kfp9mXMCFasVvw07ZBnzkJGszuMGAtUTBi
twf6OkMe5JpZBXdI0MtxeOTlkKC9yrKz3YB16y6JL7VVjpa7PFcI7TR8jf4hjwjB
TwK0bDpYxe2XmkGqsxtzDB6+fPVmm0fua7ygLD9RYJtOknR8b3fJYdCug5TaUijA
1F3D4bUR6Kw213LMveGgb2k+MYQthCxFpkIjwelw5rDMCF+rzATTvQoVJjXdcWR6
vdlux0p5DTgPqg4+FnJz85IuXTOBZTg2zjGGi0yzYUM+VPD0I+Q85uBvySmZm3DC
9Gh+/lhilapohVcyw7PEtT+OrN6NpaQ76UQ1fPoGGA2AL7IQoplm7vrEZNYHFVEG
CzFyYE+dZi4mpyIRuJKVy8UI4zOAz7Jd3lIjTtP/MGM/5Exd2XQYPKohA1ZcW7ud
MKNuaHhBCWg6asOE513If5WizcFWkuMqnx1wGhGy/Ot+7A8asPN3uHv+R1ti0t9l
E1pCsw9a6uZApbifXo6OHiTE06xNtfTjWHOZz66D6AKPEW0LUHoaJALKWC6zzgE7
BAqXPdZTaS8WPdu2fP6Akofs7tTreMJVTXgfJC0VLkW+qz9hJQjZ/olDz2FLGumA
tzFaZa/433g99FnAXQIMafb0WwtO38z68SpMZZ21OvUHqcD1nYIQUREjla1KpTpv
1GEw6jKqUq5rS3aSVnqmMOIqRx98nCsr8uE4uR/psn1xPAsxcYIcKJzj6dY3iGO7
gG5FN2NcFTEqtElb3meV41pB0Zh+xhcreSGIPV8HGXjuN1pGik/H44FHtAHbQJVQ
fdytC0zJlxPZcTb2lgXECBq580CXKKczG5CDYuLHRJcTqyKtgR4bYkJPOXDizbP6
fhp9x31UE6X5wdGpxr8Htaqkwj5wTwPOBqBtpRaoha5QkuoqsT+Ittzx85+ZrSLw
Fws+qZNk72KUU3r1HBOZWqPEyubxtyxY1Ueprmc48LTgbNw+zGm1MhaJfggLAlWl
nGd5tPfxFQDUIUwLgszRt8FGEemKOz+aLbm5KvemAgeFRtv/wg/mlP+VUHUDIABL
1f8wNZErTGwiJd7XhIuYqe+amoj4j9G/JleC7I3DYsRIDKrIzugwKGjrAkwxkvP8
h7Cm98V5BHZhNYi5lncUbGH/KPR1v6rotqs7d2OwHPR3enDiT4F1YCLz2hda9RO4
zFO5ASM36Z6ivdJyae5sKyWwcrcG6Hhs7sWsQZW5iXC8RtUqhWAJDdTUn/zYKB7x
iDS2yn74lQdkFOlWb5rq1ncBtu2ggdKarf5bdj4+6FNVb+2iQUCBxtGJBGfUuTk9
IAGYkn0ovFJz1In7h4zYbpr3KK3vSBcqA5qkwDAxKPOpfkuZOJwFuTKTpLzikLQ5
mvdCMuvU1GhoeTaHGgtOvJT5UkBNpb7I4gwr1em/YrXx3cL6tYrDU7FhIYAA9wRl
oCoD7X1/wnCmEBYDydw5X1l+k9B0Oc4dGJOXEnq0kC3HFPJUgSJUSMWydeR0cfRK
jEml/VLESLk6VJwKx7zgVy+bVQSdbMNzYI6hTWQe1v2Z43COpznotCa9nDgPjHK1
H72ricTBrlR/CZRDevesKobn2cZCKBhZM3vVb2xjjzyOPzptkfCOTf3QNWhQ25gV
ezmEcRFr0xAzwecLgpxJxxcE3jXMm0fbS1ZRyEqCCH2aUKTwhoSMZx1gGqyC8wMm
z7DW17YpzA9jk75jA8T9kLQx4MTOOlN3Tg5yd0bgYXB3Gv++EJmcsS5BpybwSljF
sVH4sNo0q+YrUTRpts4nAOv0ekyT7pefTpzUfTDhAZM4kRoCm1iw62LpnxkcEuXF
rilHqkoFSSOwDetsMFKI9+Iqx3A7XiUFfda7hrUlk01KW+6thMex47EuNcGDj3gt
G05l+t+iP0W3jmRuhW18zMElvH2wYmhano2Cc11WZI3RjLRV7CVp0IKVZl0KOkSR
1CN1Sg3WMpy1bEMu4r8lmFN0hLQW5bZQ3xTgFbBORVSHNAPiMJNRwWjOTlfq/2wu
RUzZzSe6ZG9JOvorWJK/IUirCCAwIi/3th9DPK+TOiVz/NG58x3ALUJ1xGyV5s6C
0o1oDwSMHSVjOa0rBzW1RG65nVjMcicWvkv9SSWw+W9bs7kjFmUdtQ+xipXsBasg
Hdn/KRkmI9Zk62c9WgSzR78ypzWx9xuhY47KDWdkcnBZ6hGuqMT3rsT5wRi5BPQg
WgjsGdnmSLHsORZOHZAUzJsOa1ZKWJPeF1hv0uUerudi/gW2aDaP8uCcp0Hebkmk
Opct8CUYcUWvBsp7HOG7Gc0Hl1kwEZzNxvyYTLkROpGHIv0QJjxtpOEWDMnrfOA8
lY733JaM1q8/E2irmD+GbhxW65fh/tuv7ExDMpobPuRdNB9JZj+F9eAsbi60biaQ
OXsHo4bM6/ly/T/mOIN8pr6p65+7R66pymBnBEoXJ2tRtNW9faARpTerqc3kRvfO
2MHdKk4NYt+IV3GXc28bw4RkAE98WVIN8a4umgEHdOPTE31E6t60vAoM+k3rfRiI
c/9k0fN78tFfvX/PlsC8iZmySeisqszbDxkTLI7V/Eew9sHmDRYup021Wt7wj4B1
Xl3TLW98baQqywC8drN/JL6iu7CXMfDHmCcY2ceJvaH3nqVbSPWCK7V61VYdT7mI
N1FpTEmHSjgGva1oBi8ZpKOamIK2uJRfAdzAsQQxbAeJ+TO9Hqh74cffecHJAyDB
nE99TVdtRoRYfoytUd0nf1O/s8kfeNnk3Cav4sy9qv3nkKAZnOnZuItAvcTgHFVm
9MXulHTX2Z3/wf+4SdalaqlPb1VOeWv4gZWgwJZjoGKFEW5SR+yeS7k91MJRi/j2
b1temlETG6wSJ8IterieTe1d+1nf9ZuOMW6GWc3bZr3wVi9XRs0lYTksV+mWQ1v4
Z/DEX0nfBWR5gBtrGwa3c9B5Yx+yVG39cJ9IipH75DMag3iYuUpuwbSLIW8WQxDj
TaOwEKUEwrvHCfRlJiwcF1r1BRw3zz0jDdRIvJqReC58WKrL0HdoZhFGoKAjIjQV
omQXrZaJc9ohLRV2BjCIGA4SybKlGLfdIPnXmsfp8PKyXuPgHj82GmJd043auO3t
JfeIa573/f2uyH949gfkVgYgaV/s2BzwMW0K2DA5er178GMqMYvLkKiATgahTos7
2vW6yo+zYREeVlMhByOvoJAndoJM+Xwpo3NiE3pSAgIcfOJKe1qjsaaXvRHyjV5T
T5iPRbRVvWoCDNl553pHtCEw4C8IK1ALUmA+FSUThMfmbMN3xHdAv745Oino0VhE
csAsdfRWFLNa5K8SpI332mUH1z34COayhOs+4Eq8zP2VqHUocN8PNofkg6kvg73Y
l+JSN3QVxQJrEiYegrmsTR771YBcrbMaL/82pmzxTAzZCynsOAp0+qIJeyUDzcWR
X2sg3I6Qf7+QcfHjTfSREg339zK0EFGtDUxAvvn740Xlb+cDzd4a7ipTS3tVX/Hy
uTL8lnNJ6PmeDymdmQX+ZLHhs/7WCCBfPHMBh+WSSr32YBTy4ylP1JGUadHXTarN
brty34xF1PTaM6gKKSF4+FbADTauOuQkZG0hg1nEn2mJ6qJYRl694oPq7ZVL+F+m
sNlydter5K63kspxdGiqiMWUpncNDEZD3IBJ/YcuKFscUrLj4wQE5KXcGA3YatX2
4QjkSKT68C3b3LmbBnqnvriGtihIpYpnR1vO58M3PJuEwYG1wLYIHsjPeqlsm6qp
GauK57EY6xSnNPj+ZxA7Ub3VBqOE00HrZqXZ4mbP59HnQPYUjBM7nbgBeP2YiA3Y
6gWrZDIAJI8jUF8z4eby0qvpn5735k2/rn4QBuYTR3hRg0bAgEP+xx1QILfMCG8D
2G59mV+0os1xFrdVj9kzCnH7LhlXHagEAsWfCBPzyFtvnujurxe3LiAjhcXt2/3j
VFVU3bbrCEAr1fEArNoJJyxDSLnTFWP0HV8ffYhvFSXIXbfvkNCWASogq4I0rvYN
VMd5zgOkdhmhhvQHUsbCgzRbU2oBJQFUe5qA2FMH1j/Rdzn8N7P17xIWoF/gbHFz
k+O88mNL2rwjWzn08PG3VHhUZOZN5mMTIxUQ7gMFcMtAnZSvP8uqPY7A8KMHEHqk
/Y7twaJU1Usbe8hU3QC/id68SJwujfxrweQBWujbikTNJI6GJ6GYGClB7BFlxCeZ
vG4itIzagd5aWlF4P4F8lxChBnEQL9EYLdSTGmU/DtIZPGlxEAZkR+Y0PFugktYZ
pID6E/kXeIn4JMFi75F0+QtjsTtNfMsK2hLVzN//sI+zIoJN10K7owVU71BuAsSo
mw3cTU70zadDa0cm1oqymw6EPkT8K+2RT907Q0NvHWu8UnVteuRb4I6L9MCLazhc
B0wOMTU/oORvfvG/T2N2gCQ5ffn1iqLqAPy6/QOd2vCqk6QsVQQyKlGQuJSS2cct
JMI6dmUuBnuwB9DiberJmKfxKAi4mjfCwTmoEqcese2dmCPkjVVJIqAIb7HYfDHh
VuUSAGHSGtOjjhIHJYKn6G2j6zCNnwvmTdgFCDWWW5IskX4QKZbF8PyOOATympxN
I/y6wIMo1oBhWR1SyvF5eIBJuPGYHngl0+nWooNEgjSTf42j0kvnmhQ1yQ2zhASc
tUmy6fTlX1F8Rjm73ayOVh6D3Y1U5yriGfq0UG6OZQ+myFBCA/XRQ2B+SnAX7Riw
rqE8V3UK/Ol6tZDzKdxdjZAKo7KKa6SSOpnIiKAR3A+9kJHXYC1UhHP8e03Ws4SG
iU2dqt0jKtM/YM1mqDvTIiGmVY5CemHWhc8P3G/9pKDFWDxU1lsvtJog557tZAai
nf3Vi9L/BBQI07bmxSVCy6I/mERP9KuCBI9Eq/ep3Jdn8TJ0eNGBx79XPSbslj9j
PK+uQ7lillgz9sCEuzU2yxSLccgMzjDTxUn9rgKqzYw3TwBSDhJMwg8PopW/+DBw
lkwgDEX6kgfo2/+hhRHb7LBy5r8YTEFA3qZ2cedTrmPw7rS/xUOCk3GrOeajh2RU
2suYcWBcKkCRUktL2EWn0tK0WKRuVtcWf8j9W3Ufy238WttV2asKvzEt4K453EO9
hWAoJCRuNsL0H9P5A5ExkR0kQcyP9SeEVD0mrQkYbWgcVCRqDiwdFjXqhX1x8htt
ylTCjJoZ1fOANpbYE+42Dq/O7yB0/fRTzgpGcHa1+aWwu++CRZ2ZcKiUNTQqFH65
EWGNjOURQuwQ4zVLd7Q47ZBy/oATqpLZgjAHe4kWy9O9qQCBga20KNdy0d9ri6YA
7IJn8joSoJ1JWAgV9W859MQp3nhWclt1/riX+vOFopXrIO3lN7lQ/pdyoIJCWCC/
FasvUuG4NINxAa6AYUjKLnvaPeWDBtTQYS7NQpDqhmw4oDI280a3hqy5NxWRMI81
Ft+h3/ATblim0cbAEWUnp9bWc3e+Lo560rSCvW4iq+cOk4Gc2L9Vt+kddAxWHa7K
+b461LLdeWAAR8SC1lVLP0+myQaAST07PzGt7y6WmLkcqjNNxTfPSjG2aeVHmuSq
43T/HBFblG04IuuiiHQ3na+b6CksTObVPH75m6TZahyAIc1vIDaht/yycwLgeTSb
moIfOMXCMv4LPbFQ727HchnpFZZNBBOhysO9hrCka0pD8GTMrINsYeIjU+Qb/7dF
s+Kw3NgYvWsO9ZLUSUAvIVsTDc20b17iq/jcZw6EvuFmAI8rDA4Z2w2D7Cj+QrzI
pOSvI4CMHCE5yj7fjSDwmHtj3uNGrqlYNSoTME7xWdehpwz88rzvTxZ6sy8/Dj5/
+tVHkar/Th3RW65epFkJ5fnD6eLA+xBmDC5StdMU558v4FOa7PK/pw9khpYKNcc9
gMCRWnH31gmhng2oS+M39Fo6+AAyH61wPkUqGA+Byb9dwCAY/okzFIZ9P25XPa30
VhrXFM1kHzMlXZj0wKmCbpqjY7Zvgl4Hf5tMAIysaIB1rTwoLjxEAhu5IoV3SWD7
MSYBGpTodns6l2c8zphnyMIE2E8MO7Uv4yEUeAuZjYH9mFHICzY2Cor/hcViJuhD
QO12rSnmMFAS5FI7nWnfedm39VL1undoAXFKvhIb89lcYmRCGiuYwFAFNbmnhKQr
02JmVtqwfZszzSJAX5BzccOsUWDXk4DHIhDKiJvoXjMppgtGrdiJhyfHAkbg7NJD
0V+H5JZHv1qADU/xKOyKKtfpQA8mULMfnzPsuqcQy+cBd2nLgnK356QoEgQrcolo
7rilwKiCl1abupuBMzbU17iOO0ysnjpuc03uEvyj0FKmMO94YoJtLZ6emS2Z/Vpd
IBnYo9FCC0MaqV3ORWsuvqSo3SdiGWRhf5KNlAth95N0OxVdUES6wKLp3O2c5AEx
uut8V5qO/VikgKO04lq+EmGGZax/nu2pMJhKMhv2ITPRNjhhn/Aufn/6Om36nB+k
WAxmr8u5CKmB/ANO6ye2XEj48aPNBzxDkkC13TEU6YuMgqPyvkC/cRKE3WKBtlSf
Wxue5msPXyMOA/WmNqP+Lwo4/QHDHr6UubDYucBukwb4q0OFrH6OMjDHSd/YotDU
i9Dm1qeaS/pL0eMAyxjIVddlnFD1D7jMI69BmPeBjSObs0f+sUB9EUPcm3auwwkt
f/pEixKknCJTtZ0+Yzlbt094ZNhcofrlcbxRyKDXiyhyl6anJRztn4/nrwdofCdt
A/Psvfd8HBdZZNwOkUQRbLDcgV6c9djTcOEAogE5+rkdlRXlHnDEyCBlsxq5n1dk
+cwfc8fBLeli3cdlpGyLKJd8iLtkbvrnbWnvK8AFup0x3vRg2SVh9oy9XC8b5Ohc
4vjt856Bh+DTmyoYQJzI4C9B/vrO9fF6IbbZL0pl/SNkVIT7VOKV29D9HlRTKu81
mbltTu/RIxlTGICEXXCOsL8wfMiBt76AC9D3KexMeG8xd1EQt5FOUMHUa10lxyI+
Bdk60htcSp4mAc+stc5dgw5vJI+fVw4hUgl4fCN2ZS/SiqHev4nvOqIE/yv63kIW
V8CON6IsRvPrvYbuy19DY7K16KEsJ1kkIlewaJerOCmjas5NDKmxIlQ8nznfhmPv
g1eR+oEDbwHdb+1tMoGkfJAJKZJ5uZcmpbHJOG0wDQPUE7FWgub/gyG1UgPxrMjB
Mclc5tRUxytVM1QJORQI+DVqdtfNHUrvWqYcsc3OszDd4qZmQIhr35HXCCvOgegC
46oSv2JepwbXRuBH/ijnsAhq2ApkPRigAMh1qbNdq82YMoKqNmqIWY3oQhNhCl9k
blgHO2QB42PK2SDgZoEVRyZcoLOGsqas0f6TLnxqjQX6jW5GFd7QoCfn4ox0ktGh
vsW7n05xLhzXr0dOYHazWl/rAC/YMpjXVeWUfAqExBsjkAP4KjXeOrEI1t0c+nAu
1hSzgXwqoNmvJqSeGZDIJsb6yBZvplCl50S3+8oJZPvVBQvWWpUpr5gM7KUne31v
Ioq4+yRK8zHWUMtZnXLVi6n/w4vnVxXkNyzY1RBSZLKEKXaifL1K7ZC1ieUw6SSc
PJPazj1wWp6Ilj/ZxwJntsJ0fZzd7u/7LuGuUqshtlJPmwho+sJhFhkieyugAJ+V
xJuOPBl5PBxIjbLCf3/0O1tVzEiXJMq+6/p0e4myKlayVK8TcirKRCQMyq+N8WAK
eszSkbaRFpglyljnIda/Dd/RGQsoPu49cFUXxgcDZkU2FbsD0HMy7Y4lHsET0pYJ
jcybY2RPdcnGe38+QHxATDucQDlZBVlSN5sKnCiF6lcbTvbmvK4KfSbqMwAdnYcx
MnhVSC7g7LHpkyWHIYfLpkG1N1bloSwKU0P7WzDx3wcnweLSuHYsjSvgj4Q4WLQz
PiWVpw73fb1l+h0N9z8z3kcPUbbpwhMxv3/pbzOTVS9zWgOKvS/ZS0UiLHjmoT40
1FkInCglXYO66BK3TG0/cUxtL39ml2fAGayZdMDMJiPz418zEYOi2bpsyPY1Yskc
un8a9zFLnTOpigJeKgwWg0oEiSu2pzGW2YJyVxfUlXahjByTx//KP/Sw2N1Sq5DC
IQvN5k73ts+iyopvVCJgN3kWCHLzp7HrIy6J+EMi9CFJMWRHv9tZy/YP+quNXuHS
AmUYLe8G+p2aDAKY0VjD8lbT3eoAk3pSNTKGoU0N1nPTPeGbYjB7X+Trffwi7Agr
IN+4y1Lrl8D8UIamfTVxJDW9DsUfhnpDvS30GJEdt7HTVNmdKXuVWSjFRV7T/Fve
mJyZEdrYjOYFdE288ZFl1H6NjSn2z58RkTzIOJHrSDHJAzHU9/TxgoKTWkRNwoiS
LwyB2dxnU3JolzETwSUDADfWG9nG4SHljL3Cf2hJzRlwK16z/xl7lUdkqFslMc0p
gTW8BxVRXSfB6h9vPYsjA7i+deKE42xSF7xa58TWw897yO1b+o81TpAvBCWbynHA
+PRVVGoGHlhyCP2Lybb0PIUW2O62cfuQU9BjlrHEFnZubOxXveFhIuk6XWPXIjy4
/CyrticmtHs9ZTjg+UL4TGYiIUMXfhPUOBFSvO3eucpIobU5ACJS+2KltMpfnNYe
cLoXpVOv8n1V40F4cJA7BNaYsAchhrvIQ8rDWT7rIUcbETt3zlHeYtH0PLUXKKXM
Rnp/phePQWgmok0tYCuwVGXp2NVuHYpGHuNbuv36DgsYLUchkNf9wc8uTNxQ66Pi
uRDsTznTRGZEosCsZlaQ8XZ0LNJVwmADn78yAqDt74of6gC6N4XjY1Mga6LrdJSk
bWnGQEh4Jrr/NgREkDvyeVwkUhDOFZt1RaLRj6u/amHlkP64tiaKS1px0/RP57+1
hUAz9POHSgUmqBIAKk6sWZ+YqF5hvu0dQ39c1agGp+OJnyelIcronOU0icWXLR8U
6TMCYYS3s6OTjyw/YnTJBfHUi+nCpRX2vW5KJpZcmPbNDI6ZetayliWU/EIKiq4+
92kZD7KnqzYYuRXE1bi+XEaoLIKrKF8ESLTpodn+PqyXvpY1EJcLpTPCYSIQIlt1
NHm0erbIZQvZM6CGUXfn1GxoB9MaghLDkdvC/lzX76cGLzMG1NGPZLGGz3QEnmxZ
U/9CZSHfTMrMYXSormD1I04q/nGuWTPEExQIB4i2gwtwvBGO8kB1RU6vITgsWRL+
aV/l5IYsbu7JlMECZcDyFd5jyjGWrBdra3BDABSO/HmdSDVglRPSPTA+UVi44WRy
z8/Sf0YdA36jnj2y64Wjm68x6C0+U8tl4BngV9iSCrU9orxomYACp0M8fv+Fjm2C
fYx4KxeFgJKvkyozcp2MsNkVIwNRZFfBIU2EzGIcaTwzsYhXiqs6O8ELcWnsfxtU
QebDKfazRNRWNXBxa+pGyIoyjB97I15uheZdUjxXY0cCUVYvFZZ9T3Cco5tEfGRD
4IY79NcKz7ZGzBnCbYvpYc5ZgBkN80Rf3GTPFzX95CH8puxoPdVD8AUHZ5X/0o0u
FaL00fEUoewe6Nq8Bq+KC7mfFOYhNi2BUVMHp4EN3fnOhszwi/FVfpdgN+MrR7SI
IUIpykKw8OY0WPNqHUNOoM/nBnYbtcyuFFy6D/0TYxDWN2ccshSDYtML9D9sy8br
9W5l/G/pWjPogFACQtMuaYWikz4lCpKvlz0/ty332hS/MuOdlI3lR6dENTuDMnLF
fgNMxSA8PeBLELjyS6uvqSYB5wuZMXFw1lpvvLY+fnOztVo8Wg9XWGrDqZqp+sPE
BbneLTWPO22EraPCHnNZtxJgtNFkYxlStzeCJorZtgAOENGxW3UxTBdiNaYt5l0O
YNYKgIT/aFMf1frs9INsANAsDIlNv8qsSvUfXDhAbX/4Lisck9/slliM5Hx+JAjG
aqI7AsMkNyXn+poJxN10ovh5ulmzp7+nI0deUGLnXBZLPQHragpxwBWYjB3OCJx4
F4WI+V27+HZbM/yWuB/XlpDonN7HpJSxMnN8prL9i4mG7B8wjFbyNNexe1lhAzKE
t0ihImHsqZolehuss2PRnsxvZ78DIIBsKHyYdNeMoe33K2lMNvHnWULrsGSYTwaL
vaPINNP9RwaZykzuf+cV+2C8fDh/T9mlnbvwnnExhhcuJ9ZDCMEelTTikRHF6+tK
TGmfZmuToVDQc6V6Ngeb042oJ7+fVWRMu6i7Zf9UppYtP0W/mNOcxnuQSWU273uq
8iLzxqv2YYDRffSqPPn8As4pFm2wf2HknZ9qanbjvQVOy4yEZeBAaeQrQKlGKE0k
rb4Vq4UEluZhZGI1jshu3ffrBAUu8GTYHJFShi6XxJdXudN3WOkKSGRgIOjpolHB
DB8xj70MERLUnPAZjxjHi+eppkeB3b6clTUWdybTPY5ulolzcWlJXZla1ORIV6C1
gBo1Aelpuv7xwJ8cgE3LPAlW1jQbxCyKMH9kWxqkEHgOWhTZ4bgPIUuBYfCGjml9
rdJxV5pe/y2IaUpgeN6YegE3hgFrYAYCI/iMAZaRUv58qi6XtWrF1nF0lG/rk+Yf
gw0XaEUMR4SbedkcpGCC7nRc3PbgR+XfrPoLEwGRwUdbvac8W9R/77KnOBtJozcH
V0tTBPy4oFfKem92jOn+onxyNRF9bd5FdndfGOSNEikUkQD911d3Mv0aYWTOs6os
ANkTlj5Dn6Udwz6TVU9F++A+8b9OUj3Btbj9gq324oL+goXnpEp+2hsBRDHrk6s3
S5l1N9VG1sB/2XAaUYc/Z1/Mc3Noyqfw4NScpUVCvF0fy7v+SvStAJLuIjMOarO9
za909j6Vk0RsL0dw9/dHZdXkiFXky+zifVt2puAj9fsznm+T8bXw0G18GHQTgdp5
SGa0zW5qyDVp/4e1+LaJaEFf5f8TRVcFyBNaIiOmLnrwxFy6rNxHrLpQPpvJWlZ9
FXotBweiV+QNOWoh0I8LA5O6G/J5arGno0huYXnXPPv74rsB08eaSeO6L1I1S82H
4qUUk3VmHpFwTNObmKA9ULrMEDUiRX6WGptvbM8dAoMGmOffwOApCDkK0PbQRH4q
8Q+QokO/x3JClyMw+HYV529dx3PLjdIErkcQdrQ1h52O2ShWgdrpFcx1evWJHcJE
ntHvSxoDZcYWZQbnadCfGVWZSrD2nGtCSyMfrhRc7ip1Fim/HTD3YkBfvcchBJ5W
nuUTy+ITCkCOJnWNgiR/4BBTaA3kk97t3GA8ckkCd1qNF9+IW/OJSoSczafDy2Rr
e3mX4qsCd/i9Eig/AVuiTpR/YJKJbpY7No9gri/QBBZ7oJL/NfrTLhKRSNLVLiuy
IX8V9GVlrxqiCHNTC+NDnXv9xBkqlWBnk/z3NyAE6rlnFpGJwxnWNTaI/H9uvo6j
s6uvNjTKxBmOwHEdO/hO85/ICs1SFm2sDyjpCxIFArccxfrrzhyvcvXlK9VvQJK7
0syDb+SZw1gFI1z19YoplaBDH5QQs/8a8N/FgT/GYUQwSjOo67EjHsTQlPbWIb77
FXkK9sEbD+Wlx8546hTZ3159UstO5xGVRGuCTVQl5xUNKsOA7VnvU73LlNXBcpeK
m8yo6tnNNoHG/wSkCtHtJ7VpsXRHtRfMzIM2qU32C3fU+Q0+Zy3DtCn5BUZRSTQI
VnXLPrEo5EvxZ1vBJQfA/cUANEUKYaq45pad6sPqpWJX6Y5AFf21aojgY/9FOgQh
EF9GDKwYoHV4Q5lSSynWEkV8QeJg9LgYhAQ4AY3roAcEEfLLnpAmTlNGcZHPyRbI
0lLyhG1ZWTzUE4xLLiAP6O9dXnMgsF/6ZtZmh+tFyic/6NaINZ1wfMNW0BCxxH4y
Sn7UFhvg2L0mnjXD3TLTzqNORxPcK9bnA6NV8mzk/Bc0xc1+PpdiqUfhrCA+ehTQ
1FvowtnprHmuNEcCvR8n4TjhG57WWGaf4ROBaipVYAatI8TpOJW75pM/GAAn2SGC
eP/enfjswnK3kdnh5Op5RDHcqqkTeai50ILpTwtz3haroz4Tuh9sg6m5v+pbNtFh
lPBCIW+3dbr9JMYQq0AbyHzkhqW4Y04GrOn8XqsorvHWWS6gIxV/ehwKW23oxFab
495IEQSUdEZFfQO2enAK6LIlErJIvgwaLscTpnZLJDxJONHieRvUQmN66alE700c
Wj1r8PHxPfkwMWJtGXegxZpNNxcMYVvbXLpfXFU6TMZxe0mORgZkn2HF3XhOUVap
fnOlFEsP2No+HYynp8W7tSmHC7TPnzXLGyS/l1t721otwl4iKJMPTg1ZqJkM3xLx
Z5AiANnrQXAZUoMRoZ7BekqW0Q+SsZ/BWfgGhAOvQxKS811GpAMGWxGZfsFt6P0l
u3cKscmpEFXQoyUk1l0za/bZd9f+h7FoBH2wlOXneXcxWKIp9w7GYMpqft/O5PDc
fJM0s7Q5nMQfFaLmyABdXMulkuLPsN/X5THjjSwYmCuLZI8jz3ynXwU67keIMt6O
6M9iDGo2jmPUgbzexG6nhcFKAWACmGNi1fGBo62yxgIiWLoM7lJzU8EeB9lOLVlE
XOAl6gz/Cuu6GpAsQFtNWSiAWfTiuIuMTUajhmY9FApHA5VaKLci5+e4eumEGmWm
3+Th0i0e7EBQgfR26htBo2NySC5JZHOT5fp0/fVSr5ftl0h1rTFV0KN7f2ZE6x5H
NGZx9vSF6cQCPxgid3jQefSAJwVP7WeFFBeTQQl2q6ydt7KUcoULoUOt8D8R8OJT
7lOwyc/NcMcIgSjyJ4LrQ+77TdWzJFY5OZ+koMskcHaXicebuV05uI+yWOJBpJ4k
GwzjENNkBfEDCjdAPF/4TmTu+TcSMYr4+tlXS26YUXb9PLT2S2HwL6HZqUehrnEy
IK8PgudBrt5r6JGbklVU7L6aAHUHtpCzJs/0R1I0zlHbHU1f+DkrzEw6GDsfYy57
hK2RwsjH7I/rl33sVSiqHTCBxVzKC5FxSSX7e+v0g73NSPCb3/BWW5Wh1wdPPSiL
Z7rt2EPfB/875PQtyD7nLOVzd8iT0kQYp/Jw44zIqRj3Eo5kVwp77eAa9rHQisxp
WmCobSW+Nsx47GUMtb3DJ9N2AlRC80Xw5aVPAg7Yz8EUESxrpd5t6Sm/JBcTuhdo
gS4A9dsHetZG/X/gIbs0iNQlMnttRggPnkYMcbwUEXxykPTI+/Wtt0wTINMzs210
bRjyQXo9V0x7XQEvnjczl08vvfyhgu+rdfg7nw/Mru3Z8mg7DplEM8UiHjamgvOi
7rzS1vSH1qH2vt8nS4y+DLmRCREKyfa/bK6Kx+FciQaN4y88ybhMkG/8kET68v1I
j5RAb3sszMkh/7e2MtVlX8rlWIBxWuSnU43oL77TBrRw7ZcVM0begMegkKaiPEfw
JMzX0opXa/XFWPaa6TVGSIgP7vMn1rlOI2Q5lCq0L+/h3yyjfnT744XiKfucSiuC
G8dQqszs7K3YmrdCq00T8pnlVDiGIL3gJDWdp3KOEkcNzbzdsmcpGh7zAf1vcnLV
JjNFrdX1t604HjIV1uZS3Nt4XTrd+yMdJeFAi4H2T7V5oeja3v4wzjp/KEDG7ei/
DV7hmKKILN6TXuEa1mkMXwniL1sTzgM7da2OgJhUYLKqlKdvrWMe8S4eoOJQEuyo
NaZcFlQFFV7xw3pMEDcqOhJhDC9bqXVZRLu+ZtAtWWEA+Vou1k2lr+OeBc2AZpdC
nvk+qalW811xQ9x6d9GAp7N0AzcQRhgw4X0xxMTdyfWPzf9dXv2pSNTVAwl6xXg8
hXgz2AAfjOxS/aVT58yTv+lapFdEum/CxW5KihM2YEmGo5vhXwwncXtPk8UxuplG
Q/h3HxPr8tLF6oHiDdcZCWyJEK8Do6AAnkPVd0YTS3QO4w/h60QxhRt71ypRTwA3
3Sv2ue3CjInJa5PVSWtk7+at07vx1DkLtNgp1+PqrpsaNXosmEBQuYp9wkNl8orl
H2XlqjgytJ58VuOW7jbePf067AifTK/U0twl0sv2SfCesT3kXL5xF5i32ym8jDd6
nvnZdgmcgw/k6SbwGpwdIrPZj0eQS0JHD8siQS6L2UMvekAHeMjgQ3KIaqaEErpJ
im9pnH19swo/mDxdPafHIEgk8wznjAjER23w3Wl7L0gVS5V0cNstOnGAHkM4PQiD
cVkHllt+uXa++TOLdV1aI4S3wOvqrjf0jFyD1BOZBuijkxbLZMIl8GMACu0zCdm7
ijYFFY27/TlaXsIaa1Ov3JxOFG7oGG7D3jvD6TZzerbUvl6/GFq85A/GW0x6hJFH
2e1RjGtkFrFMvxs1Cv24zEhGAUsUHDtOQDiyuHa6vo/5eQ1i2fCBQ1aahgE5Wq4W
jhi+VjsJk4jO8eiHs1Rfl6H6xvHkTZTqYQ+I8/GlK9iu5z2q4Bmllg8GgFYX6EWB
sW+MOHhH93X5rIob8LkeadeWxptiumVP1iKN/RvCllHmyvDKFqlfaulydkzjwi+I
WYObU7i4yi9V7HAC6wkcLfsYuHXF9B9JDb3VAnH1pHxV/YNgAEJGqfCLa8Wxm99k
liO5vCwGuoOdfnPdpTDVIWxFaL66CXg2WZXfuPklrDYsr/xtxivLiZFmQYKmcRX+
GfdOp4ukb4zR72RHgvdKvBdbQCQ0GUK3LQ6QZGBPRKbHffwoLE22lo420E4LTHOG
sXDqGtTH5OeTTIOWCgbCTTE9f/kQ5R7hbcufr80IOgt7MGj8ImAapHT2lB+JLHFJ
e7kmaim5cx9fZ6mTZqv9KsuXHXZ3EfzZufOzRMae5u8mVhxPl08vGoMmjIuUiXk4
7KEVxfGlVaTqZTQFoGH5ZHRT1CNZEZDma1gXiDGXWcolkssOxJLcBo2QTcujfaub
qX71P0XW9PsM75NKtM6kwnTY1zuiQ1+Q/aXoo7Yke7B00oW8d2Mv0WxHXkwv1ZKV
jKK7RieEGLymtzoeAJTpzeDt8qxjBpS1U5GkWf5YvTY7wPs6AcJOKZDz8cBmV6Gp
kE+dSxj6xASA2sD3AZwCjiie7Tgk0mK6WpVplG/fJRkVK8gWy/1VnhlIuUALiEyo
E2J5Q4QnBhiFPbG+/S8YijG9F5z9Hd8fQh/Mm7MheHKZxmPftcSk36ijhi6VKVcG
TUFZMfPPj8JNb6GMB0wAqwm7CrEb91/mQU2tZrktihQfBj9W8FQYFmzlP8C9oJlx
00lN/9Wa92EtL6u1/yCqrC6Y7OO2pv6RNFIdL5KDCHC83Jk7UZfXTyGDmMtadOZY
PE+GHGHyXG1tegw37cPMR03qMoQo3uenOPBmGVcx5mjlmmnDV23rS3zhtn06bbdi
V3GM0h2uahMeTk4ELBSW/l3eZ/ebZSh2OdV2bhjAcdrbrjsP+g9wgtDB6dt+xRq2
MDxP01qvpHUJXp/YUt7xFOOcJnmYbV9iqfBZMeJBaHypN3hVrvaUOk0Bsa7GJ6nm
tobhuFi32BiOlH8H0zz3/ebaZ1RX8+Sa2Plzt1bILHKlQKeVTYHPWhkzPZ/79tX0
QYe5eIdSgxTtK+LTVzNVCoBYuo8hRIXtrUiTJMEZ0yn4HyXjpDH1rmFszOEH7q+t
ff5b/HSNtOvSCofzgLl2B7ev1RNrbpkm6SSbXHxeMuGC+ps9nmZNO+TtnEupInUa
NYmWFM62GBk9LC2MTWwfmvotGcXbblnxsD9a2MFujEF8S8nhJz6gl5tamk48I2HD
YTGhkdhWyAU0W0xlQqIbigiyW4kiCj/kioeipNfiqOPHM0Af8YIpckCpsY01XeuX
vUUEjbWD2pD0T0bgwJSDlOdeZeJfAbnZG08NbF6ia2SytXccLhFXgDrfdj2viiDC
nsniirOwjq6FSc4Og6BhXpLYLkxfoR81qjcIgzU7J7Yn7H67UKKAfNOoLdfWpTaI
lkwjfNS43hEk7pKe9nW/+bcOIL9UGgzsfK+43BgLfYoG86QJilDYHlaBfKxpVAjS
jG8eOT6refW8KxvTDo90eSjbcS3eH7247/WrsANmA1mazjmSmqaqrvBi59ghYTMl
ja4lEi20mPOQNtdwtc05e73SxZantwuMYRGNKhFk1wCpZvB9XMKmvFSOmjAJOrrV
OW/D+EBQXgEtsYxMugn375ctPV1S5ugHsLiG9yDKoF6vnuX+0SgkRpkLuDnIX/OA
Nw2uKi4Fr3bq+MINQJAMBpv3n/NeQ5p1U53vrEKmZUlmj3a+FS94MCEuHIaP5DVK
1MeR6Jk8r+YQvd8NFYj4d/6ihbuW5TXTo8x+XM0XzhV7ejBiTqh5ekL5lih99t/l
QIovqbMxarmrMYK4O8m2O8LEinAkI9gTPDb5x0UdRne54hrly7ivLgYFof7EFjf0
y29EXzRhnTBrRbSU9feYWHIzYZYt9C0plx10N2NDhqbS+FqWGIfEiDM5e12Nc1AQ
DtOt7HCulbDMRWjQ32fpCn1I4HsDHI3nVJC/Xb4E6YEhr+h5HfqJvQrpaPWwKOfQ
Gkebcu16TuA73jNCZH/eFPXyexKc4Nk4owUO2W1ZiEgYM/eqzcQ9Fhk6fZNjbMsg
d5V8faILUaL+BG7cx2/MmxwBtmNXgz0pV1KwOhEOKATez0020WEEYL/hy6X52bvN
gB6Kj81ZhISfidrpeLyOZhnTnW/2CETZkpxmKC1TBSEG70SlSIKp0iSVnC14rSgn
OktPW//kybdyI00UeKb1D18drKJO/oCqCDDrKEJYirkEaeCPEbDixwLeaoarRPBu
Uy0n3gYlSwjB8MKAJpMqDgZe+Ke82APmFWSn9HUKOtoM/eafFR6PcKpS30PQt/Cf
5KUvGtjnU2236LH4hexqfyA9wGRoTGzkcYnJcEDqo3AqTWosoouO1imCWuHReJIB
XkHXYYAgff2LRyKQoNyWYReMVHw8rSU/6Z7yrvFJNSnObS6w9mP7XDj1g8p3b18C
QLuu7FZ2nwkfl+TkqRT+pNBePdjtJG6aDJrplKzBMPTqbxDy2pbqvrPStQcCvsg4
nKOByWrsZB6tTvQn70+E7hM4/khoNlZs/oceZo+dwOHlfH21JKcNtPcSuMv6ZirZ
jzhMzNpc6rDHU93TKpxvEacMF1UroaL/xwurxR8N+nhyJxyS2RiU7XwL0pfvpeCB
eU94HS4yzEESN3iL3mQYVIuJl6Lp0o+DY0VP9EcRVuVSVHnomzlCd9voTxDSRSfT
PV/U4HF2x8pQRAEHvSGG239vgjHpDooa9sJA9G3oEHac1O6oyorAL1pVTXL4VdSY
bQBNDVw5Tnu+4QlYrSktmAr1/xt5egRfEM/826aQbt51SatsfXk9cza16STAnJbd
CkOq0n1Gx9xXSABteECz24yww8A3/6oYcI6aNqnje4Ovoj+75Pz3SR/bl8ktYTOo
s9jLscTuye8Sitm8IV7pRY1LboxDY1wK6aNlPNubTH/fMOuQzJlHpyvR3vcKw4oW
OA3Zb8aXDNwPCmQt9CiYLSfiaJukR6X8gX/lFgfKVze9qQUguTQ1bBWyMKmQcsdz
H85EaKl6YMFmGiRtifqD4NsE7slw+DHuf/s02WW+yKW4ImhoJvit/UDwvPQeGWZO
EVQ47uN46w1AReXi4q3wylEwpV+tqrjhxvaMRopZiFRfClJyyIcQv2w9qrnANy2m
/8vafua11SLYgUy3bcwmVGdmpgG+FL2nUb8DtRIViY4QlCGUjb0nt/bZwDiBbbm5
HIWLW8HMGyC1gf09PswRF5iE+vGwkPUCheNxXbdMbyotapcCmaq1DypVtpM55fuV
VGp0l60Je1A/jbeGktfoMaGcYErKMx1746Yo8IaBjHFSJVTV5zJdj6jlM9rbdSZ1
t7XAFmu5eK3yNV0sV+PJIoswUP4ASH8k66uIt8tjbEfmLXCs36O5gKPlwDMIdfCL
buzEpuBa7KUTNnMUSX3kX0TMpDU/7T+1nmxalShlgJ/i+n1kfOBQPo+8mmFOHxF9
MGPFqZfZ0G6yq87pXFM3wTjDisy3XFwMCyuD6I8qBj2E9t6P5gUH4O/u2Fvv1iyC
4p6xzKw2nZUHyrQ8Plty5BCcTn++hTIN2nRMxQLqfZLEsIS5pJdIPmh9bvALPPh3
535e73a0w98KaArZwMIqmHkckPzs72q0HTRrxyABqGQ2g1XMQMTHKv3efNyqpXEa
FaBpd4AJUFEidsk+Q4T1EjAB6G/YgDpVNgLzE33Da48KIdjdEp2bOLVvAzclPWsv
oiz9jOBbrTE//K51Da6M19YL8CA1bACE7chHnUzo4NgckzWFiCycg6UZn3Avs1Xv
Cz3jWnkaZ96Zf9lYgUNrV29jGO1szNgsx9rc9zva9oM+g+5s6h0qpp7ccKcDFNDE
CsJHrTPxW6YnT6ySaz+rFQ2eZMXl4VWjNgM1vI2R8fIAkce9peSOekdlNGnNw1xY
db58n8xfMdWqj1JcbV1/zHu2kYM/aYPJM+IPSwqw3yWpyRKLkgtFMdNOjzBTrnew
F/PRBkx81wvr0JrlRMwAfe7cHCIiadvPxKKjW6Uu5B3/nA1EAEZm9NMN+TuZz4Fa
1D0F90j6+f74qf9WYMw7ZS4nLHrbaPwc/qTjvMwfRD9AfAzkzViKZ9XKmsln8DNo
z6MgJe1ti5g+o01OyviigcZyfiqyrLtJCauELFZ6CJAs0yHulvmIAak+dSOkUfc4
VsC8tIps7IIoHK9eKRMUyD2tQxWZ0ZzIqGs5ZTxkqcIwgsHppp/eo8zupNjptfhB
vsaLTKdzITDCNc4Tu/Aa3QcaAWkw79pICUqw6iOM1mPaN8gWTAIZHs7/X036lJWD
KauaKH9F+MtEgsIEAt8GmA9HjpWX1OGfvR96AeM8TWrLJVkK8N1M5sNDhPNRPTZP
OjK82nhliZULGPwd14RJ66mVkY1dk8/SkFQCNXg8wcTppyi2wZAy67obqhrVd1VL
K1QkQkQt52d88GmAzHrlFXxIGecFavReoC4BjK7UBRbMZTD53EMAE/u74jqGV0WR
UQd0G+GGsI7nkJJwHCNjrLlVYChOBvVT/fusImbLzFPBy+ce0XEdjKRth5A/4Glk
u1QV17G9HSPP5a25OfMeCne7KRFh5vxgfpnJxU2Evjzu94udIbQlT9IYcAkdzBG8
8edhS/GJNxmCFBz1L2D0l4pqJRL3VP876LIGLSlNlPRqizUHMmOOKZTe3J0f/LLq
j2/CAOtp7aQKWK81YvE/pdQBY3hOJNpOcl8IeVVeHWZxfUtGedLYrQ8bY1qwrzYZ
qpfdekODghBFVvNFeheGCqylDhLZFgMIlNvdyrt53x6V4nesROK6gwbqFBaDQZoD
boOuYvR9QExDgvmd5Z0n4tDSA6F8xcMyVZP5fuEBIl9MVz+l2grKQl5aDk5LSjzl
r+wB50wXrVIjgG7lWXLb51nsC9damOr5+cvWyf6d8Pba71GBwhSuXIvv+15mHUmk
TpJn0/eFCiPzygkGR2MAcidiYuEkaUMGnydFeHb/AiH/WLJ0Ex7TRHEpMq8T2/X5
lOGyEyjjBgdoDmxsWaETkm5gNcrHhhq/2D4TdM41C7Il1iubel/wAZ7N9ujRShJz
RwIIH6A69yYCjz1b2oJquLvdj15b3MpCHerb1/cENKGFBpKPWN9Mbg1jzL5TU11/
AoIKwPkxRtD2YmF2SjBpI2r6y3uTyKWTANGItYBzrihomE3F28ipH/dUA3bc5gxM
M4nGTcDq6K2PfMgsRM7IAcB2p/NbCthoY0u3+sxPz7i58zVw2+aGwDO/iC1931x5
LL3DGY3T59a04VuB83K740VukxtvFc3OsKrsqVusB0kLX4Lw/v/mUpfxwC2hMSCP
r53WYUCUqu+WM0mU21vTR1VCagQrFDehIdTqkJcurxcTXpcaNVhcaMsAE4FPEuMh
fx6VukHWkSna4jqen+WrCXqObonODO+8k8DOcb4GUXgZ+FdDBV8qbqgVBQT/Y06g
3qVCGRMEgcBg2eVsAGvcWvuYgfmOwbbYSdxBF6F6DNdhhYgKcBal62KMZwBJ8fSj
JjJqsYIM4ffKK7gCcL5l6Id8EpNKI7SboPx8eWJsZJTu/zZcpNLfqQTKichAqMLO
LucKrwo30N7sCI89tjhF+4yU8O5AbA+i/StU50F8wjLYmpEGcrvCZS0uCwMTpYmv
tgj7GSbl8GSHQudVWq9e/3VF1VmPxQL3veJi+vheKFKsUBdomdAjnQbOXQzYLEln
kW4m7+A/LCSP+uFaypW9ilk7dvpcrRRncKkebBDfJRAv8FH7zlyjkBjcM5MG2TI7
y7v0Ga5DBvKbviX8UISIFX+926u5RjsQLPzH5Abn/Cc62R+MLCogfABM/42y9i1p
H2pKt8Uc5lV0sHeuYog0xqUI7FgtUOVkP90hP3WGKzuIitHCR6/se8JpjlAJUmlF
Ogmlx3pmPJz89dbyTH+v87WSFMMGpwJTKFHeicex2h8mZKQWCjYrAmXpjwoJWVD1
e19SyJe3OXYRP+jwSXyCV2/pvZRz9/TO7QQL0ICEoEwjIlKHSy3Wyc1AGE7zLutN
Wy/Kst6uxKoLinCSwmBcw/stmz9Idowsh7z7O0qgtCO1DUFdixLeXRW+TvelvfVL
vSKcDELoTN7uez7BvCRx2ox6hm5943Y8yUfGu/BHz8JgIYdqy/l1paL0l2Zw/tTe
uOGUZPblnwdDKRnGtJTlBSgAGN+kw9SOGy2sjZ/IKhrNmNedW/p+T42d8RfHwlvl
KXNGB20i2BycbH35CEnLgbQ4CxyaCISeClALbJXvWChHcMW9SdXeVTHwm8iHanwE
krn9hNs+WSxVAS26PL3qQ3IdiNAB8dPwxW4IFVhREsxsPT2r2owYbWgmV4HkcMuo
lzwmijn/qrvWD901V8cZVSbEX4Df0f0lJjP5tAStsTpTtCWGqk0dhV7SrkVE9ou6
4m0it3FzipZPKE9xBvcfB45xUwF5L+Iu3iK8RJm644k35aOKNjlF14MebmgT42WZ
n3nNBLi0Xov2Pf1GIFQL+FaTI9pa9ZRqEfEmtiFCj1YP3S+xjrdK1NfPYcal2agn
CS9DYnqK5dpi183hvgwuJ9eRVAJVB83m/lMEcvS37IDCDvNJykXSS+fazSTr9dtv
fvWveiJDKKB5x85foTDAsNTXgt3LeNstdoe8eJP9WA/XoCphUa0YwJy7qx/RnOfB
YZhOboGjYwSB2DNFEuFz2kG6S464qe6koc/TEKh1TOsF+pDIVrPVZ34EQVL+mYLq
0c5pME/k5yB7NM2zdBt8W3lEIeBLl2C6944QW3PU1+XaLEw00USpQ9yWFsvI3RkW
rbNrcOOOzmrGNN+kQjfR1eyt/T+G3spdPfeLtD+fRjXcaS6S8B0qKG0S0B3rfZn4
/VUgBXI0lYI8MVE/7kvYRcRwlpwDC5D4VmUqUSnrzL//GECTsxBWi3kVvHLHEBGc
RngfY8o0D0upgwDUreNAr7Z41wHT1jWxJ4lLEGFbkN/7ymuDIzUmx277Fq6PNCq/
aSYVtsPVjLg9xu9kECm9HN3xV16FcotQtifxZN4PajMhiUGyUDfQuZYkibNNT6N2
7q8OwMxCV8NUBoimtQObXkIZ2yW0MMQ+bgTQQ5A5vDmc7eHBzQUaQGZWj2OlUUNm
PsV4bvdabaUg/EDYOSRUiocXtKZhAqolI9VAFh6Tl09XjMaO/f7wXLdZU6HY0ol7
O5+7gJf30VtDBvWT+b8Z/x8lEFa1u6UZLrDd4D4KchKp76FRZwCQcpUw1lL6ibRQ
v7mmNmO/lPTgtWi73pSnaB3niE2fdgkgvZ++HOpEhlKJY/6xGiyOMJl0f08JsLXs
cqqgZXfkNGfBofOoJlItnr2l93vHYtyDw0ZgyyAAA4jWKoSLK8wvcxAJFrn4cqIF
bnMiX7iW6jOB/B5ffIasM8KF+703fZWgH280AhfHmsbFbLlfwjZBtNj/27K1QMa1
xj7ddFFIVHKumoNfGU4U36QjMsxo3dmAkZlYH/veIRkjcPfUg8jvUcsjGfti8tf0
0Pz4jFIrYmh+b3klM1xLiuJihgj6o++GnD+7KPwZltYAgBdJXulEkb2Ls0xAZhMs
i3nCaoIwE/ZiRMPNY1lBs7srFEm7xLzi+oZPdrx37n9H0wKzlgPqL1pfpSO46tk8
LAe3ZSmMN73agCgsYuthDAZtt9+uXEeniunZK1NHJ6SKuO23i6Wg/e65/TSmkdTT
zLDXc9UUKRR6fDiGv+/yDrUfB0RqGUoW+mMZcvC16j9GkB+9NK7BzyuAf6LW3Lrf
iBMrhNS3YJJJOLSKDt3maTUQJmVDjfk6ys+yCpSd+H8JBSceeEKGeWhuJMpkL6WS
OLdmjb8MXFYnR487k8rWsY2tWI4J3jANHoU/RFXGT9kdjDlWkpcNkU/xiG/iE89o
ByiUjzb5bxu6nN4Vh3Qkh7TKpxWmMPVW6sMpHzyAkEK+QmQIZRXf1g6RkKPoCgDY
aZnhyuYpvOORHLOe+oFbn4r/L3LPRDr0yjmkqg7XW2zwr96A1jtNVKQmHc6LLdXS
NhVTDn8VXz2Mi7nMUDJXoftMsgXYRE8lBIXZpb/WU+ImrghnuIcfVJVYE9PGG5PH
c8V2qBmsMYO7MglIE/nMzBrWWLR5siKCCFa96p3mCSh/vb7zg+0oxGSxs9qropff
t8T0fnjloVK8hCQFgYWiWUP19raM15SRjLVlbOuntB6pJamHjM3PCGWTRacOTjcI
TohwT7xvQLeGtpGQ50ApF1ArNc1Ra8R1G4qkiaqDdyCzO45qZR/YEXVvM6R8JJNT
O6rotCm39oHkUT4Bi8QBKUr9erLXaVwjI4JhcVWAyFkv1MVXSjYb8he3iboG/cAd
hLU3CP0ffZMIp1REHzAMK7DYFiMv5dTaYY+B1wR2n49IE7mSV0HOPkC17yGeBn7n
u0oWuh76WwK+7p40vOFi4qfGcZH11i/YpXwysFeS4fq3mKdiROyq+BZqqyNd1pmr
UtS6LcYH8zhSGF8+TWsI7M0xOh6uBZCImiU/xM3s/8ANO35wTMMeRnMui34k3VgR
EizXa2YI8NCvUUP0/YYCERMrQWj7huTr3SmPxLpjWSXNZKZ7kwIXSdCNt+ULy6xm
i7EUNQbh6gg12pmPhhfVtKOydxQzO2r3teEYgiobwml69YYsNqDPot+Xe7wLpZSf
8oC7EExKPu89SsSUVUk/f4Ya7C3BwfrjLZpJVyuJpDyMrgaMMXeSfZ/Hzc8TkQVy
fgPqQW2WNq8zvSWfNR6P4CqG1oMheVb7uxOwi85mWT3RFgOcmYZaB/50eZRltCSG
lZkJLLAmb0p4zerYrqNfzukNZVyM3/KCE4Z4jVrR8FmWnieNKo3n79KVIPRGlaGW
1CYLMmwr8bbW6/4JdYw+YV0kGMBNNZ2dbrLaMImJDPTbLMMlQuBh73ZaHdJ4mafs
34OEq45c7geHMGISZK7zJjc0mPFvSQWWIKcNA+IQEHQhfG5xQ3B1RVPh4UmiOt6c
7XbCJi2EYYCJeY3s+hBafh6cMYBdjnGFL1U+TVp/+9LwL7eArSLsGzWAyaUqlF7j
BR/thulRegUvdl76t8ZV3AXFek8oRDGHQL1y1mr1t4VF/POIjiBOh2FUQCJJRfE0
vYQEZWR8GjtLKxUHX8bRgg1vZ1Msa43pX7NTNDV99f8fVPoK63PYP4azKyS8Hv61
rM1TJRnTzsIQcVs49rKsPc3D6ShYAFbgPPMFffNsZw2Pc08bCQj99oNMmadOJRIS
i0ecyNzGBC1GDLZOCU95kXKnd/20c0UPZI65H+5n68gIqcKjXnKKS/JwsJtrm67F
pQGn9uGpaQyy53kCw6XoUtlhkGYRckoajedMr43+bQ2bSoyIntEnEbQbgp45+cwe
nPVUgyWBeFJjB2SttoF5k/aCtpi6VcTR77bFyXdiVJ0bXrurX3lAII5MeqRKPtuW
/Jr9dMDFNiqdRD1STHxyn1zj7LO/LrlgkMmNW/G4QZf+oPFxeppdYw7egcyBSWr0
xpihbhQ/ROKxqVsJZeH+0oK2bcaHSU+v9D51/2l3YVwOwPU1JnhWiR16IjsiI8Um
PvzWYNNvUrzM07sqN3yzvpBry1TMwiJqxynkMFCzbiqkWWobRgstCt5AmJoN3yiH
zk5FGIXr+Hm/L+Kg7f4lsVIkXrMF15Di7DKOVFHi7D/fLSKBybLssNHD8uwgokhV
/7cEozW8jZkwVb40+v9G9HQgZV5qHnNzGuOu6Z6hB1cqzX+ettHXWvVsNnzcdCa8
Rc8XE9i3utPhZBcLNQzJ07H1+BdZJSqxcxaS1HUMw6tR8+HQPLBkWIloeuixxxhU
X/9Gr90n37bwUCqnuUIxaFeqMyP7uXK0iVe3eCc4KZHbeJeFx3nmDeT5CD/naRwq
ng/UkHoGNkjbxz0oJQd6lMun/j947bxYvbmyCHleXJZw6fk8sWIqRYSjlS/yiyMp
yXfJITIS+ZaVAP5e1V1CyM/uvHffC26ts+bktJStrigzMkAJdESYR2ubZnRdX/6u
3mZU82rEB3CF6NZh69/QbBS0TXJSkunwjyaG1hEdosaACQSb2Chj3AIGLh5hnoEE
zgdf4HYdZdSfguEq1p3mMCVaaPFstcEnG/33W1SxHKUuQ3CbB/QnMd+YYIIa8B50
Ze3ka1VDOeAZSs8BDSqrKQHTrY28pIVHPHRA+DavbQWcrVWyPakn8PZnzcmD75/a
NMQQtFPyzpKynC0LflJ0d8VybA7UQCk31qx/M0qkv1NA1yfHdC5pZLb7DTrorlQv
N18eH3KPkJzHhiUDqT3i8YYhIWt8bLIFtBZ4/ylQHlCSCflls+rBjzjJhzE5CMbY
ynXWio0pXndZjMOHklTaKeueW9wsVuh+z/wHhWw79KA8s3hfvAwwJP4XYPrtzEgK
zYpxfasP/zeSlpsfk3LNe7FSY5U6pYNEOdamZVVjbd+hQVlybbTeoG39s9OyH7QS
FQCkjJh6EnFzS9cOypZ6Tgya6CIjNjZ8k537bIKl90F1pRhqb3ELiAuhEhM6Kefn
YUo7zUrUeJG2eVv5mtTHhovE+QokI1WYHMRvbCs3rR0+cqMdv3uDpMANKnytPP58
l1LoYPGLgfuvxG5lg1kyoxXYQF/goA2ptzzZgWdRozh//8dk6sBanH6bE1m5YBih
sGeKdHI1Ve1VaVhCydag1OvYgBkcbjQ0EMi0crqjMrWLf7DQJsRPwhunBnxCpR3J
M3TpCHDVhReOaDGHXE4fQBxx2ZYKFBLhiFi1MlrRDumx/l1A5zqHKN1s2VhOiSJN
ED93GEU8A5tleDVHAd3285HsiTpZ32YSJF7Ioua6r4tcZliQMZG6oohQVCW8K0Z3
AtA74XEZhSq1br4ixYonSiEIIf6PaPhFdL2Hd6JH3flj94ZjyjPAtTZr7eIrEg5o
QVp9bFYISWjOviO9oX6O6fjQrAfFd4f5MTwHBS+PBEV/K98qnT14Qy3Aq4CPUzp3
cSoslyBGRr070fqmXx0JsOsALdI94995+2kbesZn37pWKr+G94EONAylFZG2wgdO
+6KcGuSV8RkiSaCBF0vrtCcQtutPRYEizfRHZaRDXfFuj6dzhuIEY37Js5E4I5zc
Vvg3K+qC2BTR9UaqD/4Emj+Q64HZ1zieNHZF/FEHBfaQNqkk7NDAEVMwG4shJ1Bq
VDO/8uzjf5QdNZ0u3DURRSEV64xrA5vUULzspBx94y47N0PSwBIGrM8Awze9FSML
4NjzGuUCK/eu5qoV5TWLUn+2CuAPb2HDXVYL00uwC68oqwx0ZW3jiSw/ONo6CTsC
xZ1FL4ANFGc9MLiD5dSrFjcgxUyjH6zkFbJwCeyE5jY1PHdOYQoFnfmzmo4Vfjlw
DxEsONOeiypXc9Nh9pGPs82vqDpPtbdmmCi3f/Aru8tciA8XeqboPG2cEiQ3Rz7+
iOb/afVAlv9pL0Rtm482a6Mt1mdEVzv96qmxYyGW3ZuXZZMxH166wUfLcYccqqSo
uGxmP9Owy2zcmFr4mYALIXY89+dOwJ+wdDFMZmlrYmHMn4LoCpXODPwI5y0LU1mr
PpdzU9x9kOWA1PBAWg/NW8R2H2xyc4yY7V8cCSW46/PfLt3Ngt2gXOgCKmJn8SUA
79y1tHLeX0pak8sJstbVenWy+ehKl5fI7t1aD9mz4Yo4BxBF2P6Dz+8js0dSRlig
64EvgF+jfoiFJJo6i4ZHicGraD3YUOZsPxbYLjSkh02mE93n9kB6UBPn2tMvVej8
KzNCUcVo12J8I4Jo98Lef4S6moMz0VORbKKzBTjmclf2966/Nn97yH23ZlvecLiK
DTFIfjsCC7gC6W+duqWWLAefuP53WT82TMQGZsUUg6CnT+aKeB/jnrIf5PJikUF+
Ou5kA32yRfpztFqSLFb4+skB/7Nh1mwusW7KeY+PCfHYChDVM+G17K0L5tSjXONP
2mWMSHUcXh7wxc3UlD0jn2PARwdsiirARsM8oGgCdRU/ySUzIaVC7o3Y7bldxn5p
YsDElgOeP1/t1aeEWL5nURUlGcznF7vneAQT39pH1+lkBy82F0Dlpl/d8CZcxEJz
mn//PE/KNW1av+WkV/xXwaEoYZ0FVwtJWtTPuL74twlEr8IMsrNO3eagh6TJUwvM
IqyROinDdvCsMrlXwNVDukHPwcDTpG3Y9Ny+WRXKlmCl8+zn/17uEvaoBxIueGSG
8jqktLDGLPcghEDdEveLLqlSMXxNRtaLEZ5Rk1OedGvi6R2cXTlVnjyefZV5JTnU
veW8a3hsccWaYYG/4ipSHHvLMeWfD8Erb/XOO+IFK+U1RnMZ4BtnJtJPBHdmLu33
sf4cNbKXYA+PBfCXn195uERk+74fh8ajcjYQ5rbhGch8+3rfjEUYU4TQiSSxD4Vh
iDEieYmTbOIdeY4oRuVXlkL6ixmJkcMwB01bH5wTXLA3dzrZrVDgvNrsJU9tgnJ4
Eva67vjh8o5wVU+lUGr1amdgX1lXn8GQI4m/Vy9OygoCPHbeNSTrzYGB9yazgyu2
MCEbyINwr023ThxYljybpItAdkuqAUYrkOu5IR+l7MxeJmzEtIy/vEC/RWbjitzs
0v6FI5mjGkVBQfVmQ6Qs6FaliLAFLjmvyy3AgfMxsyY76BlkV0egnOURDKrpYkmB
F5JyWs+7JbrhsAOVd12XuSXpi5xUrCRiIQolD5VakCeVgs2Bh62zPiZ6NETC7fRh
O42ISiZXiZTJJx9vnQ5lRyCuvvMkQGZ3csYcfUtu19VHlX2oZmimJ7KJWmoh4Mni
ocK1XtxWzHg2SLHxTCi4FbrQREnR3KJCVCO6en/Jak14vZvbEWfeh4R1TtpL02yo
ENcz5MyNAvQUwIzVmORNjW4rpH1FTblvOnst1eudBnGFI/pFB6jFpZsO8rhjGBlb
Undcg5J3kJqQK2ONK5mDGY6KYmLt2H3/kMC3SF/I5shBW705Kli5UmFgh6YYhtrn
mIChVEwIsyF2DMn6Iz1rnjJ+1WyIsSZzkG9w9ssyyP7olYfcC13q5uDr1vNEMxeS
EXs5MRRzQ+teVifV5AHOAebWqR7fY0HQPX72pQvy8jHK/8aWHLMMhLezRJI0RTq3
/WbjXF0H33A+OsddWj8sKaHT2IOZ/1HGvIZp7TyS42/4O74UEj+ReyhFMSEY3c8v
/qcqDsP5us/DPm+Q0LLpB5+NZEGDHDfca17/zkUqBuo5FYFKUe4Z9W5KSmuba48G
umSI3+mdblwwnwZ1mCXqRrkZgLXa+NUgPyaWywnwnu2EjT9Qeb23R/jBPIzDJ2bY
9IJ7WjiaXVFzGJMJL4itPDtyAZC/hG6wW9LZTARTS+EOz7YGlBiN/6kbYyPPp+cx
y5jq1V3j6XMC9SyyVYE1+DwHtjcJBMsvtyrlFP9Vd6velsV7BB34tcdp/1Tphl7e
LqagFqHvLkD6/3fYWE2xLtnjTnn+S64IJeWEj1enoZ0bnJV6OxnidGSgibpBZM/F
TG9T//QWoiaUe9YLDP2AxUsvxd858cP8/WSn+xiYqW3woeM1j7RMSZy3MbZDXkMC
Uw7M3fEh8xxQ4ykB7w8W6QKI59wTYxaaRb2tCuQDJjdbnX3a+ztjlsQ6D5sD7OlD
NFxkp/kXprtj28yQee2q2V0zCcSvnYYNHixy9iZnzs2aPE/uTtvf3mKkKep6nUBG
HmglLai7ynmmtExA7jKa0kjKESBtWfjLvgSxkFimDGRAG0CL518c3Ltg+zrIwmAx
R9FiihjnC6VrhJlMqlcu4dJZKzr7xrMikBSdK+9Lq9mzNrA9t/ooabdPX7k1N2fj
k3qNhZHPISItsZQgoKJU0UiLGBW5IAt+1mVEdFDrVxc2dqM5Tt4TMG19CfD3hlFM
cC+bdQcR3kJvvE8a1TKitVlaPvFw10x5vrACOQ8vMmV5qY99Sxn7K3rPKUihwo0t
r4kwxcqTNK9hN3pk/h2aAyjq+7C8d9RUlwJpYPDQtOyPeAMbnvSMm9lYfq5/BB/1
TmybHbh+L/i2V7BtgLq6fTzE20i6/CQ9vVrvtIDNuQJpnkziW6+4kuzMhLfNna7U
9CR0G1HZxKFa7puxBrxUjX5XMgPhdzjiC71FMA7Lz0ng5PBhe4CRTb/e01kJurWi
lnS7jI3K66nDGdt7rNCN3DnRqWw9uJb0ZpaFyn+YpGJjd/GAd8UK9h+9uo43FQVo
SmwlJbxkuhwilS7w6UWpK+CbsUqRFuijPByLw98JS2Tnzc3PJQufPsAdpiL4cgfi
/vQBsiQcjeEnoVYN0O4NjKzuw1Yj5jAt2tTxldpOhzrfQa8h6kcydpi7eyewGHMG
JSHUlvU7q3XJM2CFd8zgaz8wVFFZ0p1piPjRczmRmX9oM+O5yGQaP5YXNkX0EzQo
NhMAir9O2y2d/Y5yyf4AGigXtNM5j59J8zooaMz1BGKcCbeAX++F8wdbXOPIjYOZ
1DcC5zJlJ0YJ3vQjnvqkPyQCDFSEf71C6OzXgPSHlwxGujkn+KBUbzKDNBt9SYuv
Pu1WYzMVYSoKQF3WJrVYVn8iAyyX9gPOsJlJgWonJ5tlwbqWVFvl3ZOzRe3HZITh
luaIW9ua1uJ1v5zFmNgTfOVP/PVajQMkOVtEa4gStr23jK0IXoMm10jk35+8tFjv
05hS4ToBzPUFWGvD1Qu70M0//+PFYuCu1hgQEbr2FEq/JzbH0A2OSRPY9srJTWQN
RtTdfm1lHTmjELWfFWw4jwe+JDy0kAVcBti4hiLpNI1lFfQw/J2m8tNi4Yas/BKB
cI65OBt5KUrUKjWDMd3kJK1liyPwFYAMho/H4/l3j99oHaSejtu49saY6pZIcjjP
uEdXDltvzGHoiPr/tejFHm/49UbAFh54NCwPka/ivimFZ8CTzFssf3U8nCTs2B1T
T9dvwj6mE7bp1Hd+GgNgiLma/4QOCkrz/4aWXzJp7XnGuZkpgDYRYSqDgPPjOsR3
zHh7OfJnBMdSeGoe9PAMzPy9flPrZjX3mbsh5DdQnbmsrukMKA9crWNcsFvg96Jo
tWWw3IX7/8MQ/I5CuqMvr6+tqUMIsv1a3EKUFo+WZ+q1PbPJzkVLZGoijK2b3cFZ
E9z4yWydzM+mJR2ZGAbrBcCkUqIKQsOaG2flqiWelZsMgxIiCYQW5ZGHSRBscgOf
ViNckaRin2O45vkC2NVJkEvkxrJVYtVzT2XlZHiApNK33qKc9669k6BfiRbdEMYz
dLWFmTf3HKJSwXMnHXUQAByDjAQRf3DXt4ChIPasX4Ap0lfOzJk5vB9Nlk8gp48I
LB4JNZHbuM9Cxv4proSnO++V3h4yXMUYB7RmEeyu36HTgWBmZ+b7iVRnvoWTf0Qk
LUxsRe6+IvKFHP0evKkCpR9vEO30NNYUyNMQPdTYROWpj/obry4GNV1eKbJiEax/
44xUe4Yf1uWFprARdjco564tAvc9FdCOrA6fwcOCNw+t/wDvXmoRfVPzHUJk64ms
t6+Ap7zR5ZHvszVvv8qVTa0SRmOwHuW6LAFmzRPKOAztnCm1LVAyac6t6m0an9KA
P5UahVeryrVgGWwRT9bqYS9X1j4qY5VqYoOz8Xz8JBy1yYg9MEiPKqhRfoLOb/XA
PEpiZw/G8sMHxnDXJ0j3TJp1wBZJE34jvIFANsr4CqJgnqeZ2ykCoYOsZ5oLcTcw
P1jgbAV8yFBDtVnRcUnIYP9j9OW0rFI96YsGPaBTOlHG00Gk/AHpAUlVBUe2gwvs
u1pcOiPPfg3UbJGdq2zdbqE5+wO6t2eEcRCotVKJoOEk9yqvciMLmf0L7NzU0HPV
n79zBp+9zoQ6lMGNUN5xl/jsDbqB4tXq9AeyU3JJ95tKhC9G7n2WbZUoZ+Es4qRp
py4FHn9vskaNrdXfjF0wT/gUU7xsgIqM9DCfDsbUUaBVq+GVyN0t+WJ+5UwBkCWW
70YT95uRV+j4p0KoJGQAyM0fr9psOCqy00ICk+KGhOsdEjeefOoqbht/KSSmEMsU
05wd91cuEMDpoSWaz+1bcxCE+s2a7/v+XXigJUOo535Wpmv5oqiSIzD5q6KPHW6h
TAcpFYKlDZrdnMPDX9QMsZIsk6Viz7SYBPq0Zced3pPLd7xl3QAk4DnIsgnpIpzb
TvL1sz4Yu5B0nih8TEB6XghAZqml70HQyZMeJmj9RMhpNDBmFR91rFHc5xfBB2Xu
MrC2/25aNStcpOfWqR8r5RPMkOyC7QIoaoIDufdcQA2jTwP2FCodXQJkZiSROonX
fytDJQMcO0rbuOglN+FZURSV8ONO1gXMcFEk3tEKNFjC9Fz3EwkHaIGbCCYiJ+mv
4KxgDX2QG4Nr/ygK7RCFGDhKflfjRVTZ/ngY5PPwlLGtNJuObSyar1wO+td44Tcv
tKcwagHJ6fDDQkCIBcknGjwpj/mYNGuhRkCQybQrJKZcpMK4k+iFLCE6c2dxHcOt
1h1fEdnwlABQQWvyr7jNRY9F/jguah7BxoN9M/bAXMehIeSuZTA90k7ptNtjS658
UxnGT9jPLMXnXPC2QuABFrtcs0Y1Fd7NZItt4hYpGzwUsQ3aSxc5/u0oUnbM+jsO
Sg+fIY2lz1Cw8hqjOGpfbd2LjHW3X8FfrFlbG4oYKnQlZvQ3O6piT4gDLhNGtA37
0NStIOlTTJXoltIKJHfWeRCNtbGbfUIP1B3Bnqs5pWwnITdf+1bH1udgBmRv3J5y
nyvbgZNxlezGaOtUyao/83aOdkbVlJe+FapUJMhEPv9zEr1o7R/rRPtCmZ59ov7U
g1E5ctaNMvrOpQokTPEKK08PdCJ3UKgw6U7HIVDRoskwgMT5j/Sh0PE7WtdSfyh1
oQeAcISS60yy3TNWJMm2eAp08n7AzuC5L6UxfI2oq/mlYbrkxYdoZWXdMC8gRzLo
UfYdr5OnH2RkDBdtHTfsTkot/UsQpSwAwgsY0klcXktI4zfVq3BRPdu3rmB/QNy7
s9r6A6z4pgZm5+TYZMRggr0v1SLD9cYeSZYq9M1dBKbfof2551nWlzdSCEFp4cUt
iboaDBgtAlizyI+8ypm/jamqQpZV9RAWc0fO/l/19wfNj4tDiXRgj5Fdw7x5divg
HMUCPbc5CxyN+ts3WIBtb/0pd+SkQoGyJZgS3Chz03ttFe6eBNjHIzvBcCvUM4Bd
yS5PEHEBmHBlavMzWd3sWHJ1vR0fy7RiHl2iAR3Xwv1NKMxmv6OM/5pFfnnIIn80
aG1QPNILalyfNVEKyrx03cqSf82DOx9m55dGNwSb5DdZUHYd7JAcJNITpXwy98Aj
X6xUDZzPJd9acHRt0xj3UG/0tGJuDtJaYcrNcLT3buWVCOUh5YoMfklLVxO/A8nD
efEEOictoMskA3ErpAZqS8Ij8tDNB2cnKJ+jqVjZMxZO6Q2xQj221GLN6UBAbd6E
Gl0UXZETPXTl78SICDKbP1WBnN7FdFdFP6sSrSsdF2N2i2BYt9qab48iG1LnQMZE
YqyM3BFGcF3QhNqOBUgquLuZ4iIouG//ioGjZuU6RUiAyxZvJSNeN4sopP45GxOl
AYq/cdSyXBmPMlr/naERdLcpe4uDuvgUuBAR9fyz/UcML+TgWwezldq9Pzg5fxt3
YVp/hwe+1rDv+1q+UKt6acE1ZBlMsSjh9Eehj1vt/EUGDWuYSF6W+yIOxBdtIYl0
DYrz1kAYahVmX0mxP7QT2rh11w/bUwHq5dtZWT8Y9tImzjDJLIE4WcKVfb+l5tGf
65G7I6ezWCGiPxWG8HINolZtq2y3iiFLEVEw/9hKVF036t1lLqFqF95l8aOtPiBx
jPKyOzdFkmERJsVQrULYE/eDOIqU1yWS9aNtfwFngkTvCHU1hJOjtIJijkmzIL95
E0y4a60cgHfBT1ueWeKo02FsrslRaBhrjzn3TZ3IY+0X4z21t3aUm1e5SVvoThPy
MK9Lel+T/AAxYy/4+ZydYEdsEW54+oql6ck7fkYId6xJchWfUPyldOzKqcgXIb47
BN1fnGgxOK9eP26t5wtSvuQyM50YG/niPY3Y5+DWvx3T/z2uWf1/ixoghuO6X9xu
nPPRyqHG4KceNd/1X/TQVJxY70NKWbrkczi8QWfvuvci2U38v3+Vyby/MoMFKr80
CYgAokBnYb2IBEbL4p/l/D2U/uQp7ceLsg2L9XyiSXR6ZV098WDzdvNfu1Y0EGs7
owGX5ReFHcXPzAtFTsnbjwlnutX1/tRtMhDV94YsMyKWRgzCZ5hDqnLPj+pNvRB5
GXC1+wiC/X9M5ccHjsTdY8QEyOHlBCSkacmFylHdRe/7ruSoHJpK08jvzqThQM+6
RhUYHVCCmAq9xfHCbqMyT7W2CQfKY7DJOahONzH7JnY0ATVQwy5u/iNkjRLjO9k1
DhpZul1Jmkn3o/swduIB095WQoGzAfdQPrizVZ64vwAKPJM0DZxUnB5Wgj/3H/dB
LP/GuH60LOrPTxwxO7+0AMda8ZBwIEgKT87L++XOi9eNnGsmDGkUPBZj1dk0lw52
yuP2kNHMvGy14wOuFxm6UxcO//islIM7qH9cwHA/6FfnriBeDBGCVII11s3o9Khk
ZKaefgM4re19P1DL2oS8r+ppcpdTuW4quetsIXSyOmgvwCU+ZytUbFFfC4ddeugW
OJXJ/ZhK+c9ujhasFHVKFGZtrGr8uIlXBhwqDVbepA2h2MS9UavFfTDU82lsdxBO
PAXu6knf7GfmrtK5hupM7p46MwZr93yTnfH3GYckwa1965wtVHLCVNvuCzSOMhWr
VXzSb1yFPlRls0Yp+JwzQpZnc8u4yFUpLDc46rBrvcdXDIuRS8phGvVPntRyIvC1
F9QFyKxnFojhEqx3hCCvBOU0P08pUvnZhcfXEAWk0N6HB1KUsZkDcdWqWUpg4Vpe
D4+I3jovugfLyr/MVX7E2hQ4dcsMhOgXM7QqJRK+T/2MV4lCAdMQKTyQHwmaju08
hprhLW9M0uVOAqtcG+wBA/mgYhIroRboHI+YMGXlk0SsNdCA7N5v1u26rR6oNVv5
UkkwlkZcPwUTW2IuAhjLqfZbTLD1JcRYgXP3cZknOqsRHoHqDBEJ6k8QJRlVcomH
YwjigkE40aXHlzgegHJfUnE4KDjGnUpL/BxNclCtHzIiynVTJIG7LlFf7pMfr8Ge
4WOCNwhxqs1INrPX5FQFrvODARIlIf11/a2gPwhHVikIzrj1QfDzRzUIEtBwvj1q
JXDbu8SW+bGr3Vy0yuXCAxvK7M5Mb/g1/DJT/p1ljAZQgxSyGstljV2ZkWuQulpT
8PK6LJAoZHKm4ypSwSTv17SirbyWqWGOhySkMT4IPDpHOTxr/qIxcp5if0QTtFiE
5ajYVBLjdxY/mQkoe/83JGg57BJCkvl8wwn2Azrr3bMzWcl+Vmx+1Rhw98kFy5NA
IB9sS6/xrwVU0t5zAxsy9gCd9kH95FivjUig5CxC941s3YePETv9gP74kW/V2UXa
ARq0XfRU+tulWgpYvAYFknICuA37+mygYgnKYkdzlELYyVFWTsZjBwyR4LWm1QhV
jjM4WmmsoxYgOG3IR2U5dK/ndfQHkAw4TQIYkFRRwH4hKmfsxTzE4MifzgCNIXL5
GB6TrUyFiF6mCbvNTAxKfnKxwjkwfQWGDrk+DQ23EJsD62vXNMpRLfQ6t4hNGUFW
cg/xOr6ugstl5175yyjg4Y93RlBjU/9W7+JRY7m9tl9DgEtOX0IrrYYAfF/hSOci
/A+GHzan8y8a2k68hRpWB5MgML1kvtin1neaWAQdElO0Qo/8m5RosHnihsSWxSG5
j9CGUAZGdli+e6RNy7ZljmaHAbqTawnUC8DJ/82oYqAtjGdAqYIReO7wTy6XJ/Us
O+wMehxoStQ9ZI+P2YFpAnpPU0O+faxSpdJZ7GOt+EHZCkqzbmYmXBjn+SjtGMQT
G82v3g32X8ZTtWiBYpzYxh3fq5Bu+H2KcMoe5rhKMWF/izUkz4pRIsD+12iIg5Oe
7Y4iIpGsdwROXqkR9ZQGLaLS7bm27qrydHIZLqpB9LvYtI4SoAhEXew+ONM/3mQb
b9xVMj8fEuRotcrxd3dJoHaJDkOX4YCFGaUdHfbkbpTJWon86IHrfAI1PJJ2f4dE
EUA6k0Xn9DHkbQ9a9yYzTQfH4ieqljC34HuLaXXiPnQLmFVRGtPwNANV9JG+IJNK
h6k65YaOwdRPdhfLo50orLDW66IxxeXGs5ykZVYixtCD+YSVlM3sTnI7DjF6iX78
g+oKAYWFLpvm1LF524zTuQ1GH582MfqJdw3JFhN7Ra0FqRXpvYrqBBg3F2skS5Ez
fVJvTTYoN8ouZXD2YBZ/ZvMsHEqdrvaooWDMz+PU6+fnDJUMD399mAEkDxQljbZY
DaQT+CbD9ukAeeCWLqjDAvlwBcubv7XpELEMs1+IpDYB2AdzmVOG86nrWTDcgOnk
PN3mCXmcTm3wFWNLNLC0Vbxe2lXGoamBi2a5ICNuqxPgZvB2Srt5p7kpd0QQ7eUP
kDQdj4wkMEWGFBZVVb6XgqdatvczT3j4YuGFEUl3bdULPmKsUSplINfExDAGQkRY
C1iFH8sY8SidHMaTXkxboXkiyGrm7lmbPaF6wuuOBaGuaf7gmPFxcFXEdSHK0M2X
W8J/ClJOWg/4W4m4J/yJDnoGHeyLkdaCJz3vp/msOK67SZ1Pq7HF/Zj7mH0/LJOI
BXNy31SdI5a4Y1wchNCnGBxyOIW5GOkXLO77Kg+o+q3rpEdW9qayDMPRAoq5IlWk
YOPkAI3kNxg9xI53v9WYeXayx0oLOUeU4ksrRTdOwvFmBrVanX8t7F1+Jyx5Vctk
4Y36pyeXhi0n4RV3Wgk8WVTfE6KHrBg8yF8bC52fq6xFWUCegxhBf258OG0Pd/pw
kvBlTNII+FveCB9HxfbADmYtbideVcOryoSSonDoCZf5r86y3fwHhZnBxXWTbyx+
HDqpImFqU3btsMS5n+KWoiIq+CJ6ykkRpSE/1uYjm6yH3IQDCM1NTdgx19hQbIHh
mIAlaPWpuUUYhQKRySSJQqXrCIQhLHM3dQIFIuN5f7mbbo8x3Q17h6MZbt6qzXHj
J36dV9pRhtBmfoS+RuBLJ1oOkYrn2DdCcQYGYaevxrlH7ezg7Ya7dfE3lnDYGgff
r7s8ztQeGuUJl9RYC1UG0K6PFk+vnrSYkmSuW4gmvqCi9fhqBX3v67E6v3pG75bh
DxUv7NtWsLeNlWlPrxnfdlY42hHhjKDmwOSccASxtFHnOideL1KZ020gey7h/ljz
bS3RKAw/9//Rr/3HN70Bg7zCf2Z+qImsxImK64VWJwPOmCZsg8t1p49+XWmuGy+9
HmGA8bzEtyvgVgoyRwu9XKgHmtrYNaDv/kuZmUDfiSO19QglVrlgxPpbgJfAEVF0
OUCFGfylh4gQd9ZAM0nQ0uu+EqfF38PKeuz2vsCaH7IFUnRqT4jsLPQpU6CfuXd4
MM44D0JU4aACLU8XcllGQhUx6AxzjRycB2JMj03psummaKu2T9ws8fZXtf2B+pN5
TqkKXWZLQ0WbtHcbBSf/jgWgiBZpmbPv5zsO2Hj6sEZg87jcCpx/veuFwYwi1Od2
N4vrmdjxGhoogkGifNuineQ8WArx/WRdCnEUSfKFdw9Yybw2J5EWgSbY2K8/zGU+
K7/q9Mg+3JbfME2nIgCsH1zcgNeggMki8LKzSlstkNAMaauwgByLwO3QpyzCcnRn
gzVJnLn8jmSPa0nxGkq891Z8UId9ZUmW+1uxNx1KurPSXGnVqJ8QZEj72l13QOUn
s9e/KQy6JyMVgWthQLTxZMmlafq6h08YnQunQDrGjLaMZ8WiFVe0hxl4pJv44SZ8
IFgRD7nD3cZJS0U9TpCMFYZc9fbs8fM2kVz8M3uK3DMIm/RJrL+agCHixv4rrGdL
mGNrId1YyLHTyEUNQVlmrP/Fk3dYv6rGSGzr1dQYK7aWHcgMUX9i6dGNM9FYUqkw
cjiwuJfH9dE2ugjNs8OSBBckxN/YJ1EMgnmQfm6yxvWk9D+uE6aUTDlJfmWP2hGi
CN3+WK166Jpfkf8Hrh2RYMHNhX23Lx94v+bdHQh+cXWfO37HdqvqyCUID7glQC5S
QjQ3p3kgxx2MFPYcpKyJWnxvRCcASNzJvC9WETHYq/wpDD1b0GLrmPlxvUsj2bBt
nfhvwaoBSGpJXQgIO+6KqU0bJ8CDVu/JnzQEmy/gUz0/5HHsAHfO+MjPfuIIed+N
lEXy1+u+k4qFUL/XSX/SI/I8aTBib6ZLHIQOkiZgkzVSCR6xWqnJX8V4lKeIaDcz
TDQGnCJFYlZIwo+4Sz8mg+wGGgtWy//XgYbBeEBnSkIl6OQIHkJEsGbO8MgJnHBI
1OC/MU24AixUU3sS8XRlPmUsnTmALvawQTe+ehFet8CfGqVnDI//q8Lo9IStZWrU
iY1oGp/W+mSU21lLHebF0nbMl/kUMkA5TvBE79a/OiRvVyTcgYNGUDH7nLPX9hP+
XwKBb0aQbPRJvNrxGhRWGaKPSfmVWpkSq2XKe6JnO0NOmqtiIm4ak5s72osZtDJH
6dzCA1DviMuhmnuI/Ffh1KkGtx+hGcpgpUFI4boQBdsfm/vS6+pOMcPZWYaTXE3e
bqFqyDpBNtGD/V2Lm9w0C5fr5YVvtvR0wjEadwistv6Y0spl1u5Mm3mdqp9ZweKw
vTIu1Lww+NWWynC90GO5g5dbCQlyEcPRZd5ZhjCw2vLBxDA8GSq/H2F1bGa0OYFQ
+RILsTrWcaTn8KZ72m84meY2YTYAmQq6uIn45A3XWstQ3gnbM8IJBW9/3tMWj0of
Pxfd+RMbxJUPuzAFNk14S0I0DxwXCasq+2p0Ck3/xRtn+63ZNxI84kCDxHsgFDK5
4WbUkrWPCNkuOOuKlxtS/fxrECp3QdjbMO19Auo4ckgYvCjjDSaAgPqhnCjyPM1r
Ljwmd3gyNQO57Nb8AFJzPKTmFG1mK8PHx8SS/0yJba7WuEDi9GRFBtZRr55Sb4Zb
c7vRcbFL55eXnJp1WagOSz+pWZSW3nRMCGpxe0qbzUKBtRq7GBDsSrRtB+gmqJPU
tPsk6vuUc8KhEf0MokhSY0oPXcmEOcXnrAyN9+0VYYmxkvn7LcH6bG6B2xqmZsHk
5afqauMUTV65uZi8hz+jbgIOYwB7hntbk380t7/ixxceshD7DgDy2tKceGpBw3r7
YXhmqyC4MnxeEXd0KD+NiQDFNshf8/DzREIFAE2wY1Ft3WQxJZLwjt6qBbS7tJeb
qAvq2HKhuMxRLXVTR4csEXI8tm/lUewBzPyrRN0e6EtcR4ssS5H34TuBUmKmQrfa
NJEzRYaO7qpnei2g2R+nGuRpxAS6PW+vjJT9HYFPYHwIEj0jnZ5RmcM/7Gfz2T1y
/bNnMEKwTMpLqR/OjuAL8OBCxbl2RbEGp0DvWZkErmxefxLojDKrEmP3U9AQgYrV
LWdZmXW/iuP+/K08r9bWrJhY1cNR0S/ylaamziEvFR9+ud/EzGJ1Tdpk/hK2iHgV
NT2lwZsnpciG5OP+OVmEFNoGJpUJF8caXypUGhBAaN7ySNohH51hUtPD6H5SKjq4
gufFHXL15l0ynNzFALQOaZxbZsT1hGrytahZaHd00GjkrXTKr4tu5p/Nfz/xlvhD
UvSo0OKflWTN4x56vSTNmJy1F4b7QYJJhLcY56CGbKFMiNRPbi/mqbIV0rhppeFK
/MtVVre1y1V9/XCWt6rXimwTr+VC5lKAOitdw1+uM3xe7GJUs8g3fr+sqWOoaTFi
j+J7wT/XAc69cxtXFqwv5+5dIYe4f2uxHVE4esx20V0FWhmzMUSW+73pKbTMB2ig
kamzzAwZcTOMo1ESadgZf97dgp+Fa/+k1BEKVJr/ypS9O4cLdJM7d1kepTbACIeR
SDkgHNrddlVN768b9V5tX3ALldkcU1X7ifFEXIDatvOxfx4ohXw88fbzpPxFonoL
Iv0U+Fwfkgb42LarTBx63TXv126lbxf2xKOgGRKvcHVUfXZKyGLyRws3rhmlA6CX
ATb3RtD29XIGeyyl/jkLuf6kFb4YPSfjHfchsBYXqLBU0d/fdlUNAkVkliX2P8js
29af+eoc21Kkl+0CvvR4Da0SVvgBr9YzElFJy48tReggfuybL3zzK759S6WDGWDu
FgNjcRfiPYEteMat4hj971KhJnd8TmnC6k1JfFtC91eU2Nut6y1rrYij0l006466
uCCBCmUNLoaetdcrLUvCHbX+CQcD0xDppleoKOzAaA3LtFyHHME5i6t3PNHFBHnU
4QjmIViq+ZpzlnigdUK/X3pf9EaMR8MHLeEKDRo4qa5Kf3do4sHO2PMunDmMit5i
zcZsvbaIiAAiz7P8B9vREl3CSRUedxcHVVQwWIdh+iDE6m3AHohY6Ao1p4AO6J5g
144HtMvuwX8jrA7XqrtX7pNKPMJqxzI1/LlbF783y7om9DrtZvEKEpwvLS0k9S05
odcHIVZ3S/1UeNR+22Wl74w+2Ai66bGvfYTljnuzODN8DfriuFyNAjlCkQvMxp+m
LA7SUGflRkdW3Ul4AyMC4vlcs4EPlK4mCAfaGLacilAF93g8J8fsEp3h/DHTbUc2
dL6NpXB2tFHrulHe49xGF58t7ddNXsm8CLtn5W6gZTP5a8Kp1J/VeJ36bpLsLDAw
i/5XtJQFpFarc19tEHlyHVJiA7SUX/ANGBpaRFPNJxpRUsdtzcknbj2yR67S6Sdj
2A1jLj48Nm/5hymsXNcJd+ymVsMSSYrhziSz89kLVYevTYYIPvjMRE//ZjYj1VK5
exA5RSavfcVDVW3QTGDWcJ+8Jz8+Zvk27t+zHGVk1GgzqlRgktqzpTEnn4k1V6qE
wiPIVFugJcS9zWeWCi+2dMqoNCP9otc1ZN33wzOINgHMvgD+T24+yynmQmlBu5tF
2MlnMdlMykxBC24LuEZy/IdozMBtBWi9FF5vRqolWwEX1M+xBSG8KobC7B16+8v9
uqlJmuA/uT0ZH8np85GYjI9sqmfpqvruXZ6Qq/FkdhuBrZFmxJ0EL5QhZrppcbSc
ojp/o3EpRla9ovawIaeytxgFfIvBksBS4GfVFmJzE/EDplnowivaq3ne9J4FTAmh
frakVt6KFI+tUAWlZPVnkkvMTRsdv9HfFK3OhiSJ0ma+rJpdJnpAcc3KjHukjfek
CeSaTDKHmfL4SAzznsy4RFMM/tvX7yoV6c9yvbGX1Q0YRJVprNoxQKYJKMcg7Zw9
2kX8DAJbp5ObAiwX3gqgiYHPasbcwxwbheu5g+if/UAcBSau4uT9/+NFrvjOkpEv
dsSUoSRkPez/N6plDzCKu007UPs0msxPRItzpzeDdRdZRqlyvmA586Uebz1irbx8
U9rC3D3DfoLi+S6zpuxpKrzwFwMOy79mXf+srP+ocG7zaowd7rXGZ58DpaYSrzUp
YfOPvQ7UKjFmklwfloSd97Dog+l/i3g1Edx48D5/BjXHX7iErcegDqc4Ybl/vazz
aYNQZl1+D8KmqtWbTv94U6iOjYYdfRL44k8OPczB+/dhtr4TI1OgZRK+sUlAeNOH
h8b8Ts+sYC7ihfareyNBtO47VKQQoPhoqJVj4wiZFUYzC5I9on31jr0Jn1R4L6q4
oQJDNHD1WoHf9bPEH7BdMx9qdPs91Uu+aQOkROVWuglOWeyLt3xSmEE/G/Qp4Phi
aQi3WmlfHAOyD4pA4t83bSaj86qxVn3UqSW5nwUU4NxIPP9wv71Oon2Hc3VFtCHm
RLtr6BK2AKdjdAkvGITNWmYhXdP/m6L6DAzN6xa8j3xUMWQBAhhRLbpHorf8o5O6
CNsFTKiGpjqs75DDr074VEFxUybRafk/wj1TGTqgzb14miZDkBMSD1fi8kP8s9DD
mCIfU40j5pmnPXg39e/cRFohKkT4MyLsRQ6yOd4CV30l26Q7xuXMpT82CG2L/d7S
sUU3jDLTsdManbm+GTM1RmtKy3IUOOQyK9Tch+C7hSoc841ITvDiXQfH1ROqBVuQ
K6ZAtap1LvNhKPbuYdHAmBkKulYH+agaZBhrK+x6dswYkKhJQarKRkBMlxOArPOl
ZRac0CPaFm4FO0lcTzdulCsaK8JtTN5d16cDqpmWxMfT9tJj9x4Zzc9oNdEh1rly
eCjKvyrHWjzsuurhcpxfcGsTv4HKK01qHaNt3evnt/S52/jCxxoKyUJRKUHBQFN0
FIHfKhhDjG+maVop+2WeFy9SJqSdfjx6CgbkQhU89bj58FhxWsubFIu87ir+7zS/
d/G7XQADEYj7DUzDXH1RVy90gpzgABluY85BOWKohDapFHOMwQSJp7JkllvQPgLa
ZXOca2YH75OYRtzWJ8ZbBI5D/Ju8pFI7I7l99Oy8KQ3o+xWIWftw1gcYGlkyFV44
IvH6IJPuz01T+cPee57OnTvcshzlasBxSh0XX32JO0dCXj41GX2KK6/KI9k5Ju4C
1k0S9m30AE1ABr3ffAeXLaQWfRTLqbv1SlG1YgM87ySs9S2m0cKSxzfyCNSaD9BY
BvZ73Y7Q8gzozgbOQfxmPMpX8e5nY+1nHgIfZF5JFZDke4ZPKFqJ2QH4baPwSLmU
cl9asjSLEWZ0IzhTbJ1wUs2hJ06waB23rsrds96aUZkGkIbZC94hSb5iRYpxZEdQ
cDUDEQhAshNQi7Vo5rZYRPVI36FA7Ap0lk50FMwyDRCypVasZ8AjVnkBwuggEd4U
Y1JgXQSwBhDm1SPYScgNVc3JQBGLfXXGdLCwEzTQO1Uj8IT3eQ2rSLnDdW9/a8wN
OqsrykpPjOngXrDd2od1cj91A/pEeV/CD7mu5c1+H3r1fYjGSxq8HCD6jT99E1iO
uesvZij9KxpcjaViGYrrmuv7Z3XqsJkmEHZe4Qm5pVPgUcArQuYlIwSMUHroeZn5
iLUU5xZKGP9DRi0iq4coWOzf9NnbTgjUsURQNE6nQL2wI6JPuJpQDragdZFf9Pg9
78OQ9bm19QqEgQEPKBjn08827tlREMlm+ao1mwtuo2tkhv3MLeuZ4snZmUMVjDmC
y0embsu5aDguq8R9hxQFjuEjh/2PUh1rDVOdCHX53vEnPbyqK7K2s5m0fNwOq95n
suK0LrYNMR28eudu0u/msgJIA7PJReBBJC3rYZQGmzF8y7Q7iJ3kn24LrGl7wgNt
6QrCxUuwmTR74ADUXtEpYwH5GmiLjzC3kL1kRW+xDIt2nkYoKWwpYnLhKJVbxelk
hNba4o3uQFatJ5Z9gPmg7rnxq4doYGe12r58JmcmRGRwmryFTUOYPkPf3PhUVtx2
uFXhLWpGdOISdgMpDcvDkViBFZ7i8c6aDf878N4skYppi8W/uCJMwO1EWV9OPGl3
DMgMFuRiLhndpbnvtwlUjzpqjD14n8GFhjl0NTLIzcyGnSxNxq/MGuf4lRiz1mPx
VA4hCcmKhp6XExAIr6Bva3DKdYVmw70K21VJPiUFCvnDg5AdSTA/oycIHgcApLNS
alqToWF1mI5iHEa6ra6HCyhVyZ8KPt5igvid/LT03iftrc+pw9AxAiUslvgLkMzN
XmB+2My7TMx9BJVi5KxJeyrepgWRftchxMx+a5TsoIVpiFLanV7mabeTwKLjsywP
kesxsKpdZcULsD5wl8mK6otXmH7qw9NAvP5eWJDp2IDLjVVuv2Bf3rxZQ6nzC9Hv
UaA1HLn83T1l11N0iD8/qysWxE97hn9nXF8QPghRkOIhsehTCHSV9UEVepByFyyQ
N8GnknANpFNUuajarayN1fdFCkpJuaqTyIoCxI1l4irWF39UGzGj9ksCvIr3srIo
W4IxvR9PQ3AYc6MC9L0ESLjDN70AT0NMrxMW+SaLhw3aY79CiK5MvBw4GHwxwleH
8ooa8f27wNFI5rROZ5K6xXqCiiPLX1jv3cxCcLK8j0b2TIz0TiYVGQ05MGA2cI4o
dUFePg2ZRxGo6RGYIq6GUX4+N9x0Q0KoYjQeXN//GexbT1g1KZehPlDB+vpAXNuR
1yhKsFG5dfjt2WVVafK78z4ylJnDmuM/ttaSl0P3fQtZiApaDFyTk8ZCishTc+G9
ON3oSdOoeeYXici5pXq2qClQzJn1+YmaAJwyiUBvajkw5Q/8dwvMzCpbrrFtLd7m
C8kT0155bgdQzoXdT0yiAj6v5s0eFfOcRLV+h3T4pmSJXnRbSTFuWAu10y/9PTFF
nkSbW0khqwOpCop6kpWLzM+i/dPQ+MyV1agzF5eeJ1rGCop5mS1KVOtlnIiAYyMi
sB5c72yzZOGBKeLQEpUX8zRP2CstkFe6QruGyZKqnY8QDXyFiEFWG4lz01ms3Oys
KoCsXuLRexBbIizs/1Q7EdfB1TtZIJfGbX/Jdqrt2KH5/33LBUCuarLJ2C/2GLiI
51T+mds37+ApX4OSQP75KzmkqjivK+Sb3ojgYTyp0hZDW4G27KRKZkyX6dAjY3XR
aZgWE+Hmzv1/dX2o/ALvANO7tS9Uf5T4Me6Gsnws3LYcgN+KDxqxKgv08qcxAG6S
lQTYthL5q5CYsTawCtGla2Y4iYAewSbeV6W9qVhWc1GefzmQD0I+rZmezWbJTY67
uNB2FE8ijuAlqDQSmg3gbI1jovJJYc0KWo3FTB45k96r1z+4HgnOy9xV50/TxwSj
XoK5UeYY1IWPucCsNkVEJqNKpp9Xsse1EyVrwNa/5NnWAE9RWteqjjsMrsJS7nPV
Ib+RdyQwJabqLH+Sog9p0YEba4v1CN7gC+UNTqg+qFo1hPvXARs+OLVnILh0NzZ0
ZlPjq9h1mHnOqAiJPkP7hLxMMOLxsSFbv9bahxlnVT4KD+Vy7lmAiy8Q+3m6pp7m
kqgQKzWWaxgX+QKX4VE7WKXutEStpndncXSD3R2UD/CgkVYrXENzArUqKVM0Qqlw
2puZl53qI35ht4S50Piy9+gqKFl8P33g2iS3C14NlJ6lEx4xYel4EJ/JSkuxuQQi
x2kfDs8AwsVsAJMtZ+SeoZ7UQxZ+XFMz6YMcej8/aUjPnw553KC/W/4N60ghCV0D
9+1IwtXZ36Mrab3AdZ3bBqpgjIWog3xQYyTRGXb2RD4nWhsW9MYAfBDz4rRR4UuS
SifeFZCoTkC+FcNNW3DqOpUvSHII4O3Ji5TR+dbGsFMgZkexZjT234GSfZSQy3GY
b3GjZYJNYusQQoWW7Y7wqpKkhtKUSfzl2RW6rh1EjcGftgH/zjPVSezKzV+sgL1M
Lebe86J79jnY2xKeQW40isJ7sdqo7YtZaAT1BxgXX/PSYdgl9eFwgPNY539BSxEK
O1/iaZeQS+pkUEOCPdNyZTPmyR0TFU9SVOedv8RqdgRuKXx10OCjw3YNvJaLbypO
GNGFG5ogBLY3hSa7nmusi0iNwnQ6MsGZOkGZ32MW1QAPD9676nC6ORPQptzOGCYb
qNxX6eSEysBE4sKe+KI2SH0pG05m5nQko2Crbj3b8UoV5UzuT7K57knqfXsGa9OH
ThklbW07WeLoANxQcuNVL88JgYzmCir7q/1zySd+OPGVgast043ep1P+u2/NpwZO
WcMoabpxm/EeBehkbor80ZqI+zEMYSt5EHEPUysiaRxKYxjsCvY+CUGr27aEXzjt
rOr0jo3B8sPEaNqpIshOaU0WLWURiSoSoqC6+ioxXhybLE59N55k9trFMlSPQGf6
wJsKVKLrOByhAHNnwYHk4QLNxkMZ7GB+GkG/Q1oSI2wxPFdUMxMkZOiZlBL5hdbR
xoB7DZmQEOPGl5QF8XZkq+JxG+6t0ZzYYU9Po2VH5WYfTYa5/KKmEiIRG2JiVglq
FtoWZXYrZ72Vo7aClZfdnaFKpgp+AF8iRoul1xmBrtGj9hx24t9lFwRCn9qQ5WXu
OCI3jF6/fEPXiw3ZaUD10XVlbZL9L+uxh/EIOl+d/x1lBjNO3J4KLwCzUe4XVAnb
lWlmJTLWHouTspM9F7MoOsJ+qZU5MFb5QbASBiaTg5ebPqU2sxRNewc9CqXISePC
U8WPxQvqJ1brJM+r5kSW42zIqmCHfKV7YmHl14jOU3Ks7PkwkzIGsLilmD1Hju7y
7q+wGS732RGwzrj42NkOLHAUP09ZrUBmiBQVrqp0qiBCc0ZqixyChDgFu0rxqeMq
wOseQxocbOj1QVhhDoLzYyahCXWX6sx4m8vW0xmKEtPHGKUdawPjJymz7Zabnqvd
eAELHb//ZePaqOHyoTB1kdfEPASckOGjXLLdBGRgnVoHheh5MDCtttytqAV1Nj+Q
nveQkRTmhfvFs/amQI73bG+cXOZ+KBa/zI7xLpSIv2biQ6E0U5uBrRt4nGFyJCFj
/oFXXZF1PfbXGoj3wg5d1QEtjAVT0/khWr0bMT1J0X0Q+6VxjP0SLA6vx4z5iol4
fP6ZPXzRXYmRQl5qzqW94cLS74xl2fNBH/tP/0IrUffcj1aNPhmcjhMT0By21GqR
Y1sdYtya18aQwx/d9CBHtj+6W1G4L1pLOTLbhD+G6URvmtQ4q47bIteeUEwafemS
MaVnLzNWphyAu84bHke+CPKRSLrJqPUVnC8JXMrbGaPfWbx9Q5O7n1mOovBfp44t
hLregvQk6EYa7THhYJqvuygm242YdHbDBc2FC5nUj4hsYN+SkfcwXHOXgxhJhfgc
55zFfejkV2drQPnSG3DSgWvuFqEw2bL6Btldm3PZ7QGfNHohaJ2LJYdKzpW4fjkQ
fRzjtIs+0v4ijaMd85IXc7CIGz8z7341fVyoUuPN5hyiyct+0gljkT2rD6cWwChD
KDUMaQJZ+yA/eUxiemVlEE5Yg0kCyPjm5iI0XnpspM+H+Ctt77YTkw8GsVST2Fvf
dkC5q/U3gzfhf65kuVzVOE8NV0K+TXNeTCy15Kl4Nb/gm6tKIwUDVQkYPEIWxF8K
bAZ14zHwNKUcBRqqz4Ha8U8yKhHZtwyFKUlgKp1p8ZrmSwniumD7UW3c1gVd6ouQ
Z8yPUVhgUSsGn9Xggqiu/CbZVh2DWy3J/S8e9L/BVTqglzIjAtQ5TqEpDZ30ZaYV
uuOIol7Ed/5piTz8WyOgtEHYcyVBfpggkGV5XU9KWPcWvdPeX7T0Au4LCAYbfeb+
vrNFE2/UlBfHbJk4YhEBv1zcEB+4iAvOA3LTEedWPjjRb7o7Lb6yQYFIbQ0viITf
fSYAwRJet/KGL41kVnsj2O13Bf72E1/Q3ALkrtGxysyI6Lthl/BcAzRlCyu1LGc2
NdLIv+MekfB36dELfQXBseZuRPn0XWZ2Cc/TUnW3Gjx7OUH4hgquZtWC5dVNpLKv
nZ0FxApMnMly9Ta4aI4zVXBfgPbSHGXvhV+BD3fqIHhpPDv7IfuMjGhI/7idkq3h
2D/WSJeUwKvjwVCuUD8dkec7YSOGJKCSgSO0Ydj/NbL0FyiEBL4r32U7mRHFp1i/
8UZlOqYKyVf6tra+Ahm5YZvmiaiK4cTuTbpw8hJzZcNcv1TlEdqp8bE0ucVzUvhi
iX1HJbQZvq0vgiKB+/bTU7Cpod0LPNHgFvpL5ZBirCb0guCtuvaZDfPVmx8DtP5H
Q8DGTwkAsJmHE1jBAExlBZVlFZTuOXa1Mhktc0VXI6kez6Wvg0xP5kljKO+glZDX
0rVTAk63CuSe8Jr5+FScnj04NDU6saEOq0+ArdxT7jEvhHWCa5FVlzAATnZ795Wg
6OhB7B5EUKvkZvfs/U/rr3w0D2EzVcWMpxjgRQo7MgyGOBeAKkzrHpjqbc0i2AWg
w64rgiGbogD3VybpGWVJUt8ydrSyyoMnimyp7MZyvE1gf16r/8hKDAZNOWpcc8n1
ZFr41bex8bDLv7Ay/2F04fWFZKFFaf5hfk5AzSV1E4pflHUO9U5gz+m+BaFQMUd1
whhhi51A+D71Dzxr3DZayfiXSp6JnJwdq/h+EVdIpL9u1TMwj6MjG4AKYQRsvGwN
H1AjV1dw7MFM96C0FRa5tgz/GIuOKRdjsFgWZ9mcFgbktFiZ9Tr1pqLcU242FSzQ
78VKSOfuRHmR5VYPjk3LFz4hdNtFT0VWq/z4tU8yzki8pTooPaPeBxWRqj4iMfjB
Ji8H8hr8RlUhPstl6/RjKB8IA76jHP+uiBvGOjzQAOw2wRIvB1DvBayV039nFAso
W2YDPFDZBgslWdqQWkq02aV/PKhor/IWazJ3SopAupHwytrWHnTTQNSWeLWNYNEr
nlSsBbwuotv2dWOLZ7kJsmtoQI/Z0T1GxzTQ/9k19O+r2GtqQ+anAvipqKp0ElkL
vN3zUeHZ+KdNMA+MOI+XjhaOYR5tnsD/k7nBuau4KHasboyQ6JTF6zDyffOw8sYX
l5qP0uhQbxWeWVfrE3GoQacF3NCmBSuSL/hgJiDi0fdimySADxUDGx8bBnRJLVLN
ZHC2aKpvrMVVncDyZkGlff0CiE6Giamz1g8IWFRT00cMmcUFM8oiU2tc6RCdBdV8
COH04o3EB2L/eKMCNwAiFxheW/xcRVAXiQQi0NKuj7XMPtFzMc4NC3DuH6F4u70s
OU4DW+s0heqW1jTO75hzuD+kj9QAo5VhzrgPSFL3qRFfPB6fwSvCxGJQ/VGYEnzG
lhfBahBfcgtrcCZbAxtCJ7XIWdI2NFfqiuAokFre71hMUo1CtXwC7GRnp1B6MYex
7BdrpqiVLluhutYe6LQEeLZ2ezmm0P7vxcJQYlr54z2vz7YJtsuiyWDbfMG6neLJ
zOze8rjikYELBUQ/F0fJFviOe2CaN3WX9PSgNo+mWffm0VYgCN3LOCpW1ElMWw7+
lqIw48EJSmJ6GJud926Cimq4vylvnzcixZ1+FTloViJwYY3rU7LTJA9ZJokINYPd
ytOl+sA6YII9lVs1Ic+u0hzIQ4PJXWPq8msYpKcRvYWRfiMp5blsynycK7aC2UtX
VbeqWmoze5sIoFqrU16EJMWqqAn9UeDT7OOwoupK+bh8QBx2yzVGMnzlX6QQiyZY
BYy4Bh4uXuKEsFQAVQRcTq7i2AJ6id0ZbrKzGtInH/fEzZcj6ajhHudNjyjeuPDB
IMojjE5o1R03zS3sQc0X5mNvPmkTOtf0EeonAO467XOsXDAOR0KijMmLMAfhlJWq
RlWsAh/+EewbkOAMSo5IvJcyf2ULvG9F9I4C4wELpUZaTg0aGHbQxQtmKcTlwe4n
UM3umYSgLLplzXnZ0QYnt+gSoLyWESAh8OprKm6XG8bhqdOSr0nib6hPaxQjPTEn
p1SOoAE5U1qfjNhjmAgoowWSHIhYfWDFdzs/4m7MeQlR5I+YjKKIRUUe3uL3J08K
eAbVzsrVRvzH4p3p8scju/4O2lPUWy57J1QXvco426XoOnpLJtsFgna62Yt8PyvH
ufuKYY6lnulFRdNSzEo75vXZhaCRFoJuAEhyFQb80cQbIYjRsMuOpsuC2EoHY6MD
Y0i55K15FQ6KOdYoGuIXt14VOwnlHtXme+v+hXihlXsrp9kNgg2Xn2nl/X5z1VA0
ocC/pmzjwC1DLVmCGBbEB2ofETk3Jz1grt9xHqDW8RX9IOPoemTqbl/PYT8leifw
6T3usMzmmxL7PJCh1xapRdigBqkCvNU1cet5+fFk55nuF2EpLLBciMdPA0v8hjZe
IkcsXzOtPNKBtxy3w+f/o25C73QHLLnqaocx/qD0HnCzY2J1kzgHp03F8NPP3H8y
hBrxnIpJcV3jHUNCbDZkquWD76VSzkr7WujZz/AkjyF4htCyXPb1RC6Nt7gUAJ5w
knC/jbdp8Af5Lk16PygmwBO9sIHqvaReUl1eenZtOUp4k2B0kpfHF2PGOp2PcDf1
1jZxbQIVoF6WSE6iwNiSKfuMxW5BmkWQG5yVvByoxoAak9BuJwP9evxP2B0ywcAZ
VB2VLE1GDS6NBthSOosUGEmI0uZXBIcqOPtWN81/qMQQaOKCR76p62MF40y2LVYz
aevEUd+2+Xzd0m3JhmoV3WPKu1OQIfuaparuLw9kqJD4wdOHQU99P6uMxunhHK4C
n2EdI3QLxUdbCUPeh+lNDeuTk0AP1roY1X0/es1DCbg+nUREL5DyeqGb48T8QdGb
h2GZ6gKKx0a7teYcAv4xxzwCF8ov3NY+Wvq15UA96i12MdBXS2jaOI4NPNHh3KEe
Vcz7rb7GyXG0RRWSscLNdWzBPDRWn8r+SkeydoURxNDNfqTQKEpe7s6jV1yzllei
huyzztg4pOk0i3BIQqRHZfd5u5m6zel6qFPxNWhvp4Z4fmXSjaSzP4+Hf+aU77HK
haeXu/vtj7HiREAf/zv+mE1Ee1vJD2hHvvUThq+tf4LdCX4BsbLtT8sDmexoLK6d
nAJTbuzdX8cHoEHc9XIs3YzLfjcxQajQVfF2H5AJba3iKe7hS4Qfk+lBzYRJXP54
ylTeY4Wz3dh64fgsRcckoXEMpIbl7Us9G9J5Ybwy2CeO58HM8xC4NMZhQw9CvrKv
Za3pMQnqDEquu4EQFiibf2sfYi0CHipfp//scR6TGWEKAj1tqfdHMFBqe0c/6aiT
CRczZFRqiPSjdNSS9vC3Jp27yooV0uOIMmY25oqGcU+Bbo0G9PWQil2CntX+jL2E
VBBYB6lU3JzWusV3LpF0vc5NzU37m05p86VykWXI3DeVCylrfqWSzsSgmdvcdfQb
CKv9LNuzHENV3Swe3wlqE/zGgDkPVcOkeMMZJSokhR0BSdJpwgDnTpWpOYaTOE69
vvnRIK6fOp0lkwy1YCaO4/iUAnCTebrEIWVL1vtG7fbEUCtfZkl+iBN8mojkZflY
PP1OTiLErvw/TN06Qb71Y0urm8XhHLK7DeDOGDelbEaO5ezgrMV+ujddsoNMYhMg
U+qR2ca1sohHRs/ntVa0PEtTd1Zm7zK17P0VolxxiibVvdRniacTyZ0r2OXIMTXW
6dASFUzepyz7RcL92BIblxsj+c3AU5BegCseZdRL6IG6y46L0caUwd6/nWDbwAhr
xqMRn7js3C7u3MkZEDDBotsd7KE6RELa0Im5cl/dvb4e69o2pfCCS+ScHycaP8IO
jDlnYlKp1B616hbDhzJu86alO9s3zIBxR8mhBd7fk/WmlbzpaaBnpjYDAHowKXLV
XyKaaiwO0S8+/W13mF+F+XkNO5sR2fDMoXdrVtRD1n6g9aTAxRheN52cAo4xd7B9
yBJ4yPA6c6Q7VFKAr/9jLLM9ZaGrJN6G+soxmK4QQQtPQzNr8qKk7J/gGzy9GtXu
HRNJ+O7xKQZu63TPFSYqm39/gn2lo885L/3MFU5gxeFPg9+xu/Ep8i55xrKnSehe
zVQXHKaEQ7d0UH18N86eb9YiT2zkcDWMUViaeawWXt5Jmcx0yv7Ynm8KZAkQxxH+
ZgrGmEUGG5GMjVKXAE6zr5Ui7vIWH2DMz0f96wX86zC4MwNOKd54Npek4w+RSIp9
rZdNZmZdnun+ZVi91dExKvfCXRrmlL2baduryR/ATPEFxA7ughSTlXbwKy0RrkxI
ICsSl1iUN1W4JJ6S1C/oX8EyINiPybo7qTQP1n6qD1uVoOmZcKLhNrKxja7PR9Uv
AsH/eg7xPSuTJt0X2cXV9197ar+iVfKmu5bttqwsxnsoKl6ASuMi1Me+vPcKuqkC
zGo5O9ArKIRL4GZUj1cAC2uhEkZso2s0+lG8l3CrC0GtvD62AP+VC87VBhPRapdj
qXNPKCnmOojFjUzqt55uxI2vMXxb5XFaQ1CFnJNW1SIQIaH/6LdOkYCNy/zQe67p
SlJWGmO2XvIjobAS9i7QzvgD5pJN8x31i2gV8kmUD40Xt1JLVMQjLOpas2B18v/Z
mpxbjUlvj2C4txJiwXYMogh3GQaSzvJIsHDWXzoHmOHoDLbEt8SNIaLahUwSJxUe
+wHLzzausIqCjg2K0Q5ZoJFqF8QaQ+lx7749gXZpxc+5suZ50xKmmnJpO1j33A4l
ZaHO1ra4w7mCZxXBVYYgmRdUVPjPfnbxS4vrDjNwW6AbYrv/+0oGWYmXDV2p5+NS
kdIMkMIl5Bi8e6Uvk9+6zcxbjedRga3VCwcE162lsGR3NDTyO1D3PCpsFZiCD+kK
5lMwhm/uP/pzWVv1vnADeXFS4CR1Mq0p0Drs/iByvTzkdm0k9VIYKqUhA2Kn20Az
6mh9Y1OEEMpUqHW+6ObMoazfj+tMZgM3MN78B1/gDvZQN9N/dKfNr59fo58Ge+L0
GlL41uqOo+f3bDBFK0jmvSnGCR859HZcBSmSYdieMpw5VmPVc8YlD92UNlfbwhY8
Y7bwfgdU5GTZ9r7SqCtEmpZvr1W9Z18Ppghd1Um2pDfkHQOYJp7gKJNh8TGO7jNt
FXv/qS9h2F3fMJoc/iDpkOr2YXoqJ5BhVKjsQD+ZbRwW0RAwoaG/mHse6eJP3gnd
wO1bgWnomO7vYEpMyuEVoBe6YRWCnQpOFW71R4ETECeX6Pb4vcVgsNuMm3LRIVhv
0AEaGO9HxTt6e1uNIc91JP6Gb1ZyPXVNwVfJk3qq/xC+IgdeszwiKyy8sastI5C5
o0idVvSeVqAAMbROCzE+FT0xf4O9A1cja3Kq5/QTm3amxxntk0iFV809aL90TngE
fL25oWe05lrd0ZN6c/u9Nrnd7OgtakseRxYDsSLv7opE0Jyyk6BwvxtZQ4aoNPNA
Q9hjvJcFvv8B6oUqPEk/I4DzFl1+9DJhhYnjiwhVWBMh7d69EwBWB01yh6cN0wKp
goZjLiv9BWQcJGw9V41jPz7FxSsLltJ6ozHuM0JyFPUSF2n5K3bA8u55QAVodwk0
2tXeN4XtBmgxf71IyBCxgyQLB0j+41Psp8hLD+4QYc4tb+Fk+ObvMZCPhNXe2qN7
RN9vgPiMrbzllBqbTVNo5C7lDeRKCZCFC4E2C+bPIBOLjxbdZkZTIre8xxz8cseg
juvif0VINdijerCSGPYyRfFLzSyPAxQHcJ6ucpu9xGd8cQ0ut0lGh2Y6kqXCeEpI
hpEdH39c0qlHw5iFajam9Tc1It7BzJ29XejH21aPswPAZdNp/BE4WIKlLk36iSv1
3i//bMjuZbrfxOde13xl0QpPAqSVrqaeusgVcNRpwxhjq9CwyZvBi80oEMawV7Bh
RMWv244xAAMKPlBu7ZJQtMx7R26zSS6rnmzw3JxkV6LOPJaN8rQcYunUM9LK/D6c
uhDYyunllGxhZcaDoCh4FcMsnkWQ44KZGvVlaH13wqFv5Ze3HrHsOMpBTj1p0GNP
uXyxCVwQbVA8IxrVD3VeSzn4W1hcZpC3Vi5PKjvIa7ogvsJ2cIdlYtoi9RUFMBBF
AtHpLyAZnMsYO6gAC9/UAg5ZkLLz//LrsE10rmPr82uVrBOKR3TIe09rY9OsdA13
y6xO/Poif/8rld5mZaEu0OsFYUVR58SuWlfHCdhl920VeW1/N+F+8eg3UDDQ/Pyu
9DMeZAjk2HsyF+3os5iA7FcXkxSQcIbrFE6uAblxGQ7FT6+u6qT3SDArljfmHfH/
8TIAIbRlG6UVruGBdl4NAtf7VwPDL7gKYXdOnIo0xULPAUzC3uyGNJZNIZo7DR96
VRKCi7gqavlMRhF5Mr8/rDJNB9QDLfAgJt99nU78QJM6ZCAnWZb9FqaFOnu7ntIz
tr5SuoK+q8kpnO7b3dlkMh1SCOf9zuQevKCFLXVelIHLlzA3lhjobLKJDYUGdJtI
TEoyh+HdpQpVNb6/Sht+kX1rFodW0ivnHSPPo/Oj/q68KpE6eVVrR9Dftiu+aXuo
jkGdXreuwH7vKOddxC9Lnyk1hy9nxD88tYj8AoFjcClYWa2oC7kr1ZGkqfbGun8W
x2CBcww76Zk263o10umtYzkfFL+utgC1NyhXkLij+0HSnmJ9lqwK+khemf2ycSPy
K+jsFedYSdAit/v4hqQifAunPwDjM8Fmf64pBjV3TSDUkx3EuQG/OUnRW6bY1Yss
68xFccDL6EpxCkkl1lwJ6N2RFxZ9mheN0Fu2xZesPZIGzgXC+3dhQIED/+39ePY3
JCHoTO8yEXG1AI/SwQA28r97T+l0ivgOawuvsooOHpo1roxWtl5hW/fqiM/Zg6sA
T5ZnFO97eAZxyQUh1IqPc0Tul2yWL7BXVsLMF9fNbqv098YxhDFhDUTQyeoiqocI
1aIb5iEFOaaUEkc7eL4+RJufQRLK40VP68zScUpycJpOzA+JCVb4J2TlNOpU4xOu
7KybPy5DPNBC9a1jp9RJMi2ubUm2YDVmcCmXKyvbcihZvRyobji0kO0E5rktsAOq
2bQgn8ULEgClMMj791A911ut+xaf8ZR9EoK5jBpjYjkqvDVkgBjAzUx0yWwJ4xiF
jmok8ZzKvCdoiMMgj1NfW8AJM/zOlXgO9Etfr6RgNxdpZu7MrLgXuVzBd+rNwgxO
CspuVBPLK+xVolKsgYp6p2Ewsuu+SRNQnQc24+sEiFZQLm5nrYFlMjaPDNkDo0LI
AFQCP2MPW4gDiRY3HzWD84n28XKTP1t6oQg1LyB97gl6Qf3I6oGECJ1ekcW2o18c
OPzS0qBFF9aTND1XexJIjSrnGEoyo28wyQKMZtq0FG8UrL0yq1cDZ7VRcF9BOZUp
YIbk3YgHIhy8LkqDfek/bjj+blbuUacBrwUNyd2Rqfh3Xj//+tqyBnVp9n4e/TLM
1X98+zHqnpbGfv03wRc5mJDVyEET03vOyT/Br1TdO/trd7aAVuFehd+v2BPXYXt+
p6hycY/RgVHeeI5UXTXbdDtzJH9mDgQA1bRIJ2uVvfJxtnIz/rE3360dZNktU2JR
Q3+Z3jr5Tp8eazsqcyGjTUzIvoCpftlT5fdrJoC3lzFq0rW0fZ0ZoxI/Mre4Iq/3
sH4FUBasIln4ZHcu3zyXxhUBTd000pPt0WUDaUJytiMZA/HjcnEauFF5axrFSf8L
ej4e8gdT72C+z/MnLaEEuehVn5XbENHEh4qmjhVfWuz3TaCAHTrm07Zb8Vo8Ui2C
UV/5mc5E/k2Kpa83m5lha7OGqOU7JtJcIwolwIhc0SvaOSYftWDf2OHLZ7qnbd77
jG2xZoPJytMJe0LYm0WfyKD5Ol2BAambHOXeFxJa/zg4goz+tlhmvGsQoyGdHjuO
8ixgjQoP3w49sY6cFfT3O+W9aT0GPjBAuHZm2tGvARNfxnGplF/RSTq0nkVvchpV
oT4bLyxfAbqNYIlpFB0gXKGHcAiFoHVCJTA7djNH1TDRwPbmuix1PHWuf6nYyan5
jmvokXQT2Kdd7o2mNyle6mee57HpGubRMXUmD7aXilUlzPsaZ2/clAJP8RBCYF9K
5JsJcaUYsJ/JiCkUHE5dDAsCfSGzFjJv2rRgx9XfgFaLZ5L3PMH4zS80wUXZ3Ppv
bw5HcH8U9E+vrvOAnu7bay8DKGr8ItRjWCJo+cgUsq5gKo6i8tUIlFdTB6c2tWba
SQ3Ilx+yFsHnmsQC7Fdp5+Luesxlvna1kF+0ibefNB/FCNQnxcKJEn36kfb5UAQi
Q8ok1ZBomf/homS7HptD8aiRZadgdhz/qJ6cJ3xWzsIoAWBk87R2dmF7Q5rlPfKE
xvTolIMGC8CN1UUeNMw5MwmYx2YwyrqX4iSuLfiYbKoWh4JhzE0CxID1KT1mSvFa
3YSh13sF0wwj0vY1hyHNh/jdhkzwcZpCQQFO3y3oT3u3Ps9iNt6nY9mLDkGNqVy6
b7oAFW8ois16s4BZnL+d/1+W3sXxLk+qbdFNDNnYBlQr7jyJNFNhP8YLpJPE8Kj4
sZ0XK2u17gf9vHOa3BxQ565NhV8B1wDicKbmjVXtGm/lrt+JJd1JnS1GjUaLULQf
ukTbhOa9DoH/jJcKuxbT5+1asyiQCpkno+5HxhEqMF2GNlQ2DejAad1jrhyDoGtA
4q4o5q3FoVOLGpa3E96IgXwjvW0G8fYZ6u8QkuCM1UHf2pBWprF1sXyGhRad2nmw
93VRNF3cyLNB+BjYYO8UciGTKmOV2SaiizZ9x2D6e94OAhf3v2xD4STJ5As15ifN
FhBTiYHb3evKuD7+bLWLPVQp/mqc0agIdb48LX+Gj74zRNGOA9N0MBJN8RmF41op
B39w8keLSmIzL16EPcCiNlTyRD2uaWxxWOwY7zATaasCtE5m+HWQ3icDq8MxW3Bo
FRteIUeNYsHrbdzv8ijXB3bVs4CPchKmh7YrwEYplgqngPRpeCpEhJsqyjdbit5C
suqgtwHjlHF2jHj8ypW5M51XEqFytyv2fuaCXMsVXb7vJaptY3PgIf6zfnBB7fLT
7H2gcbE35WETTiFKLZS3AG8HKVxe2LPOPSaoIYxMkJe6QAptJnd1H7F7hRakVxtV
q51zWtDGmJXZs+JDxzd8cJCyo6EGJzo3xPNVUfIrtHLPwuM76oUpz9lIWfG7Dj7+
2V+wzYPeHdujVHPjOj0jSqG76J8D7W2H5hAg9w6dMAv9roKXPId41HL+AnyJ3hfE
s0VxVJe58c5hpX1bvoVTAmHRy/49iO5IYFjZZcYEgr0MXZPTZEP+vuFO2rnbom9m
Og9LmykN/l7Nvbg62mCHtLqNxhPnLpBy9PVRxrHeF/al3H2RB8nfORcQsMfMzDV4
ku1AhEVoHr68psgVK0XIi5C/yMMn6KAHN9/9lsg98Uq5jhWryw9eG40S7wLzLDVf
fuZFt9oVN04M1jRBoX8lbwZb5LXc2Px6wqutTOZqxUJK8Shq1WDbv+hlXrwtkMvf
6buda8YeCRgFiAavvhugNIcbjlgkqk/8JMbpwAGY8OAVs8SN1AYhvHUisPpGQmvq
YNWC18T2vYqhS/Q0T/0SFg5jBZ2xqo9Rt35h23H3LATSTVMD77d5ufce7BsXhUA9
4QNCwl/L3rPT+1YKJbPqxBvi9gDWQIwh4ohvV40rgIkKolXQjzQB/qPqmTbwvgXu
VcXsUMo627KMaxzk5cxKEwvzti+gAYdw7PgqXupNb/E1vb1sLgK/U9RxVlujlCmF
PP26JBQTBHTrXalRTsbSMPJVUyHGSYdoLnRC1vnBPl/ipM8Vtqwj/DQwKoFXqOx+
vRmbm+OKecnzUMRVeXmn33KNcyXGhbIMzqY58Lsd/LE/VJ4hGCnfCdAW3gqE6ksK
5heq341sFpcWZIeMReUeUjGBPEBjhyGJ0mIU/xZJUiDeG9DsKpkUMMpmOiZOMAh0
AlBaDKLvFNo9E4JEpvt4tpHs2gMEY9eYSTj1jF5zhNphp5h1J/39oh+ZE8dpWtIX
vC43lk+cQYisfpfAMJldOpmofEjofnB7tAuLVscqZ6IBGkNCiiW4Bpf9B2bPsWFH
nIdNuP4Yh/kW+wanaw8g4XA/Xd6DJKjM2h6uXGMc22RAK0wY6Za19nR3ctzJ7FTd
WVEybygDwy/jVdw2weGTk0xXUXoeapMavY+KPRATmw8MZxGgotIFwyzEtlb60/eA
zYMnBJ9Mjk1Qje1AyGQBgVfdJP04epH2SADKEvZjMm1CZYSsFmLgF41LpCU0wM5G
rhHSIYFi80WPJojxt3seZtzYEG3Ng8r1viRBVgKKGTSDHQ8b3S4RCIak6/DDDWni
MyNzXFAjTRHjkZjulax+hblhMQZ6RSyk33Iaki1oMPg7WAYXU2xjGTUYPMwFtNDb
p25dBR80DciS7mJhQkDMmHcA6ki1Vo9bDxQnkm3nnXiiYn7CJehORPP6oLf+vLoM
dMnTcLHKODP0bxLFwDfk/7MnSxPY1Q8jg+WZiGgxtRsL1VuTz4NJUu8TehD9of/a
WW3llTH+jcCLw8jzculXwLa4HNjmFxoyA8lnDFpSsxhdBoQRYPhCSjks2q6cubEq
Ym07nKiIQ8M7eWxh3QVf2Sc2Z2a0VdNh0iDt7l4fmV+lH5qQxWA1DeqtawmLoYEV
uEozMmMFOiG0x6XZP7PeB1CIW1dWj12Sr+lPTd5vPzDThe45XBY5ziUAjs1Ox+iT
byImI4yDYQpyRq2mr89PoDOMXeQzy7PQy3XTP/+b5y+8g1PYF8rdL/YrXm8572yf
oc0iPtQGc73uERQd6U4WqzxhNxa7XWaG/d+PGrO6B6CN8XbtUGMK5H+uXJZVnMFK
pvGuTroZRvZ35/yizORiIvX+3JGYCtjYTZCmD7TwUXxm/yij5gsAmpTZUHa6X9BO
pe5TAVSMsz8HBSMepwgs9tbyEmXcssYhbWWEAiynMYLt8gkSu15Lca2N1/lMLtC/
83gUA9epQSMQ/ThQuo38LP27DKBZKn4rsMf2g1FSN/5CALZ/iTjalnQMm+nsPlLr
a7YynRPAd0dli7+hNjNHI6hilyzLMc1Y0/sftTOotPSbFN7L1w63KIQTBC0WYGXz
D1h8IIBUCqYN7ITPogKkfZpTa0Wkv8WT8XTqZ0QBo/3xqESsPI0Xal4Z1Yf+ozeD
1i+NXqzYA5sJ4N0pde1fNC9DK4C1yH25E85mMRQfPI6T//Fckz9WjnY3V9K1lSZo
5+hgvvhgC7E4M4AHhH9k5pcvJKAITjcB5qnd0pL8XIhCmWyfqL4H146PzG2byTMy
iBrkk+dvfGtUD0FxU8ecZriplBRYcC4tkeM8/5KZNGv4iEfyRnCm74WRTdWl7u3I
19B/kYVLZmaoTSI8YDGlXwzy4e+y4E+Q5qflprUktCTcGWj2fkcA7c9ZNb+S3xj/
5hwE0BFfJE3wQ8IwAKM2WiPrf9TYW63OcSYum0zCrFzmux+DMl95W1Sjo2UHjD6E
kFBH8sOvCufJhLGZjgE6+Up4wm76wHhs3J3gXbyyyIMp/H0ozlBEhDM+2JaUAoy2
Pr6X+UOdHGFGF0ZO2JMI9a5MlhMbj7B67WXVa4VFb7u+iu1PC5GIgLPxsj7kM6bC
v3lnT8NCsTCW3lMJsp1xFnqFDNUk4knD4FGWOjEKKFEakF7/48jCycvR13ncs2Fn
BZx4LQOVC1i5dUof1crZ1QKiCZyAaXKsXG+g1+uRSgkcn345fdt0Hm5qqoEijmwc
Inh9TwehWbXurhRs0cur6aWsyPoGBPA0kU9y9hBJTLtonO5GBDArAvHFmg/z5ZMw
LKEWgQqFEpAo0TUWNKc6PaCktFIhuX5sEJ82ayFi4z3Y7DP3nijgvR/9QCExNh+1
4sDJyYyhO7pJKdiC2H+wOK59kgJS7Nz+ypm4zlAcQUl6QnaujaEeVSI/1BaTNFo+
30knaF9C5Oldr9enDbJ/zdEPfofvKoLukTwMZ8xsUuIZ0HbbIJEXXiKIcVqtRfd3
Ogt+TSL3/g7Cyy76EUGvtjGTbb6rx0RU0wmIXWkAz9UA/IBscTuYXBBZwPfd2ybz
8or3WJY4QpU9DXTc1n0B61gAmLPdBoBTbH7/v2P3ZfljpOoaiVn2kDAZ7Psrs6gV
o5qZjJM/cDztdekPUgc4HAebSY0m+74mrN4IeZGoeCnQZmgfccqUOOfouxGiJ9xm
fC+jTX/12u2TPCZaZ/bVYsFaewaqf6qjrAtUiIHTN+0qzA1+tQDv/L4+Et4v8k7K
i5NBfS543VpTQA5vIS+QKMCQeGn3rKD3LxXyidO9bF7FL4eyNrPG2/BJbGy7Z2lj
WEDFgr3j3KGgNGkPcWFDpVflZefX0PwLCWnlY4rovgbB/sZhenmCfYaz1eQius6C
zBsEmUMjkayRTtVpl+5zwbVYQpcFSmtSk1pYsEG9l7Q8rUHn4vIp9Xa8Tlgi4jkw
9IsobeuUgKv9a8OEUGk1ShQPwGRT5m8kjuHfD125SXw/Er9HJvRDm5LRPmrtr0zV
N4k8vugM1KEiASDNIEKzwPv1VQy5QFPXdzFogM+xjaRiO1H7i9OeCby26lZCXGhm
oK4SUbvRHfkNKdL/9ntv8XDZhTEJo1n0MmzqZu7OQnZkGVz0NlsQ/Fiv5gyMW4Z6
A/G0px8oaVYcaF/V/8aaTbhNOqE0XyN4YIq1Jm624kES3bJcIL5BweeUp2vhCVYo
JVYAZm37KpY4jvj9gA0ePskuyOgfTl+tZF8JZPlx6bVA7LSW6lcF1Y2dtb57vBGF
brZBtEYjR3Lc3E/fDAGd7xdct1/OexQp7ziYcV6efo66ISyx5pjdzGfkg4gXXvU1
xkYKUD/S0Uh+pNG9bh5pbgcgYTO6MZR5db64FEupd0wsV+JEfUIVKlPMoZNoa1D6
n8UqosAUU1LXKnDlusR5PchVn9vDKNDaDjSJLrR9pMEkhgFIpVhGMirT72j02dr9
eqQSW3O08SFVyALkYGe9b+DXpXHP0dl1eyPTbySG8ITZffG3t69r2BjwZfwXu1la
Oi+VnhuCq2amZcibMN+VW0DMJf/FYb85VMgR5WJIrqfxm0ZCOLuVejIYLx83u0hD
fg/k9olbZWzCXfLa21dsN2HXpuTet5swXoCYD8tzDlzD3aJM1IKfwssCsw5zkNrP
e7dAnSaEBmL0Rpq+1lvchwa0pBv5nVOobfGxjT7AO5jCIfLy4+HzGfn8uJ5uXy9n
JHNYrXbRMA4T4E5vjgsJGinNgy+ETX/Q+Y2TsqLyAF56qH2arBIdxi34kLaMAOB1
g1FAaGh5V7cVTt2IzGcdWoKZ2ewAYrc7wh6snfn6waKBIUJavY4ShSBL9tss0I2/
nNsV3DXwlELCG10RzNpTh2yVmfwpOaUSkcE68MvqfVehHQMb7R5M4H00ObBbviVi
9X+5lmHOc4qhTTKYZS/T6C6q+iwqPX91dNCP0b+2EczhC8Tt8Gvz8w1nEfBOCw8H
L4FM9mFLF+oxd8+AsIYaHFbw3x2hIxa15MLoQtPmicGv3usV9e5fO/pS6O6mf5eX
2Ox1cWeVDeCIylzTQboZFGdIOi3QseSJqliFoXgA/qtHRbnwwrkKui5T/8eADO+X
9ZnIbtbOxoKPGgCSPZr6pxBy0g/mdlcXSjy8NIL25ymiWauJ9SQ/aSpOFo0Smwwv
3cZMLIO+078Em2hFQVSc/gij4GW7+Cbg23TC6PWQLcrssmURcLTkn2/ePcB5Lxj2
ClGpUYb8/dseXiWvhrWqDgflAIb3tXCIzrEzNn+HY/Vnp+lX1dtswwXVaqgJQso2
t/opGsNhTFsuGomKtKKHZTyAlySB511KIOK9ghYdLmP7KaEM88gFlJmCRaOLJb5J
wPlVpLAJf4mY5cIw23GkmR/jHMhjMBKLTWHCFwleNSDIRJq7etrleb8SwRxnFKTv
0of3bG6FwfAHmn8CnvUHFeGS9UOOkSiIlK3+9f1F14ytJN96yg2o8/rhQFUE7tSh
cKPIYywrBmZDau5THGXM5EXkWc7nTQuyxdgstBtdy/roA2m7wI1yrIWHzDd/VZob
mUHkio1uIQZha5cTq/3dgIlBh6VTUTdjwcK/M2pzriJBTEKrMnOU6Z0fwf0N4M0c
SO1j051QG24qE4LzkGsLzqNIZxff/aRYb6iOnZ3YndH5uOPbE4/DYSpZSTae92Sm
EGxMSrWK+OG4DBUTLWOHkZlayAEHM+qtd+rAbWhyJtQ70aIno5mugn6mXZlt+0se
o9Wwbsye4qgf7C+vn3Bhh7GsY6oqZJcuNx0MOAQeRAvTkt2EwNMmysIJngy3buV8
nfTPKJpdCPX6sGWVyJcEBp1BA8rEyi1zvT0b0FxS6oWZbxToqxLxPj9riScIrXvC
IwsztZsyv+6yD1122itZDcppAR0ocnWxuIdPWcKnMJDY/NkSaOyfIx+zwtIqr0HZ
7bUIMXcF6DSfFLnenxGmhgL0fANZIrIc3PzJidomM5STnzioqYNOvxHcizB/+qz3
IZif6ly247J93+JMnSnoSfJO8oE24JUYNMJg9bKp7TroptumtZCpSZlWbrZLkw5X
a43M+RvV8t9CZBBXrDYUfGOB5pUnCMBDkmSjLCdMTYcWNTNCAlRx0m4A9tGU1hqu
dcy6REHUcj4cO+Gz5tIP1Z1Iv/AkHkY6ISgrWdLxqTKkoO0WlDl8/mqiSV3P2dol
aW239PMHIax+df3NMyyrsTG9L2qU1SsxFFak+HhJMSxH85YYsCeDObre8qTmV3r6
GEFQcmTvqltTdPmtcEqMUqBSr6s9B1P3NxspaK1SnWkAKiQ/u4pfhvxtLiKdvM0d
L86R0PeZE8tOlv/Q1Y7j3TaoOW5R1Y4eai996JTnPKfaJRHE5zzSomhIV4WkAnnP
yarU1/Ns/AqdQpIv1CUgPde5+t6hskOrO6eCAEAbp//n8X9EPKY4mEbvpnPlvP8E
deu+xQZktIajy4eUFWpkt7lFR+YpOW8NoL60oR4VoeHHZDkK/Eg47BX13WPRqvZz
qB+cxRGpQ7iisVXDggCO9Pht+ulI8+vRp2i+gH4YnTprXOd+Xeq2DGc2wnNQpu+P
Eh6WRy3Onuhpc3wsHKBKbxoL91Jge0oJ9ZXbh8DvT5AQfrTnuvaVgoHixDEQKovG
PpMboSAwW0u6/xZvtxB11qb7TetROShg+iD6mJoLyTVpVckswzDZVp3qYw07UYSa
eg6nNuv22r4pURNfL4BUgqju+m8RwngDXONx8DC4xZ9HV+fcslTO+k765FQKXLg1
H3iAZfQjrb1fNqRc0gXzg6GV7wfAOVW8QCNj11x8SnuvZJ6QQNsqktUIIDjUfOlE
3DiF0CkB+4mJAbtEdGwYRPUFuIWnYGmlFv/bwBOqcxLfXBvXGOQ57eikbFBEEHdk
VRibLNl8rHX3Cv9Oqlh8zNezo/11q3oqB/BFfV7fY9JWd5JgUHYWQJqUm/ir/k8V
xdlZh843wckRJrVUMwtxEe4gc4pteJmY8VfNQunPbkl+EnVUYJ6L1hzn5yOPsDDi
5GK/rWw9ngztq/N98VZg4XHzhl9Afj197vam2Cj+35pflf7KovLGRBDq84Ev8TpX
ydlRoVwvvyN25O8wndum4AG1D1SnPa4Qi7RFWls2oCtVvxsjtkN2IUOeuliRI++a
jp2V5vjhcgvuK6DnW3aOGQdfqpjSIBh82KOH6CxfWgFe+7ovJ0NGLLdYaiHz8K4Y
mvtzBUc1Nf20jZXe91w07DHu7+rjFogHlSWlCQAGoiY8qzAlpb3lBZ8TuwHpZonF
9gYjn7TCBAZiITjhgFmX/5CakiuVts1ZtN80jgi3JPNcNjfd+9PS7BqrTDh/hp1U
bV4NOZJm/oL29z57IlptJPP9RLozs4w75U2Vr/4sUln1c97wvO63cI6rBCBA/HOL
RPvPQiElK/ai/LImc/RqV+IYu+pgliG8T0tNrWIcR5hYFpA9/GxzSl4sdgSChYfg
XD5VWxpeFyFeCAuGtPim89SKixY1zS235NJTM8NP3zteVTwh/haolzz27L8ZUtAI
jlnvGoEoPZnRUxd89lLi7qqlNki/I5UdPy7ZVpgjqmtQW7ylvSy4AcWphQl0AOpv
ugSiW2ykkSyrIUk4XCpwawCFzIKjy8+awzz9HsUcD7rcS9GhPmSuvC9nUnwPyeQ7
h61MATTca7CnkZXbIXtkuZghB9HFjxfU4nnm+aZA3E0VvQj+GP+b8zgGLnROtRN2
X4CbzAdOEwjhSPJBxE6MQ3mxocg00XZbs6OEFPWGz3IGozhTlxETRq+qTDpobIyu
iVvjheNC1SCqXmI3TVgoQ6CrFIUQmOOEp7AX8aD2msqoRy70VDLgH4adJod9nFy0
JvqelvosP5+mCbPd43T5M1HRqOn57KxSe78YWpUQKjZn27da360pBpyycpHxL0O8
iSaxtfA+Ox3Z1F1N1fSUgQAu1iuWZ+LUKCo6Jzz5DXfbXpIMuA4iKXo5WhjEbRCK
0IwbQJ7itw463kSuHpdVxDYRlPGv729idv64EZZw5NgZkxfTgS6cH2rZ0jzM67iq
lRfje8edaMSKA5QusP5CPgDyRzrmfDpBKl9HFXGgQ3T9G4EXxbQszE9X/rqLFa9y
9N6t2R1/vmmNTh2LzqndM9ZKu0ZBZ7tK0cf7f3pbMK4XmSV97ttIRs2+1BLrhdso
aSmNjOKJ1EaoIPibkqPQ9el8ww18Y632V91H3EEcOFmNvjZmFm9mT9jMSTvDsV0w
e+ta6MFzbRt+mlT0W7VO5LlyhfDbyQ626UbRT396jezm5HJqZr5C789IGUgTFXBU
eV53issXWf4HT1qnD9DYuoscVqAVjP3wZnTPpFHZUozKVr/iHcYbBnBhiMnWhLA3
xQt1nW+/Qmq5LIbXogXpIOQ/8rJPqL1l+NyVJlTjjnQNHpyWgj2h0jOYnJ7FChgS
kpwrKGXyCObNg1C2m65ZoWmcOkp1aT8KhMG9eyo+M644atHXyZsf3AYz3ZmR/pAm
IvYHu5tB1Hm107WDNOOQH2x1CTZGqGzwmiuLyb0Gbg+JeICvACw0iOCYgM2KvDSV
ntRvcykKdb34Wdh2GRufHqs7wxbsJ0OpBi/4lkvHiFToeiy/vzpov8Bl+JwgprSa
Z3VZbkJ2cIni3KIPmnfQUf8bUXoZ319gYdadznnJly4DWf7DSO354H/5s98CHjFo
tNDH40Jg7KDojbKYbyVAvikhOSH5mIMXkJ7kAvM0rtinq2g1ddSXtT5CJP1khvu3
seXdgxwi5P2QOEuUy78GWU/Ff3dadS16n3GwIp6UwvXshZhOnn3NEl4N5AWvt3vc
DuK4lgh6vFTNWHSkKsghhwcvFfUmTlUuNpDe9yUNBGKJ+xWlv4G6vybHVIrE5UK9
0cCy9B7PTrDmVR4HPFf+yEidolvwiLece/QCbpknnkaGvcGLCzSqLdcyA90EBaOR
W0S1tLhOAGfhIcUYtEdoS6jTYA1uZQDanwAfYUsXk0ptRo1wscr6hFreWJWhudaF
6b8AHNWTLcR4MH4QdVaXAt1ZsSe32XdHqDWa6ckMuGq8LoH4F/EAPA0b97xqBh8n
0UxrZPZZZUgLTTKVMQBP1na+Veetlt7StTssymK1gO57hhIuT/Q4ak9wtYJogDsh
BxV4jSUX59k94fthq2IY87Vcwg6RP6Mv88+3wcU+bzUpLDoSVbPDNUFShp5o38cD
SLJ0OWhoAVWMbj7adiXvL1tz4wMFn3l6SYgaJW5MLqfBe0dDA1AnrphAhm4JwA6b
DFRzj9O9ewtwyzO9nOmKcYMsAOqTFCL6+RRTC36JHCNLbNVjA1DVGmp7DFNm6IjE
xp4OJrVyYwqMTBTgbtO9nH0N5eqdkZmppchBNVaIF+R7F2C5pTGVk4sUzYJi82HU
k7HjdHNNMsta1/E9iQAyFn0kh3U5wMFNE6Hj8Ab/CSPyOdvOI39Te6+ovSI33rhv
jiW1IKA1qaXNy6nWHbKdzG72zRDIDqIs07MNjm9EJ1cOZ/tJMcvaoJD5RrhJ8JgN
LwLT34Wj7ODfQJj/isH+7SAfbOkAPEupcaTS4Zs323J4tg4xSqZQjqDS0PtpNdX2
a3x3wnlP0wiwXXgPcRdaRp0tfC7yCf19pzqOdrSAlD0xbUPzTGtv1yufJHbyh1y3
xtMxmqXA/g/v6ofOMrIWQ775Lhj/2n0HPw9xIOXEL9GuxvALyMEgv099pPVIKTvX
DwYQC7l2MObBt+objs/1jj14pO0HnNI5cc7GwHvIdnzqwq64Ap/2xmJWNYsxrsmX
m5hyfTy/8wnzNpV2O02VCcNxE4VPY6896zEWd87g6UAjZGX1xcKok64XUYaZRS76
fIlNOLmlFs6BUzGFRPrPLA+VfwOc+2yd0bMrLuz6UA4W9QC6oj/x/4fnHNJUkr0w
6H6bS+xfeGaiXw74mokaDy10uiGzGWAl8N/LBXKuUJsvaP1qT4kw8IiWI/bsTz62
kMRTG6fn7VHy2sN3iXU3eXLvcHytvb02NkSnBEbo9Iah+wRkm+UvkoEf1RKz75Hi
wlcXhskHGzHZiMRNeFW11soESDJ/jZg7wAboJGqxAw/IAkxzznmyHgLKC0H8Zq+W
OmiWvMWq/uBK7eje/lflSwYbp796iMtgIgrjfqM+z+G/3ooyy2P+BFkfSQfs1OOt
WrQ+ip97zh+LTfAs7QBjDgUrxUSlWOTguUsl2CbLuLSnoOYpvKv8LPeKrWRRdYu0
pItoCC87AwVfcmQ3568dVVxYI9LQ+1/OWKGM3umcnZ2NV0LeA/vq3N58a3vJOqQi
Pmb7lfDDx5HU2G3NO/G1J1ffXuohUbouqiyTUSOQqtHeBDwAnTP00rJfCOyUNPiZ
AbVsCcF9D0o4FyGum7Cfu2/q3/YrWy/+E2bnCKsIe69bLniAvq1v/EHCgwqmf0dz
0i7Q/dwQqyQm/dbWKm71aZ2ZczVInaxf1ChsKN4HqZPwCL3GePe1HAUNb/sI/Vhq
63qKZeMg7cauvuFpLTNCudixD6qTRLQjFsD0HeB8OhvJ1SNEfrfeCNLuM9MxJsKn
sgTjPGnqEH8Ttypr+jQJ1RAz4nuFD+XcgsSdawYZXlxE0CjVFeeOUOl1xVnP7oil
nI8/qcXiagtc9csi3OzrBFc2JDIGNOTt2dbV4lAyPKztUHn6v67bwYZTac2tiCPp
+g2s+qMdXxoKzLCei63CigKO2VhrKRFhi5N7Hv4usLwjz3iKsJD1geoH4Mrei0Hd
r6Uo5aqQsBFl4D8VtTLEPGcVImcEMtuTlauCoiVX9um8O0TciupHM2LN3C/wqv/9
s/DyVly/wDpih0rNlF4Vy8eu5d1+lDzjd8q55Q5lobLRNOeofuYMNyQq3GXmN+em
nsdA/JkinqEscjT7ABhEPzjeLKWCukPNRQObrwnkvHzAXsMQhn9F34LbMU03QnDO
enEhHv9RA3xtElVVqVTIaII155SNhNTvO9yzGjTAFxLQ0iLOG1H3xIsIMVEDS7yh
nU75JgEFGKeBXbr8CHHXjEWoi+OVbqApWRgj+zZ9pogv+hJD2W4f5vwJVj50Yi7s
PU5VGh/q+V+rRmldyZo1OTISTt81K/JDAOIBreAJkmsT/2PHWhj4zlYAOKLMayG7
AdCOjUH1GfCNS2VyvpIvHzM/p/6dplHwioCs4udCKXLa+qo5mRlSRC7LqBmxoR+k
MRjOB4HqYEeX37Wu1i0L9fTVkc0cVafOqTjubKpqQh3HPaPzq2ABUQuqzT3XQvyj
eOX7FBfhVa0HhNnk/ENCxQR9uW9GGY2EPsbVaKH8vi5Ng3PooHgngqwesTCDB0Vx
3NT4uC/tZPrmYZL8bGoW9scu+4SQMe7VY+nBqTci5/sKjXwn6AWDzc/3vmkKpGvm
HvIguKtTtjt4XRXnKAXG1kq8YmM+yRPUXVDpQHw96/70uZwQCgWcwbr8dKm6/BPG
b7HobPBSYEMyn5DU9NkHSX0RjlUvT78Hga8pRrsRX6jSJgHT4lmOobTi6eYJtL7g
8bllUGhGXTxRXfceIMPQsx2Gtqb5ixr6be8kNoPYvaOnJ+ZlFDCLcKayL31m6mfw
2Dva3Ld33i2AlVwZfQFHFemdoIP+hRqvTLLr4K1BmmxiXsYWH4nOrCSdw8I1IVAx
NE6sP/Et9icJj849/k6NVgbrvL2XpiBkvsHPMdZE9b9oxhUFnG33po1XcYbxaZsf
GCrzlR7p7JeyTkz5MdHuFYTQoCSMw0tdFE2tAixARuAAEF2aNp16KdYzRXPg8Zj1
x0h+yISrntmb2BftaXl27+kIvaqh4mhah9cpx3dY4H5UKF3K+73Nhu6JF35sTpgF
8buFm/tpKdqqf7jxdSCVNUAHepYx/dD6aWhL2/KSVzxRRn7LNrMdCcUR+tOUtM4z
QbuHFvMyZa4B7vgl+DxkXap/KocFVeH3nFds8Jujbo37/ZE+fzVsQyuAj52icZqD
NiI1xqfi4B/TpECWwWNsSRZqxT54WxNwOf61h15LcPiMYuGDYcA54dASRNUuD1q1
q+mMPPjAO2PpdAQ6a1pRUlZbMRXfs7ZtZImXutEVpssQPwvn7N2DBQIVeoR7qJk8
1lLl/TFlsuPGIb6MxKQXzLVKecmE1RklwfvCHzMur7jIl/Kkn8By0r2FIAM8TBOa
HHPe/yIHs81JIQT1UIMfHpktbzXtgU5D/NIhYfW/YxEArVgD/6ob0LKZJqnP7fAU
4DI2pGVcXWhJwWZED9/TpDSsZZRImaeRzlrxzk+HA0CAGSJI9OV64A/pzNClBP9/
9DIbPuirMu5EvGANxhV48igVaO0CHv/2X/sGR47HjnsKk4kDTh756tnfklCkAaPK
3Sq3iENz0CCAJqzeBcl6HMmPr8X6ONl98DneQaxlsjiqcz1T64M87twZLX1NY3IW
BDndBTiRRMo4i35MUSV3D62TPr/snqPfpF3JGzPArdP6IRBL+4ChQ+m7Yn6bQiSA
Bzq5QKv78rIRLMigRehClW5oQJFMicLos11oUQE3QD8mJ9K8r0GI9vARrTEz/A4l
yyylTQTKc54jcSD6KPQlynDf7MmH8U0gUjrm6W5h9fSQiBXH6bkgVibrtPd1nWym
Hy/1iGz+tOlJVh4T664/g5MTsBF28MMoxCVdhXY5GPLpeeOJorneycW+6oqgvr0v
QUDKCqVm9KL/NXmTG2P41U+G05p7vRurBTohqEHheqOR6RAd756MkL23fBvLBCws
BL8yKNzUe/l3xVDEy9swfVbkgU8U936OPlQxZccDTr1sC83+rwskf62d/EtzPSCU
JYHvTuLtGtcN0veMWqKFCE92rV0C6gOJdhtoeNWXz3t9lzDOgriUopQU/I1qgXrV
v0wv+sBy1tKH3DubvarvqtpiaIl1x1E0LF+TA16u/vt0a0URKsG8kBDIsb174aa3
dxTVRKLAfqQikw1Da8qj0z2sIPWWwf2ipZ50Av1Xld7g2bZjT9DFRXR1neDyDVz6
WTj6lFr0LHXQ6r9lU4vnKgKpInhGW8bTDFddvjiRW/vcNS16R8wB2YM7GGCaNeft
cLbFYgYcbbHy+4UEJi4njNPNteRUk6T8Yckl4hzbyQws4j5IMN6AcZg2Fzv2vAiV
fyi5jK96qdDQnezptHI1IiCWpCKR+HSXRKULuA2/Xi+NhjVvZeknbv3/NnJi9JRP
6K7vnXwj9wSyLkFHEs3jkf9GP6+0PHgpu/YAlOkwLgImgPhcWJV2aOkf6qcZDeYM
lVWX69X2iOcb8Sv1nLiu0wIwrhyi6RmrI/j9NF9dlH+5oIk/9VeVAGZPzdIPr5Tb
XTplv+e0UgrPpYfsd3oINxcCLeUGgQ5irguZtzHRZwZgG3FtsFqaWR2jQzGxfwBt
Jb/OyPIU4g13cO9c1c99JKBr2DdgwW21vGSytIaqSaxJohlK2enfK6ok4g96B/Qs
qrMRrQwtD0UCOGOofpaVfjXetfNPM0cAfOVoiDil2mCLBXsX5LxJd7TR5D8PQCHj
qYh5ebuNI79xMFwwLPXc5ulXDAmlxkU8qMF/AvPZ5hyj5OVulpXnGExZsTfRoaQa
8ZU81YmL8C4ftweT8HldUR7evfePyouDVd1jJ14iRoClTJRAFdYEavYkVJp0YXIH
cqaSxmlHJ3oUd/IKflnIkLL+eAJOV3txSjYIHuuzBa+pQGfxQ0XASxSWqXuKGqg4
C9xXQnklZEQfEmcDAUk1kTlviIJF65UoI4taETwCUIZU4k37MdloNobnx3kNQ4WT
sbJSw9vjn69mj640McMmx1PY9kLcBSUhpLRmZR18D3eldsGpJR+zmjf2Y0qU34KW
6freYNy7si8vVzDfq8lJDiNn/LkL2DXm1NbtHtvf3c7XIqySQA65qluyLJ9UcLRR
g71LjuLp80RvNN7VKlMwfDjNrP1GmVqDkmflsJasGf7KljhMCIrXWKL8+Jw46WMm
acYeBFYDZZv1Ubt5t/Y7qbTObpTAJ6Sd+whHA2aQsG0r030ptTlrlSoJixy1p1R+
mNlPnx+XTcwjg84mqdY37a77WQmF62Ubzc4v0UJS6hQ/NrBi1b8Fbd1e4tsorL9z
CQjOYeIaRRMABNDIe3WhZpUxuGEo2lZg1MwmDUgmNUAEql9lBY7LI9S3acGE6hIi
w3kRujHT1OZ50ZLg3fs2TlT8Vhf4q9qAW+kfs/vfiCkLlo67c/cjkXIgFhcHMn14
oxpf5HAXm509nmqGaVyfs5FwwR1lgRYPj5G2EsrpKEzmVcYWJE5dzz/0tZIcEVjQ
kSUfLtT7nObFiksZOnD3MraGbc0HCW7Li9eJew0sH3D1E/94dULj51rdeJUrTLZB
YDSaMfSTLL+N0doQVLt0fbwYhqL+u28B132tl3Rzg+c8ksR6HpaczjY8N+ObToU1
TJBk8xBxW/x80T9MQcHCeHDd0MiqQ7SSUPx3lYC/wP2hLP+BxGEAGrs8xCiO7dbz
BnNLA6oNZ+GdblQZhn/u14cgqp3nIAp94VYP9HtsodaswyXDVSJ4Z/R8686lGsOg
4Ia1B3JmFSNigx487v+1id0bFXTIKQ9tx+6cX0eIl0gGyZxxDWb8GQ3aNm1OzdJM
va7TGrESObT2u33vUSxvpGF7MNrzRXH8WtAgKwqVlGXHh7cl1mhvcLE1sVW5L1U5
PwzZcUG0DvETIl9Q3V4XRE6yLF/xDVzNGQqia7GU1OeszzWrUt63MJ/zmKwt64E5
hpnqr6KjjmwpNfl4JthbribDLitAMt008i8qbhAdLHO5dO8vb1Qfk3ReqyTM9Qw3
FM7IF6AP7EIPEvQ2rsnY7uw458OQ6zV+60M+6ZfggaTMv2bvx9GJV9ArNMQsUQCm
EMKrU9ReCn+xyY4YRIKPsW98Xwi6dPzhf356DxsvEc8odgr1czJJtEJDzm4tJSpk
Vetdtcu98Cbh9Pff0mOy1P8yvdc7oY7FM46X0fNGorEsAEhlMCEyIcKO4B8V4R+U
bzBVKoAhGlfkBE040YbRmEkyMYdHbXD8xBJ0YE4YqbG9Dc0LfBxaDGuShSmtMi5r
QOzJPWM6w4jbbdJz4//THnYHS9428hZV6dLekCPsFPhgXlIHKjowRJD5E7BpkMw0
FVwa8zfO5a3m58h9dy082W7GnbSz3qE/Uitf3D7R6FROxT+0UjEqThOsj6DQm4W0
cDuDG35meZl78ROjubvP1/Z/4NBvAEzk6m1FXJiIFgav5S9rLc16hGkN9pyFheSI
Am8tdJFVU9aXdHACimaOAwQqlXpFmFcrfmqKcGBpqtWJnT7rHxczg7EM0fTrTL3p
yr7jR8vofE5z6+4vKkg/UiiufV2WcwVf8Pqu8YkpVCB1o4Z/+UtJo1ooFjWCySLW
E/5reerLKenob/OwnHcN8GfXLGUpjFTDpa4ktFqeS6sX7iuEePuOkwnLsPF1ZAtJ
DytZnCfFH5oEho0MFCOaeOrjBq6vJbKrz6WJtlhCGbLC++yUg7jAOX4MGeEXvhV+
HNyaQA/YGzI2xNt3NT8aRh7l+CHmVqtCiS9l6CzG1dsEmACGquINGs0L9abcMMv4
DIBpWm0L87xAnnRhSLi+eMmQ125tCEVBaeCQzWoa395dPIgc6ZDjCczH0o+8UCXG
sA28Dkrs18rd6Eodkf6VmDtLamB4TrIBnQAyPIMdsNGJPrNYrHU9SjAou4TDHvG8
Zkd3rx2chmkBqmapul8M4Mr3VpxRtq3rR8DgBAUoD4WpQgfsgIgZLqRvA9itK/1h
RYiDxBZTr81ZGQPOcxTm8piidkZof9lH0YHcjbchnu7zT/+Cr9hI3u3M17xiA/ZI
Lq6ubn12VuJBw+Ib7SD+IGjDF7/1/yo2QHEqoOt2wQwXwikJ5riOJ+lQg4mfjhYx
AkQBBayjNY95JQvVtUnOSieDM6rb78C6Q7E1COtUNSAgc+rwJp0l6TfLVwnEvt7n
QwXAbs7Wa3NvlQXSu72OxqM60OM9RfIlTfCMoooLeOYh91lUq614eG5Tx6G6R3U5
fHr41RFCL90k6+rK9zM6iTXipJLZYDP3QcYfv9OiTiGjWOQ2vhhYRcdbNS7M9Dvi
ZXvRBS6JH8Gq7hMI6iMQjpNpGrRDD9U5qQXL1oA7cbunuiXfCT0NwloEg9AD/g1b
HNbb+NAwrOC3lzpSvvBd9aAdfHPt0fBEnA3mTqDv/o0JSYJuiwxfBpe2tYOA4QEF
lW3haci1UzNQ5oXfAbySx1i5nU4A6cAlhYHCcHNNojVtdDzPbqh0PbPBwpDqEXh4
90rHylGqOl4aZyS16RAJLtWATb1MOHAOKf1EV4VXpMjK8DtSWnt2Dr7dap+9En8x
Wz5qRXh1Y+87Xg3KNlVIRD7oRUS2d6ZEukbiUAAu1zv/3N+/Xi7rW8TQ8gM7KaPY
RgAycfUo/Wvt+1CgtC8WFtF/Dm+hG+nbisnOszudu/ot46wprEi6L9wK42ZtCfOf
dVJQHmVyHSNam3ZR8MQRT491NmXbrlERTBeJJA/XT3qM/7uolLjS+ud5nHkmkIzw
xfvYmEyhkov2dcViA4/F8wXiMXgPrN/VGtDhiXCSRtM3pb2mRE8n009tVlkAWGmo
++++3bQ2UaSJs+6zb01r6FVK07Eh41cO+4MoPbhkPiIZh+w/PxB5hP8DI9Re/R2y
InSWRO0nnuGzUEmob+S4QK3QqWjYXrr592QdRHhpizeh8+KeZeDS0lFH8voIh9Ht
dFBir1TsBe9+n48WsKonI0NZAjE4i57t5MnNymUXI4rpsRC9X4DtMCiIOyLj6PUn
daX2QrC1ixWiZebgeMNcjWG1FmxtuJRdPcRex3u/Q8wdkwrfVeIBN7a2WhVdT+bf
wv1ztlofAIFoUqq3BCq+kgOrm22Ezs8eWnOD3qPN4sRHHtFSxDVy9HbZfp0ch21d
/6X8Cvz6SN3jExdF6oBSOnq857c1Qawd534QOp1RhcKs2kX26L3HA4oJkHc9nbuz
T4/F9koog1I5YY8S3YZq3ZJyc/ONdyGZMgo8rcCz48B5Iliru1pXzUtIOqE7izoJ
IaL5q1HieeYP5rN8d7mo1jxYqx169RYtQrDp9sti/AWR2EcRv2ts0+iAFGfcFXyY
NTRP4Z3uPLTM392cle/o4Y2+PkjPK06geYmSWNici96FrDkgm5Mz3ATbyWSH5NNV
quegCUwiyzTBXRndchq6ATqyDBf4gqSVbq5fhBSf+2+/CFxZCVh0L4m7Q78Rju70
P3MTdM8chPH3NyrTyt/7k7bQqj4eUhtcfX6HOFjWKX8bPP8AVVrG45Jc+JemckyX
sV/tVrsBxpu+BNz9mvMpiYO6bpgGRcpHIl6nJEZK7qHDjJ0IWsLNi3HKTyNgTaip
6FcMhT9yZxusJjK33h9z9QK0sP4/e3Nf9Lh28M3D2bPsUm5/tWsTdc3PJbR30Srg
x3djGSdBNaoFqgbYNyT1vYp2e0+IuqSsLDMCh7oJ3LjJEDXGWOU0UZ0UCFrDoEBT
D6fogZ+dd4TIoFP4LnBF1OYFaoCDBgN40Y61Fha2LXBa1HH3BcPbJPr0meYTZ0kl
bej7cYI2OiiKosKPonWuuLpo6xLnpxl9SsZnAatDaa1j8LZtZTTZye8x9gQSxtzP
DGszzhS7A7V6Mf2J+/QAGZYNUAD8rHLfqkPqMpmLXIQS84pmpDKpO2FMO01YU1e+
Jop7n0v7PUz0IuDPP7Mx+ELeMW/5KC0LKOGzcrm9dl3pfFYRwbpBPiXpclXaPwt3
DFbHG5YHB9toj4Tp9IvA8bs5eqRn6RF6l6jUopG5gFY6w/kAtwst7IB56onXtpy+
5v7k2bGaIfOwUgN/pxjoD/REg9r2i7ljeVrxjBoEwR/K447LPMIDwxqFXf+6mVBk
ItpLnk32bnX9ibcEw9G/nU2/owVycC6j6D8AQIfRej9MlaKJl6D2llSHyKbneNWa
QMpa+XSXk9qXO9YKR0wbaHNaSey0HI+vE+qAkiXxibHoua1/Gxf+vsSx2k0vLHly
NgTsVqHqHS/goLxW7EDMDQPq4PMSiWykek73P4Xar66CnbXs9ha1Ts6dbLslyV/K
id9tM9WD6fv1kE46gN1OAakWU/lqYngqx8jkzV83GkUqcPNfap8a1Fcq4soT414O
HKc4jaTlmEN0MnB0ub+VdIcRuIhSi2LmCxU4rhdPK7mlFaSCFymyp1M2QrdOhD1S
0ojRdDRaCe/yD4TzZTBvsxOL7mS4FJk0Ben/RvkPA5drBNzXjv0b1ief7t99JTOR
TRWsmfLa6UwCtPzC6Oeyo4+IsbsFMSOCClkZYRMzYiGU0jM+6X5w9BQoDdXR0wdr
Yo8AN75sZ4XdTElgmrZAK31k0AheUDs2Pg43Nz/ZDBqtCfH9cuh/Y8/Ftka+PnSR
EMNMhfVm8gRhhyCDCG8oMrBItrfLFn4nVJ6Qhm9sXMU5FqcTMqaTeryywbn1Yg9T
++8bFkk8eLspUD4JNXrx8C30i68ZrB+EUejZRmNy6GHxG0aga3z67B/R1fX3Gwby
6XS4yUR+9pXdWaRoGAqZvsfI0pjnW6u8ouX4NWwzk7XBZNWwBF5q75yp0VRxbdKh
nKGiSqQtfBVcI9xHtj4KRroc2lhk0VPdOhvJYDWMcUmGsTvAgA/TOUrP1CgUgul9
haIFSIU07TiwTMAjOrSTgOn2J7RHgPM7sgg8a6m6OBqTU6l7S8fAw36sCChGsiEB
7erfa0SBobDEQlfqurO9voXZs9E3fsOScehNO/ZBXAlqSVc395mVlckJqmk6fqAG
3Gum36Fgp6q8jl8nkemT8o2VWe73yfQ0lrSKpmdJSbgU8Hgi+uYFzEEscA3URpsQ
FqefGe3XPsHn8vDlaLtaVzrcMHsuHE6sVGQsVnfKRSvKZVGIMQyVCeZ3zkqbiADF
SYxVuSdOUhVfytxYh0M3dwSrNHMVKnLG7GC52ryIHyDhn22eG2Q7Ly02KMoXov1T
ZcL9We1bEKzpUqI5oNeLiKahJ8e/9mpJ5D595BTP6/4a55jGsv+TpW5myPZ9cvne
Fv4AVhbLz6QYymEyXX/RJgqRpc+kLoPsQHNXqKlfYiJVbaA2JtJw2JMFEq9VXp5r
gB7rdzC/5TFrMS64VDDgdz+dksBSpjpL54m6hPvKLyk3eJNWUu4no2Z1jEMj6F4H
dbT++DJlUEGm1h2gjYqHncWN/Q4RTrxUjLdy6HWHHs5hpsV7y2BPulWxdoSoJYXM
Bo78Y2VWXBHdJTtjWKlzqnn/wceoIRyQOrV0ffgIOXJWU4tE0yMmtoxVi/yV+bui
GFi+1XTFwt3AKFLyzCXPMSkSuAB4BUmabnKqE8yGYLKtx77AhTsqGnwV9JhoZhuU
79xgBKT8XztJMUj71laXuMM64OpA2Ji9o/jnn/m831wweTWUrWTZ7ym4O83qIe+u
k0VQ05rT3Tjl0Y1g14a4aqtjZFSXKbTRUD3imr5yBQFJuTtMeS+xx2QlfBeiMJGz
/+/sJmEnqkCkPwZKUTJTnDkU6kpUiCoT0YGb1tbQgfgAvmIQRx3fhlGo5MVGl0pX
eE0W2LJzE2OxJ9t9yr90XaEdYAqScxAaAM42NhAHsNvLovXnw31fPM2/qkNx9RiX
A/ku1hABmppt2wCzjlHb6CrzE5ililfh4TWY/5y3vwG+K+Zv6zeMikPXFjva66l1
3N5GAnAv6Tt8fpuxJNDNgWO5h18vjNDj4mDSxXfBjqpxovgfKBfHkc5BOz6EkJ/u
qIt2H27qCrAI8gioycFRPZNeSZ+WpPsgZxhKF0kWufQx16wZ1m/hxrv6QvOohWjb
SaO6dm0TCvQpHttC208TCuMP08/iTxtEX+CDzni57Y0XyDY0VRONLHhx0Ni7gz5x
tNGDLTn9ui+U2/CyHb4eOS1NtHt+GeP/JLIL+/sX25btilY/h8mhesZDk7JyA1vL
CbftrjCwtuTF3Ou4qMamNpjIZsYzpTclh9EfYhREHmzJ09VBi3YDlgWHp4eHcJ00
fm9Yz4S051otv+i7hwlp3vDexKFmfusF/RSjqEPRNMwbXSTIREKtIt6d5vR8jGd1
EGD1Jyy/6ibsjMMZCDi8yJ4zpvE/BqT8QoXuOy8SOl9MJiHLZJq6mvHIDT990GzB
pPGMaKo2k/WW530qqvHG8F9yk9BHS4JbalinDLC/nAWJI/wc2z0dilX/2hVGN4QJ
WoPNm5mCm8ZWf5AuOjXlXf0GDGi50dBiaqRBZ9fh+cncjsLFjQKAVgimSov5aHCZ
eo2rLznsYMJbllU2YVTPmyjkcA1LCYBclkFjqeCgpgP8czGQ+Hnnbly2lu5Q/9G+
xvZFknXvVNbO/7BdMq13qYppxLN04hO1YM+oWNCAB/IcL+WxIQWYBKzor/a3R0gq
vdquiA4fPj/vUEeV5BxolqBh4kg4+B/RHLcbxKzdGavkDtml+WZoS3biV4ari6Wj
wGEQnfKVhxymuQdvuUK9Ev5eNt1Hz8yPcLELijIuwc3j4fVpP5vWOb8oeezwIFcG
M027yQ/Jkd9hxf+D7VDZZlb+VskCuMaBGObQGCcCK/PBcMaGu42d5aUKtH/s0Uip
bDU05YddIcPe5Ms9/3Sdrga3o8EUJhWKkXFLWS5hQBMSSrDTPTeZzzl637CJOEqz
kNaVGiY/Bxx4LMKNe/hqT2acWwGPYQriLSMg6L6vXmnkP5z2Bsw856iyqobHHmdO
Wzr01hikOy383wSpkHEbKOGY3LK5R3NRHa/2Y9jj5C7rzfVKARZf9nkTgXUb4KGn
27rPLxYZ6qLCLT7AU0QqMQn/Puw7RA0nwOsU05vdzUT1rg03jIzsX81gdJoFUhV+
K872RK3a9l/Ls7sff37NATZ0Z6zqkgmlSWMXP8x4s5ItQersNJ0bvtEl4cpowr6N
RqGLDXVYzjsN3eauymSKq/VLURy6DEmV4XcIqmuskfcBYQs42wdc5iFax5oazbEO
lJ4vz6UWcZr0UcYelDowBO89rgSps7rFUZjibh0yZYL2tA7suMtaAEc/8tWv7Hve
+k7pnOmXpw7cakgp35B0q6Oyg+SABLHb1gkUaxFwTikxEnqoQFUN+XOvpmeY74iT
OfGR/reJGpsLHCSe48eptvy8y2iSWXkXbdkqnWSFkfT3nQxYOwfMeG6KXPJE9sJy
vKPnlybY2VAa0BP9ILWwRWZcNmZFwfTQVW31UsqMD7aEHafirSqetl+l9BIxzuae
jTpJuUMDdIj1FUZaAQC8PPIRIW6ecnXNSyczLJAIC6jLaPjU+l9u3n7j8MTNBey1
Qb3A0pJL3e0HZPoutuTiSbc/JL8WLV6M3r/IpabEQxtNbFeBhoQrirddQ/rw5h+l
WHH2PqNzbHkIITQ/9fluneIDIvTJ3HbVIPNIA0Zzd+9UnbmjWwMmLsCN5SyEFmKF
5vTcAjFgg17K8+Vu9USw61ZQeYdgeTO13KmU6ts/fu3z10Hn5bYHD4I8+LLcLBB5
7mKrJdf43v/HY2Il3tkUG+Xk4lgjvqJDSKo7pwsBT1aykhv4fOumrNsga2JvZm0g
kmghqXKwMPHM/iFW6XgfQ2otFdbpvjza4LoVCftwp5bY7E5/nzBy2gEYkJkOiM+H
PtfZb+n3DlhAaMpXj+sa6yWzjnS3zF91eOuF6MC1i+9/tbKG+4FT1Xl/WqaALiAi
kv4xErGHjXO+vVsNRexaj62JrCmI54XySJNzFwHioH1EDAQKrC2iC3OaWfiMON4p
UboIswD+HgbOmg93RUEmV3l3ywTj5EBMTVZA8+qPYvMQGXg7TgBfwHxPkSUr+fII
cgMzQsCeqKmKVirxAOLvpkvFf/24lyPIgovUNzsnynSB5DPRGGkKp/qYX8pe3tx4
sOTu5q6CdtfGbVtWFtQPwXJiLsJJrWDrFBnHWAOriLYuKpdIUSxgy2v4jUDBtaiW
iYjKTcITA9eWzSstmvyxq2AsmAMMvr+uxyrnWQ1JZ5eucWUlSbdNIWmbP6VVUgxs
DKfp1f73Xw0SZRZ+fM2QEd8fBg2NznMjDU4kqeyBLym6doF900qx7wMEH/8+PUaF
pVgNkZVCOkgmVTm3lnFCy3kKqkKnplXSl2TbGOx/xPosnKQtX5BFWkf4TEfnku1M
Iy4r6OzlQZ23XAwwAFBac5uVKeRVFdu4Luilnex5hN77y/haaQt1i5Py7pPma/B7
O2kEGk05Dw0YLS9N/Dy41vQM0z7HCjVFqKfkZ89o4oo4pFq7AobPTV9Ovsg1OVRR
RbAjdfQCoBBT7zG4WCJyY/e4dVerXKr6Mm3Wtr0lSR33nccCffvUgAPa88b86989
bYmRBgjdyVITPsqCrDb9EGP2m0QLmdjinmbewW816T/ZhakrPmBjv9Grkav2fFl7
rKYoxt3qUrY+Xv5QSKQEMbrrdJSuTIlqWdo3zIKwRsD6VXlErcOelQwY7eS+ZbOq
0CXRC/6mIOnNqVZqdWwbSQ4xyaD4BffU9KpBRYKrQ0eZMd6JtJYgiwW5l76e/4wt
/SZAVSrYwLfiId0aenH7uWCGTX3a30ZWsTkOvQ7x7Ckw1uqT6+prhEnkWGAm2uj1
r+jVBii0zrFqwvRoibF95qiaWkMCte6/dhXCu9whpoYd0twVMDHTBoFIAAyQGSeC
ncpk8qTwAex+6eu4ESzGK1Hvab3iM0ZySUsExKTgUQte3/4kVdieR2fxIrczb5Cs
O4DhPQP8fpagswC+StqSQk18Ll19NViDv/h9SAaCXg6DcX5vd6BlKye1Adu1DIp9
ae5T79P1MygwIlE9fEWqGKEqfgw7pMIoepbj5xZsE5sclQFVefdjwWPgpJfsR8wy
Zb/fpZwAkxj6SVUnRnj3guEOGVcHWp+UcSKGVzREXGBLcK7/BeeGEJTCp6iZqkvx
pco9dgsziX/h9TPWStWJDsT/ilh9/tRDy/41mmIiZU0vL3ODZapF8v0T0wqhd70e
WMAtDJkkspR4W3FlrOmvTHTEAhFK3GkMy+71TMW0mF/DD9xzug91wx1fftmns99x
IzaJE6ffwYr6NOMWpn+9ddLIjelsT1oNUl5gaYQRSpDIfHNv46hxLerunNeyV0TJ
KaLwPaoMFlQIUv/kk+qkC+7yyan23qtkBKZkbSs/HLiGEfQL/nrOnZwp7KAH9tbs
izVXkh7OIiTO8ofvVKNOX74KPqQ/o7uDDNw+l2ZbUtLrpfru7co0HzauXyFUbiCR
o2oNIgPIyOYrpkwF5wxrLkJojsXyt5Yf0jcX+5/V/oSOBwl4sJP5/hdq7+7vftmM
9J4eJLX9VnbX8R7WEDACOPMSBBv0dIGiuTU/8Y8SyYrM8KX+aFPZQ71qzBuAWWk9
j6mUkiHnTRDUjPaqncDdmqW7w4gBREomsxphk08zra9bo4vYSe2n65+WfBasVItm
XEAyibZ8FlDNn/AXgbjiBIrgqEzEIygLVITk6k/oeF/l+cpL3r70GOqCkrT0afKO
IA0NZzsYEiLaIJFSKI6/mrHWm9NXUwBqmforBFfI42YKym1OMRSUrD0njAU5dKSX
NJpgiAVjeFbUBmhZ4qi2wmsNAD7tyr6/BAXKh1MX1B2jiAfd49iGu+w1phr5ExHh
1zb07lcg0k5DY82c/KSjDhSDpD7jsU/377yBbafW8ovLOK3PFsJzAtejPjN0V/9M
CtIp/FRM4l/E/VpPU4n/4a0vd10Q2rDHB7Qz24+m/i/PZi6FIhZMm8a7fHkH6+rB
7xRHy6JytzZRufzhp9DGhWfdadtQb+VBiiRKKWQwOa5MsAcl3jB35pBQxdpQu1Sb
lHqon1tFw3bzULJFuO39uHmkZ7DD5VMzvySOv/AVkOeQqTIQIOru8cBn7R0aNVAs
2Nw9iKr5L9VirWZUzqcLmCL2iQJQUPVXiPEvkV1yHi96BOa1Sw+1rHHGKunwZBBv
9zhBy5JjH4bjHiJnBaN8EGJxOul9K7QIVC12nYnvzeBwySaNspdlCLK4lYdo/0yt
sAYo88R5VLVDxY/3YrpuD14LTHqimUGVT3ACtsIdSS/Qxuobm5trtGdJwtLN7mBL
0a1OJFtZsVdkWrqvaPfW85EoMhnHlbU9EivB+cFopB4eie8rasXqLHYo7P4DdMK7
pyCMUsSK9N4m7Nh2LuBM/Lfc3KVQ8IkfR/oIiiGa/jz2god/TNmkySP/jXAXSBuI
Lnt1yHLeSYSh+q0in4Fy5zHbyFpF9rDlFE1rmRGTz/c2MfOwOq6FsVeDEWEdF07L
jtrVnwrH4YTWSgGXIDUN2qKzECM/tM6P9AKidT9GJEfAB2WjmKFPkHekiDK15VSY
mQpkKB/4K6U1AWNo7Qqm1/Fh55sIR+5lJt156yl0mTANgSz03dMrcei5TibH3ihe
dyMM9CRMb9yEzBtYmZPP+IDRHEcvZmT8K/mLgaWyloQ6CCGDQdS9VZrm36pf0wQh
gMnOG/7dXFIknzH/t6IPKEsCdf6KtqWtee4qzyc9WhOfsiHpsXvAquVjkCjJKEA4
QCAloTkjCHvMEJDtPmU/W9qpD7k8EaFNoRVEc7akg16NY8RCwZJId0O/BY9ki2K6
c/ja9dmhGIvx1GP51Qtr4dIhMOZKA6q3wxn4rGj1zJ5uUGopCOqNeJHlafvwiCmj
NMfOL71ZOYKwJMX4257PbkC1mz/ic+Hku5HTUkwduvVKy+clV/P+KBVhnTGCEEy2
KJBPXT9JVcDKsdY9LnfZASBtxoSrA1csrgka5iE/nrG/t+jWz41SCmbl95g0NUMn
667D9FO6Kj/CiZCP7NHQUDoEhIBnC7YM0Ge6dV4T3EZ5QkxKkYe8uc49dDnQu0C5
zsjgP+ZM4mYg+qht3ImhpjxIv9T48iU4GkuT5DRjdk3P9IwLjqonSmlQDIA/e/kT
yKefwJkraW7AqV/wWkPoviml041yPCDBGRI44FPKidF5xt4TorvMmArJVhcUMNwm
uxLckVmbgBe67x0DTCY6WCTd/QshfBURNYbRV7JzyI3NRYMA8Qyq4Cy6Y8CDlcba
mg7ulBxCuaaWQvrfRJUB9aS2QEgndFRQwvEqCq7e+HJYRHG/8eK+0PPgaM2ySKV1
TarRtXlIGH/qdkzHM2dsciFzslB2ts+xLLNEiO3n6Kr8fpV81BA2uAP1kJu/cEOa
ybArHUhGFhxl8z4Ag5AmZhxXHHF8VVFRtSfxGfSKmaahp5RAUd+7n1uTosnJUMU+
L61Dbc17cuChq9ChWaO1W22K+lrrniye1SHQsTI/dodsLL0MYtI5oMG6rb+d1TC0
4S7zvri4+sS22XUqd/qijU+Dzgb0m6qa246KoHx5NrU3uN7eNa6o/mw/kMIHxQv2
tbYdWIsM098nkSQTkyo65J18q1L+4pwBzZFryzg78JGbZ2p2MyqsD6DPGoNTBK8B
QVaX1TgrppHi3fnnc3SgjSGlGztINDHpU74BKKZzsmu9TEEpUSBSrtFWuJum5FNK
PCmxner2F75IV1LpqhuqKCxzkfTR9sZ357qjB6WnAY3CTE5Lf283Jn4yqzdIb+yi
gCWP2cN+PJjtmA/xlJQvSkYvgi0cedev5o+FldAskVLx8u2FFFArkOerqiI384G4
jbcNh51IAbjLncBR/PTcpiGE9rLWzR8WOP9xlKUHdqRuZ8fFouQ38CdocIKyE1z8
vPQUFDuB2xb0yQZSMsCUALavu6/X1K6Zc/7tEoFE0siesWIs2gcJvYPDeFnkkhd1
yVHTmSubI+YBrqwxmjLjtxowlVoTiUq471DZ3TUWsiCnGvzvAfRWCWVKNzQoN4fJ
svfdrllb2lUIhFNmdvxxRrfjY+VYremrDJxJZhp2TACysgHN0xvUENPiRHMeNx5Y
Vfij4gHiN+paBbgP6Y8gy2Jl0IjFHCDjMS0bAkjvOBP1XhmJ200Ju2pu6KBIGt0c
AlLWlNapx0Yg9XEQgg4LvMfTPu1rdjG+qNCXd6O/Zk1lpaE26iL2JKEk7lTEC3JL
FXYa5HmwrhvHmZrsC39wQfR/Se2d37RG/cDt+P7MEMzTrF+eugBAxo7ZsL0SqzMq
XNGHhyftmrye6OCqIVBiP/TsyLlRHnP/65yivOReY1iTuACfUaaA9KDrQURtOsgn
WPVICi+JlYjO4MZZi4PYTNkAEde1xnsqxYpCW/CzxmcOJeKWfT+VdN0ZLhy+jOMu
eQ5pv7XNyAbYXToAOZjlCqOzhGgbXyN0xJPtaeU9g4rdoO69SEwXPYCpwj/2zGw6
ZR6OzNjFir9A9eQPe1v7agRIld+vhxak1bF6cFkThLFmA+wXtFWZHjG84A2gD671
b27WiOfeZHVTggx+/VgBvbBcXtcP5tHc4jsRY61207JY68QVJg1P+d51AB3w8Rsh
g0r4c+Po8xwjJ40RJfDuQ7Q+4TV6Y3dM0r4gqCiP4MrBuRe/6iKZbb7xFGMhYNsG
FD194kTgJ12CabXv3fcH0DTfZBeVSlc9v6dx+si4C1RWLFcQBHtU0/6SrrfVZcKZ
pZ6tS9+VIH9Ir6u0P1kPE4li6hflE0gwwzJpnNS0lUNwecSN3USd9oL3U66lZf3g
iRpLGPgJNwE0iY2ZkTkhdcndqmmmzb5sowVb+vBKn2vzYN2Cj1+SBNLQWFlpnrLq
HZXArGFibhQOGtpvRS5m5SIju7socn8ZeEojXHDQ092EHRQXt+JEApJG1CC3Dpg4
1CWSRZv1Rda1agG64ZiGrqsscUzD4gS0qXU+IERwaIs52Dt35Gm/kGAKgk9coTFr
ZOaVQtIRIpoYVU3GIrTRrVNJZv2tri8T19Ji3lehSvExbgq3oIeMEHAxj4QthRTB
kr1zCe7bAB2Liq//mIHRXUeoDqHXO7UginCJAyz0Tj3AknVzzgwAIcV9P//ifnsr
aYwchkY7aIATB9xfoWSMvQbB+yge2oMaLQ2D6Vwg+FW5yz9SgiweQSyArZycG58v
NhMU+LimOiYoRNeEGCXOL+XN//8TFROX2vZAGPAAbLebC+UF0fA/vnY6P3q24Obp
mcVxbQ6uib8TeadnL8XtmJ3wMFcJJlXDkbJd6XlvLMINiRAQ6QIJ/j3Cn6odwABe
XlNTaFG0J3C40tOHlG1RHoUEsKPaahO2sIxpPPgzJoQ03NMTW1340Nv0fb/wBrYh
WXYEv7X7VUMu2tn8/NXur/9jQIYUP03wFXivHBQoAG7l2803tQ36WTLAf7cfDf8+
U2GoDKwSRK8eXojmSmDL+dCjtWEhpjLNSdzahqiTjK/j7L/Yj+I6Rpm/I6HbHTdR
w0cZTuMU+LCsZC7y0N83mPL56OL7mAbUgwvEQzJ70Gs+KuNT3Y4ucLecaHiEAcHZ
WGNdohC2Gfa3QvDraA79FR74wq9d73j/2eiD0PfpoJJmQibVAgb1OiNyMFE2M5ZB
M/9cY0+t/zpNOr67IbGs/D3EBsIvBN1Pyhe8k1P/pWDKKSS+EhbT1hVdfVyg3XPd
7P8YuBdmzAULxGZ8eBtrETBC3UZLcqrWIy/NYtBeBwae1sGbmGIg4LhqPmPkptgI
BQOjJVyKhQ7N/ClDIBv/60vhR/gg5ZGor7dVHZNkP62ZiP1nxkPP8e1fetHImjII
nB6VulDxet0e1DEovFjqSw8FR9Tp6tN/q7TtwWEgMEIr8nHfGjs4c5emMdB18Ckp
An6U0YbG5vbepOdo+tRAfGX89ecbRa3YnOuvMcOzNxRbxUzlDzRsUyeaNaEtySxh
SaThhSLeZvaBKNXfijdxSDw8rj2Bfoe5Ya1Q42Z6vgXrhPMIO+Psve1WX3BUhTSD
cjn5F2h0+KjRaa8mnJnfzBBl9jIke0+LGOGMJl/EF/buG9qevfx4xOvKjD8uiRC6
qYCnqS7AMz/TgWv/uXpI4MltlMP/TF/n+Mw3IM8SBgahQCJdmrlxP8q4GSR0aqf4
245qFFEoik1IWm0fIoXnz8MaxjEb5JYO0fHJfG06KNo7t5CxBmOQjwybeufxBQYa
oQzBGMACR7AOZh1qaPwaCMkRP1O6R+nImuIsgVh0gy810AB5SFjv5uXS7NKyjmHF
TYZLOdyZ4R//0mOGeHfju5dxC0eraKaFsIaAJ+WF99zW+oi25MojSxBLoUsPfi1b
eLruU0jvU8/C7a6GXgTRHukjk2G+YYnxkim/8FKb/0+dSTdpeEsg+OXp1qA+yMPa
bycrJd5zxiqz+2G5Vsc85zACGZ9KoM7frEm5EBnkuRfeJCyarx7Y+tJ5rWnNa9Us
TaAJtn9PGVP0R9X5U5Z5AVQmVH/tYmEHfBzEhKWjxYdjH/em4zbZhr9ymnw5hdtC
I2Qrd1EYE3oEA6yS/YYL9EI3yvAijTzHUxssBT1TQ8TuIzPGnirgNwfJkedYg1DT
wdlmmK0IUctJXCAz6nXo2WjAdmu+VHz7/dQkOhyC26GAyBYLt7isIgBTC6px6ENm
b396yGgY9GuCFwIXAMEfaCASERWFcRldXukrKCg06QPh74ouDZNvzY+HoXIzw2JM
SP/AxcSdhtL+tTmmHg+2zkxSA+b1ad9pGHriyqfio1vY0wC8VyeZ02tcOn1NkT8w
XKu8CBR8aNwe7/fmMJ+YI3/1h8eyENoUGYuA6uhVnywZyxLrYtt0AocrJwPIMWir
XxxeQGTUSoTGav3nQaPpnGV32QlNKWvCPRaKBmnRcCDW+ayGoQbchA0NLVFb9eY2
EZheJZV2zHGeen1WFRjruzd/TErFKOK+tv6Tq3/GMAuE9VzAjCsw+1J3oKlR0lYu
3qf60i+qaLdXUI5eE88bAwu1zruVGgbpDU9DBR4BRcyOHqVoao8PAJ7AGBrn5SFU
uDCzNgVqLoUu865l9IIUD4AeUW0jTkLsoAcW/Wr1TfwzKIM73QZoZs9mFA2aT99i
ng+8g3FMdldHRFfJGEBDMDaN7vlRbG99s8fh5DRAd9+UOb93VLeFqkWo/4WKls2d
lDMiJVrhsn/qXpXL9EprN9RF0YploLYRA3s/8Cn3zNMh/qqCs6k132iIgSAR4brU
Y+cyyxORiZBxj1kGgacQeJRXy9RyNGc+aO7z/MkmUrHibRtiH9vlV2fmd3aoIrPm
BatDVp8jxHVu7MgSH7kK0YOiev3ZMZD/+uF2Uqc0zCXv2lq4RLZ1WQf6R1UT/j22
Vh6ktHDKd2+bgmrhglN5Ds6izFmuogl94PkJyjshlvsPbdCxa05kJE8pUxxEbfTe
22c30i3IStvLVGZ51ziwTQnIqALIKCeFeSXwagXc1CmR51erois7eC12dUIKKqHd
x2mmQgUH30zw1HO9Ao20SEeAlgQUOVkMH5+W7TAIjnSG+Chhrrb19fQcUcuHP5D3
REAftAoGA1YtGq0PFvV5CbbbLyKRGDn5OFlTFi3N/yksFPS9NsGe4Qd3J2gwCgkM
zdjh4DR+9XPWhQQo8jlVhhhnI4qWiXC8Svuw8yPYJg7kk65uhMBqrHijMQrDer1L
wbXi9rAsx6F87s10u+08CrDKgPxcaVhJrszogSDWE8OwVsW52CC/leY6XQTuYJYz
hbiGYCDu5/j4ALgxWGQT31ymrmndag6Zh0nwcjc3DT0yeiDB6amcQoX/Fk1P9z+G
/chFxeKgD9ocIh6pq+CTqvuGnyhzGoY5qQsMjIm6nu2wxGcJJAvNltyXPHEMP/kB
Wj/k9yHj516ffAU90ecDElXKVE/yFJ+q8VVgM+sCtqcQTulbvpmJ+YY9QgjYAkyH
xkpi27AUbQlTrx2WGdd58rT7ProwqXfvfwib0PpWy2rIKPQu+vMml2PbL0eeBLNV
WfFCzQBAb7Jkg1yQEutxFSX0zB+fHt2FMkUg6mP1u9WVt91aM8WjeMhURuBBoShj
F9pp0Mgc2oWLVTa00FvX2B3/gkGcrW3T6FhjDBF2nOHZjJjuEm4BTw62BdtCt6N0
zHycZx+tRGYUEKVHOj1MyXVj3166qq92LvxerKiY4/f5LKRDo/cjN8ccnedjFXYc
M82vc0Xz7EeXck5EOqiodcz11W+/3EBbV/y+FkZVKEcliFEb/N8w9HI3OFayORDX
gDdRn/m9ZFWe7mZLVEt56j6lfLQz4P9Lp6i/F0DyzbPTKizCKYumraRZSK63WiVX
8Pr61DA0G7f0baKFtOud+qdtlPrDhfloM6Gu4/chb3t2orYSR4fHD0ZjhLIKVFQC
MVMDJ4E2ouObYs5Bj/vFMxwJ4EnfSKy7+OpfIzzdKI4e0h0acDq9JE8QYGRpeBIX
T/5uMXI6LUbiw4R/n6DFcVdLaosTAV1s2TioD3KTN82PyvD6xHYrSnmr0wnUE53/
tyLrV6eYtnOFy26cjHS2TnKxlcnyi+aXZz/VTCjNSoo1B4m0WBBHDTsy5utTrKqr
y1PXaonNisx4XU1hyWe37Y9+4k6yuzedkBNnCDE9TugXFRgUUApZa+IbRFTvI4h8
VW/qzdZbsUd+zGfvRBY/1lxlC1en2jqjb8DsgcwDl+5mMs2nWITTvuH8ytQA+LMT
GX1iUQkIjEJoL2mdqscSDNX2BxpmDGzFM7Eo6nNeygoGrdju+m3kVNmiyNtTYk74
mf1IDBZnruAf7pUUkiNufF9APdT/Ml5LWtd7lXJFsTVxl6xcXAXxdOfy/j51bgtJ
bxB9j0fiCGhHn8MHHbIOfIGY4XrYgTBMYpo3tO48LC9Mkq02hZZorb3hLloNySm0
VQGJ4i9dlcNwpIiQ5UgwUj2uth44tKRqMcCp274U/nIvDueJxHoHf+HfXseTWNi3
5XYwuZeUpy+9JV04t67euQTL7AiaKvF0UAUY3iZ8T0/j2R1Z8hbgdlxgLeD1NDWV
w3j8IiXv7iEaxeacdOmbigMYC9H2BiG90CzzeRaP/SfMsfMhUYwhIACUhlal4ZeT
ccE62ddOZdvKaQmGoYZYDroCkJh1/Jj1AWfoCEOwQDSAtFU53f2rcrlXS4AuWREv
0CvQm7CsRqDnGbLy4r4dbIApM/mL9rBwSPmfpiuUNqBY96eeDOw6/TN6C7+XHHWv
EwHBjIkh7AZIDGV6yuP3BkyDVDXAQjT6aRpHIGvcjBNw0WMbbQ2qxWxmSmko0L9K
B9ovDtkuRbq0aPgyKuzE5m901LWSsHGFjwUy0FYvAKL7Kr+m2K3bdcvtvRFAXWQg
zLsPgxiqxdYWEPQ7h8Z442HtCnusezZPenRgWBHD4qTBMJxpfivB18k4V/GPbDtQ
+DHtYVtSL1R3CqVwRjXqxe6AOH3pLlkOHkGmsFpY/fjDX0FR90JV8SFcBJ/H+gn6
MiJ8cYUsE2O8EmOP0bGGkSEcF2y0ZtXySBp5vKnRJkhcyYqrVQxcAykPQGWMCls7
cbnG37g/IrG9cLvx6w4iKGVIgrirudlaycYHi0HzyMs8H9Z323baKaon5hnhwWD3
0mp6+kKC5VCDY7nOQotORYv14brSsL8uLSBwuwSGJcwbDp/q24MMqqEsjdnikWLk
GE/mftLigPDKgEF9e2id1VE/Md71rfi1h5Pjm7nrPiAuM1mBu2qc/yUKnI4N8GZR
2/M8ScGRyT8aLUHkxGIwkL6BVC6EcPmQeMl5wHN+bKNHraICuOb0iYC90ERKB6TG
A54hiG94dzOGq4OqJlO8NMq3Yo0TECmSpv7KLs9gy4RS82CBnEsY3NJGAGpKSuXX
511TZrtEB+Rnvn+jhQJMVYOknPLrPcCYrd1A0GX2EtLzMrvhT3Rck51OICjnlcKX
xk3PXXQvn3JRVSLHaXBZpLCbozpClduNGAM06APWy/aSF62w4QLpWiWYumcaM7i0
yRLkW7feq1PQhQBvdBpQIGHM72Blz10Bqa475yF+IDnyUNcUEILSCGDhkSj9d6Ve
SpQVKIfODUU6eccCKzuEgb6t1YxwUi9hnY7WV9e7Uc4Kw+zZkeLRG4xSrkW+t7Nz
SFsFXcNf0qnx/4Ncm8KtfHaI13TG26gGIScKm9N844Qk/S/LdLmoq2srfdoxj+6k
U837jAPMqiY06Q1DxklFUqZNtNbFPx3AJ3zZcIsy93y9j7D4RlyktLnkqSRDle17
Qaq1zglNzRe1Bc+UtjoNB9UPYfG+FgZYrWER2DNqFBMGEyDZKIcDgLt1NakJfp6y
1LedXGonUNUZtJwBGcWdEcCrQN1+t53x9UV7XOyFobcRz3Wyf/hvZjYM1cjpfKC/
+PnoB7XDiRupVnVlOu60nrXUth80BCualwIpKOljIqrKPQlA7eNcuYNT6umcuFco
9wCPbRmBxu4CKsPdLjScmW55vnnXveBdrO6EOdds+sumgr0j8nBeO+RYKB/dfwh0
0m9oNefJ8nqnCUTg3tUj2lhXdV5s/EK7NJTTfxBK3x6ueZMKSuN7FgcuxkjeNizo
nW10xXtb8zf/99ALbhprEghERc45Rj5pDZ0DHmboRHJW7oxVgE7GK1zNcYPKsCqN
GE3aocSuyG0BvIKmL0AGh4tMGLKrCcqmW79qx48uBwE+1LkS2lHMiythaGL5nqEa
C05D/lf3p3j1S6ETeHeOPAsd09H1kkmoUtScxPlcfFtcLgB5k1URC9aL1yEZ5c5q
NdKHRNH4DTEeLTTbqafyI+q9dgXgribc/pEokASiF0idrDCxCjTCRB1Sq8amQBHH
sUs6uTr/4WjLndStooar9M4RwIrSS17Af0PUEhQi1+Nv4IO4FPz84w/t8Rjq4FVM
0gXYdbPZd29lvfj2h19KAkMKhHzBvaCmUqMyhKVHLWaKKA6scNIUm3cltkgSBpfT
UA+TuPF8Z0SkVZ54mKcMs4cH8OdKGBKnUU0N6zaFujqDZfUxVD+l96XakWs+gwnJ
4pr/KfSO1ACnHXB8uwd2843gxYk9iafxcbNQcsL+qQdOcrAM7kIjcxc7cvNrXlca
FyZN4JpYorL7f5YnaYU7TBPb/tKAnQ4w7CqpJLPn253iW+XOLpP8MvHVyxkQYzOc
t0VLeoNo3qT6gxaBMaZdVkyqOthm0tXNCwDHAZ1JjM6z8JyPeszNiClJi3yrlzio
eWjp7QWMcdHiUjyIlDREmnnV/mhTXvBE6bQLjFi85yywlSp0SEvhsJzPxvZnOfjd
sgZ1OkuUjuSva4tZiNUZ8cIwAS4BmzoVPWyU5fx+xIuGA878ec0Ns5FtlpXaGQte
Vn5Vxl0ZB6qNEMJ0UEaq4nti9Eg1GTfK0IuvdDubqJ8d5chPWLz8jdBPJvFCIIdM
Qc0M1yNafovrUyStl0OucIQT7pzp+acsh/Lrhomg+eT/6Bij+bzi0V3DharOmxrU
YOGv8dT63QcMwjzHOkhdsimdn1929trZuskC3jHZak/1c1Y0F5TpfAst7+9PwC4p
jWaxZLruoxUY+BGasOWkyxNBLZ1y76YbyAxtEXo6InKPvlbBy9OSFlMmFn4N6QgP
m1GVkiBrPFffIBzokJAXjoMFyRxQmru1ML6rt1xEVgqISdMyfy8FkUanHyDQdNjH
YBRAceC9hGUSITRAnfUEWqJ08KVWsTCiQEI8KaI3lynD5iFY96tCYfEG2CVzfM1w
XITkRJbG21LLOO1g3ByceuE+/dlT8XC3NGk8UqckJyTSBHcX2eCWDkd9njmaFcl0
WMby5MblHoDLwoYgSJAp3eT5ao0mQP7TbwGAkReX1koWWsZ1GxcdiMK5USjkV9nA
DfQRiXGyE+C9mc2Ct/RbRsPaCV3PjLgdggIDkMdo3KcxZ5gUU8iqrLf35AdZuksf
nDyv9XRHkUU9ILnFCIrkW0CM5WU7cZ7S+nQXFdeSYkkckea0cwdq4qKdF1Jo3AAH
KdIqarprZn8U22prwcdbCxEIahSywY4qPU0N7iWYP70gNmctU5/G6XMu5IXnGViU
13xJmA5z/g1MIQAlfeFcfm3RqbTypungj9UxhoU+vQrptsvjoVJ/vGvXMrfcpgAj
Xa9VKKYvY+wPv+HV4jF3LHuyTdkrW6kcxMqOHm6eN+gplgIINafBBDbmuvNKkTBD
V4Te8PSvVFHfTFcMYdEp7opX/CINoZQIEG39KnvSUIm/meG5o8lmb725u27fAGBn
8u6ggEgW9DpYszGgc8eZ6UyalA83jSqmMVRBweVxO5A/UCBLEqc09MzDw/LP3jZy
WTNnPsRNAjVP3OuKYiwhJJIpFzOoARRJNih/gUmigD9RCTmbre033gP5EMNShIxl
SPxPs/rX92ksPCWTFm8EO0vQWdOzFZXxb4VfovuGU2U2s3OSAUyq42j1+WMjxgJL
zKHhloiN5c7wMotJaeT4dpQoOfIlz3K2Q6sPhOD6C/ROCwKvo9pOLMR9QQWBSJ29
eLVH8kIc1mVWE9acHO0nJJH2h/acneDRIzW+90Dbgz8xvnr6Pq1Of8ePNrarY7aZ
TTIH8pnlC9YcY4qg8Lqi/levoHKiyZABuvplr0o8t3TjzBLwTMVxEVwAwXeKTJNm
fNdPotVNtM4DGJ67Fc6i3I7XM19/6Q5+zzn/aCgRr7sMnj2HeoAecokmlV2XEVf4
9oqFBlekZnQB9oC/wTw8ztWKz/vt4xFwie3u4eYhssZnqA8Abzs36pxObkkgYNBL
Hz/HIX5zyRHtq98BQi3Rt7rtIAjRuympdXdMAhQHvXq47X8DbaGTmqlAn3HEkEbN
DfFbqkVU7WWTiq4xtnp5J3eHydvvMSPC93M0fRXjc2CeJwBnwFG4+E3bmZKY4WoT
AVbzoNKqhnJCFVqSUQPHzdq0ssePkJkfXw1H1snZ5oBO7eYQLtfbQbpAd2Px80EE
oJfbYuZq8Qu3v8XJQMQLJXyvIT9AJqtxtjzN05+vK+pMRrCKHNAfupJN57D553lt
f01YkVGb95AiEw5GzxcgB1dt6JV7dC064hh677SQf+ln2eogxKrF0MaR+oR7R4AS
o6gI8Hn2R8WRRWs/kGIt22JXWeL1E1kijjwUBJhLnjHqrBjamqWOsqIdLqjnC4bY
AqCIUnCfNHziRDZMcMxibH9G0IEe8KoM+jFotpFDajdPwh8qWpaysmOgSui+IUL2
55Ei18kIeT0wUu4EcLXJ1IhYRZMY4IVxdqSfpmY6oN2VJvjhvmRSE/A9gy3CKDPz
I/p6pHxSjtP1m2aP1HOsa4hZ7Q0VGjD64QdUcDTZovJEwgzPQ9T4O1IDe9kfNDVP
sYCfr3UkC4ZjatkTfHeVnOAMoif9ArcaY+n2iACf/zIjX/ALP7yrqURpm7oMegYq
SiNIikXqCdjOMrwKJX3F3+gh2pJQGDqfIwNsJWaxSiw7qNZ7IiFpfI4Eray/24zR
hlTIUKQCBcUw02ykntV+3yqH10WRhXMpxtxRtCId9sUTjMHIB5sIgUEYrblEgRM6
LdafTjxbYlbLPDPFva+2+fjIbKwN6ICo2e42w9IPaHARbnv9StWJPRJT1Nm7VdJc
P5Q0oHYbCJ8ikCjpYadGpaY0hirPWDkpBznlqT9GbtKHlXQm3DufLEHj6441EwPW
vEhoTKcm6M8KnYYuXyIU/JQXjW3oy6So+dMtpYAORhvqGOxZjoVCgs3h893ona+d
fwLj+LOD9gFonxCPNKBE39vnzxALffqobu6JnlqISpucKY+pryROvQ4nwHGdq5S3
IJICKjmPjXHjBth2Es5NT8KSgXWweZO2Xz/dQpY2YJaagLSh9n6rejWpDdwohlhh
rreyYVQqbRxtaWQwGxguTnJyQtKkbABFzegO5bXXy5X+jI3GBGJbh9VrE/RaMBlu
cEDJbNA6NjT1m5LrjS0I6SH/tVj7Byl7bbgLODiYeKpx2mJqZs4XTtbTfMDw/Z3j
Pv5Jaih8yx3n2wYKEw5eH4zVba52cDEujMlCS19gWagQQF45DNU9TBOThK5Guaap
rNi4hdGVSuWcc61qaevHR4QIAPEzC6exMfVJmgZX7togzKG61kvujtpAhVF2xmIb
rZjpFvvNzbhlgZDxsVIiJQn9MC5IDXecgvzRPcciF8O6UA2RKxh+rFX7WZhg/9Wf
ddIjQxg4cunTDzr03RBKC1Fo+dcy9ic9B0LaFbhB/AST+HT/kuRkBjDHjm7Dousf
k/Zid7qCb/9TC6KxYf3mey8a/mgX/XlHuziz8VZCNAHC6iVggqmCVHx6NxayY/XC
pHJfw4MlShFMp01je62NhY3b8o5XlDEtGJMDlZ6bvY5xnXKfoc3FHOsM4PWr+lY9
GXserJ2GyJHRY5yDgIZX6GID26en3Q3b8WVwQLL7fEUXpX+jtSEJZnR8fCGV5aQ2
4fEryACj22IYXcQzImwiAiVp0pTnSJhCE/X+2pp5vbG8yk4BellXzUhuWVjtIWXS
+QgoKNA4WEazKhScbulBbfue8sAOUSNp4DoC+N9M0N5X2G24suTN6lidNf4JRa5C
kz/NJeNbF8/nrSXIRJnNbM7MifTpnIxCNunmLwIFflV54zm6wkkKEdN6HldY1+3Q
+z2ULVF9LN0MORq2IP1CuqUSPkUTpJHPevHC2/9BTV8bq1wMni20HfUe8Cl/kzWy
QbCeQl1PDHE7zlyb/gWQ1dDGzge7DhnYO5lQHWm47zj3RLeZJM1ux4ywu7LN6/gi
vza2aTz1pU2eZcJDWrKmDClD486UEjST/9Xp1qKgWBXL4WcFcUV62C1h/fUdd/es
y53eVopbBFFuA4wLG5cYmE2EXB9KGJhTsE13Msv6i2cRdh6U1O6/Z0U1QTyDOTv6
JZ+HAH7w5hT0HwyeDD4q+ZIOO4az2bC9GCSAhbLfo8EACu4uI9ZBRNFzi53DmeDR
qYQrlyeH+LYGYrkD/kL/ucejlCokeMQ1G/lPnAbZayynyf1R6E8z7Mc7NtV1iTwL
FG9S7sVK1Ege/HTdDwD2LZNDa/IuI4Se7iEIWc4e/n+6NWfMhz9ftU8fVp00EoEF
6Vw/6psjtYTXOTxvFBtl+HPP79BmGw9t0lOffkMy5yt+27ZfrrbNg4CIdb0IvA8U
wlkRux6VDby8nTC2USQ6hDm5SgAl/ffCR/DHTuDG0jIi8KLzsKcecWa5Y2qcILs4
OU3wX4QZqe0J60gbs7aoeuK0aJS8WECcBvr2Ve4vIoRWfMHnrECHcu6T2d1g0Mj6
b4fXvUgtRYsSwKdS6C/XJQvrX6CYHhKkA9b1XmOK4B61vlZo7QMCLPBb/4CghmLK
uvESOdRnqA7N9ap8JAM2mjSeRucvMEo1T7MIKu04E3vYK8tVLHefWEq+3FKu8pPW
uKMHL9qMPL0tg/XJ/MnmIm4yybHAGxyvDuZkWjM3mCdcFuZSxJ8V05JRgw/g2K2X
IfRH8Zvj+rdHe2TIOhLNBRiGuprXftijkspzcVGgAAOm9ITl5Vq/Gz/oESCZTCr3
y/4F1oTl/Q7kCcVqpPz9T7R/n5+zuGvi40gKuvLtYfbqHiIK/tL9/bIUM+Pry5h5
KQiYuXfSOzMoCjKKozZLSymYawDDj7BsVGlssdRcivsv6qg0phbWoIf01eva696c
SejcLqAyocJqziY4Bf66PPEx4opAr7KTL6/G2lUtXauZtiku6EOApKrGkE/q+Q+8
Rq6Y2MMhUReL080P247Vlq9OVxh5k0tl1jmEHKyUE/e9Aye7CT6eSOo1JJawcF+f
09ygBKgbvNWLuEcY7cUEXAzIzK0W+QB1Mp5D6yXCxoaloaNRZo+e5ixWyqFhan+n
Soz4sYQ/0pl921ZKkzpaSnCq1QkFWgFpLm8bDlcp8JH2+e6kwxWa7bGfv6bKdR5o
qzMgs+HOguOfnIbl2dtpzsIrtJED7C2fBO+TC51kGSvFiv90jkKFQKnfzmFtcy3W
gfbohyCWv/GcG60qJS1uHsjU4OoJaKOxqAJ2lBZ9j5oK0MGDNO25kiA5lEG3rD8w
MA4LZC78lQ7pQQhcxyC8sriuZgFgvRbn1pXvYqXhIXh8J1vzOhfhA5ibth41O2DF
4h0NcDegPj+n6xpeDVWU6gBUsqcWfwUYFF3TYb52qN5FHxOWqnmFUDz3zxDXoVhr
Y/Zg8Gd4dHq819N3l0SVo7E9F9kbFdW6Qdy1s+hU02rQ7TMDOcXl313CqO+L2Sub
U/syPJn50lCKB/qwwFKirXhUDFX3iRbzR1L5aGRs7d/nroETTsVLbQGXSzClXlM0
pdgD4wkkNrXw1PJnLqZkcp9kR5XW5HwMglm1Gj9wdGfBChbzNc31WO/coPxwqoC6
aBZQcLzZrqqYmL/NNOnnk4oPAClZYXd95Z37+9Fby7CQqUiImlBsd52CQux+jm3B
Qyz8AopImh77/7kg0KA+GjjIR3oTcNkirlAbA9J+OvufD2fgMfhXi1N7kBJWcZZL
ijgQYF5WQ0HqgxU9AqOnX2tlD0nvJl60z8dyqN0wu4G7HMzh3dpjND8zHBMuSdUc
4tbSYCWX1FYLeI9bkPq60e+ldDNc5kogAlu/M/GE4zOGgGD0EtqE0wESA/JaRNil
8PM0rIoTzIErv9TmbcoYWXZEhTEkkLrzAyOqCmxgvg0RyoiMDbB2PxXoYU1NUkUk
6q749HlRC2bmr8OtT2i3J5YTB9rbtoVRjtdLQoqvh6yq1X9GP8PPTUM46BzXejEf
3l6rogs9+gplv6I4FKJc9jP4KTudz09C1L6bKu0sSnT0PQNYm4uLIyIvXH1Raz8r
gO2BNIo/3mS9KZfdtyFsW2+uJiYpVxD43YpP/TBDuedpEYJrKf+bY9gal+G0MSB3
BoHxQW2ThxgIGJ32xtyq57v4vfPJMlyFbMtF/w73ejrfDjflqfY7S4BaVlpV1lpw
2pe+VWJWyyfK3XtL2LHvuBD7PZGQvlNE9tyCeWw5THR0SZ2LZHQSVcuQT1Wa33Gf
m1o1EzcNTWPEmnxDBCVdgVVtsApf8XXl2u8XYTJhVTdXrmaHzlea8bB1dF0am7tB
mna1AKPT+Xwy+qnp56L6wzqaNqbf6AK4AZlK9p4hI23M2Gld0IJlYl8Je4B/C/d1
bmbxrPbKg8iO9RHi1oFRvrJia6gTeyNzv/C6HbHm3JHaniNtJzdnZP0CulhaHRkg
XLQ6HfMY/4eIXIKRb9ARRSkNlefJ25R57Fm86wSc4AtuAumrHHKmtLRi0cUJJOeW
Rdlb5NPjBE2oeJSOlXQNvEFVbA4c9vbS3pyuqOyp2iSs10nHs8kcDg+GHbaJYs8z
4XKjDFI5TlT8EPCEFM74eetcEMfCiqdK4o+0TYQUrQCGgDxehoF0+y0MZZMD1ETE
mu2eZPGjDGs1vBcuvBkTOGuquiTZJps1F6AqaR6dLsgFOeIIwizY2IQ/XtoM1Y1P
b83LIvR83IupTPq62C2lorbMEl9eI/cKX1mvb5RPcCOk4fpq7HPSk2I1FWZuHE2o
R44aKtSG2Y7VS1o1IXAG1il80HM9lcv9tfF2wpaPpYCZeZ5WhAK3rBzSJH1n41tD
Q+xAb/bBYe1e8Q13TzarC5nnp5YU9S8ndWihcf7WHKeClHPHpxpiCzEDnSBgafIj
xxKC82j1wOtUnac++FX55qXfVgLE5z+VHoHbmeGpZqgNMcoWj7io4v95WjZjDU7S
GsYG8O8PKMvT9i0Q8p6D73PALgtnx9HSlfyej4KdpRUDKmK/auuINkzmDynYw2jA
/sk9gnrDQtpAR2lNyVeyU1l0LOBPsB+r54ItBNV6g5I5B4qoNB94buux/uZGwivm
JhVXQWNAATH64Gz9zX/26fvuG0/V03hOkkLzHCHfDS9KtgWEZ/TPrSIenkIRPm3i
IIyaA5h7lRTNv3nEYK3W6Y4OjuES9ZYkbpREnVB58O1OW1jdfBG3NOk+A0KiXkpu
F3erd4g+lyKQIuiKFc152eojq0nM93JP2+61XOBmKpZtseF7LPDqTHrW8wodAQ9D
GAfWHoKoTaa/S0H8Lj4g/5f57mUq3ScB8HVnjI9upDH60PJXtFeulJJ2LvvBjR69
z9v+LLMHjfrCr9hUB7d9GYViA7FrF8e98Ui5MQa5bdurOpFuYllzMl8LP9JtHJ5e
z5QlxULF7BiGqSK25zDZUvJ6u6lR1ghX+IDXJPnrTAeq119AHLcofzcGRgeHHsNE
phfOlEWY3PKH/FSbtadhhQ6Gz2Cqgu3x7xgrdwEUN8oLrKOV9GQP/5msV6YpqXjP
uyj1/mc9FVnf0d0Q9ArsJX7SGF0zQbIO/7Vi4uU4c+rOMfzxrXjRGToaOQHlPWGU
LvR34E6HI859BMFkmZQRVXZJLnkUjjkr1BvTmDOALkIo6omXMzrkHwyrYl4TFUQ3
natmQeg8HPqkYmFtNJcA4UuYeWIj1GZoF8CuJoea/1xvDIMr03En4L+9Q1P0RjfQ
Ep4r5EfUwekWm/p/6nEpd3Vh7GcYKlbXCgnWnda8/sRE1OfuPsix3dHtaZVbVbl8
lEUMLsIGt2lunGtAZ2oOa6s2aWafQkAvPuKhgbwHLKNy9wjR9s1HxM+B50Zhjlst
KXsQTwKkRW8XfqX5Y7xPGHPEBxyjBMiitAZP6ZHomUnOTaD46eCAdBuqnpUIL3Jc
Zqxr9NG6ArVv7meJgSCV3GX7d5Poyf/r95yyE7Cl2Ya7/H4KGGF7izml6tEBduI4
b/is35QKp442YsclpqPmlCCPPDEzIRdBGzLhtQUBxlgh0pZZd/oM1lovmOz033LX
ixQ5O1EppFVLjmTVHK2d7yIZ4L8rjp3i+4EZdAJnhM8bBsZwVlYBDJCpJbg/3xuP
Sp7mHCFAuLLKg9Y/q9szWa15pTBwBmX01nXOXz3UkcrNqyTuZCHcCr55KiYsVVLT
K7X/qz9j2fB4mkyTG/uD8dd9ojRb9uqaV3DJeBKMa+9tvNRtq1HnOk4fPzBHY7uW
RjdYws/r4tg5h7etkQtmlXxgx81ORuvsmrNxc6AVI+N2O22iMFbJTdPUOmXXREz6
PajIzhnfk2qdBVj2+FICFDbr8KVPo1o3DtuGQaH5aNdggoM24uZX3yd1XX4+SeYI
yUbPU9T8s5s5sFc3lFlp6MkiphZSM4p1SzbrWfnENTI3ZwxrO6u85wriJajC1dTV
2/NXZLITwxzCQoiNPivf/SCW1TLIzkQ0EsjK4SyOz75yWUXrWWAxoky7wuQnqPPg
tYli9Ke/zBay9bW5eK+bVKopRgGPW9dO9FYFMQuHw/m6DB+gWHIKAaVynZFa+E/R
K4dyKmkWLMEiqQ6VdppXIhI87vlAWxNFqAFTHC/W4hB1SlK1nmGiwnXN97eOq4Gj
NL8rRXzeE5xgq3bVhEnvGgFX0n8YU8t/ZTFSLO+sdsHUCTQaX3u0/3ey0+j9pzmP
qBrmQacmAay/K0MAjvsTLNVixQEaN+sOIcnhr899n2my2pUlUzhWBfkOd7Ct5Zap
yaNaJbBEXS016oTs+Q6M3HD6tSyv8A2ghitPIU7NGIDwEryZG9js5O2oZymHgjLX
YHmSGhKUQmgaewmvyMjhrm7VazXnSVVxx705R1+ANph3piMrnO5QsQlJBuTXaWkU
S8T/oj2y5hXaTRRqLdSH587XhtIjqpN1EwChMFRMYOOaTfPaCfHhuFZLglmrAIUk
PlsBrsJ7/TFkc34uTp+cWyx0S0uprFyvQZY1WpEETCaXO6OLzynEhFtKqqytMX28
6uvkIKwHThtofn2NfkKoiWube2Xuru4D1IqvBfAQ6/YFKVRm/cRN8MezVny/GGgP
Ral8X+Zyo3/PF8OVrflTHxYkr6+wSsdGCVGBYPP4NuGYLV02rP0IvOrp+IGt9nBF
TVh8Dp8HrdcdtwueANOSakF/vAL9UIl4xglGyaKSdMz5gvsL0gx3XpUKsTCTeewH
0rGlYJRJ4+vh2fY+UvRXre0DnGXXEdA7zBcMn/w1wf2qvWjhUqDOWU0bLERb5Keq
dWwZTO6EOsWhI0iWyBqtAr/r+7+e1j/jgbI0dpMNLIcz+GmCYtC8d1GEnI5GUMek
JLBZhkdprCtr96H5MShg8wxMf1SHr9JfjYlcaeyr2NdqtLy0CRSB96elejWOs5ht
sRDGG05plH4LAT8VhtuMnDkSFNuorD3iOQD1fVoUcC1NE/jk1d4Bk1i8vHLp92Xo
Pqg0F1sKfzJq1+99JTukWgPVxYXmdDFNvlPLU59TVq+sVUKkJjwrNfBWfatBhN0y
saTc1naZhtkOLzB8Ox3E+sKhQUrW7csaxMnFobovXGv8+qLmk9T6KXQCKuV+vAEp
LJQqx4/s1UqmU52COgCldZsB3Z8vO8allMZUXFjYy7yK0gUnC+RgwiOEdGP8w/nk
4EI2+kXw2/i56EA6C6lHhFl+py94HD1aAyVYIKE790obvK0I2Y8TQ8ySRLcSJV+O
wKxdqJI7m3uw3P0PQYVczaXu4tfDAILECpQUJBeOfXHWZiOZPNhdNMz/lttT5JiI
eQghN0SJjtRr7rQYXTShChbUAwBRi28HeAZuqeTIRG973r5vIepOunSQtN6v+xHO
PMfwsxJJ1UxBk2L2zI0L19FpEDMAm5kts7GdLnv0RCP8MSeTZAk5wzoZIGThagML
eVFshGF6MeM7FzMuq1xJrSaZiBQURsBGq1YVnEv2wUBe/4gaRY1m7fDn1T27R30l
qMozG92jJQrgT8adseh1Z3Prtmd/Mrdkta1joShpZzobboKSqNwYhOilcqN/dR9N
BT/O7vDADIQX3G1H8r+lA4fQFSKsBhJdhkMO5h//NFWk5qtvvg3/Wfky4TW7BXqu
VgHl7l9dM01loB8yuf3Hb7ekFZmMW6O/bDpbUckTuvv4wXS2imRrC1V98A1n5yEs
ask/Y1upeeHR6uUBwddsYitJBXXCWlHEuqiaZxKVV3JviahvBtMULbdDY51VyOKk
Rh7XhRjr+NdUVYWfSN2KsKRQif04neLjpN7YNhbblLvp3ruvaB8Bs8w0hx6PsD1a
zvcsfPpJDcLJ8AKk44o2MmnwsoECFqxlGTxH48gNv8EzRdZjNGC4lJLZ6PoIau+J
geklKuI7rs9pTUorqZzrnj5OpqyuNx9R6vwn0HaGx5gvL9XG1sl7pWQcRQkLpSt/
JQ6cZlaYLJ9IubZtTX7KqrYe3lbaisUDnvbX0fZMJaoPNfpUIZqMIn8gTdbJd/5W
UJLHK/wVfeAfDMbKSumf53s0Ug+Dq0GrrQCjh3C+2o4cWdA06HU+VSVyWUqkyVVf
Ave92hRJ1D7RqGHgjFb3Dsehnjx82X7WUzrQgr7AyHrc5DLD1G9hZUNRKeDrHA5H
e+qwaibwaorO9LDIoTPIBkUI5j1TTxtNfzYvQCfuazhJotnKLIU3uShGCQqVH786
j8Bx6NI9A40l6sdDwfaFT3N1rGzNXNl/kKUxTnU2qCFcEbynf8LbQiwB9cuWg9a8
BYZ4c2go/t3g8pnNktbAQosddwZa4kLOX4RulrvXvmsXc3/JhXeVzqKZTtUjfrhY
l8xPMmIlgOavMltK6F4AHZqbLiSTw0rPjC3ycQ363NhNbGLTIs383kqEjJpJ+VhC
Tkogtim9Oe0fh+uZl5O3rN/matYOvMxPWY4r4OBesMvVvaM20Gj6ryQAkxbaNEsr
R2DPC7pUo1Aj+0/zL6QJV9lJRC+c5KHHkqaxBLjGTCRY4muEVD0BT0t+5z7kLfIA
JrsSC9KzSA6g3Lfpyd8rFggUGA/Q2mE1SjZAFxslbSDr9GbY6hHJ0zTiEejnJiPW
iElSaedoT1vYm9hV6OCPJF4BDqcXNFFszrCa5I2K4QieQELTvbFucSNIxde37qZv
rmu+LLle6sAZC3tpOKZdRYpsWxN1JkVdWQmaALIusuPs9Xp8Nqu3mdwfdr89byS5
mJinq1kRNdngPtGn5xvQcfweS8tFGZeAOFXQFp+lpGeLN51S9lT7o6euXQjo46At
vqYFFgWf1d/J0WRpMgAIAJRcPLT3olRCAKyt0tvS/bEtHGk/NaoWs/oHJMFAD6Zo
7EehKv7TSx81v/BJHNyCYTzF+pW35gNSp/XuP5SQCkdg5hbGLPOxgbWdR3FB+ZkP
tMUvZ90HFEWbuikJ+tMRb84zhLySSxCgmUqFo3wYZZXJEDnh1vqRVczZpqEbE6sp
XYPdseVStQ2H3L5BkDRn3k1jL8R0V1L3k3ZgaXLodj7xa+zNPWj9XU9R+E0cHYnu
A3VaZoV7cry93ZbRSbl1eG820cWJGxl7wfYg8bGY9H0BDhodqMSi8D77FQzIjyHu
YzQq2tE2g/4W+cDgz5HP+X8AXM5B9nn5gtqlPbagQ5ZG4jzyxvsCCCPpYVAnytOj
IEUDXV0CpQ16G1xb7URwxKy9nrPS3eYZUY4jDwPuMuseF9Bj/gLquWhOufvZFKbk
wYmc5vKeXCrkWF/ve15rj+AGwLQg/70Ejr8AowjbeGZNXr43uPrJ8tLCwiUrm2Ps
IYJ6n6SsQO5gkJ/x1JlcCi2iejgHrcjfMYvR3OsBfyyWkq0nUBuWSh2X3cjbFfmA
hruhE+XsOjoWCTJQ8+nscZA+wYBjBCFI3kLcawsgyk1Utm9coeEaW/pi4+l/SJIG
MkYEuIlenaW3PvIdp6xnnlatW0lAMo9VRPvMyJKIjMNDjWLmEkRduwTS+AYlYdrB
8xn1To9Dk3+4QqR/1MM3qwMjZC0T7yE74VOlLgFlgDzBBT3pAdmYIO6N0tQKQA/C
nhDf+jrqP/uQJbLG02YALR2fvTT7o6K0uGEPdSmy4UrrwH2KLM7ZUD18C/IkVy7Y
ZqSpNa0GtE6WeJBYuJPVbL/m7p3bmVTd/no653vlJQnAFLg5jhDCRlhqF3a8BPa2
CtV2KqmbWySpLEKlOdLaB+COMdtTwbRTRgV+uOt+qa9yZ8TRS5u9h21YBx8goEin
XTu+NpOGwm2nq4kYwT737REvN/fz6sYh1CZAWYn9QPUKfTrwRbpe201AGV14aV66
wtGAtlQrdCumSZS7IBDdnOCgI4fETciXGRmo/jbQ6p98CvtPLiXgrJ6cly+J9bBD
2PlvX9695pnJhr/N1169B7xKHYDLMsy4Ks8j+oLv08wmzWNZxY297o92U+mvlf+T
u8SfIIgHnRSBUghm9T33xM2TkDvvR8ZROJSydK/d3002YGdKz/NG8pu6n13rBaWp
wmUtep0K57GWSjHU2gdGPFiEElPX0kG/0aGWz4oMK3AQkEArQTlAu2+n98Exxw5c
o3rf8NVRFTp8fMNiGb13wE536OuOZBY5vWmZvSI1OfwF3dKBVeRL2aNHZRchGwpP
2Fu8FYhEUH/qPcFdyal1Ob6zRcDNJC41x5VKrMoni3lVXASRZxE+FxA9W/7DSdzh
WBunVQZDN3/459t+onAU27so5OtvLpRRP5GfthKsavNEHFvYovtucC8WeXh4x3e3
LBV/c9Bpdc+EHBa29c/r/I8Fj8TCAbn/EcVDpW4ksvl8qat6kqlBFxbnzt5d8nZV
a4l20uiB97vAe2yBeVMQ09dKp2KHVoYociacQMWsBcFXNKDKdTkiyJG3Q4Np6S1X
5hi4Jz/ev4KrkH7kGzBi28RfzM2xdIq5w31coHYw8PeuVBc6CxnlogC+aOHjl3J0
ty+ecnwITsBsnGQV/qbnlqji4NDP+FEJ5qSHPBJCez8XS6D/xfEQbVpaMFWA3pwB
Qi/V7wtIVUJPZc+vTr06UF3kp0fjsgduzOHqJwx8xGPvOkKIys59LEcwcPUMmX6q
Uf+3PeXknVNoogzPaWP1vBP8d4eY1gGvnXSy18r3u23cGfoJXr3FHdMevCeOrKIV
al/UF94mBp60MdkP4ZjyRxn6SU0C5bHP1J03cr89J0l+xAIs+EV4sFgQ8G/UdQKz
bWR6/fGOI6n2eVr8PDayLsjEcD3+3H1ZYJeZszAVdJ3c/vwkN8BEZevBUiW3r0td
5yqBkQSkP6k5tSB62NGv0DUP0kBxkimXIdOfNP7oZdrHUQ10cc2VyTVRoDvrgISp
BGCX+1zw5AZkcbWwydK42rhcia2Mu4r8r9K2kHkO+sAV+WTrViuSVNT87pNw+zGP
n3pXFwjEVyfNuRkl4epFd4y1u10GpM2rXf71kGYxi1EHqZxtVEREA8lJ5Gc9o3+/
ZP/V/Y/n5i4bZHtjzdAcolgXTSn2KDu4H/mJPf8kPbfmpsA8EVEytWEKa2XZuAlg
HFG9hUN4FyrOhv5C7YIRAlSPjtCkrJaU/esrs030uKcjD5uVJMaKUDaFD46JQH39
rJth+edZj9rZc7SwgQHdEM1V3XxAELenbZHV+pApx1Ymxq4JW2s/o+9exfFoUfSA
zLk94Kiq528ak4CWvUb2V0sB6s2SNaLDRH6RUTtAbynaCz8KtMpktxKo1C6igom9
OfxLiS8EfoMZJdAnG4T/gLGL8QaOTzowOosdy99jCoQaMPCFUWPB5zRvBpzjbSnn
uRG3zcHALUH7BXfwtgpKxjYr1rBpJuy9pQvqM7UXwynAPbskVGYNRU0Daomepe4y
GcT74qnWwa7LmvoXhoZgq2qw9yQTs4r4SqW/V4x0xCWLu9JJGuAP8hLSHgorTn3N
ugKp9J3OgT9rXxbqiMYQZyPo1zze/TwyHCPC4lRAwz84f4hxC8l85UpYFEEXebVp
LkGQxL3xvfnH3KR+ifCDipQaVsRMbaVV7JMHYFEpGgWKOXs4pA3RX7bmbaQVktWA
0jIi7NfLx+4iOMOiIkhjCgltgNzm7NTWex6wQVafcM7NK3pFFImmAVSF2ttMZLoq
R55HP7Q4wBvuiNirCWUIahdGLb3Se0hhlElOIyragBuyjDfWaR2UXPjvc0GTei+5
NtZQ9Kx58s4Ov3Zmmeo/Hon4Ha+nFX7tB7B/vAQto4NtlE1sAMIANdVXvgk6fWsR
FCr1uXOj0hA4hlvmcPS0DMWqMKC5m0lmRRpGibG9tuKGFtuE6Dxw+IK9CIsskn5J
X2e9ih0nb3SnR9ZSz9UQJTFmLfAtZ9TkTVdbM1V9SVFcroG4izj3nmFKlQTARASN
2u2JRVeCLl59F2C6HQVrHF2oDnp2uxKJoASS15A5hBC+r3Td6ao+CLkxJUb6Otvp
N3+gKrnYwXA2oVjilrnzGCkhzldnAxq+/bWDT7rIqMZuc00yAl1VUCA/KKbU6z9g
3tD6wqAmtN2BxCGqqx0hk6E6X/C9L5SrcahdTFIN8BkyVCfSpZSnDPvOkACuB2gy
TccvAvL0vhvJp3X6QjyxfREnIxYx5pPHQFH4U1qB8sdXeOIj9+BN+TAX27NQuMUz
RiSvX5mfJPfiy0mCkhgk7ifTmzqAMFPQKc181/rYGZ0ZRzltEa69OXXQEUBfPsNx
nyzQ6Zg61x8VnTeQ53ov8Xu8xOBzLOnaQTKCcsf+2S1nzwORedaDak8NJ8qR4Hj5
GL7H+UNOAzjlx+UT0hXE06uhrCTALwJoBCNaC7TV/AhxiFCGMTiM7fX7kh7dmRht
h0qQ+mIXDeSD1Lqx+Y7y2iknpwU6pR30P59ajN04YyvDGV7HTKHA6eIdO349cM5Z
KnNuwFYN1uwaS3Z6XYxMSvjp3EZjSTBtTAy6u3lZpxE/qMSQJQHo6TnOsIYQDNvO
4DvELkNmJeK0Ar8w1GvG7zHxavphRqH7yOqWtaOgPzcwotqlPAiEd940kVm1TABd
S4TkS31BIjbH9q6kp63DC1GNQXG0iOmV7QyIHRfZ7jexea00wdVkBnZAr9zCPt7t
Nij7OCxyunSRb6PMTCQbmArgePvKwN7O9Diw8iE6HkJQ3JkVg82DsTk8o1k5ATbO
5VSTEWfwXPMChby255E5bNvNzlOCFIkRZrGrm4xw0CD4XWM7pF4LiUCFxAJz/Y5f
M/1f3y4RCwxf10VcgewgtUwQ6NXH5NljoBZCG+AIm4U3b4sv2GNHB2zMNdW0qoNV
B2HuUdt5hz5B45Km9WLoMCnfp1lIBMtaZo8M4b+SXbU0Az9Hir1b2rQrvxUQ7m7a
SIcAMNMqAGOj5lSlz7FxS2iAFiSEuvUNaLoOhuVQo0nNxZeH7FpJCgxDJVmiJPbK
YX9lrENCdp5xiZoaJ6pyGyvF+EOKccC8bNssDmZaTtHvKbm5xqq2HxFz1Dk/Lbz3
VirGAGZiADlR6oblXo33FxnoyFckgSHUxlGe6wQE73kH5q1MXT+o6y3Bkzh2oZJ1
K832AzVlqrUDlAm+x4baW7NUqh6D2KuTJOpNB41smTCrCh9Dofa7oIlq7NAdVMPn
W69kEIuugoCUmbg+keSyTAns4vcuxa+Vmt814zU5lle+GHOIOpTMSYT2BkiYmuQG
H0BKhkZtmHBUsjWVlfkzLDlFYSwsASAOPezJ3jF19rBMKBt5hu2EBT5tlTu6L6fH
rUUeUAV0ht0kS4BJ5Lq2mZCvS61w+/LwF9/bFU8wu0FTkoeVBM078YTYsj3y4E5L
VhhzsrOTqoein8qDkMppP6IurfesK4yhQfC/DMogcd1FPtR+ucKkj9c6slE+8Oxo
wCOYXT2h5azEpi6F26t/IAggSi2iSYXx1DP70jIYdhcWdC8u2TYWZVo8gl8Lw/b5
P/ypHBxeycQ7SPg+efEzTWixK7vN04zEc3KszupY1uUb9NLyS99kP1yfiTzoEpm3
fNMrReptW5C4sSdaEGC20NIIC+iHmiLvzvbKt1hJIbn/yENCKZ+/cQCIp/bIop7+
AtRDk7ft3c0ZRhNBA4jko8cg7ieSPFayxZwsV4AqHoUgPicuHHZAKsyjwvC6cW14
3v2blAofBadhTWQcMQDSLzv4OVx1e6XuxtSWeJg+zHn7+FvC4jzJdMTNe2RtGODY
w54sR/ocwadXQI/PJbVVbSBa+r6TSSRuDlMcNtlFQSiZjqN4w1muS/bE+UZf93iK
6FpzpQL5PU9KHkuGn0zeB+MsAmD4HrIJhbMY2a0M+rExPoZLsu1uVvOQTd2oiusW
p3Kjtw1AtLu3dOMi19e67f+Jeu6oP6SzIDgwVrZQggPOaStB8F2IA+Ab5LOsai1D
DQpencZMN7XWMmlqrabrCF9l/QD4oUiMAvlrDsvm/jvpQVeJh7QBWhRY7LpWJBHX
W15L31lMCnct3WaEPHq7EHAm0NHKTIO2w85qeU5gYGA6J9cC0zewrM/SaBD1bNi9
3TJ5j3JBGCPV6w46yzETDGhCOr+gTIP5yLnQZJHdHOFhTFMOKH7I7fowggvdihb4
Yoja527xCvCNKOD1s/8bjSlX66DN+D7wRw8ma9IlnynjETc+TqG5w4kKuS1ZCWo8
NQMW88/SEyQfDqm62AOBqUdlVjzBoASTXs39DLzRk+ul7d2UGkO0xc2KpozhWnUc
fn9BdSUBHvLfM+ldHib/YHtxzu+Ggvh1bvay69tB3wLBB33OhYLdZ1lJdxH2yvoR
wfgLP3uRhTV7QzTW0EHzxVrT+A2P9k0G511TEpLvvIVTYVaWMNk/N2azh1hCKjaI
+WF9MNRuQqHF3f1mqHO9rnmcyvf6tfDUKxL4ShnZ3MF95J7WOSZUCtY3uaf5Wf2k
haOdF+1uZLggshrjF4H+WxHPQVPmVrg45fxI1OXpCgtuK4NSwQLqdSdKzRHZWmEh
+QaFf5PAlX/NSJeJws4EtnX2UlJ9hI4dpRaY6CX7c0HnTtxMg5erU9lkBU8at0L6
kbr81ntk7PRVEKwh1xdAw+zyWwzW+HFTu37itcFYVcY+HV2lMSE8dmFxMrHYFLcd
r4Fhl1LGDyUqM+SzFNdGUpae5KndSlKAXGcNixa/xH4M3hazQn1C5YbyqVGjSuO7
H03aAn9B7r3ogDLldNMUtHRAasPz4/5XBeyK88fINAgtQl/2tSuBPMeEAKDr2aD6
SU7Hp2DDsvHpt53rWvAmtLdmw5oRoaeUEfSN9xIEjPYmXfNXbvG8nWTFsXnKMR1q
HbqK5YuOyUVW3XaNE5Zjc9Yf0To+ZstdrWjN65FWtoBnFu8k97fvif60Jh8w1rCd
SBjwtqibdm+NlRZx/UsKpUfEmDOehQXdPZRpO/PmqUjwjJO6oX2YDnlJtUbMUaaE
lWOiIBl3PFDn/MIpjGBMUA/xEqyoi7N/yQP/8YJsd/R31i+8qKnhYiVY/LjZkaKx
plH9HCWDouDnsSjPMuX1w+tyUaEdsHQJcATpF3h6V92IBtDDOYkWRZkevp9j9wXM
vsA0iMFJzm7f4mGh1F5h355Tr9AH9uJHdbG6GGN4CG7W9Cxydq+gF/K1QMW7ChTl
UCqHFHBEGhIajC4l9qg8ROAHOTrNW1WkP9IjvK4E+PcGH7Flq4nWd4vEkkEQKIcY
0WCun9P4tWs627jlpATgNofwOQ37yv8bb179BRkckou7T85Wds1W0aNHzs5ZnUMF
t0UCljWFfY3Ux/bMwLshP7jH3YMlGk/mJI9cP2lRSl6Q4t1NeDTwUxB20M1lzNkl
cUnEIev0YLJcJ233xtxWfh6vWqfgH6b21rSfHpP6wtRjxzjpNmPjg3qk46CXFySp
mKXKo2L67ejsnu2R8u5GpI07qmbQhZeWm+LXQJ3ZUYgbpr3VC725Ow9EIwt4C3Xj
vHBFz5M0sBMi3JU5LZcUM5zJywUIbh+ThlkqoZvJfZ6Zr5g6GDW3sShWk3ngrOlW
Aczsxu7Wmzhz21Az9GzDx/HUXuk8hof4sesODmcOFn9RGTmsmh50N1vwPGq4z/GO
lTXoq+wok8fIfRmN1pJBTlrOM+yWQ7noBl9+EH0pr1AG0+6Bx7HElTPZhDPgDO+P
O+pMwQyi9qZlzhDYV8/R0s5J0lGLivKJyrozVf+sgoDLPICYRchDw7zRHZrs6vZy
FsUixSCDFKQ0ceEEvEyKrOslZu5PiWMjsGTAVFldZfiY74AZJMCAoIM7uHr/imBw
4LMPaKcFeXozzWzD1xj0tfywrvELye55Y62PY0BXXqVUqs71mELWDdMmAJ/mwrAk
MBCtOwfFJxwBg4EXwVqAi0j+ZSZRNEGUSU+Hgj8oveIBXV+HywhoW5jyWVprweJd
Ih4JBhdX6mRFnx+nwIHItmceuyzhjR0GAnEFS5T5IV7CawjVlV/yakIF7DbxJURI
sjfu2AUvkfzXKICdLLhdmno9VnhUZ55LaqePueJdzbCMraPnLd3upqc6AGEybEVy
kkwzehIGbSLx4Eqin2Uz9Nu6yXOQx98pFWWXVYljxQllb3qSqifda5q2nXuLrCDm
kKV6w4JDMqmKKgqCT4FHHUeuY/1UT0OWpACtnxaDESXi3t5nbun+092Tlq6MVo4S
DftRoEm6MBzcDpvN+UYHVm/o4zoerP5FvDpdr59TCGpxM7/WbcuTdstvlCJPfUtT
Tfg9j9zGnqpw/KYQC4OWdMaSW1+Hx2m4vqr3iPjCbzC/OZfxMBC5TDO9m7xTKBz1
+O6gnoOBVMJ5zGdGXPJ+rzmTyaswz/rQpuqgwK1Xe6bUCHYNK4hZuoz2ee+3tdGc
Pow/JpIe0mzvoxv7oNX91av+wqOGsXLAOY+8MMrb4l3JQLOzO3e3v29US5oNy1Ax
aHlZ6t3CD8H1437xba7j6BTCZpFo2oWLA1zbZjimOSJwsh9aWrw/XMdHSQtimkC3
crArv3UXizHNHWhp8Gv1KIgvjF7VXFQD9Kdp78DgDiNShLN7FoBJtYj+13GKZUi2
FAJLvfz88zDnGD0Qbsjlb/K/KTbERnM+FYJz0CQVT5qW/dbeiG9Hby8Tyr3IWXun
dpEM7+zDD4lJsgXD71eii1uJVti1waVlVHr2AEvDFOzep7Y3aV6//I6RAdc5jph9
vmUfXapxGCECv+lz2638BGMOoSe7/FtOOILl39cSvy9Ty8ZirEdHTYua+JiXF1Xw
TDlj+b//ad7oYbvJlVVPFTR0jN3wugrnMqJxVugtZO5vYJCVqu/+nbwSafYnVWgh
/65ut+YUfmOqrxQKCYBnEnco8WwUQ0Hcftgak5K5SZ15yZTAPELtElHkUpe9qEsd
/oxz/rsBjn0a8ufLGt8J6clF4l4mK/O22fc/6ZC7HGCF5jw7c2zo44WTodcnzm7r
VeCLt02FAa0jkGoRTv6J+RA+E++0o65DyORDTrEep4l/0qDKOjes5aKqFhdpdSKY
pCueoXG5e2c1LZ7yYgqExReQx7no1VJWnUZfev/9Xz+T7LWyq+wmsODpQRSRRfri
O27DsnKLBZbpymmGbJTzj4VeEY9Ehd/3MwiQFwHEQ0wClBT9MynsMcNQU0pA1eL4
PGT+sgKX9vvyxRJ6y7F5mOfNmY6Qi1X8oYxbHQ0zRPmHrNq3Qoq1ycnHrP2xJdcO
5R+ky33wa+/ZYKvnUXRF7dGKM/HeLHMgnb3cGjHWV3fkG9Wxc3vEmwdlMepKGrVg
xxKWhEWYST9jhgfWCHSI0HMKcsgfmtWM9NdzBwtzc1HqJ+VUyY0nxMamokiFO08H
AHsKbV+peXdgsCBXuIg+J6KbSkcvNk8CKrQRANgE3nSrwZE+9ONIZIxS6xOCwGcN
yUfbbGjXKlpJFMK70NX3nhrjPjV3arneLRNOOXiE+rgSlvQ4Z1N4s/KPkfATjZUE
hw3zmDVD7mP0DOISP2HWwaRybCxLg0wwT8lsJ3ftqleyqxPuLOvg1hJqn1yz7F1d
zKrMqA6y9XUxk+g5PijeBpwWxDFvg61AZge6x2k5kF7A5DXbBYIkXIAa7M3SB/PK
HBosmltA3FQbmHlDHGZYO5jyRKtVML3hV1k2LMIU6is/DAANy4fpy0blsyWE8hDQ
YIZnk0BmMktgdeu4iCPtyb3BKFFqI9OySGMaiyGKZiwNUrlZ76TCqOuSjEsy+IKD
jddH1szOF3P//WQM6Es+PFi/tW49MQ0OlkPgKbYyx9sp+PpacP4v9sEzBLbhEJhJ
Jds8mybwHXhgRbhA56NLP7qY9pHkmEbs2o8vHNCha1g7mjsZej2HmPX0/9Fcj9HG
OHbwdsRJyARDCbkKDqbUvjEHaYZvPJOQq6ODpDyYmV99AR5PSP/p9dcUH/Wr5DmB
6a143eIONe9kINgnpz4MXijV98RMIVnRyvZjuVmU1++u07NUsSqC2ozM5yTCqceH
O8gBbKNN0hXsI/ozP7EUpe5mm2ZwYzBXAk4OH8fEl8R2pvrS92GEC+gS6CfqkG8w
5VGe9jrMOodciM/+MyFN+e0X/d2otwJVXDEIJDVu33cabD7dURUDDRIBa7U/FRNp
BFtmabVIPJo7ouxzMwRlIonkDXqAhwhyMSMMoUorM6trVT25azTHQQfgQJHLa89l
f1ZND/NDF5mYj3qkfRQsIHBQUyEyBcDovc6f987LzYsAGYoIgRfPgmZjj9h9hDH4
FQwbI47V8NhhoJJmKqD88NXBW7Z/CaIrWZgQoPDTqWsUyYPmVcBr1VXeK0DJAOSj
X4Ye4PyGZEOtvsjfYnRTD/xmo3H0KpaZnjrq/46FqkoqazuaBFHhvenl/E+hRoWY
I8FbgoAA1Ts/0HTa9UdeKd2VdjL/axE+/izOUZOALN9mPNm1xtyQ0Fvb/XS5NPmR
SeN1RJGNqtScVD7/be2xHrLqRT/kYZc9BwmQTmCgFfKthkjoB0ErllLOol3MXmzI
80/s8MW4KsZk9XUhN6jz+89swpZjKSZU8v9a9zGebUMPS8dguaBoAZxcpCGjNLT1
ddaEdcSU/saRlFgHy4eubpEfh0AdpxcqEj5XuiCEo396s2OxKA1PP60MqCO1K4OD
eZ1GjIUI2FZ07t8m11D8+VyW7xhKQrhe7uB7w2vF65FWVrXK2pTIV5P9WvYrlCJn
wPF7GqVW1v+nPXCdi0tnxV2zrV+Tnin1z+m0Yos/FhuZwh5moqzVd1kdi/iiUmDr
X86aiH75/4h3qD4P0W4rgVSFnmBtVSvms4h5FpvTuL4Uj8YDZ2z6MY6uwxC4BYwt
UffID2CRbw81WtyJHaW4oEKVruDQLZijJL7k/DDZYCkeBA+mhFQJwpItInHNhEh5
MEneN8s7MvRKmqfezCqYo/xQybMVb6OJo07XPwuJdJG52Hu2udwwLcJ5y3hupgDp
KvR3GmV0qS7WBf/R/ot2A/iQAs4MsZdeUyxRJ8mf8vaY64Wjtk7OWkYbS+yONe5Y
9+ksAanYlmQk0bFUVvNkfmENAT/iz+MIsZhZO/pJ2d4VKMJD0FVmJqEjlicmT5bR
jW5RKzqN17TxCHZEndnvU67baaQZb5OCH3Nvi6fCk1y3c4aGlAoEostEIm+96zDa
Gwa2uNvltjJAZIuku3xdfedQz+w5RafUY6jj8xcne+NMjcPocQNa7JhoGAeku/WQ
0S1mw3dqzlH8yuzogSkWBf4AEbAUX3QurzKEJiEyhEeJ/+KxNMVhBWf+FZyxYOPA
M7Wyq336AuN5/UPu01YPLjYoMLFRMcN5ar+5htG8degDRAQy2guUGATmu5XCoftG
P5P+nO8qlO8a80/0JfJY8gQoIV4YXbF8sPMQIIbBJScmHyqe7x9XP6n0y9LhMyPa
oz+uXUT3ThfmYNIyQCmWJo+WK3fdzdoFuE7sKTPzFHC8JFdIhPxhGcBtipoHED7v
0UXvXsxOBSilxYSPj0W5HysnfJRkdY9hpAQLB5XHSouUcdeI71cxVTAsskpAX7u9
gydKvl27HQ9VnJKjq+O0keIeobdWCBcdsmy5p8SqqQwYju20BWUWdgbqcIA2WDjc
SD8pv4huv9/gAESIoRlIuQyyrgWvzphoX4Wd2n1vgrVz1Ymm17IXRuqORid9RvNe
vfAF9wWS5ipMK7cpuUE3Xz0Q0fheLChGykUPwMGb9Gmq3he9Xz5Oz8v7kFbdB/3j
ZEXkYY1jIfwPGIljV+1Xv1TIjBDPKSU/YfXB6FnMSWFl+DEP/a62hR6tcVh+QDUD
V6nokRPF5daqqwODeyFT+GX6o1ezHyabb0IW2bL1E8x0Q7RuZ1yusfe2gL8LZO0C
9yIVK4U6Zy/ukA/AM9i4FOcsmU4PojvavGeYmscQuWjEk7ObhwfbsaWVnDc75tjC
CH7R7q5SqkQsVF6/D+MCb1o7kK2RP2aTZPwWbocsutw+3CEYjwt7swM2fjsMv5dv
RAS5unkYRokmKPE25PkKu+M9ggdxQhB5M7rAr1s3VYiBoAO6sYzwQP7s/I2a54vG
imIm50nTR8CbokwnDsqX+itdYeKkQ6ZHScFVBpUtHU+FcAiMDnlKVsF8cGloEU+9
utNUhs4E2fw7RUoIbxFe6SvJmnrdKww+Jwiw32VydQEt2swy3j9u7YmfLyg4/8/m
NaOdvc8tbfo+ClRF5GVORxkDO4cjiuHi6jk++VVJHXoRlM3xbOUPjPkcSOtRdDyn
nYFzDDUda6etE3YIqdhv2Mn/QXU9ZZ6rvaTQHBgfiKbcAuuZd4KpghQM1lJDjavY
CsaQ9meeFkqEVIgCZcQVsdvyPK0ME7dQgCR28zD19wMx+bNcYruLQfvMBcmLOEXK
J6lL/PHZVIjtSUyf7RMpm8X8+6tDtiKOV1LeQ/nJ8i2y73VKRGEl3gJWMIlj6b/+
PdssHpy+C6pfQue7QjyONEKV0tRUooQtvy2h/rJEUD2QGcJJ+wxoewlG95JreLS8
xmSkl/ZzJ1OojXhck05dCvtQHGr6QdTPRKEDmWrSejcRxuI4X4p9aON19D+W5zVA
g9e0WJribkB0uKU8RRNc6fZjpSgU3JxGMFjKTDJ9XHEMRtt7fhymFN4V6NmSLaNN
xU66e3X6XWyTBuendSXQGXBmdP3iFECCeXohO64A7gPFOlcVtxlyHzNSo+jSQ/uC
A/ne1UOryNcHMZynvAaMhDPn0gtW2tNONJ3zgy/wkxB1cR0RJttXsIsVExLgbaC/
ENj9W1X/ztaFjNO/6radmlfxrB1lufZfIcKgqvYYtHzL+Orf76QWwjHrHludyZwm
PRM/4fVDXpKk48cVaiVuKSCqoWU6CZva7yDi0VvougSan6LRccVo6KtlVxGuL7ko
WzEvLQTh4mfJQJaFuP7P/0T+yhuW+hc9SBNBhB9+6GePzctdOdiYE+CKfsgd5xvz
pfdVzm4ll3IR89x7Y7SemMWlQwMqReFknBMQ8ky1PEAHARo3lbuisgHGi3/7M5WN
HbH7HBLMyGRb/otSsgh8tF9Fh3+DbwdQfGJmS9yax9Mkfhj7zeU8XklNlHxx8/Qo
hB6ejtAhY5j94tPBKseKdVTVBop/DTgQbgXxrM1NNMrKOGn6xTzHCmmnVb567s7p
JFrfcR3hV6g/Qm229tYJVH/V4eP21gw6ah6VHkmJnJl26L9Axm3nkeBewa8L7i4C
RsdG0NbrA/GaLFBmvphr6u0eNQwiQ0BVWDFW1p1OX2SLO29+qUOxnAyjjcXykTFE
dhMDrGC8dqtVyq1eBu9MO8vk777/UDELptga8K1vE7lkleyNS/0gsO4pKeOmwBEu
vCKNNQhMPPORyMH9jWi3AJWQ9eb52lIpWysURE0/H2GmLu9jHUVt5weeuWc09WlW
RW+gQ777XqqkHVG5308+Zc68Hf2d6vb1Nz3xf4IwaYU35T51m6jgbIBn0nsUd96G
cmL06JtffdaiVBNLI/iIMypKw8+6n+dJI40Eh8fx074F2CwL+6PSovZ9UN8XRWqW
OYLlLTY3jluHh3nCJ+pBVvildEtX3VSWkSgMUzV2Y8h/Mws3VF7ImuYuw41RosIR
RWlonGm9qsNklRfVGoVf+icy49V6BBv0YA6ogcCwbL7zHHeaFtZ8Sz81rnwUV6rk
bIGkjRgZIBMVOTlsFP7SXUvxMm0LyY4i54UjqfdRiSD3YcNjR4S+kTYBQ1xgJRcs
eyHrK+9vxvYMNOI4CaUJOsfBRnRb+NT2aUoI7N/jW6ieIDMYQX3Ruiwu3hhsmmF0
c8gN17fcLBbUGnzViTxD7UUZ8fnapcUTM72PiTbcBWleeeV/QJX+ddFnRM4slQdu
3I0P/6fexlbBzs7tgfweR46I36nZZsNNJ5aSXssOBc3+Igruwhew89pFOCiElfiv
ykdFVj1fR2LJgvyOx6U80gGQa7S63G8KrOJc2mdSdsmFFE5Y4CYprGNSTfMoBlro
NTXCp4qPHjVzx0Py/jDIcbNfn1ziDadeEHMENWQsdZnGZzyShpF9+cahRmpH3MG1
ZzuhKw6JxdRDbIMx9y6Wi7wahjfWMI6t24K4r0aUYLWgfex28lp2ilgTQd+HstJH
LH60491JeIFXZJ+1QkGvjKDLWBPg9WIenmIzedSCrG2UyIwS9UlkzPDofcN/B3J/
i68f/bwhZ0NU5qN+3TPn+/jvRxfT4h14hhDaFWyFDCeaqCAvqk2U68mmm1pZpZT1
m7ei1pyj/sQLcMNkf58uafweRSOuSK5N1LyGqjVU2xEmgkrhJojps61AvBodYQXH
Jfd0O3dwQOiNZeFSoCk1PbgVfupxkuNUjnwF2EQJWygmQQFGco8ZdB6DOdAmidrk
/S+oPLwxNHrHGbEntdNIlo9RzUI5/WKDmZrkSM7ks0c1z5pvfHzoClIBeHYnwkmo
OuTyUICLG2IMns9RdTw1nKVUo9D3zT1YWUilmkVrDcK+DQW4st7qoG+LMUMIgxAv
jbmyhBidTPhN+jd2uiqWI+hB4JfylGGxV1tUJAmDc/cEVbWpA4mdSX974WVrYE54
0iQBlb2RPiLC8is0HehjDK5lC4th6rzfprHh/nOZyDPpMejrGWng164CXHiBhYXa
4VM376SkvMSZHUg2aZetvSFMLw70KTC33HofJDU1KT20gAGsd87einNVBH8CNCxE
1Zd+PcsS4hK0g39vW94NHxM9Y5taJmk9nych7FjXuq/S/gL9O92K87KutIiZegkb
eFLPokXVG0MrBRm3JQ+q0TlzucxcmCRu0Vt9X2xrKly5Ql2ZoLSGt8iv5UIeG66Y
4NK0FoE9fbK3KPBKj1dUFfBwjfOW3LHNvKyZW+/84tlGji4lO6VSdFaFFAVZTSF3
LpzzPPgc2Q6uVPW/d+rlZmp+kYxioiHlGPwHJ/btaLUJH+tgNjxk7eDsNPFHLW3/
ORXvmrsk/7jgyh40hApk/0irFFPDZG4Jm05x0AU4Tq0TChtAD60cVdgZHxSlG5Q3
VDAkhhpWhTq/Hr6MKmy4moy5uBK/wFufLR2OYkE+683VNupvZ3kkiwuhIERct9mZ
4mkr9phU+vn8gJmMnsW1c6sBwiWqChtFJeF52flX1lw3NNxHRETTd9N4k6YH7I3N
vsITlXnvqZZSqvg5ZeFFypG9eK658om5jpWFwKDEpNBQcLxAirx0KHH7S3vejEna
UB/FWqjQGRV2o5EjefubVqVuv2Sjv3n0oCA2wkilMBeDIwHlOUbptu3UFdOKVMRE
Wff4ZrFSxZlcReAtJ2vghc/VaLiexs37CRGS18lM2CfaBZANlYlL8xxEMJu2K0YH
unm7uOypZ3Iqkwb0EWXz6irzSTtZRCRc2Vi9CvgCOr/Txwn8KYWWQkGjQm6HqOT9
hGxif7cDC9JRGbC2lrGPULDoIURsddvP9aumLWn2+CYVZGSRQGY1+8/CLL6I+I7M
T96WJPk6au3sgDcIKV6K8Cftx1keWthjeCPU7JnNFpOgsQ5/Sa9iPxs8xLXb8wpj
bClg/t/jd/afyJdu1sLEynUx4ZJoihm5V8dOV7T07j0RwfpLLbNIoUGy99Xu8cH6
dP9K9US1vEs6256aTKYQW3S5RlxMGIha7S0GKgMHzv82pMAUi5KfTyKP+JI7g3lx
mDK8dFOEPI9glaH62BtkC0kQljLg4u12GsDRsU0nNW8b3pWzc4OiZh5s3ICVmqRc
+lkkYZcCTbcwsqZEbgfnNK4Udey0STPXGEyxHLRxembtACcAimq3uZgkRrLjXvWO
9OhsNC2xgezbbbCjYsdlS/BN+C4aZKcM+UqMp4i1wGPao/f/S+NnKFRbrnBGL5fa
feSxfHRvEJI2/4WcYKx6ncdUXh4raFtbRJ9TfbMnniGQJryJDCfFnk3kaTJI9vjB
FLC04WCOj8jIbmaowoQPDv+d/yrkTKoiD1MKI+PfgjYGm4SsGeQpHOIU0UQcpTLZ
cCyKpQW84kJyqFdI23cb/yMEAFr9kexZrZAYar5Go5iuC3qX1oMMQq07firiYjh8
W6aSpjarK7GrbJOCuV76JEoKY2hD7ufc0flpcZHan2NwRR8qCf+2PyEWp3vBUgem
sbLqzkQdqwE/RN87aKA8GJuks9vkHUae4NE7QjRD/X3LPzr4n+HmkJUNNZAFhxlQ
DDjzLeHcCBujA7FDVcpwJs4hO474AhTj6H6MDrTO1SVyAAsN0oxYTu6t4Oo3HfrU
lvzcYvJvSPIhc2XbTHhwkcSQuw/dAyZRcSqJj8dwqrtHeQIO54D1PkPptbmqEpfj
bc6zpXVF5C5qlNqZXyk1tT+U/KG+B+tBkBqdExfYHXEGKJy0+GUtOdojhdVDFbLv
nEOw4ajJP6qgAksn9wzl72l5J61fjPf50RBDO1QfQ/2xHsWuZ7lrwZxC6o8GCU16
1vnk8t0WnfsTQ3u9QPtmsx70+45qa7qju3/+s6zLrmxRJ5FDe167hfRSP4re4Pff
UxT6pbSIIJityIZS9v2OoiJt5qmdrF/lVM3tU71toDv6Rpkm7jFqvcA1qB4sv5Ce
bqrU7jol852EacSfOBJapo6Em7uWtnoAs4UBqegHhAwrahhL/yqgl4L2wNiUPYNn
XmTgBOuWOdo5oduw3GnxeAi9AsZFrjtuUInpr9IpL/9/EJ3vMOi4X3WM/fX91XXI
i60dL2tb2xpOxfzqi4aBtEv9LLRtIjnpKhSAj45OPxpSRbyxDuP3+1DGASFkrIVS
t5tMPlnRAa3CRPFwVWTe/XVPsvytTqDdecteXUyY7vXFlfR8+kJor11oXEJqvfCZ
7FPnVl3ct7Tt77mNmUm74CgXKR1SjnQjBDLNH57s/Amr2aHJii5/iRbUfsq02kaY
Z6rWTqZJ8qYdksRtXjQrj3uXnudXkJPtMoKJI5dU9dkKmazNS2gwqdI0lJnuYkLU
wofINu4mVv3FNU7xbjewkR4vpqMkOUSCRt/lgcqqaPlzFExh9CKBUv9qnPH7M38T
CXKPmc4W7GqfbAOH09kjwH6wxPlbUens49CB+Ez5J17b74iOXckXQih+AEiRBI5q
9lnIDVrGh/SriHBpf9fdq8JmiOU0TUU3Q5PJKv/5K/AulCy9V8COYCmwpVQSwZyC
Wv3lHQoy1eZF9RZp5Uwb6V24ItivJgn3B7xzXx213ISWjf7uqW9IUi65hEAgyKTV
4oDk1GcuNtORHuT9g7KZetoEJ4fprmEz8d4TrqIH/TVcWuma1tMo66025KMWucHo
0s15XYtLgqTtxYDkpjuOTcWt0d+xfMmxsmQT9N8k6gTOfNqZoqfi0phqMuWnefzc
HBvqlcUsiNWdVZDt/9z6+g3N7nQ6SBEhUEA9CVCf3M0f3sfApoXmJKJ3eGoN+zXO
R6uO011YD48nQvPpb1mAsShXCx8GUhoi2kwac2QHyaaLCalMZvGAiAbu7ZIzy8Pt
Eq/cjhnpWz1MmpxjK41QNPiuCvtGxVYmho87HROARCEWEsVGpdhjAzpzNXzx/uri
QZyIUgreDI3w1RiIz9pmJkpZvIHVgaR1HKRTWvgcqFia2uRoL0TW215tihdypaBN
6ABEIuvGkAWWtpw8Rm5ep8k6xaF5mj+duqeq6pFZnbYqKhdDBFkU7Ea7BAk3+TE8
q4nb5KzGf3WcBYfVU8Dx/Eb3wDHiM6DJxyYVRBdPCf5lDu9QDTVLM3jfpRvP1Ln5
W/ZRsDqB487v9XsLDV4MQIIOQCXyIcLoORN5cGJmYBxocTnrfME3WfKssofUIvhB
XfPs1AW5RCP59yfMlpnNVzhn+2hQDY/bBxBtga/jIzvHjUA2yKEevhsy2mRjN4+g
vaUH4++mGRIWyrVFkvc0+qGAJejLMzJk0FO0F9d7Vl47E1IsttLCcDbq448PEtA2
zHInGSBFk3RJVPxAZaazfxafbSHH933ibDNGIucFl1YN9vi4dmarvbvvECrE2jh1
5YKWJdwjg0EjZ02L0o4q7zns7FoKUZnZLhBlev3xKR6xkdiwJqw3ongn9PBZOu1e
ABoGTPdMDUu6Y8nwhPiwzCNgAeYNqkykeTbKCuo5YvhX7yhYESx/1J/oCZT2zbwG
zAcwyPGOC3OQ50srOQTe+L19t6stZg+dzrMbZRfvoGAtz19oj9h1UQwCFu5zVb7T
4SvcckEwmR55rG9ad5xFCuNsoJY4T8b6igCAqHgRZaTELlH1bCvNctUtHLid/Zps
i/Glg3rrsGCUKgKLCIPusperOkDhoQ1JyWnT9+A7mhS2cGpvbz7sdpQWFVkVrG+y
HxaiFTh0Sp4HksH6ay5gGgBHL8SkeJ8hF17XOr7+DcsQzZ/u4ibF7hQdSltmXe1v
FILMG6ppulv2pap4fBCHhCxMLpaOeoUjls6HFeYwwsvNbqMCLSya4DQAOFGf0E8o
sd4BJKIsVuzEITmwJqy2uFxvmv/xh70G550lsUMyMfGvgu5DYUKO+kwYji16ERzh
r7NTr8KC7KcTJjEqOxm7W0ny31Gwty0fcFQdorTK8TZf84XY29JknqoSakQQxCMz
/aTzVO/lHDarhJ4Pjj6gGvKF4ncc4R93B2GNewkenbE/qC3QdjdH49qeDAQydXYu
t7iPP9QfBqoTg93bc91YUPry24NXjsY8YQg/ACpEnOX9ryWLECg1/399/q6R9Cgp
VI/7KSF5jGATwUp5C4JEfd81WxXV0anBSyXfuDgICQ1GoE8Gc7/HTrJys3GoM2O6
De+42LjgtVmDha4o1nhNptiUruuRxmSE1YT7MfAxtwyZGwkjVN2VuHm+gWftjsSW
XW8Erg+mq/lWvEhLdTMl+U5zi+PF2U2WUMt5pBa1cG1yv6r3HB5l5pBkNEFGRLru
SrDDPe5GgJnRtyMtGJdzWlel8Ak4Y42gOonYNUEIPpmAIigVNP138TMMe/PdPnO9
Vr7bgrT8Zi9RoI2w/PNyziOFasH72y+qTybeaJdBjJi5teGG61SzUVQ9jFxDEqHY
uxMfE8pHvTXK/jl4YTWLRyfp3wtBURCHJWRzYyYq8N54IYmuuHejwpIcNq71HR6J
qGmZwUrE5JguoCY5X3TWDHnoB0RCdjhdMQf/w9LKc/SkMpGawkmWyFdO0kL01wgH
krix415Vk74Zc8azn7mwuGOMciUH3KQWsHjeswRwEmDHf9wK9eIPzL4WaZPu6sdN
LrAghO64wiMZoHi1ewWcoj7FwweDI9Zt2kvlrjQYefWsbuXCDHrprHb3mYlaaMXC
W0LhelFED5FOd8Ap2KoktBDOWhixE6t0N/asdFNubzbJwsVCeFdfyOGb7mRnlnln
ygtn6lRKysL87EP6Xvcb2erE8q/XHOGWXsqo/fiNGN2ZKHg6akCaob+KR1miZ7Gs
GUQbJx6nH3iiCJaptrV2Pvh2etLJH5fhUV69Y0QZvdYmQt007VbkiXsx6gL/A4iN
pKRdheleSw503ib2OANADuBauIm0LVZ9DqZDLHglUzhEBaJkP+J9gvXCbxzQ5t5e
NM2Gx0B73lrVANw2F3DxMgq+76SqEV3d7k1wyAVo24ZII8ZCkVvN9hbyEBMvBZ1W
IldGdej1xn7i5r+jip3S67T3gFxCLwX/V2kUcQhjEDD7C2o+qeVgvmnOxNCS+o6Y
YRDAqhouuky2Xl0V9wEBNctnvLShzdsLkF1PH9N4xoNSlb6dJc9plDssQxHcPHN4
YuGhMbo9DUuUme5Gj4rJqq3L/JQjXSHiWsi1gpUpDdjya4p1Eet7plMFDsJ2XCXx
3j3yIGLdk0tGGUnOqMLoVZmi1Syhlv9Z1Yu11oBkpQvnRAKyjjd6EEhsT2ppHKhx
pdLZkGj3dUaje9tMCbpiopRGOyTGLe1Q3y8IW7IjPZpYlm/+dwFwlfu2iEnPgj5h
e2U2jZ1ERkuafOQ3/6OkpAC63C5qMOOLjG5orUVPT6BZGy2lPDN+muSgBkLL8DUt
EP6xSTiPe2POBDnnhKT7QgG6taSEiROqbGCSY5cQqlGx8uRDzasNUwgp86Ecqdp+
whJ20z9j1+0/qZbEmyNYZjQPSeoU6O77U9TLfBUrJhHL2EtE2bL2l3NLCNG6nZQG
PJKbjTM16g6V39zlVsWALDVkNgmjpamhyBNMM7/9XagYlICAYJ9lHCjnVCM8Wwjr
QYthzdWIesiWEccAZpiHX5le9C6zZ2F2mMG+pS9O4gy8xmXvEwJwC6RI9BgVnhDZ
skOyxeG+k9bnBq3/6nMfc7m7ARASNUGwyCEkjPNk7ncWyX6bMULpSPqK0mTIudG9
OFM/eWW+S/V4J9ANiX+ug7MuTVxKd6uKfJ2EYFCkZIA2a2YfYKlazk0lqSATgAV9
n4NJlhtzdIj2UV4S8MIgYRl4/WEcDIOBs3//5wSYIcHL9xlG906cNyg1V4V9WIb5
V05zl3rUiRZjR00TNPHCoMepJeU4f+fjIuHt3pBFeQheWhYO+UXS0p/rMsQHWtHB
LM3+Mln5GSTb61UiVg2t8N59L+ApLJsJCd5MCxw0a69hFsB8/noKdfrcC9xMISAb
SPZmmOMylpre3d8W/pYCwXwmfrO413LKGoisfJ8gUIsZutQm0oBOKM9yhgIPpQ94
QNOR5DbHYvCxS/plnnYFaBgwcxtgZrvnfe8UE7BFkqBpGGiqUpW/ZSFxvY/QY3x7
MKT30dlH825Fy0hVC1Z5I7d6lvRvCUwHYT454/3IVwZ3J0cMd1tdzt6MZMjeYJyr
0qy6wNqBg0mbsUuAtusCVuwA3rKp5FyJ0fN5lf+YfNZ4qqnR+9bEf9CB+jjAgmTU
EJqeERxafWcdQ//2Gxup5ZIadG8E4xUAqTVD40sREl1vGVRG319G5yP0XEk7lR8+
mriYQhzCDdJmy1uwAA1Bwxib1ZuDD+KibXt5b8j+N6bkjZ1/33eh1QRTmy9Hh/UV
74NgVYFwE2Bkb+W2R+KXeGj4qRsGAUKnHg/UT1mfLslOHHWvSxB0zyn0VMe7cK3R
ER6j8NbmrvwgvOlITuMq4XlOLdPN04IuLJjAB8GUqT6vZYjeir+UdxpMHBiUCFoX
GjxnmgWYip4pkKQ7uMpRpt09TMzsK1S2JZti2Tp3vWTua2xGJn5Y1c6OxtQbTdRa
0QmtXmcFzM+tPW77+7Q4uyiAEICgejyXr1wRhOywUj7+yyh1ME0BraxBM5yo8m6O
mvUhRoPefhDkJsXOYgZdSWmce+8Prg8MHqF4ey85dlRUhPqcbo0LU0pDZ1dbFVa9
ee4jMYZPZUTHE3l7gvsJ1BIyR7pSxcXtsPhLaa3cizFw9M/UYnAaCB+59Dz0AAQ8
ZM5Snw43B7BMOYHrPwNSKLl4R5tH7vw/T1m4gwu5Mv0tdnHyletjzHqAGDZ2HQCP
j2FCy04uInEFMeVR1t6vj+ap2v63piSVjuOFaXbJnro0A0qYrLnsZygQOHHWEAJo
h4hhg5CDkP3rMmR4miMBrK8hgcAR4og8hrY+IE59r6d/eRPngmygFoxib3pIC+TN
QB8kpN5YKokNBhDYHr00EZIx2n6HEVLGTfuaXoy6zHoXOJs9DR09cYKy4gLZd9rU
4qAhChHqy2x9M9TVImeOwZ7QkeqBgR3uuVrni00GRwMQZGvY68tKfMQ1YT3CCsbi
t8Ugs6Y0ObOzYT4hg0pLI9BRgCmyVWq532mXwPwzIb7nPwJQKdYWqamumIpBM6XL
A6mbzT6SdJoPvJQ1FGmJgwvu3cQ3Ig06ED8hbfB26J0gGRZU2E675wyEkO6le1pE
/lRpOYaEXM8y5kAGnctxKq1C4aPpoIlcfrtoBHgycKr4ApX+1ZFrooDB7QEjm6x8
YpaQk1RfIAnX24zADVFSvzo9GwNxb3QdYGvw5CEE2mIQMSa730655u2SQBJk3lME
TYsenMEMOETMZ8xNKS6qnMGpZBL/WHNllMIj1uiRjlOQf3oAYTHFqNh7foFWJAYg
AJvJZ81O7hIQ+8cCWYcounsPt7Eqvlths80IUp0hHlZXkpjV+y8XZcAWewcuQQfR
hT0HIfHL2J4jbp0yMuH+7pYrdSJ6NxhIcfQE+8b45mh6Ilzl31Z1odCoVvVL8GYd
UMQNY7ZtgVqH8maL4e3++m4Et4DACDLa0xxRap+QyzbNkYv68HWD3fy2D5ouh7X9
KVLxLoa97WfPmLY6Tp9BuFkJYCps2ayOgsbaAzvuKOmWZjCAWq2NM/c5+VHbGwbn
gGMN95c3fN0lSQSOLU6/qdfgJSqdfECtfN6nATPWcTvv9mR9BDgAmpjMEbLMrqnW
8/V2CxsHd0Y5t+45GhlCdQad+e7FhjTo+qlMYZ/wSNZR+/SV2PZfo45jkx0AM1JC
SfbXWUvgSJxTtALqsLTs0DLUHI9I2V1SZ2+B6+sRmbUNKFsKCJEUk7hseZNXgpbu
imGgB1QKu0ZYk7eiSW8KXZwi51VVE+Q/dX3q1BW5M4E4E40TdEesOcTHFOAlWo+B
bIQ4O3/MPWQGcEQlFYEUWBOjUtx7ICd859/MndMSKX27gmUQH2PduScMwKskxMNf
96JhTbE1d9lyV7qPRk66yvdsEjY/BK1LRROl47QmiF0h6RnePVSY/X/MgMVqOkMD
NRt2UYGLrRCmOrwMnUGd9MuyHkCDt9sN7G+DKPPlpWVnTwBnsTOOPXL1vif86q6F
Qj9jJ54j9hhM0/v81Cs+DlDHD0jYHBPBqFl1GHs93Y1cBP9xG73da52JOwhXTG+3
9IYD/doaNYatW7u5lvy0CaZzE1P0w14abSpUjBjSkiSxp3DS31ZfMMCDJsyroBrw
ZiF+wd/acKNwOYAnxVo1vYSI4ushDFbAnvANptm3WeHzGH7o2RmPmL2kK9Aim3iz
sEYdSQ3Pb5HYqGQOKut4G6B/ue//66onqXNcTbaBh6IUk6KGsRsfSK92Ei/f9/RT
Qte1Az7z4Y84zjcHbgL66O5S0uM9Z5xjkF0H+9749HdF8tfeZppHFrhu7b+3eZNc
sVQIa2DVh2tcAXx9tvQgQHIhGVeTQ96HoONUvy1NtZP1oWrzTOuV2gFE6Gj4AhMk
mDYdYDe21q2rLJvMgU2vSCb/rj8MopQa9E4HXfHLeidGVctH46sIaytYcZRABytU
XIQcqh3KsCEUQTU7H8LQVfdSBXVc/TDA9QwguxlnKR4HzAepLoN1aqV2scAEEkxD
F8le4EXI8rA/Y8R/gvXJBNwmQoz8gZUmS3OAY41q78ChxnA58bHP0MageEMZGUkW
33rH4TYK7FVw+Cmq8OmKFprjWhI+NuGHATQCilrwUx0yWBuH2Ur7rgvrtIX03//f
FJd7C0imHbyQ2jlC0tucGxXd26x3C/HplgRsq5/8PUavRlFRB8j1MJqYiYBxSOjY
wOsr5Z/Ls7y+Chq6UufiDVJu7vfErDd+l23Y1Me0QqSrW9D8/6OH6TIXo4LhVGAP
e9XJwNISGvOwFWKtmhU8t3ANxbsCl5duM2lqgYnKfp3yWotwBLxDa8loG22tMUWx
MRkQiWjWYxTssXtChN0sLakCs/4FKaePZu5mL6kP0UhTF1INSeBAzj71L3AxpRzl
A0Xkbo76nQ7E7SnRp2p8ZkmRQdbrRCrTvQS0lfulmfPMx/ZySO57qpS9CubZRQbl
u9fgKwnAQ1R25TJ81Eou9tEgQPhiOGRPMywe0uVv5+40b8CS0eehplBjhScSjTGR
xpMpheFZx59iCeQbfB63OCIeYeLdFg9IbLpIasL0ozRhHncyFy3H9J2hl1492moD
sRIGnKWmx+OTdWOX664tObOZXK7PKgWoXkehvIeB5bsAOFXOP9rAn9EcPM4/Z3MO
PQJBPObgpg+1SaRa4kR5zjmwv8+rIElOUemsNKryPMNwlCuXHd5jqVnlM4HXoh9g
Mx5rzLAer8qK41xH4VXtdKHM15n1fA/ca2datuZQ4lMbqqc0JkuHdck2P+ZkRemK
t9hzOA3aaeQXmW9dlquezk3IrZqK7doI3lneeRzVuxziuIREOMBMEdYZbsF85kHf
4vQw1pbH4RQ0P6Hre74kAo+5SUmk9Kbsh9la12zM4TBdAZjDXCZM6uuK7hvD+o0d
IAD9WXGRxXQKP1aupR7/6c4GliI3qLFHADFYa+bgaeHd4xSHXG0S1llL0Rl+eRIw
Zt9UBjU6Rqdz8EH+i3wEVKizEfO5XRDyZUTfuEEPEolq5+LQqadd8NmSZwvc5siM
b44latwjuSHgtBZ3XiJtiLNKDLWWbcYEu1ccLi+L/d7cnUYwaJRaRx2dPEZKbzbB
ULTSK9GfR2LHXMHeFlq+58oyDEZseNg9RBDAlpULEouBtTcDdPzLslTd/dj8mJSR
vY8X9HXgEwq7QZR3b3djzoefRQJfHtNDxwcJh1RUFjK5N7ixeOIhjw0WJLrSaSie
/P5HWHcVza06Gadk5v0ygfM3X8wfurtEdJsk52HLGfaYVup64RbFCqxzBAmaYEmA
7AfEjw6n8Qk+OYb975aCt0vEb6oeeSeAFB1f2POOp17R2MjwDvhv9Xemju5O/Bf1
dxa67HxFhnyIS08nh2jPOEGuh59MgPUBggno1e339ITRkt3WSdp4asl4ocAxt0P1
jUCpAaGhkUFwVkeGu5BWqVPNr1YjQAChusVPAnD7OClDe+wVTzhdNPxnJ4loZ64Q
JvsBucfY4MQefzKjPC3t/nQ+44FprfwY7qVw33BaSKRpCGNERx6KXM7/MaI0/fd1
9f792/3939d8GNkd5ujOPVB14O/zUSpXyydm/e7PfRqqsxjC+zfBLNuWDgB8Lxpk
PyJ+Yf84SObSzj3Tk7DCmATsczrVmqCEacLDJGCV09voWYFcfWdBSxH1JJxqd/93
42tmgxsbaR7sj0GDMMhpfZuMQDDSclqptTxOgXR1Z/uT4eT2u62Mxu3gOwWt7hp0
6cwP3ZS3OIgoB6kgOajTkER3+w4PG5RcjeUMcReCvgO3qKgBpBvomSMGl4PAXbnh
nv0EmuZxFGYHoZVB1JtA+AdVGtN8R6duN3LWzwYkYDb1xIhJ50+9KCUYn+86Xh8e
SMENSxyWOdgSg3ywi6JuH/a7p2LcgUd5JJAcRuj1NZMDqyzJXbTtwUK7ItrFvdfz
F7WSURp/38jTf5xMqjq+DoYbDtjo2W0YFdBlNqjT/lqdseGtJ6jvjNcrV2I7j1ed
ZhmEbrCeIo6xQQ2Zui6sU2wufBhj/yBPnSn8ylRCkmGOWacURcnjUstCBECqcqlR
8A5G7S7nLSRurPkKipLw8eLnD91ZLVmZgsvzSz7Tt7U79Ys8VEc4ULlDhmBQv6Um
6ECfO6cfSwXlfYV7QZJSda7R/Nm3G3YTfTWxPpcAvAgqNkfS6MYksYb1c5P9enIx
Tw7l0zU4OFI9NS8vJy9j4jnC7ngmMhPEpI7EcjgyuzdSIZHqBMr0JiYidtG4O+Jw
WHgjU38AuQvmoqBfJFMgHjRQxoJsXSAS8lU3zj9sA4LJSXIfwMciA9fddc9bbpOw
Yse5kH/oXIFLiOem66oiBDhh/ToO9Hh38mNouTAYslVLrckIC44AGgR3OOwFGVSL
56138UTJyGMOtqA5hixz/MAcPbAAsZDtqdipD3/U5199tLUC1usrolYxBe5NLF30
IyHTJZ3Up6d0AtjXs1iryIMbdzBDINas+wYDG+kcQRGs2CqOsqSDZXAt+eMC7EPF
plg+qyjOi+qxeit2HVwEdKOjCkRxCHbA5dHg2cZXxuaa02W5So3qAjia8Bi632Ly
wmGbm6YbOr1y5nL3pF1D553fB9dvHQD1WOhJlzdjJaw4tKxQ19yvCUmCWT15wY+s
JPzm1r0bDA4GyeX3hvl68BPHRX9BuNpILBBSRrdPQxmJury8c3vblDUxleXYPUFa
N7GLnaaAA7U9JKXUhE+y3nXQv9qtxq/mUoO7lY/9kjVbaIVUbEQ10LrjMBTbPieD
s8KLimiYUuMfZR6bGaxuvX/rwcJbjww6wP5C0sRo3GwqQylkMaLal+uA7HbyHNUg
pg/gy0Yd0cyufBSgMBMIpRC00xaWOe1/8frQJUi6k2QcV9eERoy2dYOlctNL+i1n
h0EKIv6uvcLyQvytB0MPWWmznoZeznptzx1slfe55keotMaMe0GgnIEqg75uMH8J
Iv+apeWyxlg/n9UD6zsKf+RSqjyMhVXgsMzVIfETIG7EH1KVcFsv97glXXiUJxTe
Yc0CO+kn/XFsM/N6Iat/fsTxecGyAEJH6xL1Zfdp3CaSxng9nkQyKeRHdzzzw3ZE
xkoa/p/L2nGPnFRMG48fZt5vQXT5D1XGGt3YjbiKwsJhp3UZiI2kXjOkIeLSjMSZ
Ca/Ej4ZLrhKzgBXh44+eek8LXyJGdUoSl8QmDwjBEg+nDpMHM5WDK29knm2TtUY+
CScxuNEaS+BYjmfXXaAyRwjWsNhjjQ78YI4Ze1ZCFkgJajvTVVnsuKbFvId7xB1h
kN4W7o1q1YkcpDLOCZfPrrBaf9epH5N5Jk+rLQAPPupeXB9Wl+P45IYBixLb0VdH
YPQnnyPHp0STjSzf/rlRF4zh0XCUD0nMaEBukJLEylPGGCuX9j5/vp6jZGe7X+Y9
NKJ6BxzpFuNSxWFo/gF6DKhjrApYWz7gyhtyp6l5+7QMGg5UhM67l3+o42VN7G46
jXik/EIN+EKWIaF/Ugi/uaplByQp8KkIsxjoLACVPZv6XVrYqNYYIMfKAPxPLQX7
HtIl34rpS0acWeIf+tV16WP+HkqKGLn8wUv6oNBcKUOpq/IiB10YEZi9EWu2yqEq
ta7WaFQha4CNGwm9/bFoKGJbcywWzhfErqUj5bahyxH9aDaTgf0Bvsr5v7Tf3CgQ
VNyhAiv9EAldrQZth73Rcslt9WQKYblmHrPawayzrMHCoVyM+V8WIDoaf6HSgL6F
ybI7j5Gy98El8pV3id49Jm+t8Fh76Hcg0mY4jsFeLdr+rvHO8rYEGLIgYvAAgo5W
H2UqWQop//je7lkyOkBeCff/MXonCFHOkqJFMqiHSOwS8FEY24LpAUZYo0Jnerg+
rC+NiFSUdOVFmQGbqHXb7EDi/Q8rFxJ2DHFH7TYt1GmKmHFFa+ZTuIbr8k8p+FaN
8v5+jvMF3fPu4fPV4vGY8QFcsrtp4pA82kfdNCSfeK6TkwbkdbmMhuAqmoS+MQhc
g/cyLkQ2YPWEH1PJnzNyZ4Jx+p/sdBi7mO6cuMISjhkJR7CKJEF+rP+VnYGCHXXd
q6Xn85HRoqQIVi3gh98xOi2LigoaDcnue+jorvwIO4Khi4FxmyMdSAStPBbRN0Y9
Pgc8Hl1zpBscCCTU1c6x6x3PDjXtSAA+nD2J6SzacWxDroQsuEgBggrr7RpajHvw
Z7rPp56FPMCm0vDWWEs/Px3mGw3S/muLM7nU2e4E2IHXVv/ScA27C05uH/e7BUZW
VgqHc/Ul4ykiynjKtw6yip7OX4u3Jq1OO7c8LK+p1N+qAG6QEhmaHw6TIH0jx/Qb
trNGM1ykQ6EOiPxx0UB1tLVscOaFDVXD4FXuj8ubtusIFptgwrwrrLkxlHx0Ne82
Pyc+4SXHdqfLWmxM2p1tY/XqJWN1M52MS8zjzBamUAu2u6mhFsz1qIuGGp+smO7C
xsmiKTI97S4lQu7eWd7hIAUDL4rf7hmjl3b1cJSCKPBRlQHEHnNatKkxR5luerub
y6VZOwBhDbv5fCL8i6AdL8UtxmcJu4jxwJE/8mf/atU+SwX57DALIj7nQKvOA1/+
FdujURnw2gj1CU9jnKY96LORreXyvVwAkKQnFZWk39H64NdkUiCCtXiBQ9/zh352
YGZoyUOd1Zi1hNvid397tb2q3E6uDgq/FSBfm8lv4uXTyUZ7FolX4fjXdeqpbz6C
v2wANSF5EfXyUKczyQNx5yfsOHX9qWU4wvQCRMcL3LmMpuQLn2MMxLesReaWmTIW
4s1VngcDZj7us4zsJB2S9Ahy6rL17kKzOXNYMifK3rbzOoeGyobt0gzogEWjahpu
OoOpoR21uiidzasQJOjbp856l8iapTSBXOlqasjk9+CwfcA9GMtdPRPgG8yljasF
FfOZE8Q5Wi9ccUN8wWZmCnsi4AcKzFOEJGPpmUDtvX39AX5jfqOrKhrFoQHHRhyz
Tr0zoGzUNiUEUtxwjLbMgV1t/0EgjSsUEkWU68pUcVeQ2zTabY7MLgK0CgCmV08f
uYtB5fwl7cXtPYwisk14167CYtOpO4RlmOhiAK88l7N8/JbvWIeG8675wsFqZMVW
TD9oDt+fa23gQfWsaTlziap5IRVj6h33vTdFiCtn9+CB7xWmPyqT8/pbvJ0M33UE
HdL5Fz/VX3mcVpX9AtGJHEs1nqYBDHX2NQjZgpcAMc8PT7SRmLg8OerI2g/rfR7N
cf71k51b5jmDDtmbXO9WyaMeYKpssGMatfUrh8sJOuo8PR9fFIvyTsAW3xRNo5hs
qGq5JL9jDorhFj4qV9HRt+X5KUnyYjvAwcn9WTva56Gnne2mqi0r/oFhG41AMbMV
IaQnBhdVXWCfiSQeAxTO3WEeDQ16vDcg8sEGJNDc73qRQXwICCYqXtKil6zdNQRL
mbDpSE1/jGy74oz2lJiixEzK/lnPHMtIBwbMKqOpN9uNCS+SPzeJeL79yTCbndyf
N0aOZwsc1BNH/2Uun/ou1g3BrDVyWPBPXBNWXJ/kGBGB7C9usoauGtym/AIwfJd6
sgdymGk+Q55XmHmyZpMRNaeV2rp1yLNAEsGhl/cUn7bQpDXimHxg8912F5hLHIti
bL/KNqisEv3rzVJP/AyZUb+oCYde0uWuk3rQ2Eyhp9xNvQT3zekCibopzWUZV3EA
jOST8jr1oWlIRi6dEjclyIQFrFeKQAbivO+Wm1t/drT7syiwcAPebkY44wUfb5oV
RKCdbZOR8E7uWZB44FknvGKRmOfadvlZQaVxZCgZaojZRxXeu3IBzkJmr8sY3pr6
QQYW31+Heg5gIejD8yc55G9vY8bko/14jHHr4R/Krxh2dRFc/TVk2Af/Yxi7j+/e
xZIti49NjWViteTK+DvZLm4WUBkRMfdj/1ZUPTBKgwxOrF54yBi+h5fv97kYnQd0
gsAkXQ4gnmz864KCe8HtAlvhOSQVPCBopwDPXUjSDZ6aAeDrhGIXpD8XRCkAjDPw
tfX6LY8Xm7A0xqsBWUcHjDpxVVuTpel7V92dzcQlD2xph6GLVT3BuKwJMAe4AlNb
nO2oZSm3EfKNnq3eFQIlhH+sqlxm2jWul2+gHhM44DJLIhEfaNE/7KlJxytEnE0X
X+sXM5eZdDxJJ343tdrwECEDFlCWzjlyVT+CmfyOakbXoAfrt86s5A6H68h5wAcT
7x98zDgSnUpwuWpEipqwQnSaArMCV1orme7W5uilZwrW++aqw10uwl+cPaqOFFKP
zOjbbn4Zlf0kpEzUvNTvvMtahjbZ2nr/GaCyh+cYtQwrRBR6jyonb1NPXyMirtQ3
ujhZO2oKLFpaUQDQpHbOnVGLV2Zv93EvEXR1Z5lB3Cu8Vs5wGVTtLvwdhzAnTp+G
gCp/taR1jR+wLQ25wSYhPShsLXNqgQaXDcjxp0Vsc0jdO/odVTQHNcO38jRFMl+I
pa1TGhvUZmtRp7XZUoieHQvK/gDhCW2xFHFX95tPD2WgKxkikiZM4I/jaaBjUvrw
HuvPxK+nfal19zKsSoBKzBwRGqykioVJde6vAPcUupOjpAgkoJfV9V8ZId1Lsd3Q
GJEwnHx/ZV4tYuQn3d+AlCxiscGXLwdX8PUtAdRo5pvvA2V6nkueDS+Lgqi/8S2M
/e9ppQzbilL0FLx28s64VOhqFFp+KGzaB/uALtejajBM27I/kO7/2AHb18izQa57
cuo09o25PhJZzfqKXyNS88EV5TSbeft3OydkEzzEkkNtPJ8IFC9D2vv1EnAgunnp
otXANHeHwbmOagYTiKOgBnErP15qNpKXBUxY8Ki98prLs8obwupZbRA8URONF5E9
uxoActN9fy6rZ6LhE1VKGVq58So/jtRlt2YzbuzqdrZgCWg9J/9UyPEK/qNXOXEA
xPjyGkmqQAuINnP0lpyPjdixJhJWJ58zJc9NsQNbOzJxRVlyP7cha5HTvHlAFt1z
Pi5WHxhpw/vgB5617sWb9PSTpw0SpsuEjq26UOhDvrl7mw3KhlfuHTn0FK7qheJv
6bg10YWGEOt88OLuYvxjBXmXrG/JHnnQMKFpzKrJnAHb089WVXz9z7MkhQ2FAuU2
lraCtAZ0XaP2y5h8AEBy+FqWYxAStFBCrXWBcTONDiq0geTfrvN1fWt2We2VOzkJ
y0hMOjn8IPfhgmZAQZZ3c7a/afgeSuRzud/w4/pPVAgmO30f7zo4PVBq652+8znW
KTZg8EAWV44+EG2QO1G6JaVjqZ9S7ds0yGc8SASUBMIBvrFF8PJaJWT8aLQMIcKn
U7KzcxMi6RAcyLP/E2u4+WkDkKyV0CL0iOxPBx6kFf9Nec14ZVYjGCPBvvFYH8tz
uAsekPKytMtM5+xMXxwFI45jLIh3GbFGp24/o8KCizwaoyISMploEOgF/Ed6jJql
SQSy4jRPySD/wT5qv1zPon27ZLJZlNqpWa+YT2bEMqnAsuaU7hKxIClnXfT2Qu4u
+H2pLRx5U5BZ9u0psPUCmELIJlltU+A+c0NJ5tpWgy+NcJAl9o9Sf+Dk9WZS/1u4
aOKkmN69EkpNOejhuQT5z7BrgGpgd6ANb9rTt6rVznFqIM6WQ8I+EsvBfojw2LpA
zK/HZEF5mKodz/zbShPBQx4UT4CWqFpDXg7pJOJjmTqHnaWH3pbV1HYNoLFJimuJ
qNrsVJ8QQNUmy/uglcmWvvXmjaSizZR61gjp/3Q6rnZYxWa80Ig5gNMm80Cb7d4o
rCKhsoo3UsZYyVQYV+tBcRFdLXyNrRVkUucn8zbM1rfMynxfWZd6ia6GO0BYJvjt
YqmYl19NVZpGj8yW8CC9gil11efU0coxSHegYkh3G6nJdbDdyIC5EUsL40O68Sgq
KZqVjrRNtxbvMX5HesRGRt1UTfn0kkpFwpTf6FscNsmEkwPFHsO2SaVKjdLN2yPP
4z0UjjXF6NudYGP65ez2RwoO7TVAvdXw9LQ29+xfe5CRP4G6FCXtauzsS3EpG5s4
DTFRFHMJlnr61mUQSPAfNtGnfGZN4Z4N93Qo5zZFehzkSYrRncYDx97K6MKgaZwa
IivDtaQyGB8jnwEoyLx8OvZ5sgDnNxYNMtDfa2lLrfvAhCuZ8Rug7UuzKPAAyZ6B
ikwReB1cphVSy0g3qdQIpQWB5e2V4jgsAK8TLlGVyvGMR/DEPrEodXGbBdaBnlTR
2dfB/jWDuATvNGjuZ1GSpokQ/ciPaApkDbb0U7kAZBKcUfe8Po5vARsOLo1cFivn
6V9h8z5ztMynxaYcxdAIwShLG0cVK0/blnIKQFHlFJNjfmakDg1499WqU/Q2LhCR
+ykEAhVQfJAu0dEA0QkravgviXpgaHrMc80rq1wrYMyCX7jqECyKh46WPSdsjqUU
EBoArbbe0qaV5ovFH51AeIBy780rrD0JAXmpL2e5MNxOSZ0kjC4pTUjQHgZT2kWP
Rk0bIrxXXAzKw0PuHFrobRl4j93pW0fAi9QB0RupOajZUpO5pSzyQSQsVn0oZjrN
LR4alRQLslJ+7q4iGv/7ujTsmRok1GZlzrPR55cBvjMKvvJvF5g6o1U94687As/l
UWlF077fayLV7vB8C+uUCIVpkHbqOmKD+DTXqokKnTBO+MTAFRwlGjm1TXcquDyU
MXSkUC+WrdoHOPE5CcBkTUw6KMb1elImSPdCJok4BPLuwbNMIh57N0f/xYLka5R9
MZpqKw6al0xZTcqViWHTyyTc0HM8BGSAB0+9lh9sHvIhs6mooP5QfoTXiAfFb+tF
HlZcyrgrGa4Qr3BwFydEnts/T82q5cm3/ttniTVLvqYU3T8+LU6qBF6UNqOUeJia
H6QWYWI2v69377EAcWC2x+eUhtWf9zDLeyFs//pS81hHq7qYjFaQ+CKuJ2PWJYf2
wxIX7Lw/L1DAzvPT1x6mSAiD+D9YYR5MmLXsnFXTwGdaPhF7Mbc6Nd0UmHM19FnS
o1FmkAoNtfHO3i7v///zyJ60Nu4MmqmLE3AuxL0t2x5NnbrQ5Bh5231a3DElqvxp
OTm+zmi24hS7eMqTu7dZGTvln07VhqOi7sAuo2hCu5QS4qKXay34cqphy9SUL7YB
5Y9IWCi2HzQiEnBx49DNZAf5z/dgDjBXCDJMUMqQ8x2LXMYDRQoc5TV9KMLDpE12
jzpGAWUPu4WCopQeet9daNlXI+sUwrFBsyTQidSpz/yCh0uzA7BsUajIRU9otsz1
AqTFmFrKVDIPewPcjqWffmtyc+xFABt481iLhn1/sMPtNdUCZwVcyDkFqg+2/bGd
ICW7f4TLslwbG/3fu6xlX1QDuFsgFWB5RSDldYhdzLPyP+OHZeaD/GdgB6ezH7ip
6HQNi5huLzXhazzji9vR7qWJ8aIZvSStWmxwdRGqXL0iyHc+K9bR7pPuAwBvQTQb
2gun5424lsxZIFpWcqCY1AQqYsFRe+4j+7DOP9vfHDGTeLXr+ic1oKYkNX7qitot
HMzU9fjaheNFqPcfOG8VDmIAJH4v9ZQ8j8O07Q+2ja7zA2T4aJ8a+eQvteeQsVKo
7PcXYZcBrKOnuLdejFHY9JASSx6usT2zl1+XS6kpS3F3DqgtT0CNARPqUPqpG3So
VQdFHdIUFx8RW8W8nALLq2pzFFq5rYSQhzKP04Nay1pG5ovxBX2D7dVvQ9QGWcD1
vuV+AcbbsqZEcTJU270U1wJgKSv8rNmiq1oVrTQc2WNGpMF7NAm3EU6XQ/oLK63v
7CzwIn2M63HDmJyfXRVJ8j1idhq73O8EKXRVEUAHZ40YMXeiOZdR3ni6cIFL7uIH
2H5JaDRqm+LxGJmM/i7mlZGKP4BLs2BrPB27koXbnelCt06vKaRDI3bPZArfYzMv
e2DkmXBLvaBtTJj2e7p5M4Kfd/jzI9L5EI3b+LnrxUUg0ohB4k98Ag99ak0cmf08
oTkjAc1PoHemdrJuEC1tcz58ixs9FIwioOa2qThkm8hhDgbcAsVWjjdfIXaZPL0B
5Rw3+Ig3VDalTA7Y9KbO+XJHF6dwzRNpuJaMVVXn94fSHHl+kEBgXRAAvD+CFCS5
gQI9+lNi4F8ei5zGN+DFU4yKO/oUiPfy0nwoO9tjcwotpvyJ+BST9VrI44Jqhtk3
O7JpAICSXnf0EeyP14BCZeDnDZwPciACXk9tbHP3z7jgn59O/KOV7+b7bE7nJzy6
sQoiIIbtUHMPABD0gPxViZL1nZY2HndDr+oIlK4Q7h6kUV801Dw7zQddpC2JHSpz
qcRmv9OPtfWSPshMWdilSfxuS/UVVTSqSVebXpMbEe8yAFGPTS/AxzKMh6rE9gxf
HV6lHPzlQK/9zohAU75ZR527iNyLZnmaxlj3lkXgS+tu6EZaikXfqUVo0jrl/guh
UJqiCe2WiIEPdpbCw00XKUZJ0iKilVzVbEQu0dReAD7nv9ooAjSg7U0wVoFJWV3j
8qW+k2YXm+fAr6LD+9EMvzXKUbkSdzbdUvql5rSWKtV/dNawH6vc0fld+b/WoRcG
d/hX2Perk9dwMNCE9xTdMTEfK8VPRoth9R9JraQgSm81jNfagN0SPPzWYiTa/F7m
lrkzBZmi90frp7lXfpMx0EJvGstY4Sq0Og47SspM1lt8BNTTfw/4lAeJDZhefiIW
VvVLbfveHv2ZmWTP9sTaljT7pCPUPE16TpmqW1czK8Q3gd0urH9Hv8FnJ76/yzOT
mAHwhvP9F68ZmV+/0kL85ZU+YfICGCKd8QpNc3b+otzs+q0CQBZO2xuV5kzFwNN3
2mJK1JfGZA4YMlwv8OCRdH4pZKVDb74hVs74jHoFn9lP1wdiXdCYEnMDBDXi7w9K
RooFbCQcOfaUbzzrktw6MO4V/mUjb6VC6rFy/6Pu5WVWbx5g6z0E7MzW6U3CWRTo
7l9d/vufoDVt9/ttDrlC1VhqkWOoRlWNRJ6XSaaoTjKeZmKZVhzwAXgy5rLfvFUo
creL8/rj/zcOqMbjmrniGToWZEDDZZ/wgafXs0hGocUQYnP3G3XSgmpuXX4qBsBz
F5cyRVQ4DslBJLKMLiMfTDoe4iltoHVNEzVUfar2ls0NPUhswsUpB4LOC4dzaQVG
2sxUEvSBalF417rdLLLW7ug9l4chciFhliT3J0dANltERuwJXMWh9fo8WQabD2Nd
hWwM1XpzSxkW+4hn+ZAjwGA/xK4H0QuXjUC0WaKpCOo0XTUptP67UL4w46353U9m
DsKIvp0ZIckI3RpPEGDv5exJmonYeMWh4AefoxQ9Mr3FGjAEFwHE4vNPnvGkZrr3
YiI749RsD1QEEIn74yQPr54FGD3oJaiFFHh/71RU6W4/e6RR0YRPaSBIPTrH5Pqu
521zc9Mphge/wagodtuYmukVl+WA1Y1zR6yNFvgUOdf4wzfPwbc+m/IJ0a7D/IOu
QmwP8QKejw/op5ys154zfQkIWdVWZ/zCbfcp1b9sqEG7gM+tndLyUrvtgKsnRzO/
bCpJEu5bo0VP5RilWR2qw/B9IDQF+wVq9VuClILqhwxIwwNFrxc3GqeNZVKDbaA2
O9PiniX1bvf8UOsVS+3kYitKHPVvplOaEb6BwQNSRlck3AVaAp9rwvgr3OSaukFL
knYgYp/JGEvdXpzNzwUidfw1TQUeiEtY+Si9SwmLk57DVP97cJXH2ScYGXWBMkmX
5mdMzHAM50vnfqQmX3nzgfn0xdz9oZj/z8Cq2RAn7jbeRgiVLA1zyVVzp0872j4T
53MnvJDX/WTuk7X3TZrUogkXBtECKPaX0gAug1/gkPyeepa0j1x8on8kKeXUS9NS
AD0SAkxSJM9+lK0Y1n3iRl7lQfaNmac0XJv9YGrI1CJzCbCVxESI/lVPC0O7Ycgc
fxcC513mYdVm3OFF3y+aQ7WMtJHJvZoCBMcLMTnGIE1hKoDM1sGDs9TDLGc347qN
TEth8lZMpDjwKhp4D0e7e/HiEa31aS3qHSf8iyAzJOC1tOXyT98FmmOITLgq05bK
vfppLH3By3awGftZLOtQweTBUuM8UeMQguS0b4OfEAuI5YDD+8LST8p81g4t3Tmd
S/4V+3b+gJa2vi9dxk81Ol3pvWLcUyFTOTaGXMYnVWWKgTN45yPG/M9oMURtYWp5
tcZ8Vof3wN+Feu2oL9p65XahbIyG9QQJ0r17GMeJaJE5ZohCZMyoyuaCwnnLNhIR
Zvi6qin4enyymx6c7/Zup8TVdeH6CTLcCVQs/i4NbY++CCXguMjtUSu5CKrNJx0I
/7z2Dn4d7gfYqK6LIr+tCDMECc3kqgZeWQIK0JVpGbV+/UaD/fkfjK12huPs6IOu
QQpIRoB5TcEmN5+UESSR0Bimg4Jw1wATrbvIwLaRP/uWW5b+CSmDPO0eZ5z+jItn
S5OY0a8ltmXmdH2b6nRB4IgPrE/4YtSdfZb2rIqzAHg69ReEJtThl7UJHP0k2WO5
fURL1eORsULJ0Ksbowq4Nm1kyqR2vD5+BMAHU51vy2Id2XkIyt/wlucvNC8HB5QF
UThgNtkBgJfrb7yYpXCD1b7W7r2/Gkuk/BzTJ+nUD8ajr6eXAK3fjv4SjdIg3mcs
b5oI+ibKFpi9LVoi6dL7jObYUqOTRV+RlDPJTanQyutMWH7nhqpfuROtjP6AQCpo
CFdiwIcup26IrdOzQHjCRbKkzPUzsMLqw5Qs3CvenEgqPqzWLFg5WAu1QwWgtV1Y
BlcOV8PD4SY5UYlterM/91wmmezgQA2q9iyWQoMRANfHRYUXzePIEbPsjtAQHawn
Y43D5qCQUovqdvqV615jzgzojcOzK8nFamLRZiTzMiUZTteb9NZLjjrjaVJ7BuGO
CFs2Fcb7gcgO4fchpfszrCa5YjK7SYzOQOnlR0MtlSynOYrMdo/LfFasXc39Hmci
fQbyM3PeSimSe5hOckBvAfBY6zw72V4PEz3LlLFqV53eaSOZUkqeJ3q84/6mu4C0
wFLDKfsBUCqUg3JL/0pfFlawCBMffAISaCGbPw1WxHVaL7fHRlBnDT9w7sX04rO6
av3NGjmZWZNgSki6+wsWvFpGUhxdFg9LnInwzfYbzIW2sCxIER3tUO8LvSxriImT
dnGY4KAFexdITskvSKQv5LQKNpS3Rtf1PuV/6PiT9uc5CvnRw4F45/2sSlIf8BAy
jwGqRs+Zx/7EkoUE4057y1o6qQJKYNYQ0fpMh4irMUYaXL7eQHAzxWA9rr9s85Gb
NWkGYdEYzSpiFDSN7LHHfVPMrC7x/PC8OJ8oJ/5lTpVyrHmsj6NEL8Lt+aZbN5PW
qAml/G1HUwmodf0mboN/gPOXqw4ASUsJe7z4ryCZpI79Ml26/BczNRZDGG9Lpxpi
oq1nkjQ1ZTf7h+/4/dbqovqDcHpQ0WrXJeuqw4yA3GNSudkYl7e0y88ZNX3UNAEu
4xKJ1peuuHcRnOp6LhWsstScQFcKZDrxcATEPwo7XkeXdxPP8kwG823f/xKxeS2Y
4yZGP+agAZbbEMfExiXdRmWaJTzAGNQ5F4to/3qwphgLWLTIzVZMyexIDwo2lmfc
48duC7a+3A9ABH4xHFfyKH2UCnJH2ac5VmRXlmJ4CwcQsKu0IPYPt4bgfeYZrlCZ
A8kGMBUer1m36TofFVg2Q5Ro4pMqg4D6PqV2NZR5tBOYOyx6TzItKQSSJelPIZkM
D6f6gm3uESegy4yXBXd0SwVQRwY9wHoL2vSD5Xw3WsRvNKP6NtvZT/ELu6l4DUdP
F2uq2mOiG1wXX77Di3kCuDpwRrs+IoF3N+o1yolM+TFf8e4WO72SUNmO/pxcs3Rm
1wlqH5J8zU7tToQZXg4iK5zUM12K9paTCLeeGUVu5oIJW6vDqYDUzCwuMmGEMY2A
b0cjDkuIJ3UKFPvJxm8u88p/WuUH+GI9V9Lltt3chh8fFNERn/sRaSSe+DnP1AKK
viMUOocV6Hre+2e3yO38sP8QBPN73OSa3nDKRmEb+ptM/k0p44A26jkK344jQAVi
XWkfByoTdL0QlCQ+XGwJ2AD9ZqA4PR4Dam0xJ5BPlTpAD+l66+PlkPrANqiWAc3y
dKl50gfQL4ExhRR42DowKJRfgmeUZU0IzJ1hQSn5idgqoTcXkArv51GPlym6Tkbt
NBtCjKQJ6/hM6to/vDYKrZiGWPkzVW2rru/9VdWHftGiLyU2N0h/SiNolNR7kyIQ
DigeP7pRwP4Dj05BZxNWe8O2ev1zTclpqxSTCGF4j94B4rb1T8QiFX92mrsCZE1F
nyVTsxciuhv5XWVG+BQaqqIn1tXY9Eecqs+5n+pfFZlyRm+QpmQnnxB0rBV6bZ23
rJCUVgYQkrXfRs4rVjeTlJJNF7HId8FIqe72RAMcwrzptySwNWijo/x7xrNU1kMN
xCZLMdmbM5Hqrpk3g3a+Vy9wJu63uXh4K+L75H3AVzf4q6MwIVsEwrqFWXGrDmx9
bc2mHjj8LeiBalQiXQAMJ2ycUgILt0FczpIC9+PJ0f1H6Qk6H4cgfV5pQ7W1mT44
IRN933/t6gIPUiwkq0nYqsvZhi9eiTQIFrz+9GNCZ/1PLfcAuztc6OgsALQ9AfrY
5jrfjI77pc7SF3Y3PnV0b3NdTuYz+cUgoD2RBeb+zC+WYnA/v9fQdcstUrCRNcpP
DJU+ngWcvIH2jNWu0/t1osUBu7GDFBgqCHrm8+xrNlVmFPb4s9bcVgEGhAl89vnL
x/z5avTSDCk2dr5HaWnqOLu3FFx+qRndkyrKln466OBoGtA16h3m8r9Co1TMz5fx
JcsNHF/DShdCmxSIuBPfdKTHrFrcvlFvh5B9T8ie7lEMSYNuboLJFv0yTglOmCe2
Xp3uuCJ5drvDWv0fFSR1s561uEpIMBB1qoWzpxUNBRxGFh1kbgoGeCoQefIAyjnx
73hfiUQqdtMiY3Wl5Y4unCffKtKaavKLxCZagePitFYbHvY4L5CwGE1Nu0ktkOuq
y2zJjFR/cnHOBiMy8AbMVfjZDqAQUiBNaPWMU7lj8EGvfVBKV9Y0jCDfkI6oBxeB
0IuYVNPHSxIj4E0w5tNXKslNV+CwR9YL8fJ5APGX2O9L1Xi9eoA2lH9htjXlmpKb
ZRcAw5ajkZgRN54JpGtHrZ33dUxKfpIdu3Zms6klb5U33brY4/9G5+TNL+CymhRj
hKBL64VIxrR+LTt5LXTOSGyw9xc1ReCcf3BsRBYH3f0Xx1r10OOpAwoRQVGesbOa
3QalE6Rn1viEzoZPZesNuo5PaIWyv9rwgbKhDIhGpwGMf5D7S/zy49dEDkyjwvYs
a8zJ9JvV0UqnyWmWzsbwLaVkKmNgzprZVPHU/x8i1738eW+ZFUItFQ7RhPe0tkq0
DlVDcTznI8qvJhpQtiYMycRNwulZsBpnQb2JFXaph9U1cMRU3TntlJKsNB7iZCci
qylRY02kGDEmj+DMmX/zSku0ssXEH3/GDlk42YO+u/urVN90RBUT8VS+881XVUJs
dgbXpNW2jXiem54eutmp4351ejb7nyKGc/E68Hh3RX1ZfYvaA+/ZLDtsQ7OtSHbG
J+u8jIGVfRUpckob6px/tOOfBA17bM06DECNhgclFQVcfQi1gjAkFy0rL40lD+eF
BPgfneAXp0uDr3XJrfp7Wz5yzSslCQ65tBoh7KQwpuDbXsFRH7oZrlJkwOqT8XbX
ctMu5n5aD9EEmv1p3N5bzWDNEsmFSXwJiXneEdE+yT/nQ3gWUhMHYxbnhQgfUo/c
PNu9r98Cc+Q9xGqjg4EvVRlOq0TqSiM9+EdhadrUlNFmRyarwkGdbzwh/104Edmk
W7ig1mAKsCflD9B7u1ZrMAIrTkb7nHB0Dlnnuui7WOC96QbXdS4RhL1783I3Gc9y
8NTwD+H6WXWIgKRknrgYV9HulrmBDXvFT3tUPK9QjuJLfw1jg6u4j0FRRPD0fytD
c3PABvvPugf7PKNVOm2xyH6dazfQNfi+R2o3u5KleCpIDvFeMBa/1L+PRF1ylBnC
krtyhNdvWTJ+P7x1iI7/qPKvuO9hmMTYW3dnHOu5QmG4vN5Jv+HOZ8cl9nm+WOo2
EKZ2ZA/GgcbJSNE+TYYFT8X3FoSp8tPlEv5JXD8ernX5uQArsCoOlY38+C1iea/r
IsqGXaa4PYonAuV/4U372NxNtBja4M0HijRk54wyhPEJl9lTMbFGkdc+CA219Wds
02DbG8CHipS5q5Tt48HMS3BxiYrKqQQo/YoykI00x03VHt5KljpdoYjHF1U/xok3
7UxqyNdsF55LzUCcpf06A8R29anb9f4dpnNfnd+GyQCI1BmZzk6TlqLjmZpEoqpb
BgnPRpxJiPCXZMCTCu7U8BJK7OHtYAav1sh3kuBUn71gOV/a56yfCk1pzLmjy+I9
TDQn6xcBieqoKP/4o9BQb9c1sEv41+6i1bM6XRowCbIe2YQx+1e7V478e1caFJJv
enC/zQTqsqlTjWfgUUZwH3PUaYkiCW9JhhPlQR8E8xF29FwIqJTRD+fgRfXNxLmy
ttJAfcXg8I1UqIB9f3/AykXWcQV1Kd41fOd5Bt7POD7hM6m5i7nCkBaWXMllJfkm
EC5rVQgvYswCwVUCL5390D3aEbt2xZdkAqTV4Hs3wMKRZWS/iXO5zXakISVsFHA0
xyDhw+bw6w5g+adLtefd6wUKj4kaDL2YPy4IPrUTyDMLwS0JaegMsT6X9HsWjeaS
4j1cc2qPc6FcjfnY9q0XJ+m+6/N+u52HaeEe5F0tDyZpT8Zg4+xWgZ6pY/yNnqZ/
MDOOThQ17lst6ubZklh7cR/3hwX1QUCbnj9YkRxRH5xLcfhVf5VC7nR9GEOE5VVT
vs5waZ4g4sh5QU8uxTxug+DZX3mAwez7H6uYs0rUKKwJs4VlXM6nBVRWej8Of/LZ
hxfIiKbyeNpyPZCGwmHZiuBO58ZtTGslGMC7FelOcAsnSZ8oIWJPmMGWxEvibGij
5/j5QWyDgq4GccbWQzGUSAGi+Ysdu2g2ngmjbV9rMMPlVc2KBMZfTJw4GURQia+9
gZQy9hmp9rY8cVNdOjlTRy6nGQywukMMhC93+Qo4WGNyKRkfj6y/WI5YJ4XNhByD
28/dqLnXBqvtWIQTre8xWwDbkqO8gRlgu5ceyqllG6mACwGRkTp06MeqHFP1R+lv
tREkvLiTsDy37YmXfO4UYrzFOxMN2LSmWKYjEF0QuhamIhR4RZGqK2G5dv8SB9gK
cBEPXmeP2fZJUbRPz+G6HSQYdd/pClVa0d4SHrDPhji16aZIvEeE6Mo7Ol4vxy93
GJGkys+OWRDJZubOYLFeG3u42x448WQCdYfn3C/A5mAa8FC5CQaORAKs6GRoOITh
6JBPED1MB6wHKkcSUC8Fbi/P+qqrGhn8tinjUI6p4Adtm6F7ryatS1HafuuGSuK+
0ZyfQDz3VojLwk+SXoEv7voJ3Ujhk8mhdYL6PM1U9nkcyO0Ti/TbmL4xzXOPpsA/
BEsO3hNmcvf9ZXnU87UHaQWu//H1kEM/pXJcGf3uUF2Ipga7AcXdC4OR3bbVeLb2
1Sys1sUFr01PO4DbA48cVunPSbCVdMac4Z9Au/Yr7YBkPbCcFGJq2P5XprmOOY7r
hGEc7HwpjOawin1woV9hJoplL9DhRuX2FuX87EikmwvCSo+flHWZfXyoPTQGet2w
RgGnvCaXafyWJoCwvC8lqUYpyRgWfTt6L3gJSSVWHsn3VkHQ+2HJYM2kkt1YrH4e
pyvgi3slnpFIKNYyLL9mFruOmqTq+G8mj6zXB9eRVFKtIczkGyEx0jWF3Xbu+rlY
FEMz+7HyGbgr5P1EhacgQpYBq41U5EU3YCYpIMxpw+xbHSxz74Fx1fXIfiwYVzNT
9IY9svXfEwthSoC31K56yDBMEpBmlQ+q2b7NeHwJOhtTsMRwO7/h1g4103hiTzXr
CVvqTm6rcAGOoudT33bw1OuYu7sB/OmQzacLSINXQYcNlYIMDHcMjvXMiT09OfLc
/Xyp3XJuhLohAJCEWY1Vf17/5kaenuFL7CzY+ByqncRTj+Dv0z0fpX9EPkvbzdX3
MrGgk/C8scD7Z7xf9wba5yhDEPzEU2Bjrz82xDMi9p9mrRlGsejdGAWCZ5j86fvS
kQZXVThsunNMq0ljTFWCqegGUoX12yDk95H9Y6wK52dJmDHvr5Of+RBrPi7y5UK2
GPEyeRCUV89B2/+Yiyhva6D4FydpVNZFzbctTbqFlnx+AnNCQLg8u3rmvHzhAsya
g9GDpFY2lt3XuUIWc2sl+jVGg8gzKSdHS5eUhU37XCckPN3iupyq0j+zyM5KCa+g
eMipjTr5b/I9DkAQdS8nGc5zGm1tpw2XZMQV3vQIheP+VVyyNUHjK8Awh+Mupjus
bfPRVwNDOTcu0T1VhzYZdoVm3l77ghZOVIDzm9FFWkURAm4qnGqmBB1/bjRSKeQP
oLf1bfMqKGrb5Wu/R3feNpjcGIj4mqvoa1xwDjheooOyX99DkcXMxHk1C6zxr0PM
PIkq87NePB5AJC60qYWKKFPdj1mJ46tqtmT6IMnUDDSsJEgQX5wuanD0X8YJfEUu
be8V5Rv0RMHJZ8Zujm/c1A9FNjCWWQ0wfJWYecjilnMILmbNQtscFaMAdnhgep7p
DDDduLSsm5sSXS6KkebfWFs7uvyd6IWHJ/ojHUmFwGv7ZLj8UKjFd5JXccDu/CSR
WFfLWBDRYX78TEV2WZBSoft8N5CZN/3pMPijzN2V0iBrmtADLGY6E5471/wkMIxO
cr1I3OrjRakRqg6icVum+ozRreUowwzzY3BPMCFZr9BuP6pynapdKOKQvlUa2vMC
1NQlosX7Nu0e3EsMQfUpjL1IGe5BNDQq87oWnPmey2PSQo/1AoHHxfc78u76yr32
uclHFoOMhyhpfyv+RTO8Da+Z1OroeOUuXXtinnNHnHgTw8xalDra0mxKGDc7zG94
P2xbeEwKzX0nurVDUYdQ2nrKjiww4puaQHFp6panxQyT9KqWPyS+KxdKU1uZJD41
S3b2IA1rZKUVWCM5+aNaKt2qVSOgvVnT/til70TLPs0ELC7fGkRoN3rK28MQSO65
ZanQx3ICtbCdU8173KexAPWaYSbzyKfDTU6nCOIaEWV7x1F97UMuGATrRT+zwce6
27Q1EIy+Lxs4hu6EZMWApDMGjjQB3xsHacjkI2xYd1Iw9iuhEQpT7WIcxJB02gmJ
ioAXx/q5wdQsemKFEsPEzoMNNhGsiJ0mojfjJolg/1MHYDQ3aSGEeQWDEGIIynvx
md5/NAOdSAVsgX6LNhneg2rrPuJmYm1nXGzfED+9gGYRpxC9Xx25OhtUsYmHy3kI
+8vPfpPYnwsVeaV3RvKlPUhAkoNRZYW2AD4G9z55drX0Gq7G+kSctWygcgZHqqet
/E5Sn/mn2UDOB1k9qtg4qMbYLiaR116buEi5/WZdVoFmtwcAERQSV5dxw14KAw6V
T8wfrXhsl+CBEB69fQDUJqvpa8jpNRMEed8oPOnZpEvqigHWFJeYjRrBQIX/71B+
NxrNcq2fYTIycj0EowhIpEyG1KiFAza9A2Up0qEa6dGdyq+fIQMp5vBsjjyXToSU
V+oHS/WDe3Pxl4K9dE2DcIdsEyxE8Aejqm9smf4W+LCZ6XyjVdjqIr9wtEUAtssP
kwwTViIWsguQxidEZja5Tg+PRiemfd2tpKmG+uLDqRjHuUGc+XX4F/F3vjcL/upp
CR5KGPhedy0D4xf8utFgus07Hf7STrP2uxBaHyfPk8RHUi5wGKTrfK8eUnjUfoTl
7sN4zXOVnaxPghBq8AUyIgqDZi6RHB0DFmnFpfNvhqgnn7KZdZsAVtIk5d9ynngx
pxT01nMXdPr5+Z+7xkbfeFkjpIsTkjUqb+5Hio+CNqDe0k5VF6Hvd2Ace1TlY1Ea
gi7oJIggS4o42Ovlc/Al48NGrCchv0r3VlG696GoJsuvEIxraWddCJTYVgzpuW7g
j/QRrRPi/DDH/os52mVHecNFVnPQGCHf9HgDcqi7dqq8SEnqqF1cMMfS6wPp4pCZ
88s9dME2dwOWXh131YXYqV+j4RM8N3E0Py7S0tBLZkCXFJP8AumgDa1gdxS4LDfY
hAMd88476fpNCvPEH/FX2vgZEJmswn2ijqE7Rwtbk/tJpEX3kmcBkF9hivH7ODxN
h8EmpWETgV79yB+XHBEkMoj3bbajYgQnuWlGrBYB5U6EzgG1RlPLWskrhj/oflUh
FH9sJQ4z/FHTyTK/2192/UWIV2JhHz9Fa87hjD7o1eO1BDVrC4L1DZVfrhh4PGib
DeCcLb3W47e/nXL3ey1dIr9iWQNmM5c+w7WavRnxWvIc+bvbRlh30pM4hWMpF4AG
H864yepIvbY17T5shXIfWnDN4wmUhFRGhavD1Qymm2smArnFicpx44rZVULS2/bU
9Y3WezS53ASzvB7pcoougnP4cpKpGPpt/MG7QPUCfVYMSROQrVOH8fKV+k4rTr7T
T0hXhaeUEkhf3hOvKjDq9v4V2MNKRB8NnxokoJilD/IS132vtiTY5U2aiP4xF/2+
WGF0z3ZtU+BBwqhWXbJyS8d29d96Dj23P/Bm367AF5xj116ZPjMBTKNuhlQy+qjt
zzKhmQumiLJUq6jeID7xU68txix0jAtgmvqhf1hkxG8RfHzU2/hYzNleUV2j9/qM
/Gmz/u16hpyA8Q78itDSA78NccBFb7a4YPfpXgksEur0hdIgomW3JexRFVEHVU5R
NpXgDVLLD850yz+rxOvn4xnrM6BBDdRAV7Jqt1ttWyuxXlgq+UsGWP00wL1K3eiN
jR5sLRReV7yYYqEqlTk+f5ZZFR/7kvKWdDZL5A4juTWjsDkpTuQ7r7f5fUq12fzt
LJc0jjhvGIRblFTdRUCOU5xMenbXvnHgnZUu0Ik0dDDE/yxDiIw8jV3LYubCFHka
bpHt+cDiBH6mK78jj/PsP+FDFEsO5K0SV90Pe1tMNgs84EXVnBtXVVIuy/42qwUA
uoh925t7aOc6r50FMqQt0MrWTZVYiYKObn2yMYKXhnduj4gz0dCbb9gGBtrL37lF
u/Z1OqF+AULCUCYkBqMEJs8wHjHAyFnvvgdqrbF3vv5jgeKjq8rTYjDPclx0zQXF
B0yOSZQgIkN/pgUeD5Mf+j/rwei9c9TISPjykwtmJTQv3xzBSO9YGUrhV4kwu4KS
bcvh5TrdnzS4Xr0TW4Z7o0xKwtEqpUPkIRNlU1aaKkypDFwLUsuk2CJahg71lDWm
yqNR+X+22M+PV0kAfB23K2xpK48PYOJ80wePMAKCT1Wz+Ia+XERwhEXX43Jvg/qV
393Q/xE/HwEU0tY8rB+OWx+7WpUVC8YlYzHU6awEUms/bVK1xZXuDg9ACkiJYPGX
Et/1aYWr44FwzVrpUFu+IqDX49bnwN8IpceRWWA53ZlUjNbTqaQbcIy54UC4jg5r
uYr4wcUsPFDnCT+6a7hAl8PndElBaS0kgcVXyOPnfwmq9olpbtkDAxt7MV7NpiUs
aNwiQojAIukKhZ42kRwlBJJT/yL7KAUGyh6UhfEdvrBKGXp4d0f9VUmJa37QbO55
FRb+0FOwDfJnUvo/JR2fJsgSb8KPPD3l130Mwo8k2CSv8gfDTK3K7yiAjH0qsQ73
blI6kRRJds32P6dk1BKUxo1bzf038lFDnw5dmsOU1bf1Zi/wbcAJgsWwodLh3Sob
rzm5jjMOkuUUQi5fmMXNjz0SVR7Enw37jzg3XCKDfp5gudtLfKQ45tH62Tqg2Bzz
5QzTn3Q+gD7udFEk0DH+UjiRcUIBYW6Z6Xwq4KB/mQ3a21TicHAzPiDkz84rHTKl
LBi89T4EyyrrQY8gpZ6mg9QCt4bVw08HDuTGXMc5WPNlaG93C5B5dHn3p9JHvIv3
aLbQTY5y15bJ0mBfoQYtk3V+PFMhukQU06NKc8cIOChhb9KPnQq8WUuE3nWrNENT
UGtqqcf91WSp/AZN71/hMUsGg5i77+efeCuGVfc6jZZFeMqkPqPYuJ7O7AOq69Um
51qK72Y75sySSRrlrZMtyiEmMJ5w91UFJUnihxrl7tQz33h3YsX56tiLkg5wOL7S
gwh5crJdTcf7QwcHy7Xap1ECqPCoXL6/LqfHYEIioIn4RmMCfiS4OITTEPMv/RSZ
L4cmP+v3IBvy3AQ8x5OhqpkJQoZGbOHi7CzkpOZ+bNPNOGXmtmq7ad4sTPS7ZtYv
+GhJE8Y7enUWhjdGCLMrda49SFuimIlOHETSOXTtEYedNRpDgrExcPKybSd7TERc
Ei4qlA9OlbR9QNcJJfgVJQ+ZZvudOcXSZtRX6Gg3ApZxJ5fcV/4Pq505GJ36uPkg
uGsM3WmksnXoauJGgTjy4j4Tq5xaFTRMmfrOjK1k9TG2aUX/9DuFyl3TQ+VO6J8V
Fs0OyNFJVnJJMuZhop8+WcR4wheqlKftA9opeBG4zkg31mdw04JyMlqKMeupY5Ow
XNqHW4lnHcM9mhB3UAwTZcKhSBOTWH7U+pX+RHWieQlXPKY4TwB7nmlVS/G8U4GA
Ir15X9RkitvKzg+gnY3FIjSFKQLBSwuFfDn9FRs0lo7KAi6ZAj0lwGxQ6Un7YIoL
f19V7WNxzY+ZNQfl+v4kSKT542pgkIFnroQ+kCOL669Eb5M22tYhni+YZYWm8ToZ
cK78LhnEvag3ftj2Cnu1rGR1LcHA3PKy5t5z5H10ZQhznvdo5Ad4YBkE3Zhz48Z2
meG7bBSy37C9VehEaxtRiCz486AHFShyYkv/NGlNo2v7eIDcqQTywmQp1kTQUE9m
2FcChbT0WXCkH4cPjsrX6C1y6nCk2w6V6cXpzFkuqWxD5glocrTvUM4LQbS7JZZI
7hLJocl8dCtTDOjmvXu+7Z1TANMCltMDPlcRwir0Tw1z3azSQBwm6JetuB3uw4Bu
h4YNCJGWo7zPnDQHSEgexUUa101vfIA8Dwk4deEv61xfdMPn9W8w3PBE76Bjqyrn
jJRj8kYcN58OcQV0Jw1yocmqkvUtLkfCYrIgr8vj2I1VRYCIWhT3C1fWUUp5oJvq
yHKgcmf3RBJR1mWazENxNtUokQ7ncE5lyFT8yWXjxoO4/Erl5hvJwGDBuA1tg6Lk
ffxLj5JoG5QpHZ8BTeWcNw2PlPF+ACRwbIWXJIVPWu/yCo12DdxRBrycnbLJd+at
DwVS0ONJCYuGQ9xjeWNmALhtioxZo7IslTZireE6e481RmzKUL8t6TrpXtGP+UQ1
bMULyMxFlFn7M2AuP2SwiHax7IoKbyhvEwM8xMVqyz4FL5PFKnp44sfa/aCUka+O
KFRSBcXmPnyKTqUoVz3u8gz+iPGhAhIlbJLeY1FroCwyEW38mc50MptptfKCJEpT
77o+OStDlrAcRDCVY+sgS8myUZW0JyOMvDhEv1Wjmme4sSEg9UouSv2hUpD3e5Oz
sygWeBfyRR5v1/xIdposTgQUO1p+1k1+qCPb8Efnd9I8J/gn2WNhdLY7D3XGbiuf
0yFdA8MzWfXEcPc+h7FZibBX6Hr5hP12t8JUI8hPGQZmChvJACdHbeVhpLyUFHdU
E4tua+Icj4sDE+Grp/i3gwkMiTpwbdXVEeL0N2O+Qda2glMN+QCU6PrZiARSS8rF
DSvNgiJEeuyTkacR1kIU2gztvEJ6cNnp5KJcCwES8I6VIzUueGXNbbCL1Qe0hhVn
FQGgd3ueik9CZtieyD/bQjkD5fLKP9vV/I4qa7n7gwjzlnSdDlxsAN/pp7RTS0Vh
VcT7JwiBLETC+FIG/iLNTJ36CWevTnxQ5craergMsG7UWVtmZkkjrCHY+Ok6+Je6
c7jmK3Aas/wQ0C3OrLIHD+bPbYsYwAGlxtmmUkeGba3cOnkLXXofKvzLbG6VMzUh
VE7P0x19RhiNWsQOkLb6R+Rh9LpY/Nm5gvWW0ehnCJlW4880+ldKypgnSrDPZoyn
nGMl3aGTI2MB3fG1oSMMeaqu1Kl5mwPyg8Sqcfzek9t77ys2T7Sc1hSHX3p+CI+5
aCgGKQC8w6SVqStz+tKvDd1EiAjGwR4zW8//+SO8BXOHejI8nHTuiKTTJbunUHba
+ddYEEcWX/zVvKehfkj9QiANVekARzamRnRcuPdh1qlRJkiq6zTQCuF2W2FXWIov
VFRlWTT7fTuHGOGTp1NXs4Zef1jJWKMKXU2yUivf/5Gr49vvzIGDMwbz9PB0my+3
YGKh2LL+VtxfPT6kvxpWP+beHLXOpzjhjqlcz631cD13Qcv5swUHpo0PwL9h9sSv
vUHaHtT0z4hvtvTCXn/wvn1Xt+i0pmTk+VflqvQzJQqQjjMRuFlDErTajRSPwpbS
OHu0qzK44CxC18WttTSRiiZSw1+AN2wNjkITfasuV6cRZ7cl0ySQAMlTMTxAF5rb
0rirzNnzyblFukjQ+d9B9w2zyhxH5FUBn7vS+ucH6O2kMM0qIP6sUjghLqdton+v
dAuwrHY2C5GlH9J69kkgbafmf7zj4welCbzoY5v6tdjiL4KhKSQ/nnZ4PWOXdKUg
1vWIOnNZ/6N7jeTWg+sWPACoDeS2vrwQI+ryNHRJU8YwvEJEVatjHkJ0qmPFPSFo
zdnSCssqfg1/vO1C87OgXjuTAxWiKKgrk7NnhAH+BRVgxKmjHBqWuylrKYw+nKey
GNCPq0+6TLA+0GHQL3McXifldUsv43pfwPkOe0SpBpoM3Ei4yvKlg+Frd7uVXzsI
0QM1v80UkLhKe2HHAycURkj6uEU2GiZUiPTypPkCAUA8DMz1TZHvtkhunvJ/zzv1
TzGu1adltaFXazXYzn+E9itesIVU4WvMoUXFJH578dfLLhA++nImRcZV7+uglF6U
CBoNDinUgJVYTaD/nTM4RPr+P+0VPNNjlN7jORUFATUTB/NRnTo7S/uUDdISXOzf
vqO7GSGJ4FryR2cblKt7wVphcMQMuHBgpZ8Eq2aWeRCCw8SNPyIo4FmnBaeJrQzh
E1ggw68SGF1g+7lKSX/ai9SQJY8WkPCLnmD5VyAz0qgr4EPECJGvj84ONCKkZl2O
ecjcGIz8aeFnVmR/u3/5QaATX90d+DXln/YdHs4qLVw6CJY/nXXAr4wkKVggmw3E
c/EMuB4vO4uGIe/8YyV2JABlnW7hAl/PPbwg4x6H1enmVr/iFOISpoJFMJJEqQE8
K0uP3A33HQl7ht9lJIJ+ua40TAumuWyxOEYXj3PwuGvX+M3DJDKL1rtb03qx1vJI
2C5kLk8Upy9YjAwJ/ZTqlpa+LzdUPcJ+MzqRlaC0dS374PazWlHTSKXxUXX6wAuS
kMFmZu8KyLmEfP6Ftz2m2z6b3LEQpQyS40tRxD42cZlj9/SVcOQB4iiz+bWUin89
rBaih9CNAR7xnZkPP8xcQCWWUYESSA2a4o4Hv/Vw2za1BOumM+XEOtlm+SWX4JJM
UBVm6f/nk6uAB/hlGs6s4IgEwW+GXZDH2bnyJOCFakBcQ5V3rAl1yGI2tNStlckv
eAa6raJutAR7+lHDZT2SRky4Hf/dN7DVlnt8nOMW+vYzxCA/UgY9BhDmEv65oXS6
t2g/4gdcRkRXauw+lihtn2R5Ql4/qCvgb+6u82J9zI+qONvKeBJindleAwVn3vSo
VHM340Ivl7y/cDLelbcZOo/nON4jVSmcoz3Z5TIUIgvVVBF6zr4+Ugn9yyA+5Oed
f7amSJtX7nCkCLWwOBL2JnupTg/4M7pCnEOtpMXtVIavEAo85yrg1UhtVmPV38/y
2OJ69qZEGvyNTOQ3XDKTJPT4QTRjUZnb24j1MFlL698n0vEtc0lVmvlmUrPHV8O4
B/Iq7MrogkCfrDqHu6GUHUnvLIxpVVSGxnkYNA8rEFre5qThTeODGOhXqbp/SKmy
bTSFKudWHjgqqJTlzSlCno3YpN22Rq/Cp++xk0rPoUC8TBZ0OZ4zcElKUB9gEsX5
VYZLkeDISIQQ0qKDkhxbrkRVPzFvuUPzCuAcA9Pas328CwDH2/5hplHuL6zUwu9F
TCs4/grCb+nHtPOU3wRwxMCGYGexavqj07QWLm3q46dm3AtRSvYz3pSJNjj+Xl3K
JtmlPpClegEPyMWElFU5FSM7ylvrkPgasVvpsI4nrJTcHAHXBNi23eUarWWRG/6w
RLOALWGDKjTWcSzALoWBJRj+s2yLDsE6TnPiNo4lwGvuIdEryP+ZuJBaDurkp+ad
o/uIbM3KbV9ISbkdjIOVhdLjfiG4UygtXEHFacx1TGSTEdVn5OhQfcsEZJjBJIKQ
TdfIh71XjTi8Q4hYh+IGc0g+l1LmGJfSuuteWJOns3nqiAPAaA7rarqlJ4ELGZS0
GIucc79fXwr033W5ctXpB2XCfnU6aye9GiwNN17i37GKYsCM+pnf88633bknl/SU
0XOS075deslZl/JrrPT0Weyv+BlPnQ4G130tDglmZTEMdbA4YsPHAPFam9WtSWaR
3z5YdAZdQKspcMVNWNZxQMM3Ba3SIory7QEutcfzrb2og0CtGpe8wGnFL7JEopu7
WqLEWvAT/3hmhrGiJSuRggvHHLOVbsz1tQDWVFG1eHs8k/4p5hA0eZcV9mh7pndn
/f6Rd+B5ZJ4ms7vj7XUPmnOW+Wt5BZ7txcdRZLDKUbkehysxAUwpoWuX+JSN3thr
ZWbJljqCqQcok3xQiIzvAcBnNxNJgb+Lf8NUotyCVHRtWSerzOkATmu0yXU2j99X
AZq3DhLl4DIlyC36rBNOh28FhXYpkNO/0xjPZnNKQYRoZiDZ+vcBxGhvEuXwTjB+
AuHWZRBbtJq6QjHYPjXfT5N7UGhuiiwWHhnLcr0gOsUQ/aPG+OQWdAuyCeLwTHps
YvRZaxDxFQR60IR1Wi81lPEwbwX3OJZQTLoH7FgWUTtTwPdiLdj4XxU0wDdjoa60
r6S5LtbQdPDuT+RIxW27fQ34JXWMdEu0bfTi2RKavVeEZGC0QDBHp4KwBwmg25Zw
Oj3p2xtR3ueyxQXFidlxiMImDTI7BQyWFIKlt3WQfDC9Iu0cTTDE52Vuf0OSuIQK
+e4bmofVZUHXyu0CTGvE9bvZaX9/sPWnno6XkyoDqHGtSGEaZuvSJtcCl5+BIt6e
Lqugm/eCl7+TXBVomWlZAe1mnLsBI1YapspngdBt+ZsUb7iY+elfbtgiamOCEwwN
HcJKya0NPr9iPmla/SkUkjw9J2usrgU+7FdVbReo5C1cDYGzYSwppgM3y33an13h
5XMBBQss3Risv4f8v5T1QSGJgx9zYKRwrk+OJEhlE4hE2qirDA92FMxGx3Y02zVJ
lUSS1WaPP3dC2x98NGbl2Qba3lp6ng/Chpe9qkltmRZTSxUrU8yY3800YmqvHMzF
WFfAoHcQFkis5Dv0lZQG2U1C2bG2a9z2bY1lM9dIv+I7Cjb2v7aeRtziddnwEo0b
1MyxmkLIGEIcYo1iEyDnisM8tgBBzleOwUOGCV3Ac0MD0b9+OJ9z9qYQBr+WMGt9
buuMFP6QH/WiY2YLb0f7ORhT2JDAmWsgveMSxsSKNvbHomTlX5siPfNlajcTygIZ
mDcrjyzUaFDt5qmPpd+1x36Db3qSJIqA2fa0/TDjiP7n67xZnPtQ2KIM02zr94Gz
rJvHa8XFjKXAcH7l9PzgzyTjMVm+hgRvPiuzCf3qHfO4B5o6Yt2XHfGbF84bEC6p
oPZV3cJ0zMs2cLCDwYA0IqE+eHJWpjEF84LRjvkyEcxwe9z+aAR6VZa4NZOC9KEu
ZTRzLA2ZFyKE896kIEoqK9EsxXEfeodHQ7HO9sqFDDXXNFdTfVQe2aPRx8BmRcQs
30DSu/Ci09Vi0YyUC6vkqnaXDJL7RnBgArApEUnv16y8R7UmQ3Cz/LVO2GzlJSzb
B92K8aEEoW5hoSJ2DSoA19RNrN/SOYtZmalJ0aTxZ3aGpS4i+QpMBwPQg3Y8Y41L
YlB521XGKEXIW0zCvcXL6A0WCWuew/x34PgxMrlU7SHAXHPwUmXp9seO69PjJwsM
3WdGVMAdL3vVYgEO5qcp0uktuuJKZ23VaRewcezMMqiVbT6xgVUQyrVdg++KggCN
3Uk4fnH1glcs1qOI/RU4r18xUKBqLoyAZSthsAmzMpnVEx735iUscV9aCpD4Pzt6
68SKf0WX84CcAL/1CTiWIRnQ5Fi9nE+g/HVGYb2rVF51U36erWpCoxoD1sq+5onZ
puyBMNSSoGcCl+GEouiMgIcYQVxtqNQY2BMl3mT+MvmigeZiIwva1d0FOUvyHs++
mXcyQ9ScXOzmVNk2+RWU+TOFFdyEhuikg1BPcuA+2RLNqjeLeFF+dOw3drMbl5vA
xG9voLvPyr5g3J/ATJ/Mfv0D2bHeWKFuGuKC2KsPodAs/N/AOFLg8rw5OY69T3bX
ks/fa/GR+otndlebvHLYFZKP0HXw6teSllSjhMxogFVfLk/iuPlN3fMi2hGts9I5
XuhwPGCg+CHDDz59Km6zpLReSkqFBfLlcoz60CyZLlir/KUVUJxVbMTD3/TiEq9d
I9xvB+VCOBOFknF84hltlnJpz38PAfT5OABX8YXh77VOxVHdaCHKBe1dYAm9e9m8
GJpSTXphMbixivfq3cbApGLyQWLuE1kV/K2hTyo8ObzKiubyLCryD9U3DAQdGOYI
hd9bEQxnPZXYh5mdJUcpVZugyVfiwadQa91ea2pblwa16i/C/x1A623Bkh2cmHkf
78CFXfUqitrCTvo87L5VNQr5NkTs3mFgBhapGHeczZj43+H8iKMC4/vCat2b6D/Y
uDBig63z+kgPsgXE46YdZhHVEbOdoxBRzfutbrtIRLbOcxPVfz8rwjxUlWOTTZSH
PW8OgUK1/07M1bHXDdw2QZLttorIFlkAyLDNpGf2SAOa9IqFW8Xl5j3UPib1hddk
7mtrY2kABYyLDAcLkUydGDDkZqq5SG1PSq1L6dilQpQkuYV4VnO1FrruFWeXRj3o
GIGPP1U/yUdp1NIpg7FDdy1EdRy6bWXBeDzTGbH9rXQVTD6in4i2OQK+5eAMH6OU
iyWE3e0g61F+sKPvarDZRB6bMRIuU5LrPcpjz96jR8vWME8ICg9Z2OVpwEJf49eo
v2qKzR9OKiUwQ7WklFir1vayZyv67PpGlYMejCNCgDsDSzlTKJ93AOPoCiFhfweR
3NTpWfoHn9lLUUnU2R9N9UIXABJzlITqLg7lfhqu2OffwM8C2i/aPVnPM5blmguX
tMI7yl4RvEfr6U9NfPbIfZBmfXNRV+gQu++yIE2pJ++NJhZGaiOfxut5A35yx0/m
V+ctAn7xog1Nh5rpZDpZORnNVlu/68ZsybLF0Bau59xd1SL4HGX4zNA3bJmm/c10
/eT1zYYZPdOoObzHPem2S/zukYPEGozp4j/qHGjWz5bt2a4viqIgWELSa6eOZjd8
oDtRD2T4WmBK8zNaiGs0nK9HBafCuShMXaQA0kgvs2qI/yCuyyuReexlLBZYMQOG
57BH787BbGHM7eMRWOfYiPNOF90LqpAUnZuym7t6NAQYBRQsrT8C/t03AUmFVhqy
tCMkwOht9V3XU7MYfKJXkCJNX2N4/5vls9wtea5npjkEKwKgSln8ifmhQ6MGw/nK
YGn0Cicfc8t6+vrMQlEzpTfMMuYYnrbM85cy1+16NBBG1v47aLGlNWlzQ+nAQ7Cu
g9KZ/GOa4mnoprIZuyanNxNoS10s9iOzS2FHYwJ4bWuZj7oDvB8k/Ed1nptwbPhP
4jO3nCwfWbDRdgBLH14XfxmzPBwgzk1+YxK0Sy+KMjj79475ZfBFIs1RLHmSYUpQ
TxJbd+1aVuy8FhtHnp8s/khkBYqfv0Z/ptBw6LwFB3161biNKyarcz/lChdyT5v9
GnnnZSkU+M/Ne4bmlp7tgW3J1Z3istyDYtA0wH8yATY5l2avWgLCruohyTh8yD1i
DCg513jXIUa/GjeuX+qXdYribeQkuRoaL5sr9GhNTLK5fH5mPNCVul8aWZWSClGu
53kRYRdOmzZHUH1QIsMLxEbouNsRQmqW8twC6NrTdiBj4aQ7oV06wW52afELDVTN
/UjHqxfo9OdfFZLGIEcYaZpPUAsbLXyjxZBr8YgCmD1MNCsPuxOPXftfGLbOzvDX
IntlibtwA4eX+wjYkQPca8uRlc4NMtlOVE+ZswVr8yBSQbSLSuUpPU2/vAiO8K70
5ietO8B+2wTqBzTP5YqlNcSjj0e4F2+o2kMmQvu/QoKLA6eHOKkVxNCXhu6urFUO
HNaKRqboYqlOkYugpuhOERES1DeeaBygMG/sAtWPUoujacDNrsEUw9AvRGawR+Fu
FqqVwQQ5xtbMvK0uTf/kkemS/tVIeTyH+rCngoYv9DxtsUT9XH+egxpR5Duzy/DL
NDFTjtq+7m0GjHGgDtlxhqbdY0YuohCb3M2E7r3s9wq0TlAp/CaZwqVWjKS3aocc
7BM/I/ZUpUrK5HDXE02nnLrnFzuXEU4Oxf9NpmaZJAKBYY/DQeq/Kl8wuGpDGvB+
QKZWKIY+yOnxsT6H6Xq1wd1KFKp6ku7N9VIktwLYfM9d9yq87vj9brbN/2O1GWEC
cz39uDXczF4L9WxdrcRezDLRSQm14d1VUUZykAOg6b2OYsLHE1sD3rD1j6MvjvCm
C6hXpkJslSrQJvcPO4eEB2Lu5TC1pHBpeWsGpPa8pScpDYdD6w1wm/SEHGSfFV8e
O0HiPPEMGBOrXX/ffObmxeQ/eGT41g5P+0jq57C5UTfvm3zQsZugm3R0iLuxYcuQ
AHn98WP0vQ/YuFV3/cBhgff6d1i1FPB2KUSxxHbBtpQca+RC2Z66WaJJkkhoIhat
5iLBaRDQgM723YPwDJqduRT+9H1o+ejcJDeGC1108YgCAU1bjJ0wpantNCVXvBVO
lVldTR8h8KTFtUpTsQ6XSk0wY2SJJs8TVTgHoc1ol/u0+s96DJT+oFr/nYYrtCNO
+iH4t5S+6U4Pd4LDTRfyxvUPwWo0RdJsVdmU2SWnbpvGFK+prRozb7KfsKHeBoPM
bsrnCt604o+j5sCWnT4jOZNN39O/scN0RFWcnuKXBS1HM3e8DXrKtI3kdv83KDqO
nPIjDh1Ao1ycF2mhJVZ+xLRYuO25P1tk9mM9Y/0fD8pS9j0kBvqXrdvrYWmJ1AG9
On6maBAUPRG0XmoQowpU9jW0f/VvccyblaGk6wx2ghhUmu6ealZKuLW2mq+ph5c2
gTi7wPQ0rANm45PRL05mftMM2dXFoEgfizI+agW1U/wWdQ7lqbfKFhqlbSS2HLfH
iJ3wq3dK0OCQClFlBFla8LNOs0SB1mmx443JHc5i3sa1fSorO/QfmVG8oHmqyBoJ
cGf5NnLjy6L9gixJAGzEYck1/4xOTt1l+kzdMtCoTuzw5IE92do99JrSvR+TiRca
rQWBNcHfBYW7XWJL2e5LpX6b/2GkHEViuXCh5TNwjuPbsbx3RWlyk+Te3yv3pWDO
PeHeUeYp75RI+S/YZKlTuhZ4tx+Pt6XN/NigKiHVJQ6Xk1V6DEbusurxyYMG1aKp
5BCwev95jbr/QaPqna0qZ3FV8IRCejWI+LZAp7niZYEALfOB1V+qVzbUVpIvJsSy
x7DT/1zLuwetkjuB2xoa+5uBvWWF2vSLKe6XNa0D2kmRRK/ZeWC4mSHg9i0O4aVW
WmWsGpU7X5aN/jiDLCp8a193VLjj51Zt4hSoMUrJsMiwOFNeURspilYG/WDsRwJ6
aI2j42TRJiie4IWrzRUpF687sLoaILMm4aHZSv8Bwo9HPfol/jghFAKpA4QosKiX
+kuvTnNDb6Loi2Rkkln3fpRsC3RTWUV+EIxf3VPuA1ClPotbPRb+GjWyvSDWi6o1
/B+19U+hnG1QsDvZfRmOhkYOsrKjCF9bK2w7Yq/ZC2tq8f5oGgiaqu73hDLLZ8VD
o/Wo7h+KSEnIoVD1fmZkxgAXQROC9caHOEET1yV04cS387YrbcmLfq942UiL05ok
qj9mt0OPoYo2QTxWa/DpmGbwgigZ22xMsFLr8Bd4JSrfm9Pt58Qn7tJQ2iaF2xz3
2HhpH7mR2aSKiHopMpxwG0119KENIhMWlg4U4y45/Ja+gzO7JK37tXAJIc/ZiPuM
FFAp2X9Ov3jeGUCWyVv8neXEv8EfWT54CC0eApBENWtQvGiJSw9F4gh6nSMwxg3t
/iVEULsBPo/vjQB7YJuMdmtCaoRB36bRgpYH0ubGApNJlq+anB/2qeN2PsgYT/Fa
+SpkTPn4H2TWJzuAMR87D5LFNfGcv6ZVvXzQG+rXEqDJlG4Hx85SazirCrfIfZ26
/UGCpzEV2GxAZJ7ZFfyRjBguwZ6m8PfiIeCpKjwN4J4ESW1xHC74ROQ3uMjNEaP8
i3vadfYlE4DvqBFS3lMajyQKrdcEt6/25fyBfcMZ8+HU4Qes0rJi4E6zl3ID63xp
RvaBjAPcY59Q6qA0rNyq5oBj12a1Or+p9Y9XepDTwaVM1lPihRBvmHkiuxuZSLiZ
Jt8PpDo/WASdaSPJD+naCQm1vsKxfEuT82JmXN7PfIZz/7i9UcdNVszBvdvN7LYh
5PO24sGA2mQDGBv0dzJ1LbKr0G11iQryvrRLFxAlMO3WR3jTjXutwNa5C/KCAyFh
v0W2Uvse2d2gF97S6semcuhczVWbn/AQ5Dx9/4E118H+NIU0ODj0pJ5h3eDJk+Yy
k5YaPI+dkJa/c5YmvmpxnAnpy1sSdU/l5a69KaMX9YF3vOEJ2+7kxxrH26aIdN0f
rVGaCBNJbyqA7uxbinNDSxactVsGLGVDPRvtSR2GfmyubxGzqA9zohUamXP0gnXg
4onG3NuF4FBsJB36RmXgUsgsXXuYimYoMdBPo3V9UAoYCR8/tMg73WycBLagKlWI
UdZhEdvlb6l9suck6uNlZtBBmtCbiZ7qN5xnxx0gfA10R4f3flI6Wzu+bs/Azr9Z
vljRS+sGYBLDHBe+44rkMHQ7eRREYP/A8FtU/Htif29/I0Fb51k2Q4ZYwcNgqso/
KQ6qgIjGfMSTxgZ9m8MqCbK64vAmB6Wzmsl2lDZX5yN7MnMflJmYkk29cf7ADrwz
gDfzKVtY/AwEAsI3HQceZ3ahXdPJwpO1cskTdgIjB1e7cWyregegWgbR9jEjn7OE
Vw3vfiRN5ZKL6jb59G7F51jVgpZNLmPSySYOXelfy2BwaipV5mybgh60ZAjeqGxW
fxY5bnkBtd2hb8Ol34GDBWT9s/FWh0XvRpfWoVSLc1Llaeo9mKxcaWCTmLdBQaX/
cNtfpjdqBZ69f+MP/18ppqK6e4MRwSWZ/QH0rJLsOTRdKgmjgTT4TUSzyxgBBMk3
Ri9TqFmimpAZILNVduRjMLmKDIP782RYsdw4mitLQFBYkVlV/d5gIT9cSbeuYWgQ
CY8MI0EL+uHBW3dnJMiP6+9dEJnYQGQLWEHVmPhhdTxmOHbSt6NQNP9TzRgooPyA
giOk+cA6C2z9c/sLKNSNCJSolvp/ezrvNxckmOagJ7x+f43NO7XmdXklTYslN5Ue
YeSvnQJ8czNjIOGOdnDH53LTAcxVrGtj7c7LoKhmPU/wU+I0asrpLpRcwFmO0qlJ
ZVR0d8iBF0OvsMMcCm+uRYZad8sjr8OMVCQr6mfXn7dL0kZLcBbxQoIJfiT8J/Ho
CdCkjTpznizhQ8ufbRl7OyeiDsLUJGxZYFdu/CMfvj78ByKHxjHr3ucjH/w2MLL+
javu6w1QzH4pdm4aYbHdJXYd4IedfiFvAkouNPpRwib1TAcz+YiueBPg6b9RxcrM
DB7VtCBE22AgDB7mAgdl1zRFv5pMXpsU5ZgaXtflzJdcVV9s6dPRGbmYmmssdveA
6dqD6KsXzVS5tmG2Cbe2jSweoSTCoetujt2tZ8jBgxzFFyCu1zlvqzr6iqlG/O2V
we7swrtYONoVkiHQV2+kGbFRuxYiY+e6R0sL79syiaf3jHP5n2FLNGIyWbCKpqiG
gPIgZaYkSe3C4Uh1dsbBgfxbcIoR7IBpIaUsM70NeBgrs9Ka/kyqgr4GiZ3OkDMC
eBd6eZmqcOQfNJ5hCiw4Z1iLUyzI//3TXPg+2J9tEHOGKor5WYcTFG8FUoAEnUy3
JkpiSi7EUEwavT5UX4jdL2fmkCVzNb8P6BNScL1Tp37cd6uAwNTIOjvuHhIkn2iu
OVWyevrlNZrPC1cP9HzXKIptnQ596VP6nXmynUe5BBUbeNtzIODZrtONwOSoz+HK
XfsalGo3j11rj93VUotSP0jLI5TPMj60NDT5D5VJ3wGD/KzogLls3DqWqFFDAnqz
XP85UQpuYkmD8TPeaBWydqLEP2yMpfOuE8muMo8QR5mGcffAJ2d/867gWfxYdYNs
3kaBg57gFlhDGSCkUbPmAy9wPgQdmMVJXU8+yuOhmGdOk1SdAvsupz8FeArpZPDf
+PsteHofA7oipPKf6YAn0caV3FDPOLRO+GUSbgvganPzKYWXkLJXbz5fS3nTcDgJ
a6Yz8QpOBv6yTEz1om5KwDytTvP9oMXmb12PpJBoDm4MMjNGhfZQ4KMI49EmUeQR
duwSItBZYOzy1A4TJPsxxDjBVa6vTy/TzUIm0bmnU9kGuPTFD/uCmoCx9rO8tZAE
Zf2Zw9djFnIMybJtqdmYqN49w5/YZnRrJvV+T/Y1TFsIM8J4E03ZbPjbs0zcuarU
pXzPDxssonbSOTOqih8Wew42TpHHAfXqyi+PWOpuCUo2wwF0/LESO8aYNO9Q1Krz
kanpd+zD5XSR6ny8Ii2tIeXafZ017dePClSb6eRqtYPqGrfPdamwuvFprxS8bTtr
5DkvaTfYBtmvzcuEtNRPfm2wskcLcTHZryh5hSaF78/FvtzhpNRtsMANu80WBhb0
dLXEThzb3deE7Uw4L6a09dt9V/hcJAXTBk0Kxa8HP7zXerAglyvro49bRZ+OuxmX
U87D/8ryNgLsIUNuGZC/pihDp8E1wfRsRnJxUVEQ3s7776s/t9K8TsFSE1BFO7ko
HpeQn3oeXewww+4Z0PN9pMHK22Prt27bKiDymC2DEXOG5xL398Gm/Fbmd28Qp0X6
Qbbn2z4+5/ZjHxfMR6nGiPA4WxkDx5oMVGmlTno96j+KqFVFyDQro2j3hc9XAtrc
JkumtqUsZUtU29Z00FLpKMmaMUA1sdxgP/ntxzrxpWCL4h83IbiZvZhIJ0sIPk95
zDnR3T0TRWGmXws0B5t+j4GtS0LvSw0AT4ibnKchCUuSEUswVcCwnjPSmdEDPQFk
THG+I4b6XL22jHXsbbX1+f7fTK945sv3TYQjsz0fRW0U8ogegny6wuNvaVZRPKg5
oNp+dY6JLWJGcf6/4dFnqikhovzwsSiikoG3F7ApTy7aUC9ARCwN3X1lQFVzjLtg
3Ht7GHJGtAVCN6zQ5QggWvEeaEvjFYLCy5Z8+eID6/TT77EcGtdd/euv8Lf06pCS
4yWWZlRlQa6E4JYuFHSuwa/UHv7MpB2FKv4iq1jFKzgu8SsKoqQXnAYwYjNEVAcl
e6SvgygEqVuvRMTt8NGcgI9LaNQSkFPYV6oRYDs1IQRFB3ESh6w3Ue1cCuJx2otp
N+Z98Y6CGTFlCGms5T77CCWr2TndLho93p/kkmuOsFAyoa3gpo0Dq3iTjt0yQp6c
w6cqQtyQZ0l1FdgTu+xMvzCHvCX+sxdH/IjCLit0+Po6csS0fAREqfIwXWCt4F5a
ajzdCo4JTT6HUI1JWlBcnNz1I6qxMZOpoleDGSqe+l5Xqw3SP5cuesW71V/GuM9w
KNp5mAyIRm6D85bEcvxZ9QmMT0MtlfRySO943FMqechUilM7QcrhugvoQY0qHd9H
xet+HgqFTKRygqOjL1xSA3d9wdMQTsX7j/4zYXOaIvY/mZEfsTGhTE6pA8s2OAjB
oogT/UuMq3OIuXjswu8+c5dR5eJ+qPwd+yhS07JFZkPLINwY/Cg+fZdE3TQxKshq
ievPe5NMno1LnYPQo7VrMXlmR1TxAhpKBjNiNkBvvz5Y7b4kdzdMjaT5eq99k3Yk
5Z0Bds5WEI1+YNrSRkP/QHyx12b6gkKDrLhxw59hd5HIxKHqOSSevJvzp48UXkgX
3kUSuxZwemeJDrgBfhxgHWBF9/HxFIaesfq9UCmkk41TeihPH/R/gItgoD8GOjo6
RR8KR+hulTVxdHc8/peKof8KnNq9xKN3wbi6JS0irQJvau0f9FFko7EXmC7byhPu
TZ9moVgnU/PsW1aj1v3RdeSCwjAz87hH4ZqHrelVLWFhMDZ0h7mlG8sWLE82kiLc
MWkJB4F7/eu2cYInAQ4qlaDUos+O8kMO8FGS5nQwCqQT10EUXJ/JXn8DQnRY4boi
+4EimWO9l1iAMru1AKxTRtVCsom2SRw2P6swd5rOqUcRqch3dnhvbIyVIfVu63La
UBLcfJqenVvoLulyNVt8hKSySHVNCxOWKMRGIcWtJMIpby+AoLKMfrwrDSVuNHR0
WwaKaDKbSHqOYwkuaPdNBWPEc3NuLwSJTHQcScebXPHQLo7duW6ID5BfZKOhQ+vH
ZT81WIdhsMhOQjY4+os+3D5NNylCQ3YN6ZytzrqZlS9hLKkWKb288ccjl4cc9LNO
9WCLheD8KBlsQXKsv9p+vcQSxMdmFaCCeAKUXXqAwwx+YgEJ0m+IOxhKnuy19jQ5
dtDTFAoff9fr5+7A8qqKBYrt36vNIuy5gUV2XIsA6SDp3AQaqUECwgUbEGk9xV3p
EgTIT6JiGC0/C5+1tHSkI4MxOg7zVNrz1REnLBB3c/TEhp4Uv/QVG32A7IoDpT8g
fV5fyba4rN6AskZYBUr1lR4OGtzcDt9199hMf5hRIef94cAkhzyLWcqyr9jlZCqv
0fhn46sqbZrnLMDtT+R4+kQinoV6VKRfu40oRu0N4V/d0obqw8eY2xL4D9lzFJj5
0HOzBSwUxLmflYj2xgSPTmHv4Def3acqeYmbrAg5ZbTLEHz0k7r8MxFQN+o9UCGr
LrBwevLauEjuLvLjePf/oPsfZSSmzOgQa/1It9dtzCecIHeNb6G1bPxUSatGA8Zz
7+bBqfI1LuU4e4A9pYUnnnUBRhT42Ufigqy5CMDOgrRumYfdoMhGnjYdl4GHg5yT
Sxptju0p/Q1nwBuGXuOLsoNUt9ltlfGNm8shZ4WNwohfHCD4OVaH9E48R3NLTHUp
NxMkedd61HF10DBDUKwSuCV2/oDMQ3Njzz4J1ic1jQZ0Rb/BEw9kkA6+NZwDtCQO
AqJu3T4z9mmExMTcCYnA1ch0HHiLHW47kADr2RnGJTK3ocbadqvOxMFxZQ9/jtbG
g/WaG9RktKfQ3mCGsA5Nm/lypf+SPrgJjOjOFCnkn9RQDCFqvXUpMbB9RxNVzhnL
3Rjn/4Ox+b5tLIOWme6pGBSvn0yqfiKKNQRqCH1OPSXA3nIaHLJWfMy0fBLI9TJL
3wZlP7ZHQkyQTdtfLTef+wnBDUT42+5Lz07dPBvPmNevJhgCPuJjVmAdjh4jbehF
Br8lELnSAtU5oUrKIcCKxp4GIgEFtls9g0YWWUlQxIgEGlRx5relw912fGbPEyTa
p3AiJmEgjGR+Ovv5pba3V7W+/8JJ5JYQT4B3CMh0WsUS+KO13RW58SNRmtA1RybF
GPvy+65vIdtPv6hQiQxlBG7C2bS89pxDGwAT+RipMIFxtP6Fc46WxRmRflMyDGzN
yUf/xKl1fLxN//DWEJTG9vH7G0hBaZW6gYigo4l7b4M69BAa6/Z5+1HKAsM2+wKi
XS68d1o8PGTrURMIWdNRrTY+rUgWrm7GgY0pfFk7MZoI/G5VktnVVP9tqeODWI2r
q+AMJQWyskUYG9TRFQ+e2ZZaWuNEgcLnTGce7SeqFhf0rZPbcRCo8c/ZcMzw7hu1
pWoUEyDU0opldIV2/cG4BQxNINyjF9U3k2H6KSO6QmgDd2C79dRwUYPDDidWOA3+
IId99XUSd4+JA2PG9ktKiGwLcstSFw5gRh+W//Wo+NBH9Bbe4Poqq9nF8CPgyHDT
YdTD5dOZFlRDBfxe8xbmapH75nKp4ymf/zASvALWPgj3j5J2GQY//WdgUGmBfz+F
aIGGKL/8n/oYSd5XbEwwwqNOWvE4ISQwDyBnem8dsfoc27inldcz4XOboA5nlsgs
JkRzpdoaPNm00zb8LZ5DWi1g6W4Wx+EGQ5ZWjz2DeNWqH8DbrLU18C9njdsRJJMA
7KDRTaVXSILQEPA6QE6aDT4a1bFq/8FfBhdN7MFAjisqroiOh1FZJNGd2r5OJapG
z/RAHvYTU7vN9/1hLVbNo8jggSD86/iZIbAp1GzY/RdlOQQMbcPpmJK/wb6Q281N
nY5AZO9dWRAzpGGJvPDhuO9OpcG6y/Pr3+gO2n7IjKJq95QC0l3wA3HMbYDlRf+l
l3CNZB+IdVQjodUrX2uxRpr9N49t2HXG7iV9RUd2XMJInn4BjwiK/7gYFY0RdKvv
R0iTbe58eahHEfcMqtqzxGfAOSH9cFgBN5OaIByatPgVcfgWnEq0YsYhZf8vHvkM
rsC0bWcKJg0iN6YCZkYYdlZaRFecuquEY0QZwICkIN+u+E4y3RAyDMImDbUX/5/s
6eDadB+D3Ii7O+2g3F8+w52rSP9jk/WG5De2OCfHc/aKYmu0oBTzy+ZbdFUNfUNH
1UDS/ekXFVtSsP3eZI//bRA+v63B/0oUImNxZD0YrefksI+HdtPfMPCmSvo9/FYr
BYuo6HmDx+VWeEAabIYjls5q/UiThcBV94EGX22IBHEJ5OsFOZARlN9KRxAkhsJX
ALsIKI+hpFyt0d05jY6z9df9AazuhuOPWxVtXsiTJEd0NyNqHoOXjwubhlcEGkp1
Bez3JVOPYDEQe10bu0sfbUup4YrARrIX+gd90KF8XT+Z7uaviq4Vk3XG+CaP0M4h
GpSySgRWyjhTIRASGPI3AiY1uSJWfqcrJk0x0pjgObX/2IpDfvcIZdzdEn0WWBXz
lTGgrcY7O2H6rkhSMQoJnMtVDO6dS/u7OmHC5mI/j8x7q1j9euwBP4uo6fWiP9rM
sUOXmiZLY2nYkoOT5NDujxFRKkDuhzOUvm1GwX8BGOcozx6mAbwvrZ0xdEYZZ1Re
BT9Y8iIvsjd0FirN/CRPXPVIlQplHVB2Ayc9LOd84+rdmvxvGO4cRg2VJqUtX/q8
OUmvvS5iLBTpU6NZQ4uJobgblpSnk7MUppKF3RmNE/+vvnCNd6iRNORAX/UOXHmn
CVsDN9XjCSL+ZVL8R3qz0pDXiC2yO/LNRWCooPl2ObsBURItMRWcobMWu/rUQyV1
6oK8Ivw04lxKjEgHCozAtmg8cNFXT05t1p8k7Unn6YaWOXjqzHs+fVWXxlUpKcCz
RETj4ZlGG6pHvfK6Ay52IV9bKCFGWpoS4UnBcaAzdM40dgI4UVprtpZbdS14vJ6b
kGB5EyXvkONW5rwhPpoF3SI6P0H6trkRibSBO93msqyF+20jY47Dztz6OY9RKLXk
Mlr/Ma6YtN8BJiWzyTxkWJTwzkrD0PJODe+XjGG2745qOLRbEb3qBoYbKI96i/nb
QvJIfSV93iZQAZCJoMWLFhxRDscy0v9uBfToR7DZgkTL6uiGNZKFqhXJc/lwEYp9
dEkrlgAagSV7e1HSVITGE//4qDJnaTotRzGp0H0GqMwbIUOsXaWyrxMtBH6LxC9M
iii3FlHQbecpOxAayPjNGdes6agW8gOu/oICSAqHw0GGdoyFFxQwXeKcMgAHiM+X
4ZB1CZAcHcuAKmTrKPhLrPzkZF1gIDuGTXqM2N+qqY4mDOo6UTEKa5Q88AajMkSn
Ct3H5j5QeKGXv8WIrnv/g6KElsNc8q2SAzmg9pb1ZlScpNXugjlbNBwRZQvtnlDd
P9cjPs4KFmOBAy8FPS0b0dXaNOf80+fmD+FXERbbwsMozNjtVst+d8GN3s+jXHLW
BSoHby1nr4UpCbCI0do5Qw5M7EM6Fs9us5QStx+d4oPshjIicckNNTS0A36K+Kxl
BmyouZ/7YgfzjNaPuGH3zsfP/oJBj/ZQZ1iewn2qvRl9EKY7RV0bk/MI31jGuk1H
gXKpobbZulaeTtjBd9sX2hfLQl9lqxTLzgTL4sxdVOQh/3z0pYXVchQ6tydZV2Zf
To3OnA5gNVdHkzvaWPBsM23K9bX4vYgDV0M78BMrufSe3QAvxNJ4Ah5YTdL9XzdW
B1NE42VwpCrWGbaZ8sbqFHqdtcMrHPuBC9xMo37QrM5WWT1Git7yc6QG+OqOPD0L
OEfR5EVkWych8RkwUHcClWFZKA7TOcVgQ36D+g83had2RzvwLOQdmBil8lo4eRfv
Y3YiC2eE0bbpF7Bf8wmIkhTwdeZo8bF1cy0LkXOTw+9sPQnjyrpQLl1IRtnv5r6m
Qpv0FkQ4+mEpVO6KVXnV4FK3m6y9ftoN+TTyAc821b/AurpoCroBsrIkqFm5tQS5
l2dnb4YtXx7ukDcaQ+TGIgi5B+ZrLMkLFMLvVrV/p2US411VlVwunR6rxD+3ciFt
eryzlsShKJDmeMgEqwGAuZmtT+ilbDvUrT/SOVs+YuWtr+mWsizxPJrcYazWJl3O
AB6aZFpNG46CLJ8FLi0ab+YLc0qhBNlzY+TEZO6zwcfbGwT9K3oaC4Sy6/rn+EvV
xFzeJ5g1J6haDj912RQ5a9oNM7m4jfqdovZSVryBvsYX+erupqepHEiVo+/WDXm3
lWSQ0hWnXkHqYLdeywqPMo9yXclunaUx7XJVTEwnY4qVBDGOAQX3LovJ6rFNEEaO
OWsS/K5TwbNWULx3r9QsmxuMk4jPLDcYT54IxxCejv62IlksAjAH1JMzFHD13/Zn
bIG6wJbeePOEhkY0lI3ixk0HABcHVhy6HnmKQnY5uAQT76M0t4M5hMRDtRs1+mj0
8zrC0CZ9Ua2LMq/d4R0+6D2D3EPhem84B9mLFl0AdvKro77kFLZ8qglz5k0MDSJg
+N+B4mk3czJvAY8rYQt7pThGPaXW2SVAMvabKXwE0h1ty2bbGF2bw4oTFfuejYkJ
+umTspIMSvYR9LAHNxwxSLSnFDbZ0LSz5JJjY4YYlzxVbPlq5bd9umeC6OcceChl
z7a1yzMMBF1mOztQ80TmB7Yfrqi871EVqGcP/BkPhWUJATYEDY4d4nR1WJ+qEPHS
yk/P7M7OowvtjmI/Ovx/MhAyqf2OF++awPbFmCN2g22JqhPaH78/ylASMp8te9mC
iZ6khAtti23XkJAiibBhrRDpEY3V7Eiz5NAdAvT+HDuMCGBV2nAUCog0Zs9QPAmF
sS6+1ZCGEbYfAgRzbQDeoQSuvD6zJvq6MGdKAPod9nwWvtnXE8gY3PSS6S+XOHpE
IpATfJkTlkPOYa/DAYaGoqVzdxK88EUQFoY2B2BMfEXa+rz3J3zniDRaIPx6T1yb
cq2r9E6pFwOBhByebkrvPGzkkbgzebeWxnDWX6xHPimrYNJL6xWxj1Ialb6jqpML
we7JiRg3zyBqu6TsNdi/ZthO3Jlu4Ud3vBXUDQKFl9oKi98c/FxwDTWENZaF416q
dgV0GdFP75gg7AP5KGZHlAuzQpc3io/p+EIEcSBQc/K/6+Iua+98WwMqK2jZ79cl
HO/nPJnt/i+ieoRlQcCjqjUQbdvvDR8yGUox24tBRxGxIGAJu/Cz+2zcbE7xilPA
BTqoNCrJWBGPHXF3Zf4lG18esPe57i7aPbC7tAVRRNQiU5VW8EUConAkacVxcAkv
JszUX94S5LYUMwjRr2gNPl1SmLrCdal/cIWQKAAUi2PVsJtT9sFzF2kXDvI5EC08
bibzSTfnZDwFuj9M+tJPv1gvXlPt+w43zbUppS4Qt7ZpqboiDztDpdYc7AAGgL3t
fTgkXqomi9h/dA80Ai/++XHT34D9f4oTKd2K9kV/o3MkYZOSuQro0JMTLXbn9WW3
Q1znpHcOKxfd7Ap9BDvXQ3jK4jHrozADotCP5A+8dC6RHpOfvdH5RhmSXuCvkXzf
BQQHIf42MwoEBJwMBZqzglYJfLeTYA/wv6xTYp68YO+52eJRF6jHtNqTVPY8YFZf
WXe3LwB8gHhWkUE4XZ/2VgCeWSz4RLwVgRIKiqt2FJCgU14Ct0gK+I2CFq5o+cIP
Le0MdRtW/MhJwzZDC4VOSeJcgErCWhhQvlwLpZg4ziulX+Jl70q+Yv/3uWWVkyTq
jqJNWu/KXoNRm+ALonkBWjmDSgpzAWMytp1ify31/NhQJ92EEIFsxIsoW8Qod2iv
HyslXiGQx2Glm8v+WCD88g7mMUXeicY+pbFQrddeWRm6BRjnTSGqUsj4b0eVD1l6
eU1ZaEweC8etkmEXxnrmvOcUGKpfi1ozpfrVSIPw5XCKCaYLV97fI0vgn291TU0J
hqi1cmeul6lMrqEj4CAXvaFxTqk6bSFbJUrEn+RkWropSePTIF03T95nioVAt/cx
ZZY/kiT7oRLUxpCe+OIpTM0jYj2GJ5gMVONtvFNMcs5VHQ3lwdgLATvgCqir56nK
9xgUDzqoMf/HN1CfIjGDDj8ltPNAbsre7jYIPg7kk+8cEsZapIEC+bQ97ArdpoYo
2dyYNK4sOSQZ9wiUJrazr0LVVpBkgxBjk3VvtVh5CtrzKgWB87EhTGP82QC4Ndp5
nqHVyy1lpNqpeBYvkMoSpek/Ap7L9ATjzC8zrELD2giS4v12Pud35Ng30xJFlUmo
Y7sTejdIvwl0qeWvWqmCWtqeGuyUwI560A+1luDt7oy1x8Ogulzjg8szl1Cmb+xJ
kwC4B8faNru7PTzYZ4m6WstlMJL+fZlU77Pqf3a7iCJtcekRq2snyHBrciCvYLGj
jvXRu2KEd6cRuia/nP7cM8oBblmIz/W7xVbHM4iwV4iJDnjH5v99Jqn2QCXufxL8
74QNfRBWute/0AUoe/fgBTxtqSyh4jsDZhODCtPjc1JjGhrzwHzkZ9ZTYOagI9/3
4G4D9fUnmmxcHsJUYSFLS2JEzT9jubWxfZR1EJvjaqRe4AYsot2SuhI7metawhHk
Y5RAzoZ/8gw0EFF4TlTPN4klsQI+Y7WmhDHk5p+EryjBggoG6v1MYlDGTBE+uWlq
fK3HamliqPqvoZZvNsTKmmXXv9olSmX808RZb6C0KL91AlkfE4YI5+zuEUoUt0o8
/CDMIN4OtujqrkKO48zV9ihwai5EuFtVehbldnMmbyBnnNfGy1qGiI0CfWpLflC9
8Pue+XDIzPonKUFwTHDBFHVG9iXA9OHsRlk7dLMxE+X1sk+Jc7KKy5fSrIf3gfte
59GYe6wOKddrhcXeMB4cgo7bgUmWMdz/WcE327S9AEeLHFuewkBprWuryLFNKaJC
AXk8VXLB4Z/vupVANAyUXTcagp/FaA2mOrgDL1NcAcpUm6KQDp1qVI+dZW7lZaAa
hjvRRe1VfyJViamCDgLoIk1Iqi/Kxj2i0flsu5nCE2/pXKkT4a6er+9HWYl98FSb
3fzo87VOnLObnxW9RYxxsuFsNkh589WZo4bZj4b3rf3vBPwaHdMaanbrERmEF1t4
lQCn5vNs774qWjPipz89A4a0ovTXHJyxY+F0l4KDSYIcQfUSdTMavbiHxyamI/U4
zXPS9ORpHY1rLecZx+pQEEQSkzWgsHYgbh0f7nwk9jvIQrtSawRXJFudiC9uVvKt
c/P9ug2IdhXUEwQI3jxeJtvFtt1OVx1ZTjzk3ogJVJ6m/uaRfufGBA5USTXSPO8B
GLlmysQdao64FBPNXBhBhfyh+G16p6xqcP9mOZGrjf+xoMvKSg5n+Kg06bchE073
/+BW6AFKqkO7Wn7AOfxyK+VMVpU+yRrF9FO4uRHwvRGyVHRH3Ez/pIOnbY8KcpR7
Klp/kn1QOruebsXQPbyra4RcORRfW6d5wxeNaVbDFE7kvkhn53WVgdQ7vNm1WoPb
c3ib4VVLqYjlBiU6fUm7GsVXfh1Qlg3DmXzr7/LCDbsSLNEBZa//ViYkmHfcQKrM
UsXVVKqsXiy+BiWdIxkVByTGhPict8kafwORiEYKV5r7FgRh/8u5Iv0g04D4Iunr
QR1YOVOxkOxY1TuE7vkyJuvFZ3/xpIXH+c3wF9BZCbzriyb4qVOeSfQb/qguUq0n
Lpz8AwLzDNmGf/gQQuhoPf++9g372gEPTgeKa+zsHiYkovtHjWZqADxzAfPnPTqo
GBoumTSj/BKeMlyc9RqttJ9WD/2Pz94eunjq2iw1F15laRhyzPKc1g0Mp3hkmJIA
pAAEi50xn4ya8Ay5YwdQWsV0efxnr3VMFQY31YDzcl7H93wPcxcBIVySrqutUIU4
urb4XhBIILHxzSPlwUiks/GmqBCogheKqeYNyW2OLcJPb/kTt0eoJMtJ0zcJyZtf
nSIM8EePUa1+wX09ZFML+i8bE8jvXzt0RVASmUUMCHfKGaoGcy6YbDOw8Lrkzkdf
jQHlc/AJBGTP8MPWa3VcOHWtw3D+ukfWAItrrH9cw5pNpLUztDzcX3Dq8zRjSKSE
BhrsZlzDyyIzBZ7JBCFmukKTYmwB/82T+EaMx3xEarQugTP6+xXhkV1MdlP+N8V3
5EHnAQxacAVZQE90gu1Cy3sIX1jvK4igYW5JJsOO1u9kZIooOgPbC5Od1hoii6JX
4DhMRB1cnsEEQUqILme5GXJvQE1nHvKAdJr/G9Fwto5KgMUh7VLlBvINZB77c4N6
J6DzlWe0dlDJFmK/XO6qYC9dQGG1V2IB5E68VqQWTWpXAbU4lzBQnX5EV0/KGAbQ
g/PONphHwTKbrCwMv0NBhpLK+qHvSYARwxLkux23sGESkjLbwxp67a1r2Koo3uek
eVczInJqkwNe1yD1kpTove0xKAXZPA1snTHurUCMgvs/S4lYfNjBKdNuFRjiBeaK
UPaaIIyncGILXf7bIr8h6DKHiiK4KsOB5/0S7+HH6NuuXQqaERB0nnc5AroMqAku
EobuAwJOdv4ff3qgGXQePWdRA2AgSWWi/t48DNPtk9PazJJMptZWv5w5eQLxPDfw
GLjcPwEPSFgDnev3I3SxdcsYS+kBF4PhnHdNxOy6RMCBO2bKwRY0AgQMxdjd9kzB
qh2Qm0HSM3EFH6uHWVw/Wap7TwLe/dFE6FiKHYYqUN9HJhFtItScG+xir3vLTwbA
m2an81IPvdUwMCt3zIFgAaU/M1X2WgSa0n6iOKdDVU0MZuRYJMHpsjDF8UKlax/c
cPOx2BrN9hX3L3VXkB98Jl+iNxeNFKvRsqiJN6N70MJ8bhs3QthCik7wMgAD5RNy
7FgtsLqmLJMd+d4kfUxEpicbDTKX7/jQvuYxTTfhjJ9gI9BqkHjFeZmCL+2w/wII
Ac1FVI9sUBqn7CvzinuccT1vWLlR5NRxoaJv8cLbAXoPUdFpUA0Jq2xoZCSnnwvc
X5Ei9flcM6pv0/kJs2+lNEFVF7NABTlvDWNHbFx4NJqwE62NG75+ljXRvjvCJA5n
VXM5tiblcpUsL9bHSEHqv57GglqSXzP/iPiqio+VVkmuzDeOp3aUR4JObYnMb2Xd
idWk7P5GDSgvDiR+/a6YAhYQUXDfuVGMVJuEU0QTmozMAbG+q/fNy3tb2IivusK/
MgLIRHZJpu3wiW0dDIgsbvLsDvfVecQfvDy33W06dkZxLTJ3/3DPosDNLwk3vWX1
J7eZhIX9c+n7aXM13FkUGxqL9ztyFDYuwA7isbufp8zFORdh5sv35IEtA+ort71+
6vIk05mHvSv2Pd3xAGe1NHC+3kHuMEAKyjZ4l0dYxjfzxJu8FEN/uYGmrZwdUGra
ttL4i0xA7UBlT1yPfiAdvYv6qq+qktxOQWCFBUS1h2aP8Qd9iMWIn8K6siz27iOQ
OQ4DFeJrW6fv+paKvH8P1nqdUs67cY++6hKkGcsUD4Hv0l5hcxuDRrQqfuEpP6+o
VM9+zIRVNu4GwW/90VFh5RTg1Cv2sXROcDmQC8NFdJ/vUMMl+RUuvFepipIxaH0U
e+px113TqtBDtnEMHgC2f3lqlpnL8c/SjBs1FpL2UjsJJ+Nf4StdhwHDwqxTo7cI
8ETXLQ0hAnKg+7XGIkd0HQfazTA4ne0CGBzphc9fvnzKy00phwgIdB0ZKxCwrIub
I8UUhGtzN9OMDomm1lN9IlbfGvcIOVKEpGtTLN97wBlBBNeIzfgEBqKtCTTxpI/6
zxuld88Mg7E0etwSxk3hrLOs9bB43KuELacPVpBKiypIR519TmfJ5dc9Rkc3LFF/
A7WAStLdvgsG2OBjhK1WUIT1rC15cFGb7OMaDSZb9r9IV05tNL0c676K2F+IiPtT
7Rn86MzvA/HRGXbDA5gHXE9AkoXTmCE125BhyIitWD28ESaavb6N4mGFLkaEqC3s
yxlo6qHttrdbLQY9RfrHO2mnVmVEOzMvCTlDQCaHXmCzx4+CPy2gFDnxVGyK0cXC
V8XHrIJxn9CpJ4nKNAjEB45XaVj6j6tg9YTlCWXSidrY4xt7++WobHfCKDknGpVT
VGpQwHashgZ9T3WqFImb+tTeAxwqVw1pPi8KYzDV/cvgPHoRbeZ5616bxikKO3s7
7DCXkg9Xuc76/thhJAypat/BiiFVMQR414piDlovsYGLszzqBNOwHV15S86/m6Yr
oTT+6v1D5iup8Ho05uP383cMFpbyuzqo/8Vd4d/VwrWQxf11/bFy5wJPQVCvuXcU
grHHYTP3QVGqjMB4s1ze1voe2cnO2ksKRK5e82XyPobcqknye17Pnxtxl3hBJRcv
mvH/L3R8YZJwto4psykxMhD5KuaZ4Chvsi3ziyoJLghePo5C+1i5zSBqRQmdkyR/
MztXXNFupaF9P6KLwakwvJll7Ad1X6i4OM24qNyVbvS/a1EKf+AlT8Dz5EPnmZ/o
vqbMoME2Avww9CqqzMpBrnLxSv4q19b0izk/SDBwlA94Ltez+m+Xvbj1D3cF8Di5
6vkzi3YyvlaslxJP/qEx4pbWiJOw/hnAmqGMs1x+W6TfljKeaGr+vALkB/399e6I
cAUBossyLoXoMgO+Iwb5LCg5v/RWmyhJhAmkMTMasbRnbVO5yerrW70o++cC1Vgw
GMce73KNadJE/vZKKttm1GSJzi7NFw77na+/GIaaO/FTk+YTUf80Ay8DXpJ1eofY
25mWm0uKBNxBrrYeTJVVGJuTiKJ6npi7V97DovqOIVYltVxUYoeVt313wcjyFzya
GchtYXORwRMdedHN+wzEaX/3bc8bs+/A5UjsxHuzTGAo/n6wuIJRiFdyD/iE9X9v
EGf9/3psnX52J4LcIvunEgkTyb084EdXF6Ao3xZudZ5nsviFyOCMiKg7vRRrNiBy
IFdcIaTMkCuEOJ5r+zCjbVVfg26xzgITgITCpJKzNvn+0beBmxxKxqyxCvxriSOc
z1r9vUBrmtb7ZjGbfV98rcLQeS2YS0rcZoHK9fVGucHa7jsEKUgusu3b4TtYaAD+
qpRC8xJdmL9MSWAUSy3ykTbAXMZJMod2MTVG5vgfQjW0he7bL3mAzpa2tITT3W0g
9QhFD8lCClSw1Qw3EX26UJwVwgURRvNh3RCxJ4I0PJwpxmgk8pwN6CytP/GooL11
X+gPKOFXzAs0z+xwtMbDix5X699up3i1NxwRkxsLvRblSlFYYaSd5J9WMHsowy4l
anvUQQdqJKHovm/NZmzXJPl3NoJMqnxKPSbvUXp/VBwdTEM8rc9nvvNbM/b6UiJr
A/ao0sPrCusXcacjOSkUJ5IzaLmRofFUOhNnuSoaeGtSdxcEZZfcIGnJg7b1V0qK
m5TGyRV0jbcltLqXvPloW0vKPIevTXP2ilH6VBJRVqYezVlkgVSz79H5wiTQD/TV
n9c8lG3VEV895Gz7fzW8d1MrXUkvZz664m5EVAWk2F/vSUBZtxqkhthQ+8n7jjif
649JBCPcNpTdRCEKHe7LPKcCyZ8HL2tiKgXC17NTHN0oSxEXBYX0jv/TQ7KCo4yL
Z3Ss/EXLkH46vLU8kj2spKwq6kmHS1nzl9VY3S2CUs0sILvchuGROoJqA0bc1gyL
GYxEYqbPvBJtthflGnEbm0i6jW26lumcZb0ErD4LN1Xonls0GxADWv/f2GF2wZlL
/ykPaE4aAIgq6rLszAoxZtOeL//YEa0y8VSFe4SInw8FB4oQ10VlM+BWUhE8pYYQ
tk4RuFIt6UC4+LpQ8tr0Lmk1OpM5Ss+reW2AhYCKol5M0HIik8gMtY+5EnHi4B+T
4K26Eu/QmbVEhodArsMt1OrEvLDImSi4AzdJFO3VFgnddWPj1phR6oLidjojJtoN
xOklm5Z/rDw3+Y6KvxN0HCTI0BhhXAy64CMzSxAcn+2q1hcBfGKHn+sKpBWjMc1o
uQslEJqhQ95lWjqYiBXddouw3CBSVpA8pWsWEkjm9A5ILwTvXms/dF4lb73kwWIE
ewGFBA2h7PMsrxFbtigV1kdpJXa2jtyPEtsp6MIREUHYVmHrLXdzF9VicwJ5RDAY
5cS0olOni8cHipBfqAagE5csD4omphUvWtx8+/7WIK5pg8hAXVEt1kCXNIsypvnk
3TFeDv6X+daioQSV42brXSeprMlzj8cC5Y5L4CQFJoEyJhVDT6P3NpTVwYe16H8o
EKoweSfEad1cLRi7qBG5uOmRyadknOEpzlk20UMkZQ5aF2IFnZ0t2zLWxtTaLPby
HA1ca4yCySgz8llye4kdqESRNWWOkZr3VeYH/cHOwC4YYL26l0tdw/i5nM4tL6X0
yIqiK7nlo60JTtYv4OJ6aUHTcPFWMTP+h6ILXve0k5O/MBz5VFimGwpSj5A4DDH3
7WqqlvlsmGax6ce9/MO+LzhMHYpL7oHgLS5qUSsV0coH452jssLp7XIbI5RD8sLy
RRq45YMR2dNIPZj8uEMyDHoX0Rnjt7AlraqJRTefXiFWBrukM21zVG31+twzA23a
rz0GoxwafDIfINGNLN/Nyqx654oxpkykhixtZ/9yQ2hs04bQrmxhYRdNFE+vRYYh
XPdXu0ToEfBX1nQDbAiLH8su0SAUkQoGIi/7oqExVBwaWGVJjtWdkk59yks1uxjd
z0QXyUl91NyMJhmauy4nlAC3Yx+ygGosQYyuxGEgnVYVtZu1YCycUU+CgQmChDK6
RI8mR+f9adoRef/jg0+rhWvVqD8S7du5eM6SQYv6AUbu5K/8CqUI7wJVFH8XaGWA
s5jRGQzfJwpoMefqQe7NeXZ/MC4ONr7z5AQovJ8P3BKdPhoxfNGDYQOoWiKyKgUi
3URse2zzmGm4hTVd0QDHzn4sFvkx9oRdP4+f2V6kJD7sQ1ARZ2KZBS8mOv1ohQnq
dA0u4NgJsve3bqn2Pqv8COal2b3tJI3WrJzp68pQucVHvqlUYMDn4ALQCDe9IQUR
2WScgrVarxbe+/C5c/F+YrmOYLE0GrZRX3G8OaKjnaw+AZCEskjtW49Im5Km21ul
XDzQvs/K7ssuTnyS5CNASrjtMSFARfUrWU+4m5YrAD5v46GbbqRcvNqcXMskykNw
i/Cl8Nga4mAn6SbSHKRYVksLqYXQsFf7QwTKRjIQZ20je1qwq5XiqBt2nIFsNYR0
QMy3p31ei3qu/oXinP8IwOQR+lttrr2nJ1KGlZBYfWyTe5I0352Z9pWFIb7CD8Bw
b11z+dUF6hakdWtTOntbo40HvSfE0ywiWB9DFH0pBxPLI8No1ntwUz0bARirMA7B
+16KjxvslsnY99alyBv0t2WfmyhNvNlg3DZhs2wdGfIONPgpzQLB3WiHEp52Gw/U
dmecYtHMoVhsQCNNiAhcx577N1xWT0/W12j8ibIuxGdvHUUIHtWQtn1BB10M1dWO
T9IoGHKPi7DxxZfEeOQCHrMg3eyAxmBibstrGdDRg8gzXUb1PIG++FjVI0tbqrtl
yRCcRU4iYyjxPu+EHPB0qW00GEFbesZvgUtWRmFdfWNzOkguQUjPI80YpeuAcxgX
KcySICzJG2TE8TdAJlv7ZH+qSyvHNtkxJH16XMvdolHwEql2FljFURzAqS+jbo51
4MXLPBENID/Lb7QoftNvc0vdXCds3ZmZgGko6Na3sJn9msgAYKVckQUqQMUsBa2T
ttwPrD35ubBRZORRFWLn/Ety156A/jCj5LEORHbTAoS7gDLf2UiRv9VOHz2gfLFO
pO6xwofsj6qM3j7IP/8EeoxesZukcQ2uXo1nMFMZ4iygMRbD7DPZI/SkiR/I4HNN
t8h25iiS7UVd36dF9oWlkqvrRyg9oLC6ycdKiVJdhPeLGLw/QYSJnbybFO+h9nmO
vEwxGGatEFChB/KpdLDblXi4JLUZntEtcLH2BdPXS43bNLVQ5yp+2Kb4AGLmgU4p
OhMxhZ+lpumnoSn4dunfFT51kd3zjQcV9PHkGlOKXPK2HOUiJf7tl0oA0AfPSFq9
80V28ki8DZEAttbeq3g3ehNzGwLdS0z1Sap/U4Nsq5tOeke9pHPpdUx+7ZyD1A+y
kG1i2CdGlECw1AwG7P9PXTbDsEo6s2Baowi+Nx+B6xjBGpCWGrqAgC348YsQDFSJ
T3LTPRN0PC3j0lQYRaV1EOx9WON/vIVpAYCQHuBTduaYgC5oMrKuGd5HVxtAy4EW
7O4HTKw0JPvAsXJqOLDQFmHjfMkVc9qMeozjreudcJ7MUlJf4KBE1WU3oeS/NhFV
NOPwMRu4NoyKKZpdFBWpXmeZvDyUPK2JLZNhXimCbdJ1nf3v35khERLsqNFcxj8f
ITfLayI2+XXoKJAEd0mXOH17JDeYwV+AFXm4krG/Hk859Gd5/xal9WwzBzMgeAuu
odtRSbladHWLJzGGeR0RnGUCEOrWYbvQMSAMyrXUHiRgYlofJTyd5IN8ilGpw4DE
zEwtk5HTPHA+jerXQ7PXWF98/piFFtoaktKBiPDSyJ3zdK/PoWz5FzD/L9ZoDBD5
zj37Vb1Z0NquSBtJ3u+E7dCOG8udjebbVF7nwwijB/oJtAu2ub1U/f2/VctAFPPZ
Htw6ICWP3CBovlkxyLpMCLYZkQPGAZh16e+u2z23IU66kNsnZnU3/hwBGXQzeKPF
jYtpOQliMvfIEVhYNjluxHzapFZ14IV9a1HoR0HbkIrHLSm4aDImlcdnADINyCkf
lSN/QMrhEzF4aaAWRMoO0JtXnMvwtMDCZq8nMZUfJU1ZjZwBNf2jHlq2z4/7pWc7
5SjS3BTRiPjmk+gQ0tq4XsdbR9AREzZtu1VwgvmpuBo1sLg6HTCeOWNGi0EcEdFs
2EbbN8Y8iMj9H2PZf4AqHpNuBBqW2vPDge/Zia10KYQySk8D4ELy+hs2OSUCiNP+
n0kxshhwtiLHX88ceFol7Kz/tiFTdwqd41oCER8GRJ+YNp2vZUMTgXxQytd3vOOb
zUFwmG14YG4jQF9s9VWj0CnZN76w4OKVZWA76sJdEDPHsAzAP+WxCI6hG0dxVgAH
/CqnZAAtbSaWDcpguIdDQXYBYoLPGkz4jJNNVQhSYXBZvjzhrcB0VWHkCPC21KyV
ZQRLqNz9cuxh6VyMlzayRNKxqgwtV/tcTBmWDekPkb7kbD7/HzCKBfyN7ryxh+Nm
8AqIZXgY2taXWII6w9bdu9qxGxHNMNkYu6JlFJWhCIpsz8ZIk0ioL75xs9LISC4M
XoZkUHo1InLxuo6wDELg5ody5NOCEUZ5AhZUk8yDEXHL3Lh8o0lRbM9KYh868EcC
I4Fop0NPrtwILM88gPZiRt2Hiqblt5q93IP6rDxMYtYP47ULDiuQQgPdH8Mz4Kwp
5Ev8mTb1Sifpkl4JYr3xRw2dg7dy5wgC2OBRvINy1Z2uL4lozSlKZsikUAu1pQou
V+QQudEHnRXtk/LuCjDnRwy7QFzb5lz9odG9HX6SEv4QTUHYPBWYEx6nUQGLJVpf
N5Rw1vLkrqOPTVaZ7IHkacRX9v/TGltAF5GXx3gctM2zibwtn/5ktDIfflhLLDid
IHkXNZKye3hiDQ+ND9hwkKOKy+BxcCeiokLQ7DatYHAZNU16UnOkTRwYjDw+Qc1b
EMkDPns1dLmGh/8Fybgg6IfyZYkE9vYTeGtHEUufX+4Fx3BXHvjIxL9XSbODKfbI
LbSawMnY7ESoJRiF9smeME9Qxco31oUg1MkzhAWfwEVVIZ+spK0RsoW++1BUV0Rm
v3qgU2WNYcQNTMGoHIp6Ivv+mFhLZFu7yziMY51Q0Oe6M43lQWezweIihsJk5cRU
QC6dUhZWvDkHpowoNwegZ8/ubHWLPirUbBM9QN0GUH1jV0R9q+Ah1wLec+6vrJbO
3YdJP+zhZUAbnVqsua2YiyIRAbQzfg38FGu59NXmmYan/iYv82eJENuGfG2mE/5M
A7FMr7QRiAAWE1AFC6Saq1XAqtS8oO4Wpkz0GXVhtUezM8X9ipaQjXVZb2KZ4oUw
TRsRnd1GRjGcI5810EVVZMkQQsexIOZspdd8/vlZhaRp7IwwX0QxRoQ6cmml30U8
9IMdnyIg8RMI+yMh3179txPQeEuYSbx50YBK0H4eYgRvZe0DBh8oQnwzIcFbOnwX
RrbsX/MEz3Lf+czyhek4Ap8cew3RwdCzGnIVjX9H/d7M7mf7ejgKmUXlfKx2h2JT
vh8PEUs375Xii84U6Ounc9ED9IDXJw7Xtgz0lxLmpqyT6GkKLey5uywZbLF6704C
sMaR6Hl0FQRmtXCf3yuG3qwajkbp9nVXmyzbaCNmi1xuk1hkdVorIXzD9l9KddmP
nxKYtG4UOlLGBEwiDJyblFIBHcL0wgMp3n6R+Z4ySjDQk0AYjclWkoyYoOOBrlBR
J0lQBxqOuRyNZrej1c7JpvX7VLchYD/133YMilClRvouNn9FW+HmLOuZm6HgbWCy
ntlFrkDvmG7GCcPYJywJoyakdLQ8eWscAWvs1gW/QrzKSOubqLlJm+rhW0NDZIBK
8pidj9Vf90u+NkB9DC5vgwJPlwHhbS6IbpmnlR8OMhZ/PnWa+373fMw8BM4kAh8h
fvhRy+2QHM59UziYsjaMoYYW+K+ePofFgJonSx+zLMiJE1MR3COknDwaJf6xvM6+
xow3tZeCRentn61Les4nkRKChiYQRmn/h9OLuP01U/w0Uly25oZFNkZZluzCvbce
CtMbQNJN6T3+0b5cd4wGJphhngN80MNtmm9FtZoe3VoGlq3+4DNUamXmMz3fVqAK
HGrxpoUfaZzTezkxLAPsutqyRnr47+jKdtp3/bo9qYFsH5Dct11BAiesr6WvngvQ
BzQTKSd5BZc5hNYBpEcR+Ur3lIzgClCujzYxfY8YKpJNaFYO1JMiHL0NrNf97bRM
kzZkBgRMwzMXTk+XzObdJP7pN5P/su5K5eVJDL4llsQmwoWnSogyRIKokeSEx8AF
5UqCY5rQfUeqbCKwMdPCSJYhb/g1QYrHDkyhccMCgwGFs7HFsP7luhl9yS5ZL8ed
fzrgO9Z+GbvLiwP6L8qoE7dc1M2MsLRHPPqHwT0CrG+nOqZ/80VAvlXPvEscI98p
4QTOheaAKmz3cWr9irZOZtHAHj/uqW4lBDe4RCCPBbo2bseNh4+9i/KZ6BajigMl
iSto9KmJh4FI4EYtXV+vKEeNLiSnW+pacncUMRYgXnzRc1fSUx2jksv58BZX33vr
TzZd3FcTNmo3BXyFxecYZKUO4hDZOwQDE9CT6U7GFZ8QnpiUsqTpAq+FPX7cngeS
rq0s9VHGkYDY3Pjd5jE4gSfBKrfpsBrx6IW3PERCRnEb2SkMJCVh2wBpsnjzENDa
Tb5ZW9Hxrgh9iYF2tM7U4s25145RgdDx/MyXWiZMAycGGkwwFfekmAvrgKy8+/az
v5TgXiJ007y0FVerd+ZX7zGOhvIG7STAmVeUyCy7Lbc5PYxYNARqLJMdBqmN5xhD
F1w9TGmQ75bxhlhPmvN5hEDafDdVkiUURYMtz2y6rP6ylHwRTmSh4KO2BbSkACDb
AUGc9t6E0vXD1Z4JckrJSm8ibsgsdmkGAP0B1VaAOIrj0C85DILXpqfGwjeH0GCN
vLZ0wT7BwkPfNAX5QL6uVBawyNf8EbKqSlSdMnfrqTzBdYEX3hhiG1k6t4IAPvcs
uhfQGxzn7g0vcVQcWMvbUvdeWLHdkY2RgISqUOhPxKtAeglCbOTSFK+NMdrBkMGA
kY8yyWgBRp4vH3IBvx5CPh+PEaUJZF8X3ZWxioawd3ohWd9CrLo2OQKK4ONN67Sf
VWAW8/YPZ0jsy9D6DhCFVaCjQ86HecgELgK8M4xc3O10/bGv4ipZ4zikmjyb/EFn
bVlotCm0Vze0Np8KShBkhZhdrOcRnZgruv3D/38HvgZNvFiQhz0njrSCEErDiirL
oizHQmCEyKiDzAP50Htpl5LCP43ysCjMcJrdmFYfH0wZCNZxkfyAsjE2nfIbR/4f
3GgAUQu2a7rlkgaMvne6F2AMEVLyzvTr7dljUmJWs7sx8easD0QUqTxC0CSV/BJH
Xvjcn1BY8bl7hl57UR35FK1O9TKtS7LrA35MIGskfGXodo1otypDOzjWSRqBkQM4
nPD7stICAm/C0P9ftcCG4ZQ928lb/aAtJLiwNgRsXRD0Bqpu8sMGuUoQ0/gykR/1
HyszdEdvq7HTR6TJD7Cr48Btt7ElDK8JWblPY07OklHYAubfUdv3VlKIuJj5Wrsb
TKdVRmofpfl5qdDN1qb+rKLYiosKPX0NWPOoIgRNtyXFF7BnrPyBuZ9y5UajW881
5PPM7i11BrkooqtU7+UgKkCbTL3z03BcCnlGNHgupq9SNc/M8UXae92JDT7arYyz
0O9bASd3nfopKU1a5+Wp9pFtxdJyhW3jYIQrnuCT/MK+hEht5DPYXjyyE39GIU04
u4HZopVSkIp8bfVcaccwTEQ8IHzYtRdvDu1K2bMJWE3Wj55qPLB53nG/AcjaJV46
0nYYnXqCZXIEoDp2m9xBu5oqT66RofDmz2t8dJZnvfGWRN4P6V6l+kRiMPPgUhwH
xTgDomGTHCm4NcQ5tl5woLeQ3K/x1KykAoexm/Zizw1Q1tGPkrskWU/ajrZ1laBB
Z6hen2MDJk83tyk6EzqA5ggTxyUmEhuLJ6YaAuUOFWm1m1ceVUiOTmMfmFPJhlpK
mL04MbRGrPp7JJdi4AU5AbuFP6dJ8k4BStFeO1eMh6i17w/ww06kJcdYl+njK6/l
eHx/g4GIbCzRL3y9y+8vrEU+OdU18+0IuZ1oYHfjMNY+/qYUHdjFLKmxhe/nIOwP
OMngFSgN8Iw1zmmre3LqKxI2F5KrwK0a3K/v5imDpIJOBnCSxdOI5SlKBNcg4GjU
KzyRJ+uPIR2kUPRkk2cYjR0R7HPUzhDoR+ZBn7QAs19tHdoUa1wGpWGdvj9T702K
khdj2fnYm+p9ZgsLz0qjTnefzNxk0ZyY/CuyhqnEpW+hpq0xfoxVi4MItOnlvT5U
0geOWCudSdg2e80fNzJ1BLbw2u/kdn4HkDLRRQ4yjOOfCpuFllgD6kDyoeWTxP3c
v+gYJJf78fntn49cs07FuelQEitwaE4+U4f7SCjok3/b9+T8wjH/gziAttAksnln
Ac1I6AO0qLMInp9qWfSg9SvBU66wu8Qlrr2joUmxStCgvqtV7cxT0aMj1KKNK4mz
hzngRXz/yLER3pqkYmHg+EXnADfM4jMZlYC7B2aK8gn8+g8XwacdPNVWagLtXkhr
ffsxGKXAR2kDX8q9dP8C98TNjSnbv+lI4jTxFvaJ8WqiliKjLi4ImhKlw+LTOBGA
ERxklOraopAzBsuMrXZ9qRbH7fPvKN3Ae3rifEFD7+DE2zeXQgUPn7LQc1GQ+Sfx
ToS5ZEMy/O8gopONf2FyBVk3QYxvChjXygJrPawXNUSQ7I1QgrxV7OwqheGpMuHj
Dd4nVBZuCPQBQTskiYTrUKJ8IkfNCq/qYgE4sUEhvPgjHR1oX/y73t7CbTV65QyM
KMHL5bsnUkn6L85gPHHqQRImd9BOZ9rDXpf9xnD2UCGrT2+1BB49OtQPU/HhgdH4
UfUVBa0xLsTNYnHwi5XXWs853Vh1xiTXsRjbrsstQws9kTifeXGDnerXAF5w5cC2
sU0jN+sk70jtBOHHngG3P5TUTJIMQcnjaoa/RjKOARZDXKKeOLRqceHextoml+y7
LrHmgZZ79ZqevUBvEhWmBAbeCbOE0gWwDo8KzOqDMrVHtGGj9XrxoaLTgJplUonT
/j240tOwO9gfRT42Z7svOpW6QjzRsxcWVEOUubokUbAYU7dbE+GQVmuheKIZUJvB
Bb5c6XWBPgZdaV+y37QHdXZ40fOuB573TrzixqRDIySsiQAQTgKhntcQxbt6T1fQ
fuiu8wvTMIlxhLvx5RATdxIa7/tva0/FK727BCJcB3axTxMj6w609n5GSJClAFYB
SpucS7yQUPfstxpf2p8eiERfm1YrUr6v/2woPlSb4AXISB9SiOx7FPDxmP3ceNqT
dn350bptrUhNoPcYzRvHPNapFvxT0UehEKlXz0ba2BViAp0CXPVBFeVpLO8B3Rep
ndG0w7zfXWiBxmGzyc2KZrCOkB6dWSZrOYb0pFV03Jj73l6mjBjFqIZojP4QYXON
AXgLBJisi9S5Zw3uVyEojH9AW+vMREXASdRJwIEvFLtJwzZJLX03mj89rSgcG6CQ
muvqDI/K1pg2x1YM29qV5ku87IXriVkUkOcy16hJRQaoSNn9wxMpjMntree6vdvT
dXjijs3OUqSFvgw9H7KfMijnbL3PLu7DRZEhf4yb2xFMJFwNcNTRVI+qQDZpOnxW
lBjvsYygtblZbzncn+zkJfdCbOAZo6XXCqtbTmZBN2Zu+HyXsNbn3Zd0OgY01HJT
a/J5757Y9B6yikjuXxlCedblxCU/lhWpf4p/Soc4XAGHdfz5vyfHN990GR1DYkGM
BbmZHuMgY9ig3+yxGcINPeI4ITu10zzkl/LGCwlxJOvvErzGuC5tpIUJotSzG3x4
1xGyhOc8mDHmL9hRoI9LHkILl0/CSKwTik8EqQ6TzzivgfdGH74U9dweOug11Yib
F2RGzHprSBsIBhttFdMnumHTGGK1chzKfMkws6G9DFS42lhUAXiG2btlZUkkziMs
BUmj7fAmRXDv666WL7N3Y2hPgTWf+LEnjQC5fU2zLiFYMTgTjGuQdghRgN35/Bpj
QMRRwVhkprSqH/FMugD38MICRI89eubX2H8kIgUdpm7cTbLBQLCVIpw2tQ8Cu+JI
q2yvtuct0PMVSBUkdYwiFj/wwOx7C//tVBDzriy7TOkcBTjqPLHYT8PKBbjNyebV
vTH85UcPx0eTCJIIH47s0IzXR30aP8D11rBr8KzHJFPZNpYiQSSWl71KYayofq5G
u/QastnLooOoQuiw2ZYMaK338gfeyc+VolZipY0A+wmF8LYyvURDmLnL4oHDW820
dPuLCp7a85Z55pTbvDVN3ozTOT7X5xjtUgaoy3zDOH5HstmEVxtNy9jHiKkfJ4a1
5W9xPAg/lU9lMdEGcEjoH1FOissSNTAS4zj2dv94ZhEpTlzZ1WnC5S8ILWDhfLHi
3kxP/OncO8X1xbe6ORSfz4PSvI7XuYiyPJxxXiQ2x8yGC3lVYvNbC86+M4WwIpnh
lSlb0GZsijuBTur1nShVkXTOwCGZJJvZkAhedhzuXXILxcpTq4ajsD8nHKQDoutV
gPMKVuypqW/UTFFaw5Bk/Y4PmW9Qx5UmTAS2WhjgB0t9kDypOZrEBA7HqKuXAHaE
UitQlvzAizMVfJrx05k6+q5pQS4ePQwwYvJFGEtQSmSyRM8haAMzCAQciPirPRPj
6hYKrHRK7HpFdijV9kX7Au1ARFH4/Ya1r37BA2vGlOkN1CaM8shbRRWkgPO5VXaM
7kFps/Zj3uwxdVCHVoTFqkopQaKR+No4kuoWSVK8B+sBnALZ4c4JtihHrfPgBnT3
n83amnJ+HRdvpBALSpIuOqni0pcimPJJKska7FnEKUlsBlQ2YW2CtwWn/u7e+nYS
0KjUEUOZqj+c+zZEqXFR5y73/dgB3NlK/pXXpTHcH03S7SeTODtXLtkxerPJ4NQz
P13t0mcIGrB86uqiL2NhiqMk5hhP5YhuUMoZ0lpxO5VTZLHEGN4TwH2q+VWc9aIa
24aSsth7wCTuV5/Gek6DGNAlae/kNCwtokKLlwqYF7+MwcDW96uAPRa/CxCIY6ir
UIWgDqVDg+BUGxbBsaXSKGlljz3li6iRcYQCYqCv8J/2yFi7y+VfIlTDHDd1fRQi
rQibKLAkBWGvKOpdYfJ4sc+IbziyCfo9xxpFpx61YglAoo0rIuDby6YmA2HOj+i7
nOJTcuR74HS93X4sNsIuDjTYsJDhGOwAOANIwxAQbTs6w9eUDoIv0J1xcxS4YcFv
u7BgCbgEkNmjHoTp6L0JBdXBl11X94yXuL+KKYB/kBVHvMN/Npy7FB0aQf9XQ76H
EhuzH/Q+++QI/FE+Y0FNcq81wdHW96wvcMfm3DGDKN89x53dbpscpgeM9Z0nQMJd
bu2/PWAqpSNNhZSrszQmdUHxuGF6bdg8aSLlXZhCNQGV16ZirFdlWEu94yk/bTsr
OKjQbSdrdnWq6g7sk+SEZ5tgrhYjq0mzJ9XwJKxW+s5owVWav6lF9h5c/xhk8/Oj
EbMqsclcjjp2XssQl2D5phYQap1o0itCWawih7JeojGX8GvaDJa08CyjWtOpiJM2
EsL03gB9fhSVz7hLl8f+t3tkvUEIqPGgOoWe8Nz74a0TaLy7agf26GXcfKLkOtnr
eZ3tjtSB0ZoQztgdrkdhv1y2FjZthhcgopG0/uWCD2XoJTHFh+ldJ905xB8Q09Ue
ESOVCGKI5HJKe938cW/S1ioOH48s14xJSFZ+b6Y0duEF1REim5zuMBPGDer78EKM
u39XKWuoj7A8ImZhvGDvUEmT3r1osoU4S6rdtHCQ3u7DZdPzH1g/PapvEmsWAF7Z
ENj9uCj26sSkiykhH7NXS/MoNRofiSOGrP3ZVSDRj64JSEYMjOphAV8C+rQV+dlQ
1UtdTiEqk0jyYZXvwr8hu17YsElPXToixmGYjnCnX+pxdea6Br+XgchPfhNsglAm
C4rwll9H3gTLNC+dsUq7qxoSUjbI5RhC0Jdc/Da81VN7MAC2NASqVKu2ijkZImas
MXXPFTMuD8HfNLk+J+PzN/XW4USBAB+jG63sNuVIzas3qGOWEP+35oGp0aqCzFWk
UyTwQ+X6yEvXoNG78XYVazmKwMoxJdXbl9WTDkc0WxBiiBYCqVhWipZoEzvuQ7R2
J7zlKpILfohMg1LtRX1+cMpJ//4ojErRDSYKcRZEBhR3w0qaRrobdYXk5GlaX081
Ti5E2UtuYgbryvOxIHhbh18MBko1c1DaLNLi4jb6SeZVzuUzSknGvAS0Eob0y8ho
zJxbtfjoJXXV9ORmAwaOzJxFfiLZQz0mYd8fIHsihSDg3Z+LvOKo3c4thEPTcVdn
cZrqmuYWcTitgbrCUqL9C9hU1nzHyVUwvRw0RjQvWLC/DqBc7Boz/OOO28icBDFr
Yq2TujIDgiwfGkK/S8oQX2Bk/LfaUG2JllS4pSrUa8vE1VS59pWImtRoOq6jz3/f
DwMriuTEmGsfdk9tjL9H6KvqtJUBynC3nxKLyZCqg2jDLYD9QdlsHuTXzcyQ9g/D
X9LGFbKIhk+rbhDNbwat59PdJyHiUvtzJL1BjMwkRdzF1xTEJEHgYY02SduR9N1y
1TYOR78TMBn/VPy1oNUGdzL8qB94bRTuxoHPdfs9L4dJ1w+jfwrRwkWAulpvL1GC
8h8RXxFUxNnKxckz3PmVG+z6BxOyavmWHVYptysX1rrrmmYkmS934xStP6gXAJOL
ZkXVd3EuIDOUX80SeLm1wyggaf77apDl3ElwU4zkZdyPlNALoShrQUxzDiv9a+gI
FOYFAtht8rMuVfnqXwdCwNwwwz26EppBb2+H97bwIrO/3vG+L9WsjQJwbay2UOD9
FpdSmuw9q+Igc3ylVBLlX/FHAo6SIy89uOHuMSrgYXZxy0q/CwZQK4INFAaz20qv
C9UJKxTksv+sS2inW1tcFbn2u0KiIXLzuN7l9p/oTMQRida1Rzpro7p6n45ONsHs
JX+7SrJBcZ66KIvbh6PQ45Q68fOReV9aQQOLM9j7/W20f+KmKJ0O85nFwZFEmwaI
iCPiRK9IeGovpOq5ud1BEGaZlLG51Bavxa3ZPwe/oqNvKGkDA2mP5mpcpd023ER0
hvWHojJVOSlgmYPVHVtrKLXybM2b+xaasj7NUPnEI5pmb7wDdOyHSOjgYNyCBszo
D15wfUQgFPWSlflwR5UGhHuBiQfBi/RR51g1+TS5C/SzGPZOWIOAEDECkK4q6TfE
vsVxn8NWTb7wOz/LxMd6kII7BWLYM8n9w3B5XjVy32uj5CIzgamtNbwYUiZsj2SQ
WuZKtNSGWnp0f00EHEGEXnKSjS7LeBSstYY2fRFB/rxad5CEnyIex8e7auEFfAWP
/qYHSpSKbXqj75Pv3UtgCipB+T5jOREuqh9r7chXSAB5HObh237YmE50JHxtfAOy
ZgU52Fr75g8YrHVUDND0jRdmeWPi9Ih9EiEs9nTs0bVZAsBlebDRlt7IzOCZpT8H
esq/KTNq6xk6sHWSN0YnVE7Z22HdihKUXDR/GQHk56QhDsL1EPYChNOzbxuSd2JB
xd74yhfE0rfkTV/Js+JeKwxG4XCysOK5j9ERuOwdeblVgef89Klu7/zIJtzuEHgD
E2EEez2fw/QGp0JpnVNvwDuUKVChzdZDO1me5cMaiMqlwFJEbsts3MAs8bJaHkGa
GUbF+1eJS/oM4FDUrnYYlyrKguTA3J/aA8YItvWsIjSkzo94IcTBpn8elfxS6GZg
rOY/G1D4dU9tvrAL03r5bfCEMQLzRn4lVDqtQM7qyc32+nXlxRsyecste1bBzGgu
rNhaFLj//SFTeDCXoehUQXTlEHbvR4dHuGHX3LzPe/L9EqbLgJ8nRHqx94oEzhFY
K+hy/yEz1+jzm7cGNGxNxwhrpMdFTjEcX8Bj9mTW0r9hQVYp6PWGkF5Zkq1HHYQ0
9AZPFQYnp312bfYzXYciRnjPUHoqrUmurKXNfRq8qLAHC6qn5naQfK0vryR2QrSe
w1QVbEUW63ARqiwaC1OJHcwUGY9gHUazI1YyjisFuukno/4w2RvPoTkty8/w0AXf
I20J6GFC+KEPuJKd8vQOJdWjtagLVKNjKYjRg2VSxC1C3Wc7j283Z5sZj/J6rqzo
vnsx/1v0+YMPaZz8ZtE3azGCN3ZVo5BGbAWumjoSoXW2IlvADu4fEhkP7UCvWnL7
S5CpbNrSO0+JLL9UM2z462OS3PQgdZfc3AK6a9ohL4U9UKShTbI6jfdfvSRZPBJc
iBZb+q+ut6uoZ0bnApbPTgpmOPC9RiqCZ5okKcHgLnGP5uw+lWUH0fvQZcJE/3IQ
QJ5pbeDcHt34JzJJ1qmvJU8yTNqLPbjHN1X+FGUpvgd4vzSqI+hFyjko/nI29pDT
ilCh5glGMr46Z6epPc24qX/HKZM/9HCLaX7QaMsLn3DWs14nBweNNQJEKKU+GnsV
iTYORlf5R4fVN4kLp5/ZvTDmdS4e+W+z6xTB983nGpnn59N2PhddR3KrAaS/wK50
NZeLCCwJETNVu6a5zUpYvpuwBZkIlma3Zm1hDGlMyZwsAnBslZds63HTGyIAyr/v
CWOca0ch92CT2+3VAfCsc8J8wbPo5JeMFVWGDvu1FMs1FhO4qjouH4iEqKolOHWE
Yc6lVypXa/fUs00N8g5wLve79CdgfECmN9CJoc+ijdcwUNEbydc4GvfmHl2a8Eq4
9oLKNwVfZlolaP1PN5BXagxGRL6uilBoUriTmcGMpiMAnqPtX5zlC9GjgAzWwsC0
JAM7N6yHo+LmaNy3tBo7oOuseT9ZlPDTuf8c0merGEBjpozeltZW3QcLMPis8D6a
+Mj+b/2HdqZMoo+TKhNbJkv6x160TzJ59u5xFbmn39N8BNT47E9v7tuNXsOPVFJA
Ro9yC2uJODZy+EZT1exu0ZGQVvddc4GLbVjVSVSbKs5cSRxhnF9s3Tq1jnAx6/CD
k5J+r+e//1QylC8+0NojApmvjNzlmZs1lLqxUi4XpMzPo7ky54ON0ToheS8LGzeE
81YT8QLDeZdlP/woTm7kvDvN6B1xMHPMZ+Y5aB7pHEFoKRxpmxsZ0Voa0drXYurY
6nAvudNbhcBLJ0QA6Wdk4nxHgmo2ta4AKRc5N/pU0Vs93bbDsZtj89L+Hz87O459
od3CHFqQtT08xhPj5iuAvDjkmEkT+qqJKN+Uqva1/E5Eh2v+Ra3x+5AhcrjZYowa
Uj7IZdc7n8FhjAPX2zNcJGRo4K5ljROQpMY5dRjWCdo0BxXSqU0My8GekFZLGKc7
NeM4bzrIZYiaJToENO1EnR4GzzyajnScRP/kHRMibZUQ/COFtXyyxe1RJTfN5UqI
45rVgXVuQC3d+4gLoIQ6nYw8PJRfE5Ddfb7oOIoTlybuU4fYlQMJhhCIHWJ2u5Qn
4gQmqWzmk1H+MIryGwEIPricB1huDfGw8AvcEclQXWLGfn0A7PjlyfWs9XcZYOyX
OVNHj7ooYyHj+cVmT1X9TujSEiY8IxT+7rHHSu4BgHVPKAvE6R8Nw3tTvZ8O2v9M
D9Z8AvOLo0eyMz7jamSxxj6gfffQE6Fjo1j1j3o1ecfYFD36t5CWmYeRpdQBjyZO
+YVWN2YeyoCKV0HIgdNpaJ3+euoCcRaOVi9YX8Obz86X//qD8kUY/hu0O46BscPs
4QXrUDCVw6c/0TB8JHbkbqqDnRNFV3Zr+jH67hsPcTv+bXAIn6FE5kAK6+2Krq6c
Fmk2ShR0fkTtZ2MJUSaZawmyQXl0mZ97f9ZuNVpWTE1HnDS9mu6yDMPJgyb9zMWz
HuPOj3EikSWOJrKO0IFtxO4whhI6iTZaSPfMZ3NU+3lNUKeSymm6H0GPXi4rki5l
EmtzvazDRjfuL0veUZ7Nxw75OSRaLyhEnQLbGeeroU6WjS3a9qlroqWJ3Bo1zGha
XYDABqMT0j9hQ2WOm7hpf+VJJp6duC5x6BR+uMPb6HXnjbpDSRjJBzA1Abnf4khd
gi0uo/tnOpml3kqYsS+p/c/S+t7xOyx4Aqg5aYC7/RVuMnU9N+O/B1AAkEePVKnM
A+XBuZevaN0Sxgm9VpxKrPZ2XDVesJLe1xEAWG9gr+fb7GyxTY5VLhRW7GRWIYOp
fMU+9IwO9nmM+jOFcLxFM3QjmWy+qF9fR0sgiIIJeSeJw2zSAA7ekaoqSLdsq4ej
bTxMXiER9oceptN5XvDknSlckE36cMyF+t4UA41Rg/W06RrGXIVO2ww+IfmkhRdb
bU8X1RKlLdOz5N6SpCtvAGUBoRY4kkhNr9P3I+ukY/UOkSprHRfEdGneANY4e5S5
0QWhDvFJnj+C5Q5Jz3gs1V9ij76MDMde/oBooLLcjfwcAc80u1O/UQo69e5ZfbLv
rzZLADpQTwY7h2LLGT0AtfhJ7wRxv5jemjTt2PORvVbRoAauHzP+hFue89UNaRGI
OdMveyz1bihNTjNFf9j2zErwIsd4z8xYBe5V0HS3aJsM99l5Ou9/kY3sTHATgL5m
pE0Sj3YZbsSLqNY8Eo3r3spsHAj0GxnAbjz8Kw5Vi83l2ZgDVtmkr9lAZE/EImj6
4KWs8T2tXC9hOzgYdFN5Gl3NB+3XPR1AU21Sst+YZVMakYHRFBFl4rK5ZZx02iDT
pHdoSJGDiPgN0rxF3AhQE5gbsOkGEbs8d6eOCALwSSShTjIF9vMZUvPlhShFJwon
iwgkkHW7+hicKS3EzoABl5Ig/L+J7tH+CeYJ0R6wedg2yiBPl3KbKzaZo6CoaEI6
RGvGOVpdHKmcHcLvJ7et0LLsjR/hdwSptSOYAyo1FutnVOS3o5j8eKhbtPoTozAG
WEl7ZVni1dI9U8lLly1wKVgUMeUluK/UVRRGLBps9V0kcQ9BfiBij6nKfdnVj+uh
GxfLTh541/ksYn8lPLFkqQst5lMDGtpP8+E+f3VaDmyO7yXSVuSujjhKQSAphE+y
jte6LazlvkJUKq6rsLUQKtPGuQOq9tTnia8nd4zwguOWUzEoy2BWJF4NP/SSwf9F
9I2hBCz8+kvEpUEYjOjExWrkO4vJAHD50m0qtJBOKOhne+80JatkzYr07gz8VeEP
7LbDnuF5jq3W20OCiAy0nU/pWc41ZTMDXb8XlPBwLdFGgY7gMhibd1apg3OjVjRm
B44Y88ABbQk/lkdAaHTIdaSeEDXdQpiC6RIV2wz/DGvi44wo/C7W+8Cqys3+qmrg
c3eIQdA62bPS0EMdnGvI90CxVhO35eXEZ/oIA27CkpuGZmc7HGQh6t1BWSgVt391
pY5F3kva15tn+YrX9jv0HWS6+XjXEFmRs03rpe8mXS0Qs1UliBW+lM7wywI6Mnxo
7+7jQ2GeXCy3obnNQqQ8WNZCWYvNqfrlF8fjHlwh9qQYzQmJbzXH0yBoLgTwwXh/
AH45eDxM/iBt8tKKT2dU+JYVfNd0TB3MALdWtSlM0yO7sSR7bnNzHiM0eON/tozP
e6V1BkPefO0EIyDQyXEwF6dPYto7OEyyKu/0VfcCQfevtnHLn8XWHXWyIrNvbBUq
Cci3oCyHlESfjPyNRnPsiof+LyZvo777/SS35Q7+/YVyfTZjUSTiAvOWaFbMjXYJ
egQltaooPwtOzBlDOwsIv0zXTe20bhE5zpmMKqDm8/L+gI2tLcFkxJNfEfXMeuL5
qRfjR3SOoqAPkYYqVS2aHeza0N7j7rVgLt/Txk+XQsY6YXIUQVtnx75gJbIEPPrX
4YZQB3n4SaiHbiNhEkHTxOrQXbgZ9zM8b3KiYrSQyocWAN8Sr2zuPP3p4x+A9+nM
AF3135iisOKl8wiRAhiievorW4rpC8a48PEc1v6qsN+goHPE/uHpS/hkGsYF5tR5
9lp7X/GgUJXCe/nSldFUqPK08sJ2jH9kMMYexuMjaft3KW4PQg1Bf3/FhLAZS9j+
KP6LWNywqB+8zS2eSPlbNCdeulIU2X5weOjsd3T1r8apFrcyvp047h8B99dItrUB
lI9G33PEdiFts0vfrEPQHFo/kfdyTPSKwzRvxd6lB/fsteYQM012cY4rOnp02efA
MkQD9uQY+HRAw/HvgMggP2ic6BcHUbjaZt62Wr13i5mD37Zu1BoO3cOlhubEo3Wp
juZM8/sCg9PE7qekoD/KMZlvVyGadvCAH2nUInvlXZKAK5o5WrPDl2upnM9RdKlX
8VZs1vKnUXKEyz/rb0ZNpxN3YjUcyIjFTT3LEeld+/dAkOycg+1bRq1mbZcQYARG
xiRzU+GM86LUGdtGzKoUpck/sgBUA+U/CUfrSTZzjeYYS0gIqQrcspFL+T14dhqW
lYGZUeyIjr4kbPSzAWk0pd8AiflzxgEgM8Egj9bUTtmKyPSpeR72gmuQLgdhzb5f
8CUYqLr+YRYV3jbN/UTF7ROt+BdRynyixv8wF/9+xq4PoU+Sh1G7TAVaJgRVIb2w
S0GE8yfooTfpMpl6obWZtsbHheygrlKjizoumAki+icYL6CTavD0jmiCtYqENMWJ
eE29+xoA9Ag4qZ7q9oUtsDJazoVFm676rXmkU6ZQb83p1m6xElR0kyOmTQi1yRpX
A0NPu9AMz8exVF8BishFwYmsON/JM4kRPvB7oSJrEp/LcP/Cfvon3AT54QfhAN35
sYfMR+KBn9W/sVcYACyNZ1fKKY7nDU+UXMQMcksWQISH5zxHYZwwQX9Uf1KxsXs9
n4AamYBPpvOLH4CqhKGR3/RnGCy3CGSzvvNAyPxS1ModMNiL+yfF9/ZfwfOh2grx
omSEj23BGjHIsoFQFADEtGIM3u2NdqAN+qvBmTI7rSRgYmavyNtyfBRezGYxepqK
e8SZQauemnO9avPXqYInaHtzOtEqRrNLT3Hel6Q+dGKvDgU6VS+9HsYFM3an+GVI
tEq2+yVCHZVVMgtem1yZ6Cpr+6Hc26bYBNOGzOmNVsI0n21fmE5x456CFIT7kIGV
GnHNCXT87wnnnyIqWieNitdCG91ehZWDuG3pIvQPtkzLTP6T3q4nVr7knF+T3ne3
79QG+U0N5DU7IRDRxcDGalYU76w6OXogVUeM0eSsSZcrBnfVgDLofeapvagfRQS+
9heCQ6Z/ut4bqdpZDMX8h0pel93PA+HUXW9w9z8A5GeQHo/DSMtD2gQ5vbIR9dt4
ohSW1l9CCeTN44f3UMhv9Ddsd+0wTvbl0HO2N3+vzoFu+p//rTum4ni/sM7Z7Y+D
rX0WTYh2SxIcfAvCqHqmy5l67lebGrmdwvZAfSm3zJBr2K5W07wFcDyoYnlQBXiU
9H9qchyQc93FVhMIWqdvPFDxrskjPSxpN02RGU7Wjn6pvoTp0wUnoCX2fPQG3WtW
FROjhc4/8TGwyd8sH6JNjLCZvL/qNrXNEBvS7IhrebNJ4lQdHvTwGZ8tcvdjrPDr
/pXUz+MABQ9RBkHIR7aOOz2OVqcrJatXH7s7o70H59bd8YIahzN/4bAYRfZ6NQhB
EUdTWn/iiyvxzX4k/+zP1v/Db3DmGA812kgbSdLdVicUt2SgpB4oba8pKj3XSUYw
FtEngMwGM15PKnpfSe/c0w68hCUefAIaDSDz1/L+aO6G2tnKJtVaVFAy/zNkAyq8
owUGPDHOBLCjgPeDj4el5sA74TKh1hUYiT3ch5drMzO6twMf9dyrlc3FzYvmocsL
PO9O0mAbL0pTuuLMLTi2+lNf3vtbxFgMO3cHt3LWS55eotyBFaxbsRa5vVpy4w/U
7eth3zMfFfej9oVtxWv2P98d/b+sgZdvbQ4BDkaMV4ex4pXz6S8giICv/Qlj7mJo
eV9qNNLa4jW3yutsq7lXnolvaqnqxNuyOWzgBxrm70xIIZ0rA3fo1+pcSI2pxwhu
DWhKHXC85v4MU7bAw+Z/WODzoxp24dIhbvVRKdpDDnt1Ihe8qLyy12CgN+gzbqky
yguvZZ6E7OFbSR61y+KRHJt+kPVPRVampb8XfbBGmbYvnMZzQf/s2nBmEwH4Sdc3
LFpXx45rrcFTVHGcrRZwvtS4Cn3zJ/e3WF/p5xPCLWBMuPXM9jdajHma3VfmFeZl
ympAI4/GYw38A5zuPnfOSIy1GheNQr+twnTovfYHljm9fwVB41qMwCxs4Yoj+XwO
DtzgrEqDlLDS58T4rWQ07VcocDNnonXNFC9op/BCvt//MF1DyZVfmERcvKWnv4m1
kqm4x3jE/OGIlVwvqszJz+ddE9pcPJ0lZWU83IDvQwln/rScKxapKR2v4yX6IdbL
aQUw1fMdgnQutydPm/65WYaRxWcyfOsLXkbiBj4OQClvF6TaqLRXmCezHWd3K0wO
p8LWGnRUuMFTJXwLLiIIUAvOVjHrknSNYeSMxvaiBdjiuoNvtbpWFEpHklDk+SPA
JVWYBbkARFomig73c+TdxBecdcw5cWIeeJEHbP9lE66Fz6i0ZwR8BHBU35Q8+qWF
c5jS1KAY2lYx8xKvnEJnFYr2jBmvyoV4rAuT+BUTo6OAoXLdFIz6bYcX62jCRgtM
4Dp7yw45IL2h16z5gfWzXAK8ZptqFTYJ2UOJb71Rc9F/ZoxSVdqfq4CJ04HUopxX
FUWorflM12vYuVRBCiSnKqklaanz2CHEbCfHfulD/cG6m3TOLKqLU6AX/w5f/Zce
2Zu03BARS6muJnZMBmbXldaoBc9/ms0j0qVs8K3m8MsEP+2KpyAroQI0/qR/2DO1
tiUCEiKUgd35hKTEE2zZq4ZjWQN9AvRdgcqpUI2ESVZHY3mgBApb91TR9KdYceMe
ghg8WnIeBHEfdhsMsS8YNr1budcFYlDKDQ2d7rjBp8CNbrC2BSUF5VeCyCNY/1Km
YT7KOqn6Uq6tPfFejcwVFoBjbP0+7NkeWupQRa9h3Ysr8tqfcFB040DXe61Odkrb
MvtSsnn+8J/7ZjrkcENtKEt70bEWsLUyfhxmLcoZYYZEsdzlx+b/0ecm56CfDHfJ
pNUCQrziTWuzWIWb84Mg9GuJK3kvxPcV61qX4OT2f/k/iqV89v0sHa5Fzx5q6akB
hntan/i89LZ/UIrv1p3X3uq3O56IwQSJZB5qp8hKr+8mXAJEg2hWNdt2B3dayisu
rjQ45uNTi2QoD/h23N5rDV3jOhzE7NclwNbu1i6Uco0G3oB6Y6QdTxQC3sZA2pIj
YbpADzxl+SJyxUjgOXb06ZtCDD8VVaMJYWZ7CtIRs4+77BOZI0bBO/5SAmJSs4VB
MKfUDpM3Q8jY/sdUmm+S7ppl38xezW0Bfm4hlTGo9rDupVq6RyddonLsUGTP9UiO
062mOkKiGgjdvvdkpULecDaRFTtVxvfwbolLEPTmL2wMPJK+9Soo+uB3wPTMW7GV
OGW0vAvNw/bTVlIAIL6Ig7KqwM+gGqrXBL3JoGPtgmJBCJ1KJTwku5Z/hK7U9Eb+
1bTIaURUOYKq5ne+DSu2RyQElC3F3HhA9L89zMmJSdR+MCATbiyGAtWf/7idJvtu
LeWG7UELtO4nsYLzDYy01mXAkX70pKq5s46CafzIgBAqWGogTmn7P/90ybVuP0OH
ysup/OsIzaAIQRnM9UfAjZq6zl6lsWhHNZWdSCP2FmE4LUGW+qJssV33lSbOszq6
LzTlWXv8JV5RuvvdPWsh0koJLeANstTQJzGGPb1mz8OUIuWhGndXE8E2mKKtPwGP
nqjoXbklb2zPfmbRpkyCjxt5d39gW+2dTkzk87SZJx6k68E38XmrZBmE3aQdWBan
LrUHJYd5SOBaMuOI3I5YtBfmLW4MI8bVypDazi2WcBVFVbPubnXdrCtuAd6dg3IR
mGN7wg6La/WUIzewsftp6YQF9ymeCI/wEjYTYTjKvtPq+PU3TdJqqMQqZW/VtiKQ
TF7B9Yq3DsIunRIBXf6A//fcR4+OKQUk+WmyCOlv/tgIZE7XvkHRpcbuVF9aZEqS
e8vT4nXTLQ42uNkduf0yjYeeK8W4bIW2arQ59+XeSMDxyrq79K35BVG0gGY2noDg
uGlZHpMcvPsozjjDGjQBbPpF92zmKUMrdRG80uMi7BuBkwiU6SBuH9xzpYenR61h
9Tjxrh97+t6cbu3Y65HBqMv2Ws69nSGMJwVkBFWk3iEIDU4NqYr+kbJDb4/Ai3mx
tNRK01TKGmkZg9e/0CwlDS3ddJVOMmXsfdpxn/adVQCRp5t6yqWR0WGZapMc+sy1
MN4BTqh8DJEgYfihSrZRm+XNgQR5IskJk1OQCf1VcZJwVLK4uL1PHQCZKD9XiIbC
6zhdiOWgxipstVHC3MvySVAYRHUzL/gQDO7mDcOp4cJ8Zm5LpMkP5cF8Txr2c62Z
7ag8myoNPwZMerHPG6dmi22iFhyzVO2KffWGxAPSJYQXGMUW5wIl3IPqUkID4zxZ
gm8CA+uCJ8DKnP6yTS1DcBCZlNhxyLN3MOlV37wNOZCX8Ii16CkI+nOD+bkgVDS3
KSc0pFawvpwkB+O22cYnu2P7ADffuyOEfiv6sCJUILZlqgKnMEHOIYtQWXoBVSoi
8XjO+y+o0H48bt7GYPHHe1OC0JolVtvdINAujcqKCOiX0BTGV7wegBuY+LM0xAJv
gyazJ1wgOVOIXzmAGYrQjZ+a0N3nSLFa1gt9uOimWzQ4EJPEd6uYwcwdS2hVfw+3
1aNmlF6FgsIW0TlkCtRNx9JhWay/6IYXJmbcsjmgwvGlA9wZXc4T11iXAP/+DHJy
DjYroJ7eTOZyCGwlrbeLRgN5XX5vPEl3BeDJVPMLOXevyeVBXMvCo1MZAiiG0S3V
bo9waqvd5tKNB7cZ0pPAdcaxqQ5m2Pdzjv2OvKbm5zW55LD2xZrUc1AfWqwgL6+y
3XM7aW8pc1p0OEt9ZNaP1R1CqXOA/g0Q5HA/9XTFGFKYaf+injuoR/XdYspSRt9C
mfhYnpY1zp9JLnHpC8PjZqMIwd3YqaZi304LNQKb4mo6w5rLui475NZg7Mvb/2pA
3yFeDe6GWYnBsRuunVbCDE5DsEVcj8YUcq5LhQrG9FgX+aGZgL/DXnDfsOMdnAqb
+G8DlbxMfNdoq219LRDOefpiaFZd4dN5q4wtzV3cG39KaKuGLuSLtki+jhLQU8fQ
Df21GOxShwahm+ENVJz7s/If7UZuru4XY9GqSb4umZ9tWoKJlK8OuSzPaK2znRdB
hLXFG/ven8glsYQwcsBE/zflK1yPDPkQyTI8QP5meF45u8VvuHlhoWNyVgu/spX8
S3nvVkjScDtYRBig6UX/cq5u+KdBeR95aTtGJKY2lJQy5ipcOR+Z+1ObDX9KDVgc
4SKwplUVysJNRz7YmWoT1jojxglhFOp7ECKZ47cRfa70R4rrZLZKBKYOq7K6l4Sm
/cDxhQvWSdmyuGU+YzvIITqkLDADmQjCNympb4JvhuoLvCj7QbDDO32plawPQNAO
+cjs/iPAWTD1RQ4bA5QO6v9q5w8Jc5BSrIIl71rFjsUCgNXyrDi7hBI/C2qD9dTt
tQ81dpdU3TsttfJw19XHw1mf2SNgyP0E93IBMQKpzEd8gY2uXC175M611sodfHOo
NyB+4KVpyH0f+mr6aO7CTiSSycPrIKJ57922W+vH3Jch6kEn+uaIJ3nXppGbtTLv
PKCiyMr/fzUdiQervjDaW5Sa/yY9yzBCVcSO7op0K7Fuhkt2JLnZye+y0HvqIuBT
tsNOknqUIs6KaW0a5aHH1aPpcBIqXGIEHrFBRzM7oCBKQMDVs0oaacDqIeTaPdAA
3kGWV0kyE0smxOa9q5q+07y5zTIzDL0LBcZqeO1+7km03Ir1SdS/68tXDlKDYPmM
Jz/ZHw+BJE3JlA8YQJZDG16j8QH+SZFDauvV9g07H257erWOiYiiWy6URwTm4Mi2
YyKhJ3y4y55hf/mkVn2zVmUbLWZuq2bmzvSMOD2WA7ojC+KQ7wOIzQvsh7p7mynK
BZxO8T/x47gt6Dn0btnLTKXOzSZ8u5JxQG9QJ1wG+PMMxXIGTn0MleG/EvUeBwgs
CBptvUHjbfAUv8/U/uYcmN047gEsH8zzxF4oW6XE2K0IXgL9tvIlbPeILQhto7pm
YQIC/n/TKp3S8z6YEEw1RUd4OiqMajkxoOGq2lauuSZiP/aEgAAZQ9hOolazKHBN
3UZ8rVi6p1FuAfXpndm549Jlaf2jZf/DknhODlk0kHv4/6E7D7P8MbvuWB3wmPuO
Ir8HigWCpE2Xt366DJ8cxTSAqPAKrp7fD36DPYVaAxjB0xiaJ7R84sYsa3gMYWtN
SCW4OgVKB445ldMpyWmr+GYKmJ3H2MRYy1f4Id3Gm+XDfM5nMD3g+GyzmCZ+p9pJ
VA5v+et6OEjm3GrfFUBSouX1T2VZ4EkDyPObT3JCEtxLGkUxh/d7hWw1TWA3Gai2
p2chSMPlK4VXc4fxXC/Pwjzsd8A83vXabOhbo1eP1Q/fu1+vwXxer6sOMkfnVrP7
nCTsJ+CsWVM3UY+nLcEurVOO+4xw1TyO4VcdR8I2BAHzhGJjRsTaI+xe+MMebqGr
UjOMWv7vK3CaZ6Eq99r60ExiYo40xltKUmHi8LtoqEo3xvD2y0Zi56ihqANv+xhI
en1TM2IlrJ1qcydp8Bz63JaDO7n6Cj2ay1AGzFMB8opt9MNzWq3ytOIiblzoVZNh
JSrHLAjiBUiB/9MOR4GuSJcczInttvTbdz/0XY/ETpqTB4w1IcNb6ge7ERZsdsre
QUltYvPxKOaxumE4CrpARY0ypAoCeOoi67zi9Uwb6AEsQqGzFuggr3UYEqssA2qt
bUcXPrqbIJDeDcpqR2dIi0d4DSm6txEq6YSuteEMHuvcGB9c4a6wWOi9JQRi6KdX
51S0Nd7u5z5TaYxuw1Sn253VHbmOykMXkdpuWeFSn205Odr9muRoWRH2oizuphgQ
o40BQztvq7Wie7N7NQ4bfljEyoTjFgEFaXrv2/7/RXz1qo9GmoqfI1d6H1X9T/5s
SdmIE9/OioBeqvqfkE4vJ88qlIztx2ReLQTsULF04nZxXvlFT0x3cIoJcsYtUQIy
ypW8mPIoRCF23SkQmQNodNKPjD7KfECU5cAvrhPuZpLXDX4qgfQgZ7nnC0ZLrqnJ
rRv0afH27Onavoukmioa1ka9YpoCQ52V13OUXlS929pFTEEpDlIxSDvigQ1Aats6
934IrJjJDV8pd0tWP2MiFbkqp7OYqPiTIVRGM26d0Au0lBvd1MItRePTSWUzc3hE
O/ACSBGlMEKQEKSrgq8JArLOysAXyRV13qgT877K2ECG+PcTgU8ZN3QLovtE5lGL
HknjZ9aH4fCvRqh2hg5Kr7K6VMwjo9gsOY9eRdIi+Qp+jxTbFaQ/usENS3ZzQy73
NXoKF0gRmawbeE6rjk3jm/IC8WV4hGQ7b6UfLuSdcktEs6XTaSK0xbEpghmk9Llb
sU6DL3Jb5jlPZll+9NlRQumAvWFQeuWlL6Di6pTuhFX+3uWchS9dTnsOUCXw0Vsz
drHBLWxqYbN0/wGZwslsAwK5co1qlxs0J8dPBnxg0F6sH6thg2M2vIzaXDVoNiCj
tpxGCPryDede1DIUA3b4XRF5UzIA0Y7PVW4C/AtVint+6SXuOwy83l7aoC/exkb7
EK+tLwpsQD9Lj1iC3nmNaqfBJgQe20OgPQJohvSbkQbJAGybTzpEjjjJb2ZZidwY
Rct3/8UEqZAil05OEEh2LVyZbMTEFnC1t8nMsaxLDkEh5PPY5jiVnJVCNKdzzFRE
Wr02A+oOB8E5CDswEeplDlZ0ZxhQfG5hlR+/VoDxBPqrAyc2G0IFktsSqwi81uBJ
b4CsE8VgaQ/rhC1dr57iQNR3Q5oCV8DDb10250apN0siGhLU0STDHRvN8x7GZQ9z
uT6JANbY7DzSM2Veglxw3v+bUYCJ5r8LjLu3TS8PmLORlRISWDMJ17ESK2RzTTl3
TlXQI8J35B5mrvhuIWWwLvxb/DSHff5zkVUrzaw6Gp0tysFXj0gFT6g2f/9q0m1L
G1VIgoQlsf2oSv3GEKubiNTaqzmeqCCK1dA3RZSCfplxrl3WhBI685Dods6M2VOb
piL1TbPyitcdjxSlM+4QeQUF7/fPlnaCL2BF7jMDoFBc8m+dM95PmFfn+ozKGxLH
lJumxqaoZiatSBw6tqA3hSQaCgfb7+unJBpv0+ieO3ZbUIdi96IpEr0Y/dBRgr5/
d5yFHV4NXrFlMIp2r6PI8gqfd5x9d1tj8qcGyab66xcLCefKnJEOw5DidYIE9Psi
tuWtRuGOX1lfrmc5nj1ym7jeHQSpbL+F2+IXuDGimpB3bwzbCdsyz5w6jHmr9Fgs
ZdY4FxsMtHNsxp7jlXOmw2EOkLwCAoiy+C/R1U6d4qWDN5fQWphnO7DQ41gJ7sPJ
kVAmSZ315UoCEwGPXAphkK17aiyZ1waOxJ+sZQeFYizMIEn2e5DaThNMcAiEOBYD
rO1ALdHGlD1v/zHx9gBSjXyd5wO4F0UDTwllgmNrXKbTFCydXc4MLfcqi9WCcfz3
k7vpposjuXDaCtwEG63cuDNfNEBbtAgdSBw3opFlGzcWXkHrP2Lo5MIhlphWLpsZ
uyn/jqxChX4mCMGyFWT22xFGxPgdXiJY5LWlNq2Cv0tiotM33Li96O7CBLPtkDxj
DVlGTxZO1m6tSVS8lCnvckyC+ft99PqYYJCyLrPhviTRPMdGVwPh9HsGW8qWLSQ5
50jyMIrxVgxpZsRgujbYDgz4dY0Qf30KfmbhNfJPVrlgoDnh6b4+bKxlGkNLP9rY
th4z5SW2xLRmA5g47+sK3dFLtyPbT7v0JgNGgFskgQSBjafAZcV3S2YFx0uLoPQU
Wd7AEOd1TK7Wcb3r2lGasESdwGxG+gIoZ8d0+TmZ+MTVaGRnBD4XaO9vrY+NFMCv
eVaLxwGLQawMcO9J8lyaZjzqZTBfBjG4sGOgWpxJzCv8HA3yKi6oMuT6fc9Afmj9
ORT+bzRIS01tl2F1BVMch78zBSInIxoAOJrpm6Jg2F4Pj/IFOLUHI9ZhVYUbVEC9
AkRPo6yqvf7LlIrWO4GyjH7oWRhchLW/5pDmnvvxVpa54Gw/F8RNNADEPD/HkNGX
2mTo8MzX/xxOLROEHYrbkn1Rklr9JxeqxoHN0CdjEz+DTq2klIF0q7pPrTAJc6FQ
lxBZYFxtGg5kc52C9nKYUb44ZshbsZB+NHvkytbIDZgmc0IKKu2vgq89WeMQOGlI
B0yUft4P7F+iKaVsM1F7j+NOm1isYOA0VrO2YzkHvWaC7xR4qYI343WO6JFcWbd5
Shpj8J9YjkIDPJbsuq8KlKY07aQ/rHHvMsVLbQsEIBr7s7D0zEiVNcVYsLSqX/7k
fNKD2asJwFIUyGi6nVbf1D1VEv7k0Is6KGxUUyy8CHGmg0EMENrEJOuLofOwHJbA
9hYz4T37ymF7FfzQRjkzPpq3yT7MJdS5mEvZ3kvXiSnPFd1tvGBvFbxuZagJnvfr
QBv7oSvMhkzHOrLVfZ5P/mk3Gv8izwY7rCbzXUymhHyJrctTECaG4juSHScndmsp
1bWnUz6DTW6zCrFf3PKneeN7Y6GzTElEs5r63RQfp4BUc4ggq06B2hirugI2N768
5g7n+nWqnELApn1SHdCLgs8cfwgjWqrRdakHzXiYkeqYrJYANRJmt3Qbq24vtOTs
YYjvN3H/VVNLVXSMw7/lyWqnOl2x8EXduj7CPhPi4s2OxxPrGAMHOpuCW2I0sPFO
c/CK7pfPI3nu0gJGGo6ROUn7vEgCnTxKgrsi8xPRj7/bSm7BNcgXtNvDE7RHXbOV
YzcoQU0Whz3YfvYsUmWmT2fuxoU+x6ryEaOsD5e8TqUtmJjUPxrqVSj+C2vgW+rM
e+QoCn4FFo1o6+qH2G/cWdmdgB877271KMjeH+erWNJiYwFcv5UQQu1AILUAwSkv
cdwJ6ryl1YGsuEqI/evxEENLOugo7vbyRT1LHrgZar3VIjaEl2Q/jO4q/sZiEy3M
XcaOMOJiyyb5qJpd8JsOf/eJDqjH9n4AXhUCEegYJxX1XjRmQg8JnZn+2mb1hjpr
IAeinc5Wf8VKxmB6nYwOeykCKTRO4y/xerc+i/MoDAU0WE1YCNkPEsP2H0yfkFsN
HwsQm3AH+8ssE+IBN1v1o6QX4ZI7XZTD9FWc2kRV5FcAJLR8uIzuo7KxxNk9hzlI
fcZEyIP0KGSAnmL3oYbH0rPcvVy5DMDEKeXRBCSndqy3m4bCWUou1leZaygkx94D
q3oKbYOmcQlN2Yqb9c1S2hxFTNLliPdjVzT6tVPLdu2C/+k/RZ+YRkCzmPLpEN/w
P9XC2AegNY+gbnCTT1vdT6P4+eo5xjUz+vM1QQb2pDR5XxSBgsPDR8LPtQcPVeeJ
p3f/HrFqZxayhpddsokf0nmHiM0vLL0L5OTyAGpYHg8Lu8Nqug7wjIhKcMcL3zZc
rtMGPGaPbUxcMbWFrujJIPGINkq/z/qVNYfzJ/r/PiGlw5peM9f1eenjXKusaj+Y
agKUREDqqzT+8dUMvEgINh609buVg+ereoVVwkEyUEuckW3xYlTe6yJplbOTFo2Z
uJvasEMR3q1Th9N8DLztQG73NKUrWUq2Pi4hGLF45eNRALcc6Z/i8chUYUngoN1v
GB+0DYEfX9EjQjHenvK83m/kHmhlsEy/Zbs1USQ+lrq7irNnjhmJgfcSQlzWBGNB
qHIlxu1NYRBmzKzMvKHkyJIFUrKx4i2gXbiddQPdBBVWm/PFTJeH5B89nV9BQCab
NzeCs0BdJhqDCG+H3vKzH4of3H4i6AHSN0YV42zxavUC0C+G7hQitd6zOy3aWdNT
T49pHhE625jbsYPeuVWBHfPDy0zKP0AJf1FLCU3vbQSLb0fQ06ALQQ3ym//gQkbB
mAHf0Y+Pe4SJEXIPnOmOeVKiZietvb97zwc5YDKAPSfWG0J8J3090kzMUXaI1cx9
grNS9CTCU3ME2lr0s1tVlErJEFrQgQvUinaTAUaqVPHIQqK3uC8FsIXv7MsuWoJo
Y7lDhtV/+n5jqQ57ianOS78qNX9elMMHdCrCwdkrcjdcRYCQMR0oVsh9VGRkt96N
wgZguECz0wVKiEEXSwz3M/F9iJPr4WUBB+5jIvjRRVcnzdGzXgW0rhTUxL7QiIw0
7ccOKJjhD0lznfzGMoOIBTNJSimAimUCZG31Bl9Y1WqhG9z9ecHLMB9dc6LNRBoe
XjPZkV6UfymIS8S00YYQtbi3jcFLkf8KBx5lCJPmsXRoD/bj5TWaDUd7BqS9m+Es
WCnbcyUnk5LZsNldc1j0J9k0l6X6EHmoxPVwbKhuu+GGEuKkDlPyiZP1De7fK3We
ipVXbBSWkh7d/0RO7L6mg6Z93bUphE1xXiR5odlPWdb26VcNFxbpWGVbvSU/UrtB
1lQc8JvUo/oro5Lp9quO9wHtTS88tt2ElHsQmCoPxo5kewBRYLEBm/6gT5bdXXf0
n+KgRxZPIg+y8nV8abLoDXgrybkR100p9cnx7HEbVnxC+7fqTxo76bY8kHy1AM8G
GEzNxjbb3Xx+3PAG8M30IH9nBZhSZZehB8ksIB0Zx5d8PXZn/rpuHjA1QnUOcI8R
fHi5PY3vrM4fluS8ZSo78IzOqsO0cKDJB9JGqG6/3YuzLFAdfVSVJqr0A7Y/DvTX
ymAEybx0VENFh3L82EufnZgixhl8PMeS3aY8zltzUX2LxT/Jlb2CFyhTo9MfmK55
+hUet/F8+DJqxovEtvHaS/IrmpvVSxVbbQycDfPv5cgyAcIGG4r9sFeMStqCL8Wp
bNsR8PK2GTj5Y4Ujpbl1X9JFDNUaUekmpTSFeVEVpi3ZtDk9PZBT5anA1fSrt/8M
19nSIi3v38fJSWZjWqnyu5murH9ary3h6jlg/RH+3BCeCdtVmickzWd+QAVaia60
Efv8sIaoC0jQYi/vz4YCPd/slfexLoU7In5jXjHoWWxl0r9zJoKr5rqcdl/8fd+Q
tg7wHo+yVhHYVNW40LQZrm6vS47EbUDuYS++99mrlCR03ui8MnFfj0oZPZ+Wgo3J
o1pBj1P2GfrJ7Lp/AltlQnFYxnHQfrCKzgFgN569gnz4YXsWhYmAfDGJnFUqE7LY
ByhY6p3YmWYiYQ7IWFdzwW6n2YWtrVZ06ExOEMnPEOeIXQhLA9zHOtJMLQJCukcl
+zfoXPkIdo9o7OEWg+BrqMTjvxoLS/cXH+ROOyZTGAOgUtb0NEUVrjluDM1Xfxl0
1nD5/QuyXwxlnO5yohnhynrHnPSvZ8yth8+3YT5xpFXAAOiL7176xHQghq3pBdwg
AF8c8P945Em1SdQU0gYRvKY3htw8uqtAjshZpeUL7D8RU4kPXjM24azHs9hrN4E7
gNnuWntNP2I1MTQPGcs/UgBcCYnffJOeLRGen/lCIIfZUoJdAI6/oRcBZN6rjZEN
dL8pc3H/0M19uv73YPVZL/ehvX9eQOZkMzhCSY1/cbkYHgMd2gslkAZNaGlgk93t
LAEeJe8SIeuqKeOC47KZL6qiP6A/0QsrhmEZuvEv9m7IThjdggNssXN/fWAiXUOk
+FME+Xt1i9Wmr3Ui8hBLlZ0spslEGlaTj+1sEIqxM0Pzwwb7Kvi5EwAhTUO1bbFZ
C6jS+DISUmM45apHWHQgpOFa9NkaaWaVzZvOOO0ckXN1n1SOVS22hogqrAeVJssz
z5tgYb60C8pPseHlyOgWowNy2qs9pvULGYmoHe+NNz7U6I1V7+8OJ6ITP8MC/wBT
yyklK57+HzaDYRBeaUp+MLQsVrHWWFDzrLKLdP07h+3BJQon+Zz5zRy0jsAjiKDG
eC7KryO81X9xMs2Z8O2stJpKL+h9khnKFXEe4xFTSrzc93tzTQ5dMcaUbMqCfg24
9Z4/tRJk6c5QUHx/68qyvcuiGTtHC5QHPqQle6z9KKLz54AM92eR1TBCgOTXzvN6
JjguOtMM7C+yk6NVcgVFql0D/2gLea8CV+MPlyn850zdDErHNvD2lyojFEvwuxby
jS9LrlgtS3U+0WnAPqmoHfJkPM/dJPWyOPzIEGCsj/3uBFYLLWNjpj5auCS39XaK
bN5p77o3+i1nChdRqeM2s9FfGW0XQwL4dp/PuvpaAKbJtN+buK0TuYprRfgXgL6f
Rlz7DgKgHzdvjBQPrXUvksn8uRU/ugMGPMLgaj41eITNqqgp5tG6XkQ/WRBB7yf2
yGnthWvscHuNj8GJrCJ5DPvU0xSSXCvr73V8cdqdMPpWtzwdoLPCmojer94oBygE
Jmg/7WHkqPjpTGWuCkeRKS0k/hIqFt7wle6Beu51zfhYj6M+H1xzjFgEPHEV3yJU
NiHiPOZvSYc1OM99xaZHSxEdqepCPF2K/o5UAdfjyI7rrc2yblOCVAb3ogfRhLt1
NVl9tfstIoUUjkEdKdlqCzPjfP2NT+k9zyGhO7jFfhbF3gaP4vvMUxz5AdPnnpFk
Qf4mg16XpOo1cOXfqxFEMdv/ka9kKvBNjBI3SEdDG7PRtAcUBhz2u/a19H+viHn0
5JKEignJ/hu0ipgTrKdkC0CRoLY5KTs5Acqb0G33qWtAfe+2sHYnbCTM9vAtO+p6
hY3HbeSd5wAls+UDRf+dG0N6pFaP5iBfNFze4znuQTXChvUfiXqE1qfBp+EtKou6
MBnGFRgrLb9sQwMmQeCLi1oLwlM/F09zQ+G/pgB0T4h4/gYc8FIaYb9yr96Zh4M4
EXOst9xZu9KJeQ7twY6ozN+mu9V199oENTFRWbkksjr4HpraQGg9JLyUO+g52ZrI
abMsph3jVIQ7nrl9wVJNoRyYt5hjOBWoUdfLLDNARNM4PWINVz8ee61i1CWY0IKK
4tVm3OewpBZHIZSh8XdMcwjVNokqoSMe6ojUVfZoe/h5bvyBctA0AA9rFHhy0674
E5K5MderdEw9PnfZmR1+qCV33MrfNjaxa1N83cnAquwc3Vhw73mofxrifV7WW2y3
zju0Vg6NnLtBh5zrFQJvDuL0qBDQtOUfjCrN06VwRXW5yUlG09UWdlzWN9mHtJEm
eGIuQb9rnO6VzhhgmotZ/8WHQKlOSKbOjU15Gf/eMnHLLGQXjSe/tCXE9mM6SQvw
oL4Jc+5XS2K17b0BCYeqmsSwvFUniFD8z+0OxGAzKdZBCI/aJAk1+sbFUCZtgiJK
brRLU4jeh1zW0QlUmQ2V+c3XYHbHT1jVxpHbY/yq4NRm58ZBStQkAlAcNG73OEiJ
5WLwnsTZbaQ5u3fCuIseTVeRWvKlfJlzGLAY/fPubbGFuP6rOlrq9iiDP9JlDFOM
2n+/e/D812id54m6/MiTfgrx0higv425DqgUhZs2ijvedzCqvdJjzwomXEhItePh
zVmORyxDyJyNZR//NphO6iNRsScBOvkRbJHvzylflYm0i5q+vBlpI/vZd7GGRFa5
+qYlUTLfULCvMftWW9Q5PmjMCTXSQLIOz2n7YfDLLc06WND9TF/h9lCsFz/gR2bM
EKVZjD5o+bQV4XPqDY6jRG0USB/Rfc7sO2uErhmNjXAArjyMo8VKPP+v6GMziKpq
XT0KAHuA0DoLiDkM2VphMadvi4TjSNcLxQc6gohBxjLSqJvDtJdoI3gonG8HTXfi
4uA3m6vNk/e7Fe298HGCm95w9Mor1S+EmjogfSHijPZUwENJqpOQNtu5aFG1yVqd
CnMaoPdAjHHFmMjzcOJDHvoKcMnm7A+28PEUm9XG3qPj9FFdaOHqNn3c2wmxAZ2s
QRYyDbcl1d6fAMDRyWKBaJtlpQxX15Re8qUC125TFSnM1IWFe+f7oCAN1Rj9NpS8
ECRPPK/AgGd0vlUKAA3Kv0SR2UPAe/i0QuCJCEKbru11X7pS2NHyszqAT1d0A+Lw
rlSfLqKGxRLhx2TDpfVW2biBkbl2cYCl5hEBuR90393yoHfJZYsIJdACcGsdRMJl
s+jLgl4bbmOfDboaKNOmQ29tjSR4+Y2zozFlo9BcPC5mvRXDNTxmiEhl9NFh41Wk
6aRbaD6SJPy475yNBr7qkkrceWoUvfVDmBFkZjAp0PvGO9jdcdLoAnQmZ9djktS1
zsyfm/o9W7O54c/NLREr8bkl7RKrnhmyZXwDnDv0hseTDU3bbzDnIoY8v9puXiFg
0TxO+dk5rNoQTZrAnUQCIpZId+Lxo02UM9PDudsCSVbYvMFtkfpb/3ppSXeyjqB3
ywZrKy7tSD+xyAoDCsqwujy23YNvnCZ8PyhLR8bYFSVbfziMbUCV8I8uJmF2gN+t
wK/mea324n2sJjjTa7DYpCWP3RcjLu1IYfvPDwHd8Yx7+bYw2TcxviHYGM1zjo98
kLg3xiijxIyajXnunp9+y934pruuQDwmOEoJGIZ5hKhaulSD9UjgayN/8PkEZUbp
PdxAM4IgArFrlyNPFjN47y5wbDeLfZo8K1iB213tJAQaoqEqgOIfaeYhgVKT4taW
S8c/gKjMeW8M3tuTylu+5oJUS+A/okklpyjd3zXGWnl/m2qOQbTmAiTFybLxy/Vs
qGpae4WuJZmyJeMotwLJdEpXE8VQz0t9QcFT6eEdpxJG4wVPhij8AQOksp7QgQCB
cTsYL8TyYZMul3BOuN20TAUaqr6wVdcgjayOVCbBUZLJN4DrAFWoNvANW24Arf0n
lp+3blmg63V6G8ZLuLfhjE6f694xfV41UprLlMNLacC/TlZfnSG3g1DzRu57Oe0h
0smpfwGy88/8qC/IwRSmiYqyijWrziqYHKkikMFG08NrGvT1w4qsVK8/u1nfRmQ2
cr7UYnXz5lkengIzoI56O0Oew0WLj4td3LQ13MV241d2+DdyARsjWLCtmcK7xbZm
7HIVyZHfBumm+7N3+C25GYHS3iec4YTZ3GjcCsC8scAf4/MxqdWM7qWiaQLwF8jV
M0v+7QTcb1V6Oo3adJI/FpLSiqRoDkt+KaYAGuNtYpZRbOxK23rS1GZizWRBrtLL
DTtKyB6U2sUgVrVsFYBVW/OZfNIVEbqWM9Cs9A1yxPFpbEPoLoeqIYxc5SvyPZAT
PcNHOYxHZsERABTuIdvVM3uia2VkEGocd1oCB/JdqY0Yjpv3uN79mcE2jPucPrXv
uS3gwXu+UlWChlIsdVakKslbz0buSWj8gFQo7e0dY8ozaSQ62StfpASOgAU+Cwn+
ZGZF+N5aFpoF1f8aViEux2Fp9NcgnaOmtZaXeUkZ+Q5unrJkwlbeOi/LwbQrPkPH
gymMDhGMVylK43b3DZShyBZO1h9vvvNlZ0CkF80SaVTfU8f4Uu3cKOUjy/4KzN5a
7S2biTE4tjdGjWcJ0ok9cId4ZGnScfs4Om6s1OjMXPbSXgKfkxtog2l0jQAxHOg3
5ZV34fq5BwPi2bRpf99jiq3q9sxW0P9R7shW6mQbiz9ARRyuyfD06zOjEzJWtlgw
O/y3bcWhmvNp8bDDmIA3kOpIb1n+7C6Qj0XZnBqvH002ONXE2DyjPIJq6IyKhW2A
P8Z4as21fq0WWCQ5RqzjIPWb2OOS0sgmZDEwdOJRyC6jPGAEGyBEFCAPQKaRJuaI
MNjTkbmiOizAm2VRZIlF0yO0oABWC4SA0xyw0eZR0qZbyT6b8trlPoWMqnJ+zPbB
RH3VOWvcER3ffOVCh2OpAuTtXlufYtfPMqjUaPWvLCretNh3vN6SKiMzVeWSKt65
5VzWjhg76nrmFYmnkBGAa/3o9eU0pdD6AzIMD8eS8JkMtimse2B6F48dYM2qcGur
xQaCcQc0FNb5tkOKnqqf4tocPGKd92bh5J6OLdVshyYvvJizH5mGEcozI/K2DIun
WSRt7DalUy0zAe8jnkF8dnusY05N2tzaX5XAnrM0PhQUTAe5fyqypgTJkjPYlMkn
J95EDp+nOgp5SEg1ga5UFBKko0ihhy2K9UQJCBz0Jsuk7i7ldTGupnW6onz6T3zI
Jzh2DUyBZ/yt1ppqYTzieC2wSEh7+J2jbpbP+baGpQvFJnO/RywGbiz5JUP3jMoq
7+cFMJUgK49PT/ly9qZFYG1q8NLSKvjn9kfWsOAvSeErduvwrojGcl3wj2TLAzVK
CB8Zco5+3lE9DyCcCPG3T5I3uRvT6s02LmCrcmmkbRyl6OpWc4Ekywg1uf5cWARm
d9ox1qnuXpz5/1NsxWs1q7Bpu73SCCjf8tVtpRusF7JyKqD8cmAKJJkXhXzTkAkC
bWju1Jo8fHm95/gAG2ozYq0CQdGCFH/fPMXm86TqYbh2lFahH8SYA8bKvixcnJZB
WwNIcFE8x/neNZOK0E68+T4AJj/V/Xd/75COaVLpqHba6BzvhRvWnm///CBtGHUq
s9x3rPtFCzYXflTCp9GrWPLp0SbkjQaC53Zw/5deto+wfNzam5cLQHCUr5CMVFbR
0zsuaK0RXRLPsNPWDaB5M4WFtNltewh7m0OdmtdEZR95d8lQdNNxVmly9KW5WP03
h7pQxOjq9Tin573LzOG+adkW/Wu8Qcxu0YHvhdBsryoeI7VJuSuP6Csa+FFGuZe2
2J+RYpeNWEca05CMIRC6NYMa1F6lk+rdIsk9tXNoNLajnbwB7ETBrGOi8ZsYm1Et
fV8qlCqmYr7Tn9j0NiqBF5l1IWRoDUDngNZSlD+4LWqxE59Kqvuq0Oxp0U0k+Yxm
o60CyaER00T3kSq6AxAI+WSzhIf2xv3hbILofzLy+iaIKOMWWfFgw7ptI7AEhrZh
cnCNv2n8+yVAcVtd01MMdfhLXvX3RXuIhpbQ52GHaI2V4YY5UokSqCHXUDctkBX/
3xfq9IxAKjiUR/08AYqnuVO6PyVizUopVKi08fK1P+TQM54Z+eVhX/wahfEf2qVZ
KulIVwochP7GzyfPzY+Ta4wtzI6tsi75z9zHqyGt+sXHpjMwbrumaeD8AodpJxD0
VYvg9jU9ugkuS1yZd0KYfILg2uSlNmzYCRX6So4AyI1eyWONqTAUkh/KHhGTKLFE
6l02qGBqNao4ejblYDo34dFmES5PyqnwclMRz1Eky7QYEdtz9ggXY+DWiSr8aix3
hyiotXI9n6NiwbYoqvsEVI3lyMzOUL/zpFpKgq3cMrsCUfa3LlV9c1w3JsVUHBq4
JRDTuS4fP6CrxinlVDD6XRU0VaLeDduYISqAnp6CpBk2eRY/fb6nqD0wOZDtCv6u
dKJFWVcp3laaUv4xpNYRDL/PvtnhemE7rCQBHR7iEz6/0JNDayW40PGnnWvO4HsQ
pRGRoUtUFYy9fnOl0Q2Czx/2uNPFK4C5nC0pTSL747uionplJtavmZE7DjCdYVr6
ugequclGF6mEOHF/5KS5f03yb8+1D0zi8UgJEpWUXYXB7NZrBzyFpms7szKgta3u
JYfloTaXYP77WoTLwS2EVwyvlT+IjZvaH/z55jUvcLyjp5Rf/M9mY3+8UnsRfPq/
sX4jwp49IBzgDc+nj7Y+ySGu0lgH1CIT+GBJwZLJEbhTzkJ4CfOSn9GhCimnqVnT
u6UllktHRTdVM6n1KQ4KKjefDVqD0eLJko/ePCebR57QYl8tIMFgRlyoLAtbEMXY
Fw31RU5Cb34WtCuh/tJf99AcCZ7yIdXCYS1wSwXMzhs7MtVWJhfrbOnCrtyDdhqg
UvQXja3LgQ7IW5CCcKqcdPZL0kWexksf77VBxOs+/CwrpG2Y0tTHJ4b4dLbBq9Vt
xOgWYNhI6us9fOdeP42xGfyZReRZKBF4y8wYQAYbaCVS8PHWTcQsbOJCVRZIZYmN
8b8x+YWJdvpwnEM46NA4xR87iCznTdvVT47iOHAEElWl/XOWwzUPMmC4KLccuVwz
DxqdKeJgdUTi0N26GolsyH/bbn0FqTYk0WnGahyzigGimyUtyD7+jnNFEa5KT1nT
zM0Z+mUerb/1PGI6PfUCrZ70yFlOn+XGzZCZm0Fp3qY3T2ajBlJReWVamiHQFmqm
kbOjTRZ6xINS70hdjrA7qESSHnBYHVcmcNXTyad+oDAtmzRhqisP+Qa3WaobHZv1
RQ8BMk64pMCRuGpGJoWrPxLISrg15mB3GsrBx2ahw9z84PBbNps+KRFPbdt9Gxgf
Tu7oUjfG9TBw+QEqQIAYfqqx18vqerfASpJelXWu/rCGHYrV2RUy85RvPJLzRLmk
mTu2quLUAaLroHngHOVOXJ+2qAxVBtOt1r4XCblZSw1mtR1SW7LQh2Dtf8ABtFKs
Iz5aq8h/DkkfnoUaAGOgqNPRWrFut9nvxi4p30gaZt19zwDLRzirlMgLr00SuIn7
f4l4DhRjdz5FEeTIXPBJibADwmxwKzVUMB+Hs39oA1YSqitgE+RcSkvXMgPd+HTb
6UMGTXWjQmcB46MsviRwnepswCecOawdYkUBZ3ORq5LSG/kjuo7i1dRSvkhwArSh
SaoO7ZFkMnD6w8QtVg6lwOt/+VTDZHxs8S82Z5BKKVW1haWV6mN3LNh3PKQAKulr
dSw8f4Y0UO4a+jZC81MMZcPn8hjZfK+HoAbxC1UsJJortMU4FxJTwtQfz8NI7bXP
vXpBB83oCi4O5klHVNdhj6txxD97Kx1n/6+MdyR4j8t1tNlCqAJurHIvVH82Gt6V
NG3VDKYV8sEvTk2O4yBBtov3jhx9gsr/udTkzjmLjmbMkjYAEP4ajdEeF21XX8CL
ZmpzIjrn8BbCUl0MbTMZ2pQcmLQC+g4/TL4OjrtxwG9FX13K4nHVqH7AX7vhpTs1
1BvmLmMtRm/sT3+3wjWrZ1ZM6EtfmZUUwXvszM8XoiEILW5ys/BWsUI6l7dAZhj+
nIidyjdiTj4wfRN2gD6fIHoDNiQlXxzG/9gYIcfHRoBWnQXuz+PEzB0BmgDZr2O0
xBQXOqGEwb4gjb5l59b6QlNMqt4/7SRlcNbvK2CL/ffsMOq9Ahl1Ebd+iDlJnnKS
gngb+glVfkVIYTaFDV5bYra20pdXbSitamGuKmynHRSW34ITT9Oq2c0WVaOYYcpM
dnqboJM3l87Bz+xJ+kj0/IF1+2JG1MBEW5pJ6tzGEDKeHpbxCQtprWD/04ypYeRv
pcRwkB1Ezr/3Pr1okJ+1hGyL2QEC70HrPTBKuCyGuMXbYml/CbCt2w54m3ylqTzp
qB9aocEIbHh1HKi/kArAsXHFuM4f+SnCR1sYpKL0lqxFMrRInAVfeyeAeJL4se/p
QxbCQVPao/k4Z1jThKPm1c3MWxFEwQsPJHYycEKkEH90nQuJaagkz22QpzdP2LUQ
FSzkirOQQvPh69IHGMewr5lhMnZqJWplGNDxUtSGhI7WFacDNzhGzIlsQlS6DUEY
blkU5UXxIzWa/fm0Zg4cH0wU7PfbhyqIdkS0XPN64h6Hexzn9FXCNqLzgGPwkexg
rWfTuIVzKgRkMahFQySm7FCxUxVVNbVn6mUk16Zp93ToL30B1aamQh87w1yaO/oi
GtjQi4KMR8vjSihP7ozX07kdlLpKb0FKhh1u9GA/kArAjaJ90L30uxjqdQM+zeSo
+i0jX4VlFUYZRpDBw6GNtB49ucUBbuA3lAf3BolPRS86YIGGA8BzCUzjufHMArmo
qEZpXLIWManh5pXrg4TmnnYSg4egFH+isJfAc3OcxC471QWKo0UP/oI4GWQMg1yT
uRI6J0jnIHYCY4uR3Jz3OdUyLrpKnSn6mypcgPV2GQreLRwQ+LdB+aO/0YdrL1Zt
yiF/Em1DRbW78FkHm1JOx5LgZl1DLuMq4fyT8i0XBl9dXdoDfqvA92DgGWGXJOVZ
j98ubWqGDD/jUK/jf45lhZLCyRybG23m/L6MQ9DFtkqWgMrTSnccbwXdtRqRBsyH
W7hoSV7msHMyi4q2n1sBYXyHsCsV2DmTVnT1yOagGbcX0CowwzFqrGK4XAxyt/s6
yXerIpBhJ6rvMx7qggL4oULrgnV3XigBDOUCj09zAxNF03dNanl5LCMkL017ttu/
OBCAqzSXintL1yTb26uWkEvQPddcY4qhbbWAtetQoTdayCfPS9vXwrdEpw4GSS9L
tjriIwcIl0sle949yPoZMRgE+8F2I8ClwnAb6WKn3w79MjyGpKZja3q6rcMmgI/a
RjHq2BFP1Z2W9+dHEbEl8mevfsYvIgFiFn6SP3yCmycwcSaivKE1AcmVDzjoYjyh
rH4axJbdQWSn5vF8sj7aPszDgI/k3rqqcyKiNAgG0yyOyGmDFx4X28COjQjRnRvg
kyc8l8vdi7Jxwhz/JvvJfdyIX1nkNp3TbqfqH8pes83M6bM6F4Xy7AVhvW+THnx7
fEF04sdic4g2K1T35gbG7a2cvOiTJ3vWFFuL1xavdidok7Irh4z0oqTChRYKrj16
xm0uwiBchCN7sTMQjxO3Q2tlQutlVCRrCVO0ParZKA/WWYrcTb5Ti5Y1h4bKvX1U
Q+WswssPzyqzjL6xNDZfq1wojz7nXfdtnckGaTXPNe2E9ibmJXB2DvtGxDvpHeWQ
3274KbXoJFkuHX8uYypeNZgXJEsrKCLQeEGOT5mJ60r/5RRqdKIZKA5YDuqhQ7GP
LhnqVq4gAnMmui0Uo6QT43wG1wZssyrqZftT5sUdpqj6VBu8p2CCPz+9YOFmpQO0
WA5cTcNCKYx33VCCYb+J2m5C+3uTNEWV7ZpTT1qCWrcGAW73oLyabJZc1Ppe5HIN
KupVuKfFjWbkAeo7U+u7YlI9QtNlWAA8kFhMAjRbtjfp8k8NhzUWDsWTdMt8rABw
2v6hc1/Ugodd0+kBKUA3L1zmKnqN6HiGNhVu7Yy8AuHjcIKL/y/634Z9A2yoRhTy
63ylIg8VPvXXUEkODg0/YLia6FZbaUr5a5Tz/UzDgOGkCgfliy5+ECtHuiWIHGcF
jA0J4LLWPRl36nj0e9TD+gba+9a60G5eJ+AGyGgL2fAX4TOatShmYembz0yNwP/Q
j0JxXs/775USC6jXZ04ldqU80uWK1NnZnJevuLKh6jHTEREfkMrr4bxbz6PHVSQg
c+058LcuRU8DUbHJ0foSiCoJBTR8r5lBkJKxWo3ntGYM5x2zSJUILcH7FwCEk6rp
kFxokgvGBiWKg0eg2V4oQd/b/+QUMISoNtnDQAg0j2Ef6pikFY4ZEqGN88uggyNN
SH9eeU0tUxrA0AtTh8VQ1eyxtiwux41dsHRlwezS5VAE1SR48oMz+3bYit9EvULZ
sihYO0KXfPYoZgnEjM1rzGIxR8KksoKFAtADA94GQzBRjXxvVJq2djvYtqAQw6Nv
WM+HhpvhDftI9NK8PdvSLUghW/IkKe8EJyCYKiTEe5aiOANGcLxrd+3dybw8RioD
gTAYiAbmcTguNK5cj3KzLvCIqEwdhq6RdUSMFdcnVMGU5wjeyJu/MqPJIws6nLNq
Dkk3CP4fbvGxaNAerHbOOGLK0L1wqLVtrUBMoyS4Ay4GhQDu3A1XAmqhXhpjIzW1
8e1iyXTZ/R7oRto9r7Iwpw+gCdNgzznEN14bobs4Ye9v3Dgd8V12NvVVIEIw8uUP
9a/SnGyzg8/3pc8+KI+sIqKkwKHvw4AHnBmVNqJ20Kmmci5Aq8ebw/besLfBaZLS
vf3w3+oFajxbI3zBOoVE6c5lieJf07cEXfnpo8gqVvhpzrwYMrg76Sq3xtNVHxF1
TtF6G/rc1Hiwq9N98PZRmPkEjxTYpBGcNME+QElHHslw1d4JVINCmURtLxqgfLmk
7STbDLUvQ4ksqXsWUjrOoZt2njLUMI9/7uPYiZCN0Lz2Ft2hfkVfhPDAEeKHiNYr
nATAxgdKhwWWcNQyI72xTYbsV/rZO53e1H7cT89YZu3aqvSeJOG10t2/OaTWtnm0
t7nlFmYO23R5++nnlEsbukinWseM1GnSkRKB1ZP7cD1QIQPNSmu34++ZPctlLA/r
8vSvBg1RDyKqHeBEhmpMjpxCv985CKH38j2k3QrrZHpYwEU+Y1p9L5GnyXwNan6I
QSSbKfnyDHFYealNJaJ7gW5yQ/2ookaQgEldBuuTVA3/6CQv8nFiU5yeVs/g2Mhz
uEa394lvea2tQyE/Mf4bAFeBfd3NXSUBxJ1KRVQ+2CGvJppGFWpGsOUdowJtKwWb
fzngYLEqKSGOYNzrzH5+GMrxfPPV/dZQ38/qBquwo43HTB4DsuW9DEDsMHKYGuIC
KFNffxUvAO61VphhVEVUBOUxNqkkK/kb1FF0J4ksz9S9U5Awx1Ox8KThpcww6J8U
nq0zD6po7GnomXq6YMBNFzQ5ihcFv6LaZi92+qDTKcRA3vbtjO/FoZ3Xv7oCNDRh
gBMVby1Wiv5g6peOtzXbItCHZdd27lTxibINViaQDl5uY4ZO7nzJv6Lua8WECOvm
eiOmNetOW4HRhQySQLp2wgwlMuq0Pfpt1BBXUqLHW10HFgktQi9h0D2kd9n+W7dx
VTl9KdPyDw2aYYg2QNx7kpad0ZFEi3fWLNXAIT0xMbXswDlCdgh0MCt5yeObgXPR
tkNKOKgT1G12Amb1rfa32HyMai+DImTKltRtHjnHenA07yR3PehXBuBY16zxfJDm
T56rvUKoKvtsBo1o3tSauflDrj5NwbL2xDhwhiIOvZI5eZrMEFmHksjcTyhjZPiq
9Gvzb7WZr5uAlI1tb6xO2GmCHYfMH2/DqLDFQ6LQ60ZsC90bLVwyCExkA8QCCkgd
0Yb7KpwAwPlhgUHlIqeI1MuhGQ5ojRL0H4nDZBhJOvN4qAVg1GwpyG5r1YGY3phB
qiSYo2ZqG17d9mbX3HN6gtWzhxNbjlEJJoSU53vn3TD0x5CSkt4671yGt+SjOvdN
FbL4oqb4arDr9pwp/9TAhDTFJSWnthsi7ljKAOjnj5QNyVZsEVAXJK/nFTbBG7fR
+ZuoVd4VzT+2gCpQ9uPzJsAE8S5c241MrzrFhWWgkB9lDk3tyr+UVnwtI5PM0D3G
CkMhuw/W+k1j9JxItkn6dgmTXI2H6HEgSpDGt9OGyp4o/fU/fxYZhcK3tQn6DReK
L0CwX1DCBUtbACiserbxxvQTzd0G6gWQt5HOWfWBw8E/Dq1WQ6ujdInNfGfM+vkF
/HVVFsZzXddZFL1K8vPXSUeIJkL4BLLvFRqTdLu0YkhIKcuH/8EBmur38WZBT8DB
PkTKmDtCxgiO+9AfM70fvdJe7zNbJS7MGVPOXRUmN7kRyt+/2mJ+xYSz7Uq/Xlls
Z+38za/V6alkj9How9OLzyx4/fO/awGjcr+4gj2iA9zOSnS21OOcB7VnZthCnA7N
72OdJrOJy4f4kalU3XrFTo75SBabZosI4SSX5k7FYXZrIqoOrrSfLJSYl7uuH72p
nXuiY/t6bTSgObGJUm7IhDarz/jwG7ELuhinsrBU/H2/FGbE06aOPdjejS2RzyWu
dLOHxhaz8QD37BsGkW5dxpuFMti+6L1oDIG7mKW3lwHhlvoF6LklO7WUZeMZIioG
6A/QngcvHTwpcsIaspaMAZLDXFK4w5xFo/9fueYrSucqowf0QWi5u1WR7U3VMsRW
SOMl/RavAxxPWoFzIFH3wGOloXSkoSH7RVoBErX66/2YanAhKmk38azG4h+KUJ4l
qb/196W2BaI3to07gB9vr5n7gTS6T2I34+fOutluiAcC3Ol1L5QBPponagDmiIEQ
Rm3jPEfUAhbj5EniC5F+MUF3xjGc7hgyIc1HI0fa1b0e6h5NycWMqVOIVJ/+FOzK
aFDt7RcE+2PeZCDFGpdr7JV3eJn517DnUIctqiZaEQ3lWn8599NW4oDtfiTXs/uT
QIgSkQdpkBqEBzSg4Lsq+DmcHfJnadABB5cT56K+XUwVS/Bmqh9xwWHHr3l7Wk9d
qBl65Txnk1q68r/U69CApCZEJRG9zdQ3JbKNvjufrw2+rWenAakwW+mt6+qkmTff
cpNrXYqRUOz9xkDDkzsg01y04K6jlE9WaxR1C4XYiNXB7R9SRsAVXv3RJzZDBGiT
UaWKWiHiTasObcdv2lrodxm+hv7SGFinKEEDQYi2+mMK0b5qpZ6IlUpb/2QcNwD6
o5c6cfvP0o9PJr1Pkq34dRh7GJtgM03TWaUBffh6v6oB0aCY/MJoJj+eFDLDvsRx
DF/NbSADyLALVIk2aXSE0Z0nvHyAhNoQCexeS6CdUw/BfKhJ54xhLKD0o94d2wj/
P3RyBIAMwl1fTQkMkqHIEShcMakEBmjcS+dI2XuDrhiTvMqeRFHOkpjA3qA6cGuU
9YR33aebkjAekM6q9EFlauxjTuFh1rCGz8XnkD44qX8J4DjXbTmn4SA2uxD7bwQb
Mx4xNijWLCsAE9hSjZ4BesDBC9L++VPveZKa46iPf2FSA8+bV8I6rDLI1XsRdId5
m4hcI2qRnAA4K0jgCeUYg5XRb8An78shrqrbWRGQUsWPZtKBECeC7JQlEM5iZ/6+
vle1SvOlrAo4uq6AvSgj61KcKBSReDHy/TMnQVs3p6xDUap7XPz3OUhNgJkhY46g
FLMKi3CwUvjgEjk0yHdHjLcSExRolVqvz4TwRHLDL6bNqYog2JZE19uNMkKqRuTz
OsVY3z4HG4gIppIhpPz+8192hiAxZkVbWl/le9udf9w6RpcCkFI0qD6J+/ydscN5
nnxGrg82MU/2dcaae93wQwUu+mJ6i5tTOSRH18zom0J6qh6yOmbxztibdefORmi2
LJvF2KW90yzgcV8LaycjJcIZ4H3wXlHd8y0UKZnjFXy8fvJZ05ih3agwanR6V4gv
ZiauXsC39bCHHnR02mJvWTOY3EXkxqjbM+ZrM8MCN5vfl3ho1Rku8UyWvOkJYoF4
WyWKHlFNhdpNmyXEEQc/GE2bh0KHcMv+EqV2sEqIEgdApl8TvcwTJcPOOYQDwCky
6M4iVjEaS0rCEtG0J/yA2PWeAE/0cphEl81j04c3Wgm8QJ7PcnQccm4dw+fTgbNB
6WVcg2IOBlDv7afCLpsssEsYmcQ5Q5zrs5PzqAoexqHOB88gbDoVepmjwxcXXxA8
99TLGtKkRTOiBRYb9kZIVnqV+mKkDQ6teC5Ip5Z3AMzpjnlbxaJqgBNIpF3YbAT8
Jqo1xdY70RfAnEyKAgcpKODieZT8ywFgZVFyfD0nRT7CoogEB2nESa98Aw7HyAhv
WFXVDiimsu/hbDI+pDd7Oynwf9vaCJ/80Fr0iMMU4lScum0Hc5iGFWkWBjv79JJk
y+ant6I4GNSFLDTXbbVcqSkKiyH0LfoazFjZKJfA4dVu6yllizL/QYs348k9Atx7
c+lG2GFjLi/N59z81E6ML2zUp988OJ/xOZ1v5QOBDBnO83AT3f4T1QXIYEMzRlrK
tN9zITbiKzyariW49Ga35dwcCAIqAahDmzo48ztt7gmbJKoJRMochiZ/FuB936xG
VduMFURcl+uQZ3MxmtdUdfaN/OF5J1AyNBQqmlmVTqMpLNP7m9TWgd/RTlMa+qZO
T8SKyjgPr12L/+bR77l1Kb+2g91meL28VJM0GxmLS6kzAgzfD3inx8HtcEb0VPKO
JFcqumFwN5IpUyu3XWjlbA/8sZcGGH/h4a9ldq3W3vzn9refvCXYLJyxUmOCXrnU
M6ry8Gnv2TEMmi6Tk3dlrJwuSPO/1NBFhIHhv/wAeAk4MG0emn41DHFBRc0IUY+T
jDc74fyMw0hPj0DjPmJYf1Zu1MGJMJxepR0hQS6/p7ZiUD494TSn9GljJccfafYm
FNOO7CPELpar+coZ0Idf6OQG3e4db7zoUz1lVNZo2zbwa0AYH5tol9WAvmrDwet+
9ry97Z7pBjJs5Q2ipeNM4uJKr6Of/HskC0VlvAyoA5R0yV4nLg0iqIwoOj5aPQSL
cGu2bXZm7PRRbhHvS9g2tiqK/g6XiAm7lTif6vBLiU0Y084Wh7VCdknGB59Fjrvo
rZidThCZjfY5yxJ3EpaaIynkR8UKcffk0IeTuaBFiQyft4VolBaL/c1aHeIG7ocu
6xrC6F+LuE1Hp+JaA67slXQRs9IkDkbIpKI5pItDX0tdExh1WksbSM428ume6rdR
ajpz4FiTaJ0mt2pe8zfrzbUd8AsP6QyBTGWmwotvtTgcwR0uzjmTR4E8B69FB3Aw
tiu39YRi0oFI6cm0gDRAcKhle5RVgv3KvtarA2kwFzFNWITuV36mXderA+KHD0To
nyioNc5iTsSgqAfsLJAIb4AqrqsVJ65/eo4rNqgRDT7PILYFjleTwccAFd7s3D2g
nZYzah+IqXw/JUlD1rFEwiTKSU1cimpGLuu4SitpsyTmILeGr7mIZJlxrPJF1Zga
vIPLT1QNMFXC1scH02il9oT4euY5U+irCebT/USi06spkmuycy2cpz00uTGzfbfA
IKUrT503PxGB3DKutzUeTP2D8528oV1H9A8r/ooEAY+4L7H+AEKEmx9/QPbIrIY3
pclabxHXkE8goKJPWEVFMoDE/cuTrmTP9zMbhVw5cdaKTp8QbqjT9/EULcFTUOOL
b5d+fnkpynxJBDJTx5+p0HtiJbNh3N3kOaiPdRHa1lbQth+neTdweypkFvwbVGGB
g/StLUYVY3ok9ANRaOptlRNoGPsyjWT6G1+NdHtgJh5k7coFxJCB+tJl4aF/y6IY
dfABfGgtJq7iJfZy7W2qUnTC9d9l+/XYFD/mUbYN36Y7+woyG20Uktg3whtT+D1k
pMj4RoosbPbpIVBt61GIRt41IhbvuMXQ2M065G0PYusP7um63yMKHfumQKHD35LQ
1DdzCvba+S9AA5oWnyggjlWynHL3wMKfYgj4n/kd8OpD+l1IPYsqmm9P2Bjj+zpt
qx05mhK7Cy71saCIF8KnpeTdgh9bPPqvPwyt/l1GZZlolFTztoeKA3FMwA3XQR0A
6R9SdKSQI8AjYjhAF3rEbd/D5GVa+78q8TD+pPTzd8vzWBuiTGEXs6UmMnB6FrRa
vXTj2A/urReAVCOPv3rtttTbyhPMXzRNDgAwQwzd7Zh3Tvt+V3jDu41hyjmq5IO9
JTW6Z7eT2Cioa1ChxHGcbd/tXYklUGjdMT44CxnZWN5EcTdmbftRiU2OhudYHeEb
YmwAOaKpaTHhttIGHVDI4AfY24m08NRTIu69STVeK8+MHW3ppY+SrbGGhYH+cwqu
Fdp9G/dx387EwJCrJV7e6886rKE2xQGCDBOcgUmy+F0CMmE4HI6E3/1YpgaGGS4q
+1i+VmQtCqCI/W/hpa6wWCac8dl7ZxQbP0wrs3vR1XRZb7I3TgrUqUQrg6K4OaOk
jU1kTNBKGPSqk73aya3ZuHKkK+Dsf3FPsmEXqdwBcFHqejVta0sswx9iuRVFDiGl
6xUF8jYkQA9dwTS1ESCkQWdROADAKUaHw/+misJ4ie5yCaLCrEERFq0u/empo7Sl
ZyPmFZqVWSJE0qJCImWtby2MBscHafXwao65+qbixoETSyXT3hLUw6q0KEfxQubz
4pcQk3owrDtKceLALMnhG+HSHe62at3Z9kwP0vosqq/TuEl1AZYUaGA94HeiGSf6
JaqhfW0tb+vvKAULhSMGnJfVfWOmkEhppmNEHnASpCmJQxWZYuOHF8F/H1jevtD+
uJSm4kLgkT2TZsiS1vwNYhNraiqU99X/u0fcSDi/7o1SDUwcpWcOVwAt2aO0L7mt
kTNmi5EoqC1dNIk6eIvqgw1GriGJUA6h2R1z7j72wa3tRNdrBv/s2YS6zJnpcefH
BSGSgh2/Po5X50zrfZdjWL0GjhcXVEajtRvbuFItJtYHsRMFYtqZdha3sw+WjK2l
HwJnwe6595W5Yq1y46sE8K4+oc6h29Cd0ZsFe6vBu4jdw5o6Am/8lrdZCB9GOgEH
SfkTQcdrWwt4JEVj2OwimOQUrvLjzSmu4xxTSP0gxdP5ghx0q8Wf0UBtiNAByyTy
l3XCbISjN7okiCqmEJWFqhrd5zbenbV7A7rDQiPDwtcFur6YruT9R+kI6Y1UNfdh
CGXwHnirOksRhs8R/v82xEXrAweO9OuJ52osgni9ba/mY9QR73s3iTrNcI7IZmtP
KWUSe8ltTxjdRRblA9L5PzhabmrT8hCRjBUUk31nyOg2mnZqnBYgukumJPM7dTMc
PnlpOUbn0CR3xgI+BM2sB9Z5zLNGYogK2D/SG5F0dWqt9QP9++JKoH+M0OQPabvA
jiw/18PD/VRlYGNRxP+rJWmof9AS3I8USNUEDjIQ7lE55P/JcwHBenz86wiieblD
hjGc7N1YCFaaXmVV3/AVUlIcmEsgv2RwsTy1AZaYzN/QcVnlQ0VZ0prsVdlxztIN
nMM2+JSpECnGdY+EXPPYvcX/DIcBsLUCwKvz+aV4KNFFGu/ciDXnWGYeP5muvy/W
12oKOwuDFN96fd325zJu7jz6yShcz6Oqlbeadmvhkj6qksgZ0mPY7rjmoWAdqySo
iu+/tXFKFmujcHfIr7ca9c/qGaVWVS1pEXwMe0NvdfM/C1YGAVfcM/kFA4b4DCkE
OeRogmD8zhKRHzMAWMS0ZXEEs8Zk2+3fnjn8OY+FiZzOuLw/2dkCO8dcLS6ywY9/
po8twEjKH5Thj4t5+6zJilt4E8dard7mg+OoMFAPih5B50rpuEPRPzdemZxbn2la
wLTy3KyAgWzYa1m6x4Ns8piM93selQZCVLfbS5t/JmRrS08J3Z+ClLDu35VS55c6
a9QNiadrCgsHmrRkuHasXHFulN8m74GmydXs6VTR1Vn5TUAFo5vP1z0lt+UuLF08
U2ouJTQJdQ+Yd9wwDmNw3LEEMeo/GPZSq+9Pju85hrBVHXs2HRbinBzIUhx1ZHnT
vhbTZj4K5je7dahggQe6rLesimNxx7Yvi0FIRY2BPfejo0wqN+BAVP01PppnDKv3
mq1SSac+WWHhqRooMs/Fq+oveWDWinkoZPu4tsqsjN6YCkI04utWUX1H7+diHjd3
nTcTOne0By4o3QGgzEsxjTWjk0CDZ9R0S+TSsSbEZJvXCi4Q08jzX0ZE6UUXV6Si
gW2JwEFMQa1R9s8aguCQVYEVfceMFVE7m1wIZ06RGOuJ9OHA4VBWYd0PTmj+c3I6
gBlE11INmuRbUwJ6djYgIRJ1a3mr9LOlxoTAqabi5+wP5L6a7lTOK3l/N3TnSMfo
kH7Btd1k5bFgEVE7ql1OLGImenxvUWdQ43i+nTvLqFNtpoMxYm9vN2Oq6H5dmdDb
d2I4Ye9fK5+wpujS+abMSNR0bLt4qii1QivQdI6vbhVMTHIUxz+VvZxEe/p1wuWP
kkmVPl/Hp5RJdYrNJuFXm7kBPddbuKeEC6jPg8sarMCR8P17dWfqUgsegs6JhwFu
6wEFBXdQsmeztG26//xegNOwknReMssfueYXIOv258rZvx6/sRiU+KQi/dkP15gb
L0f5wlkW95Vpy73E0rhYFmkciGz6vdy8YJZ9INVqOzScX53SiKIniI9A768LHZbI
31s1gxaEUZFRt5p9E0T2E1uWhoWKhJmAW+gW5dFzvlQOL57hPRBgGTdOEnoanYdi
sIKs72ml/5zakOMFvR1IbdRSgINSItdm8I1M7zhNfr+9VAbxTVv6ZhSW4Yb9fluB
vWGF9X2iBfewkS/ZyzJm/cJYvyC97KQZK7Cfum+mOEXDfgKMIFmOpE0m0qj1QLan
pkTk+cSEfwI6IPIQPPrwH6F5blEQFsf+m/6GKNDhC1eikF+IzCTtNUTnkirm+FMO
c2mOPYAvUNRgk5dW+5b0l1CE0rgWvOOzqcAGRAaYnmUI5807iEK5c891R8Lan0VS
jjvMbDA6lH9lIUdKWMz7sSr/hbzajkCRE+9n9K/qvaUMhnWtANAV5hKfLlHO9HhU
AUbTQgX/qejRNmeTMDtd0cicrhVWcotcsekeC6GlJITancbd1nVc1dWLBgf4qWn5
9Wm9xbFY0+hjly8xtKm5TG8LNxJGt0zgQiPa4FcEJCBRG60h2naDQprTZrIOaPTc
X+uS6AZKCl6D1U8ZHe/W1dGGzdeo0yJiF02NJDh7kViRBWPICAlgGTT09Bua9Tmh
6u+hR/2tF1GIt1qRaX838MBNt9sUzhaoUk6Nn+J1hY7Foecez5uSzEKYMJuiLWIt
Xp3b8WBbUb7n7uUwPzCthnNB4m15woavoj35Nc1XinKvjpyPH3kkXktYgnD769gj
lUpE9e854O8JohT8muUm628jPkwpmxvR/CrPOGuexubNum5oW7oIgbEEr4qOTuTd
yE9vHA41AXxRNr4qFQ3nQMuAeBG2yvfaGwA6/Gi27j8ZLWrOfnhdo7DGJKlPxbPk
51HFIG/zdCiLcgCXYLTDKODw8dG2IBqbvSfPIF0/xHMpWPvTYF059rJDLilKpoFb
ukrXN6LiD2O6vWQl4/66mcUC12nNUgUJFkeZ06bgVNjSVQEVWz0MsSQ26lUQZcMi
XXAwjpsLOhbTz55SfSLxWR5QPvkggpDLexKYjktbSCqAGhboymGWo0w21X2naAsG
fOLzTzhYGw6hbsopMXraGrZpW7ebcwXczL5VSvxM0w6wsXOcfh3pz9SjA1bUjPuy
7mj86itUYClDFUQRvcEfSVRPbNmY5Tjl/MvWRPKgEUm0nr2L4BivnWgdSrugC8gd
63X/Vt4+CX9qmA/UEqehjd94JItY62EGaTm+2DfgtUR+SW1c8CPWSyxei1/DYDQ6
06Wm6R5bO31Dq0rcgMI1TS5Tk+7Cc0LrweCAjrRz75uPRZrXyn1BLAxyEp1GXMvv
qr9klkKvkSGfnxQE6GyWyY11Fz6WYH7OTsHMOHtsMMAK9+qsLY/6qK3GYrUP2jxS
r5odOLtgWxa0oqUEUQljDOMKP01EOyt8xViK0i6lGVgvLC0ReiSH/80VzMjgPwbw
BKZqxTOsArGcwQv/NJCW8/xrvWUcUR25s39lcL6jfzuK6R5/gsxQ6px3AAeCvxCN
HJ6BxkCwey8F1Nlgan9LOZHdTW7Sd1Uq2/CEeTCWMZdBl1awObSb5Cxt73odrKHd
CJDl83tHCShUmOhDmmPoW94EdszzxC2fyNHpNFP2Xw1AyBzRZc5Qv9jiXaksZEEN
A3w3llI4YUg5L03QjveYAMCUyfIk18CYW9xl12ThUHXurxgc4HW8rZtlmuBfIoWi
7nBVWyCFndPUTuCLc/AA3OwcqsyhInN0bKp6zh/jarirzbatByJyvMOM6w+hh3jI
1IHrEIA40fnTXHjlPIVQ83Ctuy0L3ZZ7vJ/LdKAwNc9LrVsVU218auj+sFkR8Tsk
0GmmQhlEv8fsGiVX11YNdy9Y3rx0UTSK/Arq1Brh6wV21nSkkQYsd1E9OOkS4mie
jLnEmhDaUVOVAJfKPJVQw32Ejv9b5f06nkvYQr60kDBVoKW0m2GDk31QbXW99EC0
hurMHYFsMaf1VUxgQCHCSjIk3UwDlfcWYayQeH7uecLTMVnHQBMMWVnORR6fxMdo
Y1RhE3H5hOqsxlm8mjXTxqziXAUzsDTH40ZAC9SThzxSCypLzdx5kvRMEP3Ef76I
jtaF4pr7PTqicP2F6OY6RUBnA+QfwRyMPxcqll8QTTY5NGtnwDhL6PChDIMrd9VK
yetcDh88sb5YkCycKkk0oHnvGvrkifZfx6ew2y4yCnBhe5fEnBXehKcZEaCAaJTr
GQRfFQZhLYU7PMQpuyDltZRyTETVATTwZ6prtFf+aS+UukijDR6DXAS1KnKvHFjB
vGXKfK0/ildKCHznKuSoCyJEyGBD+bIEVcgudCDUVxubuxKqc4uFLjxlU64wgzwV
J8UmnTad49M6AL+JlrO2FkMAmcf+LtCw5+PJXBUPyOQ+SqYdXg3MdPa4LxdWnySJ
TQLBzwMbG5KKHQildisoaSI2BWzDXIwZSquEqK3z/vB7V637o/13Xw5kft67MJ9W
f/uOtwugtGICC4QzC/0IouTCF0ypkN8udzpwSHdKm4JS7xXreYNj6WXRz92k083U
HPJbhDsgMjQAEhHuz6fy5sejfi9yHTpddqYYd9Z0nNEYUaPKgq+8PTnsDQB8Yjsz
N3djMx5xyc+YzIieMxOsd0HNpYSS/P0dG+bF5/yqqdk3+iPocqUiSUqbH5CsXnZL
mfimJ5ByckeQDbpLSqV96Cd0Q/umckvrL5pWJWzd+ocZmKVJsJldKYqq8qMA6Fr1
BbdPjbxSjmFihoexITwa6HXa5wGeIO260Bzw8jWB09PGuQasDsKvNRYC54sWSONg
NPlJnL+5KYBIwL8YfcrHMFsjk8HpNsDDxSuddmgSfoqWfd/jEa8CnzfzE36MQ8WW
U0gjXfm98VttdiwG0uLgJu0sNTgdi9pNkal93jWTK3P27z58Wqz+Anb+LSSlegrK
wd3J9xrpSzekMsdrbwmRz8qR/cQDo8rhb6J1IOubbLXex39g2IFqTtkLnpzCvpbT
ctF28Vxy2j9YFCaNJkOBUmGvMB2i6bTNFnTbAjxRrIM8LE1MNfKxZ7DoDtIrHvpk
4Nm6UhyGedC9M2ct0Xt56NjHwa+lolyqT6z83FXS0IVEEspGK4qBfVfFWAahBDrH
eP3nO0JYJXZBnpgyyRLtMN5LnKYYQ8bfyZTcBAG2tAEf5BQR3FFLdeiTN9r+4Azk
FozvtIM4CZyuo9McsHDG0cHIOdkpCy2ZVcjA57EulwkNHyUWSIlEGRiUpj57A+5B
EBpTeTPpmNLJFBrhUaXOTm2+nud3kIy22UTn4yHPgU2wQfdTQ8m1GMSdijCK16rp
ghryH3hHVxgLIqHTMBRstd0vkiTX3rCH3cQ/+y+SAbGc081Emlkn0rSUgbJZ0+9W
iV3NZoW+aGqxQKR++2zbGT0V9qU6G/sJC/XSdWCDOrFRiEPXdptgUacBTd7M/yms
gDaEN/8d0aVQ9D5Ab0FS36KMdlRCA9pCqIu/7dEYDyB7FV15ZV1QUM9lYS3CejMP
YdIZRP7ryucKdEDa3tBa+Lg93QxMV3eKljjf1P12yfvcUBea7UGP61ULsGWLCyF+
0BhlYfgFmnnp0bHZ8JFBlF1TwqBrvUd0VieMLIfojStN+WCuQAX8EF4g5NTrtecx
PeIGr5JJSiKinjM6hcr3WdJmFLVf2O0Xfg/490atf9GvKwh4Jjn/HbHB5sjSpV2P
7Mgj35RuJFpFwekxPGQzKjlSZfzY06pvAbF7vKDgxuoe1hcfuQBsZb2iPFmBppPR
JPYaj3P88TUkz4yx3aezxK32PkGY7+aT/lRCanFCSBPGpq/2c1cNGgJiQoAJ9kgv
5qPNuu1/p+YpZ1idolmXO+3bAX5TX3AsziXBLhoGnMF2tEFcbohtSmzYwLN32N6o
YiuV02CkuFVYVzJCT+urUsn42aarRJEeOJWHCbEZHl9OZ/64MyRzc1Q/VP0K6Gjb
YjebXK0GxSoOzXmtroxieYUxmrp1TwCbQwf6Q3B2R5UjGy0FT+hCrQT8Y/iRdg4Y
3hvAvHga0Bbn3pGTqb/fxkdbXizSE2vJ1Q/xPF0ATqGYhCLjy5JRO4TBhIManUnj
Zj45neJlAMWatmN/CRLJarWjo7B6QKTLTP867B1Mek5CZ4vqpZ4bBeBnwIh+TcT+
AhdAtNztTXrqz95GreK2RV1Dge/jHuv61XiewD53risvv576bBTPcLlAw/fS+xez
3mvXJE9c35nq0w3XiK7FEJxU31ePMWdHKoeaAX/9MM6XaIp29xJsKeeeTD55Vbh4
78pej9sgRDRckehjFzLpep3FELSiqNbD3BMLwBVxITL4N0NzeH95xpLoQl49qWFL
iHBG64Hv3PzctXydwjNSRsizQqbmR73shh/ZH9Gdws5Hc4GINDXJrTBPD1qPrAey
Ht8dU6GonNaED6tamQkK2PJd1a7GRmgSCjvX/RFu1aTiuEyEv0kiPBuOXpR/UxiG
pcAguYhUJ1/YmplsNsNSMAA3HDm65uszTCk51lXsQcmk7LHtvLep+boH8L6tApa4
OI+rp4hQMle2h+CluMIkKZ4f9RgTWTx66o6sTZ3ahhenlCdmU2eVB8/lpy6NqWj5
x7nLKqVzmwMQE56ExnSi9WbNdPv4rFHRqGWEDrR9Oe0gbOkwAA31/ys4lFtTD3Jx
qOXaGzbBAlmrGJwDBsXhF6Aa9ge3mAY4dFXDT8NRZHM9OtxNABZ/SDUcc4C/0vg4
KZkYC3vlpD0VJy8OTnahIZ/+OwicUK2nFYfK5dPV5IC/8sT6w82KmqIc/DmP7Rzg
OjRyv0CsufKaCtb4OlH+NSaukc/S/wgOfJKVGbWYIl/cH6Dhl/781BkbX6sam0aJ
xEH7zzUv8Ghz+BTA11ywitmP8nmXcL9vTlJzO8yNHgKP1r2C3tLWR1GIwXDgYjdd
eNpRHH56YOntaTcdpbChXs+wEchCcMAWoNiPaHE8ua+Uhgbc7qe5KgAE/iW1Fq4Y
KYNd/amAoXp7pojkK730sNFWtU/OabOhf9C64npH2dAPm6BAOZ9fefqE5UPTF5VJ
WllAGLGvg9k4nncUzbCDvHBkaaWQsFSRXwGavHPpFd3YiO5PMC6jloFfqUb0Z0QJ
QPI69YSZVN1nuV0st1Go6szBIMyPGRFpfz3Bn03gI8XEnQc0owYpQUDbmqYxTEBw
Td1XFy1iPWN2idEM3SUwsYxn17jc0/4s0Lm8n10ApVj7dRgCCIJsGqGyB2NqL/tf
S+cOZ9wtCa1Pf9K0JnuiRq9f7CxvNzPojfK52tegaUFGiL8nj8AGAz5cqDHjx4jI
B52SzXaKpbxzDTY9NRmOOguHPshPgI53Th3OLykTdAAUejFS5Judstae7gIxJ7be
+9q0Fml8EvILveF4im9N7tO4Scp/azhBmnNVnPJALZRVMCx66coxYeh+E9K12Utu
QHqN0MRDFQvpJrNyVjOPWlJwHGEZMy20XdUr20fod6TgxOGTAwRbgzpPTrN2iwjO
MCI8rupKQGARxta7pIJR35LMIjCjmHliRQaO7pHqcRJMiA371kkle6MepJGCzvlc
PytDk71sMzQf7CHVsosDnD//E0rXUC1hlFDQfhiyt8PcXVDfhefXtx3ruz9eestM
WWw5RAsf+20casy9O2RBvu7KhIoXn75ZvsjWsujeiAkd1gPHL054ouAcxydGN+nT
i1SfI18Apo0ztyeAeJjEsBjBrP8yG+iRJdcaK6620ZYVl5nMx84HUC4TFrKBt5tz
TW+IuhPGPQnpP6ed8SgfxJGc3l6ZAbJKPb2h+53vn86fNqbhoil96qRxfDbq+Fx1
RaCEkqywXh1AyIx2sOpE8zlnTTWVq7uU/YW2ly2PzPiwr4S5cFBI9AKU+SqSI+0j
VUj3PCEu3vHBYZhmMLwDvEv48TMB8kjCmQqN6bHRDTo28Ed7muChbM+iMX/fVe0B
Sgeqp6tW9OoUZkkFMonS6dW/5Lcc4mANRspK7k/UmpAiXDsw6XSp/sT10xlX03Wq
RK4Vw9DxSUHy+hUWHOA2S7vJo6kPjYgxrWuLuLXEK275rD4ogLhfWwIo//e6CsFK
eVJp23jEAu7NOK2zx/Jv1f0DZqZauHs5y4GRKyShq1SRlVeaozs2dqql7wvLqCkF
hWjqOHDo3YIR4OKPO6Ufwz//egx2+thpwMvvKs7kQs/xiAjhA4v+KmhH0HqIX25F
/FJrv4OLOyZT/swnr5gMx3YYqN2r91M7gsyX3eFdfVvRiCf1zVYPHbW8/xYpu6Cz
C4C8yvGAEcxoVTB/sYoEZiRTbTgskYvkeFDd7Swoogxghcth+881R5R9CwM7yVMm
JffR+CGaYbeX35bFl4/iiCW4OTYKnd67YwMp+B+wxx2oGB1qnGIGn/n9sqS7zWGF
61o6RbpmI3REv8H3D8XtkAOpf4b04a2eaWNS9X6rbY5ZQS0FpGIF/o/t0SxjuX4v
Xs8dsrTv/Ei5gOjMUUtJ1V5sy6jfw6VDs74G+gKcCSx6rNYPDFRvX5ElL3NGeM7c
k7LWHzltDw7lDWChiTlGzQp9tktBILErsXFPt6T/+qLMtozNSoCRst6z1mrnjZww
jmsdZvLgXIzqtr/xPNB0QnUMr9VM40Hqn2ljNGmtUG73fF+/vJ7B03XddOUN7Vp4
cF6i7/MIlAB5IYxH9yvTCeRYWQrqKCN3ZbemwGbFJDpiRFAzp21jh6kgIUOWfNWL
fQyhr9E8gmkIHiM0+DC3/VaKD9+YXgzYaKZ+hAHJjMgcA8zhiX6OTJtf8JaKCg69
KOMQUItRlU2bI7X8b4J+2TGz5VWHfFmSjrqyDGs801DYhrGtk9jl6BfEQm86y6Nb
40R06XS/n4Ze4JUYHH1/9x8V5sQ42GnNK7PpS5Xwe0P0pvgG2Ng23cw0zU4ygpC7
JMLw+fNYIOCGTwXT8KR/1T8GN7bLe8zMQ4ytE3M1pG7GyOGNsxr++vLYBf3JpnZh
5H7RiFt96EjsCADIeWvOjsnSZ8NAz5WggrJ8/EfqdzJNlribJH8BJIWzGusAamVm
2DgtJ9gSZo//H960+OhWmyhpIqTtZE+dVQ8H0biMMknuEtNoiTwVEPRoSWFle1q8
anIuUFyFyJiXea2y7dpW1Rc7GvSh/WYvO6p/XxhLntk6aCMxWDNmJQISEoxAaTds
MkUldrkUxAZpZBBbuSyDqCZNelk7Q46UEFhzfCSjJFb7ipU/06EgRCZ8afqVQxS5
I67Z9BmvYcm+Hz2lgDmwkn7NXn6Ea9+v0Jf1RYq/DtsoQD6Q/5ewWNdoiknszY3m
P/aC1yd8WFc72m647n2qTOMYH8OaHmFTkpjRYJeQZrwrxg0tIijCTtdYFMq4Q/rS
ClFAdbPDnGmS+JoG6/phbhe+UqGaz9ElUIUmlr9SRpgjxWjPDaqbbNmC1Vgz6hRG
/QeekS4WtE6Z+OjNUyCbJgblK933h7J1/1kKOJXP6hhDUcXA7NJG6iOa53iiuQY5
zzFkxeOqGWYHKxdtnbF0FWsJpdBmdarCEEngOvA4MqZ33uJswo+XwiCJXKGNG6sJ
0/mpg0V7GJ28c2WyZWUZdj6Hbdjgf6tlGvYQvmxUs836pxAUaIicsHmrfutwxI3H
r/0r1mYFJr9487SQAGtqdJeGT8Mifcz+z59PyOk3OtHnHs4JKlBi/vXt/iJo9lEp
CihEF1ZJEUdu+VCOTPj/7h6xwS4V96/svjxVk2oRwipvgR2cI/b9gJbg/MtsVkQy
asp0Ok4k3JagVWkgDTlmAo/0hHFKG+u1d9NA24H4X1yA5mABZaQeCSEhBGKkHbs4
dBu44IdFTLeFENymTD+1U0YYxZzi+3BE2oypGWLSU6rjfMc3/swt3TSLJxlXwuWY
/zUfjiI7HIOuvO7uznF+Y6jtewga2mS+07c8lzFTlnG8fQvWWxviYRsdhRog4GHR
SHV1veM2p1wkYhoktzM8rY4aKhvb5mgzE2QJ7e2h2VX19CVo8OdWNhr2rpbVvMKM
LfmhCHQmEVap+OG88ZUX/ESbHA/BejrMtpCpNJWtzfXSTkAuZRyYniIUHTDMGZQ+
oQ9sJ4/CXXfFoG3E6K/PuJaZwV+9+KUiDon61GivOp6wYlcFDNqH/U3Px6rE8Nly
FHjq/6tpBMGvZNwd3mihvdi+alqT2tCkaz/NN8fqAGKxRY3+U3ppJrb/4az5jse1
fUgMhZ+P3dJzFib7K6IhkqD7kzXInSUxi02k5K8pNmiAwI2kf/1hCOfqorWgW8Mx
acBCq0bmf3RMX/rOz2g+IMDTkwxrhLpDY2dS6v1L9rem3Yxf4aaKBy6e847/2046
RDYIzL3ZCDnRxtPWluSE0PaicF5Dd4zudvNr0+D+CcV6nruAXM9Dvf8ougD6apAL
I1XszxXWEom4pxsUBxn/kQDISgHaBiX8JPF3LBa3FswQL4UAk7Ya1niW91iQLwTb
qqAmVtBYhH+pS8NcuKfMIl7jw6vNb59QASPd32Y+wsPZ0RPOgdaOK1l1RhA6g/tP
CpEXOl6wFZbXm4rNpDZps83gkw2nCLsxyKUVnm5N0eGuk6cqtxxv7ktIBBe0MSXF
lAcjY33Mij6NtMoU8tUvan6/NySZjpm+rFwAXG6SXAEolH6KtAnBSSoY8Iu9gKx6
5nNsN2bL+nFg4JNa76ssoj+0VINsr2MywIUDVinMUH1ZiUxM57mnwbCkvBL2u90V
sB/goUzjAZqP4yAoba86PdcDtQGVT9KFEaP1h/pGTYiKZLKMqAxDFahQ1nbsyZEO
ONS/j2G992ieTnZdCHfVNFN5K1qPyPtzckED5ozcVLcBBzdA4Rn0a97UL772hHsl
MqQGiE/s76dW2f2a4kOrxL9Y2xru7C1uRQZeEDlPOiC5kHTo/oquTp4/W3Y5S1Bi
gDdxUEdts9CszoJu3vldwnp1xx3zZjyqMqMyrYrTTOfSmTv3thk8EyyC/IZ60cvp
5MU4yEQvDl91bz0OJw0Y2MqrQXhNH/ENhZeUlxpU9FbsKhUWINwiafGfPdQ4xjl0
tKXcsg+CY8+rV/IisjpD84ZykCyCp0KKxjpH6v2D/XXTIi3JPqXppHHdQR/o3tQt
KOLhrfztLiliaD9irfLxVcEffKjou6cjMcTGqa0TGZyoR2VjHFr442UklwrjsenY
xKY6pgWPUtFNu86MCXJtNOMCZUWaAtK3FlCci9o4ZTk3oPlq0DY+qcboM0McHnYu
VB4gJ4mPqXYBMs+GfHTJT164diJdrMnWXyZPM4UqsC8LIJYiV+SI9Yis8tWDczmt
M6Xzj4T7mYqxqkzIxScgv74SMnp64ISwg/FtSPx62mKEp1V5RDKZ17XZTwqHcpLq
W6QFgiWOjaiC4h7CewfKqKkTW2Pu8t1R2/P3PP7u0V57VbJiyPCxKLnX5qOy8rS8
KxoImM3gtkGks+vDehTKe2C2XXcPMAd3kPgfL6x0IVf0guVGZm8AjKSePxaz3Eye
35ZMWPX81osuxoo2GiMQTvgT/yWWeMbr8V+u4qySOxHGFAC2OMv5JUwvt6FN+vVi
quszjiFVcdPBx7vxRKgBxthMRZXkXcs8HbkA5S17d9t3i4Plr9tdE2wLZmFKqHPf
qHfJKcxjqZaFh0ChRvPKhyy9RhwWDXYqIw6dvatink4GnscHTrwoppz28MB74qL1
mVXG41/Cig/XhgO6Nq6EO60vKWpelDzFvgRwx1lHDkeBjuunGxFQthOpcUjM9DFP
4dcd6GV9B8J+n21+pJ8P0uUHUAQ2SGeKFrfJFPgApy1YRxm8+RieNEWixlcF4DXS
z/a1VzT4P+I326QDIlMsdJjJ4g5I4FaX3IsHULh04slAqaKmaHGndc+Z7yS0pH0b
5T8hG2Fc/0xcAZq3kbQhOBQj2ms5hYLaOEkn5WD5/9gkVuxowc6pNqKA0spi84Uz
UhJVmCWPCfyMEs8M/AVUTwdrLqi2z4+CsH8rLsysaBaxaM2Svq3MoMIRtwXYOPMI
pW6VNRmUO8whMPtGG5NWGtEewM8Y/bpBI5ruqUnJDxTyRJYL+YWzrbMc17THQ1II
cFV/o0IG0T8QTGA4UdP3eTT0+y+4O++Fa1XMyutRyuashr3YcxTHR3DszL1z9DTE
OrwheCKgiV7x7jdKAzFh7aR6OIAtxcJrhp86xuTX0+eemjIAMPnJslZBgHL/fVHj
O2tAjsJGQOfR9OVvbtMNdszGs/cpbsPmkw8txFmuqt/viRL9rzPOf05uL8A2GNbB
hd7FjZOQDyadIhjN0XZIPk71RrR8ORL29SQNqLBIzeGRSxcQnwYYfx9WAQ2UCA86
WXAy4qyWvjsmImEWRlnx2jvmqrU4GNXzcue+FwsPcJbHYg/xt7tZGEyicbcAGf54
YVtHBJ74sDngrki5werh1zZseTBdVVVxX+nEmyPuc2FUIdPaa2o13ugG4OmnEHVe
lxtVOFlEqUSFjDD7iSFpFmuaoIMmkxE8PtrGZZGsKkyjNdck2VY1YEgZoJTmw5Cq
5f9MAq/ZkU3wNd6eSZe+srtZfV4EbgjWeTst8XZ8+A1cOWXoURDdGUIpTypD4uKU
dfYkrFosH1SRZa00UC7fNqQR9n04psTxY8jZyr1nCR4Ktxdu0K+USA+1NdNg/VbN
80/C1SgKWhpoEf5yfNSnpOGEH3FDjgeN9n+HBBO9y7/gGcBi1+jkrwXJjCIp/JbM
Rr9+nyZ17vrVGl88CM/Z5bWhdAZNgyOKwr3JBRXe1HB7M9nRYKoEeYLPNc0HwduG
Fj4WEz8b9Rcqtz362FMO++ceIcDpsXDXn9Oy+d89VghYDIgjBCOU4zjE0hhHwedp
KLa7iT5ehdTKjIGB11cT6HoPHRUukdbroNXUYLJwoKu/PxZFEKCX1qwErS84n9A2
vq8D6lakonTjlskC1Co8b5NxbRBcnSSNtz1525NRP/Mno1YtOzN2jYZ2gUPJHYdZ
p0CSsqag6yHS495J99LUZV6eBp6NwSCjpSovGUGRHrXPt2OoW+RiF5a9h3HiUiuv
12eV67puvPnjAZrDJ33bAASyI121k5c5HG36XnUMkGC/bLejTx9R2GzPOIkJ5b8+
XsBLxNe1Qfg2yBDy1u2/VzQh808Ui3lKvJyy7/rDUs+K3EN1mlJXRnlFLpH1k2Un
vWoviAEN8t6rplcQImor/NkaR1syx4Za/FCczJoYr30KcDAOnDykyMjOV+sLVbZe
rOIANbU6K/413XXJ0vhGEm7eyfS0E0V7D+I9WttxxkDkI6bpuNifDXRmBpvkCJwq
M8AeVQ9u/MtP2s9raasYi6UHrkI59cJjIje2oaMfBjtZ8SR9dtXWVCmZ7felATGg
qGOfANEwBfNwsSmxRGeii5fyB7NgRQJz8sFa1VyzppEaHufLlVBsTg6WY5fKWj8X
ilIqpAL2XfqA2v8PlbYIAOhpbt0q/KX4oNgetcckqlLxCi+Zu33oo5mfjbvIqihe
ACHy1MFMc1oKyV++oYVyI8gQPWStZq7vCf8hand3BBSmFTxdZ62vClj+Rdigbpt2
LmXvo+VWd8xrCeDh93Z2ilz6448r7nyeU/t8MNDHe51ryPdpNpRiGHzPIO1VIJ7d
ooFeJUhyx5xEcluaqzmQaWzdP/2rwfXk1uvyzk8YIR2UIts7QLsEzgiWeM5LF5IU
U3iOBXnuU4AH8IvM9G+ENlvm5V345ulRk2ItrLgJ9fe5DM5EnnHBt6sE29vfavlH
ox+wPmUuWlECviu8M3LEUtAiATEu9o4InJW/2CaQF5j7s/wY8+QBSCcGktD2Yuk1
Bi4RWzEJfPdK8TpvU2u+ijRJdAeJImvnJBjtZnLHOtZaOoEJG3jd4I+Jz/FQafXC
F/yaRWZk/U6oTh4pJV8ByANkiFNd1+C+SA815hSAVDfdm1AoxfJYWY8XRuS3U3BB
gbeTUbYWQ1xiwadr0QFBgA==
`pragma protect end_protected
