// Copyright (c) 2013-2016 Bluespec, Inc.  All rights reserved.
// $Revision$
// $Date$

package Readback;

// -------------------------

import ReadbackDefines::*;

// Abstracted from link
import LuminaServer::*;
import SemuServer::*;
import LuminaPlusServer::*;

// Specific links
import JtagLumina::*;
import SceMiLumina::*;
import SceMiSemu::*;

// Obsoleted by the above
//import JtagReadback::*;
//import SceMiReadback::*;

// Not yet converted to the new abstractions
import SceMiReadbackSSI::*;

// -------------------------

export ReadbackDefines::*;

export LuminaServer::*;
export SemuServer::*;
export LuminaPlusServer::*;

export JtagLumina::*;
export SceMiLumina::*;
export SceMiSemu::*;

//export JtagReadback::*;
//export SceMiReadback::*;

export SceMiReadbackSSI::*;

// -------------------------

endpackage
