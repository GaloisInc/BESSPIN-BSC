////////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2018  Bluespec, Inc.   ALL RIGHTS RESERVED.
////////////////////////////////////////////////////////////////////////////////
//  Filename      : Intel.bsv
//  Description   : Intel board specific libraries
////////////////////////////////////////////////////////////////////////////////
package Intel;

import Arria10PCIE ::*;
import ArriaBVI    ::*;

export Arria10PCIE ::*;
export ArriaBVI    ::*;

endpackage
