// Copyright (c) 2008- 2011 Bluespec, Inc.  All rights reserved.

package Power;

import PowerContext::*;
import PowerPrimitives::*;
import PowerManagement::*;

export PowerContext::*;
export PowerPrimitives::*;
export PowerManagement::*;

endpackage
