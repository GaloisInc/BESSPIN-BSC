`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TkdHIXKu0nk/D2btNzb8I6ImfhTsxZDFLzfj6mKN8BIcT4AZqx7PzaOuGQek4Oyc
gW+Hi89Wt9dCGoYNbxwTtHe2kFv3wXk6nuVD9yxZlmt0kO3b/gLe+nmYq+bNWqvt
qOoeuJyY0NLPND1Uhyo0KGeiIPzECofwgh2K+IOG8Bw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2992)
kLRvW/9+F2azbak0ZEgOP2EENBEmJTNWhAKN8cvL1qtz/xFVYxNEKAU1rAzYDJ+v
UZrW3WdSCIX0ROl0cn2A7n9EUrLSI16XfLlzeW9zq8LWGtTUCTiQtpE18qTv5n8J
dLtMwvfj5tUzoRkxfM2VbrwUu10xN7IY7y/QCb2aVBB5tqugBOo2aFI6dYUnO8L7
1orsUVM5P+MiSKjbyJEs9kQz97zh3Cg+eSxQwpf11UH4U+RKGU/GSDJWa4Y2C1NN
WDnphDB4ebqCtG2AhqHg2Wv156EWVn5NZKWCIwYNXTXunSdggw/GHPlDTDI0bRW3
sm4JOtqAHY5ldaWth2YhVFjpG5D7qUXQmJUj0wMDaQi0yPtDAIoc/kH7dTE85W0M
SqPkWGAo4IpMwEOOTFllGzMNm/mJBg2ufh8xVKtb/y+gp6pwcNhbg1YdE8mCWj7u
8XLpYGKUlSwcKJXihfRy3ppkv07SsGoxQqX/6fmx2ckeHzT0asC2UeaVTWtvANdN
PgejEh11mukQXgbX5/9fcY3EwcuAAPTuQIVibK6bWdJGw8jtbzxQlL4hivq8/iVp
EiOtOQNnuM2ZqkwvtYNG8Ts6CSdAGyTO7Wo4Vh45eZ7QkdZATF6yMyLoDQerOu+d
vBkFeOdQC7GdpdusD969XXgu2sgfeDfOU5ZaGw1VwEE4vkBTAQGq9m7cd2kZXw+s
3tiCUMK8jRi5tFc4EWb9+cxBTDudvxDf4hXm3Wbe+lNuWpdzuP3iWiqcN7oB9HrT
YGoKEY7k8nd/p7O5YFvbeXbVlcVNoyxwwShc93u3iHxokqFoGYreb8zhtoPqHs2x
+RZDBxNoXuCGQK2HaPGFYF7VEuARL+mAj6bWYCVFARQ8gJUVHUN1xk8/SMpbmwlZ
rCmzeLp/bA+ipyZ+cwp3ru6ElgqZ8v+JhY3ThR4KpMmzSqMmmh7BRRMEkmHlvorr
8EUsGKvTRTa8OycRG5gZUoNwvq++NnLnA8SpORx/s5nz/d1FHzjrSFaNccpZ41n6
GR/6xnVS2Yw005CS7tFt4gAb3wY4ldNVJKQvn495XKN6E/8K5KRoTLJzh6shX+tw
ZtUC2AAOar02bzmVozqaOs/t/kBSUVlI7RBNTNgL9YiPpfBn6ZjxcNzV8vV9bRAy
NVWWo1E10WbK/MFB0YQpdmFtBrWWhdWzjENnbYvEWnYI+2uDCWlFIf9tPUHcj8Ei
8w4j+HgJ9KLLqUSg8EYwNjMqvHuwf83ndnQbjkFJJS7c2A80eT9DB36iFQU3nHiO
zk55cW9Cio9R95GGfHEgAZ0TMG4Ir+IriJOYFXYVLNJoU0MVjyal1zQN7372hJTr
0AxQD2sAdAwJQpDBS3zu/4u2QzYzLnV6DPv1UJ/JarNor/KwFnNOvUJWjArFOWW/
9mkUFdD8Yriv/4xVIEGcJ3ohZVqGpOFQznIPiN9yXL2mmSh7u5oULIAb7VSolVe8
oGeQtlwOneo0CVdxxk6x/0CkEti/daWLQVQgYwaW6kEu63752DRpx0oYvDLCtu9h
el0z6MbmlqyMZ1tL9hFWamodTZ6Usl5ljX1VsI/uGSG4uujm2QpGWfDXI47PmD1U
UkYZ/T8LGNMCRGImsbBouR1fW0XeoObp1VgkfYmzR6cUcLs2ghvzsA+PerBee7TK
23lPzmpps3B/GnaLRArWYF0cZCImNmSFR6JFfApYKKtPCKZ3Aqre5KZkxMbVfrUU
HSeZafncuicirwvAg7aOkGg1lhUbSt/LosOaxQuLg70THD6k+HE9PpPy2DdpvGTt
hmXGkEtyM60b56n/CtEzoedwDHTEEQ8yybA8Bui9qdnGkO+k7nJgnTonDnB2Dn+M
TTSMv5NZ9mTLATr4Ylvhy2kO1YKJZr+vybQfhuEjmOQPmDPndMM2Erk+H9N0MDlL
N2phaxCLtcPRe1P9HMy1OwhNGKiKKHzfIX4ClMeKiuEaozEsePq0SfCzy9BY9I0G
Myt1KIrcR42SM6/rtnMVeKbzW8zqLNffnmB5uYDP3qPcKcw1+hOn0MfUuLUI4+UH
k5OVyI5pbWik0a7zd7h5Om+Ls5XyaGluhLWjzYByt3iymuofSGlBxYCB2r0pd0jp
KRFVEELN7L581+L5EYVPQPhv+bw7bWtwwgIn8pFTFBKvkEmvvkpwrm0lmBpQKorj
OP1mE3dMoFb468GstgZa9EjA2qsLNqj2Y2xEKG3Ansc8fwgWe875ub5KNzGKpFOb
iEdUEAcNsi6VBtedgvJcB4VxSJU9aR969Qpi86buPFoITzgVz0EvJApBBzsoDg2s
dEK/rH86rVtoMiWOwG8EbtunxGf1j749otbSMpBUMG9UXCI2USSSIPFQxtSL1Nno
DS2/wc+UfAsA+b1vvcwdP8lS6rntmfPE9hCPHsh5ghpUT5OE+CZbUe73nvoU6e6j
fAUkOdxj0G52EmOpoioiQvKWhSzGn+L8fOmkYpa34bBnVmB/NbPAxKBZoxS1tsWw
OIQAJmYWKnB0PWDtOAnn53AO9X2AmCsmsUZq2qWR43mXk5djVSJ8+O0nD3UsYREV
HIagogJJo22q7QUN1WWa48SDWBfKacTiT+o5zOKNAfTYYQmYK9GtYlQOG0Fs67Jv
+1vKDpPgdfs8B4/1EtoKmgF3NCNjIk1XaGv1MwoFDLjtSVyih4p7kMQX0WYvD1L1
gYhzyB1nDNf5qjMsp0AIblGgFh+tB8tZclIrfWCshRB4hAlPJjy7PZehzmvyqay7
6kJTdulww0bqlLeNxEYGLtR/mpHlSMrFex5Q8h021ZAyf35wgOi+UROx6YEfZUC0
5REy3RZlYAOkGidx0F4Phq/9w9powEZRjfCMzorjmgwcpO2zgr24Am41Ur4i9pJl
1Mm5L/csoVAnrHXo17hoDtcrntQYKfb+rGJDC7KQNWdbo92cQxX6qnUp0SMnf2aW
dj8Z684guTMoSLVAeg/1i2RAnCG/Eh9UQYn1xVj4OzIEvZr3BukIcC+ByX0TizsO
zGYdersSqFu++ttN0HxRnRfW11vhvUBqJORdbsvyl1daje8RFD4s7Jp5fpFB4aP3
wef8N/6CQv0hUuzSpRnv9wgyRe7xn/yAg/ZYUBOMkOLJzYse5FO/cQV0+N39NElS
XUqPKczU2B8f2R5GtnSaspj9Zu6CV5coRqCIc941rL5EhfhnvjO5opSmsX87Mcb1
lrKdQHkK4AOHQYYlMIRebMKp1sP+AOi2REk+hvOUWWUKnItzQuhgGLLSBDw8UkcE
dPqwgTV7lxmFNWpvPXXSgzqm/IL1re0aKNzB7LtuEhOp4bEiwDip9dpXBiEAriEe
8SWtNpXzxl2RdV2gF6E2CpVvz/bmZbBvS7SYvPGzNp1Fq89WLd/Z/IBEp0hjz+H8
b+btbv1RJ6G3/lTFcfH1KH6qByhNxMsvaLWmqjDCt1FgbnM70/Iu02WsbGga1emM
06BNbXIZiZAspv8OQ8xJS/3PwYQvX+HscJ7gQWCo/qvXUFvnjAayk82NVDw2VWbS
pFGCXWLMWK4cSyyWal7/6SP0JZFsFHw8P22irubYufCxT4WSjcHN3AMCg3lBu/1n
wjKyWUz97I7MTY9obrwvn0GT1ahQS/M22DCOhPO8usT7IHyMxOy16t7NeK12q8+r
sKgoF0W3U2AT7rZbotQuPkDmImTEr9lF7yGDxgL/xbI4CWWJkaMw0dClNZUq9o4Y
nEBEQMcVm6Z2e5F4cwlc9ED5EFXiunSKTYPGn5VeEwVtFKK58W2bZ8GcHNANbJF+
J6h1PikyhBoCV+mPnR+mgxQwB6daoWB2MZ/215JsLfLVZ/dBDfOguxHyHzFbu0Eb
oK8CBJqcMilSEi38VRc620YBx7GR9eDxNh984F0MoJCRz4UxxV5FYC5fiNGzRRJe
PiezcwZIfepFzZbWDeHuuq6HfbJ6ak394sFxlomSOx8uHIYkdmUuLN36Bj6F8c+3
btC1GzNrSHgfGEj/oJTGJQ==
`pragma protect end_protected
