`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CLK0EU++WqV+9wgBVJAbF9zPEfUDxwxsxkUUPsGGAnLeyXL85vJu0RXxtkFzx8nx
VwMwVspDrWqe04VwJmgxmrUriUEVvOxj0pmLWgCxQP3Mcxfvm0+13fSdaiQGZWjB
0gPMt6MLU8ctxgbzbSGor0XCplj9UKrQrzaWUhvc+rY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 749616)
pI4BNbxFnVknNKNnS+gLUVJNmm0nJxtrwftR5qqpfF8/osWJqS/ZGHTB1XjNh0eg
LUR4Qa8+Ed0dnyzg9O14YkMnSZJmodwQDiVUXNgCjagRHbTz/Xw98iWM/bSkF3fO
ReZhN7XozbyyxLzCj5cHmw3i5a6wbVI4qJe7gk7ZsANaMN8OC9Qzk92BPZV28FN5
sm+qfSvXqY9zBB9RzpIcBM6vVtDMdZBumPzxGcSR4JEsUW1gXQTL1jvULnyeYGQy
/sbd2Y2VnZ4uQuFEv7AA950WYzOgphEXintynXXckT7w1ZUWkdwI0XHZTF97pVeK
qpYOYTaCMeFcDHAkxICBihdCr6Kf4h9X/f/V+He64jTaU4B5D37nsCRwIj3Gbjte
Wkc6e+rR53RCzP3Dm3W6ipm1svNwvgHSCpL1soiKsehzUSpsdYo0KGIQPR3Jmzfv
6JFNp/loAEJiq+XEZMC3fR3Zr/nY6LYWPXLtorbAlt9EqvRePgDD//Xx8ha0elpe
qmzQiT9DMwuD3RigRZWdV+5oUVGjcrxrEoX8e8QvEVGTnbk1QdnW03Yg3CT5R4vu
xjETwNoCOq7jKD8/MXXlcOq6syQVdsKZYLgYLAT8bXmrU0/RVjnnuLWGTcUxWRub
lZMk/TOxVA+1EuogpnwSI0VKs/5NKf1o6UDkQH3xMsDabYqDl8QUOJb3H03OdwOg
M1ffVbzT9ltu0vJ42aD0ic/sq841240XYPhUDUrs3S7bDRVPN7O3h6UP0XTJO2Y8
4M4vVrBXUDeJY6sBCbiTwy+oHFIyTbY9pw1oXu98Wa0wGeXqHzGt5vp0oDxVldvd
CDWhIwkgzLXwHwEYiRxUcXIriZGS1ahaMdU0a8wiuqDO3jnW5sy3D4EFZ1dg9zqu
PWaCrgFlawwQ1vZCcMEeU5TcJb0xKzwh1FsQMb+fED5BbJEarNfE7dOSHaVr9So4
C6zlujF8GdnGHaRAzlEzqkfJ8znNWvF2wg+2vA0fflgE/4eXRffYnXr59l6Y148B
aSQ0bkkf8GFHh0pPB5C+nfUgkChFe+ldbtWOyx3zl7DunOnj4BKdjKrRulz4HBk4
rupJhJXeKBWaMhXDKbirnBNtJNnWJsiyusQOdJw5Wd2u8MFxIW7swA0ND/zQC0Am
VuMqWDb/zSe0fDCbYK80fbmcr9HPfTBHxv1lVRXoFvCVfUNb+RB1Kp863wiGxwC0
lZNbmvOiWbr7t2pXF8jBhxr6QAYufcNU6/fc3XDaijqbuy8JEl0rkMiUfTl2jdE9
6NWDlQbreKJcCsnMfbYjIGH0ACNfJVm37dyFGXRRn/MUTjVdFiC7CsbQY9HrxRrs
7KaItwILUhYzGfL4QmVjzj8Q3n31pOKYz3L2SlZJl/QaVQc8YlJV9+ukgtnfCJRt
jOkTgHeBScyXuFGh5Y98X1SSts3dFC/jIOzP61L9Qv76qnG/VHW1OBQgKIGmadlN
DElhFq4pGJvlDYEy7cdpmkFFhftH//01fJFS82+W0FoWZHkMAjJBn6DBQAl8GcIz
rGcehNDNvk91QqH9EnqZVTsm9tJxIwMVtKrzsCW+6p+52wGw9qxNVT/60D5ybNH0
OO9+b4eB1VAHUKwQVHcYwOVXK4IjhsblCIF6gBfCIZF9sVuSlKz2dZeHy+5H7w1x
sjc2W3/AGdqs0O80baQX+dBtS4Be3yrHONanyYlvXIMc2R6UBi9hkmxNWkA0zu/2
SV3dh4u8gm/vwPJbAx7LH7QvqnfKAPvtQG5neTAhyAszA9lV1I8l7jxUIYGH6/ab
GpuacSc9Ztix8CQTQrq9K/8ytJNOjABeu08cQNwyYT7+n2uNgYY81jDhv4unAuB3
5xklk1wrPSbD0JqVEdzhH0WlnJRSEs7yJpaSOmnMebQa729BasA2Tz0f6P9roPTR
yXrphFuYM/ih1+4U5kloxm/F1ZiXDYsE2OrGIKLNemjXmIsru93dy0f9W0ItuzW4
7LG3GjAAGyqVwzIYY7ArD6lfQDaEbx+3qFV8/kci6x2a1+t6b7Y84T/VyIGuPTOB
nKoQ44LDQGw/UwZNcZxI4kz0UUA+8ANmmZ6M4g6N0cyyIewfM4qAYfw6NCKu50Z7
g0EeaeuehjFZyLoBZ1twWn2LDC/wtDiN0XV+TRA1NHy+BlRYngpXlKnzHWWnayy5
WZbcu4C9ft/9IVltJWjN8SByZdaaAJz3/M9kzQ4xhVW32kZYdZi3eB8AAatjQI6s
eeWiSBDfzoTvWkST2lTkEvFawih2bDq9QZhbYSAzYopC+nxvWAenTex+o507235F
Do1LKzmwZffgH9fI5q2uXsoTODIDkB9dQhRDi4/cINMsSRc1v3Y9iVyBxpL9oUIx
NeB8w4ZLZHG0y1GPHzWmf6i+VZmBlWCXSrA+bu/jaBZuRH2rF2DxwHBBRSoVvVP0
B58MHG4Z1ZheQrujTbg/5ow/ajri5kkqKHNO+1rEYFs5WReKouG2qZIdMyGa56y+
7+YeTCa0M+8bFgAwbq2Vuq6IvFtcFQm3uFKVGr7u23G1a1CvAfAoOsAg8xm/5NED
flu3BMR5/73PPEz2V7Sksne0i6P7WSEt0duVX3pC9VB4+vT865pgS3W9TZUYJoB8
Q+VckxIB0vMLeoPK9dG8YasBMGmTFURsgEMNSTONj2HnPs3L7C5LdS0Mz4YRUH61
j6MfUJoImFZl30F2ImVm+k9+nUGnZEjsEg6iqgXfnYzVG0bIHMPsIBOoJZDBm5H/
v7zfs/12GKLJm+pS0/d59/EkDXAabQrSViQNtb1OvnvhwGAZdtfNH1uC00VVuRSU
dCk1SeIB7P7ndkKMphCh5YaHLbQrnS3LUihLzAwXGQ5blRfOsuEbyT26e3mlIkGu
Lar0p0q2pq06kZLWY9+zjHWGyzQs6djiioB0O28TAl8nsQLkRMH0yl8Cw9/pTZ1Q
i/e1huK/VjmrIGvOG4HCc+pfwYVXje+ur6c/VRjqPDKcThjRIzQ2Gos8F9oOwjva
1cXMc6CpSN38lh5JI2NV03ARSdpVHJv3ha2K09pG9wgurVNAWV+85flyWCNe4q9q
sl5Db9Q+0oe/IVPU6QjMhmsHP7Or+tdPWGKqHgNhFqYb5VEK4eEHOGK0XmDlN4kW
9IZzSo/jEr/1qmhrKYcHk5K/5cXKBlZWJ8BCwWvSSjaqy+zCEKTns8hUNH1vmfRg
CrKZgQRNLTTC2o63RsIq3qz6lzMAhQEPN/0glVCFmxwWdO36swMkkP3nmRHk3EH1
Bt8ZyBnTAlesJyRl2/Ta0X7pVbaiFXqS+3BbOBkPq8fMaAWghhlfM2emZBUZSBlJ
GKHxee4xay4W3dg/AgTm0kGhDsPoyiCAXCF19cSAY8xC2cnHhOiVI8G7naQ3nO7V
ac+yG0ANEKlB8wdWmYB6H8rCq6reSwMY3Z7flsfF9bxujXoxOZ/fT5wlG+yLF+7u
zVRUg9+Ecyj8l5s53SLRmRGPf8JBVBb6oQBPkrDvU0a56pNvalxrASIL99H5ZczT
nGWYKAVzAwja/mzRwVOavD3wzx+DEquoavAMTatXiA0KWfddFgbyRUGjzlirdJN6
uLm82NbD9tGAcee+3EHuFJnFxpQ3yKh5iVzk3c3ba3aDLIt3Oo3xZixejeFaWqik
UIkufZDaAj05QVQqxEuJSJpwXj2hiBXT5r3JHYuv3K5elrVObLg4TPj29YNIB+KU
SE/LM083tDZstuC3KzW5aqc0kQwdwKDgReODwIDXUmDm/jFftVzbnGK4GDoggrYn
f6LM0drOjEDacso77PRwNU0GWkGYkcgknVxRA4c1ieCfHlwwz/5bew552D4HeAdt
AgfmBhAk8Dkf9uKSa1bEWHiPt5h5+oD/Qa41aD621ZY51DEHbE9OMLS7465CMmXS
uK0WFQCNmniwScIFLt0fbMKRpbluWz4xGbZnMDDv8e7+js3D43BvWB2lCzxE4YDV
Bjj7xWyU0fhW6m1n+6eyyqvEIv1PrnhYdZI9k+5zdELkv1AuLVx/6BcDlEAHMaVQ
kuDoxoXiTiW7zdwij2HGaTf7t0w07MuKfep01gQ/6a1fvt6JyORm+p6xSiSwOqPL
tDok9Ee//xKpF6niesaE4NgowtJffkTfdyEg3b2SGeI0hX47IKTC5xgNUrCqniSg
nW6ek92iEl1OorSV4BvtGTXE0GW3udZ+WYOoIaQwb6/dMm1nWKowHAZWSgylzkDB
+xFxLcFeld4x2zpvlOCWioAMysU22fMhlkOTapzXvmwdK6J+d6RXJ9j2SXg9X4ao
vLL9aAH7DbFhaHg5p2H9yUfdkfwq6qZo/Uksw+2Qirf14iW0L65dtjsrWKiZ4sxW
RoANxvMgsuE0mteW3APWfxcW7OZ58gopRmFRieZSdc6YnXNjDg3eUYcj3J2hoR6H
QPlENQdq+lejQO3FzC/6k9Fz45AvNTGydKWOivxG2MfxLcvmylQ6JAYE1FBW3FaF
Bv/OCTNpYoqVgti4uGuDPu3ZOPnvegTTqVZWrRn8cAo4vhgtoAJCwuTAg9GwnQvq
92VRgycV5NE2T1pF6VOqcjSeiaiwa0ukKee26UrI98+4oZ60DIHc97W+yGETFJhg
d87OqrNPczaggOpMG0YRPxFcSVsYfeYuqUmNtDGAmTsoP1sWkzNoUg6vO12+O3lQ
vVtIYEKPUcf6Lv7VwR6XmBxsI79JE2c/yQNvG6GX8++PpxjcWUHah7YZ2x449pj1
e0/Qa5jLICNHN0o7njv8VbNHr5X1wc08FKEfb7hRUi6Aq/l09ART/tNhvC6w/k4I
GxV30OyYqZw2yFTOCoO8CWhF5zy+hIU5eNzTLxnEqRl0Znr3bgzMpYlKbKV4CknH
ipjp4aNo3/qojDUcn9knMIRf1ol6drfg6i/1tbAmY9Lz+O8bPqy5kYpEMrvNPiLr
RSuz1EGJj5+QJ4MwU/sGZR5IBaqx2hFQ4Lo1QXXjwjXrHIe1VLkThmqeFo/oad8C
s+5sPfrERSiHt5zOHacbRvZeRdoey+nw5tGEekS1d/g42xNtIMcR+rhA7192m+d7
4tQoDglgLn1Bv+5luc/2So1ekEU3VJR9RBOUqpvV/mIZYB6EQw4PUo6jUz31sdK4
QQ+uxXYdQ3kTnL+HtEUU1PNovjL++snrfg0w/9CZo9U9JVcV7pAmKrOBiLASWaeg
6ym7JuWJM50n0X62BLv6We0RZaVqIGwG9sqvUGKcTzpv1Me2XhL5ZSqpET4snAkw
4jAd8+7wqFttlfx4vzSsQh/gTOmy+gPLe5JlseP9xAYsohbnlD3CCrJZ64d45noT
xN3xmZdi1j2uJM+sXtF5I09PZ2MKQdwNWQ9oHsYHOlYtRqW3Xck9UelQhfocl73d
6UL5jJf+q/hVZhJFuhl0Wm0nGsFTETmXp3pKUjSdzI0sk4T0BSdNSWhrzMnXBOIx
PTGCLioJXwnU9cVTVPwqBUjEae2kXUFDT91EyJEFYsjq6c9uiup4a435yx4pboJd
6ZaW4Y3vxH5y09b6PuMmia25VQeXs3Vp0Sm4WUEvh6gIdpPYMcUOyjKW2yG2abs8
OOGm44wdGqlYREpc/hJHZ95PCqV2YdnTfy/sBrqIc8ivAnltswo6WaG7YCSVtvin
K1GuPHPpb6xdDlkCy1VFDMAHzFy4lp/zK9y1b46kJAaaEZCwhUHZ/C12IGljusoB
6+ILMnuir4tE8H4v5LZsQDw533KKcJLe+hQ4OGlC0ykXmPq2ds7gI8NexAPTREX/
zOQJsuhFiJnnNs/gsE253TKdye1RWxRLtBPZfrIA6HbGihYcleSAK4Gy3fV/UojA
IQhNZAtFc6xShHA+X4GuAaigCRsksB8FxSf1NE5wIR+gstI4axfew09etAmHNTvj
5nh8my9BxuXmHNYRK0co7Ec1tGeJaGwGJmms2PStOsFIlFNGd3B4aVnJcwL98Knq
TddlI9u6bhVeGyFK0yrvLZDOdfsj8J4X6uvZaaXP56fYrnz1opM3kNj38E9DZvbE
h7KoWmesKU5iz+DN6HBNNg2jUVQz+p056FR4d2XKLO1yJp09WJHGxJ7d4ptDZ68X
xBVgIG9rBYMV+gUJj5V7QOdwVGV4IAumDPa3Hb/B++DpqXu5IW0etRqAYyeMBw5z
q4cngstxM+JoDwkg+ZekDlFvASBmt/RUsU+n0ML1SLZEECxnkDVDDSYJ6JM1O24S
zAqqsdnYoXX1DZgkYlAcgU/BayyCjrsBDxsJ9kydEZ8LJ+TX3MLmCgqGWSQy4gyS
DJWvIVo/BPeRtjBu/ImFBQuVvAjY4ktsZHJ3IDUrGbC48mAyExf2FI9fWLmpS7x/
60sjKmWr/1JYAZxHC0JUtLjKRoCf0qtugmt1O2DngE8uT2R1VAuzq20nOgHkxmcH
AfAOZvgAKY9quIS89jAgGm1ctO1Hed0uHgqpddc2ecX+CdP+aXIAz9lkxN+0IFkv
dn4DBp1cPVVH6D1vO71cb4tV+qKCHrdSGF+hP2a0zVsNcmHfN1lAEwdepprELFMV
FMqXLC7WrMrfUielFsvlf/5rUzMdYq66/tp6Ah2GYWoZiQM1SkwbY1+kkNU1A7IB
cuLblPQHeJ7sJsDWms2U/vSyqJdTwh8iJbLoc2NUGXvctpXYX8fFWZFzmKbbf16G
0qlwIepNDlFEiJqYCQ8E4Vo79sxHPvZ1yYqwJ3ptN3nmsw3y8yJ6/YJVMxq6MDQ2
rHDbxECBbmdmemHybwlnKflKehvoSRDw2OCuZPcfsCUw3AjTiIap+XJRyN5ziQz2
6PhyL+KXZcZ+03omGjus0yqoHreOz48epuq7oo8RE0E/QAuxchzrCQEqj/YORrRb
IsH4E4facoE8fjRxnAhpnT+ENZlnp5vwJdQl06OjbmRfLQ3NDs6LSTQH4vCLLMEa
rD4gvkn+ouOurTykc/4JVhrLMZj1CE41gWrb83QnpOPUHsT2auRtUjIEKgk/Z94V
5BRQPVb11eCdwIHLl4tOupUnKvX7S7rumAjxmCiYeRtyMzk1hE8BhfpFZgKJHzdV
kwhao5/97FeRuJKOj+ugdx8DtyQei0rZhgeYhYi4cCMQl3SGFaMF+5eE7/78JUvl
74qj6FaobvIT9KYv68sQ2rIHDBJRA3oGYkwzM5cJtg8L69odhNhEbw1E9diEgVre
nbhkaTtBXRhUvsa1KZyTAObkd++GxPTOQqjTCKNiwR+x+btTr5OHInaZxWjN4+rY
DMMb8gmxMbp5UCn8wKOtOUD1Yoqe1lrdDvxli0JF3xLgCRI4W0hrUje46NJWBj8c
xVYJpGT3ZXEZYbVlWVqu2XD2DFmChHqgkyCUM2KOH6tAiDLLhIoFoMHeCsIJsqR2
iCCpdMWhrjG1PZhG9SAtvbVBtHG/IWHOM+E1km+9JctD4XG6Pvt6HAnlvkUz8Syr
jrinLKnw6Ez+8V7dpC+BA0z87hV5CKzRQ4JMvNamvIp2IGS/vkCQDeyejVQhvlrk
HaPSsCdUGXhelEjneIiNsf/rlU8jauB88Qp5cf4FLJLCPBwqqLqVOdmrFH0UvY7v
mKcwU8Rc0pH2EAe2UWjdGW0W+hx+DdASfpF38mEtAtaIT40RqcQCkZmXenFlbZaQ
K5fYZ3R4aRt1cunBNm5pDm+pqP4cX4FDQ3jLB5F3e/fMlyW8J+uBwBJDcWtu/+fU
vNc+RSv6X9PnNUPRpRxhFwYKFbGjMEZ6b0nb2zDQEaMSFMJ9usPdCmRtfobi4ACc
zhttTEDCXiVoRzKCjrRiis6U1V8uji3gNS0Ha47JNXh8nifptUALUwBgsG2i98xn
u+J7dWV9MOP5dM8/3eOq3amF9Emr7UMavI2+pTlcC2qs0BjlnOgjcR1NoE91ch89
tFLEBkHJQTsCUc+wsmgFJA9k3o2DOXrX17tQJqEwFs8UpxCwEH+RoqSZAp/ptkg7
sILGQTU4CckEZJVFqjEK4R+M98uhAR0c+tYJU26liq9mrFvkBUCu7ThCha9mhJ9c
h12CKDVJPe/OO8Dy13ER9Au+M3F6k1ZfzBmp3RmysyZ0umtIB3FIGu2JUH2zYzZd
v+HsAVLtdI/S/DFc4JYgyMtN19GyO1A8DihCmQJ1wdlgfXdluKMRd5IS0fLqxxqm
ks1ahWWWkfWXKJeaZVbD9tNfEoDAIORgyXEgJVHxZRNUHPkxih7fth3l0I1dw5ZD
+0zxFUNTXH9bbIFJDE6kxjcVoED3/baDEFEClwEEdbqb1xjfEmqU45mKTE8NA9PO
UZdKifxfIJT6Uz83YVM4cgE1qBfyHRIiIa7W890MflNuzO8B1Zx1AIR501hs3bbv
Zn6CH6cPUdK7d0sa4u7A+jQn7+zrseOReSf8Xx6Ros+RuMEdpB+g5SzUwVR5YA0G
o/EGmOrYL0/D5K51uWCxMggm0zNqAnCCstDYC9O4Cc5fT5bbnGuwSsa6PeuYueFy
9pwY5poRoJwUPUGCzq7frKfgoCqR3t7A+uw5YUAao0dPcLMOho34EhlX/cU7mkzx
qmfKTMLz+kCvZXxbU4d4n/Od11+iQC5rnJfoCUpVe16BxkOxFOTu0xnwvoxQAZ0T
zc5cc5saqCWAz6k6RCboIn/PMDniPFQiFkYnkcHd/KOtX42oDP/bSRY6W9VgFcXb
n8Lep2XvJ+EYxyT/enJTzV4u/1qkEAwqCtL7psQ8Uk8kw3SKiqI4cSw1x8xH1X2l
U/9ChzQbY6ShFxhqZDKegfEbyOwUYGTZX42nR8XlwHM/GokZl9XbZtaDQtx8UkJJ
YeTAA0duZuVa0vn+jSP315iBuS69U3dJg3qjILDLcnRO81B+mBNIDHrHZN3Vk2uz
92YXaaDHdXqiHTfVRIdh/yuFNiiX4z+1FguswssBHdN3INiNTBBmC6VUV/BxBcNb
hQ1yVLmchWuUK7B0/i6vmfTnAKq4IdFcwlgIEyv9rFkgxWse1xAX4FtIDr5YDvx+
cP0wz/q154BLf66Mqj4tIWRxo/km9AfjQ7O7B8eYGKomdee1y+X4AhelFr+Kg+Hz
4CvbjajtT6KsE1d84veBIC8C/mnJCmHuOLHtmm0W6Dc2zeb9yBJJE3yE6LOXDKdS
hiy7oj4tiYPJ2x/xUO5HsfGWJj9Ppb31/wgI28bR7qkgdqHYgZUAiAhOjvZD8YvY
L5jo/SIxclIxnnwNnu5E03nI/HCPrxbIr1j0j4ZvT6VAQFMh4gDDUa5BXkUJ/PPg
PkRIbs7rfpZ4MBaGcyg2g0hO+LQnfE9gyiMlW7VTNpEdFutdbawMJT0vhPnDAq9B
+2q9KAbMNgrKj6/lGSnKA8+SHpdQoTtsoNuIEU6CyZquEjctrajBLQAyvjkvlhR1
0qH0twZDOvYW/gHawowIBZrRlSO9WkhJ7XsIZmAMcPC7nEyHk5MVcm9QIheLYKvV
nt189AtInm4PmRVjQ3KC1b7MC7iunfQpY2VvAm0mrKHGPUAa1avapHMTP0bmstiy
d1prXH9RQhUtYuP84HIlXAcZvG4ELH1qp9N4IUw0DakNh/L4vzkpA/QnwHuquOqI
wFqJYfndS/piAoQlLPVQ9h526/ioVBfXeZdJv6nfLjRJu9op9xfU6oW/C3QK3Yra
HB2cMZzG6dcMTxDkJOV8YBEIJc4XbIKTlgDz1srtjcqPSzD/HWvbkqiw85LobbVw
l/P3t0IWwToHSoNfF7hvOxxZLsu/q+aQdWHov/+SPH0qWb3r1Yr73bSRnyNskCit
xDXNh5cvmaHQmy4SF+Ianxf0iRTaLO8JhvjTGfUXvxi/FlCa9O+tvvHocvuuBlMw
ff7P0atqV2WZY645kq+cPl3IGHDRdnt6QAtmsekwWP0k1E5nQppFRWqJGD5rsiJz
vCYVzNXO2Zn+rvKTGgSsZx2mFOnW4AlZfz9I5bBBNjYPStETHjPpxgiEJcq77SfT
y45eWS67L+4aN3Obn3qa1Xp7+wqG0ugNoidD/Gu6QrYtjMX1kpTI3GVaoJStiz2Z
MxK0aD8+1NsHIRN66nn5TomtjBWCZSrtNl/sXBNgDNBa7kxJ/vZBb8ud1+jJuQSV
VBjuKjo0Sv2Fl5uZ133RgxCvqIEkRiaaYAzD93A/7/LjxKFyTglQQxcTQQuITN70
f9NA4qNu0OQ2BCsCU3vxKr25KRL8wG3VbsgQpqT1V+NHrWnLnDKXiYsPlj1V+Psy
xoYIVgByVg38l/OE4/73g1ap1VcjvySY3LoGtwKRpSqMSYUk/ny9GfPTusGiQOiN
Og2hzOVhM/qgPrq92N9ZFOBo7ROXNBZrUBIMjf9XdOhVtso9rk5tldOG3p7pJ9qi
epMGiSuuKI5YRn9yUYbrxftEMBv+XGejFGH6ANYSLaSwSxjfCJMckRKqJ8+vP4ML
nGH748ODcMsEDw//cDjzdjiG+JaYrz+O+3WyAjuZMhqCJuMCMoOYgdmyC9LpSTSC
jDhZVJXXHtPadNvayid6m8Ivbnyng6V7hL9A0r2KHGZT/nZQ1G+Ain1OirbROWvm
lQdMOglOIIwU6uo/2t9BFzh/z9UitBkeFYOXJFsNqhJDnsU+WzKvWQdLke9KGgvf
YZrq9CVQJbioPnChfMFnEpzuwkfMdfwfabOZaNycG1/sXDqeHDhhpiW9rSb8HUUP
DRL3Olqk96R/8jPViANSu8uQKzwosinFI2F8eqTKxZTlkoER+9/WQgYWRMy77Cf3
3Bk2zw7BL16n0MSItwsg6fXYBbGlSLxVtKeOZWLVXk6yxG3koVW1TndworfL4M58
2rfESKMDnes9cEoSYjYlVvY9Uzvz0XyZ9DL6RgrbTs6ZEfxQECXk+aIabBaTP+dO
gim+ek6Kx8JtUaBh919F0m/u9+Ob9HU9q2rPwpNM87/gQYtefzCJuHLXUqZbNB5h
QnlAMAQUkzXVhP5gdfMHnSP4wggRyQyoIhyLpdbCaSgmKbBDkDMl0CacmToBjhHN
w3zhxRLInzx7VgsGfXsj3yL201waB3HyvecXTYefzaLT1jes8SDt9EFzSAHBt4Ka
CMtVK4FKrDao6L9e2jVm2qS60ltY1Rv5MjGz/BUXCpO5Gtz1LaUPTDSiLKys61Wk
gj/H4s5eRUNvtoQ3yiCcuaK9R9CoKlG++KBEHZSRaXZb+zj5AwJ7dhvZanRfVTv5
oSJvUP4CHzxESnUHbkt+7DPaxW/okFRBmUfB65ZEtXjBj9MrqRMprM/VRLHmvrU8
vhUx9gmx5FPzCwPe6RkeyWVubf6JmnZXH8VUjqx4J4iN23eVZIQYemfm8ZgFkPJR
lPgxWiGR0Gv9a4A7oYSnAnhWFWBxaO82Xr6Wpxsf8KLDUbCuARpJgpBOY/qMSEkN
7IUhMPnxCTKymoEcU2UepxnZrjeYKZrtsFTGaQDJrdvOgJOqhuuMpHljqPMG+j2h
A/kDNOjOdXzG4gA5SMvCDh+0XXOE3Ev31Uj21B6sxMlGkI2pw+G+ihpG7lPKtCx4
kF2+KTr64TH1d6P39xSpUayWF4wFGdJ8WhtO+GjPuv0eYfi6KnocQp92vcbwRl5z
ziN2uOVwg+2zqQONy4jmqLPEPS5nJDclYTXvhkBoiiBdtMZCzRu39B398GIirq7W
IRhQAr2XMTRn8OcbJjJaT5CzXXXHqostGCgT5Qp7wEfS/00ztev/o2/X+1O2Kjl4
8Bso4QhbSX62zrz85C5Lsmi2pbvgpH8xMuqm0h6AT2FuNYQRuUogdQQUY5o0k9wD
NPlStPcsNQum4aP4JPiJAleknGdVIUAeeb2fNKG3RU8Ow3KU7YL4ri+FV83mgEuo
vMjVgKJlAjdhApShnWGZEOMR8GhJDudDC8qE1jH2vOiqhAJTZn95TqWBdAQ07eT8
UCIEw6hMWtgyfUxEJKxa+1O/N9RXVIwP2bUmVQ8wRFHWTK7KV92RCD82WckH2XLq
J6MCSSYMcAIxMLHuYavPbbfXanh3Ys3u4zqZ4zbkyE8IVDwIS6mE05Y/6ZRanpt5
HO7WIeQvixidVYyTOUuyDFdA8t5aWfd6m6PYg0pwQ6c5lqVE7dUrrIqV9f9HowbP
wwNURh3Z76whah5ikicNASDe/ai4nhXzdChoPZkQ2ZnQWNVsBJDqPS2dFJd4Haes
aTv1O+7nDAjPdHpH3U9kY49IDFfDarpSZKatYFwodErt4VnAsVfXUMwH5wK1CyyR
pNxjtMe4F94bnXnGkc1QHJBfIo1ub6uvAsp4eV4sJa6RAjkbBCMY0PHJTBUaLTDS
6MmDzzi9z0ZwJRoLjgkicm90qt0JGMy8bUsvAFQoPMnPVGhQGS6x3XKJIwb3AfOZ
PF34TCGpU2/eCBatLXgoVS9xUrWqguf3CO/caX2AAXao2sxv3jeAHsnGnW9rSx6p
4rQ+oWvmQc5T9tQWtTK/9BOLZ2wQwoAj7K9+U6apWLzCisZJz+3f0ClMzC52gf9K
KbSyBr/bVN+8WNawsCEBboSLLt0vAAFnIIn2vL+pTmB69KCfk3lFAoVLWAw0smdX
YH3fqaJLOaoz3OfSmabMAfOTYcnEMIanR54R50OF1QDVc62/CXt0CZ1Z0YOocSdZ
GQvfu/HrueYpX75PQJnRZptl4iRHf4a99Y21E5uI98vPr5iWUnAMVXpIU0eXu5ue
4+A7preU27fnDVDiNFdf21x8e43G9gmY+AEp5zsEHMLkhrtnAzasfTK/Rd+3qZo5
yfIY/VYcBouqQpptSGCyMSJ97+nwOOsXvKFBZ+ArHtiCUR0xZhRUEZ9YgDwFfN7T
h1R8IWGCY7FUZnPXg48tW1rUEzwMF2n+z69OzkDjtOuyQqDVVEaBoSqUMq+ReBDf
73GclgieK6SV4LuQQ5iydRMoQgESNf+axesX84w+CAOpQlChXJRQ31QW3cVxzuwm
sqguQIMc4C0Ww5tyfMZjDac20krwzkDXV8bk27qZ07pH3oVQxMQJtXrDmNA12UgO
4PJGOuCJ9xTPm2qFUf2LorwVZ00rjMSlOD8wXxcoxAkv7rrd5Lx/s7zwKti/mDWN
Qr8fJrs8dVLudRfpwRIxZJ3hatOHhY/27TC/WJLi1BmqaKL25utkkkf+2rp7ci/G
HIyRMwfSTrbOwdMaxk/VLAgn0E/QKvFYyuddruO3I8jShqGi5vV+ShTGVOh5agwi
CQpSEInT6lQcWNPv/6WVfN+jzLpg2ImM/lhDtPxvXOFTAhXcKg8B3e55aAqFgHzk
PJjfZ+HkopApPq5nrtLy7zs+mO8I2ioZghwyDQ9XLeVBYjjATiC4SCGs4zw/PU0s
v8j3PWjXVLSDtjoz0E0GN3EmeSd8YLEl/1ed3vFg3l5pZUmGnJty0XgZ0BBsBhMF
UI7ZutcLOgDvNNRrjzeYAmyvj6N+bxUtFqmEDLa7faVGqx/0NezXe5+4GTPMmPF+
opZsF3nR4jKhhZEJpm2okLDVm8RlV84BuANufmrd7WRGSqEazLS2BDGiGoWmAC+a
TiOmAyVY9WaW8OKmQSxfccP1LlAzMK0J5I/QEM40fsLsgoFPcSQo3hMmlLcS8Avp
zylgnkYzusKdM9xiaPahIgsNoySb8wS4P3Q2LxvCDsnuLYm+VKLB1ou4fdXwa5r6
dnGXGVBUWnLT2e0IPbaLR0LnRsrwYCE4oxBsL7dQ4wlJaNlv868iAtapkoYWgHKN
OUlnH4gTUdVqDcRKrE1zmigitIB1azVAN5Lx8Ea6ypxrInhmeZL2mAR7EZCUrsri
F11icqRd/pjJy1/QZFxGwHPjMW50ehHy+2p4Jufgv0uf+91Lmt9VQO2kZQYEBE8s
0kenpKFTFqjdwQ84T9avC64fTAvpi9wOxwQ4If4ZxCsPF4FAR3GLsEWH8+4rZBWv
Tbp9x68WdjMBM1aRcGV5bB7elk4fIf+MyJmetg5WlhDUCyccYrmxcJbW6D/OanHm
KpgN5j8dftPbvMt/y8BrNPJ+Rlmg3217hbJLz4Ab94MJ290kdrHrVDaK2iwdrMd9
F9GtNxNYX0KeG6138Kcuj+C7vIAcdXXTp6BOpxxaYIfZPJ5/nPl1BRztFYRX8bVw
3R3OCiie5vIU5HX+blt1PBZkQYup5AZeietq9624YFUhD7u8w/zQ+95WUle0hNjJ
Tjerkhz2OklOtq4aL2lPc/zhsgGCCxAWdpbl0zJpEptUSCSl3pZm6hcb+/Uzh9cp
1fQpBpAYP1p3sCG2njh99YinZ2GDJTxebfKsrRzFU+adn+1CjT4xSzVctzE8ap4X
pWj1E+fv08zSWi2XKXlCV5+U+ezEtApD2dZqap30GF8j/pYEnpsN2Gjstul7ve98
T7wAvPMP981oY76E0fm/awe4zI2Jbnfj3OiEzgspGafN0ag/GS8bXi767p43zvIf
JC+tjBby+gzqEvwKQrFk5s9blQ+e4pdaPRm5Lae4phqzdvPzlbUa1IANcOYcwWum
8uY19N3NmpTxuKUKk85d0KqjCyrP31+41Xei+3LfP1h5mftqXqnki+EaBMqzjUfX
cpEdlTqAdo8LSBE7Nr5PySg1+mDiRIhkZdqbZv1LfGQWdw9MEpbmXcvwQLH52qa7
wLzTT7jv4gxce2YV5oosE9sIzaKopk8eFShjR9cALvwe1kSMe4Mcb08ClkXKY4/D
8bqEXNvcTGAq5RL9MVdd5IrJnx0bz56UQIIPYP2LGSmXs/uHUmVQgQue4kye5xvV
OUSe5dvInwvhPpTg1Pjwp5uvkXoWob8/QAt4ElkwIdnpaslY49L0glUQvYQnbMAG
TajZd5droG65dF1ARty6Wn8ejGZ3GddM2GETRXX3+OI8LRCf2R12V3vH79kZ5F9U
KB4C1pwj3Pt/qWS+LtQVhF/Gcv1VxFao6xj8WAXd1FP9+Gcg4Eut6dC/NxPqLilw
cWbUNTUFF6tQVEXQBpwC/1VXJkRDgfYRKYsFBxPhmIQxXY77LPGOnIhAzYjX8fXt
Hfssr1lr8Rgeo0xdqIssoX5rFtNxM7cpu5z0WxyZ83n9ugJdZ2GDFBWlCB4yV23k
w/m36muuwPxznn/exewhavFdxQt2B18CI2DwKr/KCv2QYnlwAvnS7+39xn8pakvh
J8DgZDZoLCp4dQ1cFg/857SYDyFF5d7lUKLUjshpoUK8yczp/4QIcazgWp4QTQhW
QmInMbbifvQ8I1ytFQBRKyPFQ4IAWMrFirgP4l5cs7csCfCy9GWn/qBfCmka+ZiT
h+eFCTdnSqkUrykI+jH1i3RI28oRLNo3sqs2V0uf7D59M+Qxtj5jJqFW5v+Cnxzz
jxTSQHdWEz/S/8oDXfw5X1O473Wxo6OpVk5ZU8Qn15kfl2+zsdO6JCeezNS4VdpO
iwlWA4ofCF4LoloB0kss/ftmalc+JZSvy3ECDrUzEkoNF6+uH0MFXuBlQb1LWgQM
qNvVI9lV35Tv9H1ffhC8yMIdiKBicTxBLLxsPjKlklA01OZj41QRCVz4BaJW+HaV
GzXqQtH8V8ZsyluwH6aMzufgt6VneWinvXQjHufL3qh1+m+U8402HEEgaM6HkhAh
joo+YSlUp6Jc0UTLNvL5gsKjPlYF7Nz9HPeRun0wFKXgL2tRrrEfmfiIbN0UAKUD
o87YkcTB/VKChYEgA71dJSUE6zSPosi+uBA7bo1EHWuZdoFUdWB4o055hZJTla5j
Z78SJm4RFdfOi4yOJqNaylTmUqwJzzWheHyLs1ypxu4aEOZ2jd3Ttfq0wL1ug2t8
ZxJIXdyabs6Vuwkc6vLhxYdYbQPcTOwZnvLWTzme2wKbbfE3/GPtNxqejH4efvFa
wpBd94Drmqe3eCYdIQtJzRFtBZsOXb9OFKrsHZznfHtycT9NOg2SqcEgZPqZk0Pd
S6yj0kb0SNWqlJQv1L65ceo6arycKoef6kmFKGIOd5K5PrQM/bSZs/MlDwYJORjx
6icx4BvbVcEPmrRjwGO49aIt6ikDW0MOjOeJ9NLatjwNxgv0BOiHm6h/bMReMLUF
4/WLsM8T9pp3qArmZNtsLGHR1RVS17kByaNwAGDcGtk7YK44ca3ReSm196dA1kMJ
YyM7l3jOXQ5w6FtYwi0P83SVyxp7+WC18o+QsXpzsF7s+XQcAU+CR4G/I/Lmfvdp
KjBqLeUtSoSjSIWieSjfuZZDJOycF89xO+tVqUslT1aLTAxaP3mDN/13FRgAiU7I
89En5jId1cX1jkARV/pr/DeoLj1+J51doLkQXxXGiyEAXynQv8kK+L/8e/SWQ+J7
UwH/ocx6CAA7YU6jsZXR6vH5izjNsysDrvU+UI2UXlMZxaPMtVl7+HYS2FmNfOhi
gJV7N+EHVJ2C+2cXv6zriw4NFDUyRXVwEdihNGQaVP6pDqsEiSyEyvlfNHH2rRHA
tvw3nsurW5tBOtBlaRXdOx0ZomH7fPg+wF6aSkcTKInjrHeXnViKUTflky7gpcl2
1ViDXVpbGoHebY10p/WIma3ZtCTZQSPuJ2/4YTcKdchoBp0uIobDRhPmI4H9Vg+h
bGyTBppje7sk7uaVyzDFBanB0ha4SmeEfMuIt4+ZOjlJ4DRfz7Fn83f0ohQP8p7J
uwRgS1Y8cApjRVERHV7t0A8AvSNKHA+iydGppmk6yWnCKVkoAOlv2huF8ikKVRvc
V4XGgCysaDMtnBxFdcnUYz+Ru+QxHKxkZhoBZMrtfhM8GpCUyzMNRIKbC86KtKMF
yMTabcna2+vpQZFL1kcnui2YT27oGJ8fjz+Uqm1Qylku6gkf/+MnWiFUayJHqNu8
VebAjjbD01+P+NQyeeSxmS12Ym1unt+27QHFuPNWX38939mH2z3GuFs6pqacVjHO
AMAnZ/oojM6lNEtXpP5u0JNwYr2Qmon1weFYifJ3fGd8q8H+aAUy2Ss1MwazfoC4
vo1+fCAD7pIAkrY/Hhy3aYDj+5GxKyEjo6Rz2w7EHYhviKlVeckDXbiLurHVeDPo
01Q6kyrK7AJP3o12VFQAeplChkkYNKD+TMulhmGVPCjl49Iw0Owm7uwGQS+Lt4j8
yDs977+hTVew97e8SWxXCI6eNmEmKk4AxiAC7C/AxJUMR95e6sVZ6t5hzK4AMPD0
+bVU/8Q+qCTV00m32az51+p1PtOQ8a7MAD0nY2Bv/zMGlRQkPRJcYDyDniyKVc+9
DkcoQ7OXOD81wA3P29NYMgKhC9oNdnPjHgVcqhe7c8ZsUx4pgKJrFHjc4ZG7FAdw
l2ZQ4TSJaPjqf7xo85eBlHFIYZN052dcrg/gJwds+7yagbP59olvPoVErVU3WGhi
F5hnosy7GlkVnWDrkEPj6jSEkCsrg/IgpqOkk02uKXZBe5yHFEs4SkxDRD1RdGV5
K4Cpt/pjeUlNOpkofRBBYhbmP93u2b4ntyXDIcexeCkxJoK4ygcngVxW0m52El0h
IyXP7LPuvI5ybcOJT8gOxLdukYCln+Yu+pqbgICzSD3Ec3TWaCzOqqscPnDQaZQb
jHbfws1WKp+1TU6j7IL0rRSg9Ujg99PLChuYwJkaZ04woQrFawcCPYflOIvrJiKf
Rv7THTgE8yXv7/aKAs1g6o/E4N4VEpNrGacJTAEIjTZxN2wkz7lB9ZTwjkYnb8kf
ekm57WghiTQP0FbmlY8g/GXHz46spzebpXHhl8V6O57CEujZbNz3Q8cvbvsARbD1
BjT6m2T+LAmDhPN+sWhf7M/KQk4SKu3oiduBzeJ7WbIBI1mM5dvyJ470tXaBeyDo
arUDpq1k8F0Uf5RIteoixUUY2Tj6VUhAOF8Dq8D4gblDq2QDGoW/5TcDOT94mEeO
dT1frYHw64d0cigUfjfsyI5HxKS9hv3mJfakt0b3iBDIC9AfyOlrLijwQToIHzoH
yeTrL8i3aYdz2Px+1uq2ubZX44RVIMoFP01jLQsJckBjqqiWnAGARVK0rReHdhLp
roLxt1pP3ksm2pk+zM+zG+cnERevaMhvqtsFL5j8GxeKgrIZYeHUwXk94ZCtI9Et
BNWgfTvy1za1PZWrgqhPiJjQUEwWFswbVQNcjFyL5YXkabNfdNJ+iEf+sdJ33Mc+
4WJIYhYyl/CNFeyo9mfQyNWus619UufF0MORbhco04z0bA7LsJb+pVxmL3gUpz8I
zKALwwPZkaBZ56EBKMBvsQLUPLg8KJeYQnwHWvQNGV2P1yAij4pnHCk5QHmIWsgy
EsEjDs9/PxwQ3Jr03r6oMzCJFxpgG7oF+4noqo9tv8U6vfTal59WX4gEZhfxRQXM
GEUv6pHS50lyXQ7YwSfv+jv3F7wuxt+NaGiTTjIf7fSWVb51oPqKJEerIbWFeMhM
LT+MInPd4dR7Xia0MIVkcfYOhHAeHSZeHvrdrI8GF9Z4vMuBeWMrRDHAnQoUrKVO
b5E1KUXQZ43j3c0XBnc1CpaJZfcEnbFdXcMdw3Ej/+ACT5zaTD/QD18PNJx2mHx2
pZWGqeC+qLU1z49P9LkjYIh+GSI/mjcP7RXi2j2Pnn+XlTjtFezsjnXrvu1vmT8a
KAW13QaaFsKmM6XzKZfgCz2c1DnQAg30ZSeAjhH0AYK2snMiTBvTYzUxm6FiYj3m
pSi/2sLpwB4sbJ0WvniXo8/IaDA+L6XqfohxTV+JHgL/8nAqnm9yXuJ9/QPmrK7E
5hzLpzjrHn36zPxYnfjasmEfrrZpp4q9JV9MLbDRlvNRuyPQN2D2uOkhaNbFb2cY
YYS+7hVr+pFIDcnmew0rwrTsV44Ej9oPjwMdda8uZURPWSbYimT71BfWJa0l8a0W
5PdY580acMxn3czbWXU+3AW8oNCo5S8GiufvtgAOQ5+hvZS+dx4FPNjGeC+eLwqq
WvuEVamzkLi03eUH/O0MxzR1MMK8gAauXjbHogfrwOjbduCfNcKBo23STtVgniBo
X6wrbcmcb6OKsxiYkqCj1tJSZ2FI0snD2AuOzg43H6PXB9WZKKN6brwSeuMIMAvT
Am3cT95sy67IPoA+gzBcyJalNj9uHtJ4shA34qzJUPG8uRTI6YZPr6PpJU5Amjiq
xmjg7qNe7RgzMC41tENZh7MD3+7oqFut1qnzb3M/eXquhoxK9cV7vZeHvEqIdT/D
xMb4CJcNIwXuLw58UAWox0Cph0DSa7BMKSdMKyPMxlV4oUQvrlMovlS3kmGpwAcD
LvyLPX6OcSmpPMjGjqG+ceYjEstd6BspNGZv6ntOlenbn0aQuH5Hz2TvY3ugvzxd
HTt+YudUOzKbnNX3Zqw1Ljq8Py4hlE5myKoa79WmUN5kKfdSFRVfid764ZYI6u/H
tUrxmaqWQn2cT7aeAuie5skqXLm8C7xLyy5MSaEieBB38HG3ulmtQNqWav6fBt3A
Q6AiKR0k0vPAe4G6nw/5T5kzeCFnBCOkSaPgAWg1QDdSaqHOjUQd+4yv5dDLg5+R
hhPeAf+pxIMw7PuWf9oXa13Znuo4pqBvrh+NoSlTyUsObR3dGsFtoAKU09EXD50A
DNa+COdXSR4TsCSD+PDIYwC4cX1X1l73Zhc/rD737WOWq1uW6EZqk5jMmtWE09pE
oDdikWxtyr6a+/qKatpNsqiY12oJHbkC+N6hD+6vImx6ZdgNrB8yX9Ei+FA2blAf
clviTyxmZgcYCPIP0iovX3w3Ov0HwUWaTTHMOcQ4fn0duNzstmsU24uoyWcQYcSD
RjGxVYix3hrHv7NZ3mImp5hvfKkMU3ZneJhOwpilUvDRRu36+iSRFDvVnOGtJeAh
Y9jWzNa5CiIJ6fCZkXS2SugwkSfYZIk+R+K2Dz5DnQ9zP12tXoTVYBgtI9RtbeZs
SrZO/B8IoKyIF1mvjIGDqvo5vX/KPZ6H6glALsfGSqLMtCd7f9qUy7VfSyzVH17q
LdVPy7zt80oO8YgM+WvBojsn78ZC5DqOeDRICLT27vo9uTEsWABgMA9O3h7TZDop
G7/V5/AM4QW2SmDtLi1o1LK47uhSDmdlTGL9drxjec3AgpvKw8pL7esD/yT4C2X0
JN03MgqlqqW8Saxfi61lH1AgfL61FBCbFdXedDFcOuv6nCLphlID1lA7mjRa0Spu
B3JTI31FqeqZQ9RU8J9skeHFurIFMcZQIzKby9On1mCAvQqMmFm15JdV4P2+hYHD
okxhuIhaHMMogRIlfIS4pch9GZcY61S+G+zci+4+dTvrrk6qETMDMLfsmGyw3sDJ
70HVGr8v2vtBu9HBG+W2ouBWz9Gm8U9Ya5flEecQ0NJbPmPxwDsfd0EcSmiby0X3
TBsCSqefjzVfxlN9ilPB6jD1DVthivuyAy5M8Gco0ge7bY3i9WkaebGLs0LCNO5V
62tDJHILeGDOgHpld8Zc1RkuoLi/A7CzC7lrVmawrDB3qcAeZhWYbS3cMdy2JG/O
bTF4wBXoXEjt4WN/Quo6DoKuBmMguUjRvWTkyk4ee1L6siyCDYHWelhvkRKmaVFN
gE9LLzwfn1g1PfAsU0a99gd2s4g0k4/xoEOjmYpPaS5cE74hkm7VF1OF0cY+opwI
+sdS7fXyCwSSXKGof8Kxw5DlnXrpU/vXEsop5S0LhbCFMEyiASTt5X8Qe4tpT5Ck
/FNyNlzQ1Z/NWcTTA9S4LtGemLPd7t6rxD2yyvql55x/ndQoP7y4cmjwyzOGll7v
Hl490yxzARTz32j5zo73GaP/GgXqiAr9wKjRHtEcfV4chlC5RkgSdw6/AktEEPkp
WgnheI0Opn/v5m2C6vF2NTcRDWL1B8bf7S6iJBKm/Qf2nfeeHb0FTJztplrzVjPo
22nMG59iqNpyVrf0cg8osZBpuTlUMtxINo/IfALq4nOkJ8efNG37QBhSPEgNPUF4
oQdIsgCtLVJbnvhu+8wATP61aHA/EL5e8xEUS/AqNU3rfFkeVMCCjoHikF6lAS0Y
6NKlQRk1s87v2Xn7d4EKkvHUTmRxVDR9Qj8sLAa0O0/CctzcSqv52pwypynoqevr
zi1D2UH6oqo9sjQxtFXul19dSxWOeE2mdejQe7hiHBh9uS6Y/F5YqW3xuxPu/6/0
WSPq/k05GHN8kJmx5ISMwcyrYvAAMjtjgPZyX+ikHagvEYWtKGlmah2tdXWu/m0z
Isdao1LByCDn6grJPhz5+MtYqbukKWuUroqm8RJkfkXHiJltFGBdH7tzKAlaWLha
E9wu8MwnjM91T1CVhPbztflIyQdTNrWZlxzoJX+x0BzsYVrK99cw0XtB1ucXxLs4
jh9JYr/t+usa5zzqZ8DrISvwB7kQPYollojVn205az63lESjrStg+K0OeXboL7M6
otsMuHy7sIscolsZhc6+3AOPoMp4OY6YaELqZ4poW0159htdpvh+7EUPQc3yjHBC
jo5+IDWLMhiBptF0pNNEhgzEcmd9Hlu96VGkudrPMAifmPL8ZFoEyXXZGQ24se/W
I5uzLKUIcXauAh4VX120wbzK/JlJmqiSnZKLeY9ABQ6Jbs4xc80y3C6mqY3xE3m+
VwFcsQ50DbGsggj2vIX9ha3KpB5L+SbfydF90B+njNQF3CLmKHQP6jDRh6Fhr+GS
J9dxnGv+hTnLzrHyOR9ceu7igxacHa5gUELFx6HAqPsEk/358gXl1I3yE8xCG2FP
wCIeA8lU1I9tsbKburIkwRBV/KHDyM5wGSDn0iDIdAPswL2g8YXMbMDrIEvuxiY8
BwWKjMsmSLPW+WJY7N1cy86uZePKRwnGlWcvcx4lu8fa7efZwf/OZLrnQCzSHpwa
ZyDxeojyLM71D00QeWHk3M5mMW9+fdR9Oao+kZSWt+FyeHx5DDonOSKuegLJigcc
Cn2P5ZLr4+YQ1XUFtKj7heUWdZZf/qm/Sy/9Lkw4UmIvlfzXQBaGlbzcOWYPk2ZH
mKk0xjB+C3IRXVDiQMHLlm9raJh3ZmG6OGskcWFhjdUdLhKgKvawo3fCcUwAiuaY
vRTp9j0hFIFy8Ff6eAyk/V80IvFFbSF9XIgFaBskj5dZztmpj0/udhHlRMOXv4RO
5QFxhN8XYX9AtFoXSMju20pXqmcE2PndY2hQ/fKMjGNZoX+naFp4bKxICbaNcEFQ
O4erQmYYU3vMJfHz3yUxf0GEJd60XaokcW3zlxhrTN130GuWQ9Vef6I/2EbROGhi
I9KAC7uump+EZwnLbifLD4AWYKU16b1Rzx1DknVw8pAb8txkQlelg4OE9epob6ZD
oC0TrjCaZ18ie0k7N8YyCF+RwJTpTHlNYRcns67VABZoc8YRzgj6QmVKhKblbZ7e
CFANrzot5zQJXWENqxscFR0h98pY6pPk+xaIbh7k0UYPeoH34nPo0z1+9XXXk7GJ
2jsy1ayy6ZaNJxdIFTyp/fm6TWmp5SfDOXR7bUE6zZ5wKgUzmDml+YNe+IYVarHE
IYa0BJWJ+x+VdlWfVIpHLgXuq3IZ570mvnlp6SzWPiGVyhv1GvWS6Y25rLJg3BLW
7vRKlgSyusNiYYR7d1B5JYe6D57Q9r5CI2xxYVPL7tG3nB6scboGCzahP5gy9LYP
h1NfBTgQdsbD86M+r6+Tz0E0A98Yz6ZMAeuKpBuXQ9RxtsSDnGXOTVyTFDe4isNW
x5+4wIrRFK7GBCsDoJSS6TvVSLEstZZ19u2xgBbHPCQmnCcPUj7zd/63hvFL2Zqi
ZGvTVOV1yYoFu36NRE4x+gBJjpytY/YmNPQgRLCsconIYKJ9a53kXLnmFByulLmL
C+5IEu6QxP+OgbtaG1GBF0bxnAPauT5WWUx/T7LlniNz/zM93EiRAMOX68T3kpD7
+B9zBjp+LMXgevGOvdPPTCtP5K3n00qxnPuTw26TnxzICopA7DFKsEgoR3bPCZy4
sZaDQ0MLCUUGdgyGoYYv/n1WtXyS3uQnawT8jDTHYTfn2xBgz1+Jhs7JtXkn0cub
vHb2Vo0hfsKnSnRPC2TnmowZO3pFxZf/lBYhqfoxSIjwbg1A5s+5BvUn9WUwpo1L
fjA9k9AoQjrFXXRPYEWJquYtIdeQqTmy9YX3bvzHp4NHgBbtEdN/5HGOtvQIddWG
0p3O2kGEubtuu0TLdxOXq9joVPL65i+NQkpO4Ex1XizcI0Oct+LNCcZHQW9MxcBF
+mrWlJydv0+OK/4P5Evu6vKBbmDaXjjfma6SwOSyGesByHBfT2tQ3Puh+HyDlOO1
blUGt2QJg0WF1GJ7QjO8VVozTo/gLWMiVNWXB5/8aEDsPuXYr9SUxCVA67iN6JcL
k0i0UEKr0AOvc1pen0K7lqRG9Tb44GiUN+eFbVqPciM0cDYc95Aqnl9uCb+OfKVt
txVtvW8NqoTXPQyFi68bbHAqPcqUwVpu4iwhNW8ymVGBGqApzKvWUEhZp2YWW33d
Cg1h7zrkNZGmcw0+pmEm/Wog9Sms5Y0WMsM7BvzSODjdzdWeXWdUqgWSmQBZlVzV
8nuakngU3z6lyCUt7cJWdrA6T6/QZFBCV/TWGwquoMxB3dO3k0bFq1jss9VmXIcM
zmpjazmXG2bgNXMtnMLQqKhufXxAcQUBpiQcoxHqPUqxu4/uwnJ6vJwrkFBitAfF
3yo/t7weXGX0l4AP5n+WijiSNMq5+LkcTLUhbFiudLvQU9Xbzi77NdU7GuFcjZ6L
l+gqgqgmWSTiWDYngy+/lqaAhZpQY8Sr1qaVMZ5TwYfyodS5KmZYGiJJ6EU/dwP+
KnvG/+C5rCAbLHzgaWMkKJ5N/z6ahq8NuMdzXaxAdLkEw15UT5hthI8/UWxrWu8T
oASj0RX90LKq5Vz8b3Yo/nQJ3w3XfsRdhJ9Uwc1ATl1AudYBHwGrJd0wnf2M5jwa
fQFfEPNWe6wfDZoQby/vCU1S0AzAzaDRAmDJgo2YYGj99FRqPa5RiTNK6Od3QPrQ
dmkiFbplQyMS2pNm/Bw9jasDoOmU7wAa3ayk448MYaxZeQW7zgw/7lTSVmCJAOqK
VqAOcdVih/XSTmwdv6ih4MCSavtRLWf69SwsYiKdfcUs76xOmSiz1S5Lql8um6p3
v8m1uUu+Ob7rrsmoLVUzV0EBsok97CxxyhU+wdI1jWaiIZSSD2w2Nkf/ZiqQ24d0
0xbcZVxD5fyB2T0D/PUkW5U4lzdDQajUDTrVLjAoj2zwyxbLYdiLEPynC9GTqYjg
PN5uvk3zlIwLtQZ0A1GgFhQfgk11gfMRzqyhg5aUll7h53bsSXT+IIxEsBSueH3r
LR1eF3kB4426bEHNRwJ/6CD0LzGYgCiI5fl2wRxcZ8RPKIf/b95ADvZ3QQOiTyTi
/w1N13kfH9TlLSRKb72ExosI/yL5aWpjCPO6KEFqS75bYHimVyaWjZZRWURauP32
9EyX+VELIigBlwMjyZPDnospa7Thi2O6FSEMiLqp5Ecs3zLF3Okw5uXmOwD/0wUT
rEMKzZeC+fQehwPjCQt4D7iEwanJ1VKK31ezVo9MLjzHOifu5cD9fhjKLrHNAz8D
18Uh25yF1Fr/MZlqtzHJaWSpsMIh//ZCRVvAFUfoS+Fz+z7BvL080Vq+Nu9TcWPU
kfIQDpaR4vWuRnYEre8p3zumPIKShhPuqB/1VFoBaEYVClRdlrb7tUEBIMLgZY7L
QJdhQWh76e6lry03BKhYqRLQLdGW1CFvwPuaNB/1lCU37fUkd3ZRs8P5QZpgJIAv
0ZMqLscSGK5Kzt+vHAU2jTgaVxZc0BwzUIho2as0bK8uoqm5zPuSl2IGqKbZDqwv
pgr88zf8xNBqWdWVWmIBHB4K+pykJMa4Z+H6wFJPhgXAwGZ4//GV0TX4NnbEHWRw
Prefa5TWUpfitUyjZLNzUCznpfN6HjGrGpQHNK6uaSjnV4P60gqF5AR+QpX67nPt
7vP+gfRfdXjd3oVJoaBJqA8M1B31+vGw9PUgdQ7byBhHcccrRK7HuzVw05c4n9kl
YvTyetLXR3/qqZXiQKFcc/Ci7rWiqGNiKY4hiw2eCNdS2LwA72+Q/h8M01mYKcaa
pYU8I1GsNF7biT68kKfJgWHai8xxUag9W/vxcbAgnXmCTNNpFVKL7VPFGDLKhK1j
Ro71y6B3HyXoE3KLKMTEIvCR+/3nuoU1LY7wROy4RtaX07gBDng03t4oyNo/WYgJ
krAvS6yrqamaVVuyn8aHIiVqkv7Q50u/CMW7mbQc8wQD/PfDsz3JczPfnf4O2Sc1
e/ZnmCbYdl/jOix7vadnGZbOpouvfbtzk5YawBYZ+98l7DVABlMQ9R0xZnpeji1E
xkWwXox0XaKjwRChl5EtXrF6UYXvrlLCwuKVsArklNetRwDlNqPNkuNQ8t2m2BS0
Q4W7LU5hVxi3rx/PW409Tv9LhVOvteOW1EhYDmBMt1rsjTSW5D5lSmAGIoUeb5jk
lMw/IYUL+or14OLIXdPoxPO7S4XCpoWV8Ho4U4nKLhjXZz1JF667dqnVEJbagDU0
hZJmNgiiQiTX0aqLKKnCtwwe4mwBtQOY6Zj3Cc9P8mChfZ2VrEK+9l+Y7RxtUPp7
HVkjOVMi49b2sbMmNsc+Z8bsxxWLwSBGMC3uPFdxsJrwxZaPLlFZwUnnXEcPkS9T
i5uboEn45ATyPx1WJmEhpnubgNGoKwBjn1p9dnWr1ClXZKFRDI92YV1NbkYAcWIr
YIQ/uMBVviRrSnUI5cDqBWgTmaPPl6Nlq2v+viZ9lWqAoGZOiZ8gfIrRDUzKTSlU
AoUNWmS5SugFl5+TtUjWSt66h0uk+POgAqdT/Gj8Qj9lfBkBj77Fx7FSd+kgvC59
y5b3s3qOTcTsUrUlmaUREQp0+SWeYVpqDtijjr29NZKhOKgNY3phMIobVPS2hIMb
MrqeHD6YI0TOOTgHR1qL6hXAGqXVHAHCYevSh9M0RLvfQ/xu4lDX5kl+7n8EWiIj
fj6/E+ZbSQ/XVl4WpGzYlQONZDEzFu6BhIbpOXIQBCA1ZGA5hqoos9JhkWMK/kLl
xcKYGeW8Y41TlprPXlbZltXWIkbsqVGTjYziTIwiw8Nohp6pJXQjldJRU5kVySTt
oE788ynPiTsJ09ZD4hsXXQ6EJRuVW6tQhWjkYxr4vVP8YTmzDc28ae9QV78yMrHk
+e79/Ef6VaPXQ8M6+s2zR5WhaJeQHeWsU9ArjI6k6ZnmLbxW37yKXHe2B/WOVEMp
3bkjiSHxYSkXxiMuXvDGX/cO1DEfIB3Yx943sGzeY8gBxWUp0Or6KNJq52e45jqR
9SfQ36imszzXTjXdGi/uSBF6VH+ZnBEpDxApiIbEkYy4m+H5fiZroRAIY4Up2h4I
0hxLr1q1GH4EkCMDipE9MXON17LfjfzxJ5ZiC9tfP4SnuWu1RevDWfQxACcrWgT9
668BaJDzXYiMCTx3EK3RHflrnNAN7Czbjd+MPQwgnDw9G/MW9u1FpkTK0DdwXaS8
truaAhJzWDeEB8LFp4SOYNTJSCXdeJvCQVm9WeHq8rkcLVDP/6wK2yFFyabaqeU0
al1Bme7aoSEXOx9zeOCFzy/OSX1k6mmi/6L5MT5tbsFiBFr0xZKInvksEGvq+fbJ
S4p+IR5YXKSfv+CbrRxgA3WtkSocJYeOQ0NIx84ObRNR8H6Mpi0ysy8qrHJQZpPV
lVTU+si7+9rLcEmhDu1mK4lCcSGeIREzKB6EEYPbO42/FFWmSTkrFmDv6+XQSYjG
DS/BmW6lTT8RBl1rp+rSSWLFRhP1yFrt9wzQq8JkYL9/4h2BVk+hDZkDSvd89DdT
d73VaVVe/JVmxsphhMc3I/E7wt1x/A4hPymCfM5fdZZ/Eim+Hbwo5PPEXljKsFh+
SV2Xwb+xnm7V0SMxcgKj3rEx6hY6M/6b1T563fUmHcX/Iijkk9i6PhAOl3nY7EE9
PCV0BrZgcyEZXHxdqPIexlSJyhCrn6t+ewFEmVl0Y671JWC71O1PLRNrwGZIT69I
VW1SLtDRQ9oVLfebrwD7SX829yln6bDC040uZUjeOUw9BSCiok2HpicicafvhdOI
Y08n7VY+rcfKx0uoiuqoDyBNSrhE599u4xqyOYV/BTSr0lGKnt13ZS4hoa616t8J
bEvxkyk3Q45eek4udf34ZU28vSTNM6r/voh2M9wIhrWgfuxlv0ufF1F0pO/ZJ9EH
gvEiACZ+Bf771UNRLjQTRfCDCV5ZVriIYY8ZAk+DaSwx+YCQS0ftFDExwz6XDUMr
DwVOwZietJuV7kAYI+hJzE432dg/EJM9MuaOtUM71ruyaph++1DOrQJnx9NoOgA7
A/fjss58jYsxb+wa3dBN2lK0v+ee/teB6apLGYZirCGoQiUQ9XOcJZUx31evLXb1
Bn2j9BMI6iq/Faoe781ZQirp9cOOcyT6mUO23uIbliNGhQ0hZDgbJGV5sQQvYXCx
rGcOtaWUDzcLao53OrLb5R1O9FQ5LYwfpSgblVvhsu8rF+EtEOl/Xm9W8HiC1QyX
NGdkaMTUZypv8OOB3RHdd06FAbrZ6Z28aX2IJyjFRyPgaMQpp72545eDgDCFrcW7
dEG85X/ZlrweDCfpbaMGdri22g7n9GuNBaOr4034af1p3mE7tC40b3RMvwy+/yfU
2jScu1z4GcUiRr2jIfi+aOwA/OpFQvvFP2tLKP/Xf7aktD9MSUPZOXNvy/Vk8iYL
qMm/EzJRgd1DtO6qWhCZtMb8LRcwVPOD2+E8HeMfcV3UYLKaQlRdXNIeTe8k8cBB
Ntr4PkCACnQO9ayFDijOvriGVLBA8YtAd6qANDmz+QNx66+rv9LmOvvkzG4nQOg/
Z8mhOGT3UKKI5zsOwAGVHyKMcNVLkjpgiAjdyG1NZkLJuCIkorqkRJ75u/lG1X8p
OdjcJ5lAWJu48A2AvJSK3U1+qhi5AJxhBcYHSXp+Xw226E0M4+brbilWLAdpOx4V
gT5de1cJANPOccPrgaKopSyDiRM5wH+3c6x2ubibjJIEe/u3W+E1qWgBoYdhFcne
aQUroVFd7QwWXoEk9yZ1R7e0SkfvgN5Y2elav1vAIIDTmHXR49TuKpuPf6H/dvX+
tHwRliOfTpnWoMDIxaVkK1Qr76gmnMm2qWuPz695ele+aiTzbjxfyviW1f5aot6a
W0/gZBozF6wWlF3xo6ShxPCwY7vsKpPoUX23pJVENudu4CB85IwSdWmSmg+NNJf0
Rcm15N42USOv/hcoiL3kv/uV3akWvb1jCj/2Y74m9ulN56GbqUDM87dLdVw9yKsO
BZTAQwiw7bHFTeahlRP9s49gjxxIj88V1QGymjKOozRUTcbxHI+QrmOvk3aZASTF
wLlEk/VaCrJxh3mlvT3tnrM4BsFXNU3PzS8qCGOpukIg8S2cQ2K/g9AWXiFfOMXR
HEcMhUzWk2OYvifg6Y7a4aXAFELoXBVVQBDgirDDdqODtSH7nR0zQ3jLcbFz971i
4nblzdEJhWLtvlRY31ov9u9y2ukNoBu1k/Plcz9FC0hKRVFqQf2yHU8DQzpZBfSg
PRBLk2zGnVV0w98lg0z6cTybbGE+QjB22w3q+CvoEOqUoHHaxqllkrPPpYkIzKfa
U2hzR76EVqNLMBgG/UDGY0wINf5N5/2Sph1i1ZwPskGXf8v4rTWH04A7X0sx8bLc
OjUof5Z9PO8G2fJ+Oe6gwy5Oj0Ekk/pmidQdtMReyQTqFFtJYuQ5w/rIjC5Pjo96
818xkAQ1zo7Us2x9iyIcFzuQRMNBeYWnvyRPo8Aq6SF8ZIV+xnmYFtulctcOQUdg
+Qt3EXKIwvWCDMe78RsGa18MEy+gIcACRG0mBAR4Eyll1Xsd1fR1cYAMLcJIhntf
UZE8mtHKkX3z/2j11vDbCLtin4C5++fGztlAbPYMJ0C7ZNmZhDxI+fAWEadtZn/x
QYYPM8lwwmhMS/87FZfzB8m9TY/ZKGKLK4NED6uAB2XJVbGH8cgmbRaN1hTxG9yT
wuI6fo48BFHIksTlagM6rX/TXg03Dt7X1tY7eSnj4zJXCYEqjghi72TshpJPDbsS
Rl45i3BonfKNi76Xf98jcYzYou7XbUK9QJ4LM9jtaUmhFA9StjKEt23Xx1q8uxdj
BwsS3NYto1AM9uQhm2lbpMpM1r00jNdqavmSAQacER82v53a/08XdAXF5mUsJvxf
XIx6ZG6GJITWRj7iCYqZp1nxvT7fRsyeFzm0KibvEbtfzxDi3obxlpUBs3JOgSsr
sgOaI003QdJVudT+YAhM+m3ejzvDa55nYmB0sKoZdItOM33tVDcigYCqaeY2iP58
sufl+svJ5AnDUp8ahZvLHBugPbww6cnlAuJKKCbCagFYQvNORjCdfM9UWPld1SXX
7hTC5Gcyusj4MqcIlH+9ZuLvmtUY1gri3MlkhhKTIbDj/DMAtZY7FXMZtXZF+O4H
e64FHPY2RFu0uHfRhFqpyKEJnpPCif/nUldFTEirMknDgBC8Ah3YJzdy7jS4iVKH
eFGKwYVTo8/mYTTilVDBzByzRIjV3/XlOD9EQZqmPuD3Z+h5SRRm9WkY83Xbwhct
0DSmBBvRd+K67i0mQJJm7iSR9kE8ylH1KF/JlPWhzaDKErfxACeB5aoo1BCwUByY
GD48pwPABCGQzb/6RLEqyKpbdIJE13QWOzO7sTBS4Dq9HwtBWnbFAXb2Z/Nry2Lp
tid6UNVAwKQcVQYEZ7OL+IP/rnzVqBvjS6QwUJd+vSjync7xzaZBS7AbrKEcSs90
u9wDDFo0/bCWYSnVeaJcmmpTmPJwE3Wnh/mZOcLZtPjxwgJ2uh9P3dFKykvtXFxb
Cu/YCZSGONP9tgC5WC19/kZloxiUaiSWi3v3z2dIYQHTkg64Ylp7Djc+gLRQPfnh
8IT7oGLeGkj/3EuhjwjnC7yAZ0vT3ZXAOC5RZMvvC4G43bNfsemgQgp5Emk6OwYT
ZT5c/35kZcOoMonX4HPpzTN+HGpxVpk1HiDWuZMwquqM+1Z59PMmluDkEHLicoPA
QV4cAJN2yWFq1wjcQhHSfcffTZFXjHhmyTIfW6uHtOhKiSGcrWT+Y4wuJpxYlEDQ
d+pK5UmZP/HhN53ZpGrd3PGQ6AmBbuzf2MbzZmr+xj+XPAt2Si165e4434Un3kKZ
IHfIKtWgcK1AlQzVjD90W2UEUHAyvZ9FNuWLetFCEHkAs3KRAVPJ/H9wjsyqP5dQ
mGfKYx2gDyP2VaNSlZC3IjPngnlmIjEGiKnCKzrs12Mf6YCIRGnYtpUS+cTXmTp+
ZDpC3/9ng9v6KO03RalSUjSa5jT3xczSbHSD1vqiXyLR5jSI8w+qgNhVnQIlnF0K
ZPZOxwwSS4AGSjA++yUI3e5utRTgOCd1k9hOxRq4VYH33GGhlLTjPqf31wDL5Zjk
NhA1OHWlC3yGeeCLFxTan48nRAlWyuI0gsv5qsWGVdmoPiiFBGTOcOyoRvlGPJA9
i7LvEPXqMGy6d2x6H36FHQOveR5rnz6wjeUVKd+9NJki5l16qOzSg5vbCucKQXLw
0lXz/kMRzyvZSeCO7js5cEno848xdpgfwdaWs6k/EOto4MOOVE8sn0Q8ntVrWKyT
vtPiMV7/8V0BhaCY6Oeb+dL9E/y6yi74APR2CM4xvSxcslIWZ7ztFJ/ZQR9SCmYy
hKi51BfayU9554/CgvcuZ0findRfb+vV6NZsE/PBFkKKx/iRdLCwTjzMaWVWZekZ
8fXmP6pmC17oOqUvc16oUsqw7uuZo0QY/RSfL5PYMliclvs7ETatN2NvbjWYpsWC
2dvijorMtg4soq8j9rV133AHURhoGGr9gteSW8uuzeQZ9BOVuqs4MupJpCYeYNZK
7T8z1yiBNi2mQFmA4ffq+6Bh7rMdwuC7g1FrzVeOOLS+jTgKpu2HxQ8gjWnrLtRH
F2fRvfwHutmqErGZs1xJb0w+A8ShEUtu6EJxg94CHZ2jpAaRDd0eUjqz5Gj3lrws
tpJf1SCJMqCmGhPRzFQYIu9P17cK0YfH/o2V7VSbcF77MnGzY059wKgpoPuqJDgV
nyzrbqPmwBzN5YmFhoFFmdgOGVO3c/FUMdWOy/ApshbqWmBQc0Eu66Jhh2SytYKX
+EWh0fvNcG425WDf3udiaE/eWMZlX6Mn/Wf/wOTL1bZJuNEC/jdoT64Qp4cshPh3
h2Sf5y2UnSH+NCriZPUGDf2MJnncsvXgZXwymdI5amPHVilbNW88FW24KqFKaPp0
fen4YNSvbbFet2CckbbyCzUaSxKlfoOxDr+CUEM7ZqynDEOTeGpqMyuS1WCvJSDt
nhcwvVA/FTIk9uYcaTpMJfjr1CNfrlWQ4RmKhdzcC0uYCTE8ulP2qf6npBDTUeIr
JqZJA6SNFflNm9a/pLtl5a8H8EVM68ln4MFCvGBmbsuzZjibQtmbE3nEZsUcIh65
+0KfJ9Au3opq8VqDdWpgx82eI5wbP4AuccrW1/HJV1rKq+Z7r1JO0niakeYwDa8i
YsebDJmRMAXFMUVRthu+9zPSTwZ3ShiTXfIuvCQ5zkeWKQ9aBhiTPAjszv/tyiNA
gbJWHjtyWY0bdfKX61jUt99m0DtieBn5o86RIbKh+Ubm1Q8e6rgLiqqvORBf3sEi
IDkE51AFJ9d4wIOXTfnmRUhNfF+Vm2Jy55Tj46+jaKZJt7SfdvUfXf4vl0BiCik7
z1347iZvRrN1pzpX/EgQVC7EQyVVpFbopQNmXn500cpL5/5iqXbUWfK95BGLlq3z
QwewpmXg+kVauY/2z1h189YIHelT/XejKn9/KbZv4puPxXwsDaoil8Qh3nHbm+ln
fXqZWwvH+3sxCaVhm5NZgckPHwibfw9obfMUCyZIavRbeMfh93vY4sUylHoXhcHJ
QNJYFH2t0Ut9zMd2JSjkvp/A6dcZvAhsyCGTact30w2nS0Q3/O2Coh5xYeybPzTy
q5i3m6d0UbFUA9owRJmyasgFz68mZHMNy886csGCIFl14EUXT7Th164LfGFCfx6F
9Ll3e8DZ5UfN4XeqE5busqMRqW7otPHKayEg0liuPJXxbMGRjwRY9gm31Yscpt+n
kWwLCKaO+G7MzLEQw8Qxod8Awbcki9kbKFGWMJYLvs+DqfDLB3kTiJSyIJlruLSY
nua37+q5P9BzZwG/qE4HGY3uI75zIz8enh6NUdWQ1+7Q0UBHj1s/zZnzs+9pdhSH
OTpoblJ3P+9nvqpo8YZ4qfHCkEKKTylIbfBWnBtTrcEi6DKAyBqjC8TVxxEMmRdd
g3TxzrM0nS0jRjpDNV5RGdCaTQZfPVd8I6ASXFFc3m4erxF8SmM4Ekiy0oLFu9sH
55kNSeqkb7kYjgbCNejByzP38bJmdjbZjYI2bVp44eNiX1vVPMVBeppGLqdDyqNA
Rivm1kZ7WBwOM3V3UWnBeTmaFVPQ9byOiuW1aZoFi3A+bTD5x3V9mkbHooGqPzPL
EpMpxkQOWzKf1q8Li5gsGxqRO3a089IxTrwJQkIAt3wlv8LiWz9OW60o2vaCLHEe
IgpAMQGlGhS1m9OFCzWF+1dvfkuRTN7VNOBLz3N2WJhl3eQkRACQNediwFkB1pMh
eTUzxiK3vvoto7wo978mqjBMaPElw7BLBN/Y6uHM47GoI4Qs4Y2nOcI84e6z2mmu
L/67Ah7gKEKGK6VJ1owDbjwK+NE/s8b/MAvpC+13sqUshPGYkR5vlRt/BUZFCMf3
tZXl0PTY82iK/2HS5Jt82/y1g99joTg2KY8uLKiYtx4EacWrr8Th8ro+G3qlhixs
OeoYLG7gTTYEqGFvOu73194opEeejUcWzuNVSXI7XlRQPQ1022IJ3FNIbsSJstj2
Y+kBOw9ZJ8jdrgz5M82UyvCBtnSbGgkgAcG+XCeKZN26CclxV1my+SymY7ld2D6h
skkOCSYcmUk+iLxsYQ13FCNiVe44QgsIY6tzbzKQYv6mP/rSozfbweELlrlnzi6V
fiqgIOSug3xbCPcHRHq79XbF2X81UHC4izunjyAvL+5DkaRXN3qAlwfa9FVCLxsz
o7qFkT4vtHsJqRZ2T0SUwxbaNDoz9OS7+AqaZTGF1OyEOIP4NuT94/t/uveH+SBm
buaeKN4kNcHidsr33WfbcDhgckG2ARHcm6DM8V16HC4qKVWsplO9Spyx9VDBoZsK
8nP4d/oZgZEaTqWeXJwgJLYbLZPMICYJO8wBFDY3yoo1nV6UZWwLGjkd7IWRXS2d
XBTHbcDy1dB0A39gyQdqcaPl0DgYAgJS/2lA4gVbuIX07t5GuhIURWAws+vmodA7
YXitWuTSxbkBY+E5mmdmSlexHh/CXTYjbwBFV3ENObWoFumwBJTapBgQhz2oozyG
d0O7SIEN6VJa5Wf7hwLEL7n1rU172lGYZgwO8klWF2FzRJvZrNWM+kXDRZfAt5qr
cy0Li3RfR0Fx01fiBwNs35PNEcz9QfTMKCk8wFWGFCV670xHhfpk15PwR2v5Te1w
T7R3TkdH2hxjr5lvZeGb4ajvSzRovQcrJyF/1HdleN/ew92zBd2dieVQCFMrBZeU
WNz4W5INk556w3LRHSiqxcwTA5Sxr+QtMe26F3h/xd5U2cUMGak93FHsEvP2w52F
9TerGMUDFUEOwtQ0xNR81d4joan1/f1GqezmJdMoqR7zEf0zmVZOZowU41/5pDpj
5/rdMxbToc2aZHFBBSzqoZAF39lX9daAlaz5juiw8q5WkKnqE4t2ZCzWJIkloF/3
N07rHoLg86m+phEvpzqaEYxPMXW2ILTpFNE3IduuPMyuN6K/eA2Hz4elpclX3+0F
ie/FuLrMC6x6Z55q4sG5fcpOsOBjRmGtBsvKuvuPdbr2BPVZppQXpLomAjfROGq0
62q11PK+PsANhNEEM6g2miVDutxhtfobqIPUBFpm5dPkx93jwvahB3AbYHTCO8fQ
JcxyiCPZwiDKRdLHmhap41HAIrx39U+YcfQp+h/18uTOSODngQ2TRkCCeIb11Doy
15xXJrBLzZJhx1ltQm7mjYcU3ICtsVF9FbPZuH54n0GQru8FlxE1wRV6qyrz0BDC
DW6XBdnFzRl3i0ffrOShu9JyKPtVASgTOgQfjAPV1aRyluH0sodP86Ev8PAXr+3x
+FH+at34FgNOdu8nHxSnJ8KNzZb/CzhPKcoFmPg0jc1jxht99hvPcoh9mnsM6vVq
u7OY1Q67/SpzTqWOU5etsXQN1mifh/GKtSeBro5jU7pw4dGN2wzqh509mdC99P80
/qhh7G2Bu0KRilCLdwpGdu+1VJO+E6MrQRlUmZBQXnIgK0xS1C8yxFI1tHaZuxpy
zkuxn/zWTI09uhg3/3WmTlH4Z19rqUCi6TfKslRlW3ApfnGbzXN98hVmvCDh8iu6
49E5gU2rarvfqrTL/MO2qtIzuMYuSdkg1jhHzwe8I/dmBcgMkyEfSg4SS5mfq90R
Wi2mETQMHVSI1YxI2ScYJ2KlgB5iiA/MujxnO8Te8dYBZSehy2xATw/o6GPsZhgP
NMdcijsdo7tIoyWpJ1P7mklOGgEc7oJNeQDQMhKu8/FDCqpo4p8Es/6xcPFn/l0B
NCATQDpMYzTkBC9RBgosVigATwoU++r7IXkfnvpaz5Y0CzduikPZsMUfH44AgR/K
kXFU7oGhzN7FYG8n1ebf2zZq4qC3ORwf+hhlydEXX6q6dTvYs9cfImx/quV+260a
ecVS+BMHFXSNXwsaBR99ctWx/WfIyfkMq6TTPPVXmODTa+3C4NOabVN5e6YINBMD
tCbkTmU2m8Uw/HbtLM9ud2hZody3IxVlqSrEgbFXZcrbFmhU1iwpvF2jfzPZ2l1k
t1jCSK0bZvIoIs1MIS6l1k8ALGJAaTtnOaV5faBcrNgOP08HCHYCjO1OHHQVZ2D7
lhdKOCN5ODzRmnzdkcCPLZpHC29o51x8OupTEI7YsMzrpjU4/rXq2Ogbo7rrUehQ
JlYH0/SEgbB1msdSiew36IUpDn19wUuGbubeMFdm3tX1O1e7vam9UfAGFKwhHF9P
6sdl6zCQY3TcjfVCn9f/Y65qZN3FnqmPY91uB1oTPj+BbdkArtLkpkog0bBU60pm
j0B1ML//ZEsr2AlTPf3rQFysTDrTCeFKXEZi/m+ts9GG5SHgw7fUxFT/eEk123iu
e78GVMSIvWBZaZlFno7Dg/8i0HlhZOEGoPXrXp2QRvb8J/uyLJ6cuPL1v9Q6Vxoi
C8FVX7/BTYYFDUrZEdYLQOaP3v8MgTgZJRiSyR9YTSLs+vS7/0zyuUKDBt0rO6DT
fat+/LrYfaFHK9XEIOIKqky0Y83z7bfHmG4lNlz1T97UvjSjJ6skbE+f1e8wc0wP
tEWnAYVFf1AQY5mPhbFmVv+ZXkhCCixCD71TGgq6TuiBvYjuznVpcDbpbLg6/ppu
Y23eRUQURGlK7TQFXSXJdK683EiN/HRD3g+Mj1PKVi2Udtn3wyum7Ul/s+iZ/6TT
L/Jn572g4CRBmmrWacgdr5orpnt0tfpR/gMg3Hk/8SdzQx95WC+vmGn229GCPwAu
0u7Ql5MTp4jkjviCMNptHJd7ttxyGDp8vr0wmQrdXiv94CaysOK7sFaLmCnG5hlK
L9r/nGOrSU424EZtUcYuY70rhIF69N4t5GnDmGG7xH1xXR9CdDFq9G3xkF3XMXa2
uX9A/2E4zg+hC+7s+P2y7hc9kgPOCBSz3ACX1ITSEjY+A04Ccrwbpc1hOl6NPw6U
9L1yn16TXb8QPtD4ChSYeHLzhnPL4G9okvjCpu5gCDczlwg/cGZ7vgtDq8xSAYY+
3gmGsA47jZ2zw7qOwUn2gqDBDdpJ+cUAW0MtQffyYG2oLZ043vzz7Qkzb+F0iEvX
fhcPSdgyWlokNoz3BV4XIwoR3RvUyft8zwam9Fios4FMKZaQ+Bfn4nAssUw+a0i4
X08zCjzRbTKcApY42EeL9y4VAA4DE2NN8ZICsnxyqe+q5kxAk7pz9OfHA2h4+VUj
xsFY0zKI9aRtdnFjdNAtBvEZyXz3zZhzecEVttr2RN0/NDfXDXdltBrdtK0fdKEk
Lf7aRcRGgeYiyzCTZJuNb3v9qvOdv1yeBqElzwM7It/6tN+XFZ+afyBLoGyac+kL
xea4CjRtWefGtMIIO1hBbFK/ZZmGpzHfBP3VZd6D7YH7qSukX0sh9cqGJksPYNqi
cSgIjNak6hdt/4BM7I9ZILODH0AmCNYbQvVqcgtVxgGKzxrPrjdIZChKGJz9kRDW
m8BhBeLkX9PpSspdBHQ3mprx6bZYu3oYQYAyxC+w+c8LDOT+17m6Uuhh13fKIr7r
hj8MP+MAwaLnGOqzVfVe9XCan/CVSETh4CKu/S9I9tZtwyJLRDiZMRTIAqxn4INY
fiYA1uN8vkk05Muks6zewtpV1gJyRVX5qnBfi57gGqzfDFTL5W7Ud7VYwkdLZkFh
SU7xjNt1XdfP8LkZ5eRkpDfIuGY62kc4lGUL1w/T8gGSjEMCe6USlYJ9vlntBuhg
TnM52//BLfgjWqQSE/+NR8XrefFBWh3KIzMZ9aCv3Uen9OJdTK0RI62OzS4u2TK3
lpgvGtTUqo72vBGhyFyjmb5wL0eM1apiti+FQYzxOMeyEaWIf4qd2B3ORWSFLAQk
wK29lpbLyQw5PRLQw7LzG9IWlS2Adx9yM3URD58Dt/h2RkVxWSGkAwWlVQlXe6uS
YUFThWtyCdFtxTfzOKsQKbrtZ7Ocj3GGJ1wyVaSqsekf/smghHtvbvskxkJ3JXhT
EaRQBcSRMY8dxl9uz++lYUJUaEvyY5NSqU9xEA5PB9vr0zKhSDSqz74gdTIpyjv6
jxm9M7eJvjWea/4y8CJh2nDcj0eqmBpKY7Nh8h6Si5eUrbWIwxrnF9AM54pJZMdH
nM34ZDXH9Qe2hMpoPFodVbnN3LTtiKDB1DbByX9pq7oC5FarMclV+ztoAfXBNFc7
6f3Ma7LyBuGp+ocYniqFG2RaLu0ytvMeGh55Weg2j/Fh5L/3AyCgsqrfoizAISYf
xn5yeu4p24NXB1c3LRA1Ri4stAC+sNIfl9CPMxOPQQ0pHS7NtdgnG8Ed2IBxcIEt
sTqNePAQIzYUNz5dvFJQItqqUEcWe65E0n3lXtMWzi4DRwGTOXgAZ/jISzMhs+dR
4MkZTp2C6FcFouDBA61RiMiRrEb+nJyydtzq9ibsbHIg2Fzu4lXCxT76YTDtfXCy
rSUKFBgdDVeI03W3eV7jZXpblk8m+Kg356naDYvNF1lyVONjbOx4pi/6iNAI5ArP
qeXIN38V6PGOIczt7WrkdbJrEXpPE2juPbQppbJzuL6FTTslZwwL4cE3pchMazVp
n0gbMWw6MmLjc1/rqkxAIekHsDOmg13ikAb7fUo75VUPx2hMc2rAcPB3/BjfwGz9
V+wvfftCbXHaSUFT//t2WhQini8F1CxRZHgHXcNczq3/LopHCrDHYZLHerXpwjiq
257kdp0L7WfBDUiuD/MDX+dDe0EfSR+/7eoD0yxO+CkrgXGe+boKosH92vRx+b4o
FTaCdpyP3Zvz+KjBnMNl8+/y4qY9x3eGlIgAJ05drnR7NMiSAaYk9MmK9xQbEhFc
42qLtkmkAPkPKZ8EjfDPJ0tgkI7BW2I+qIVcH2Al6gvwB2maqaUgE73vYdKQee6K
+fS9HrNVyw/6MJYt/knf15nlPUCfpKDkcdI73xe3kxE/tm85d6woog/0HQWZqsLF
TAnnljf2cD2c+l5KLVXlRI3vmLUrgiMbpqqua0tLvqVG3O8e2sJZVzX8grbce8M6
wnrjYHp39CjTujbikEUsE3w6aFqUADlRVCoFuclUr4ZQGyKeDPyEX9Ow9TP7Hali
O2LPwMhrss6as/bniUPLNKXoT3uB3fTKVm3EEr0WlYR6APmhyzAoecG5Bw/u7vhT
UL4cP1SI+VsZWbFsGyZVxHlbDlNuHVsOP3metqMds4t8J+maLIj+rM3h98yRXvjt
OinLCH+Cdz1gjryxH5cEERb3PusqIcWFhEYeLNgIEubKhrhvaODUAau59wk+++2i
WPLrYQ8dZzrkoKDgfq1nrugJnX7zIbabCwyuvhDWwckUO+pkU/3FOtDOfefy+Bbz
ND0ap87FQgUERMJzckbdeLhkgUA8fs6IvyygPARlLnO6DOZBLUR7uAbhXONxPMcI
TNUid8zyxJN3BjO1CvP9LEqfQTinhG5vfdvzCsJL6FdQR/mR6h6GMdCbpp6No5aS
JPip4wW4XwPOo9pPl4jIaHsiBCj3blT4uPZW8SfiXen+3BwoPldRGLNr76/iUB92
2q1viisaTTdRgWpWmctekwkVuLqfCOQgSZcmhsi0EAPkD84oHo4eteoBaikqkJLf
BvHr5wm87Jd0PURnhwGvH6BGhjste3zKLfihfkosMY+mTCBc9p1TjegvLg43Amrv
yrWo+8c6IL7vvxDI1HIGYyu9Rl3GB2qPGdYGG5D4k8lA8XkJciBU9IGxBan4hQbL
iRhx4nBjEAYW1Aa3DKA+uM9PjXqaaUQhOBqlJHgdrGs2o9Id/NFRF8ZZXJG7xjmp
44GMa3nD1RBDh8KkaIO3FF33klhUl6fQCUhAbWomB8XgpZ+ppioSEsrLF5XtAEqr
Wvv1DBPtykzr7BD89aP3cpP6l0k+CEeUtSstWksxnaNmTZJLER9oZLbhhzZCbnN4
tiBsAIBQF34Mxd4YJwFMIITjodpP1No0AMh8TItePNuRfBygOV0Gx1TdI2OodtBS
wEOAVHrZcTfbYGPZgEFLEvahgBVApx0uCyawUerbij4lddLVFSpzWjTAOPfS76/D
I6B5mYadUI+/IYuakl+EaRKKAekz3lhAlV889Wg1ab5pe/7z1qWsP4g60r7dfJuI
/d0SdMq/EqUMlEFXXGT/tpS3E/R8UJH6DaDutKv2U/txGHTZ5XhQ22ySAGftw10Q
Cq/1Z7pi3Rx+S0/uS+TZyVdLNS6Ybykqms2beBhdTPdESzFDISiKnAddui2JkeYM
zRha46R+X49Ebj8SvNTrSc1jQU/K8ToqRaVezRqyN7BpHF+nwG8oSM9Gjb2FoBKV
jDuqc64x7Ie7YWebJv8SAy0b1QNJyNEnOQOGOphUXREy9UCrhdi6IJUA+KchFQS7
A2O1I1xlA/ukd57YIvubURjebzWOzTVOca1wxZO3ejT1xscboSCCTJri9LLRB95e
ZqORT+PC6108fqbbWj9P/lAZVEGfUzXZJL2cr8Pw/7/QmA30GILcLh0FluB91j95
CcQV7iGPlqNYL2wRmTmWiVsbCfAN98SKqpFiH1DfezWEcbQmPUCluUPINuWNNQFV
3i9FCrxgMw4OFyUTLotIGZPxPHt/khI6D71atQPZnJQM8X0WTQcxdgkt0Tyd6s5X
oVaJeuhwiczuKvrwf0k911wLw19u+ij+WIXlwAVE6HnhibevUEQglH+HCmaoK07S
de8QW+S5tvO2DwjhZ0VRQz1nxli5j13FUB7EOpdlQrsTFQKdgKUsLVmJDDz6e4aH
RTti8b6NTQ+8ir795mDehdnOkTUTVb+HP2h5R9fyddNOX5lUI8VH0xX4AgflbuoS
NDBN74B16gCVfawJS4UBCl5HYmuD+zvYjoguie1se/63gsIITNXWNXcLrnBMR/Wp
7zoRVBYekjxr08nZ/njd/hUSczSUYZv1w4dKNlXgwRhC4cDhCVINJX89REsGSXlV
yqAMVxe1DFet0jeU9tYPIgw1myqEk9qSfDaRmHWNRF8hRlgqaNk9ykgnyW8W2dxP
Fi25EzIU8kFrv0zOU55htb3gVKEHr3BBc2/h1GHBeI9Y50o2I/CL0YcallXbzs61
R/xUUD5KyrRShYpcM98sGAQUy4CSoO22MSaE+jtosHRXor+vh624taSCd2UOBsdX
02Emq3A4ivjw55dQxh3SOBhZ5Nfn7nK+18rnigLSogWNT5p5D/qPdAh21H09R2tq
8NbA5E2kuTZcasRkSNdnSLmlnfP6oIvIN/SMi0fw4/dbia3EiS0oB+Dws7byKIYY
qduFLFs37iQbmkYbbAsq+1I2vvaY3lgzMN5P8+F2hP17CHInMvDRJaEAbA7FHVjM
i4Kgl0/WCtCjMm8Hkpm3YvN6rT0hKYBH1imkaqNA6ww83sS3Ah3NJB0KylAo/uh2
2Xjn97/VX78UWku1MmEITw1X5OACmPHLYjpKGqt5e4Nr1EndWNpWpK3WTJQPZ2na
wn7WX4wXkRlpA+ZYl3WgOMSJFaiFEsAnKXXGQplIIVfcmS4RpjlwtIIdyFh0CM1i
dMTwHkyO9W7udDFRotK/wwN5yYOhhB7xX8dObwk06g8HK+mi2omCXZ8YpZbgSazN
56OEtRA09/EoTjCJvWdiFzN2oFammGNx0iedgQ0JayM4F2Jl9rDHZbIcMeiHf5u/
xPnF1kTRRimwqFG2fqtbOYatUcJiAMUu2O8NIKWFkTas2REiDG0evV6rbBiEXuCx
Dpsjv84lEu5vPPaI50Nb2/8PVj0MJW7BtzFNTTNEgQghe1fhTyKtrpywCggwAQWy
7VQzW/+L82diqUTLILaGK455UhEQ3pU9oH7Apkq4IKHwbvxxfs4bwUg9FxlWucmJ
aT0IbNMj/KBw1SjyeXx3lDZ7upN/yrrtQZFUa2E40Wm00dJWwQXTqhSXRf8CmwxW
CvgYVoyp/zagcN2vwjKxKsVKlXVdxvgyNCi4h7y3h5eRG/lG7+dG3r3q/zz3i109
9vQohDE8xqw+bmv8g7Dx9W2QE4cQFk0ccFnwf8Iy8I84f9PycOjW+Aq1fuirrYjZ
hHAQKaqaj/JsFLStjWlk9dC2uDMlfJP17rVDnxCwYfvxjcc0zdmeTawrhViHRXZG
+WhN5C8GvV0D5td6hNX6gyIFwPv/FKiKYDY9lUGnkZN3PYbHezQ3yjz0va5fQKPE
9CZ4hsdb3TQVkvXdQh0SpiFcE559SgnwGKugtwFnHihL+Xh1KPtmmGnrtxdGo2FG
jn80EfNcrtJ2dSRsoiHbRW6WrWpzqCsVLPesV7guXPn99G/XUXXMMKVA4N7+4Aq5
S7YMkdK9f1aEN2ssz33cXN/ZDbmI9HOQGPhbLJxBD1vmLNxDNGo7oLCd/Eyay03w
n47T+RlDXWtars0OJLGDHmGM189WR+GuniZF8zVWOC2eQ4PWcaW9hUAKWk1+7w91
upXZLnyJIjq50xtpCl5F3rAvNlLSX9aNA0S0x3+rQRYa8sf5EJLO81IPItVY38aS
vKczoerA4zTrVWAlFTmanP6AkxMPm+m+X5zpJpNEK/T9SUjMQiBoNKlpAIVBOPat
dVHiwBY+xzxBtZ0dyOUSJ6p0jlcuG0uRYWywoKgkol0DAWKbf4eiuaAGdpCV4tlL
LckqdOTE026xosIXfmikGz2hsfpFuZ9oG3iobCBh2oEVVbPsloKwP0EtZduwzKX/
y7PJ0Fk2pXhuaUcfgFQqdhqOcP2wrSm/ledSoRpbB5mAqpE/4wtM5V4QzwiGhFCC
LHbhYXafkSFFvhOGYjlW614jhi45/x5quUfyO9Q4eHM90RSDZqAB1Pe31lXyOMxh
Js7ThPUjJ4W19tAEnWAUZXIPWOCQ/396Upiyc1coJUpHFsgDZMwHs+bec/V4LbZ+
DPOI/s9bRnztNENADzcO4Db1YEUHO1kT8XxXV4Voy4pC/lf2N/Pb7a4FR9KaixA7
XnQOoGIkSbFk8mPYHu3zOjeeH7TjbPnpEegJxlVmN3ydz9iOsseEGCuirEVLydQY
tXMLILS7K/RlFa/3lgr0dYGB5aCJoyIForAUPJ2E8ZU91QM8LKGg5rGU9HfpO5tH
ZSMwqKnFcI20vY1EEFH2/PxIBMevyQQ2qjmtmf+stEecwkWI5FMiw3Jd11ZLeBaL
ATvwtdoKpZ3/QcOgEwa2UGdZaBYCkv5zngaTbKh6m/BTsFEM6dmc/qXKiNesXIxF
EYsEnVjG/88Wlb9DWQaCb4pwG8M6X+4Xyimbsp5ls5vDkpfwgYF5ZYwKwJ4mC6pQ
UL078xbpKeA/+EwF3oJIHEu0/XAMutQv1OMygssoMAx4gpsf7/FtXH0n9q6ZUGgH
iz+EW97h/IvJszISYRjM5e28xN72jiHxmjI7/pcOaVOiw1fRZd0xkdRdsVcZcbQa
CfoXzAgq3l1Fm8NbQP1I4snYRiALMWpWU6K8FlhSlkRVk21dgqQhJwM3llrq2/m9
8ZNvBLtV3NVONZeAdo1tco2XuugwOE6OrZ6S0uTKkZs+ocpAa/kiMWSesU16TjTX
TmIZOHuUK9KziHX2UigoZ6TypiiGg6wwOAAQyvd3fm8APB7tqKIU67gtcCYMhh4p
xxj8EiTvhzp6i/FNXqRZHn+cQR96vAzsCYpdoYUEKEOqqwFw1P7ImSZNzSFv2MSm
7CZGN3P/EDVKiJHHFmGpmIbaaRXLZ26rh/7MiFETpsZelOBNtGhhBDzEg5AErKLA
z7AZyo3HwzXLGWcwDaDv+OTCRE1GvBY5K5a5hiVkHRgfn6UdkgaGowvtZ4jep5ic
o1Y2j60N0VnnvdjSn+Swhui9vikYXdiBaB2kDG1D0qwBffwdDIQKEX8X4gsCgkuM
0pDyOFzOuS6SntW8LbH8M2JA0XR8FFNWCfI4ZRMH7LbETfbq3WDXBnTKBiNsWqjA
SdaAkUJ48FXwc3jYtxuBzAlMcXuPcfPrTKSu6sgD0SriT4PAgXMnqsqPBN2hDgmM
i4/9YIYuRqLf0HlhgG6K3a/soOQbEgUAp+CXudX2z3RbZIfNveoI8CFXwZnu5lBq
VxgT4ZcUHX1dzNaXkRyCVGxtc4UA5Ie3dDlWSDXStgIOJ+9kQJ5ggDCYC10Y+MIh
eP6g0eB6dfakyGS2p0noqk8eXBexzrBG2s2Cjx6o5zbgQe85KYsGmazpoVcWcZ7M
GjmlvN319semJuH7SbZspwYq6FZkUIdsYEZo4ArZYg0/b1Kp+fmRIqRE20mmAzPr
2a1dbLcY7HGaoRCP75rqLdPVPu0WnlhOd7952+vpbGYsz28GdrBGQVtwLZJ1hN8a
tIkmeHgru5OJ3lnv5Df37SGuDhZHyqLezgkxiVnqlZRhLfJ0PZKZ06OLrfcHWtIb
eYq21c4HALkrBmeeMpyhL+CoBRaGDOpkvz3WSkkvVCCIVWnaf07L8TuMXHkY3QXh
LD6fLA1qH7ZjfiYlirixmwOmAOYx8HdPLelSwSGEhNkahA/NKT7BYW/mgY+2yR3j
D5sEdP8ddgEQ2gn0mbS8lMQTpQxYS0vgxv4H9ZOiVaObEtnMXgy3WtfCsZUZXbG0
AD6jGNMfFxOsWdpU77olrzAEHp4E5flVFE5Qjoh3EXjzTPLQQMXiF77VBBC6Xqyj
tc3HUdaGoC1AoVwkkwMWKOWL7v+97YpC3lVWUwxuwjhdTOfrF7bZw28pmxIVd9W+
rGbLyRPaZ6e+flVpczgjGHuBOqYzFDvzYCtlmde96b1dhSD3VO8BjGxgCofPM/ze
JiWGD9rcuodxaydk7FPTYsKBY577WnIErVEL1BLj71/6jYq1IPinshBokH1d8DvS
resaam5jVhzLESvfbfDjWAFEZQ66QJPE42Q64oEBag7lf29sR/5X0hZGRiKkIEGe
zWLH/k+LTn6RgDZ91U9Qwb3BYS1UZqPVa4EZ7HaLckql78UTPzbJSQo9Z19e9hHR
6Gob/+e/pgQvSpxYLoMBLILBHUTNFaXVgIkgh3Ajy3VuzgIfE0gEP4/oD7NwLePX
Kq9izbivQ70OAYgs6Am9vpU69diSD2bsHr/V74f6PFU1QDNpo//SSRh7XrmCawuv
aDMYlzXABp9O4+T14gkAU914vACEGgg/0Z8OA7oQHK+08Ld9z8dm38xpT5RzwT3P
7doK5nKd6etbrJDDj56iJR640Un9TI5Q1DGrlUkbm7DyVS72GmniNRs8/UChlz4D
vkdzM6UUOcOQuC0zexBMth9FbM9rnAwbQrtI/ZrO2m93sHk5apvvGfBtwDAKDfOR
btGIrbXC/3C7nDrIYto756JAgM6/W6uqRUWmSlfU1mhGsZRUGqDWKPn+20wLtf6s
70zxeSBePO2JJI0cIUjELkNDgwcf35SVaMvOIVdhm4RHFiCnku9EaTqnaxNHXmw6
j4D2Zfo20Pxs0XYRmH2HnBMNycaIalbIDr9cETsNrepDobKwyiYA70EOZyS+ac0c
2bDTjbkXF/0mPu3Yadj8lefACMBGLOahYW3dqUKijfXF1lXEz4czNKJ5dNmNLN7c
A8biT5qO/FJDxuH58eZx5Buuox2xi45QfoEzkE/aw+6lSpaiB4b6O81qVv1qXcRL
iX6ILNFhXU0VOMt7ZODf+SD8NTbBrwcYFf+6fiu+wJJSZ0gLC6Bj+a/CJE6v2DTX
3ygN6SDidiT6QYRRtShOe4gEqm7wFB67KSX11l+eBEmZbmYhBv1HJkNnuNNpE+YR
dFicsmtzPwhfWp3fKREdaJTquYa2sPA8st1Lt01e/0uWQWRvXPwCQkvm47bKYEJr
jHQGAKcjzuMeIpKFvYYFuHJ8162UlO71GHdRMy9LSyeGyGtJ7Kn10ROpGYZAjkEB
EZ70XZFMVAhlgCvOIUyL55/BkOlWGGAaq7GAwIukmQKlZE8vm6N5fVfhlWzWsbdF
mUSSh2exAqC0FG6ZzXgCaYei1H0YFcfinGX8IUTnuGyyFiLyRxbYVrgVjwFzfQ92
i5XIgOkmEZtR5gSmZ+WM6MvY7Er9pK0LFHc0z7Q8MAFk2oZfy0qGTnN7M0PijB/I
MP2rQeWcKXEo0AsqyaSgGnWRDauB+ivCQDFnQbQydPsR9MFkfEUC7ZBp7tGjNTwg
eLaXmp/l6dTvwSWRVkdSb8iE6fkRwgwx1UbjI/c3YLSlndXBumtdKxTVm1SvsE45
dxeXTstzoECebkBtGe3v6SJO4CQ4VXJS1vse46BDn1jbmQoXm5C4X9f4kgQ/ma97
CbCny1K7OhtgHQq1gRIVqXvfPQUZGJWV6/xxFsbQr2eonsfmf8b2GbooVSJpZQao
AQQgT6XrT5ge6sUfNeb0noD91uoZMPGhv8KoDqeqxP5YH4RNTTAlZWIsxHUjNbl9
2K6bBjIuOOPIOtTFOXRTQmMuU1clSKLg6elDvtiOHJt5mOwxUCDqZfM7Nz1rVgW8
XOKg02mlEbHbM0G2CRFUdxtjpuUpueNKWIHd6oCO71tcKhPLPLBjOvQHREOy2zH2
5ArytGietyhPipCul+7uWDedGpfVRmNzfMQMU0jR18w63JPGnfzNQkKCwV00Zmc7
tJzrpbc6/awfBTesypPMLa3KQF72wSQNUMS3BePgLtYgZq9/PYNYTla5WCdMlz8e
6uY6J8i2fF6bjktKXaSGm3DDP0TxAbmBwtgRcQcDgezNt01CGlXY31pIkd1L0gW+
zAzltmFNQ7wPhaQG5tS3y4o0NsmLnbCKfGfI519lkFzyg/lP9UQTunbrXEnY7WJx
iwCAbBtve5OoDGmWYknb5H5oUekTdcJi70/0yQ26mCeMphebSRdVDvi7WSXdJ3iC
YolfuNeJABMdeecC5iH5KYDKO65hpHsSSqEMsna8NkEW22tusiJoB5Awe5N7QKk5
RfxvEwcnwSQA8OvluBZnxOqTNRw0FW0MX9RM3KceXEUsmy3ZUgBfx+NFkk6vpYUR
JK5rc6Td1r/Cf3mL+dVHJs/O2R/xJe2CGbsutr9fAUFDuCqLV+tsChD1djDBUSTa
9vHBGAaMFRRWDM37Lkbvj8izi+z3Td7HXVP2kkQ4gT33Rs80llC+oNKFL9CCeY3z
Jlavs2k+AnyyBARb7CwvbilbJLCNUXbdXSzWDI4yroLZL5WdF5DTszlLuWsAAkRY
ek9GSp7ZJQ5kbm6nl+0PnkBtVrXZ28rtLDy78nUzwTV6KSEJqW1Is0/5qb2VxqrZ
XWY25dIaFetgN5S8OMNrNMv6iPhRFBaqhrkeX8eXHCmt/ay4Jb5Os9Q8NkFbBjaV
CDWUqIn2Si2Gbk1wk4FPWt4Ci70g/d1G5WlssUFFGkPKXyYJnDEnPiShDCjRQ7/i
RRisVKDBd3kvjA1MoawcnA0zdA3rPWwqgJjrrs7VStHioxkUoYwMIp+g9UE3BzzU
MdI/sF3RpD7Ua1PBOjshNodMRuTWyoMbubsGjns+hxllicv9iJ9zodhh9M8iXXjY
OD27RYFl54b4NkxtM10TABYMCPxhVv8OWdbzKJ+EJnp+lsgGnatlw6aACOUWB4Ve
5o0SUVJo7Jl30EFO1dRv+gLUHvNVv4ESc+mOdMo8qkX2gxA2KldV78L6RtfO0bgn
OWZnxn8KJR+LBP3eeG3LOCAIkpBMi0EvL4NR0rWSzOTHzfj57dhZOhZiA2j0xVvt
mBHJQmt2oSjcSy7SRoSVeABwk/jIyJVHJHzAUgw3kzFi6VipOiutZqoqxSO+ACz2
0hNxaOrbyiEwD9fD/PKBMgiHrBjpnp6L3VPRex+GM//qXpBAdziQht0N0hs+LW/p
SGFnULgD2JAx5BeUHCvg5ROtKFghL0azOaIqEt+T4nDNia+pT/FVwqUhLDezlMY8
xXnFang3WTUOJkCyWeMW9PVr3zA60FD422BIWu9JCg0ZvLMRYqwICPRKwBzFomvg
UM3ITy0bFUs4AINRxohR29NPxsVl0+ZQcZBb8n4cv6oBqlMh3l5g0YZ0py/lmXLy
RsyQPrYEQBOWRjN0a88O8u564FQmhHgUympyq6LQccIn+doQ7jnl0EsMKyOF06BL
SbrOJIf2UVCb72eslOoYi3hkliVEmonMcgHR6RZMpZz18rCnb1fZKy1/2ncJFEWI
q45FyNn5CT9dzrK2D35NiOBbduvsUoxdV4PzNbi2P+DqP4UiZwjzjDIOnxpbnSdK
JKsrP191faWG+zNLyFKjkTUf7bJB0YDbAhxUTOUm7mCgUfMIKukXJtGlqCFHlpfu
8BfQN1U1AkzN5GgAk0q8E1sGzWVSKzaTQw+lR4O70bJEnPExo5MtgTP9eIAv7zPd
G40jgZ1l48VxMS/880MIchKhMuLS6fdkQaf066lbWi7YYh1SQp7t2xeQBwSXrzmN
3rCH12lqTvRlsaZmJ7mfV60DCLu5d8bgP54tCkMm+lsDCE5fXSIJLpL24aPIogkx
Su9uIlb7waGXWs1D4kOSxfijYUQeYA/Oat/59kP3GcJcCtym76pyaV4oV+mEhIOp
WmDj9KTESdXQam+IIl7ETDyp1jvvpipiAOzO8RWCzlPpMoX3pGDjj+I5drAunpL+
bgFJqhhx29cvl1rVRFUUVI1C7wuKlRAPYqYnmm6S0S5nbo2a8FvxKeHrPpJd2Uao
ck0d40tsRvtFHDPdrJA1ccxDbpPgm/Y+X36gOGn5dQLIz7E0ooLx7jDiQgIlPg3y
v2Jjd8eZtIYv8qIgC5916U2a6P82HIUeLgK23qnL8aA4hkjG0tYZOmVk+t6Ne7Qm
7KIStt/eDj/mE7HvOLux43looIeyGgcVcWqEzeILcnuNM7Ex23Jp9+U6BzxpHoMj
aFMHaTRsWzwYXpfbPrVKwS/Dm2LMivCEPCtQoonBpDHqlZOqlaPwKZhgQZYcJ3cX
3S7IWApwLsn7s/eKYWQOVbgEfgZYfCB8oxG0R2YpzeDlWGMHAug/D6GOmsWo6tD2
oHx4mW9YLgvZKbA0TRVDmQz+r92g8fOsgUgNMDJQsECP2d2ZsXAyRClGycPin/5t
tEHMJmt3TOjiTRLRA89539k9s1AofCJ8ctO23ngYAUIiOzsd5xbSoZQUswlZc6qB
YpG4k4MrZ8qZzIJJa1Nwz98zKNDFzOaCm8Q1dQ2Kh1aT+abXsZhOsrQHaEIqOMAO
rG/PfZFQ9F+HCOwYNOdKEDkTXZFvbReeGKYkHgoO93HYHz8QxQ1yuCGR53Yjkr7B
cmyzWgZKmfxMQzknm5M+SHT0swXmIjyiUY4ir4BYF1WHQCSmkbYxtpiSdY9Z2tqp
oyDxQyL2cnWAWOw4QkbO/urWJv8AZtEFgC4STBP37DF6xlxAdJg6Cc6y49lyjb71
AjtmXNn0YgXLi7zazo9Lnnh/b0Spc2ui1SbVbrvUFSd2SfsiAW2nQGPaMH1xUQGw
rOw+9yvs6uGcoD65LRS/MOjoKCZ4dGTRP6CmgrT8pyt3K9mj2AtlavQas2gcyBto
f9Slzg5C0vBzUyzbuNTjacAh1FmIKk/6ypS1CYe6fuLuFvix/PJCHEBYenVv/VpP
2xlg+Ccig2u8EFzlYQKqOdANTXDupIQuU2+FL2HjdtfW9O4C7MntUPP6PP299hFu
+SA6538+2sv/nLboMOkVlLKeY/E+c/zjLXucvwGpkX+jR5sb+iZEASfXr2OtN9Xi
gz5N5dxVUXJ0YMVliAx9ZQxKvGm9yQdhfgfffdY0ujS9gIB5sdJXPoGpWmekzCTm
OpUsvfXv1G+FtECrj8iSy9ghAekt5vHpC5ZlQGtaE6Ev1FnuvllMU5DtpEAUlXky
FR+GvQOK++jWCd/Dq+L/AuxrNaBboVGAn/T6+403InjUoKZ8nRiAh1hHQT2i4E0U
RrGRTmuDLpDeWdhK/KVIHXhkdbHTbe31CjyrDV60RrRTTkj2TszxgW88rjFWee8z
oWpkLWzJwlukLP7Jod3WGE83zU2oxuNImyF1tgcl/NGky2xQEfmVOGUsE5W4qQKE
l5Kg39b6JVYIfLLil5qYI43ia1Ea4j3MJHyJMSH/VVkxCMowrW4ZSdQnBDIf3m0e
jHuIDNP/AVkUdE6nPDbd0mKk2HjJYkDWP3endYD7b2arKRFea45RcUs9E9jWIczh
cJKrpKwSVw7t010keAGTpuPPF8PY4bGyrMdLgnQCkkPaScbu45J36WgmXzCkgehL
NZWNgb/PmIVAvxU526cYbggEdeRC3sx4OJDnQU90/TPzkA2za4nekugG4QCW9EkB
HOl/bg/P690wPIwj8j/BPhACaC8afTgdRoV6TPqEDWwQMWAa0coGGAtrcfQMJfbK
/YRFCmWIntRdAzB8mDVprqSgzjg2MOGyzCJ+3ye3AjqMPSlq7X/B4sAhS6u3gGrK
zOtflDfaoAqUPLlzA7ytS4Q4pyjBU7uozDMIKeTjEOkx+qD3o/xIwQDOJz2fDu2q
5ePLHM4zarpGXGxjhmkD2rFpuK4fF3/IuBYmYQvlOgLR4dRtp5SVTGeV3M+l4HVo
UnWzURGCg1xrLMNUpqWj4lCuNSQIe+NcDgiSIdFMbl2E8FexG1E8P7OjupIRzUhb
04mXvRiZuRMCu7fVOU3NKfLtA5JdpK0gqmKlBLt4gvgmBsEUz/2D62JRsqxVPuWT
4ZJ1DJA9m1352BuxEeXCsTO6gXM5k3Lpk/MWm2PJdynff5LQHBDMaky+PvxUG4F1
WaXiLtQYCKn8H6fzhnEBHiMPIcto7kdSfx1qT71JNWZQfp7Rxz8asARtTGQ0x6Mc
iCDSWwcWYz4dEj1qdEdcAjf2ID+wTmHgp50TG7aS/CWd55el2qxmVJyAtnunn/K6
5oDTv684osihzpLzd0pptP2FuS6tdppkflwNHGy1gs+bGQRQ4lsAjQGTVOLUvO/A
v/57Vxa124Wul/A3ci6t8m7nNkeRs8OCipLORq1PkT9UIsaJaVV5BHz6B5wOxspM
tjowRLuI6W4ZamfuLsFGIbCIx+GTx0oK0Q0L8Bsh50F3p6yTByQsdOUkJrBri1MY
V49nj3rZ3oSjXuvExTjy1YywmzwNCSwvwg6NYkK+AYt+FZSwu3Dx96/a8zty9/p0
qx4BTHxZBJHYlk2yybJJA9jRoj4AaRaxVV3MCJZk40uSzKV2Q5m73WswS8EFj6ok
Z2ffKBkrDTw60+QpIQEnUg1B0sGO++f0tf4a6rIXQ4lFgEVjVWgDiTv/mIHhxR74
el6YkVJG7TMB56Nv1FoTUQ9VWLtdCUrXROonRfgxfVhv80IbTW2Q+n42FgpnH3na
y8AkgPDaPgbaw16Bo2BX+AUWrEYjtRA5fIu8mmkFvdGa1PpSXZozDEYXWT+ledRP
ow/JDwpNlHJG9+K/XoQEZHy+D+dkBPaCYDtdkvOsDghptLr0rm4cBOT4KY6psJRn
tdUOaz2bdT+phGLd4bXAaexWGWGBQZVDn10Ur3BRb8KmjvDJUfBasV6kACSNfN46
S8PbCoWXCqsnNMBh7hBFM9oFd2TTtrdVrlXVrzvrqvGVxtd9yK/+7+r5fr6Z6ekH
dSE61/Hbq0LkBcWqKIN6LXKsWMHQpvi0ctc7VpmAwt1YQq/wrSH+/rUFE5ttDG3B
MV/5eIeDhYzZNOxCjDFU6sRkXiUZHwcj7o08Z5lV17nhhvVJ9RTEjIUtDovCM11s
RkINR/9PU8P/jqchnENzB6UtYzHNeXPPVzgWXznJE3SwPmELZdHzVCZ/bHlFCkX8
YcZ04XRNo4oxJh+RBhwcJNOzi6mIGNCy5+7D/B14JulWeJbteMFNrFlySjk4iHc3
0jCT/5byGPygzOPRbVIEjhHHWNLMSXHwfpfLdKw40Zs1KwOkS/3c1pjjDJcGiXEx
rwlplVmyEIeTSBitxMHnW+z+Fdl2jakUrF7DxAf7u+11/nDIIfzxYqJV3iSyDBO0
92p3949Zo83qRGYbhNDG1p8ptSKuUJ6eJqEqzgJ/xziO3Un4HzAZ6V1I1pjCiuAw
DXmSi200ayMkclMBJ5fQRKJ2fsVaquLzKTfw/ovjG+azdkMWZKV61AvS4HeNAu2B
cINFlFVKqvaDMRVHysPp+p68y/jvLwUayj3Pe47vJToUznknZnSpypoahXTi8Bj8
5fvZC7M9AGP6DWlAcb8+YiimYhifuXkwSEExf1PSgRQt/iSai3jU4ys8GIg9uLdF
DzS7OGNy1QrvbhxvYcWHDiehbsVpi2wk3jBVSG2moMdpW2b+FSFOVZPJ/0XivJzs
xa1r8s52/BR87bugSgA/wuCBnXuF91jU/ujexxojJbNh5G0ABsZlSXbK1q42TsJv
9btTzuCkfNn82RHBOLWxhPeX8tiQ5pJE7Z7Y1UpozSvw9uIGX+xtqxo7dDMC2j8S
9QHdvwlgQfhbXnNzceSbySu4897WY6JkNA2cDg7B6U1VP19XYZLIXkCn+2yy6N18
MmGU3A5p0TB50tAiSkQsG80wrd3hFXuA1EcFpqYa9zddAhpJwjPei7x3N5vri/u4
pMZ//6zEqqtScuoTG85xHoVBQQ5JfpmewoDGB4/v9ipICcTs4SpBmmsfYNnt5stx
61kFjB9ODkgjgSosRxiVuoGsc1ppGqA4zvA2xrj8225qhIfwTIEpBed757Vmc2Vp
+bD+Tc607bhCNcKpoR8TbEYgF9mxRyY1EUADkK/unN9skV+6Et+uFukEWw3zBRkc
h8eil3X1QPJywl/AJiVq2xj9WA7MkBTneZs1GdpN5s8tqGeLNxjnfE6jq9DldgLP
7Fb/b3GPkI9OfzZ47B+q1Oj4F2hRjhZ8ffhGhzl0MtXVbum63W3t6T9AOH9qxJsa
kkgqFNH29bhqv733ImM/zDxX6lmbFsN2bk2vR9CHDdkKmaMBKrS1q/hbg29o5+sK
HWIAjaxI2Z3mk+hjGz+U3AU5vqpOoBvozVoAZ1GOM4I5DZn4/NupTP8jy7JHh/Ll
9agPamWItylV596qU5ECScPGorT63V7FdNgZ5jVPMKO8A5Mb3g5T/9PM5JkNcNKy
zzSFg95ID+d4vz2QA0nezPmB9zhC0C9DFZTDrqxEnHW8SI9UHAo0fg7UUQ0iwa5m
bwHD2JSxlnZ+6bQI8w1xkJxXOWZBBpvzLl92gkNKidLo8xlZy7odH/MRAWviDjyJ
WF115HaH9HV+9eumPApk/2Ysp+MR7w4PuiqCLWzHQOlOXQAhlpURJlh90Q19Iayl
omwyONwLm1G93PrDYd7J3Oog6RkOvusCZkjYFHJf5qS4V913oSczdyHYSARGotJ2
6drwft/nA1gYEL0+YI13v/F+u4qSnb9rAqcH085fd2f3VjIDpi5ESDsOcX+OuV2E
QZSHDY2dMvhB+sCyuiuQubOU5M/2sqyOYKWne7zNAPsrk5enUEvDZcN2Fv2Mp+bp
GrKjUCc8piBwmhmsR6JTOmNuj5R2APpbA40s6o3HYtHpvpVHdt3DCdRPzdpXDCiK
SimkgPc9GQu4bXvgopGcWtq8JJugZkPAjS1OriMPbb3okaXU+c+xXc3TO/xagWOP
9Ga1ENlwtl6lPjTtZjricdoPiSS4rGnbC30DAY6yQwsv3ZkN+H17P86vfbDK/CoC
DEWOLCP2jRvxZutDWk34WMqzdFRDp4PTCCsTsW0+6vTLFYx+O0T75G740MmHmZOo
WPW3GAz5DTDxKMN9Djafv9hJce4vHl0LTSiHtt3AXhzmL6wk4WtsucdlWP69suo9
qMeVPx0XP1FvJhEs5OmMVRd6OVL9Nt3OVeBeJ9aCM6vM58aZqAO0XJoiSVcUlziA
YZ3kzPqxx7GbcwOM43dRGRGWtThSi/YopixSxx0XpH0UecwV2Dcz+XKv8C4yyGud
Hpq+o/y7d1y7MkE2dTM2nVE5U117zdUM8QHxC1qyrV9ufKx7fsiJS37ZGgx2JrHy
0kD4eZKedDgjCGnf185zpdFVAutnUE8v+RjlN6NmGPLVj6hB/wivgDOixqa0Uw4r
0zXJUEp8P/GMBrHG0xkMrmYXg3brG1pV9bBFq2SSSFTEnDA1vqAtG/Zw+BCIqoyX
Mnuojm4IUTcRQ1Rlj83B+YnyPvuw30Fe4jC1TNasV4TAorHrJCh+II/xVxXvCf/U
xMaqLXY9Hwr9jfzz7kGuWLfmQrk8uz8G4pEByNCz6g7W8bHsCzjSzVw0qf6NknEQ
ucHVzvTzbRQDkzsZyN9bk9CFanmAYXvHCQQ9o/S6FEhmx1Ze6GKuR/c0Bm8QiwGv
5BI0BVJiy4OhyvmG19yveQjjZExl2cCKRMtQ/2ytuwQtKj8Xc2+/kuPLKgRBiQDc
OzQnPiQ+s8T4veHVbfPHDimXIsI56MKpHqpyocCUb4I9rRWeuJW9yttWr5NGoJ2+
5d6IPKTGxi0uWrZp3K/Uk8rrTAf2Q3ZLc7XbSmhr109CfPQ90oU+3YNU8AnnWODm
Ce/H4oX1AAGXqX/Mk6h0f48YtQ8ygBc9KqJKAhUGuR5vMbrdDC3pQBEstT9DY9Bz
OQn12LIRpzjZk6ztmJkE1kP9XvQGWfv2WrCJ/L1mBf75MXhmXAb8Yn9pF5fnMwqp
o9GmN2DXDPVEr5siQvT+Es2IMLLb66cX6Eh1Dwv14aJpZkaOLHKVpSLOeDgoS7JZ
CbGX1JWt3ckE7vX8Y+n19MhXDL9OLyTw5DZujTf40vT21q12GlrjRL/SDFM7TdMn
W8e8beXStEWOOSCg05szHronCqnrka+a+yOpnlQV5+mRNgOSh4UWcQmbXT//0y9a
MXRSXIjVQ+3LkvssMbRDZyZU2W6mkPx73Qfu8IBFBMcMhoLbAT6sRAkNPO/msMCC
u7mg9H5tYln6W9DBPONp8SKgXlqCmClvoDrRalx8d3jgvIrc97EbgRZkQ70RHNFi
HZzIoykCAEonA/YQU5LKPXPDbiAjt2oXoAhs9QK/sgxJO35E9ppqOS72i8lvWgR8
QRkxBnVXWAZ0flbkb7CnysSjp75b9wrMmBOQqobuTszZ+fyqVOxXU4RssCRe0lkK
cXN7i2zJMw+dl79t2nseyvNyJjHF/U33iLZUj7EeJX0494Na9PYgg5Lj4oF8Y5rr
V1AZyhKR1OuuB+cxOEt5BGdvxfkOtlVPv5H+pHIiEyHL7WJIeRlSfy0/2+OEuESn
/bhSyHRvGLfCpEEB8kM6rHdAZf+MbBA9fpdbuwlsLlE/azylx0tGz+WaluWC/cDx
YmLfAIHZtq6SiD5CGhGeeM70vcWeNwX6ol+Crm+r2pdaliE0tTMEFrxM/tgoKxaQ
qOVzLmDyhJ9mv/NC07UJ9dQfDN+9zz2zM0ym8QtsEHyQj6jMbsW7+xPedFEZJVSR
hwwF1Yrk5PGavv/HDyGiWHXnpmNikBQXt3hmnEUh7lXDtjebuRXhSjzqF7yH+aG/
7D0vy09Zk6M8S+vVGgPSjUMgTBn6sEvL1lGBvwcXKsoJF/7ZNjwiLXaMApyfRtxe
5dGvMB3ASWnq8uCOjrfJMKArsDpv7yvDwtQIUU6vpclZ8HP4Gx/U0q6bpiuRIK7q
jfSKOus7X2Qt1jWHhSyov0TEEcO+eGFuWR9GOgTt6qc+qzt+YZYNQ65XzpySMzK/
ZNMQ3qt+Pk83Ejt/5SOCMr0rUWCTERflwU24e52SpXR85nUammpzlNFlrAcNUV2P
Ea0vr3wZdDl8az3DzrLU3mxTmmd0AHWiCo3KnpOugLYowEd3nMSAmHKQtpWDDTnl
YFl00huN2KqAKaqWTv8T999eAaY3pZQvam2m32Zqz0/HYRWDtpDFWUfK7crkZfl/
2Wp+EDSlsUKYq5h/N7D80yx+RKdOy0udVDq/BCxM9emNyPjTWkI3WY4zV4jyuGGv
KSzyIvZqCuQacb4yM+pjQvRhqGvB0ntJkUQHWRbP8+1feelReoGCgjWAA5Kw/e/E
ImGap5/A8iXXETUb4mU2iHlKzVPMpZ5QBULFCgx4NmuUDO7CRmwPFSwMAPi9L0Sa
4EC4CqjaG3FSN+6VR5gYqdcZR1M09drd64VkXH6vKUbMXoi/zuPqyj7XvEIBNoF4
lT/GHRuVPU6xeFBMnE4WadG2RQpPXtJ4fOrBe3A/d8hvjjnM6gCMU4PJZ/Xz9EJz
3uCTDj3bFqnCYX60M+bIF1k4hfpvqtBEeAJjX/ygPpIu/eD7WZRm+2IyEEJBgDLz
gOMALpt2n9Soc+3hnbue1Ke6LpD0xS0hkr5pmpv49bqy8UkXQYEXCMX21NFn9fgd
Cm41BvcLVhg03U/aOQqjMUgpNVbKh2xztUSz60UNqWDaoHMX/PROqV/h55wKPL4l
0ut8CSI4J4PGwp/Jx8yFKrTA9deLcOoYPa+OiDxXrOAwkYPE8KRFh7Xt4i9+qw1v
xoo9J8dJ8gvEzGCzrLlQ0J3JN3QDN5/weSfotUmutFxxgu+dsK2tiMR7kAunOw3e
cxFT5IkLZDuEo6QI53rCHzhunWmxo/sXd3xa42IUsWUMv/q3DfAnwjDrjjyWl0vk
3zudCoyhzAPajvaTK7yrTLDWz+e5P4mJio0fC0w7Oq3sENAbz5yaJEsXatuwqXZ4
B6beEMJwEZx4LrO0G+g7mhgjbVe3maaLEkvAf0YeL41mTexAYqCQD9b78B0E/hfL
a055suQ0iR+gmYftRsyJT+OE3hL5Q4ZYWFKyBY+bXdlUNjs0rDcYPX9lwL6v5IL7
LcC04+tdRtTQDCaZE2jfJLxP3k/Y7fwGyFbjzeIMOepW0lSx+Gw0z1K9Jjed8BTh
d8a63mPzxme4HG+kgmpqOxv4s1/jfTjP7l7F9Sk+UWjZFXoEqt3SXX6vw4kc6Z+5
hQfw8Yyknab8jKjAy0d9+K5DigmnsLNAMEzXjwyvCCM8uXbAZDQhs3aeRp+AjfWW
IqHi9XKC+gBL3GoCSqGgtlWo4lSZVEP2LjgbzA/9vmOQn3sDHWyx4XkKZdRXl+NA
jMNsXE+BnXyhtACaE4h9M3Tnak+7yYa1DE9wsqpvb57KB521s4E2v10guR1VMk/E
ZFAWqHedab84qZeziOOAYjMn0CGtfRUgZLzopJ5uiOceTPIMEZH0vyJ+7MZ33NZs
hvv2ZFXVxOCiVA4wbvcORTxTPtCEk13TcocOgD77F2xQFsgAo1XnqHvWPKZ0KcMd
6hL10HGyUi3y+M7xuvvioGmN85MnZSnyMOhhEyZZyvgFe0Rw7vQWPZB9bXTHJbEC
SiZ6nPf93W+VZ4x/aXA1SWyw1t1ih2LyUqNd4s9gLUUx94QDvH0Ax88PxcDnRitu
Hc1tHLD+a+8EiGFE4ltjFEG5cfqNl38QUWeDgmuBl7fMcdK2igjlxzLaV+wSiFF8
moZ6A/wpfX2otxtK/XnRKzg/pIQlZJiFZ0nCiv9EjtUi5fiLRRh3tl4Cq4WlCLdL
sExJPWqELs46hZNGSH459+ebLvmuOqIf73Ct1pdrZnA1JJkoFRoeaVWDWFMHAAjV
exwi1RH7J2LHeveHaU3Cn557clZ7atl/5OfSjcyIJ8hh/MGQAX02PxLva3PE+Gnn
w/sn4izam8v1HeC207e7L7Fo4vZ5oChtYlSROgWsTC/z8o7tWItcTobib2Pj4tQS
CHu3mGH5ofPjAq93bwQDDJUqc6gSSgnsZH8TLTEJ94NpoYdVdJ3yX/Bw39dCRydL
E1pDQXf1qZzmautUJIh+h04kNqpALsGp1sGr9fzZOuv8l3LtcJQc+i6GpHJivzTJ
PlIKbqzx5SDbVcZH8H5FfY5Q57Q5kolBGmug9dqohSUW3QuARunjve6+uz3nGYLd
8Zm+0lHdUPufkOK+dkJjP/3IFX+O5j+9IlXjKSFOBmK2+EFfgIq+00eqR2IpvHm/
L+0VAlgXuMe3PLVr6FFYlDFM9hQrqD+AdDJOQT56as5CyPeE7IwWBWMVQnAxUJhO
lCL+WKl/h4TbxzNUJm+XjhBiF+StFOVDdPmKvHUX+KK4TLeSD/SaBW0Jl5lnXv+T
LvNPSJw17oQAi9iSWKRRIjbC16cLrQREYWHVs2tP8PhgVpBFNeViDjI7Ob8vrtG7
1rDR7AqwqDwa7TydT3JarqwBfTzYxhmelPa72LmtaUman4PMTB3b+iYyftc2sgSX
P6w+6ekz5qin3jng//+2eGuxh7pGlYMzMv0aC8k2/8wMTbtn+SteXHqSxmEluR3E
PR7eeDALAYZQg7M+JePG3i6+2xsO2dZYGHXkQc+Z5PjBor1urbM02QirATJxfBb1
qpPOfCcIPO2EQCxr/IFGM+jDX8KnAEceREgmRAXrNhjtAP/6wnb/4JUbd9OtTpVy
qVqInf9q3jyM+gxjNeRuViA3OPvgsokayWHrpyMydz/odv3eh3HqQ+lVOnduLj3p
BokiJjk0QiUBXc0h97MZU8+hfR/mSnt4+aGnO2mbbiWnPX0RY6uY2NzYK6xO0ALA
oMNOUQ+1JP+9YMFPaJx5CX9P5iSs22NtWPMNpvXCPfMiVpe+oEWBF0KvarHAn2vB
UmL86kqh1Rr7P5SZD8F9yMs0DXTT0Gd35rkHUxr0pZ8t9Of4XMrjG5rTEBQnpkph
XGJYDXY3dWz6NpfSQoasn4jwAa0J0tTJ1P0P2q73qLu0qC1m5syYImk9ztUOSuCb
UuxWTGEpJwxmDGE+7hbWqqySmY+nKCCMg4T1IOVMIKlW0AXn8KqU6+O4glvBU9/0
F5EqWXQCLaSJ6paHgdGkACkZga6upB3c2xl8SYETT+hOXRjhI9qiFZDFwlBmTz3B
CHwkNeNfwrCFIs1GS4QeZgprTTnplsCXfrzqktpow3bdrGt0XwbghWQev+t6XdwB
iYcvVlUdjPUlECQqGQmzuiNuFt8zC6dm7bMWJ1kfWkPD3tFNxIO5AKp/u3/81GU6
Wm/5lGmG82M5QHOkgWgx2+MPh7/elic0qe8YXns9IGfMFtaQII4xOzVTg2pzO9gL
/ekldBqSfV+TvLeXH0z/CBHEuS7TS2eUw8K8eju/VC3ngmvP9VSoMVVYZEdVPlXD
zcDvRYfmGQ/gSHCY+5nuiijCpBhXkQEP8mlnDdHlEVzw5+OPU/DVyRBbswk1eu8O
aH9D6qxdFzU/8HDP9cgGBdF6X9RwXWU1SjGwDQq5x23tJAv1j1LrOHn5XhQc/KO+
FD8nYyAEF3zfMU+X9oVlc++84w6NBFCIxhCIwpL9ntIj+BkYXAT+zH1CX4oLTw8w
GpUvZxOFCi9CWOABJIO847p6am+M9Wo73OZMNzSRYVdIzhcfuJnAUoG7fXe7H2vk
Jh02xSn0iCxxZqIHUP2VeURPXFj/Yi3Cm8RVzXzfhe/WpOcgwrCe+ae6kBAegA8V
YxBbS3GM0a97ac4s1mCucLAjxlo6EXLv50xsWMHBc+qJUy02vV2XheDPtlq5NmIn
R3W56fvjIP1y8vyeZrNnVOEA8I8IKOQMln6rVM1NmLSF06MLUkfahuSXh/1Ym228
ZFha27lSu/xeDN8Zph/DcXbJWfX4Jm7Afwm0/kJHA2OMJaIa7I5QIbIkTahVZxBT
spEgbPaCDhFO7k6B0eomSgZ463NoXs+tP5aiq+TXwynA8zkMQkb6V/ZhJkRDOfNG
iEA5Mx7uTHE6RbwIKpYXMPt7eNiOr6J9BYIQ16J/Pfg16LQz4j7bUpPPYtG9uYmq
TLJEAIL2sMvbWuR16/OvaN9L/V2ajxv8MpugisDHcgizLc7S6lppfMUEQR1xfvHJ
IQBOgOCA6p+toDYnqFoiZv4Nx6LVSncwFT2yN8EdcZuCyPkGylQ5gpZqAxlT49ER
CPm1iZnFs7ZYwtOqU87cuO3xrSnRXRV1LEsCBLM5utgPghI/FWPYRV7ZYh4Dbih/
geOKEMEy7fMkTZrZdGc2QH7oxNOYGZZb/Yb8fm0zlBuL1zxVwPgWJx3SENqtm186
ePnX3ToS/LLg56URD6e74m+DqiAOL6XV9HNSmhlRrRvXFGpBeukNsGkRzafcsztp
tGoTMR2vFv7jdDRFezl0jElbC/xauzRTJ/nN1dD/il8vX1GArC9UMRBhc/0XG5NA
fnnpKgREQadWNXoflms3nN1QrB0zSShDbullJGERtF84WTAAcE9hYTuKb6zE+vN4
ee/CEz7+kp7JybqZmG3JDApGY7KBm4xaQ3c3FxTPlwW1Rh5zJhor8tJQKKGRURem
8pLwxINCT010cesLCBHb7Nc6XdEc7iFOUwdUI07VZTUrYG7r3jaBV8eHUXB4Epd2
WrS99nZ7xoTwPom4DwoBdQCnmFGHWVzcdCW5ipu058RKzUSqT4o3K+wEGzknhI5J
liAtjOGd6E5xYx5a20vxNHNBrcjVOBYD0f7z2boi1z8bNaQBXcgGixq8BQ/TEIQq
6fhhu63kh6z2qe2ZClBJEWf9xt17+vQSYuH2xjChpMG7Xl0XvdN9BNdRWPv8Pg1r
6gTqg7cv75mtEQOQDp67/z73vQ8jOvaZ7DZtIH5hxoqboL0tIQbeMrZd0TOMucEs
VoamSALaXdAwvCDlP+gIXy1GGS5N2KTspFoOJc6smLGYK++mKxL9Uq95VwBhCcCk
kgXd8Vx+W6qptI6FdIQNMTTFFddHpFnadw9prJEBcqCz+HkA3/Eb9KYEmM7w7ORu
WofUKySKOvfRBgxhPibv7MVAh0WUva5C1U27kHxJyyRbED7ctGMcd2e/chl26D22
kIpkNM18x14daEB+QSOHfDK8G9R44xSve5PoOGaArTuOPXCD7Wpz2Of3bl4SbVUc
AsYZC7iFMdKKzah2UzDcYGEjr7N+8oY8C4c/Bbicpn5Dl5ymhHrRi0FPhbUSpFfL
oDybtKXdpN7ZsWG/UjJkzUEdUkgcVN7iyMxdBjgDeUwFaW24ZSEO0fB5Ox++icyu
i9xJcmmF7b/RfzyACqSmsvNgKuq0y4RyrQ9f0eniDvv2jVM4ATPlXWSj3h/azQM/
wyqFwj/e+auRpaqVFY7FxmN+BvTQuLfArmFyRwDMUMhSrtZLGcveqd2kGce3kKxx
fVXJRfeUqLKvzNqiXIh5CWTuoFuXlrCjMq6wWnnzfRA3e3RNv9y8dtLfsc720cxz
UYWjL9uAXmD9GNF5u3EhsAqOvHzupm9SD0rrmwSjZJvSjBeU/GaPNH8bmlt/lE04
lBH76KO2ryv7yIzmE2eRpkVlmW7FVvhRV7stiARdB6UYjCuhmuEeO4pLkm1fTrq9
VfIODvqfzhWpXo6B5W4kzKuqTCqZ8qwLzMa/U056GLH8MEmX0pRPVBPwYZ0pKaDq
/gQwbCI0wtFQUw1secFD+Dnx0007fg8EmVVf0x44G2WnM3V3UaMyjmK/Du2gb2gb
qgLd7SkRfv8yPogWjt2iFHOSdIGwBj72TMLhNGNjfw195pjbB0X5hq9bzUCa2jyg
djj3APhVdfxhrFTP8oN5ew/liQM8iwn9+dK0nkBpzZP5KpZWYwm5huu8BvcwEak/
EXaOvu3WPjX/vCjuq54nr7UeUdrD+y7XfLZppCUO0/ejCATRfOfqsovaloUWQeFN
4WdqxIkBdQqegt68Ql2B5qbdQX7zsvCbOceBZ7tqmflyaSNKB8DbaP4Bsv+WB/6d
rNzmOgtg0DAdrKVrfvsZwIakTSt/ps4f4bvDaQtA4onQ/4dSsU52Ch9fcVacmbaF
VhvZI6qmfgn0mhPby6KF+opULFJA9/Kfogb7ZK7OSPgk/zCaIMLUX/Ol7GeocMBU
oSqhcTehi9ecksfAdpJuW7O0ouPAgNmKEG/V7Cea9AK5ZOAQYRggvbJa5Fy9NfGl
tpDmdyBZW6jkvPtLJ/4jyUGFGGHZmDZN9r73uqrsIhLaf17srgIdSvldy5Vw/biB
uF5FwtkApuBfIUaAIW5A5iXopTNt5Ys9zLnBPz1aEmaK9MrjzHzDcwes+2jhUlOK
uexH8ONNE8Uabg1PisNvOSRjgQJ4IFbf6emBgk5wk28xo5CRMhpghJHD2zUEMQz2
oelHEQqvozlrwUjIy5azX0xWtl17aAjACLAVX4VCEGGFY3mcLgq2FFhfZpn1tyla
xmfV9V8lGijGFaxlZ07NZx85oMqa4c3/7KSc3vHTdHnc9iRSX9gUxe151AfhPBZ4
tQhnzmdVhvfjHR+PTmyLhyN48OFA2ylucLbmDKh168bvS1z9YF0AskRhaVV7ZhcV
P8SZYzHR5FaCqi7eSL0YhyGo6pY8XvO3zlmYW3GMnBAFqtmuZPSWcegzwiCjZJ6L
kqf7CEbeiKZ70sn2+WZkNr6SssPyZe2W02Ojb+kt7zV8A/lLxTIOHv0j4cs79zi6
zGicOBiSqtS3eIfy8sBEEtrVyOJ4ALcLpt8J71Mrxmh+yr7mSf4jw6cjPzuv47oT
eM3L5kxIx4A7Ld9Q1YXbjACqvAv5knD+8Wr6cn0WqPdlF/YieehZCePKYrwhBGGh
zfHEMoTOkgvMVa29nR/6y4RlRsAnqnSKKp1Z10YTZcJD4T7/g1EEHAqmxVnDcmo2
cOoN6B0qOsDAZycLbvmNhtwcVLDxlzcUwLuYkNYSdFQvsxBuwfx2hp8xupyPOPUm
Pxlg14towKrxwpB82SUhAL9Q8/LiTaOQ+59ZMAS1L/33szOAKIyKc1BGlvTU4Pms
yyfslV5t/54+h9BJwS+0FgcxA1TQipEjxWib8/6SD4UxZy4RuUTWxwPm/IOBNO/L
nlfkKKjuiQDk8qYbCnmfe8Xu1cT2jhLvycaow2rZGnd7w8LtJnmNoZmYAcs4CaVg
z/YF9lPxwRK6dDUXfU0VTShJ+XUEDG/45XaRcRO3j9hfSdxjje8qw0YAKts9LXT8
2HPBk7tq70da9LAWmh6FbwktyWhWvwm6BRDkSH3qKOs+DMFvC+8FOPp1WCugZjEQ
Z43QGQGdvSyysZF2jPAnArwEnOdt+GY+Mr0eGt1tFJtNI3mKH+pShxLos/wolEYh
8BypuTeRgQ85P+WtV4JpIM+lWsIArHAadl/1GL6iWgXPKQXc/MSPBBtgFXP/UDDm
utP/ZSA3H5hOUaMmLMKPJlqil0x3MeF+9AqLN+g3d9Oq6eXctLY7VAZ8pkXhkRxd
+fuJxI120J9TkZIn1HbqqQ2P2aUgdnI0np+Fo0J/1kcBhhigSd/MvkTibPto8nHX
4su0gt8fdKaMZ4Q9RqzZ2iUTMrwcE5vzpw2FmC13CQ0pNYJAPMwxhPWzyD/gsiah
VveMY5u3bGHjh5xy+VNFh+YhK54gdyEDZDveSWiZqCvEmEn/M5TV4iRdTgB+AiHr
tC63nI7grH+E+DZz1jV7B1fKWw/3yx1ctLr+46Vzk7+sip6ov75uXPCtVwwpkiml
Sj7SR73Dd5hqVSKq5ZIX3GbkCkPOXuk9FN7JGgpqX0Y9HtURiEWlR6nN6dgXyS4G
eKfrBccOjRb5CE4+xAVI8b2vuHz8NVSCp6dDRXxv7rYbJSOkQAlEn2KF8sOrUPLf
Zj2YdBWznWTcJ4PGlqS2dZoLMY/J2v7ceaTFDVmWMyYjH4163SPkdYksJburE3Ol
4BfLrQ9ImdBtspe/i/B4b3ue0TkV2kJkQpuOG1LHlm5mz3VKR5KAYbJHBbmLI1Qq
Arog5zyVyTTBB2+L1U7LoBVUrhJk5CeIsCck6D0NX1SPKS1ZOpC49GW5F+wM4v5y
Z99ahqtrtsgAPjYaTcWjcCt+YPc0RlgQNUOAhJf+M6Y9hQDM/Bwwvw0Zbv0XD6/G
F4WevMYLs8F/I0ozhggMLRLauYlQG7sWiKHZPY/L8skCEdlfTpx6iFjTo46St4LX
NWT8ijQqYow+JFp/k54+aSHa+9mcJAz3FAkX+JpWOUyZZUd5A/hA5lPqBhJKPZID
KlbmJR71wPvfdlbWvY5j1v/fbAlrNB5T2qrcdp8ku561ExsI2kPokaweTdDu1mVQ
v+zoihPLv2wZedEZUsszBSmcnSu3PW3nNVdpSZhzEDIyeN5q8hiHRvVkrpoJrJpr
weqJd/M8TFZfGCbCiOeUzi6OqKMcKoBo/oa+OBwzYiOXaWWh9Fb9kFZE73cZnJz7
4XJ8wRWTsp9LzPaJVKP/RBe0YIDYsIT07hcbuoQWxsE2MDdqYovTxYMyaVCPLZ1y
UsGmuJlwuaOMT/r3WbeZR9rIw/dhm8EEQFlXUfUHBL6ciqIVlmxhMPDGUh5M3kHP
dMADsPOrPtAvnBXynXVft+YB+DNeA8b07BraSRr+RSnxyqCoSbUM1UfRl0vNMnLd
BIOxmfbd9Y10kaYwpQEVM7KWwtmjGAHuRLBrkMgbpDbCQSS7clIYbd7R7TOZxfZ4
kU71L1tG0RceYS3XIJ/Ofrd36WIfYsY953D3IddExNEQ3K03rOF1OgLYsdZeSxWs
wA5cg9HUrtXv5hOJddV/0hoUTR2a02fFJtz0CwaecfHaWNtr17DRUuIptqio1oGA
P3pemm8LQKvJSdI36IRZS9NtOSMsvwd0YnI0Ls5lQ1MasS5kjT2j/KnVgLd/C6t3
CICsBCDVuacSVEl7LDoBHV5y2Wh6HxSf8oYKd9QQ95qA2su1Sjvg/VV/QeJ6Srhe
C3DYqCZmTDQntT+gTrx9GPKTur+eZIrgup+FOR4t0nWWuglmjWxxGCHS17d/AMst
A5ePP6DYJPUbhCOUC487iv+gupj3c4oU/c7SHUMGdWMsZGRes5hERoapsbLMlzL2
qGJUtDyK7U4tzRrSB8zp9IM8wcWaQB6AmCnuktkcSKSEZfL7ldNFF6nbWSQyEBrP
zejx7e9n3lpWAq4lSmJgURaJ0UNKZrsx+sXXWPrsehrcVdI568JYm/1rTL4ZdsdG
ZUnPYhcTO1jfYksO84m6YPnO6/QZaXNZLc0mjv7VzPNrKmIwOw0mIDfs+l7kSWPK
FXv7tgzKVoDndnIqrsbDvauPzidHVF2FsmcOoed/5dLeXGhD6uEffC8kpFojxYH6
PGIy/3BGT3ywlYpnRDLZ1SYbmxS5HzVMpom+OXj90mLsmzOEhDSlm5CBstts9JjX
u9CJxEwI93dYxPqLNN3gFLXs39jD7vX5El+QDI6DastCCzyLZdZ4iF8SUEMIFDB3
ZarGsVs5WIDbbBQQZtYErQ187LKIFr04yQrDGcXZzG5RlkYQFpCUclQUheH1MDJN
CzheXuN5v5W8PZ5xekJRycJAmU+4/iTMx7/0lFoJGKdNgTHC4mgJPvFn0G9oPWna
FXPVAJ3uZ39UmRJVb5XYViuMLhFSjJXSpJaKZvbboBFs8M33+xvdKFbbfzwxmSua
E82FTHg+8FL5ly0kcq6JH5aq+us1D7KRpWb/WnTyWFmTwq6kAwt0nVf5/3hCRK77
tAiMS14a/bnyBMWu6xb7s/HHMvVfEa+LLcUVgtuUTa9GjVh75VK6KYEOidbcwlF9
Tdz9vUhBSItIgbkZhBXhoNdlNaOunYSfjo5/rSXjB98fuSXJ1o8+aIpjfe7RhBC6
LtQ0q+RPtWvjc4BUB/ZA2nKjOYI4hitKsFW05GdP1REEdIknbypct5aCiWPhk8wz
KVvVL64i+RB9r3IkhM1S5MJXI5TwbvUgehOOcgQGtxjKg1E6fmg5x+C2itiv4pu6
xjbE/IJ0uqhiFRuFsKSRpvduBVugzGgMmFinUOyXkpC2Naeub6tSrB4bUv01M0gd
IcteoSDmg8+61M8hsf8zptCBDWyZd0XalO1QdewO51Mob89PWdJOiaAOGVX3+jVz
8sHbtNErEttO1jnuxeMpwWJIteUpD8/K+XItm2DyhsqZoXwj3OlFHVI+FwsECxyh
uumRtsJVO3DMZ/g221jFr4DbQ8Zs1sGJ9huxMCNDSd+F5KIqFuqxuBdAd93IhWJt
x7IZIZFxfcNdAFN53I+kyTA+Ur7PxYAfazX/hVwWvM3iEKIMVomF0Rvl8AR899Ef
Sy2iN7kr2OYKXjKU9juh22yc+LEvYWzWZMMfZij7xUQrcwOm3bd+8ht10DC4o//B
q6U3PsqGcfMy94XPGy41AlvIHNKR9MtUaikPNSvfwRlE/rcGl1vg9SuRp9xcl2/i
ZOlBl9oo6EvljfUSjI6GGBsowoCm1FPBPsxDZNC6OcMHdn4oiumrpI1QiS+ShBEZ
DhI5dU2mScr+qbjsOHFIsCfxzH0ST1DOxDZW3hsaevzn8pMzvhHpkrZ3Yq5OYK5w
BLXupVjuC+nadWuParehI4FtKlPRV+WVM6aup17lLBg4G5ljMeh7KKxtQ/wa/lRQ
WhMEbldyLTMDQy1y0wAlqnbRZ0WHgFJmEpAgNNAgvV+aeztUSqRSvfaUWFc9nHvP
VoXcT11DSElDk1lDC5TS2jeHlCkDXJlIMlj7X37T7JyCjmqQVvZSvaJqwRx+wA9T
hiLtR5/MHdF16yvJuTr53vIeHg/73dqulAgfGy2SVQs3wRGNSpb4R/Ns9Xlsl161
4mQhCWk3mvJ/9Un05zSCsBJA2HB+ZeseGny5njVDqK9jw/3+zm4/z3VgT28OFLkA
yYjD2iuD93el/htUYEO9vQ24ktp6nBc6JcF8VoV/VQ4CUbbb/ZyiLSQLZd9Is/mG
HWQbGewYYBG+1sGDkCmh7IjiLicNsrH+1OydmtkdMdKzyKeCrTAF+eaUcTb86gzO
xG5Dtc9rmzO34uFDBuXTPENYkRHy13ma10za3M3DAUUHG777eA1T7i71IJzBcYVj
uJufz/vCS2b6kiSm8o40xaPrbBJNOPcdUkjIpyjhYgw3Arpv7DXKS6gS4Ke96yMK
TL8KrOBWiL4ZnFda2Hn0SOpw208t4h7dAkUgaZMls6tdJPdA02dhOtS7+aWCpUb+
XdduB+OqdwvfU2tTIgeVKXrTMGLOWoKETTlajvUwX2HuenzffRgF553qHq4/7i9a
mG9u8jKrE4oXNysVnaI0jbv5kteYV3izn+cj0C7ESid0Gy6SGo0+/VlDa3BmzewT
eR8z9JIOVq9J6QVhKiD4drEScNlSkQncVDgUTiD/9prm9dVk1HW76+JVKARBs8X9
WGxnwmIB16Ixc6yU4Az3IiPsvidOFyUo63pAw5LkPiXJs4C/Z8jTNohk58xqsvzE
eY3Qb2sgqPDH+E57R3IFAr/zGDsut+otbKkZPkZ+wr4l35saGb+08IkYYv6i2r41
rDcTHC5X8Gbit5Nrezluyxo3PCS/aJLWs9ZJ63MB+N8iOZZrd84y/zneZsf1/pkG
c7IZJF/lWP3/0Mh8Tls9m1ipCEXHqSWx5YCwi7/CgEgP/25uFsVBZxNYltfqlb2e
Y8+1/naOU0kIQb9IfyiaeF27LOt8PWv2ZBfdY/a7/7peVKtXGoRfSXlmpvZT2C5B
XRwlKZZy8cJV4zv0xOzGmDwA32lOH7gj0Y3eAcQCz1CiKEtRL4LxsXyZrgJA1WT7
YnM6or/XyzqYoZNIRGCA96B2nHkm7FopKB9C3e6scTkn84Y6WKI/QLaQKyHq7q8W
RXASG4eeMYi2mtQzT5qHkH9xr2W0MRKpFHKeCaLPcKGcEhXWxjVt9J0HZKzMtxfq
VywTRlzyYYi0ueyBLaAfUC1qyXp145Vwxqb0PjVmMmIfqzq1/2S+K7Bbf55Qpgwd
M53dpMQpmMmc8pvWYFU8egFTeTdHN2MsAEBNXuxo6HaPcIIpYzmwZ2NC8vBST9Vz
eRWTL7Xq2S6BM7gedvBgE1agPsictWzZfuHJIkbhU6PHFTtevIr9Ip8Rxqhx74Ts
e2gq582N4yEJe3KUDmNLYq3YJs2vLwwxLGHMyBqYw2sueY5HnUbDKWUWeHQA7B4s
iRojOp/Pyo25WDux6uUS23kntOzxufLofQtFsTECMbNc/DD57qjNx1W/XycC1RR+
JQxlWz7Cx05Qozp3JmfxeDKDOMWmryWIaLmEmphR1JyVEDlyx/UGb3ol6FQs68Gu
MHI88gulq6vBBiZIKsgMUgW3d8z5pkGBPnehky1urrpGgMdFvek1sip4glGFggev
awt2sW/l9tdfE/mQBQZXtDxoyITQVSqjhVPEwTdhv73m5vvjh1BXhMQnLwedozP0
az5KNqgRjjvMW1radM/f5Dg8cQZMF2xyu2BOEE/9aA6n3WjUGA0vNryTNcHLDB3P
5oXOe7BmHwLDGLKajFQ9cCJTi4YafsllTb4T8mDlxLHivY2eTHySRB30uRuXVte/
UNV7sN6HZYcZ8TuO/a40R2xFo3PRCnlwOavVZq+MKElwbFgMTX0D5yn3412FqxWz
paWi3VDlVR1Tx1fOascuaS97cJtVFoK2GCvB2DsdwauerlQ+V8Av4DKxaiYha9lJ
jOnkY6pCIvFgmO4cBp0gc3jLJ6zb+MLD8geLXvUxb0TVg3NX7yXgx7QI9LTiWScy
NqMpm+qdeRSyo/JHJOfix1Du4NW2ggIXJ/JGFnsRztpOX7fNFUADvqu91Z/bYigE
k0r0hF63nfzR9BD20h1g0WkGPybVBOKZFoOsE3eqOKUC7WJAEtYsNT6gRA2Y19Pa
hqB3wcYX+2VesEe4h3rDeudqb/JxsoeW5byX4804xmRTZsOreqt5I1sycrXg5HGq
IlESYnphkROAr/wTybYKJvmkXPJwdZP2d7nOLeAlO1ceevmeeSHJvoMCF+3JItjZ
sKr7ILvrmIjGXf/sgVY6PckTnu/FQ0sTbnt9OWPlO+/Hig2GEenOW26obe5rmhBf
/NEwvr3lEPNrFfrB44PW8rX1J1fulxJMXRYNK6cHNgHN9zsczZ5CclWCqNe8BwEb
gmBgZZFqZYVTFiCqFYGkSHfuLdE524vQZlxAqxvKNN93WZ7dVm7/SrLTgQyTaaOs
wEJFNK6fd87XxrBx35w/bHXjs3FccEoBxrbvoGQgUiHxkMEl7JdMdLLdsB4z40t9
9bJzSs9c/XyeC13BXGz8eUQzblmXCX5DiBCDM0lIsCqiKA1CZ+eugFkWGfNVRBtV
PuXIX288PhvILyNqy0a+eW6q9PXUKvwo9sZIIjgVVEeL8WsKvqjEGRGF8VB1JdNs
fTVkrL5DlFfatiOCNaY3fd6FEB7QBo+PXUM3RuRknKgEsdvUFBmd3AZV3GfO9Uwa
nruwXGN9q3haUvwzk8VsRBPgrC4WzCnWFSkTSGLgzexw3kje/FZLu5qneJwc/0XC
vC6zuXaZKOvPbMohmKqGh2IU/1JgUA1DNaO8i+uVFt+TAU9/urP5x96QolzGR7cU
u6lkKb8x+DKuqKciUTgopYen479V+ouyT834/xm3OidkYx1XDJz2BerXxZscCaHx
1aLHhcCy4RdwOtPv1rAv2P3hiRsWQ9bfH/Fgg2m8w4njt+0XCkZJKbRcK4Dz4YzJ
QaaUomEcSqBUeIdQeoZ7uytB5o9a+gmvlJ3i5hjHngTCuK2wfftTGZmXcnfQQVsq
XZxyLFtas2Ij+1tfpba5XSHksq7SrTdSCpQhopr0NWaFiuwS9lMlVOYcy7nIMUt0
FRw67Zj127Ro4iFIkyXCr+MyIYdlBUNA6T9s9c5crMcJOZ4KhLb2EjF2TZbGFbbS
7MbnTrNfTIWndRm8OeGklIPoMX4z5gc+hU00pME0AOLeE82iw7Fg0a4M834UVzi0
voINUIknhb4ydeN2dZIbErXbJ+jZtUumWKsb/M2atB2Hpx+uLKlalaLbG0VfN2Cu
/5Yakyt6h/Usf+x0vQ1CDwhjpZlXNSZ3zu9IYx36TSCGpTC+ofYNQQy2hE+UG1e8
za4KEzuOcoYIffU4Upi9ijlh0Eb/+7A0YHJjzT/FT4eZ8J2ERPP6pHxsPJ0OtG0R
w7yqw3nNAA8TNU8HllZBwTUudNMHeyra6z0cpjlltt8AOumCITJZx2fev69Fml7U
3eKlYSD5f+kEw5QbeAhXBsgOwe+GyW2EVe0X9qMqey+7eKqtS6nsayeix+VhBbYA
dkeYwQRwCZ/a3R0RcSqxW43JpQRqQGYWauKz7tTkf6Wcg5Bc+iwmAwMPsSjFB9Ss
f4Ur65GmQuplO38X3lJbAYAjt3Jv66nRcsEEY0hX3f5eoxTiv67MpQ0ZU+lsYAgb
ocmW5PJcZcvsfylYjfcjJm60wWc419heT1tnyNvE1ix0nuL1etGKUj9ixIvbGx6x
bD6CcS24qxA2SDfspaVx9isRMgZen3pJi1051Bk1S1ReYBtiL3Kb3LsphCQMK3sj
8hgkcOPEs31CoxXQVk3ZRWLpzQXHs7Ge+R69BS9A/EdQQyKqVUolmxQ0GWFK2Uaj
fEKKQVxp2vp6wQb0/5M1R2nSP+idIl/RpNw6i9tdJzWNlB0/y1FIiac6vFbYbaVG
npS3CugKlguKsiG7Pi0Ajh3Qfkqgm0ShFGZsmJQvApqqgfSaUi9GWXvAHGSkPBy7
MSa6rG2ryzebfOtl3iN7EUdKQTg687URaE8lydBnroa1WN2ZcTSkaiL8IzRakvEG
aDg6b1LyDJJDzL+qNWRucQSneS+Z3UwDmc8BOV1z/3LQutwKMe80odEXWKy5Jyxs
lirWpwDC9I7WwgXMxt7Byp9d971V4ZukyBa9qG0zUFCnEZUu1ln9IUOtRSgGfFz8
Sq5qidNyQs6hvTXz0PbTyWJ1RhTK35byIYHVMeg2gFMALlD21G+6miFCdjmWmlAM
NHUcZxqapu+PnX5r+jlVHI8aHN5LxB+Hxr+IR2QcHLt50aqYvvBZ8uiy960IgF7b
5jsEpfZ+d8QpZpzzljYXLVoWL75cyix6JKsyiO9N0UCltn9QCFPSfESEO/zTzPET
ee5VeK2ZM5KMIhjB8qXn/xzo50nze7uw7Agobpc09N1cY4xIdsEEA6M48Mhxg7iX
rcG7YD2uLmLaZJ9U7tsW4qkDoQnTR7Z2qphp32hJXKkvoR69+T1QxotTgRxr88Wd
ldd/Dvu26SWqGXYnqkx2KVjpjma6+DRlLbtopgGk88rjMz8jFU/k8iVgS+RH4mjt
WCKsMX0HVOspOayeYXMSB7jE1B+WqIIIgiiHjaYaSdku37yHtIzZfEhOHkZUGlMt
Za/9iBBPqGfCmMWzYUFZHfy9HCGE92nRpSuQ/cJvvZwl2KOhX11je828M3nyFVjs
m51Y/N/b31LrNQEnE7ntRXloIcCf2XqKobYG3ifnxblrEVY2H3Pe6e+WAmLg3+Hx
3LfPYpf0TuFTQnWpgf/9AnzSuXsR9MokryoWgolmh31lBHaGYFpZtgq/Eqf1huCD
Jo8DyXk/vFINqqpQvBaoOtnknsOW6AQu90VAxCxSTXzhLgofCEwXXHhyPG/f4HSZ
8lOIqQ7AJmoSAJKeiu/GyMycEInRA7vBZQOzoYohLtU3rFgBy9bGa+CW4yvykRAy
+JD7owi5iEecqf3UJGNtTNsVICD2sfpXeyZh0e+ymk8H5pusICuCR9VLMXb04i6H
hgU3lDhvKMf4Nk9cwIKQeCpwmt9F4UNxfzPH1kH2o/MVT6J/MHuQp7qHis7Q1rsf
PdbLVtCPx3TBHaRpggrT/w7QaRQ+utkRS24Yz1phDJ4tP/SBPRQcSETF4whZQ8s4
dqWH70paPKSRBlsgBdF7TensPRryg25Cd/qPEBoFp7yIqTEbxY3a+vnEQW6amwmn
EnWOe5GdjpP8Gj1Uo1UQwgSSFuXwrZP7rUvOhxt3lnBbJToTsuig1o0nhwSD8HPe
fRTJG7cqYThM7kX7MwFZbzF59qWx2iNk3a/wy+W4eWAwGZ5NXWxkAhUlg/y9lF43
mwOW0dOTkY4oi2L8Qin/6aPiWewuiJ1wznFBot8NfJcEBfva5apEbxYfhP9XUobL
3G3NbzBgexu3jSt/IEuFt9g1y745J415ZBTpElXR+ArLip0+AaZwUNPDBTZrRpt3
yTkGq8cLh1T4fvX44Obm1sfILezY8CFtfZYIL29LmsPRYhZOAnYN9wsuvJPEsKC3
XxlVZVKdnUB8E/WPxCsDuX1tqf19H0YC1GknrSDIibk9fpD84jfdQ0V/bCi6V2mk
HTWPLETuwmhpaPc6zv6gFjvcbG7c1Bs6hMgkdj0zTSUtlcJG5gH/MeuIRJN0gsso
nRRdQWFDT+BxctoZrNo6NJS/WDtat9Ouqe+59jGbBIkk8yy+VjZjVC/SI8fKoFsg
0dbvVpjT8Wvc8WAebI3/IrPPUsvWO7XuTL08V4Cuhy67gjgliyCVuca710LTCPv0
SqCUCJeY+mux7WidZA2NXkn5bTfmBplXvH06cqOFiRe7sfu/Xmlh+iy6AWUXJnG/
77wMTvyfqgKzWART3tAWg2rS8j79QuJhxgRzfk58uUGhfFFCLOJsP0LVoFoO/3Vb
82f6vOxC6hAlmFGPHoNmg9W1NHE8mx2lvnrpMPQ+UFNC0gbt8kjeHiLgReNVW7Vw
Eb15Amxf9dAPUpW4cHJxxq7wh5aBAw6uK902YEfU5L591m5K4HfvPMxdu7cy9xvq
n4lyEt5oVJemlb59CaBCjkzCxm2oMEh3ChvASvrFC417Hrt475yb7My25eXkjA8w
2/e2pA01AaE+LpNd/25ZOuWGnl1E+UgmaH1DtdpOlzdBVfdFODviBQ6egVzasBpG
9wbsOK7h/kPI4fSBaPIl3Pv4V6F2b7fzypr4QMilEntM6rKtOpxJfchawJdgpvts
eRBxQBGimYiLYQmajNW6teBKbjdqSCtgn0wPsClkn/+ysLRvW5XloaNCkC5jD/ya
0Jikkhv1v3Sg18S/ifMvuoNF0dJQSiKrxPV5hsjwcbFSOwRHN8fslBydjep2Dcyx
6im2K/w+MY78Ld5/vtmN4mLF7Mns1/AB66VagbGr8i/EphKJ3RT8EIch6JKZPPtY
1UzA/qjhAIRWDY1fWIY/3ebh/zPDrmHCOZTjqa4lCRvxWPnJ3MmaDUqnQaIq3a+M
MqcNVoXnEHrH0FFwEVuByyh136wE8MB97LRqHOEfAOS+iANwHBuhCY5Ltp3Go565
6OyKEwT78RDodtxNEYNTqpGuGztqQO6gcLXWOJjde0aSJ+DvTiFNj7v3TDtn0cR/
Lzs8u4LYQ3QQ/pn32hs/5iOYarBgjIGSD2NYtQYywHxvujCs4Jr1Dx8LRxg/X0m4
RMLWXirItzfOA4Fv4nxUpkaxi309GAXypEXpZpNQNWobhjDIkg2Q/HDWuumGdZvo
yK7q4upnKXgYmHseZSOtsU19cRoX4bn3UN5baEyl2aU8PhsuAMBKLzkEO1auJrT9
VXpl5jFrziIrewJa4WpFMlpm4GzGst/9n4qVmUEnGtx7WNWcgl255OVapqeUXCsQ
wCuw0yfdmaJQPo+cUN9eKCnIqTJqMpiZI2YzBbqZsFWfuQnIvoFtnx/fI599AETN
r8h4LCmjWxDNFTdcO4Ycb9978dBNbtVgj+A4ykjzohru/vpwJIxUrybTiFPFnp0k
PH2O+pUgS20MnALFKVLtZmxzKIyCgLLaksmPIYiFl1wUD9J1iIu2Pj9k/HMlddzH
A7pyCAoMEJFfVeSURsRMsjetOR4NCYIYbtkA1PysoE1dSp9+aeyeBGWwd+mq9n7J
1jD7NT+p0POX6/3QnmUoIi6wOzUjkL7vcGTTuSIADSe0cG/OCKvTbM7SXjLf+M/E
womahfnOAGpNxd236vr6cQUVZa2El5oxyDCZec5dHZDGoUQSZK+jVTOsoLZf9BI5
JyTi4v3UzN6zmHPIwiSG1niONmZK9Cf7f2hFm432o9E4yR6zUnNx4K1zF9K7SDYr
yErr8lW10EspFjqAaasqCe9SbK6e9hAeb7l3B5y3FL+tElVgdQuYCxxDlj8It72T
oTK7uDk5Zmxrncg+IGP5lRJQRoFSWd+woJvwaNSQRcu6+uPVHfoej2yFO/EANT0o
ddIWWnOEs2OFD5r141uGDQhSFwTZ4Hrm3D4F8RX5H4ioXp0Wpbw4jT7ySXUIyZR7
ZPY6GBH8l+5V9Hzj15ZBlFNvGskfgqeIQ/VHaAtOlrARMe3lFOIL1HCY2xDK9IFC
oVaIKGQwpfFiuD6QVGCRISClWhqH9+I81+LXhS/06lNTWe8ijJxeYU9MGuTUBjdB
KS5rzcefnAteGSFENRHFooMul2aOtDllJ6SXM8d2a4NoQg6p161RJeIL8q+dDEzr
eQp8o+gJp83MMbsdRY1caQginLQqb+XFNDFHNRMo4q+/uKc4Kj6jOriaY5NgJg1V
3fg/BlWqFAiuOvm8u/LarKp4YDLgTp1+hziEtawz5kXsFk0XwXIKYYVLmF49ykRo
rBNyeBV9H4tWqPMdvFcLh9W8sJQTFB/VAjSn2rWFj2avQMRK8mM+KYoamCHOqwOk
S6K/bBGxX+38xPI2joYij5EF8R/PJnqTUBJR3t4sImExczewGA/b626eCrpLSg+Q
h7PUBp8dRgjNyNQPgtMbHPymSHK+T8s4ZzLN7FmX+eq1L2nD1BWAmaMiosdydUxo
RMr36ea6cEB6NpfhIifnAiO+0QgTbiR4hC3/Tgqrc7Es6bVwFmzmIPX4dkCLNEG/
mlCMyJVlUX6WV1qtEj10jKMm4ss8c8VsIHiSwOaUvEsz+qvmMi3+x9NV7BHDKOHq
iKoaGgrkhAlkuO3MM6XZY+SkhjaoYmq1HrfOscLXiPRC2WKo7VNlSxTnOSU+nOOR
StSrosQ+rJYMpjBRB7bwMQ9eSAKjOqJ9EeLqSnxPysBzIR48478iAb4AvGPEdssE
g95IXgb7RCtm04FoT7QpZ01lD/s2Fs4EiG5tSFkPb41i8hs5OuqrcUhL0l3CSsfR
Al6bgq7GMaOAGY4UOCtKgSEPdfQ9ft2RXrWbhGa7QBqlf2NMUmBmhUrK0V3G/r/Q
OUl/OW7rvPgsCuJMHP79YCAo0C4k29YC02T5iAXLTvwreJo3rK6XiMvNijQdju4A
ARE/IpQ6Slz+BhfGYA1dM/T68u6ce4o5diTaW8yvP1VuX5dW8+sA+5wdRGx3u20q
3UekceLSx6SGfz2OjRl7cPoNc9c+bHX/hx1adfPoTjUqMDYI2hE8WtAhlxJ4GAjt
wva3LXnHq9oANMSn4VvQKnyyKhBcHUAKQW7or2WXpZwYwd2QP4qJknNPcuE7R6WJ
Ovan+uzhYq6eh7oM7vncbYDsblBhLI8YnMg4odeK0pXoDk6urZxkDoLXULpBvcSz
M1nqvcpCm8G+BikrmSvMvFo2AlxPS2hJwfHTWc8x/bEBFYYiZwJjyQ9SMWIYv0qx
UnrajThjrlPVE9QmAmOpQfZjiUQncG25Z7qoYvW1GN8nd7O6AR/HJOjYX/9eDXXx
GzYNls2WhezPtgm/h0lrZR7GP6FIX20MxlpuIjyFJUmTS+9ln/QkXmXqUt+iONvD
WlMMzk1A1YCCQMRI4ZMZPdYKmqGr2kFeoNxLadPBxdSbBrGaLZcMNUB/uKeZ7HvV
gjeRJ5QzyAd/txPpNCwNtM/jA8NencsbHUJ8C4NsAAabpNcBsAWymmV0vdLcHjOf
bQi78bhLx2YGlQstwaJU7K0oChRMHAPpAtuSvQgdVM47DcIjEWB71vM+y4nRXrKs
68gJUTgPbKV/8sZVZ0ieVNQrqoLSuig1yNapvYI8IAGeILQ6hIGWXX+U2Jba6CNk
Cd6hKgSm5BqO6R9QVk5A2Wa5PDhC5j9dgo/q784nG5FvUzE1BBF+s3beHGBC87eG
fLn/402O8VovYTxcous8Uzlb6/YgbdwyJStUl1V7XY/n7+JHpGvCtD9wKoNQlCX6
9vI1TbDccJgdLYTbYyaz41yMArpuKOu1KO5dvpc8lghi0Zw+t0BQGAkQBQ2ozuLX
G00yadAbdIa7HiA4tzeRUdCTy6/Z8mPOKED57GCBEjTRmLkY2xXHzFz3r5dTP8P0
5QhNOlmoa3TZ9z8NxMmFWpwVee0AP4u/KH9jxIU/5oLFDYbO2NOrSGMlT9rd3d/d
A6A6A/h4/iA7GlfLAzJcKC56jYnD4SxsiJPjrn97LcG6rlIV74/+8gtYJmR3R4v1
AoRFkN5E6iPw+iJPh/ZhCcqM7Q8pE4+kBgbnAQa35NytIA5U+U/scg5uSBeci4qx
3IjsELj/xCrUkFnwhCkCj5owHZF3WaEnDGGJV6UPM7JHWMD96DSVjBFvbvwu6y6E
D7ipAW4oUY4XRaE1f3KTlN8PEf4bcV+Ng0qEZJ/PdfkC2uz/9lwdHLMGGUvo9J1s
K/gkEuqwnFSUdw9ORyQ1dngNNJ+cGRE6SW29Q5Vo9F1E+DpQBhwgcaAldtVVl0yp
YbPEplWk22qs9c4LVJNCRIVLiVQtr9zzzMF+/VpVTVSZzj3jlFC8+SOwKm2ZkU4k
StcntLXDMlApJTAvS5gqTMLdT1LBx8SIlLAyfdyFeX6rqN/KUHNbfBqHiJwJ2Arv
cyNF236ri9AF1p1+Aru1mUXh3ldH5kBtMi+t2vT6buFQnsDgUjzy+xw2TsbH4rPJ
AxUVZJ/gBYLwv9y0TfNcJT83qydFM/QiAsNl1YhIkjUSRPG7/ypYkywcLHBf96l1
SFWrEiYgZAXH6BJHifTuMw9S1HLG6ExVw+CaygMgNyIq7hRVG+a+yFNvOfqM/VP2
sbDGhxmkCpdwbbQ1wuvebu8Z3yeHLzSylTNEzMGlr3x8IF0SDdIR6Sy/EeQWv7HL
yPzgwqRYOGMHqesO1k0I3G4rRCI5uryEsNWXZffNKlxyI3CDLrK6VxB+YLyxIgbP
nsPCdI7DG/hwKERgI9NOkgMaunJeAxdU5e3odZv9TtC4auaJX7UIQ+D8GZ9Z28k5
WF1vlXv1GC1v3+ZD9oouEvHS94p9kVosT/6hq+AYpI7r91eX9lYnOUBNXTVUpmt6
HyAg0z4ybK7zoZlojstqxcCYpO7pALELIM4lIQlM33DNB1kUQBQUbY4D3Z2enwzb
TjmkQusnno1C1hGj4GKDJqjsmbuKU4S3bD1usWETzZVMuXcOLJmowlz8qiLI2pDT
EfyNOB4UG46egoylFHBmvzH7qSrs1HzvNLlbdpufwizjf0la5hh4LV/Xxo8HmTa1
orj/BLmaEsaX+IAdoZyYZ4XOZ8tH8/rgkE152cBn16yTfp3L8ut0HdoHQVwXit0+
cbMjGxZvwoaG+d6tk5OvrS266A+WvuKEoqMcx/wTl0WJWubyrwNy/3hcHZZUIX04
Gjr6hxpUYI/zXLTG7psbY7wLgEyfdcmEpIWIN9EabNn2Tio/vmGUl01vlCFTRi86
ogV7krMsfY9qMVExEkE1wxRTi2qmurOQlra3jQ+8E4Mb2MNmqEMexT0/vAT0u8Xb
6Gj8fm/vJVw25RgS1dLOfx9PqwYOmAKm9RQzeTEfqQ+F6aVoMqi9alrDZO95PlwT
+4JVfAZeAV7Ly9QUkJpIy1oyeWpPZi/RUI7p991jFBUNCH1X4zx+pwD9F4/OFm6n
+/15byBl3MkPbE0OCK5S/j4dd1wqGXlEPmIT4l+Zg0lNhC+EJ9jPXl8IqiI8MKxV
1qSY0VeEm9Lw88o6j89Zhzaypa8HomW6iFYAgKypoqcOHXLSDkigFZPkabyeWo/Q
QQeCghAxBufF9JQtQI9ydDtdAOgBf9MmjOzn/4a08hplkteUbOOXhcYdxYvzIe3w
p64pp+6/Rw5t/6rKAmc4GZciFR5vChuJXKTEz5h1EkMUkCJIFdL0tAC9yFdb7Ma3
6dzAEPSu6Gc6LHlg09UwtDMDqcfpsolbRb9ml/hXhHCN/1e19JPZ9tR3oQHzCj3v
kqeo6oubp+WvyPZc7H+kdD9AzU4ZVJv6z9lYtQLAO5RcdS438h88IAbcyYojbNsE
8O1kZHFFm88zpItCfiiyDdDr+uIyTYcVKM2EWwMh9q3m6jjFHpP3HWcGmnQqJbML
BdrV+2Pm5LUWg/cz3tgebhptFCURPNi2rEuVE+oP8V2SQ5nALuxX5GrNOsGYPEex
hYIxvd4ctA9sXpRvjtWLwXN3ouCxIbT7AcSYtGHjAWuoWtWCBnooxhQfmjtw9K8B
hiX6fRnq/N+dBdthhoU9ITwgrdbft7cIIU3l3fZZbLqJRmK+dfXIZjqtDSobyNYi
PTJ9LI6MbQH0BvbIyoB/n5OIzZUJIDf1CJB5UQ+43GrZc43tj/kxGsiDotSO3RKG
Wg6zuZakBUbhoXaR195Degl3LpSW5QITL1KHSD3mbamnMbW+mtNBF8OhzNcRI0Uq
bvV+GOPBUU2vUJ4foz6HnTJLEWayyGSPj0BrSngbidKhrVLEziJul06dxi8AVWlq
ciw0RN7HJUEhVvPHRo3QVrwJwDf4hARoXR9lO0SMLPGuThHEGnVglYRtO84r+1kD
5y5Cmh3Eqylm9uTgamM9YB0A7Tgq2iBl4Db3ExZ5Tqw6Ta85Y1Pn1t65dMgHA2ER
RzEafAMQ5gfpY8ZC1koBLR0eOSIMIu1lc1OJg81zkIxOSTWrDAwAdNMAdu5wWIYH
cp+C8xlZZq0lBhDiF/rakd8Db/nGx4kMwkta0Z+AgW2Yiw6GqXC164rJIpCypIrl
ar8XP4I44a3C5bop0QP/IuIl5H+IvzM1McQZ+j8L9pOGoyqdc1wyjUXIb7QAbPDz
AWiCNi0EnIHSkkiB5SmamCxNodDYAkfW6kvRaguJApM/sZ3yV25wZFDnk/N/rtww
G0X8728weqxL+LW4jk8eJONmUw7XtJfVG30YmAhDE+3keulvit7FFwhzDqRyA0FY
gu4j2cC3oUreiAHlqcra4ocLQamZCkDv1Nj0A4QejRw7pGYFLGsmk6EKbAbWLT7G
GIe06QWZtAOww78qJcnkRVaj0C5SIrLLDPea+5HcjI1/GufHsP54izGJj7Ocb2L/
Hx3eWOdvxejFzcvPtSXHf8D/ZZJXr/pazB78e5QENce0ioj8pcQIC36TfdlR1X7d
hPRiKjcyyKV2uBjPEeGT9TtZX3xOoPdEi58csCCON/aXPmB7gmNkwzO6qIgt/I5C
WdATRTY5Uxdce8Ar4BpmG3djQxJ5s/ty9v1isONLpKoKZRiJu3Nj0Pd6DL0LsTzB
qkh9xccUbpZVoaXAX7T2WR2MfGlDJ9aBvV8UBDqzaTEHIkIXpE5RQUHBceFjNaGA
SwlORnCHa/K7s8M085buQy8yxUuccfy6pAB1SYLNMQUyXcexljbWtbPdlLDzgDpk
qlIPS5B7tJSxT0B8qvpWR4l5EnrIDgHxNkSvDDCDPPCvYGGSTD785785uLS4952t
cqL+zaCtJQalBiSMZgWyCHYBXn2Uy9fOU8nK/6LzWaz/qDyF9jNTem/BLS6A2Hj6
LCXwAiGWFlLzknO5UsCtJ/FAAJ/6c5LhFd/vvtk7zeM/jceTvRi66Vqmd5q+cz1p
QQtvE0gEZdeIbURUdudz5XS/Y6loVuownjJ/59G5drdfqVIvS8oWV7TUJuQDx+z2
Rth9EwS745w1ieAjyqUxSQySA4KtgAXj+RkBL/mKcj5mgtmd/OUVMGfCRbhkC6vl
0urBova0jdexR5p7mFhNTQJWyivaDgXJ4BOlGqQ+pfobULxoplAte1yjvPdFVK64
HqIJn4vd5DmN8T4BtKqTo+7cM16XaeLxYj741a1hDZof0K7uvLEfhDTqij+kJuAz
K2Ut2kJKpSI49NWU913oJ6Fxi43k0nsL8lShpHYpH639jYuSYwDXj8nCAzuLNufq
nr4wZ6OhwtxiNoLq11O+nO6FBt/n2mf4TcCnL6JIcm5P09XqI82I1m9qk8mvYzkf
CcZlGZsk0KmUC8UcEB/dRmEaSGDslhodRz27e5GRq8mfyeecdsg/RUTV+wtBqKE3
SwpRv9nDF95WFYXY8hkAR92Qa4Vv5LsrGxPuQvKRqSQ0gItayPbsfSDoRM9ZwW4Q
Tb/QF9pce6AvmxOV7tTmCfAFJq8GX3N3HE+acJeT5/SCuWvbgecfc96Hu1Dnl3zX
wNCBmrM9TLNiITQkIEaGM6J7xTh3Hqkpt3ssyRlF4R8hQFohp2yxpCAFLh50ladv
nc0N8kRzHYxpYSxdc5P7f2bucVXk0H9cfVKsEHzitJRwS27uj5IOel+hMFNojBWD
3TVlWe+iLG0GB9pqZrRoeTeVUvj9dRZ+4eJyAIZnLlcjHahPDqhojl5wA6pB25va
AFcMLkD8H3jziAyXmoeYR0r+udvPQQ2NArEZQGxcgGV8t5kOZVQZ5yuLPBHYlMxO
BaGCVR1Y0TAHlyB7c1EVSHm6Cl8J7fVruXe9EMXhag+GjaqXK5W3t7PsD/a9bMFg
BXcenXnBifgVR9VblviOisxmW2XFLxb+cBTKz5zMN9HLvU/KMK1VRpWxa6/w116F
HC1scZDu1HcbkTtNn+OhEgJKQpJWHTu5rFfdH0n43XeZ+EZTgYbs1aDp1Wp7FaMn
FkKPR/IImEamtF3/1o0Ke2H5EodzVTzXQKKxNfoh9Wo1b9bgJklcTvQ3YqEj9OgY
72OU0e0ESKyS9HwH/Hu7R+ZwBJDeZamASK6zwLshxTNX8y5lNRv9vNJJ/vLo+85r
8+yg0Mp6onoPVR82xFsaopkqx1uGDgpCNLNobWixJPWYEZEDjoP4O1Fpf5BVw2H1
WNfyWzvy3AqUcbB/MQlh90A2Pc6C41AYe2AokA8eB+ZY4d6kZ5xEaczMiJCM/e0z
KGNS2Erv0d+rFWFhIDFotZpk+xHVNFwjCmQkM361rj2oBuslGLdAUq4obNv0GfS9
dFMZi0E2cRJdOZctCI3+cMGUJoF7qy4YGUE/3ZYgOwdtq36kjh81sQve20CG/RFz
uXhxyuEHPCbCm7ZQvQ+x/ok1tG0eBSF+HvbVR+BVQHIYvQ2oXO50uZTrtx71IQUo
5apRGA02s1J8jtQIzp/ZVD/zYHbLO2eG3siSsT/+cuvJkuuTrfy4pavrlYbpqkjY
EcLBiaOthuPVW3RuX0GRKK3Z06gnlPe91SqG0HVbHccAqhEpNCAzNwiPD1M2AEm7
hnNQVfKSAB0n1ENPhuWH0E9dIWi8YDipk+b8UB5ufUl+Xo0fb9gc1hObvyqsV144
E8/+zv7QSlb+5yWMDRog53UpIYFk9YNUdJX61xu/GX7TL+Zoo2+4UPkQPTNu9fnB
qUoJNtVS4Y6GeNRh2nrz+M/r4OkvVYTeMnkT8tf9zX1VdOLE7zdz5dPTAYC88RJT
bOGSh1UTUnnN4EPDNBzt59MbO0TMu9GE5OuRdKwmD3Y9M7SIrflriPTcKyAgdv2c
PkXQWakURQh0TDHlcklSYz4qQ5bK8kcHv15F7Toeu+Uhnr+7Vh+3uwd9FoEnlYtk
lppGtr6kcAgrTrR/t3JlSKZZDeLF8IWkLzYL8DoONlZt0fawASor/u5XAQT90uRy
B5NTJPdyX8TieyEnUs0SBJusVx0rWdSjrEXS0JSNve9ZeBOd+arBHA9iAo58XTq9
8MNJxIVVGuOFylmHc3X0zgAKcFv+iZkAKXCEZNieEj4IxwNGwDcFPI2SMmV80UnY
gLIdDG/cZT5/rFfHPObWSTTfrYW2Jq8R1va2hq0ok0Ef1UVGcGOb0DbkGfsf32pL
e6U+aLh7flu/r5eKak8aYkDr5tpjKGWEVaB5bCWnUJbxe17MILVxnwRCku3EfYgk
kFa0hrcDs7zqzKabyT0notZJUPiJhKgaeIyMIem89urUhU9pcBT4i3Fgde1PasPp
EwAX7DS4kTOYTkZ7tzokivzXRZimeD/rPON2z0t5J2IkpOhhRJJV+NgiLAxXyS31
8OWi902TR91kYrlqsZqXaK/y6rE/XJsqNBQAbsHFLe/uR3jhE3ovOYwNVqJiw/IF
/dfMMcUtYUVVH06r09ThpfnA2vYmpY/+UFNCPy0/MCiZMluNM+bH6ahPUCZr6Iep
pAcIIKM6PZoKV5Y2PtlElLxluc0JAcwFpxb4j/ROip3zCQhk3imrurHpT+Js/uBB
2QdmOrwlHc9zieRHWCOQdakpu7KMxfyezezxb+fkPzHpRHsuAyw0EqXt+jwUYwr8
H7vBM9TEQFtqFzO3lj3yI2oN+ZckSZ8xPmIDaU1qmTo8guiTzubQ5J8J7pgaZ2Hu
1mDQZFboecniwKaWc1sMTjCoEZuhJoVnxpfglrR0o3UcsqUdLicMi8SfcAwcnfYH
GsCL+hqe9QuJuM2TRS49m7y9bD+G8dlHciLrh5dkNMphxFY5K3tdanYq7alNmAH1
gXeD6A6AtGt4cV7oHozFsbrjVgteIy+IRGyCVwNLIBQ62JwR+a2qGELM+dT6wqNY
/K6vgRbwu5Htfe1PoPuBomcgVKXbNIRTOPeH83Xqk8OXiutbB35oUQDsTpR+BgLV
rE0Sl/J8un3WJnSEMHjyp9hop0GORTHnxwTv+ikeUIh9SRj12KtRM7R7zdau4Ap7
+Kd2jq8jhF55SE61zfKLP9jklqLkF5/kinfQ5R5xC1lts/8WRZqUlRVr7GdEETai
n7MvzH5gPGATf/cgnYvJdLrxuVg4KVh5A+fQb6UJ06anlFp9SBmAzKZvrxvSrjg/
7aqZtw0C4Vs9UM3+z9Sx7h4dOSfKYcQG4SA4vkFbRfK+OhduPxdAT/N5r3ETlfKP
MFgBqW4XBWhe0ZPsITV8RReFXHJxiqJazHTtuptnkrLT2OIjJEmnRXYpOhOfJ3vD
rdl31SjYeg5FUO3v9sUtL3sasLkmkyA3ODX8Mpthcj3UHAMHou6GYBKb6LtBNDXQ
AETH+5lLBKf4GwKse+VnpWEXx4eFZPsnJLJyy2lUKTL8ZbWxbJ2b62QoVQ0gvlZn
3v6YG1oTEU7FbDOE13beza/Iy6CACCiEAzrVqgl9y8JLx8d6Y05xcRBWz8Rh5zne
RJega/4bDXMjNxblzFPVC2lPgaIOhaIbN+wd7T7p200OGlSjQZBC6fgKOOKqKTqN
U7RABleKWjY5XKT5RcBmsV+k7I3oAtF1XuOlj4NdGDL3jzhRU0VkmAdAL/oj0Ov9
RhL7KwP5g+Y45rfoqnmpOY1Ouus/uEA2NGwJaCeCmhedlpIxQd06DzP3oJsM64td
Us5klwJdyMkm+526Z7Sh34/vInG5Nyb5WZUL96Yj9Vh4WfMD5rMSH64XmtYZHJc0
ofPlj+qBzbexQ8hbfGVkdhTo5AeSk0Gb97gnd4vdAxyvBA4pRrVTbm8U11lrf2ZQ
vNlgmSyYHMVv4+imetiFgkiD/bxOKB1PaT+BOXXqyhnlsq+HcFP/MH2jERRMOO+j
1J6sPhYKciNMyKvNoy3lUqo/CpQmSKYn8fFtLCZwvl3dgqqxmoDyWZMLNaFSjgcU
eGfKi63IXhCEHMtmoRaoZHkTn+ktTwFA3qMYdMQi0bzF3JgejUEMrBT6ZNNEO0HZ
5rfOmh2ymqMp+vr1XZ4tS2fQ7Ja2W7vRK4X1bp1dcEXWWDhCUtXofvrwQAwLe/bv
VuWAnhvO4PtvCKsea8o0DjsVUM5ED6mT8fPzVC67FGmPLl1GmGaRyJ2TEws4hH6w
t17/KBlh9xVeJafPDW96Boyv7yOd2KVKKxO8wDlj3UAL73J8/MrTXDQ9CotltW/w
HMaLe/pEAadtAD04JIpXI9VuBtzZbeJJVJLA961ulke5pIIvksdzqHZR6i71X+oC
IVZisGHsSyJ9vfyzu4aNTUZPUpSL1nVmCccUW8/JGthxyEOAFam1ZXNW9r0+bxfY
fC0XtX15w7EwTXt0Ttg4xbl7alsEQ5T7AQcyeXjie83twOCKobiXXlkACURRmORL
5aEoTJYKo6AgEenQCBzRjUl4t9tDzaMq8xPnl1KkjZjGolmoqjz2i8w1uqoMSAnr
150QGSqiNTBE+mkFhfEmnG0qf6A9S3WzKW7jfHdSy8T4w265f5jGC5odrLBWjfrp
4FGsI9IcKiAKi0C3ghoMCcamRs6MJ0GvRHSat6puFsMfwlin1h2Yh9CUVH6FKxbY
zLlt6Iqeqrvs+c8glEw7NEyO16cbTMfXiSgKsXmJcPrBs9VuoLldGl+HpnPlM2Dh
4nkcrfwB9vyjrtIHLcxLD7cBbgplImKK12DW6m+kxY7RW1y0+pzOiITT8hsmwPB2
LWtEj7a21OVLZ0OkH9+qKjp0UC9AvDqs4eacNLAxcv+cg7eaS8rIa1J38ZtpfcrS
mEZyUttzK6I94b/4j6+RQARVfomL2KND9xBkVDRjXgMGwRXKJzwzdagF8te8YDx1
sEtsaw0dF9N99+WS0OAMUxQ4tcBByiiqQH7Rqp1LzxsiSZ5bdqb8+ke/XU8scoa/
MlbwfyUxx9zeGQOroWVxrjhM+cNigo//psWiSJTYlpxGSShgJz6/hpxV1XJa/VF9
O/2WoUJlaGl07ey0P0xq04FgWUqX0nKpEJvp8cjxrNs9NxzMxc8gOJvySpNKSfEW
i/Z79jYX0nvPbezB+EYP9PzlRj179jZLeEUniiZaO4bBbm6GNRv1RSWBo8S5ScFc
gnYCrUQr5zl0LkctIIp9UUnBO7yN5XYvVZRQIt3/DsQBmLrA+zSN9NGKPiK7/5Wy
yY+PGX0YwH2+041qsstbSTGoKVzsXKS6tCXS9ZgdXqYSnU6A1tsLp5zegLYNmktl
TMxa3uUZxMHCRYBDB2VNtbIM0uy5cYJyN7nHH7GOkqYAie0M/g03vs0vXMP09Xxb
CUlrB4pOGdXrajhENCjKsyY7a1lN1BOk8MAdm/IIYNyPRC8TPL1qRD4VclXGtO1C
o8lPHzUxha7zamxjdT1OqOalVV7vS8HzSplr42TipdikHg5CIW9CwExBEDN9FZwI
KSImoa7cfgbKfTIS9HKCGIWKuE8LOQbhMBY8ICE557vIVhvHhZRmvqR+Vfpo10l+
3ew7QlDG8Pu26ZEnDtJ6npXTZ1B0ldCl4ljfNxi7t6AlVYa+zf91i1uQMYUDf5zH
dWnB/VVmp5yZcnNzfT3uA2FK4AyytyLhQjdZH64hSKEqsHpoY4WQEQ9VclpLp4Pa
u1tjgep0LpBMOx79uGs8vifN/Ua9OlyUVb50VOBn2Zqwka/yXwvS37ZLjqlQ/RS+
eZbCIGEncZYj9kREtc0MPMXS4BgIpisAW+j7Yh2eRF8jHM+sIZ1sgjVNUiaU0SCV
E48qgBAxsBWNcZMW1MRMWg0vkK07dovCoAhfINfCRF7YhnpGG6Rghy5Zbj8vGA8s
zdTsGmlRYMA/rtPYObgjic1TMfzvLsu7riUBzFtpiMSN9HMSNANoiAEFV8nHPgP4
P9THmU844B1rO0q7ECOf+LEUkKQGzr28rBEoOo9x+isAx31isudxzRW5DZdTphYb
fd6vpQdbZPTF3Ckl2ROsIR7vHgPOeHArvByAJCqiwDgcnHfePLLTV+hkDDRklahR
iIvu+2cyqss8DMMfuy4rE66jB0wDkyGE6kH1LeGYsj8nuLzT8bTxK3xfRmgT3ZxM
VxFsHaJuiLObkT22U4mHFyzOP1vddX6hUxcPqdq56AYn6fcdaf/0f7zQNATjXYGJ
fkReyujm57AYeh6XhlBiLD+TUKh+pZzAtW+6sH1T64xE3JGA77FwR09FUOIuSnpv
dDhYMpOsWVdOCRW5nMG7Z/aQClFDndr2S2Wl/ofeUeNxBhJoYFnqwMCFfpHveWR0
FbOl5U4SEWi3EPB5JgXFoyygHS9Uad2qOrLAmD+JUAI9XIpt94SNYeaGa69jwtHK
JD7I/+yOOIkZZuQlbh55AmEg8RyzqlJ1vJfWBH0tLWPONu/8d5tAFjpTU2oA73Gx
APl+OE4Jo7oUEameb5oduqfc9pNkkPa6m5dlfgde2So5StM/jhAmEtiTLZHV4a+I
9kHLylx2QfntB9gyIYl0fSGvd8DbMgvdru/sttpKS8nk5rsWSZFcFVgKHymUCx68
4TtBoAdPqlkD/bWPrdwYKiJJ+0KTtwO7NYqYpDzBll51UPLaplplls4rL0kYZDQl
2SUf4ODOPzvQQFaKJ0PxWgRJn68jFYxuVsbVsfeXqXJShBqYQCiDptBmnN3fUdlc
E9usH9HAShcC8DwnjjJn2mcvg82lNW7kAZRnptJZ1lpGUblqwd8658r6H2kcHD/X
OgpoTRTgyFQLe6yeSrEvCgq7LKHNADzA139LSdqJpEtAk6UtFYcUFcBDb5s/Avef
pnRXQHh6WVMgN08CpdhApZ7o1wJhtkkT6hDibF+HCfZ6QfHnY3gfQx22YJurYaaE
ntkTQZlSg7jy+n9PJ+ECeVMfnuhb9435kBQBOOpy4x9HlVUqTW3BxNwSXGJc6hSy
Lf//j5RbQ9ZACYt8+QiRncc+R2ld+OipAjOCtP3SnaVX0UjKQAe+2Trrc06gJliL
xGPKjl1zQR5qRCglP28lYspY51RpfEAAF5xx+axnneYeT1XghMzXwpWbRDaxL/cA
oyCZ+lPHq3YiaCZ3vTJ7bl3G+mbwhQpKNCP5DGVYpT8NfOBWYrmhTVmSPTRiCF9R
2LVZ/NT6ei9kbSLxbRvxfl5OfOVS6Ik/MNBsHn/7CNwOrVrXTz6bb/1gx/epFrqe
F/RwROLSbbx6vGo/XgrX8ZZhFyUhi3PGVDMGnVNhLiaUo3BjwxVuWxky2ElWqWOY
Vvw/jKzM8J2I5a/mG6otmrGGxvkL6UVUKsn0OCST3WJtFzugPT/KS9Qk/WS9bJ32
Ol9gsZ3UALrOzyrsH90gyZ+MgSHy55nS+Kj7PeryExx0I0W2/wrnBhdJWmqPVP9b
TB6+Ha5lROVJWXk+38u4FGry26Z7A3AmIeoIhHML5UNdEBFhxxoHJAkAFFY08nVj
1zui8jmt2e/Ta38CEckOA6PF/opXvF3tps5Nj/5XG12GxzXk3yOLauehyaU1/wIK
cIqYLmVqJa/f0mZ6GnH2jEc83mGP83iM8c3Mu1FYl5/KAb3SkQ9U0da4PfbNc+Ky
oS1M+EkX6xBRK06GamFxXaf3sIYud0eSbZZgp738GnPLCsLLg5S8gTv5wdTxQUd1
U2er8pGQsAkQ0bcH7BJs26uI5U2kx09tBI9DfK0V+Us6Mw93HH06P0880eOeNXi2
fZj/97upZmD4tsgEBRpBQmHuoBFQNK+xV1ughZlmg+mdDd+NVpJJ/JOi8FwTFeze
ERZi6wMEIMKoXj66N7heIKPCnWKnKH/8W0mBO1TmRkJ66NGH1E5I39nE8JwPFnEB
rL2Iz6TKzZ4k8duso2Sx3qOf+FGOfNxMxNLJP+h726ZqrTqJ3NGTDgkYU7OcSE0+
uJRTZzBuEjenM0+ilHNCh4S3wJ+PULtfrjj3skFGES/MZK2pALwgJONa1z0gd6Hl
MfZbhx/Nh/84TPBC3PSlhklX95uEmEdd43ZLGE6uDgGWpCMIkfLxTF8Rz1sPSoCj
XKBvj1LrMKOLtcXBMFGcpIylEfB2R2PrZ0/J4aIOjYviZN7ByncLPg0MzOAe40/M
TCc8iPgRca9ztaznljgQY1LaULioAhI9gz829xTEyxTh1C9R8fsoWuM1oA/KWxD5
E11TuA5hpu41FzrKmTOfFKCbB3ciXXYrqp7WDGsV9uMFjWFo3E8fsWdmgtrxntER
EXok9GzbA3mgM6IBi9IwSAiWetOPsf/ECVUxPULVAwBwbNBOJ1vvnGjk5X78US47
OFRflyQjeeuGhvOi8h28pNPJKCKCSvtVhCBFN4tYZzZ7qhbUS8w1x8jYBdFJFF0c
PcaozHp3uMOZuXHvE8o/aGf8q3fYmGawYKG/BdTN6weznJzgJi7i8U2XE0XHEBWX
bAD9OgaxJ+rUu5GyNHiNBH805UwAAiojVhdISPux5PoYA8zYP7pNx5khBg1n0HXm
tfeJGy+JlP8FPX6LDpLQ3XgzSYe73rBI2EwRIcI2PS+M0af9+ABxuVzK/jdG4aP8
Yv+8GlwmWHxYABPqn7njJviOY4kUp+5geVZ0Ak/enQ7wfKjBqDpXCFFi7GOXKgA1
P+IlGV36zqDFujo0QuFXd8bMVKkPpl6iZeL5UA+39/s4wMCcIg+Il3ujTdXWMhcX
0xgQ6YdSq56OXwjYa0uz//FZYWV/kdA8CyTdRvxAfmP2ejTzrOg34RbezBJlJPT2
uN9jqTs0QeMWkD9zW4VTjFSMmxUxNLgB4a/wlLi40LU88JCrjrFYRyIX80A5ZPy5
Rusvd8gGGHbWJkxPmb2xU6zvm8aZhbvmqeBMsXosmFybvo6g7LUThAZ4rOF5qjHe
6o3Z+lD0SWdbjQT5nCLn66KmBmyZ23Fsp7MnGgHW6uUcDiZR2omF0guA8k2cUPtH
hFop4HkD4xD2xazf7goRcnJGSKWVRixP5OKH5IOrHq5UD1SDIjg5HTHBbSxFRZcH
hrvYX8hJUFFK1Lc8AiRnGoNm6eyfLPYWlDX6VV/G5zXmbPh4tY6BT9gwnSxpC6n+
LxVO1A0aRBk2khLpouqXGjnKbmCk554qglZoNQYmC+itlpP+XY7kB4XUiG6ffqtl
8YqmHEKWp+MrRi0bo0eKedrAG5zto741ZbYX2x1pXuIIpQuWEeAuvkrcnf4erSGD
UQAKcDri4biXEv1wpufKkzE55pLhXvp2TpN54CcuDCT4kdZLomGSBZMnzfHPhVWl
JpRO1BN+OYLalLl/Qe9gDhuMZpuXjMLzS2/sePVbADqKpL6YIPXZE0yZ4u2q8ESm
TOq+7uebfW7PEiqCnl0cE3FeRQaBjzjk+VdrxepjurYSkDBlGmRxq6RHgyYAhyrc
hjD+t8UTXVP5ViV3qn/OyUbZVBsF+Dj3AM4YAk5eRGK9iuV8GOeS2x8AewerilMJ
fjnkVWcX7I5og6DEtwCbNzFGXANfGsYbaE9m8qVT5BPmMIfrS4jNfxYVWRTTR8tQ
Kg9wszVqYYqJO/sk6p/EgkzfLptWyJsHVKdSwW939GOdOk9GjIOLVAC2fV5mQP7k
aPxpqAZGThlG2iQBkUvDEMI/+nePZR06fb8UUMrDum+MgrLiQL43GcCvvnzOZH/i
kpDL1h3iZlGY30bp/X1aF6Bw+twTt7jDAJuUHwaaZ+gT9iVPd/oQwuOU6iF5sJeC
etH9sjAO507pdj+B870M3PZKJ8wiJVMqllGiPvtmBfoArUonVOEmm3bpLMuEzW8x
YDfXiHDY6Ie8Hjza2OFluxdoYDgJIQuIibUh8yDqf5WzJnCP9SkRShcDtC0v22pL
dxenK2yEF0NEcjld1eEz2p5rcVyp5gxhSnhad3zXGw21+LxAHiQKs6oFPcBqyb/3
IU8kgYD+mwmZ+5mjg8flZaMP9xSCwZyxIbCN3ZSeXEEpEQ77QWleYmABWxyuA0wH
3JcBP0dch/COf5vm6nW3IAEkDsVVU1t/KxWMECVoabmoUIUjBmqsh/RgjQ0HLyGl
JegYHiLPxpW418+QW3HgBU9m3BcWKVN8iwiHH8N4+VC9ybvk6h5QGVm2tP9R53Vx
34g6IWGHG/oa0IdQH3uAXgeZmQ4KkoJEOz22gBeFQ+SbMcsNmEksleCm23f++wsQ
WwIgjUdJHXkf+HGXHDdYb1UZpJ/D3ZBb6UYRenfDvTLXQnT8vQFo2E7qm9DNoEhz
QbvH30zGm7WR4AIjOGi0/7FSJtzHHDIbHAUqsynlx301hmBTfCdO+fj2eUuDSIS4
6aJvtaiEjGhEqEhZkLd08Xr49eZJThMA3s6Nyk5I/Co84rKAI0hOzlQNP3iNjLjX
MxSl4jnjkSXs6C4ZgL8X62J68CaCQ5d7p7IFww/PgW4Urw8y/ObTdzk8d3heaHi5
EyHqICYy4DMTrG69ogQcf1Q/dXFQtSlqLjbpH1Um9jJoHprZsakQ35PjnfO7HCNs
+GZluV2geYuObbyM5O/IvdtwEa8hi9YDwTDh6Q+leP1xqBUhPDThWRpRy5hhf0YW
fnZ7WUwqYlSfDI2lfEJikSRqazwPsoFEn+BWYTynryAna11Tmc24pREOs/Rj0Kxp
/bk8M6UaCG+Z6Nr7a3o2vmNAqRQy7r3iAwJR06kZU4Met4YdABmjexwjaQYW1JYT
SrTBBDCKg8Ope/Sj9scpIX5+U2OcJpl/oBtktOgbIltw0vzEgZviqCLeWVBOv/k2
V6xjD5ZqBw6d35sCag4L+68+zV+MhoCwZhZ2yOX6N5vxTiZjGVvudSNlzBMds4/g
4ZEHzqW/9dkcQRIa9dg6bbMhAfZ95Q4XCyYBRwIpG2/FKm1liFsw4P85I5crX/xs
BHjF7wDeT5+1+/luz9YmjVh7YxZDX+sIYJKhvpJJcV/kALYb8uDyBb1BGwccElUS
JBWH8omjUQPOlLS8Jd/L3VK1pDXzJxpn7DireB6hg+9+KbRGzf3/5IpCa1SFLpCQ
XxSOToOUmkPcSTP2N6s/U0sCpj1DB+u5y/ugwxEAJ6PyYfDGsEPg9cGhaJ5EwKCh
HXsRhunhdxGdwWaS6nvyxnArgIzGywuPa1iko+bx23p70qYn739XqKA/+dLA52D6
B9XhgSgJr0OqmjxrahAAHg6+ppPtC1bGF/IzhSdTQIwUVJroLoKGrUL2iH0vXQEv
7XOEGtsfl8dk/w/PpnK5wE7qi7Qqv5zxaGbH498LMNlMLMCFIV4YutQ/eaWdEM0y
P936qknTbTnOMqASezgd4uzqT9tCqMVck6J32Gij6ObcEzrZ1wG4yzg8BudRr0Lj
O6PCJcBtRE3D+c2Cf9xLL2bYHCjDACKa7vOTaxBKu9+pqag2GR603oGBX8EzCQFR
O+D1IadVXBZaAIbYimcFU1zcf1HcKOpY/pZkeZRevgmM4w9UZbx7k9HI5fjiavu6
LptvVY/ABcB+NK6BRVddV3weyctq8/4B3bhDOGrZbZFMOCuv59rZRuPpqT3R1uNa
87v5Wt9gi45STmIZybDwcx+POB++1jpzBC9uMStWCy8WAewlB9dU520kbf30Hl76
tfr2Wszr6ldTpMBRLycmRpPg1Sy+M3Q0kK/IfwObod8BjeicwUWPeBvc1hMyYoED
8fKRs5meYxSbuV6xzGeNJbGewJkMsRpnonvhwf9kM/43Wd/dckwlwggFEezRzj7l
N4nseMVLr4EIjEDEmzZ/6e/51mbIVQjIIuYYNOUMpConmfjyBbEhg+YPX3bOOQsk
aI5HSqaXcAN1myQwksE5adamOxvSCcFZN9nRoqwfpIuk3AuAO3Tkv8vZpnl/8p+N
IhZwEAvxYdUE8URtcvWu5RjRHGaCT8u+9BfxKXGQCUx2PbcmdDA89kdZk9n9hTkH
3BajVluhBwV1FKk/4o0hxG0L3MhZQNgMuLsgcYDdD+Cp4WLNC4jcIS3QQ1HsE8nc
oVXq1yT9UHksX4XwCgaacHnBs2zH+nzzPDqaO/ZTT37EiRQQq6rPJ/9NvTC0j2DF
ZbzBEf7RPSUMFXE5BxebAYiQt76CxJfnQhinNNBnm/aPDx92rKpG38X/eGPYjuAh
ozBlgTQb/v2lNjNfmmfi3ejdrC44FFAb8O7x5SjNFtG6aAGlQR9yKTByMoBujXAX
gVxuZ9oWsuJe+stoe0plcXrmxvJuUWMQuxSmN3Vcs22oSzHCn8CTSPiViBW9DiWX
DRxZuyYl5yV4AkH5WUQhkHI/OaX9MZkafs6rGgA51JR+a2A2XpRSltNBOWv+y6hZ
a1u2AEdRO+4FJ/U3GcyYwEPS+RwrK05p1Xk8PuiWq8H6Y+MzV8iHA43AmoR4lGtW
mC3Rq1ErBRL4AKxd3BvJXkFmYLXMGYWZqANSUTti5ZMWpJUnyBrBykMZpPK9QWrK
BqMDAWp4pQBrl2k4Hx+4m1OCG278vToJe0WdR/1/xTSAmboncnjyj1XCN9fT7043
mQdZ8Y9VWEN7ojCQIXovBWKlw3oZHAezbm3PQ6FaN8y23i4Vr8lCa2zChmLXJQ/s
uCRMJtfz0Scyn2AIEHkvA+Tb0Pg9HLqq19bpjlc0ICowZwqk/rPiDFf78Kdb/lOb
SFUZrXB9CpWu8k+w8+a7yyAbtwtFJTIZ4+Ok3wa0F3E0vcrr99g5/mJqUS32WK6l
4nnb+Ex+km8mcy5ZjWBNXllZYhrjGZJGXuJ/0C/tWqrpgaw82YL3MbLWKAEtPgZW
ELPE0GEzXY/VShs1WNQi9Vo/+QwoMuhIVElsBG4ZHXG+KGEXWJBMSr8LpfY3FZ8a
NSkIBT0hinNSUnnU17MLEVQj8nMAj+eFijYlurVxnDaYBHnWdaXGv5R8FDGjYUSA
bwUeO8KKpTPEuffZ12mrvzQ/woqcIfZ/ODOpLrQ8ovGQpq+eBnnyqRHbVwlcBPkQ
CZ+coKEusq2Lxv5XaFvin1NRB/kRk9dIGpn1xEFy2cCCOqTtl1xhl4VmlkBDiAMI
ellFz2xdsvX8yH2RLynuI95DAExCOd7MrLt8Ewq9Ax/JMW1ipwgtDHpGiLq2cEoH
Bi48a6YU3oBd6DilLl4URaOev1C5vDLp5g/WZ7gk9ORU82KcYes+sAdHShoc8ErG
lq8J+34cMHc3DqL7Y+T540Co+9C2x3Fa0bNpzLk/P3haQtTwgE5Se4fLCY9sYqWd
j0xYB5NLnc56VaOvZnQhstS1A4RIJAkk1RV5ZnJDNQwjSITfVUjsCWGFOxeFQz6+
dE4Bt9UfpIkh3vAdq7gOZKfPLj4ZL7TjUjIb8qcvRTdLpszlDqhG+N9JArdRFxs4
JrxcYtcGtK+0/AbHSsGyMhqOda7hVd4qU/dYOub2g/M/0RQBuQa/xtvWbhWmHKsa
b5AfI6gIxJNCWW15BKHvVVkEwOyQoSTSJ6orLjWW3eUWgMwJOksCxTZ1WYVfBNGS
2QZKFvBs3nbFTXFw/ck9Ely9FvPKVAAFrHl1YvcYr8Ub9I5OEOQQYNn+DC6UdIxW
c7kiz14AhlyAVjcNkeXtGZAnM1a6enWNX7+pwlrjfUkxyiM4C6T7EpTkRRBdR+bO
hqugLeO6lhdgQofznhcDeGT0EUbEMwK8MoGNVcBbGkPS1VvBp9rCfnjsTuxLeorM
UkxEZmGs5ZjLRZaiyrL4po4FFkd8PJ1NghKyd+iFxgAqFhr1nIb11Ya6zlT/iFlr
WF4rgj2dwRvAuBbfI3qH+KIH/pAW0+N0hjAa7XwwXtrteHd75RYix5jf0GkUwSTH
KRMCs7kj3sCqLHW0Aj4rnPPw4Yb/j5viI8EtoF78f1D+jNG1MCRRXh1yK8dwGXIz
cQ13DZnynVSIaKPnFCyJ7XLnz5SlOHzE0OtH3MDhDdN2mGcpWkVJYwewOW+J+H1j
uCJH/r7dz705H28ZdD0T0diNikIY8lmORFuf8XqgfmSiUE/PJj+cU47H9NTUHjO9
M6UHXKvXY0F2+V+eQXsqkRLE67MjUYWk1ee6cgn18jcNQJZgTbUth2nglGyJBdbo
kHbps6M/DO+21sk2DHpY8hgMsIas7eNA/RuLXw3uxqvKAaqVWjzS9ZEmFsm19oxi
Ha49nxVImkhjDXKyokreKzx6+PJwhxTQqw4l16ryJNJDctgaiUaW4Qfx2fp1vtk7
7m4ymUmiKwQessISqK5El+Fwq+pCiaVd98v7TfGpK3Dbnu2gjjnZIbMZU+7RqmZX
x3P3Dx3zsqM7vrZp5KkmKKne5HUNXO986/EUj6H0Zlb4UmDEiXE+UXL1bcKh3zj1
wDTe/2mMElTb6ABbEKlrAwGJvNyJkjhl3SSkrWZ5IdGldTkdoB8QqMysYUjMe9d6
aobwXJ8eTcFhLyLUhOj9jzb2Cbx/M2KQXfU9nigtZujJYlB/Vgg1WNXSXXE/SFqR
fQHPUBjCQ0PoOEVzQT9Az1ezKMRasgpWpAQTb3ru4ym0B5qj+Pgd1mmPIWdz4fnD
uALTVElDkSnm5BkxXPqXSek/tJtaBJV8mDesO0GvBCIiEBgZbfR7V+8xGidDCXpO
UwJLltPOcHuJIHBwUWq6I5m9Y3V+xp/RVn+wCHAjTOGW4yCcoSAeUNZGCGjF7X3R
M8OsfnxCR7HRIH+yZnJBHSQwzNJrblkYIp2As8Nki9JDM5ARb9J5eahxkoSThK+M
qCzs5og0DR+yv2wg662bxw5QwqQ/8sEdRMJcH8NRB/DewQqwMVWWhCtay0iVdwZB
pmo+SWkpNvFPhXkuijq555QhULskqCJHpF1+Y3dfOfBwxjHVsA+cd9BFQBHLpEBA
58f05hSGXN1w+W9IBMtWpnXmBD3fbwcZydOsnCP10xKELJlDfSTW7jb+ihpDIKLc
7ZVQIjV3vh9va8GaN2qFiumXyi3uqwIxeE87sEYRuWvwki9NqXRLwf3JweVIfDe1
xlMeudytfEKDcWZm8iQIeAlTH2wMthm2lixdylCYdAcoFGIqnJM0XTLgJAMZiYNx
3C5XaaqJZpQOtwVJFaCZuiKrtOluLxX8o5F5LMSAOcOPdRMBGPXK4LKnS/bhtAMb
1kzGYZKGXA9ul0wIHjPZvzB4fqA8Mf6yBLJ5zeSisi69FtrtZpHUsZP/qoNMdKIG
5LMzZ0A98SZ3kQsykyfO8L6Ag+zuNF0FaF3qVZ8JMElPYkmHBZ7cTic7PwJTltNW
2f5M5N58gazL88YTzQjgV7waTg+wtwHOFdphTEEoBg1VYp/ZYYiTXWEW++eyv2Th
/ZJAlH1FTbZJLNhAKGCCayMujfDGDkGD2IwhxKc3RRIwVNFrI47IN93m5OWCvamX
eOKDhVeCfFxAtukncJjLuQhtZzJYwy0RxErwxj7ovrLahKM0x2t20bTEZRbOPIAY
dOe0ktzfls2eQJn9Kb+BDW6IuO0Z61eqPWrV6gXdRMH+omhSE0JtaZwUlC4CXV48
Le80dW1gdmMArO34N1FQJYMXIGiw9KR4bGpxa2qxm+0q1fVxBRwWexff0mUnr/UH
mVS+j3qot6k+4YetYY8F/Terb1hfd4vAM5t89rvoqSKZ18LUb2p41vAQmYo0DTEm
ZBJzP3iKN0tNZkOa/q+LFV2eXmj8spayABOUfmk4nQmjGK9254w7d2PuuPV8qUX8
X6NtRge+3eHyL+9J5RuL2QRGmQiXKxAignHc2wK3Zx14QLd2ZNtMCnKjyOoYXrnN
HHOXp9LpPKTlQRWZPAsN+hsRjkjSUd3dG5PgHG7XoIL7MAF+AgJpzuhn94b+FHaY
N8TtcrWACKKRCzTL9tMtQ6RJ2JS86kqM8T2t6VR/ZSpHRvhy7cx9khaP4+PoxeSI
J5z+iGudVX8NwZYVQUS8Yo6hHrzLRJpdh5eDo/BhRVUr2eKyETsqxSbQZUwwbUjN
FIVOlxThkPgymaS/t16Hd8GhV3hHAw+EOZ65KLEFUGIYgEAqWRzOh/pMjq4MhtRD
xi1OLWh6GMzRZTe4FXKB1I/VwMg1AMHPj8/VhBrFK0V4V63bmQw3+yamKLPeXx1N
D9LNb81vgUwJMXJel/8oWpM95JDOOJ0J7OK5x2AMeX2CkKauSR8w5xxAXoHqmfXX
Eetaks16el57/21OsM/QDtbXrpamQmL3wivbIYZaIQmZlnaLEbCEsnnIDC9bLiiV
UchYTVPtsFOCWrZSW7DCjsR9KWQmrEagC9X7tDGCYuCqvHawxxL+mGDZPyPB6SSG
T97QCT01CuN3HdX3tphkQiCKKWcAqJu+4bv5tWwFNFhGHEy/Q6cZOpxs9vqcOqqM
pqFLf5k1n9gsmv7oUpPDfCYia8FAOmud/wuFcl6Ezux5QC4eK/WQaMlU1oLBAULS
X48Qso/hbX/OC1uUFI0D9bPFibSG55hsj+7o6U5uzPK5kJnM7gN/UWUYhD7o79ke
bMFDZypEYj7L9xJItlEyQXcTHMXq6D/fomq1HJb1JNbpbRkAmGCHdZGVcOuGVfMG
RNolWvhq7idszxqCdhYilrFngBzl4Q2gx08+1+9gVAbx5fL08fpFGqlsbTQF1u4U
GHzbVA0N25XS/ImbAc4u9+zdJPsVfBDcVzrjkkw0w4UPPQ9qHlP1aAWJjGOJk6qY
4rSHiCM7qopOgIByXIuPTr5euD92EIqxc5gkaiyfH+IZPvmPLU9JfC9oAWkowRA0
ilxFkavAWTreAElXLVGII6gVCUexf33m/FWeq0GAdFJ6MRwIh+O7dJryTSXH6Evj
1TAq64ltBtF0/flHAk22awK8KWdOmDP97eY6V/qVJJnt2O3pWSpOmSWCbyztJNw6
l/6AoYFOpA6LWZu7LtBYGIRaWWrSfcagTUtF/+SxZg34868/KYzW5BnCF+llNjO6
ufS9ngsCO+pjBz7rG73HnvI3SWQzzcdvFqya/ZQK0Cz42mHwWaIk77yHoO8ecvKU
cJ/NVpX8qSpjQ1+1sZihcj7CS12JoKEHI7cBGq2JbBffnK0/aN3AMuM8+4UY5Zqy
FOZLDAlvPm26Lb7+TEEpb3uSEYOpl//MpVsoTt2Fm+fEqqgJP6QB2b/4D0U49UMO
58AQSqZQFnrzwyQfaBOhzSH8JifJTREC9MacQ/QbiuyePr62RfKY+Y/bnhhrButh
kjSxT7fkrKW2zIWNfpqmHI4TnO62S2Vou8oh1H9xM77mydorUGRNZFYjSelS/DwW
GmeSod+0y2AdSouhcw43kIGu7diOEPtd2kep4zi51zSRESSDkhq8jDZyDkg0vtgz
T0ByY0sMvDdckyTo/Q7d84ck92h1N+799eKiEvAw0TrDEEqDUrbWOfrlXxj4hOnh
1/FgNhwo2c/YDMVYzbjGOPDjYwFWdspzTlrXstq7NdvctDtBWp8ZdRcoNkrp2xD2
fCRkf/hUzTYymKRU5yTENGxMAnnVqIZqS7owE4IPPb+Bh6a820aIe5F1IjvalTF+
75nmLPc0eUDRzKosZiyBkn26Om+pzOmCwtsYPkQU3oekCi+FuaDmo7mSnw09nr+6
vzsNR2/7vwbgRnA0LlNrsE/IY3uOnBuXPJ/wOh66jXvqXQit1T2Ggte9vuSsOXhR
m8H32d9DZkQ9SDM+E2CGNZLJVx0NsnzGb8XTfOwxtsuPsF6cIA5ZqamgYTX3NKrS
SmDgaEXZXCnb5Gx6cVHRdMvd4Z6D73N6gOixmoPWDYpeFzIt3hHjNWwhrvYZb5dD
RHAnZIxoDJhm1ZkQZOGB6X/9mQ1eJFTvkyBT3/Y+RIU0vAmYFJYNWcRwE02TqXFi
yAW2UB9YB9HbMhFXXBd+Z86M1ZfgOxtwhvkuhNbd16JCBFTwHy+lzqxLinvZ5uzH
BpJRs3Ls+9aURFLlivKweikelMUvaRMFw6SamYMV/hraXp1e25RhKG68iNGpTKmO
3d3Ufnby6o7pMb6JT8WxZ0Lfzh71sHUP7n/gfdiTolBPM9yPd5AA45kQaS8EXoKV
EV7m5lWK6i4HK+OC0o5is0sDl0ckSy1MpRhPohS++fVLv7Ow5LR7x1nWbH9nutR7
trxw2PkOEfEAC+uwh3RL8rKpZ9CKBNNn4RDXdAL7GFekC3mfOUDyQTrwBSk9nde/
7/26SbLauOGX667ocTT3XE7R/OLqKwPIGBZWMiOLrrWtTfq53Cl0FmlKWGdSDSUm
pQqH4j/1RU/UYxvrI912HbgiCiiouKB2HgN1Q9Ba4YVgDnzlPnL8HATfrp8+w9DD
ZhTV5aAVYu+KK7MXpmq33IIIs5+K2kR0Ib3RCSXSBDXVlLHr7O94db7oov4Ivh1Y
jypYAi6TJJ3o785rtngV2AS7iYmtu6jQ8W9rlDFIqAU3HwGpK3PT+y36FBGzXaq0
ko+l6fZNPIJOHJXIf5GNwXXtG6hRwbb+Ea1TDVXBcPJH1EmqNqD0myRGpVKUvZtt
ltzG8H8BYElI7Z2kLWQPEsIHoTALFcW7bZJkWTcUMDXFrmzYfqSISI+29xTpIcw2
Z25kh2j6K7qQLbVWYWxKSXHxCT5/ZdU0cmOvrwM0DGVvOgpqjdQC+Q32iFiJIe6X
OIyn7oOfowgbvGklxvcIyE95Dwg94ZWZ2ZsG8dphotT8LiZLovY7q0qQwCaUH1Gu
RknL2xEmwAPrPnjdVV186hZGKE3MAeQXvQYCxJ/rurSZpy0wF8WdGykZ74+zcVyn
OeszTBs1/qK7TfsRrsfyPuIOhlpy8bTMGDmGx2rZYZmhzJTVh3/tpU15zkRDjO9x
fJI1KHVQCkQrxPkGnFicEcayIY6VE4NYvxt86zNA2LiXOloLbJyqrX3Oqg3sydHn
BDc+IdgGj51s0+qZkNi7UIAbbsArXLzAd83IBpR6aAylhjK7jy6ftKw5kloeGYKF
CoRTO88tl8QpUbRzXlAFWrer7KcBT4E+lnq0lXmn86pQf5iGFg2UwxRAuzUWoHWY
I59PngGSPl/YtXBgGtDhJO7PzvziCDGEDCEYqouYBiuOXXjCAOiln02x/k0vg/La
uHKR62EoOS19d8sZZRJlp6zYZ9M1FRph270woF/n85d2rtVKBhiPeOGE6PoDuzWI
huwndTx1h0KQ+ebGi5hUKbO0l7cwX2Vdz4DzNsry4obmO6KXhRr4uEmVTOwos3bY
/YoA73frA2R6P6HnaAS1FooLav2IZxQrS9oy1FApzt2+4FXXB5vePgbeXykRFjRO
c68+ZbcInuY81ARLoHp9mWGJgUttqgbPoRt1aDNUtF8mhk6WZHSpLlZ2fgwDy+rR
9kzRnagh9h2Dce6DfHNDUtYBMK0sEhZ0Jk5x0hRiHeLCHMUNMyqDM0+dEYICfaoX
yWBRQM4ve9dK7NxVe/0lE1896xrG1Sm49LNnalZ26XX87n4pazZGWdhdBjIp4Gza
doozgvxHIefTVP0tKt18+9gaD+BG/cCNDepFR5flO4adWGuYBvMRm5HJdCKgGPzH
XgPkF0ytjcfIttpn2lXO6FjOkv/NZmmW6Ax7KuI6lz0IrpA/OfZ38Q5cXR1NsFtY
49MTF96QNcC5LCFjCYXeD+kJ0jMkKRrnWPdaSomu+0c31KhnucizktOy7GnP89ZY
zsHBfuyR/MC5JgT/UxuFg3h4UoCNhf6J4rCfQD+ziLWq3/D1tCymirI+ZRH5mg58
2Mg+8x/FRejzKKnoa/7TyyPABT7hAmzDB1RqedSXgpquwEpuV9nUFuBhtiE1yGRT
n+Zr5VKko4NeiGfL+DSSuU00zS8FHRuo2x0+0tH+rOo0yqHLzuSzEntxUjsvhJr4
NlgV2+8pzoLMZ2+oLTps+4zQbHPJA6sTv2JJAQDPafTLTx+j7l8PXNQof+1cqb/V
qL5gm589E0bMgaxz4ePr1hcfCRV04+tB0nKMgoA0j1qGes5pZdv4BGxwlxCYJS1/
s+SHt6athu49L/kc0IDoG+HjHRGbd18p7+EgC4+X0UFrgpUQOZuBDff/dE7O3BKG
VAnEnROEoSNWkC34F/6Td0r1dJo9TS0HxF5x6Ls0mtB7n1GXZcE0KuJhetWa1Dm4
o/NCWAKqkZ9NtOZbUsgKGn/lencozEdes0x5sUidDo+xS8jP5JscpMpQKqyAzIMv
YYG1fXP9csSXw8NbvnsH6UJCiGcmytFW95qASuw8tGR5Z6FUdvmKPZBjScOj9FAu
HV1GrWaOzOcUDRlSJMKZY0LqEakdVno1DZ2GKOza0nqMEmiZX7aGFbee6ZVfkDlr
wx9TktRb1YLT+PkI5qX8qPMJ/HoygseDx/jHCZOJ4da7Y3dI+8//cuEzv383fu76
Zf487MFZkrZXhLb8btFfJU3chjefyIjoZA1xZsFxC6Kd/dTd0XGXdVXWCSjtcObj
DkgChID4+ymP4zIjqLBHjdQW+q4KuQOwKyKkbNV3qqN5EovZmhpktwkFfv+qXwvP
Ou4OFjBZNcKIsKXPEjeMqKF6FBXMmU2L6buH9JmO+gd2/TkUPNbZHGgvByAFiZdl
PUTU7lpuf3N8xk6S0uaeere2H0v4CgZ4/hukkwDxpsX/F+gw+7u1sXFSSXvjw1Vo
1bJHNm/IB1FnRSAsG34IYuX/bJBCJp67AB2+fShg/+TXZOVTqguxsVvWsgNjSTYp
27jC63OpcUHEnVDbLMG2OzkwYwk0cjtk/D3znGT9XYnrRCMikLJJZzKsFpg0eTO5
R5vG0HdbqzppHPjhNuiqo1QWfFlGg5kvB6JgrkI89XdQRaJizww6/Y80flHHvwfM
l5JHCn0FsLllxSO5l5fD73CQVetHEvBUTOD0mC82Rc3l9Ser54tXbiXCcLmi7BQ6
7gik2eEDKKLIkU14Mdi0O0veJMIz/eRttCqUhUh2GY1lBMQO2OaFqlMX/FJM6BZp
FfoWRrSwiqSM7qqNgtXd62ImMAKWxOrY+A962OcVUnzRAgw08Edl8Mc+rhcEUIs7
hicoNt1ChQGN2zfF7bDP8jDvhH9+t+3VxUPi7z/Worg5rmaNniKJ2FDMf1u/jtQV
SNvndGQI5Qo6+NQ2v3WZphzHT/+4Udc56KUZUg0HsHli8+3u01hnETwu2tb+ZkcH
C9rFgfoMLJLRNSo5bnMOzT5MAA4QWWWInmxJT5UiWUdPMTAWz+lvTXMvivuZivhj
DMiptbzETjpvPvdoA5Lv0a8UYVc4+lgaV6wlsDNoPDh1R61zT2n/FQI7prJ1lXEn
1wBT+XmsRNxozSoeNZT+7psmV/7fOhGoDpB+XZwUoBGMXxqAF67QuluEEdYPneJz
TAojKsLH4GwTXgQzlqriCAAoSwRjEfjwlNsufAI7Q0vubQ7EoDCV+g4Yqxk2iC9h
BCeBdffMb/2YK/WuAt6IUwej6vO2fQaf4F8onfZtlvAbk+H1Hhcth8c1gXt5zxmw
LjQUwENfgVAHZRYTtbMSBvTXtC+FDh0Bk/Y1rWUSRKPe5U+XvhtDXbgCIub9ylD1
XBulZwGf9uz4bFOk/XQsYcyOf9FIvU/S2g4vKf+XpNlgQyxtJX29ANALGYEy8DOm
1IPzSr/UyTDC7OPV1M+HuFdEggBCJxE9KSLotdFcDOKaSDVCPbn20Sjghn8/YIO9
U/wcQjCWuDPPXHaEDB+qWOk635cAR4BUNVQ9DPZZxqboVnI/lJ8XkPM1yK9YHxda
ApBlrQvMB3P71QrT8n5HfLAAfCriRN6FxJEKmvEylbsKY6Q6EJG2Ar3qihQCoiku
Wob0KIZZb3l1hhS8U0Pb5RETV2ODTICjcdZKf2FhmFK78ynWZQbUV4IeM3rpseCf
m1xgWf+ulK3RW+BvEInEYD3aMLQokEABQtzgvxxrCOhQRQzeLcZqgLMgNzdPNBwL
ObFr/69HCkAJclV9E+busVvAkFFVpHIJ93kBciPwQLfrVZhveJEHrI6pRE6RV2xL
yAUNASLi7y9cmfAKcncaezy5tJb2u6mYUyNdzswnXSKddKIFU4gp+tH7v9JNab5t
fG7mqaDEan0ggGIBvfRNUhZe1hKp7mLuhWULp4DkH27Njwa5RGL6/yI0AYm0TVIk
VJcGSAXLqjgCh8oN/Wv/5whzS/at5FMjvKzIes2VABAjZAKwpF26GXM+4n8qAyPj
h86kVqLRBUmYw0r75oSAzMWIkyGClBD0TCYb7DhaVxVaU2pJbmQdN5O+3crhbtnZ
vEnb6PT0KqAo/S9SN1eMriI2tJPEw1YaSYK/gY2kNAnaNe8ADV8ysgxx/Pm1knmX
/oEG+StaklwvN6WJXl7PPf5J/c8Dio7/ddc549NJtCzq3cSSS/l7KoZ33gddf9be
YsfrCxTllGvXtGQSxyWZlpviTUs1m7Sayx/h92Xuo9LYOwlVROpB38E0fRr/jvWT
6RyiGxY/PTjiLWZLCDIUOtV0V287zT0cbf+cf8RlI5EK6CxmrnJFS+txPouqdhXV
Aft9dL3U+v9vS95lq9tGUnul4XXEiMDJ2KJl+OfB+oVBR7mGsYDq7uBYMMVZcCHE
JSUGZDjFuWshWf/v9Qu4WQQ3lyMkJktN9wEoxQUo0XWTc/OmocmUIdx1pmdDluhx
fub1rCdcKFTPS3dRhU62a2lS2JaVsZNdlskma/Di9/b+xrpQCqb0teKfw1Cf19hQ
jO07COTVqJJXLGE4s3EOYLsyUz5Boq/lDvb9JVUMoQsGwztryi89ueyeIPw31poq
AqHe3MJ7kXR0k8CTw7FqjhmHvN9zhpNSv+SG0qg5jsZ8cnQwHM+kyI2ohZSpdwqm
1ruZyyCiKZKkG4A4p04q3OGAmJgegdpAEz6/9+w5hoMBhYdECeF3R5o/tOT4rxoo
qk7Jy4XbNpbh5Qh2Ho5ZRdLs5d02p6kILuJfrx5SsUCjlTGwz6QIvm/UHf5VLM9L
1+o8d2UKOlcsCAI0pdXcQBb9ZJ1swMC/SXlMXQGXpgtIog/khtnCcgJndMVB2atF
fg58iQj3aRFGYX1DDMrmo+OzAo9VNW8fok93boJlSAd/IJMctMqvBCzi0UILk1vg
sAn91Jv6rl+HsjrV4o/cjO6ypYLOe56uZ8CxrFuM5xy5t6/wXO2vdGmTkD1T0YkO
6FEv67AyGIWH7bwdL+3gulv/iRzCfbyJNA+UViAfHkoMU0jyQ6RwxG5CKIwNOcSU
nDlkpwTy/xNSzCURyTbkwMNFST+sDklfBxoAEvbTqs3gXMamxmFG6ETX+htCZIoc
AkYEQGDfckutk62lwIssPrBmcF3H2/+bniqzGSLpQ7lezhdIjPNJfDU1AR0I51t7
NXutKxB9naiRIAjCtB5dnpDGJJIT5E+GbISmSFWg1mB7cuyYv1TykDHk3FnvHElh
oOHCOBX/NiZmmpRDsuR87WFHXBUnSFyq3IIxFv8i8Qwhk34gquHLVL1OhsQTuGtI
0NXwn6B/hg+SEqZS59LnBfvXlB4Y194EaXqkbeMqwUNDNd1yhH9Frxo/ddEgNDM9
K8UBsCPEPA49PsR6P+/fAfw+eF4wVBHCVyzZq8K8zoG6g3sfSDDeZQNlJawp64ER
pRwcCPGfRN885Ff7UR0k7ZIoJqKeQtwFwHYX1r09OZU9bXy27Hff58PDmnIENE/j
DRpJngRakHZENXQhVN03ryJBpgQupiooSZm2LEneYl9E1dR9RiamcFzqe/h78xBv
flbm2PUtkekXGVxFaJiExtRAqIO8qswaMqJQNfeD2SzWwKeL0HLwmO3XtF7OGVfD
DPBOthsUjcLGxx9QyC39Njpfw+uETwABOy0iJa3GMmbBnE6ar6h39NfivOHkKXmM
9uu61lAZPZ4I0KhXViljTTZWMBmH2+L4t+1WMgz96Wp31txBF3ztUyQbfq3HqYdL
/Ms7+RX3MPW4f+LZzxouX9fRh8voTFZLYCUxj7ART4M1/NEl4CnhhlUOGPfcX+L7
JDTWLJt0XEztNjNuV03syHWUdZ7PH2ql0W8gxBQ+SeNrkCSOq1zoaZkIeOsFcGnA
MHaukYpiB/8gxQFCRGoyTyFE6taQovyer9vKAWmFp0osO9vNJEI4hTeCqZO/s7lL
FAecD8yrwdXd1oXLN0nId1yh7KrSkZjyPpF7OYL+9JeWMQweeu1dnh6Du8PMpjbf
tFWXW6wjkT3u68p0mmeAZzS5CNHFMKeptroJBx5I9aPlX7tfAW5+Ax+1eApzAmGM
DnlHYg2cOgIDxg2mbRnlt6rqEFI9avvWLoHgiWd8c4d7lDncxzB3yBxGEQTCZ+gB
o9yOP/S1AI4LEBOipHAgYedBlgYzBySeK9mbeyKyZTACk1tvWUFYgzPFxelb4KgA
ryoJPl01RJHLMNszMJH8ifukTV8Tuw1Kls0agp0Q0ZH6/KK5NxcJKScGX13X4NbF
x2H8JPgOP7OX7aDTXUsP2ZLmE7fvgat7z+szhpTD2H13M6Wqx7N/Q0zu8Iuw7H/3
32ldQN+M4ZjpIshMWnM3xa8Lni7Q/zgn4FeHvMoMfGkvN9LWryf8stQlPSZcW5OG
zqZLgRgQLZB6gnQQ5UiL7LkDP0H0L5Ar59KY0YtYHrthHS+kL3sCm0i87cAkly5F
cnO+cQDDPeyqUvpaiScL2c2/BrWalzDj0RS4YblJMsAMkkzlfoAP9Qj9Mt7WX6u1
dFS70VswYhpKLSNGBo1Un8Ltvbp6q6a4ycqiU8fPM4hiCXYhVQWwwSQrlkXLKJA3
23k3MCyOIabOb4dS8VbRqmWwOC+3kZTf8XLbNFBKfXOMR6C3CjsaxSYurzoXfPU/
naRlwppHDLtp+0owiNJWRGURtXWCaYZ8pCeTxHuF04IaKVkjPxV9U4t/NCJJtCGF
jPiEqwTDvoFoQTRXhtB2sYv2ZvpuK7r/wGv/DxbHcnLd13anyGkb6POuBIKZle5Z
mFn5UyN+IVyXXNv9gzAAqKMxA78dwPUHm1VTs1QdCT6bOCpqd6JCS65AOcKgzm4g
Csc1vk/ieUK6N7/Vg+KyvZm7DVTwLvjYU+iOOyhIhpQQfpGhPXcpB1v79ZquYK4+
V4IF/zNWjg55B2qKAbwsbnYj+cBCi+W27mW1imS4ect8ltwj51s8yLyp/xsO+lAI
9cgH5M2f78Y4SNf47m/ZUT18xhkBA0cOmJI9ejh0gYy9qAp3x0ahlX9JmtY3bI6t
BdjyTArqySqJY2JD1pxUZuJovPn1OJj9dR0cgHrUHXcwyTmF4cw3YXBMBSXJTgOX
D80UmDwDeHgulyHe6aDdFCE0ZzOOhtNJx+uMTfzOhf/8Mel0yEuoaAcECOi8uYjG
VFSCEl3Bh9MuHWdoa9GI/K81Yvx6mwxEeVuc2H+39lhH1DuBKPw7qxShonVwkazc
93wqN+/OkpKsZxdGbG+ZqLdCWfbwX7IB/B1eVoEguh6cz9d7HuUyf+gedu4Cm9rR
MveDxTiS1LyNwllzXyXQFXTtGiLv1SaGtTyp856dDMwH2Nz/+Wk4ydkFLhw2WDSy
MPP3csvnPo2cYplUWU+FRE2RgXV1BV2pLyuKXrCkejY+ph+muxNzvqsHIOiFFOOB
hzCGTjZLU0y4BSYiMKhigeAOTMD9aqcaZ9iXMUxLdfIXV6Jd77Bb3HvL35PsLQT5
2qIHbQt1PowPKy/0K3vursxFWFIpl5MTeaQSyJq5vOraMLQQGmagtj7p2Dpghv61
4lowSY3fnjvTmMPIK+HnH+nkStkiXaYYWFvtkJdyoCqoykAdNRUpXco7F/S0V+pV
ZggQDqLtulVwG0rI1Nh+covzvs+rpaavCONDBhv/81fo+hbA5gUZ5/5vr5fhkw49
m53m7HsPGuiWvT7ucqt66dDpocp5ToXFkuZueA324LfFqjsx1iR/baHPiwfnzE1A
g0RkqNw8W3AYCDNVGBkTVW393bbJ3qwWVKfFxy2HwgSewMmTX7KWlD8lfdcLADty
/49XGvCFQFE8Kr3L1COFNOuyhwivf1Z2eER0wtHsfuBcDOOpjoR5u9OlvSGxpTXY
7cZAZyS4FIiK6c0Ec+B9X6tCUl4I4TXKiVPWykUy3aZ3KyeT88+yRBuTbtVG+EHg
QtyJNoEZgDBFB/F35hqKkb9wNZEVqr8+fIYMmywchxt48h7lbnFYXOM3TqG7nAfN
4c3yWQL2crkfhsCiOJ6IEe0dm2T3QTOTg14OJlI5DjLCR2ce+JfqawNcLt2FidVb
rGNOqyjw1/Mbo35j9tdUcps9l9gyloYg0BdTE+iul46eYtiiIuRzDw+29e41zaHK
NGLv0xeFBIKuLSm8kliVWhUosiooDRc9yK4A63f/NoPqCJlo4unKr5nzxkd+u70r
upztYYB6d8TsLnWiWXXYJEmTXTTOptfiibovPxg9Yw8qbpttr41RS33ZLxYsY3hc
2W7Ez++POhjZxDcfm43PgI1P28FRwi0QPTPyfIxnpEyc36H2bO3OXgK5KBbXscvm
IC3pKLXTXJfO0wk1Amn/OTPZRYL2xOayPLP9V0yvyHufwJLyQ0DWASCJkgtGr4V6
sJR4rjFirhOlmdJeAu9CryGTVhTOUoYUco/BB0sAvM0bS5FuQMosoT+Vj9+NqRv0
MgdssA45z+m7QIvIKLgWYffcDWQ41gscxIBkkiTqupS4SiAC7lAs8NDFYHDkkgZU
hYr+eAVeZ9B5a1bZZzM7/kV/YZjDc3HEJoRBI+iiRy9NC6SRI3A/UD/xBvoTPzZF
oF3Th2m6luN5kgMEFf4NIGxBJT1iUpH7rsL0aOd+qEGpu6yjMEZhUDj0vV4+x/pp
hRKvxVGxpbeN4pi2R4cFCmThbEOaTF2ptCT+tbxig0RpIC27y/CqzBHR5YOJuz38
8x0rFaIoiwGhXc7FjC/Zu1qaKu41h+UDfXylmiAJLD/tQl0RBt/2YJlObYeBTQ7W
lU5wpO5p0F0WWFfrKyx9MvFpKcLnHCjdkpwT+WRhj2/5miRLY22p/0SqFwjBcjth
/X1w9l/acSnyZP7gEyvJjJ67ppxZ7if2r8xuUmmINbLPbXwsopI/yDaLpiV4t14i
XTY9smsevxuDYCk7KnyhN0jhQaL7begsy9ry1MvHAnvlohzsL7WU4nxZE/FXe6BV
UYmV2tz9Bdgaw3AdcLb2YMRoNGRZXCP4fX0Ah9rbaXXG8gg0t7SYxZOQEIqEC22e
Aihw0wB0SLVBU4DJJBP9hasWYK05zr244y+DIdxxPH9M78kwWJc6S3c8XN9I4at7
HWwISzDSKqI266cMX4EEHGGSmdBmcAe5hnSCnuj/rZEMavwTAAIGLu33uLpFP2nx
FnZMp/SZ63P9RrMhAx4mzQtJyFRHaXj8JQ3vmtx3RctX1LVh052r2LMLOYzkTIt+
Ghl6/pxgfQXmWqLBfsB3ra6uEjM0Ab+qt+DENWM9wH8bQMeTQ1yyibJt8tDTMmei
Fpq/eRhrdTgocB6Vm4QIGYxbMup8iZWzrmhXT8/qJUTVaDtD/poc8Ih6I/zUdgbA
+bKvw6pGDy/mIFfxz8cB0dd3DMUF/I+FjrI8hfvujkoKDyCCsOmepdb+q3CRrMnm
95yYCb3BrPvrVAg4GOTPbAi+iKYECq7Fxdn9ScQj91z2X9IDPkbriRZT6NtLVdvF
xoJBgg05u2LHPTqbMtvzhPVMLJJmR6DTkKOtRme+bH4JaVFh25TlxQOX2rE3jvJx
5zG5oR8CrWA0mjmVvjk2yBKVYGUmcQ2+xRMyDiO2oXfLmiZFPkXzMRAlV40Gg5KA
NMoPxTuRm3HGGhfDGLUgw/Oop2rfdHkgEyEadT0wIKo/8PG4N83ULar7b948tpKH
XUij1CYs1tYO3UT1qn78Z3Cw8CKYOlXLvjNbDmRE64JwulR2BzsXVHAj7cPl0B0O
C1NoXsSrNGAQ66bTZ/E5h7MvsNU5058Vo5wMjEEAYCaV1CWsl4xh1KlelfWErrXf
vjlX+gkBnKvrwBVKiqJrUt/B2LChOB/0Puoe+aswxqvv5yorfNVorwhfoBGgBhxA
mlZBzj24vDN5OPgExEkpAg0XZlDpW8WNflbPWsEkiwcVKUN+UGxEJQqKDIZAEpBE
KU7EPMK5cLqfBq2m3JjJ5dQwSj7X9i2tH1a/WgJQi1nlkm8S6uHrB7Tn5pK4eHb6
XcoDUzHmg4Lb+hW2Q/tHHZYm3opL6eP87Y2UA/R9DRGpY0bdRdennHeenMVWlYl1
fc69YffU9mn8N3KHcQVwlm94eQi5BKDBchavhz7kj+TZtGotn/kaaxfIB7B+slIj
JjVChwWh4V1SjfQMIcSIV5z3cezPRLjONTZVLhYOHuIxhZY4gAvW56CXxw1WTtER
gzpgR3sedN2pJIHgVZpg++fMXXCYODKY9n3BKM55lXPjOKEvR/matQc9/8sKpIm/
JIM4bqrHWwMgF0t+tOOE43+bdsvQxAvCP5jE5plBxnx9LtauLd1E3wLN49z9/Bgu
JcQurgQv9tuyBI+UB+3J/STPHiFXTcYh7LIeKEld+/TDi64N69iw99yZjDLGknLt
k0ybC74Xv13jePdA7SHDhLKlSWbnLwgayforkop5R7z6KHcEyiJCLFklSRpocZ+4
0W5dtoTiUPg/GZkiGadqbK8baiAiskG1BQCf2R6pJ7EV6D6aheVajZ5tw2zCluve
+nmg6Sf73EfOuIZTCK6gkSf/j/V0rFxMGXhhc940q2p0nhiUXwIxKjXXfuzHw+2T
USRdE1mmAWOBS+Ps5VQOrKx6/aBb06f8ZcVBRKj6HuI4xZ6c6CP/aBlb8Lx4+vaq
bBjQoYH80A4lb7CAacvJkSMcylmvcoe4yYBcRIMHywl+tQuCEp9SnKM5LjJpwpsF
13inKrJ7W9yVRlnEPls4Yi5CJEc8NxA9l75WLWcCfvXAYJIIR9CEbkSO/UQew4P7
O7nqc3Gf8HYtT8lEchV5O3/TTJCorowxyIngRilX2PFwznCESg2cejTs7lIkGUzk
70Yux+kw0BqpmMSmgUJBR73o4xcdYWMeJEqipuQuqP/y5m1rj3xNarPYA5Zrf2+l
CppRbFVqcBeuyEUhOtRGNrmTcCuwqwXw+NH/1BSN0bxLMcuckPkkIUP6ZERvGq+h
kKR84oegWHLnrcVfpXpNtx2iw3CJ23LevvyLT82FnLgA3q3vnOcsg49EjnQERBp1
tdkkjc/DG1LCpMTpVFQZvmKAGJ6hvBI5bbhfadcoSWNKUYljIF3s6K3JvqvkfRa2
6XtYXqxGPk7NhDmbA7hBeX6mZt6ANARprfvADlwKKoPZKOMiwv3rhf2FATLGhJBQ
/Pifk++41LQykyVK/md4o78mcHNvQKkCBwSBmgU85ZZ5PLwWO7SHy21jIQzhrLow
lRGbEUSXNpg+JHxOLxHqT1rimkZwnhuzcfrLbMag1pj0y5ROS+Y19Fxq9MEvGvty
v9qPCadnAym8jrmqxfjFe3f1/XoVW5+6zYepe6rLqmAKLQET5NIttt8+dRcO7Kq+
CsDdHMcqDMleM0QyWTlRL3XIYA4yAWVCCK+aOwdIC5Xr4v58O7UxaObXphwHINV8
z4V+OHoSdaTc4qtB5j/ir2BE3Ak1P7wANNxlhvDtwmE/LGtI1moqIjKJrru0MRWg
r8UdNvMR6ryz7Xr3eddN00foBSexDIo7Or675Pot9PZsAAoEIZz3XUhvqqHJZ1bB
bE8yvsYumnmqIT5SdIMw0eICDjTcB4b5cdlf5uV6WgLj84ldmrvTX+/5S9RY8rqk
rx/BMyn9VGFn1Vsn2poDzMJNx7fzeKOzPuZin3DRPTwQEqfly8jg6k0yFaYtJltt
wmE455A4zrsOFCnGCJ2LHFnHgptQlB8mKPto/I+W1UUhKIvvwumscr0c3odYLP7F
uFhF9EFo7YrjKa/wKAAdtl3pDAoybs+6kzzt2wMvR5OQ5thXN16sioGSX1KT2VM0
2OtWgZmKpc56fzJa6vBITPaq1rMXUlWthll6QHsq0I8GESNYJr7+RAYtvfDJT9Xn
e/CUZg/4+p203Pnm9zo9rixBVrkid0EZyDtW1843iad/N5mtm9yBtYMk1XIUfREj
27OD5B64eZwc0CsBKT5rdA5rLDhHEx8E/lERYdAwgMEiCh2/yulTfHNzOjBR4MdK
5zL9YZ5WDRgbwtq5j5jqYsTM0+4qO8c4EYYcKfR/KYWnSk4jdrfu4a6gYE8QwKlN
2QvtLW0vLrhJDS9lc79nP8VEKYyIzZuRlonwbKMqYDDlsfHZtYlcB5q0jAHHPrYO
70ZPt5HSpKsemeWg0K5mVQP5wOhrPRRm6TxyIPrUHfzU8l/awWqPPjBLJJmK0T5l
WIxapBpmQfkdWl7KrAoqVzU6yoS5Y/s9nAjTNZDAChxxRxOE/RsaWjPbR9PgfIJr
lD+ndPOH/8gtoYcKIZzA6WEO+dJQBd+74C0nHiAu8C/nPROzEpxzZkcw+Dc6FbI4
bZjNZlhamvibsCsCLHxA4rw0n1P0jU+GC//vgm06kLcH+EqLWS3oPoDsQq+wAlu3
ybtW8nDntaPS86odN99DptsdW57b1ehI8GX1QG3KA9lpnWwqGbxNZFeVaYqw/hhL
Y+w+E94eVwmoq9WOl7Itv2GQHkYaf/fWPCSD4Ax5G5vTpSf7X5l0A5v8VoawDaae
1I0iFqdnTLuIDsXeyzD9TniQvREB2z0tqGaE6S/gKbSqv92jDoS9YqcIKJuLo4yH
4up9R4LEvlbUXLGE+3duR7g0ds8+HJ0oDxQ15xpswgqQmaMsqrVlLfG7GCaewq4I
w/bW6cs+tTcx5Ur6v660cPqCOC9zdL315wLVruRIC2ODsftQ/YXsSBzYrL6MS0WQ
5Ax8JsDXqzrXzY9sZ6mWQ1b9u7QT/1LxQ9U8Oyef8glSr/FMhz6/1+tqoWl5oESk
0v5521ZOQYQWK43iChUx/lUan9xYYMdQbjuLeXMIdUVuDD4xCpEQmFQU95pEZOYi
9uTVcmmod+nmvTnoDsKKX4T2fFt2Pb9GBbLWdF6Ej6yV7+vz4IjQyFg24Gak67Gf
KZnaS59mYS9SivtkhzmwrpgVRUl1YlllNDSr8cceQUWTlh8FiqAFPuhQjk1gES6Q
l+LORhrgzGfkmXJJUkKJocwsXGPqo/kispKRfoXL8g9f6XLoz8eIWb6f5vk2I7w8
/eod5/3A/dl+O3UTdN+akY+yBrBW73t3WnuQlxJAn67ZWpnPZY1WRLb3rMK3U1l3
O1wO+mQYKp2FMzMVxVe58fCSf3ZOwTQALBS5m0jSQxOERc28EMrCnO+is0cqCdE2
Vpvbdr2c/F5T6bd8UgmZ94s7RlTqO/IX6btBKvXeA+2O4ZvyANSlqFecjQ1qPlgy
ieyTUgBhCQ6wD+9wrYeHsl2nU1cG1ry+PHHGJIXxQlWfOQn8OR/sPlTpibMAMG8S
szSrSOxuWCOrlwF+0wd8i/xMOeGMs1F1EgiTcb1DQd8M3YZDUU428RDAp5cKpr+G
uUBGeylTCQO9A6XJGnMP1OaXSRgzW/pY1buJqNDIGBHq5HN2eUx6twabzNQSC9BY
VvgO1YnIpS7/F/Zgr4RTs/2WiP9TW9N2J7lyuBo0Br1VwxrAiM/f7W9Ihcq/BOrg
Ru66gCIqjM9J9/ZrQAwo5dI+mpZS3piEjBY0tbCFX8tydL3O4r6UCn96419IN3OD
AAXfipUFULEfoqPuG1BntPZwGXD9QB2TvEvt3hfpIONrSqmgZ+8ZynQJd6JxTdB+
bPTSLZ4iJPohJOyGR3IYHLnty8oAGV6/w/8V7GIuY9e3r6WdcXCmQldEzb9548gj
Rq2gASmebjEoR6PKkEmy7FZlufMniwgiIvPHZHY6+ZuYGFJ+D9AuVIzv2aU0rYBY
ptpQoO9gKUPAZXW/F8PSAAlT2i4I52kbQuthxpqt0sTXP2tY517ymPT4jEWnK2lo
SeVC5v4+Nzom7qNHLVmhxs0toJ2RwEPruMPzUa6/hgTAfEU7cepgVoOUSXbUhGYp
FcaUGefUhmFSmzl/ArFocRhyBQiTZO0rk6X8koL99SFrWHKgZuXcXw+/k1fnbHd4
7GaostmDSeWn4Omp8wfMumBZOIuY+zP7uXIaJjcWzk5Ghp6E/YV1E0+kT6DAMmbs
Rn6omYSw8XIleU94GYHibmr7lxrOWr5MG6PJdvRUK+Vg9fK7VKfJEOPTOifraqBQ
iHLOkVwf016d898q67YHM6wcEIgVMW2wfeOnsIk3DjB7HdLHurgyaBJlnPu8Z8K4
z1il4Psu3caW9/i//eWwIiJPd5PKCstEB3j3DceCKNuqEKZP+eTotXMxTfRtKSKc
WVgMkRKd7Nw2okYyoaJoc33Ni3bomJqlQIUPwbcDEZoUINP6dEqyfNGPQ8Y3iQ3d
gECIDcnaY6OoJ+jpn0X7evmYRqG/naF3GP3gHP2JFVzigIpFPUB5gdoZ1W8oSS5V
BXBnjSppvLVMdaWuJGGTFectgtd5CmF/XvXqXPzvkoiav/2BZgxws6g8ACY1nlkx
caYIb3ABryOC8Vu/YbNiCdQH0pfQvDNO1ol4nLjNoPzAFEUtDxj+RUYXVlYO8j5Y
h0kj36pZJgig/u/YVXjDtrC1s+lRz2NcozKl64FYmBbg0knaXfBMrwtuX8UMNXuX
4hRJ1IkAjSh+VxLNF47Xk45W3RmCNuh4XhHqutpiEVjNoDBXYc2H2BrQeiElHoxR
7tiDMeFFNSotz5M8d5q2tbcxxvHuE22WLCAOeXIokZDGIU58TrZiGkOYszYFXg6m
2fEt1ORwMxD75WSsD/6EJy+Mme0iWptnoENiRJWSIjuwi4iij9v5rolbVMtto0i/
ViBK/7d/ede4WU9K2QpJ1oFQo0XmpX4u4czna353nQ/5R/F1lH4+Mg8TiKhlf/pV
iEjU8cgxXIDp1hc0Mxiey+V4NsRV/nxLJxLhOEZqNOInXDyMWJhkq5+0wCdIgOgI
SoZtakaXAvdk0JMDvLY8+MN3sHX3lq0vPOJYhrXeFzKY3qajrvyeHYxe9g08dbzD
LePHI2t+B77T0yuG7VGY30xkAQLZGm5Bef2kkDtF21enoTq3aUc2Fu7MUhRaTT6r
VGStyY6HMxwtSSvyPZ9Xz/eNduyCkMJbHAORDQ8CCSIyBeK4TuZ80tc/PZEZ5YlZ
KynnA9McIDfye2Qy5zlekGzypXM6JP+RoSJ7kw8XpBn1tWesva3it7ToGKuLEkZ1
N7LIs64slcl57VfdqQSB6nYw8eLcCPC2RZlA3j81EPxv8hnqF9IFUGeMv01lIlgf
bEcIMMyo1NK0s+DTb1mt8ps3e1CT4eS9Nas7VyPT3sN5sXRYwjhwjV9pCoEdnBJI
H9pjHZSkr/OuoF7fIEiE6h4ES3oMsEs37WP7mufKgp/g6wAqouvZKVRuWyHL/Nrn
SxEHU/FmKUIS1vq9qZCz63dGhJ9tp1l06+ucWUeA/sLhUeuBVidAV0hPUGj/crOY
q4M2wjbcHY02R35iC8ZPUWRvHTjn4Ccd1bbmw0mw6v9jcUS00P2naulNrBCZb1+m
dwI8LFJmQYkUKSVEZdVskrCmqs2HEO3AiwkRcI3YeNP1+7oxtkf8xsXTmsFRFxTv
d/HkijWMbEUCeLLw2HuUE6sgTc0ABvD17Q03v3RM254pN/Qqf3M03mLEBvoT7j0E
DjcSUm/bTzSN0+9nywJMhdhxnaKTma9PnEgtDeN8g2VKS6ujCWOSryhwJ741r9WQ
WRIwyId9CFl33CLNoRHt9ASYbTGA450NbRQ9K4UUuMHiczwhXcd4as+Arksy47Vw
XU6PtAiktnNpBQQJ8bkWwyr8f7SirJWWFYnz/PWIqLX1rQkrDpANNpwnpEMGMRm0
Gb08CFInvYDVV6xVhFIDPtaOYibXKKTa0osRHa0N4Nj5jpkkcSiQM9zb41RLlxjJ
BGc4o4PfH5qYeIKP/s5i1VgTM1hwqGYCyWK4fkb7KxaXVOWh+b0wctTBTP6SquwA
Wnnf95xUsUOteckf1Gp+qWJJZuUUd8PZQ/YZStMMJx4zmQ8aaYVcC1XfEktxVLrH
M7V3+B3LHPGtJNvW6ia/MdWm3L9jkg16JQFJeGb3XEczRejEEoZodS0iAZtnhniH
ntqPbpPbRwc5o3fg5dW5dIV/fLaqrnyLNeFUkJDpeqUHea3a5FSpds0PnNqoHG+w
stGw5N/F1aaOdkCe2uU4S6Bat+VWktZgKIKdAHQG9A2/pYom1CqPpaMkqacO/9vb
l4GDfpkvqWIa96uupexnyaGg6xtXSZ2lgCig9pd3QG3/Cw8XoI87E+KEp3QRplSH
jCzMdy8KxBeQ6r3Z45v8d7rxLDBcPhR5XOpP74yUqPBBRP9ryMN4SJa9SpJH0xx8
grYeCnZduZDoaA393DbgPQKe8c//J0+7QcHKuDoQvC666D3JMf0qsKbFUq4AOI5I
KqpXjPdaa2orIBoCCVL4HvJXNlZNmgG9uziTegfSlDYZMOmhghpijJiaXYaU1HJu
nyXmc0ksoIKehjWVJ5qlHKqLulXpe7hscAYtfuiCMcsEk88HyFr3ormqe0aM7TMl
AmVfW9BEEOmopvsVmtodAbeCWXlynXpyIr/mePabmxylj+5SoOa6jrMpzd7aXTIP
G4VK0l13ka6nyS/r0zewSE833NT/X45R4loVSW60Mhblmr1slOg3MW/8IYgdUcqp
JS9fIXZkqdlSe1Yntnb86qid7zGcGFjIbPW4asMly8bkS+CLREgUfyB+Gkc6zOtz
SGhPvXL3FtzbkCZdcdU0rTFdMfA47h+205k2SeVnoMoMKY7E2O07E4GNyNvnu3tB
KoXcOFn9ZypciNNOLVZv5RB7G/dffvofXK/LMIl/dMygVbj/9sq9jkIa9kqbJ21i
kfr7L1PrO9bM3HrmTUdhl2AAapU4AYCL2lBJOQ1/gButFwtQrexFOhu2I5n27pbY
5Bi6n0NzpH9u5ky9GlfXO+CiZ9vAteS3HvRnXYrlbRtSA6xrATDW2cE9GszM6oeE
KfnSmH/5Dg94DV4LTkfSTGwDlLhTolzg69Od9LaQazoUpzsU2GR2HNVHPIu/PiEf
199Ledj9clHHlqID7YJXp84JO39K5tJg4Sl/3joBu41laK1wXSn7qnrNeBA8TXbh
fsvGSngBd7dDZKP3zjXkHKQ4HORZlvA6ZzQWBvE25oqsX2xWNvmCa6sdGy32jQmC
Ugw5HkngHHTjFqFawYFI7wRisdMZClC1ipxblmE+JHfnTsrDi6RywgryZN5Eh6Kr
VfaSqcBlA3fgzy0hEa5yE/XqQ3fZbhKShRVLBKX+I62r3FmoMCo1lhn0onUCkex5
TqUj7r4RqV+sYiZ3QrL3ZN7xoEmgtxnHX9AhePIAq45lZm5SLYtds0Y1PFnNYu1s
nAAiCtwlwxCkhX8FaDRm3KZXXSbO8DezYgcK74sZO5Oc0y3MJGjtbij8G8XBJzGp
MHitPWid25mhQXg3VMPvAlc08RPT7DtLSguvvYUdB7y2DohYK1EzRnIf8HegTi8I
VTdO40ctF7qIgRXyiRy4KfnOVA7x+SeEPcu5Ge1Jf3jeT4yPkb9jrNkkejysoiM3
fUvEmCVt/WJ8pe8Fj6m8B/zF9sIuJxVjpG0473Xdmy7ZS+lL3j+a9ZjqlvVf5VbT
leyzrlPkAIXvu09jy+OtOrwICEha0T8Hn8nLD0P+5i2M2NVQwY2kAI5a7yXS0sCc
XnqVKgbNymAWC3Zcrc2KDsWbjsexDbS5dibD+v7cpXqJbGYtQm4/iw94pYnS3nGO
jt9RXRjq8O8o9Iw1kMdhFAQ7a3TeDculAevezlN9dVOQorj3dbvPvGLOVEPGjS1r
rbSPNzZhvYl+9IMGZRR1lbthKZ37xZj4BEFFuwYXO2U7L5fYCKnaC9EC35tAsfAV
0Etu9tv0GLwJ832yuLviK07y7xRI8NDcr/TK9DW1ifMn/iuXVsSG0szjenOZPa2q
V41gbT5i+tvGbHFo6/Itfm2KIlhRbEfm+tzhjzwtfIZwklcWwHt2vnLsEIBhqJpo
rVwsWPCAcyNgeCEc0OXnWZ5A/RSjr7cKhlDwenXYQiQF5az2gQBhkP2d0QbDqK5j
+dHdlz6J+wqlDjpTgWwecwZWhOaWmxaLwgzu5VJm4FnO2L/9HIhp3uUeCYYggOHA
Hhdx92kYvQJ40V8k32xhFX/ySpv+rjGByjI5IbNi5s2zU/jPz0IBCt1Unj8B20wU
b13R0Fe6k8QsHYx7lLSEm1OBg3kykzRmsANIQLBY7J3oybNyY2vbxH5PtqLynraG
mDoP14lGdwUZ4NhjbiAc46ySRvDrBZKGx5T5HugkfsbhXpnLmNmjY1rZmeFfyTfT
jKyFNzJvdYqoelxuaghvXirBvRgaD9MzskVohjRpc+T3sFFOOPZrsSKVS8U+GnG2
9f79FNqz60O9SeEJ7WcWI50LRZfvETuSn6EPlDisCuaKusKaIqLMH4YMUivz+TpK
fGPaS5bSUab3tERni1FcHw0A35XkFLnUCxHkkHmK6jWEEANz4WbFTcbrEOxyl8xY
5N8oOcpBXtKcFIpCQ3i+s4cCEjjcVV0pgzRFnN9LAUU+krpay9xW4PKNyMt5FdTF
P0VC1R8UPrd9vsXvADoQKe1WETcimCcngtLwmixblEsnREPeRMbNObl8Y4wdN1bC
HieiJ++Bfv5Cwnva5NAFJ+7ae59DwRqC3iuyENF1PE2z6Y0e+GZpCylbLPy5Hxzm
kHmkK0LvxEbjjOsAedQY1tZAiP+8+ZzNStWvlnqEWMBD2V88LoorkIhHvQJZITzB
cX3sXrBO75HMQhViZOgoxIXE/rp6yVhcnBO65t9EZE13Bdz8KyEeHqrTo/Xpuv8x
MXdnfm48NTHiG3YQzDkwfInfBXBbglWlh9GF2Pan+baPx6Aqmd7yKPgAJOOrJICp
kiwuRTPftMQFBFtiNRrceywi64BMgtUF8tVbfB6MOmMEKLexdmBlBpdbCQ2EXBx+
zSgBN+jyE1xrRmL3XmqZYbJhby7S0fAQ1zUNtUYFPKGlESnNPmUSha00UcgDjRah
70KYO79dL73GKAdndfvVSMnQyb6FW7kK4WrycPd6+J/5Nam1SGUE8C+vNWpjt0Q+
ewG0fdpy7Oi3nynB48rfz5ECd3xEa0hVmyVS6+a2uuy6hr9kxQhN4leeDHT8m3U+
ID10Q6OEnUZSKQZPB0RWvyD4FTOprTWtAO6cQ+rWsnFYt11Ijpjw2pTmuoXbpS6b
4KHZWGllhDIK/2dJbldlfBLeXar4/mFK1y3JTFAKIsZdlDTY2qIyPZg+pL3z4RUp
aT8rGuPsMZvHOmcfRK63xm0xr7emgz7BZ8sZCCLKs9pGgBVNcKKqn+YU7A2e16gb
UxZPbvdJlOXGnH3bwnQkgyTw1+el8NIARt9ltzmUaDCbIU5a8okTxOoT75aCDy5b
KgVMgy3IKq8JyHQIjjhFy4xptTFpQHhszxFTGiUazgnCf2GsLbSD84Y615Kff+j8
cqk6coUp8AuBEUXDDxwUzvzDDm9RG/VcRLbl1WC6UsOG2bgGuo3Ny/7MvUqINBYR
nI97r8WseBHHKXohb/aHu/Ehluvx6ClIr4CySFCSVN4aHMcZuPSpUWLBgTcoDYza
vFRzSrK1E7vgPtL5vXvYR18xirNeaJx2LnBgT5ZAqZrTj7RXEV2Cy9VFkiDIQOOp
+la1mB8kuwK58UDkRGigXC8eWnkmEErirh3XEbcJyFLGZ702VLJ/nJAIQCgStRm7
YLwGs3DHyw8cSb36Sfymxg0uGgXsqN07WbGHZlfgVLP7YRW07q8iShx3F0iuVqrG
tMwg8Zts5XcuUaHL6NnPwcPd1VJC2olIGSnZi5yOQTwZgtOR+C0V/DfgteBaZ6Sq
M/ZDpTdaK4yVLJ6dEeuPTWslIQj+6QT5YNjqoN9A/oJvl1Hhmsw2RpWxo1X0oU4z
N6uepyPQl14PDMxAfiCivhCkecVtEXFo+zS3FdWBN/tjU52Gm/CETkWQlXhvzR2A
QFEEhwAtLYnbinF+5DDAEV4i9dYeYZXoRzTOvkl+aJPgb4RXNUPy7JJ8vqEnuo1Z
dLmiH8XNCq1+BWNW7PrkIRMDCZLxGTC4szUWJ1dGuP2KakZ1K/9jgiIKDjDPqH/d
kjgxJZcQD2QSqXgRujPZtX9YdzQcgki6o22ep5BIcU0Do0wrLjAj8TFDSM4BdqLx
/NCaahw4dhAdeYbPGvzgZ8hc8pXicZYFHHY3LoW1zRKGa8crcEMouSgM5LXRZBcK
QkWUMPPuii/n8WWYxtteDOiBcy2kDk3HFohaeEmcO7MOG9tD2MV/j4Rw47K8rpmN
KeOnqZs8wEHhq1Kz5/YLeH+IHrP8BAaU+XzM0sT2unzEdtvJJmKANx2iSZXxDznQ
QGvZmecBYbeGWe9LP/UIabk3UCKB1YvvTqCu0Q0Dym5xsWRl0JnZX6B3oVBiiiJV
dRg3CgxHt4Y4cGaHWz66aI8Fu2siqsC4sVlGKTPRWnZvTEXWqqA9FP+b6I/lagek
wdCB3aU1gfptIAQVSfcEjJrwUXM25s2AggoX1RdzfYZsqfm8qE2WYR8eu9X3drGe
vkSgRuadVywQzjRamC41nTt+9nZg10IrK89gRn2psN/eLILj4UXkIaXh3JFxjhw5
aDn7T0cL7egZk16ryY2kKDs2/g1l3Gah7WxrutjhO0EL0nd6CgWKxfxJQv7nSM1u
m72nvrTQdwqOSP+vVh9GytlhM4uL42j646tK8i9uF5ctFix4ur2vI6aLRMZkVBmm
HsGz4BCz8s69qUcai76qmHjaJpgCVbjJhpFIYj1zojy9FDrYgvmdWfUH7Ga46iEL
LBr3eFyAUH9nKQopEoECV2VQ5S06wMoJqYqKwUCVWyqBuhnrMs+V1Yu3ocNbx5Q2
nU88QaAccj1tNuswek01hD89EUgXGIOVoJbJSwRn5xUbu288MN1qEo45kKGdofhX
JNejvNJfgs5YsGj01+v6eH5nJbCZhHeVe2mj95DaJr+OR2ocXrhzhfmDdmvkBfN/
MjC5CTjpUbybKEUfcjyqQwXQAq1AYmkHpZXwoltn2UDjeIOl9eaxqHDlHIgrpT6n
kifHeNowmjl0XDsuQ/EFV+3EuRqg7RVv36dqigZsF4l+30XrySHkQXV87j/EmXn3
UV8L66h+KYW4sCqOHBEkB5qExSl9KOBmDa8hkG64EYuhbNVxISPYROGR3NWaS4WX
VPiNQF8mj7zpL5qBayIUu+TTnnl58uuQB1T4lHfQzxNnZgS53RKHHqx0Z2qHQMs0
DNMwo9RM8uXRem7I3uxAw3D5l053MsHJCWiBWS9PjWvghfhtBNhY37iPxQRgtdu/
nP/DSFQBKkoPYMdTEWo5t5fwxP5J6t4v6N8owrCc/SRtiKVOyzDaqluU10lKjZxk
CXd+I27EO5RZCat17zEbfphok6XVr637zpayyzn6Pxrb4VvzbbGug4nXyecfNGgQ
TvimvtJ6bsJdVB9PrXZ//JonJADsFQY5TxEoCGm2B+UplZkvfd/Z7lUw6At59M5M
cv4ZL/HIrqQ8GfjMQkX/mz0R6SUbgsKFNqZlzCXMU74RbmkfJuWZbOMCYaP8krrU
HMUTA5j6hQ7yDt10KYwJLUWLdLEKN6bOV9yoP9xQP9KOZrbXvj+X0FL6RKCGkHwj
Txj1u8xXZHwK4Ft/5M7RCztC4FdsDW+jIW97QWKuH3iarD7BNh2dDoilK2kLCQyy
lzRactEBgWNPhG3eKxAQcSPURFSwb1UwoEkqtmRjimZzfTdBgI8iAlzvc4Lv9sFH
vhe8IGZLz2kH1lCCcHK9P2DjLvUVptc60IK1qOydD9o3gy81BVFEhPqY2HPecwaN
8Sk6YxU77Eo2MBxNg43hW6eIjXVbxEl0lipjs/QhJR8Z20JWavt7jqCJcdOo1e6m
lKQJ4gaOam6NUmxdKBTmQ8kLNc3Boo8mA74q+S12AlnkRQjdNtolVgBYlaNm/h45
VVwj7vBSNrJD0cEP4CpBQ6Axha+ZriQlY8VecQkWGW+6bSUK3Uw4XDXZhPzpg2ho
AQSNBqUDVFZIywCR+kiTL1VQhyqEwfgSVajivXyEEN1KK/Jvwq0c9i68mZ+2UqI0
UrQsH2ZzF8grKcbp169YBwZN5elgVrPCYiiqpRNddGFDtn74XPyzwLtfa8lm+GjR
Ll5FXjPRQLOoNBbHpYltqkc5wK2NjuS83jN5cMUP43Mhl06TO95X1JCy5ewfTM2m
Tl3wb2cOIzesYmQE4Jn0+ogZcxDJbmxWUFMZKiwkBZc9AjtTOBURGsHjHvx21v5/
M/OI8iGoQlphMcqkAQc+5bdcQ3vYW0r2bfaw6SAfhvBnA2h0bP8j/jkmebayNx2E
DSGM7TEu3DEhHZZXimzkwQsm0sxPRlkRtuq1URAQgvcdgtv4w9AxyyPzsngim301
YCZZzkZtnGJx4gxrdhcMIXDZEWNzAx1/6fSNOnliThZe+JawJn51Jwfp2VcOqbml
0UI0jrWT+KLQdbe5OkfPbWYw+K+kAd41xtnRf2fvHMQIUNuK+ppZ2y1sKarREYra
oh3uzEtNzmgmdDPSFH2q2SngMU8ZsFXhHPeTAP6UcUkDv32Gu9pN8IqLHQ5n5GpJ
AaCNeOPyj6FS+QoJyk2l0RiPeV5zb1+m/k1DM+5zIw+TL9G8jyA9/5vqz9d1Dq3t
TALE45yBdIsw0TrpSVagtKbKM6eh6lpUfBzsOQ3aCkK0C1+7Oj+kqmAyTo1O10cC
qVvY8aFjc8qu85KRxXkiJa/nBueQ6fM6HS0FY1yZA2ljFbbrGpNaHaWgK6WxpuFO
vnnQoEnkxXwDySqIveQ7iJ2dy42IPh8bW+nft2rr/x/9TepmMH1akMwJTi1AJcEY
vDQzmxpAwDxIniDp/6lvgNT5qsH/fjS5lVEXN4X5gaA8z4P0Owk2byDnDz5gUV6w
mL2/9uBDLQzNtE2kTdo23Nt4KXiOnA/5ZpFTDkQ7Egw9wM0Ae/Swmd3PQYAk+0Dv
wHUr+wysKYWMylIcAvBfL4mho73Jfz1amYd+17zJVM2mUcOZ2OFzmgzbld84Av2E
HyxJBq5T0P/JdR30Y6AxRu7AOl3F9XuvTtn+2nWXdS5bt6xsYGEcsedNPNPe39Wk
5n25yjyDc1ifjr5z+g8w84cy+EdzeyNy8t1i77AHEb6uVx9VgdtADxBzIeF8h0tc
gPSDXPk1/HIp67bfF1RDYmrbL+PHoTyjCyRvjKKcHh6HMaErX17NXNg9Htn2xqTh
x2Xy5hXNGWz3/6LoYdapPhUXzwXTzBEHeFMkgZe55ACNzqbZCFgcMFVsV5Nrpnxk
xiHe4IgEx+jp9QuPh3hKwKSdEZ8hPWMPj/MI28/HFJE2Av+G06R4Fv9juHyNexBv
x/HWA0affoC9kqgW4sYp/4EwDr7XkQ/45sl9LOPF3ekwdWQaByoIVv3q5IT8rxrL
n0pKhshmg22DbbJtZrEZ0NTX1CUUooLkYtfcI0eISdPJiiXYVzQ+q69vGy/DCGUt
RPcDhpth4MULNGnEEYk/dV/qroV0vwfIgLIt2bI2eSisTWG4r5LBvBIrFkqPgkZ7
zZaVXrzjCaS8k2Y+OiXGMrjIVwwFrclrrqJikvApIOreQ3Pb+8XdW+2gl9YVdGJO
e823KEl9XghCRuL2aHtkjQ2Gmx5heAJnD78DtH8MwgAMj2SyhaNPln8Xof0RWKoE
IgFMrJ+NZN/FA6JVQANjbMADhX1Be7bQksUr3SkF+GnDQgDy0morIumBCcwj1v38
psG1f8UQMwUs2SAjnaHUF4NbJwVuTTnZDTDNZNvt8JTfZU4Y/N/Snmx+tNAObi6r
7hYYpq64xF61caWZrnXpyDuq9324Mq0TBa+VsX/p3wbTrjWu6ADaVAhU7lDodAyG
x7k3+FemXnZ1b2r3agOqMomTjWPMkbTzwnsBytoj1AGYuOaewg4AloT+3+XVvIZI
O494ggOPWBs+4XBY2Xl+ZY9ZvnwlGkP9KfUW7H9cF5oap3wqc6pckbtFMdW3ijbd
M29tdzrR4Ncx4yox3YcTCb7EfJT+QVwMh7OE9F1x9J9EH/s64XA5gUTCNaj8yPq0
6XJvy/dsF0DgMHkhdGXw2Jtn4zgp+yUQU9cO49wxv0Q1Z9/XlqDadqRRLBa9bCfR
zQIdSDYLCsFlFSrQDv54sWsGp0Rh3yBx7+6TsAjgBNWP7k8p9BAu97XPwiMGOcuS
HwyVwzeUf6IOUrHJY9YxyIvU+Kw6ZFSofXwWhPfHmsDGmYiTeHMH7DoZS4+kzapw
mE2g38kGqe/IMEswEM90aNREIkRv01/8obhot8wQpGbvzePkKv51AXCniA6RiaOW
6p2nzxB5TnL8ZgPdgIrtmZR5pZnLhH8me+alJoth8h/Q/ekyGuCw8CG/5NVLe8j0
Mmn5J858rA42nODNIa3j5xqhmlo70gyZpVJx/CD0IpoEyd3CyCvBBdBscuExy293
agMztqNa0jFMTrL4mP7xrEu3E4JrV4pSwiwNRMMQc6UeiTw5k70eQZYvFwqA/d4E
jG871FqaGIdJ11IR+1DgzlrWltWW/wGc47XYf09mx/MNV/OhxT1d4GUejRltW5dP
5IFqEe8A8nCRlA2PWamlVbp08/IpjKticTkxMJuJ9WusEtu+kUuaWMg9G3U4K57z
sbo9BOXImMzczPsWn8QZmCUxO18JsVXw57e6uj4GOcglEEYr5J5YyqDrUO3iW1yp
VrS6EdvuA++egt8HAHoBvl8dJjPoEDQ9nlz9fbuC1Uw5JmlaFjlDnmiek4LouEm8
J17SdaZD8n7LNb83icdycl6a4AKy7AUyVo/SsDlMjCpxFY6rCyyHmjajb9YL+vE5
2jx8PyvK/rbtAaG/gmbUyrx4Nnq9RZitHaQU0utN0SUQt84FS80eJrDKRAVVjXjH
TA9+KB1UFpAbeA8Utp8yvHIJDYBUe5dnnEfovgJQp6HsJ2l+mvTjwjNI6+I3s2nW
izJ2ITVdhEMTRMQEnC3Usgf1h1h0oH6cFbgIhlglNgiPgmG+kbRVrkuDiSmKdrnl
WdLwYPhjvnHjLlKDsgOrUhcEV9MrWhuSxqQewCY6lgQ9BIe1Bv8XkaVtvvsP2CGJ
CBOhA957Kmu3gwOyrKR77f3CBHljIn9O+gaT+B6UVEbn9NGKG4eSIRVtiCYs3n0k
0ANYxUoApuskq3cys87mcKrgeSzyuYtmHZlXNQi1ct/LfV3+lf5RJe7p1IugddP9
yId19+Hoth8UszOC//9cpb2HaT6ekmWEesFj7M/en06ka2KrRfuGVoPVs0WFhsPu
T0f9ARKwRhBqrJy45g4OjkrNJr1TQx9bmEH+oDuOScd7ErKmnFnqmB1q0r8yEVF3
64BK2jFk17NMR5Ey6NfPxJlrGGYrwepM0m5cpQcMRvfUUUUzqbUUoa35yJwE4quh
QvZaK8sQUZQQ6cE/RHk/aa3RK6/2FhqeVIZgl3RGCW2pbqhNt9yc5T3fbcCUiF0h
rmAc0jKn8gqRsWzeh7Sc93qNX46xuOXZbuMWk64k8claejAr1rDip0DfGEfkiNjn
LqwKXxxKfKiDtv10tTetlV1rzNRWZfxKWkzpQFBIUdQkALknf7IpZSk4Od9PZJDB
/4qBtOZG1WkSFm6OurxchpxuZbnp1SZfPLT+CVZ0i3A6W6yRGYtnvhOWeUSKyu24
QUbgXG/gByovFWah5Rf7vHMe8IrNhxBje9bExew3niblPP/JzMi0VtVxcU/YyQz4
S/NohkqVT2gsH4nZPvjinE+F+CnUtTUjMBfG/YRNPlOZYWI6epR4JSjBWv8oFWl1
2++WEs/6j0ikzxPmNqRqULBOBxBp/zLp679Z4kG3zjION3fDtwj43xNSvEAu7imW
1CW9ayub6B3lgvzwZTy4GfK7zj0D+bNKyVxzhm97ytFhui1K5uv8xLQrRSSPh8OG
eKyXf+EoWkpoe8OG5kdZrl1HgBS9QnYldd/AeAj6Y9TAmSY+RugCy07mDTZbbspX
nzt6LESsBvCknLoiHIeGj411CYK+g1SZl9L0FKF7n9cB4J+UcIDxEjflflEL16/k
6mH9oBtk39zJ/jkyv5ajFwwV9Z0dJr4ZXXv/h8cXUCP/+r+SnLC0xkrHybRpOUGe
CDshxLReLTTZkXrIHz5OeOU0IgC9nfVOFzIcWGExHdIrUZlI1NI32KxB940vTD0j
TzrwVFZMRlLFsU5jG9mkhYETFwXQb5JNDNJ5EpbCfOLRZ7cOpdBMwBcsc3CvhCCw
iercg6Cc3+rFznQY4GNEeJ2dFyBXnz3GbfLoreY+DY6+N+8p/j6ZVoM9npVsI/5y
T93CUbOozdJQxEcIByWlHtz9//0HyUVmbd622hDUXSbjniUZbvTcDWzEz2DpuDQC
H30c3xwVXAJFt6Zv6AoCA81EBl+0eJed/Ge9/dRrgqGt8XVJFVrHlMue7b2FkQCq
4MAtR/UsAa/LG7SLvaJJUJQrD+b0b80NBsge+9CJhbr4Gx8yb6OA+BS3Fehye2q6
BMGSdfjjAKGTYkL3CchU9qr3FPkZocqCxx5nb9yNVOiFyx8Wppn3LOgNkFRcOY5h
vcpsaEzmAilGpXonCc4QRZI5xo4gozYkcRhUFL1P1bIgxLHGykkiyUIfXBhdbGzb
a1jDO6uANR+e07QmEYu8yAbTxTfd6K1/yv90bywr5sp8lEtxeQ1m2aliWU7/Kldf
mksdhwNramOGYjndEZ4PUpjCoybOg3b9pZdhSb6B/cgoVGyVqZhJG849YGxbNl4P
oCI/m+JHrR4DFntvw6O7m0yIKIWao/wyV7/2ikrC/Yxy9/h5WCoqn7JbcgDZQZCh
ew2IbGCFDW6yNfaSE/5qI2+V6unurRAr5b4Uxh6ro1k3aDzl5XQEJ923Bu8JBVoP
o6QK3MawUgTycunAXLRZZx6Fvl1/0IhNnvwuZRapJBK1GuVaXKcX1iASUtH4qnfu
1tNHoLCcBVWC/mEfiqDmvajmy5G00G0B65Fda5dD1GRtMbxzARRP8j3Ku9lDyB4R
rXxh6UXlqpm5wq03JWBwE9ts7Oc2c16rUZ7iy9Qurn0i8aBhZMjmnV6XQTEBMjQk
Pn2UJfN63G4w7BXnNAcFsc418mpcKa3NyJLzn4OFRZQQ4/Py3hMeVs+73vXFLqE6
tpkjtKXRpA1o6rkfSPrWfXROIqxP5KP99Sk04JORROhpmF/UtccYxL5aF+ZirSqd
9vy0JGhCFeLo2i4ovS0ihp6MsDbp+pi8HY0vOyre4tYCHuSDsWJJuzkrkToR2s9N
oM+vJ+vlmd4z6MgRO3CHEjxmdrfMrsg/WbS2okMrGrPK5Ggb38YHVrcthGV/46Xv
WUUFqb3Jtk0fm4NPZBVRpKlc8gBKiI0IxrsMQcOtNTyY6p1LY3Tx5XTH07tfAeVI
ARBNPH4QUJyTyK09wya2A0My+BnDkfJbUjKYYZ96N31+BhHCOhW4hAmAoFrVvGep
xKs81m7faRtQFhRq9l62T+l7S/UhYscah8VAKkTVXtZG+2RbYPLsUqlJ5lZwaWU9
wtt/qPOHYFH5yosYGCOplEFrAG0M+gg2HjtzgrWOWSwLLdhZFpAfg/coTu+FJq/k
OOjMzFmdRekKVvPWIJ+wcKNap2sR8Tw/XV9eFN/+PJDsaL9R5+b1V1C3ApZwJAH1
2dlPb/QJ4OYYqLzrBOU5GfdcacSKBKndLztNoHElSDX9KAUAyNTWQHYTnWDpCSUq
3u9Rn8nI59rOBcIdvN0FiRekvwoX/CQJdO3xcCwvPaTQDst4OoHC1KABjNCKg/+P
bUjCgAVoTu5wU38aEBi+fxbdcuabMDEoGhZhat9uBui7uCJQtT3/4xGArClR3Ili
EKL4OYvqSEVkz9J5qhJ62mq1HVfcPcUb2as5fpUH7MtWaQRntD5m3m5cKAkyaMw1
k4CP9fVEDXT72jCBejwXyUAPo/ILyXrPR8GvVmQAnFlMWlLIqMfPnLK5Jd/bIOne
WnBUSqzGuD6wUA8akdRajNqL4jet+AdZC89RRLEUIRx5W7D5buHx1ssZtbsbK8ZF
NrC+UoRV+iroAodt26DDVkw1fU4oK4hygUWXpuWwmWzJ+0ErWEdJr3JGOw5bF8Pz
Lv0n8d9TuZqrh4DP8ItlTYvBaSdKUIQpzVBJg7yvb4peDQUn+HVgRe/mD8tUwKf1
1TkBUbAMj2FW0AKmfObkbS8mlPsD9cfX92tgIzZOpqTOpJcjbyGo1y6Ca8xIRMRZ
lTe5bPI8dAJ4ksnLAl0gFm96TqDFstZtmtR6xBj59cfQKJi6lYhAWRfpZQWX7Enw
ASNQvKYuVkEgg5dFMfkFNxIKehIIzp4hEkSq80hDi2sA96V1rpnVVfLh/tFNIlS5
tMiEeqZmhltLoDzbwK4J82w3+rFubbt5hhH85GBMMJRkDAegXNw0MH12X2MAVl7k
SBSN5+E+v0Z5zHLOdLbzpA8EmPob2lbxKExvpbaf/QXuyONRh+EAOdNuho3N8d6d
m9yKgWdh+Z+U2D5L+SMnH3Fyyqz9Wer8r35FLtnIGW+Tqz9yBi8wgYi3Jfs4CNOg
qYEWmVi13H3clexkYHrMvmVFoky7OuXYk/qCaAsv5HaocOEydOEMMrCa8qGoh4JH
Pqu2jZZp+zSuGSDfWnj52731ry1yZzF5/Vx/n3U4S2THh9GRJDh83B32OjKppkuU
k8fw9z+1RDIDJrbfngtV995d6mCk7l5F2kRIINlHNoyCFwfWDSzzlbvLMixqpi0p
/OW4JWaQ+GgMsB89vUGEhDxbsDjxgHDKtb0YtVKt6Ov7eoluCsFCGIaC75fvUatv
LSj2rRDEMEYfwo1jI+6ns7QsB5Rs7WbFkNbSIy/J1O5E7y0faj21Ns6FFRLxLiz+
b0IIDs4/zqyQUyq4LWdNy2enN6bilBzhqD3+0w4QbLOYUV1oUJ8cYT++x9WZejOu
mR/3SazXibcYd8QAqQN5ZF7lSDS6YuVO2uzb6FMiu5LOSAEjE+M2Av/cvmCNBze0
vGA5xH7fS+boeyun6zY/17ajrIIY2pRaGWAp9ygIB0c5YhleI0Aoy3tOTq3yKi/T
ueWC1UePXp7A+zCu1EpKzWZe6cZV1i4L/YXewMfW0j8mOA9qF8AbCL6OjrSuNF3u
5hh0slB3KrUXKT87tzaiPa4MPHAvPTLhJg9L8TO1w0lfY4/LmpJI0bQzS+BCzJxX
0YI8XwjnXoLt2NS2PvrqatbT4bZrPlKaxCwzUOS6SGeF3t9i1yzTEgBOZyb3y2Qm
58XkfPu5vMNnftNtkL/AhUh67pjiyHiB7UzSHUlSURwsxFoxu+DOJKLGZkFtWUAH
GWaMBdCANMwTT5nTZm+kMWtr8iMTrVYW5/nyqrglsgtaO5OcXoU1svd01Fo5vawy
v+1/ISNB27dMgooexz2B4EiZDVE8kcAfACMswMajdWqqwwQwBQ+cgxozJuU8lYEu
xBeFObWTHuDO/D5HPgV2fe0pZx1eJx71/1jIoNpM5zenbLu3X+HJRqA/Y+ucnmkx
13aZbWnl+udcwSogQ8FsgTLC+wEpGDxaXZO2HJAW7419FUUwep0VDa443SAhmm5p
+827mpMLq1pXOHqBAzFPJE2VlWA2s0pWrCR5yD4cwoAh85rUbnOad9CMRivQ1kBx
EVTlVtlffExOjJ+r3C2b9zZ+uectwbwl2o8t7SJuj+TDBIRP2jh2hAtztB8yWzpi
niuhQIGYvJxXCG7KvEA+E+AaAGZtpCF3IJNoeRWYQrn6rsi/82RNZtsg2kJJnK4B
+iBkPcBTmk43zDJoqDurwfOcE+eWxRBki/CUmWaAg/W156rEp1P0sLS4PcZIKqAU
MOujw3WCRvRcHCwISStTZGPUZ3Rv4N5JqieKqF9xyLiTydmgXF5WK+A6TrFHgBhr
aGKBoteAsCrPlw4ncJKPeBdvXXwz4TZn3OgdmiAuFjoj8bs9iDpQThWRd1pK1l2F
A8AkYVSHmZS5wIyFWaUin/ZCWEXi3Cbo2Qs3a7/XzoJvWRfLaIm/XBYoshDo/7J2
feNjX+v8AobEytilvjmHx/fNt7egko77cybLKukpOgTrX3ofwjAziejPzU3WPkbH
/xA+LwKGNlqPIenaK+b0eDlIzSYnxRKzt32suaJIjAlBrVwTiv1KUQIVTLuqJ3Oj
TRUNld7ImRQRyAp7q91frlpS+VXCLszrZ7TYG1tRR0nUIPBUDWpJagGBDfMUjmNw
OpoRzC0wJAAAsVXUkh1bQ3AlabgX1SPL0PjbrQTCh9QI2mpmgMLi5rkBwSYNbIyy
1n+eSplH9+oOfh+55OnMzZFAtFrXPUnxGrNOyI/X8ijlwE69mvBE89AsCNK4a6Fv
TWhocgEKz+xsnFdGLnZ7niwrqcSh/tp761EdbJP9FxFKJEjldO+ViW3VR4p0v1qI
7/GF3nmHRyF8Z/waYD+tKPp5GmJm0yIJiBqvlEJNLg2bansJGSnoE4KvFhOiKweX
xREi15ufq6jymjSSFT9NNORbcW89RVE/R3S43QOgmR4QtbDyzIdLjq1Ssj4trYMn
tl3P+8yaENvB2zTd2Gk1H7x6/rEUfVLyJgan0uQXaRLIUI2TqCjdyMZ+cqobyVaU
Q0wCttUfGPIl76Tn0oMT6h/uLKnMtaPAB321vqGPDjqw/d2K32LnsYzEQ0mnmfVw
tV3kIMqX6CJKiVoIS76bU8VXVlyK6Z1ZyM7/XfPrKcANYwl4WzBvQxhzZOfBi0GW
bgvLnn7LTGqC4roq8RLHFecC9aJ+wxHG8KoqUxPu+5NMd8EjqLUI4Besre1wCvfW
KwHVMNCqm1tycnKrj9f4b5J4f4/BIlhRqwvbGkfm63U6mvfi4m+Z4bmi9aXg9DCJ
f+May0AbMhENtQln8OniOqAW3KLs+3Ip9T1Aly+Hse9LfyzKnnttrOmvsi6+yNNA
z+nT3o72GwtqYG+eSH6jlLfZd4k5hA5fJBaPIjry73ixkrBUNyTw802Pn2l7WqLe
RMys4aIWNfaf7dWa5WbER2TzuKLHkOqz0ALQfw9pmhHL3e4nQMJmQtFlDonFfxok
ryFDpNgJrLp0fqkGUAqke4rUEQv8KCkOsUgQQjAOcWC37yiDF/1p9OfLrvkASaBw
vVWyCf5S9PVKxgetlNONtaYMMY/AqhD5xtAUgzfWgez5sYhcvRc7ZIopD1m2ZmOI
iR/cqJjo6oDicRJ1FQdaVtSwUPobVxeaPEGyLjSLvzudgTHzwl8FUzjb7Mp0YmFE
ffy7Rvjv679Txg0Ahmz5ufNTCm8xpN6xQ+9KsEOPngLVb8w6Fgjawdgas7/owHpB
UvvPDuXqHWj+5pOA2u2ADy6OPVVpE12O4ccPHo2yMQjnbcGWtVFYtSPFrP9mbmlE
QarJTfU0CAFGs4T/wXJZstIkcEZst/ms3zH2AiyeVXG55jTKtCCEZ+F+f2f5Lwvv
8ugQI9ThXeH1urlwVjOCtdFv/Jfoqt2fwtMceSUgJ/qguY5dyoIUBkpYikPEqjd5
ZuoFbNVtVwDuMQ5BgHa0Zp+DUNIUh/QkX6LoAinwhu1yy/uVgRexSuYAEu76AW4M
929uN0LV8kutVOlxzof7n7j4gqbgYSvigGdXpadu0Xwoo7X+HCUt62IdB3v+Zrms
2OnlT2oQtSneqd78VU0ChJ9NVVcWrQFQNI9+LkHGo0v0RTeN6YBehCZEX8OrRIC3
/1uVd1IHRAjx+J+UqqKLCYE1sxa0No474VBEF7+OdvSWEMU2lLV47TQsNALgT9vK
Xlg8HR7ATWFVyGW9ZNZEqTKzIf6EbROXASuAtUMiXOqpg3Is0Noi2RqGQjAFmJ0f
rMcURumtDunW5c+12+j7QYW/qDQ2j4YbOll31zinhY8bEsu61sJEtNR5Q4Y87MVb
BPygTJxAo05gsKJdpr7N0cu8XSHWIR69Q+1VTinuzHryAz1guzXFSBZxyLDgLaA8
LTDTrv/wn4LiunoxFvHU3eWKek9SGH3p2fZ5ZgeWkYty4KVhgWS/v9MhZ0FdbfJp
7OTGXfPQKqw0tZTJGT7rjKd0BSlFI9JFmYS0rWlVQNpNmjKEeH2pAhZYFBmgShQf
pB0/YABO4bAX5LZs+xHsF531/niSs5VOMkJYntelhSVTet+8BGaac22bO0iSxEKW
WodnoJCXWlO4pOKn7KaCs3PixBFYcwZqyTt1zcIpZnULADmoNQgMhX3Qme2QW2Cx
der7JOVB51nqxv9+2ng1zNa4KMAHt2j+5vg1By9hRRTA7t+Tff+G1AjM0170MYkr
NwNpZAb3bTLYeujF0E1jEO9BDqT3bK6JePih7mQIEdHeCi7TDH/5JBGgM5Sh6YSm
amhVkhsC2KU9SFOdrXnfHiTok7S+SWmxU/GE1ReMvhMA+CvAXG3wC2kxYj3Dt57L
Agx/Cp2KigJUFC9BbXHoqT3xcDExSAQei91Pj39bbsHYWq1ieaxVUy4NLoeanbOJ
XLL8vBcgZMxGqSj7TgxorIzU1PgqnPxYjzWHOfCZ4X6NQYf03J2ajt4bWmUZkCoo
9l8WwgZDuKkkEN2okEcE4i7D5+xbh935FxQoznDlN+fTvS2Vt05hPdwYT1g3PLH0
B67NEbRM1rycXARYl0nLyUgnPaZ0ab9ptefzCo/w09joaENkGWZEXp5+2UDmSkjv
EeQN0QTxuTEsqMKGg05f72Bk0hm4rK3lYOk1o+XKCEfvHwRj5Dio4X8I6H1B56oU
jEv6eLJ99GAJuQe6UeDMVkh/gOXLjN6V311OrVqW1q1iJJxQrjJzgmswRLja60z+
+3iYvet6lnN8ZDr53OIOip4xgiJJYp5y6QQGfnr2pVD0ZFAhHhanRKpIOOSUqaOJ
GNw5uqYDvednS3Cv6oolB+S0bxso+L4wZkrjtqKcNls/qKxo8b2fLdyXCUCqOJSB
WGuG9Aq9wnhrgUugMqA3Wb9Uqr9LVLcGkE4kvMdCLbJsgt5elsTuV30p4VWHN6L/
IINHHToSTN1PDYvN+3o5/jqv0rYwDLn2IAbD/N6U02/JY11pak0MBG5JEKbEAZHH
O/j3+xvYtnOuvKsLDNhxwKGuiyrlek0PnriHE+i1+IDTgYaU7gg/kbakbhmdKApM
fTotHCW9hdsA6ZS0IP4kKxAVB2to3UcGR6xYUNEet/asQmLXWkmfVYtCLc3a5dd3
FN81acFYien/OFToJjKVa9Q0wHOXb5vbQi7KA6HC9YGt+09RUcHSxi4ivHC16HB3
80/Bs1X7KzRywWbf69UhnxbQxttb7qXqQR6Qtt4iFnDQbIgEOr4VeApOAZJKhD4h
5xP30X0k7xFhDFI8IesPZ1tS+pzFxt9GqC/cnRqpAUjLJgimJvv8Wuit7DtWsK5V
Xq57CnO0D1/vDXE9DBBE2xY2V7g4YP25HFBDaoctWFQGi4wN8umsOih3ppjz5koA
zSC4duAWi5qS5xNZoZYJma9Ds95j+lIPWWfO1UBjxIPMtDlWrJSkPksJhU5ywBIV
f6Iv7UFU3prUyKAcVNPovLfvwXbyf3etA00t4LALDlXKzlVO1VgQkapz0bBqwlJC
GpYtyO9Y0XgtWaBgyLyoIN7m4X9JGoout+aVht7Kjlcqb6Xrca1AGXsjYvROk8xj
fgNXUr8lFWOKwMJxMFWeZQSj2x2mZZu9j15IGj2mzceXt/WQN8v7nD+CVF+r3G/B
HRtbWUK4QnvPUkAmoQfg2OaHLfusSoQyFoxn2QAeSqlkdsMT+ef0Jz7cmACF0Jqs
hIm07HvwxgxqXPOUbT5t/OS5h/TYe88VgiHB0Kimx52TzrAU1gVIr9K4et+fvP6a
gZnPhmhtw2GVyeQ8msSYwYY87IEb1Mm9wAEt6k9jyvSwkjCXLyH3OogEViTLtuVY
wn7+vEVuSCRUclozmx7k0+y4GeKFg1BX72z8eUlPUHY990cg0eeqvVc5ovuux4YN
FO5+V7/YO9JlznSyzO9MnzRhje8zxsg2eEB/IgWEdBIinzoO0IMVF2W1K1cOMD7i
eTEXplTY2B7d6ZZNT2OuROW4Mdbps54+MukQKSt6dE95psG5jZWGXZg5OPcxsLHi
zjyQ71YiusTu/ie6+dZBYmTI4e9MtteWfJEBt55/hkMiDFSlyFc+phd7gTvhSWue
d8Bjk8/LohCJ8xH2TXL/n3NV1QqfZpvN8CSeAardWLCmeB4X40AENtR9b74/c4J5
Mtnodd/bMUqmjUJYMtpAC4C0sEKTMpiOJHU5eJtIP+mDI+wjfNzcHd1OXO5gY/Rm
Fk+EcemMlzrv7SuwpucAuxF1fEW9ZT4gRHZSiz3rwAxeu1IB4Ibx1k1oVLlwXwH2
nb3b/xCXVFxBfHtrU6OJeZwwtskofxeegxe0u36ESEGi1/gKGYFPucYENZpl2a+d
NpkkCbIX9oDBSL52hXEy/MXbJC5uHl68elgwbry9/jliuLAqverBOjJioIc3BQAy
hN0+mfQhKXXrd5zLnRwprvBY4DDw0sC0urcx0g2p6Bk4fQaYHHlHZOXNP8s3rozc
NT16+RWU3LNSRc2hFuLdxAvuoKWNeZD9nRH2siuPSxa9j7ivQkO4aFttftv4NsPR
IIXebmlDElLEaZHkoaClALUCyEwgFZ1XL8IarduoFsWkQIgIDvljpYV7b/OrDVOI
zB14qd+Hqo0FQ9FLRtbHR7uLv7gx2oM8PcD4H/vweCmL/VKTT0IZ9Lpr5tsidNGN
MqUa7eI0KOSJMzW1dTBv7MT+DgHcYjfb9eL1+qib+VY2N6YI7eQYXDkWHXSr83cT
WNXRe9gZzQsIoWYG9AfyJ1ayrJLjGnycUx6JQ4Lcc8DkX3kCl83erEaZhQDj8ICC
Ao7qowzUSJowXFhSGLpsTmQjIf9Oi1C1pmOLKI11vM8i+/cfRmxwzqtqbKEaCvTc
+QOJw0MX3+8d9kKzcZyp8rpwSQYlYEdYhttt2NYuwJVg36Ob1VSGqRvrqBkRGZWQ
GEwhs8DJpOhg6dI4abthN3gS9lIpqCbuImgECKXZu4oKZg7qySjub3gyJuEoseFc
k8yPu/j8A1S+OakOvA8WozTsR/lxB5d96d3XGX10tnxbvqdPJQkJK878yMy6nxey
pJDrushd3F9ANLHQqCCsjCUdAfqVgKTyqJA58Cf6zb/RCEgr7UGyfsRiJA+pw2Xc
naVJj9hCHQgu55sDMFZfzXtvayvifExAG61a3qRg5KMgI9+hpxawiYswaV8LTxVp
f/b/ytuyEeE8bHDyjYrxJ8D6gz/Pd+ZRVMTyu9EugZmJa1Ym1iyqu8fmxBR1APi8
x7rbmSqqaOEj2X+r6hJ5g9F+dTCLa2Fnrliirwr9ZKI+vKYy+i+kFGXBt2eFBQgv
mV67b9T2aGOOgGLvlYY+gqfd3JjMyfjpn0rOQ2TvSRtBHO14xa4GwMRIQpkU5WdM
D0sTjUcAsuKqCAPZG69gYY66Q6pvsMDTfVv9dU14J49orN1l4wyAmzJ61X+nS5P9
2OeVAP6Gu0Ode97jB+cVhu+2b7OT42O6hkere5vLzPlsduKyrY6TezSIuGxYsTgS
LZhbjEeLAJxMiR6CdrmwuMK8vOKqhai8qdHkRjG/micAvVqH9t17YUS+ZD3DuSkE
ILWFNqoxeGQx7a6u5zU2N7MC/6illzv+CtkF59aE/8skh3LOfXDkcgES7thnwDWG
EOEMrORa00E/E1ysXb6UozGR0LPsHM4mOd5sWKi8OxO00Ddn+YXebwDwwq1AFruN
ShIhP31UJD2MNNpU/ICFMJjYvvX7MeVAr47ONrRerY7rtgkz70CIwbutH1ZPKAuS
gu12E/XdVJmFgvC7IE7Lvw/Auf0/3tAC/x0qsiHhDCwJqZRoB9srS2QpTUF25DiS
KIHvwAxiZ35ObljC1Un9c7Gj45kwWxG0n8S0nwa0Nm436zk1N9ZTFKCmUfxklCCL
HLueGer5ztRkXHPNOrIv9sb8iTS8TfTpdZS6blC1WHJu8XVuRlBlbqjesujHsq7i
WP9XyzHYTIj8ZwFAcoknTGKQdefoM4UE+4ijihvEHEdbP9KtgL0wpR4KTVzHjHA8
hqg7Ml9aQMfL9sQB6l/K5Q8aKD+wWyFwDzodCOczVdHSesP4RPuSeEh/7EaVFwWs
zp5d2RZ18pnJ6T1j8L7+qFRQ83dIBiKpjyoIT6L4/LkcMkRgddZh07+X/XjU3rfQ
sT/vBhgourbZXBbxUkKFFFupXYCDyNKzZQk6sFeSdHjq5ghn1e4SBVwMdKyux3Zc
XJRkn5yS8kcwRyfMUU4trz1UOoK5yWW5D0OLVuaKnOAJa42T9kXnvO9ID0hYac87
ehx2CO+MDEimwAyTOdgDVH0+LW55MnyX0izqqUXZZfBNWwHKBnmm0aKjzr9et2xR
ELV3JsKhKLyXPDo3DA5op5Mgc7hAekyNeJ1z9CYrq4RHOdJNpSNK8ab+LFey4hMz
NAtaHnGrIh1xzsAPo9dFm8lCudfKJS6ISBRxcXP639Fh28QfKeqy1cpp1jDqU06h
7ZYT3XcDpwXFYRmLy2YCJ+bIoS2WNuqpYcniBDOV/NuVWMckBKFQulGbraJiBWu9
qbJnkHoav9VbUHXFv9QB22aDpft1HSfIXYhLU2qWSlHwRaQ/AgegVWz61P/+YC1x
oS0gS4G7aqFcPCR+CVyvpMqn0czzBf8prKQFsJoxGBWpeVzXX4fn6Z4rjpTPQ0lw
+a8hh0jdoYx6XaoiOMHROhCbgbshfaXrDpHGdZ2Loay6HF/7z9nr4rxmpUkoIa5N
3WUzN6Wf14aB7VR9NF5em5KXxzH4lAV20fSDVY7tky17F9iPRbSdm7cHEG//caeM
nHCdmmUHTsQOZR6s2Iy+xp2VU3cCdWaefzRnqw0wvpiax9l6NZW3WA/7VzuJmVIb
WQsel08azgHaguohrGyVeTAq8p8+yCtHEWCI8RrPlphpM0er/RwaWdm+jgbNLpo4
l4NNDCiEic0uPX7uiUucxGZw34oJAUMtUmc4EPBgcvsbC1ruhtTB1C1m6oFKt6TD
iFU6TW/O+NkqVUDX9Mbg7YHpsmtRMAeitHSdEvKnkaGwJ/vvNEM/98BhhupK5xy1
+O0qLdjxuq2VTOpTsm4mVZIRseqV5hQ7ojQkdrojnYiiYR55qH2V2I7CF2iD405Y
9J3yYcF5VvZ5d5siGaxY9ricHPsgYFIZtdWaTjaVnuHa8aauhlMdOv02EgmTX4qI
UmVKc3S2hNUUpCcaTsiJvvKcLXjgIPHefvAeo/Pf31Hy3DR0BahFO8qIiVNTtJbL
CuiKxZbh03ayY8vFqNWnFW5vn4aaQadI20JshKozFO0HDL7SCXdxZ01SBGnGAuQq
BprRKIEfxSp50VP89qKyBM17jdRwjAGDqSR3mRoahKH9TYOTIszAifGpgcZuAhD3
V5AckyD6E1nGo/tDfZhlQLtvHGUEmx6lsrWPdCmGwMPgKBRP3Y/le5LEN859tuo4
WJbC+eR2Dgwe2mVpZIygS4zhOFJXb2+aRCfm8kg9bnZOH10L52mpYgSlu7PSiU0y
q9Gf6tBQTVweJxhPOmV+8Vc5RGN466rEfXogAwxSzMPXyxBcx7zpuS+3fj7GNPz3
0fL9tKkHgoE6bjvWTBR+69uAggBTlWkSYvHUzAMfOUaUCzqQpMsxN7h421yuoWvQ
NuVxP7SFdif1Prdmmn8J1hzNBSXsrAxf16kVp02an4MymRp9glhg/h+G43uBInN1
fKUHnamL8s8q+fiVMCKlBF61SKd85oOohz21489SjhhhRIzs68TWgM+nsx7ioDpe
I32ZF1LcZCAW3sxQbrYE44cgKq2D5XlLjI4haFGalouEXwEid21AUAUxqvEYUouZ
3Rflonsj3tISThelNWpiOzJXFU4w5bz9uXvJLga2zwVCd1/xrA6/mgORdqcKbNX8
FwTJGfUw4wDBoSbOwZyruJJ3DA9w8nQjRk3tsgfMTr+nPkvLO04CkxVN/dwOevaC
8xIFk5zWG6vQMqeWIi0WVDcwm/nyl4yncubf70fnZiin5LID5fIw5SxQXKcWRcG6
WZlvO0CykHbBtqaRgM9tKcL8f4CptLB1fKlXkWqBo3Tw0yqV/riHHO0P9orCZVuo
4VJ57IlICfPqMqPq5I3amtFG27D5z5X4SNdehEj8dRVTocNxtTNRD0Wx2KK7P9ZD
Vbk2j+GZ8XV4fnhfvvkGagC/XcbjJdgKLtSXtbsYNadzG7hkxiCAgrq7P7BimoUA
inWTihsZngQ2MKB296T6X2JSTWx+jVehjVHgjG50awNY+bI2KtVs3g+o277I2K/2
FshVVlEkBS0DHirlZBlq0AiEkoO9JRGeveqgKpzgJpogPiINUwyKbwnsfW5oFFLP
cHbJY3dvjhL9oOnZzv71gQysTX2r9jdKLMzI8bjtYkltzT6T/A5DVFprkvbaQl66
9BIvjDWJqDR6eibZ5n4DSivNi30cBjr58EPsDpF3y4XiQhTUphZOY7C9WXfxSDal
XkaLBlimtTckMeDDOh7CpBUUrQL21RquPw73guKhrlQ0po3fb9ElfdAt150kO8vJ
NYnv4JXLvVsGgkGfwLDRpJ0v4681dMGwJXNYQTjwC/kZiQXBVN0aBLi8MAO0rdxK
/VVWKGhS91AFqxL8m9s5K9ffWJGiJ5kYkPV6Wl2fdvxXDcJUelrNzOh/IT0GhdpB
Op0VSEtO9Gw5yPGf30EAl6wcH2rOPRxV+ZYz7HIeIEH4t74pmFeffvy9bZOxO9oN
C/VZhUHF2v/v+pbGOpDtEC6CrvaKJFZ+bJN1vyM1txNxkwLa1JpKTdrxWsUlc66+
FVeDzxDQ5znC4qBKLQnrP1P8pGNdEvQkZQnBMqAUzzk099veKK/bgQDH7Z7EbSk+
a/Kk5U6IlblmJTdltYPYS4UhXXyDCJ7mkCdrG4ks7jmtRtkL4wkNGIu9NJKcx5II
O0eJpBuZ3R1eI2uKf/aAW9jgOJlFcMEaiTdZftNiUQNiijIYjxi42+ZZSo2dMMPk
uw7syO6DOEtxdfhJ0BrAd+rzJoRXTHgjJX2Eu9MJsh7XlmslSck2S2MYkHI68f2y
V+S+lQgSHLiWq1NlvR1xpoijDtnJE3/lxyIvNVC1DhL+fpjaYEsjUr0A4GNSuMXj
gQXXMWVSFoLmRnjmlTbZqLfJtL37LlwJrjcl2H/FFQkJAdgLP/wzDLWbi3w0U+nu
/4FHdnTezbG7wGC6gGc8YlXH2gw2P1jrouULM1xcCu02Kcmxq92vsHQKfrBRQ1Wx
a+vB87OS1nrb+y/G3XCxUX45J8VcGde+I4r8Pdn6GbLdEiJDG3jkFQHRRvdfXkZs
mYJGrktgDpP7NfsQOwkNMcEQcd4um4ba8MQMmzE4a2tdPlr76HZputVWsaJRE5j9
BqO1HOvvBycanSMUkwbrWozaJyd8ZgXOoV6iNjB9qXsyjz9h/myIuM8r4NdQuzJs
OsJ5RcmBXleeBXzyysSYtG7hEb9lOw6e+KwEktK3D/BHGmsUPVqtypyYY4L6Y88k
NNMH8MbkezRek4bDu9u56l+BgG3cRuNSZGWwBLv+wONSywu4HysgoodusXZy9qAs
Bm1xOIhOYWfYFtX2Q9SDe3lt9Y2bm9bO7WmDyYK956ojfQTz5PrCYCPeY5tck83z
BY6IuSKiqqh8TBBGvKOsdBqLrSa19PX0TPRs++TbhQQIJmPvxywyGQq2B62Sipyo
pQZIBPUo8geHSLuohHcmH3lhEYnFO92anEvF1wCHZMyPhRS9qt6XlLmfY+T5Rm7x
Fn+xmKfom7xU1iU/SI1Hs1SxR41XoopSjFCLmtE+fiW1l+atSNksP4zS6reyZWFr
gSY4igGqyZMnc3e5EVYbhIOsbRI1jEGG38NCkAO4f1Jz67VmH62QRX9ldVMB9GEm
ZdjXAJ8/L+Fe7aj3mKohB51TAfQuRZ0Q3GAP7BjDM1rYzCTNrPLowEcBSwxSrwNG
fBf72gasaSyVqTs8mQvpZ658VjYzE4NRaPPZtU1AHqxIcerSB/Zf0iIn5e7GlJKA
E84RhfI3Dc9JS1TRjksuL/iUI74W2sTpnFKXdVcgwVlYuW34DW9BGiRQzX6XHWAX
tbLYujtdeSFB1DPT96+1cpdOvrqbTJJZZFWUozf2rjoQlBh+Tgxl5zzENrNNRZwu
LreMphKPD+SY2EZr6k3Gy+PznzGw5oDaQEgj+IfpCmrlh66qcDWXBnR+V5BLalup
d30MwtutNG3bxGgWVgd2z3yUBMN2TwHPpIzMnqMoJJWvUHM6QdGhSlpoA6sj0yPJ
55idiLiEyaMlPSmrr7ZOodNTwHwv6I2MCFi07KtnMpumJ5swSO//MkLWK1TFYk7K
kwU2TGL7Iy5sKkMqwRs+HLPu0tCVhnv+C/5VEDvpwET6pxZvHR95bfa9T3HOm879
7Bo+m/GMqk725PGfxbqD0WcRtj3KHZt/egxJxArgssHoaATbsVjlw4OURDyP2kAP
s+LLaeWDNeAcnt9vd1/aRie3bJWYMe0L5gv+wccEQmw/k6qU9mUhfyWtc4HxYApZ
YwjpCrtkyQt0F/K3l7co3Vz3YPupZVslTS5QHJvcgWPfFiVnaz9WuquUtmdaeTF3
dTMPERYcKSOcstlOquEEFeNp7fbAvYl3ycLPCCQdIezDxP2JPyr0GPtIGx0yKqbL
2fXrq5WkdTqVDsBfLPeg6kAkgyLXRnWmhSKUVzcNL9gGE1xVUCls3X6hfWQwZHls
BZkISeE7jzzKx+qs+OKYz/YUXJb758gRGqwjlTuBiOi64/ihW8tO6X/hKw+bckpP
rt8yLFeyxDhDPVdTlt4CqeQKPhgWUIwL+5bHowy4wNKE1EN1QvM5ZH650G9g7RTW
hc5NpohLD0mjNEViPaCve+u9sqtuVT6OruOMHDWrj99Ert79s5Wo0sdpHUIrjydj
31E1QsBOqF8jU4m6o7HAJRmKosnbHh0rYNGK8u5mo1OynBXNdnrTzte/u58swzqV
BcnspaR1+nuIAqCC0P8cavkXsrIkfMVaQ/xMk4whOXxGbGVjpbg2iHKdfv/WL2G7
w0BEGCxEKRt/sOcdwB5bUKxdGqdeSEawAptiNruGyXNhsBJa8JLXlUZa3sFOdZjp
5DCxxGoAmLtBNEf3lDtOnCBVPz2JV9knfy4KP2aZE69iCWGNkqY0W5LHB7u3kKfI
BDGK3MWgRCg6NnUzvSlfuR3eOth0WEd1u2hdNJxcMGABjzp7QWWNyMgzuKYMT9+4
2ZCFxUKgpXzL4+nzFuNdbgih/eePzB6MSRoX0+MmcFHSMTD3PmXi3yavSqbYP91j
cfHywNRHgVO9z4uPFlaa6YIgLsNXky/nBx90oRYQHI/CFcxuBTI2VCqEPEWH5Np8
m8FbS50sdO9iXL2+xpcoV8+/8UlI9oQz2uwH8a0Jd36tY3Kdi4fyhGKB40AFP/lh
mm+6z6p58Ovzw/eJhcthfq5LzNgIAy6qNaJ+6KVkpQetjJmwAQmcJ/fUfUW27WBu
aT8dFfxu9RegiOfoo7I7FRn8/v4cmoyKeNLBZrbPzCbm9zCoH2G3M4b5xyCij9Fo
LQny32Wqo5ESG4+CA3JvwwJ9MPcgFYD1gCeL0w2pBpgvFWhKk5w9sWTzR79ISBQ5
CPe40K5vhfpYnvOUvAkp6fcX4NHMLQlfAvgP5XS/23F6//3QgetR+vvkX4X67xyY
1Ko7+7V07/JEKf7kG5ZiwIpPvqV54Eml0NyHGjuP+ojF1cA3m123Tjq+atM0NvkY
fjxRxVZjlKrR/h2eFYfyZUr4dPUb3R95HrHShqrr7u0cgKiMgNaQ6+tl5EMlWhwb
bKotjeiVF8EpmJ8jS9dUyYRZ6mIKsMtRhYy60bxas5cEQOEPvWF/6qxMB4TsYxB1
3LV/frUOkxBY/0Bw6/++eVSmhDotxGUHsWfYF2YIQ9sVPHJ/Y4LsCYJuqTAJ7IlI
SvJvU94w3dwMSjkSII1knfIEPj1suKcqqcQerWT57XAJMmpbv1u3ekxzukonykXG
hnqWLWoxAnn3N9LyyMkfMZkoqvlYKOmqpwZaDPnEv/Iy6r3lArJxELT0E0kHnd8F
S6S8euJuS0YIW1H7/lY0lgr2SpEDTAibdvoNDp4qzOBGZ8BA+6bmil+teTDZb/oE
abEYtUX0xbTITnbeHU7c85++neAiKF5QC4rguONdLbstxmZdfXODCrYt56pFf26n
QWOYOuuzP3c5+fHcHUWnNEXI2AmkhdOdgcxt33OdddnD5sDUUIeBNu+8HbbSVYku
jJxfm9XEGOhAyxcBWU2TveuyFxjabmpesSwPd0k2B6iBX/ycV9Lgxu90H5OjmX1m
G5mQ/Y42XtBlFyNlCYmBOCIkCn6XCWk6YR+Q3VAje208qAUJKiZ4Bo+gWCnaQSNB
WRUwA52rR/q18TN1D9fwZtXEc7CQD5EradvcpVNBA/vjbSdlfJncWy6No2PG9oHP
lfLmbqgt1yypBoIitsarYsiJLsGURmU3J2KagK/WcuXApeAgtgdbC6IQPTKyxL+1
XDbycfsxbvThvgF8iBofj8cC73w6f+jLfzyr/Ou4ayyEIRLE1TgJMR6d4AwjpcWg
Kj2wQ3HTB6YT2hzNEONczsgz7Qr2m5c3s2VpE87t5Op007Uu44+eH8z5nseedHTs
9NtOiA0pexqASZ/uXee8okbYXClL2Y8m3IAqxeeLsn5YKbO3UpFgLpPkOLp/q9Ar
Ti1nQxJDYNhuk63s0ZYrRoexTqvfn0t4D4FBZVifdrUYDXyfMakIc+8FIKKyg4R3
BERK6Ofq0rWoJ3TP4miilOwG1MRJpAPKXC2Jq6vai+4dVYq+tL9YU+hPX0pQo8pR
vmb1PPVjh4SXnrk5umffZI43yH+k8U/Gv+YJ/xg7SOTTVPQHINiHMf7nK0tuxEH9
Cn+b4er1ulzMjyWFn5jXA6bFEYdyuyHLtK7SL8U1gtQgGn7WphoPVlvgaWaDSoZt
AztAaAYkip5Br93rH9NHeJQMpCTidUz7BG67O+tJckTo3cQsG6dyc04MRZVNVyv+
a/hrh9RR19RB0I13Ylc7et4ojM8BLYfsUX+LPIFc3lVwN5JrD96NXlYms1fRlHlQ
fxo4I3Q6+Dc11zXnAVsIlxatny2jw3+uaopfpmxOSJBWdRa/H49gs+EohBk8TScZ
Icc2w4D+GzxMC0v97p4z19fIZ6fU+LJ9ORdck7J8Xb/sZ53yUoc29yR2fSJy8E5e
A0KMCT52rbmalMbE7mykYQu/5UsOhXRfd9D6aYaxs04lgz3rNiAbYik11C5tUo3E
4260qus9pTPMHwZHELZ7n92KYPrA7exma6Iu4MxmRQQKoVPR1XgoocoAz6Awbuym
tLwXhfLqGAKBd+cSKBGEH0gxj5KfTvpuTfPBWutm6RRMVc73N4T5RhLulbZjf1jC
4v64/ZyYR1TjRzCL4sVFoKXQqBUNUxY3cA7yRSyi04Dr7dv69+Y3+ZtA+T+mXFil
J0ayoyk8d+f6YYVzJputj0YMl0LMq8HXj7ahfAKyVvBj0ebuX10zGK4/zCh+XoTr
1GpIPs5Cs5m6qOBTe8SBgfjUh/ImoKCAQFka78ekhGc3Zm1LbVnZvOa3LfF4Esom
LCgV+43goFWYfoVyucpztpcJ+dZ8eOXeQH4Z+pnm+hZtEZPNEphypJLQH3iB8Pwu
2UIxN3yQB18pvpIGvanMV/OOcZi/G+npVnsKL/WvgwH32PyMy0++VeiMnxEB5MKP
NClUNq2Fdp+cJUqKmk+jlrXerDd84G2apARTM71dQa+EoGitFdytfhTr4cSlegFZ
nkR4Ytek3L6iRyHdCPPUQtth/GqdWJE/rMoqT9NZgTBFDm3pInDo8ZtV0gvgm2zG
hwcVAujyocRFaf2t5PPTlUTBQG6Wn/LIk5lnvrGjH2ke6gvfqxYoMPob+F0pd0Yx
f/AlI5An0RKH2pu8rQgp4NyaeE4Szi/RVZi2UrjbVMweKZDqcF5GIPBUS4d1LYEi
OYhfx7xhf0ShB7qmjoaPxYLKKWkqLlJ6ysWf+IOaLI0mMqruvAMO9pZHTHMraADZ
9RVNm09Ln+zHIJB+vYsHGEJc4+q6y2/qLcvWchkOOVQ50qm6bLNTrHY59yk6TZYB
ibFaSpEjnVZ3aPR7LHmRMfDFuyDopQuEp7b6VxuBswCoHIq+wvH6iA/E/WMxr12N
MKJWvYB4GwlrgC9kkpISstYdzSeSBv/HwfyedF8MBUvk2kjypOY8wecgpI+XnNaz
47U1gMYzxjt8z+n10Cr6/BZrQg/iBdb2m2RZJP+4dS61+L0EGIXIdunDrPL6gJ5m
zA4q7dqusP9zSv6EeAaLV33AhgDbUTEWyXCNrKur8X/5TzuYB9M9WNY4318RJT1+
/AEzGssiU4KPThnspo35PGnWaNjgk16Idcwbb92HJ8A+TkXxNtDMQpXk+nUaxGfE
nxQ/vodcl96uSaQ/VlpFkkFD040fGYkILIuLppZRJgIspsTa/i4GNnO0/AFk9l8I
WDrzbfcZuDmtoGcCjMeHsq/XQyJ8/LS72jUzrE70B9wq58GJnugw+zQaiJ8X/8CN
g9jBf1RRSY0f/2Ayq/p3rQ94cdO8L+RgZ8ruNQl80jweuSaBGW3QS86kCrkdqpfa
Kw9x+wIQmp8fTtqaVTZz4BVh2bU8GcUPmccm3OXbm1hoCm5SOJ3GVYGN8EB8sbBU
/fzvhrx+JhXYe/b9dDP9nqFqMwLFNKZHFYlaiDKmm1bwjj1EPYThsojGlnamSgBm
Fck/bfefJPvRMD7mhESGuIK1U7dajMgVQMNXUPqN4a3EtQPzXwPtl7ufHlLypeIJ
9Mtr8YBIB6qbkMiiNpGEFO5RrRTSLKaCWer9NfNqVjBCrJMflXd2/sMJuS3+LJJB
hzSnTgDWrqMyRuKaQb+jFSlROy3GkDsZwLdkPieMFdWn8D0ioLNtl9RgD3rdeQfR
aDwQEQcSk/3F5bty03zFxvx55wx8s1fzkDqQ0a1hXZp5Z/oEeEVocA+2Bu2NNoQz
12tyJ9MSD438L+Jy/Y7iZ5bcUy0tS4lMVw4sJgvGsTxNFVNCmdF8IrdVLx20Iykh
KSVrUTgPQY4nV04PSip/PSbZa8sYL95Xyth2PrBOygP/vpV6Q4fVDosPFJ+xBi3G
EestX8oWNe8J/7MQxg9k14wc+SCEzfcugAF/jOJVFCc3ZngkeSV4Ssqx3FYMkOw1
myIVdERw1rx8me5pGApQAYcZBJSbgdWk9PGPtIvMVHQ1Srdi+C9Mgg/13Ek+OBT4
McjlnVn4SZopdbq0za6k3mnB2vEJXoU2cUGJDjAfEz3XeTPbwVvdnszRoh+rDXbW
ybyza4HMH8aQFcIWhxJSzI3TCE2B5MML3G3UqWbRs4ydkHRldLAxai3B0ufr5e8e
5GfwRcF3UPqDgSLw+dpJ5rwYAXlquS2LC1d1IPjRknRfJkFPLIuyWCmVXUQkGwf1
sISG54SmPkE6VdEqrOeHreqSI/qkoLmpuoa/mVplWQguXbfEc3njkPNRI4SCWfKE
o8Y5av2yeH8Z0d9Zr0t9V0vFqAYQwwpPC483xkW/rq516WF2fg9iZ+t8EN/DafAd
bSs1/QK5eWD2oMi8+bH9f+A0Sy+FtI3hV3RukFKnjLeojp9AsjVU3+TMwFV56QCh
2+cHquxO0+1bpiD+g85ENu9nM7SL7jA7ATkk4i3sTpm8OIABqvSTfgHJFkxL0rlW
SzyO3rUGesVvef57kvH2pZccxMko2kpBGi6YL2FGnb22SOINB6LjifzvzORh5zKS
Nze/FOPzNJk3N6YNIeQ8jS9/B8miB0vA7/+wAVqSz63mq3ymX5HKVnAG+ZZZev2Q
PBa5TkYwUrQ7ybifF3hMvBgwxq8qCWFAMuunyxVEGbmIiIw1FG1pkMOixXkpnP+G
z51Im50DNo+GoA3tyDyOpvZpKbWV1kALBvjWK/Ud+Ic1r5vSKW6eL18JFs5ClB9G
G5BLQXpjcwlmuvGl2PxJSjuKsXQTT03AhlqRsRDQSb77ZAnwOPLJ+6pMHGLHevCK
xjg6ezv7KtIbitqoIu5ro78FkWolzgAtq3DMoCO18EIhuDEbDomlQyolRoga0nZR
bA350FIiVgtY9aR3XXN366mEJMsi+riC3v7ZitYFjodcWoshKrouBx8pw9Ic+gsQ
dlOs1/j9sI/aUuptO5RoevHNtC2jM7apfMdr1viSSibbIxYhaDKmIR7eja2CyMg6
oHR4lwm5jKvsUaWw77XyawTxhUYfE4O/AkWixWk+DVaZkfByHNZwQtC0kSuw6ARH
W9jADOelhFsmtJJVqsmqIO3GF/XkJLdSgp0noCa1X8++pPBshMqDqUHkNUNmMHO+
RQ2v/NciGK65SaGAbS/FICBANFixF4MK7rOkB179D12j+yG3ZyPjtqp0zWWQg5lE
mKFBIAlI2F5YUUlz4Ftd8hKuqYJfX1IY4M3n7mYgZ4y2U2fS+8tIc1gtQbC6GBOj
G1jL9Y2+sL6j24OB0yaZUIGIf7ixILLG9Sc5d/etu3trZsL0fHswhNWm04GdB+eE
XlJdiXG9NimLSAAN15czl2n10gzMhW7R5blGrbQuFBwTvDDRMChNOKT2F95gZgFv
osRR5CxIDuR9CZ1gCTV9rLbLmdsN6IuLdhg3f2t7Wvs7BQOjRib3OuqQFaUZhtcC
9RVBwGHVjfiaHng2aHSYXhDLrd35PkRpglq964rlWtLm2pZLH7+8IX1cQri7WsBB
o8TGW/GZVCgZghvfaDOBx2DYRayG2NLzwHyJVRsR684lY6s6wvfrQhUZKYvp3LA6
ofhWgzxnIrvLwPWMXV2scXnoDu37zF2mJp28s5X6jeIdvYmiXBnndE4TCFezojfr
lNujH3Sxujm+TNkZKPdGbnnieEujyB0lhOltrQYlj0AHxhIQTt/KKGOEscJbVNFO
u3nuNpBBERvridpEy1K4tqug9V1n9wtwLXxIEeX16+XwxH7gLsyqeEa2jYqWUr/P
JZjy+Ccsk1JN8lTO3SwzxKHckDTmAWovZ3L3N2KA0c/0rkhZkBNTL3fF4E/ZaEcK
tQ/A+rtzDy0IlwdQC+0VynTVKICb3+G0jBDYoEIVQldp2Jm/TNyMYTexQWSuxvwr
6h8gZHS5L2+ElwEUx5M6qQcSCXeF8FbRSknjv6IMkywl+tTAvWLMOw2y1xuIajSg
6wTU32Vm9SfNjWxbiin2ySrKhueSiVl8npZJvJt+eKpU2iOoJiZwBqe2JuYx1Fc7
2wvVoqhWbCXN/Y8SA3LH6+VircmAIjd47D/0momIP+gY/ARVZ57MlV7J1MsDkVsG
vj04kgIfpK5/UblV2/z5ihhdZ2lYqo5PAfWKRdgqJGeYKHP9acIng8lPvzY+GgiD
Fym2aVyjuhnfhmU6Y4Q2mv77vPvRPT8NBWVpEinTF6K3arZHvqoYxin0mmJQ2CD2
x3HhHzmben6PoK0A8sh/P7N4X0G2BSDsdDmn5m20Zm07Pco5Gr90wWAa25G/0hkt
TNJ6Gvr+Q/lMNEo8t0tK2SdbSyky39ZrzL1ry23mN7bikL0Po0lh1167JtJ+0XOl
nW/SymmDqCgVLWmzMMmH3YqRo73iH6q6Gjrtjwjzad8tmfL//SE6Ew0vHvM0e0NC
VtIR6uD7Vw/6Ib2SH5Q1FjQxEtBR9es1iyXtenjfcuhbbYnzTPbeA1jMn2GP0+Hp
lFQrOLKcmnik3eZiNlM7AALzR1jdKpgSC8hflRiHpmynHRpzuiuMUZmf3VRP1/s+
FmrCA+PXYaFAZvtE93Z2/oStZajNv9+bhH6htZXhDZBKcegcKvDtHdB6yEa0cD0v
klZ84XuZoN3frgWK5cLKTksFt7leVdqaJj8UXrTHkHg5jI+5RlkwM5sjKGCPr15z
OFIffHCJIlYm25AAeyroOufjseBHv2rmVCSrJ34EGcdyA2ln/kW6iyRGI070b801
J6PGm6zZVZRyoOWYBN/tnQbvCUlVp9/GdZACevOVRR/2NZcSSsgpM09GbbNqrx+H
wwtNR1pFDf3Pqc4xriEE+iufdAVCVq4KZcR4KsluT/ZToI1jyR0PYqbGUrCCN1e8
476oJDhjtRV2HhHHJ+QtjFGmw1dAHONZgJs2yUjjsX+Sq6ZLQS847GDiq+g/+Hwu
b5bYghuKxymQOdYT9dBmMpvXtoq4y1BkAT6rbJlY7LoiNjoN5Vfpz7721nY7MM3/
kF69Xw9Ua0wf+famQ01B+0HyAiqtrlA20cYV+PcP4KKHHLDjOWKHESj3U/xaf1lD
y5M+KGRxihSfDVRocuOPDSorPSEyhAzA5ml0plC293i3v73XxwP+gZxmIibF7Gc+
n+GppUB/uO8EHKOui05l+A2TPZTzwSx+TwynKa+EsrLMJMl7NxNhUnFxurklFKCQ
LasXbmrHUX/XDjaWGNVjzY3CLGbVY0kmNI7FnxSuxwZeByyQfJ5uYl7W0mjpi5o4
huxKP/NC+QKShPECYKilODBg2n2cCcuqptoK8jYU20YXvkjV3AfE49+z22AzthCY
mNrQKrUq15dE6E0eSKtKPkC64JCdZBv8TyMZb3JWD3daZamQmQ7jopk8XTCGeSIO
i1etamSjPFZvqYE2V1Av6dAFn+ovIYu/AymJ25W3wz47sVPrEEe5wBs/REqmiPXr
N6weBKvn9vPGmSSGvpQMs7L8AUoqthaHIk1qrzvcCUeaGUQaqZi5yCGmmE8204wS
KGgE8YKon4sdlUR24zfVOdP0mmlk3BA19UhkNrfrcGsZy4GMHjJoOepUuW3+RAzb
wmkBXA09XPULvZ+7BKM88AAEoXgvgAs7fWYHPDPnp4N49+QfIdwgyAFt4ouTaXwi
rmQ0F4+PWy29cmOtwKmiM+tse/7RYEbWW4kN25A/AhIrqZurcfQJTq+PG8VXcyIO
CM9tPpHvZFhhivRXMhxPF5NlYGrwMdFcuBQp47AvWW9un+Iwd+pIAUCgO8QYu5ZM
BueDIACf0aTZ5hFNUjNk9leY1RWNZ/flFb4gviF/KBbyNoJkebWfkKNYxgQJ3JY0
MVrItR8f+BfnMHxEynTTRWnMOQrpw7Goh5DVvVbUPBJaFCPXIIEiP4P6/FHcxGjo
KGuyXkN8MSWzdRlbdqib7ddeDy6b1/cdQff4Eu14Q0LlnZtI0KVXaWjRLRd+xpnv
Cui5DewTrrYx6CeuLr9eRefDUvSxGS992v9xy7Zy0K2l/aD3QkDgNhFX1sVTlqzh
13Vbi5dgGtFxBm764wyX42nHogrUeLDqzxpEFFgy9M39suSUlk/UTeTo6ed1Mehw
Myb43tisXs+o5tAhEynC69IhBMxaG2NNA4AzT+ce4MWqJmE2HLu1xXQV9OFVYWun
CmH9wvjYYAtockCKH7G4o6TqELv6qjck07NvmB3sOZMeqMcrFGm0/hebWTTmH3lq
7HLL0F+4UUwmavgCJrceZ2U0cpq6JvbzCKT2MlUb+5H9Yyf7RUt0BnH5JznYnnzj
vFUMLEJzNjuApk321yM5C4DgTsDcUaZRIm2MUrUGV97qtjcVWUtwfTLVtAXnPmkM
iKeiPhQM++9B+VYadesxYTd78SLHKjao5fRdHz/FnNwMkLeHuRrE4G3Z/OMHQ6Nk
GRsjj2uoxzFQTkB67P/Nw/8v8kURVApAQtBDdLHVvYxHKMU+JssBDwfYZ80j389W
QxN02Uow3+9Uvqh9ZQlXzaIYnT3Ny8QGnvYEbNWm5i10wwAiyX+MdDBu87E0Gj8D
t7ZPoUS3Jz8cQoEwKIgSY155ZuAP2YH0XCAxclddxF5cQinf2MhpQPyMh3Ugguqs
iwxo7MlD/EtAq5G811drW/y/7HmjmM4wgyYrT6DAtm7sDzJef/yreM00fvnQOCu0
HdZ697P1ZuufiLoFhLvN45g8RpynSNMFAQv7xDGs/i3yybI1Akk6XJjL6ZYT2BYK
7du8CinEhTHwgSaSnBsEYA82Io6hrKBdgmVl6Idu75KmO4xDoUR6GJH4rLECsQbP
isEWZAhuJvAWFU+OD1SSoacEeQIhJ6CssUWDK2kwioKtRhU8FQ52S64taHENwTog
MNu40Q+JPHWiVuWB4S3XkW4spd1prvOkknJ7rqxI+lMiVWtY5XQxem5jW5Fhs83C
FH4mCQY9DPQbZ7t6zaTved+alrHHiMo2VxrkJzo5DZGrlRbHKibrWay9wWnRZdwZ
8oGsNT/B+n/UYbmFrWboTRUAS44O+CNNOGaL/nRYvairTIdcs5QuMwbe7iIoKV5m
grDBFsr14DB/XOXwx20hYMKrWxV9gmsl2MiBVWpPTrMOyxaaR1d6Uh3BorWqgXJ2
qd4faHTxGC3n4ykIQAGvhssXNhqDWAezNSz7OVvEzS7BQyIKph/AEYBkBvmo6nga
xl6K7P2iEwepdDwgRPZN6eKpJgjeplkHq3DOkrgFqLIsIsExHChG6NS/DDYE4g/G
3BzVJ1hUbnP1goIoWdYQOv/5OjQKGBJwHSmtGE0qPtkkbfY2zngPiMcBsOkg7RLa
W4ssQYurfiqZRhnO+ViJKNeWuHtKiATarSL2zVV4YmuwE6XPRMdP4MeR1TeavSEZ
pfQWcR95UjiIPzdXEMqa5ROh4M2gvwF266bpe7ka6K5kg5VdaVOtwtoCRUDPRXrA
+BU9WCQphnJETznT2WB43o0jGvLgRuNBkvKwaEud3OTCvEKuZA9vlZwLG2VOKq4A
qp9S9TKq/5JyWtQoZsoODFUCRFRlHmzQkL3Zm8S94RcXrdCCnj/SVkXaPfia2xMG
FNC2NaVHENlMQ1PfDdOfxOH4q9RT7/1/GTWM5xHcbR2Hz/0XIuim1oS75gHZubZR
EhCWQnAiMTZDk7UhHUMzRI1bLke5ALZOX9AUB8NDwSskMCCP0pTWyyI80IoZ4yka
eAnUWmhwIJf5+vRn1ixGkwTJGnbZqkMjbmzEAI7kntHDC9niOoJ37ffL0wmmJgKh
AbQbMGDDJqJJ6A8lnpE49weILcccVbehg5WqLwuFaBYaXQa9bjnN/WlKKDUekge4
28EihErxY7LIhGJumhY1wEoBMg4IOhrTMSKW72y3tHIJsvk8aHGiNXNeb2Gxo4bN
NcgHitwCsOL1XIfiBAUKVd0SVc0M0RpfrclfEfhfYP7Te1+hCHFPpVYF1Ufirnz5
j9tR4cT85BXgRo8zRaaaCxzmd5JQlD8CP1CoNgHFAOr0AHuVyNGMqwUK1HHz9YMx
0NQuTVP9pMPywM4m9JgV9pU5jnWLYsKVxPwNSKiDnUkL3TZKIbaTPWNv7nTAtThh
s6GnO35EeP79MdGgpI5m1ABfzxbFEYWVmv9hFLgRmPhSeN5h8ZdrcvwjnBiHI5Sn
BWNliyl+h861HaASHrBnW1BODgB3uH0g5VObc+RwJXbzk+Cir8LaDWuZhJ8ITXVT
ma6MEdb4n11Z8ZjTz84Z1JJTDb+k7w9GhkJuPrI2Rgc+BT8tqCJ4EC0l46RW8rY8
SVQYyXjYTMeOnp3NUz68pM+zcjI5FMFS1zkb3mYDXrTYT/5I4hCceuemGdf46Okf
lfajpAcRNUXLgjlU7fAmR1Xq40R4Tw8Fu8qSGmrO+rVfFG3jwGMSy1EEQrvU4our
jOW4TIHw3m/oESiJDV8TniupDBXo01aprqsXjTbzTfE4WgqwfOPHw88HXrs65C6i
02NEAnVuEwg0qv+a9oRYT+wtny6Ww4I1j5vWscn6cYcCVBlap3GLXhxRJZL8PEye
etxJqBcWcuR0P7gsZS03bo0C3f9yqwCBXA2KjTQDAxc0m+2TfWTDg0VLuJmqnkWp
genZcsQCbkmPoW4mpsrBSlj0DAm/XVASOClmY3MblaJcFm80/0tPasteTLG/ZjTY
PUvPmFUtfG/GovHXdCdh8iew9WClgymiq3CuWaOe8xj8NNwEYYNrZKwbHj1mdkhL
ot6GmVFN0gN6ad/DEpjQVycu1zEDsCNKddYwPcgz0mJU9FUdiDcn9vVG5ieEGWwM
qYJwieD9mLx6fRrgH2GqVNHWFHKj34tcRSw0X8n9kZgA+P2rysCFWqoxqC8x2k13
YbgerWhxYX8vZLLBbLqMkih4Upvn7uVHdHQDPyJdWQ/TUTKkV9fwANIDelhd8KNY
cCR6bygcdtfEiSd6zOcsvUV2i7jGYCu6CjdR5mZobTAszv9KuoLbEZrYKDTVWtRN
4prqjyYaaaejtiuWWxfCJl1aT7RBa2RTGZCHVTG80HfWmfdqoLQeW4GUhxkMRUzP
33v0NkT5sgXS1DYhfA6wcCyhOps97c32dFkFK12YNvv9O7S5UdhY9Lnz72z6thMF
tubCUjU8Jg6x91AqJ/d0wdTRFizrTIhky6caudGElFG+0yHR9h7S8ZteZ1NZlhub
k6k0VU+UViGupdYVPmQvJMC2kekbfbb9Rqv3co296ucgGT8WVVfDYTwtjwii2UYy
k2E2mW3Zm/2bm4C/ZpOGBffkEvhbLZscobKwrvwaQApxq9tuL9wrNZ+x0hsXQzbb
Npmwxovw87a27dNM3Ab1rH/7gA1/VtDh23Dzi3g28fVR2D5cZ3GPJbdQxnlImAZV
qrOEeJA2Ztydcl4bejI9J5ZhVtdR9H5nSl3iRhr9Kg1xhHMeuJGkl6yVPNWdZPeF
s65BS87q/U1rWV5XEp/ivvCLBJ+MUTRf3fDADYVzYLVMIL0PBO813QnFDIEe5bjL
+AEw8bLJaIM8XNDLtMz/PkHy0ajb85s3ylqHC6eeROypkmUcKqxjU7oOjdhzjV1j
UFJBQT9l4sWk9+0aEXxdK39j7bRaJ6bFzUCpcKPFTFqJ3zkWG9t8yZIqx0fgwf6p
kyWuyOPH5wsw8VyJOmbZxV/zzdo+pkIoOW+f++FwQ4hlBZ3qzflyLSVchc4Cn2HK
/jaCs/5FZlWCxNFmwANfZ3PxC1HCWW25CCLPbJ9vNhdDw/hYNMIpn+kWGpiRP/v/
eAg39GzesNGG7fvtdvmi5AQwbOP9reIj0qpRKDVQazlPxJHYMtc+eScB+5aAXQ6Z
fGYZ7OcKUPgwO0XGqX6cndwdSY5peLal5RL2CTjMg5b9fGsRBDqOfBaZJeDjqclQ
NvB0Az0QA9rdt8RIgi+tEQnGgw6hIRQLcxMRoIubfP8+JB5h0mwEJLr4mxZCwsPM
uLHdLcZG8tp7+qA1dTb16amQjesPh69Yh2O6BiDUOroLz3GZkvKj2wZrshwpIjn6
kqDrBoT3gJj0ZWUIwPQBCqXUeWVW0bnuecWALmsqGqENEuc8ofcBOF2lh4bl2hmc
m0gGt/uRArC844vOK+R4c9mS4Mqb/61sKnUzaQvmrAYIpj1HMIGd0pK/23YWEOfK
aQwmND9feDoR9ud6HbpHQNm7ISwqDnITCEo5cZSub9vsEOM+26kL1RnSSAiUe0IO
o1YOPxrTNWA89u8wbWG/142AZQCDDXj3KquEmA64pRby5nbJsLH6e9e6DQXfm8Mm
BIdg5JLuKlWLQQ8XeaylVio+W8GkO2nUNaNu5d/SvEUNLjBqyfyeqbIpsYZgtlKu
jiImFN8m8TokDz6xKPjLINB2bVpd59NGRJEqMjMmvhUEB1StiotyZ6rA3xnDUDqV
6S8+0f63ltQbaZzaWuqzyTYx/x2nfTuFskdyKs1B0YfFpt7aaVuqYOKJuWlPN/f2
BTi+lI1Gn5BM9xeOrb2IGZOD6/SSl2Q+qNUra60KuA2z/gzHhga4n7jOktqkuMBt
3PUgzUvqrDV47Fwe8SLYUacNzj4UFL4vXNf+NouByXuwoQBy3pqtJHUuAVcPUsFG
qr7SXFzhnwnrF/SV3VYxdeAf5xYOhl7rKLT3Jrt/8BC700K0sLS45T1OHocmkUES
OaBc2xnclz+O12jQ16CIXLO2HlaYzESal3F9+pkhFnUUo2UqJ8OdGWdq4CpoTwOJ
fLLWCuuNtF0xEWQJY+ZHmMoy0Vru2KtSbV8JrGARB5+AILRU1Sdh16Vf03/4b2cE
AOwZUZqUK6vKC1vq1E4+rX+YG8+zQqTv0mBR0JbtUCTQP1z/eD/nlB4Mxxw7LmN2
biqoIQq2hLKFZoZmC+jglHaxRgrrmHUwtWdIXAIJqwuYJPgREr6MSW61C/y4xv9/
38C27EEsjZbrObN4BHBzttuUMHye5XjGWvd7zZO2HUXklVORfhcsOPwc/iIFjKPX
NfIfLtWm+XmfP/k5AuP6hEkkTkVMTZdScOu+SUzXOVdduuB0uZSCLKbwTjdykvHV
hISBJwmuJxdGbAInObQBc+YQwyTRXkuenXUjAai4OVNX+ttan4HGlz5rgbMr9S2J
nD59h7IwhH42kQTCTGChG4kFUSxj9w+3JtSC/uHdtZkIVb7j4l/urK2euenEwT2u
gidZNba+hhTWMRgvA2yGlFbuFjW1p7m0uSoMKPFy3b0kaKKZfQp8hB9JsOikDBKg
rMHiPhWx7mKaC1nd27bbnJy+SCsIJBm1YatxRTOcJyL2GZhQbj/Dcz7ruM99SF8+
UwTl3B5sDFbW81dTiKEgjsYZXiLVURkC7/ZEmG6tDFcomMxnxgVF8VQUvnV5h6e3
Z6KOOppGitwDvActjS5nAwxzz9WhS6yK/upswIwK6fXRZXW6NpCLQZpGOESNu6QD
Ug1J7TNMwV7uKeZdiXEFHd6ltijEOcaYfq6zdme+o6vUaNbtPBOUI3hpG6vbCzcF
yHzeQjQMpjzvL0QcOGYvsz3jM7JoA3+dUZJ99JbN26++OKzmDohoF9rmbkb1cz5C
2KmEwOHUNSUe5YYYae45XlweBR10gRjJDbmoltNZ+ZA4vRqFIuE3F+Qxq0dS90Hu
aQxgFMv0CQVPLVywsX5xHwWRJtCu8AGSNdEsti5NP6b0wLlVz0A9+jskX/x4Bd4C
bf0BlBeQslqGvAB+YUrdw/odTGbSjBsYnEIgbSRVZ9Dj5ow/p11MUkPzqAs57a7r
CiIsrOb2T2PAjbVsFH9FsYkwE0Lsn0EUmTsFKXFYSgq+MWCrjkFMmrkboY/Pa9qm
6OyY9Kg0rj9w4Qd3vnK3QUIp/DpdGT5S25JpZwGsNZkPCt5nwS/G87aZOgXKJq35
rBRMRhB+XgQXxenLKMt10YP0U3dZOLkmqHipdw74oIdOhda2UeAdYFo0GTraxLee
iQY3Uedz4YrmOmFXyWSwr7LkSfj/X1lEmhzB+xotqcoh3CzMEpDErzwBMRw5lwK8
rs1CEnIaLlWwjIQh7jgpwPv0jv4WICGME1KMMX/qnD6eu8Ei6D0W0TTpQtvrdc2z
zHfwtcOfa9aFZeREBm9uFugzG/ISYqWfUd1nEgQZdIdR5BuQ330JJihdMgSdUaep
4RvQ7Ji6ethlZ4maOt+uDhF0XVq4kUhkExyy8q7laLI3+yAT1wxzRcRE8T6cNd7H
GQVvoyeGxxpiPtiMFaBclBiirJs9OZq6QQdUJZA1CznKxwcGUki8sxALFWZGBQ0z
KGMpXWI9znoyJljLc3rpQ+uYaRPQy93IKnzwmXrNwihhm5rq1p4SC+3cly2vzlPk
tIfIDh/s4P5z/Nn80GCTX47JgGzL+e4CwcstTmSEcax44bAZDycstQY4wqsNEBie
dj1+AiF6MbIXenb/yH16KK1LuzA2DXyHq3jblxPVnhTO6d6Rutcr/rr5Wo7XYr8/
V6N8/tT8JU2yYtkKtCfRZi6VWEIBWkrC7RVKtvmbQCNtol7+719LVUfbCZWMsKnZ
+o2RGRCZkRRoURqmO/S9RhBznJSBvwOr4QVlRhciShtWYqF+g83d/2VRS3j2W/v1
1+wX8v+gUfw1q31gJbQ433R7hZO+dyasga8mlQEsZV8sCc51AZwuJvYaQRttHiD7
W8znF0STxRnPkglkD82texDxATdTzdxJf47CDjP7kLgOUvVmAlxu1W0lAInc/cDq
pcBOmnRAUdYRVkph7ATKZt63rBYm20dJRNyFntfX56tfKzHkyiV6cv5rnrLUgLYa
pXEZprvKi8A2T1VVt5/+4SE7plho9PianR3goaGgrzQgBkIy/hFEmwNI1SRnwU69
UYY07VIgsLZKT+6M9nETObZZjccRyTvu0PJObkAg/cZF831bL2wedwLUcDkd+zWd
JCnOtuHq3A+5g/OquMa22AsEuLF7wtT2uV7C/7WTMPla3dGdzX+4qRTtsemA2A7Y
kOytu45D34/WcWAsQlU9V8l9gZ97DkDgnD0Le+8x0RAe5OpSyMERrQL/S5Hr4vTK
OHcEAqUzMz7qNMEF4sY8FzBkbs7eX9lFTAq2V9AEP1GyIhn2IFz6ocRdGhIBzPt7
37mX20VdWs78dw6Y6OrditEfOpIHZisqhNcjsfTOCt5pjpgjme3e+I91zm2iqVMT
a+ZdDoqfRC4nhp4t9xKTe2z+1J7GJGy0Qzn4/5T0TNtY0CZf78wzrmyj0ob0SpLr
HK4oUlCh8R/G7oHpwnL36766GNmwhjhGro/KdBAtWuQ0mvS9Rnfx9cU4kMWa8AKf
nSlpE9jf938fKSMnd16u33slPlEwz+OEGRpq4uyx31/HlMJ0570KuIeFTLcUNh0y
/91Ul3R0FT/fgaAa7gwe42mFxuUblER2paGT3cSdqLskkLNvz1VD1wlETHEbCVuP
Z8Xtp/HpTuNzleQ3o3TOQFCgG9LHmYRtQwjPAGqu3FJsOW64Kzn8h0dgC81q44Zq
JJ7xt09MplvRt5JxgMWuT1RSe/392zYOXXNDDKZBaVNgmznglw+0heV/uSwKVp7f
HJQti6PFpI3ZsbILO+Pubu20yiWduNgZxbpCznYE2T5qqod7DTexU6duU/+r59iY
DQ8PrGZnkgN1pobfK6Ge5/cdmoTgVyOxO7rldEIvefWvznwnatmiZrSV0zH4QhiI
m99EDJhk/jXXIACDi4W/dN1fkA2Hq4UpYk3UtQAm2VksSa+YfuIdFOErM3K2MW6z
RZda8kS91hX2A+D7N3xB9RsSTzhG3x/vyKCY9uvxfU2QFkoN5pjshuuYIhtW8Jmk
oxJE/l4PbTSqWYENkUbC5aIn7CToAhGSKcxQQL7NN6Xb9JtbojBreb2hG+i0atz2
NPNWcKG/THUAojJoXwglzYJiHOy+dyX1mRiAfWyaVB8juCxJECRMTQo5jn+RzPFL
vOVFa6869wWqcrSmBr1oSuqdP3U/BL7w8TcPdm5DsQ60jwnMbTEKsYDI+15KBBHY
HmeLUQav/lCvsGbleDGywKV+sF0F7+j3HWmLVcZ4g1+Pf1tzOl4kCdrV7ofwljUd
oVwmsYahgu4bbEdRt00y/dHEIKAwwP1WL8redXLROHEHIkxAPdnXrdKozxfkiTdk
yc0wc3inAiVl1BqpiNffWgvys+tdoPjTHdaNdwIMIS2ZmKzW4A2ThIqWr3Fc5TwR
u1o5ue1tz53PGArEE6vT6bF37gok9vOWwDrPY52z61cJj+j41BJ7d7suAxaf9XKI
dLzvwGoZ320ds5gbKL/jovhRzobYR4YEDxnlaZ1rP4JhzdpJT/26UwqUuJXcG5Lt
0ow+R85I5MvA6DYC8fDhWo07bvA677BUVzJAg1tRNMrYDcZ5nb6BygaaBQdJzNIs
4xZpuuOwC8Gp1VfEzGk451ponc8sFMEIx7qtWBtiPBuVLrb5FVVoSiy/UApxd4CG
rvtwHuPudvcEnsEFTEbVT23ToVqc1fbd+uBR/qp27Pxbaf82PevU3yNKsYauU0L7
+pf+cHPTJbc1CW98uKMKsjNDgqnNn4/uPFI56fZG4PmaR6dRLzE96pxHsiPDHhBU
ra1JDwW8KRoN53Ip8GlC420iCVSre8M1uSkemm07p/bp58eAgPWnE37pIwxwE19t
RO4Z1F9QW5519w1EQXfDmALqK1TGmSdNUTBKzXMdEnKxc9dV8VlNeqiCH0CaenED
vcBqwW8EPHx1txES71lunDNWmnA8oi3vItS33awg2Ive2b2WUsRFFp8ibnYm2akE
udws7L7tJ9X6RghRTUF+3t7Oa62CBs7wwXc1+Nbx++LEd9+9PYF6xsKfN98EPMxf
lQR6/CCMFxK2ZOjDR+V5ZUpB8bFfpKN26JVHDppLFVTVUE4NQvXVVuGUybqD+Yk2
u7zSB0ZG7QHlKRE9PfJJh8AjO8LAxOwZm+HgR30UVcOvvhtlqgA94gWlx7CQw81M
ATzz4r/wY4uli+A3SzXybCaPHcH3r7bcWx/2noHoWKNuDV2BF/jlJoRgRwXOSclE
Mgz72eFcCrwhwZXfB2WrYCVTgr16MnHjdrhq2y8dmLjcog4VI6mnG68ORKjlLQkO
0A2Z0aqq5IJmoF7Tb4dPwPckDOaBDrfQMutoyYesw7j1EpYrLnVrpFUlgWV8egl0
Dr5L0S1s2+nZETR+fpPG+5TytOlex0PAOqe9ITlGj+BgBLzhfFPTKooYl0zyXhdx
xJfeTSlQTeM3iaBx89iQmo5QcMEgFKP8QX9cn03QLHyq+dpR39XhxATmABWtNmPa
NlNJON9EC28xtXalHEDokoSXhAU8vW1tJk4om1T223hn9fHHElsLe9NaRgmXcltg
77PrA9KmuU1QUl+rslpAxgaz0iEGWRBCbJ107lUzjbu3YLc3KpXoncbWuAbyWvpP
vwtc65cxN/vo1XrDdXVtyQcU/FNgsZ8mte4bblx6u30Ho7XNq5iBFXU596GfDyXz
A36DSiCGio+ecvJjn6bfKoJUyRtjsvsoTXXHamiIp9LDoVotGEK9w/XXtwqWXBhS
I5D1USMxB2Ye1NGHtvPVDaARdUSE5H3IHeKDF5BN4WzHoebJRV7IIxAqo0GQBicH
jNeuXyiCok8RudfJtdwAS/fq2oyYcg5cRN53ukuT0rbky9w2VVeu8Wq3UjNNwrXM
OIl1Spy028ddc5IMfmtwU2jj5tr7ep52N0k3G7wl9iDD3mz4XRnn5W7IXgC31z5A
hUZjdRG6uIkg6jpSdnm7gdKanzbB5oRQoOA+/54R3hUmm3OGc5d7MA5ePSGSSpca
W3MPE4/7nAfe1lBM+f+m5zAiwL585g2pFtLP7PPfLukIONTHrHR/gEaMUwN6dF33
trWhCDY/mKEeOMBXmSGtapMTLEyAtgABu6VesGOHmSvhuCT+GscFKwZEfKHMmwtH
+wY01BsylFpqBI9LhC/AAaOCRi+k7J1B15GrdXTbn/fQ9WZy8lzzWXD+ysPg3KuE
W2i7kYLYI6uUDwbDeEM+RFGf50xyH+JTcYemMSKx7mHX2pdILmUsEILjvEpMBem3
nJBiB7wDIcqgz8TKNblWt1CbVOy9aY5yDwJ6CFyGj3ACARZZP9MaA2dRb1kB4bVC
8c2EkhZaNugWyTdDnkH1WsJGoZ3ENwjj62qlvTgH7cWZAfnIL8dPdaYCYcxnNiIO
b4wcPNrxOqiSw1FUCOwY2OXrHjgwPY3s+Kg1HO5Ulpsg3/QD1zzGad37RDBistzG
EJzVtHY19IWdfstimY3S3xSAIJj+aiBwvxRcKrnmCPHVr+3hfPj5tCbvBx7g3hP7
+DRqQ/JztGkaO4O+WygWPX51zUTk+9rabIe0GUEMMgu3K+NkP80udYN/BfXiIJy0
PV+2CN7l0+K64bvVfGQJvv0Sfs/wtzjGDdolzEOizonIx7WDfrp1sBPoAL6/9Dp+
AM1iVbm9JeJPS67TFdD2YfHtZopvQ5n+1UxKq0uaNluxnY/EHEpXpK9aEuSGAIpZ
x1xyQkNUgkUP/1TWdSUHhAk02JEp+OaDC6S46TD5TUUTAgsa2JnVEoR1AbIIRzek
/HAr9XTTh/OfZJhKGZ6Y2c5XB9t+wVbQKJdUFltkoOq2T62hz/enQSt79CZsNDfG
B/R/RqAXdF04xscUWghp2GRuG3pc8pX+I5Jnt1LQfbWX6gj6WgwUPEI653PjZ0Ma
j9ZBBQfQlWPqwH8mLRdPCBDNmO38ox2c4dyJwSOoC1jnDbIwqU1U00OSep5Ie7bZ
b1+PjLZKT10vIZhdctBts0a68+D5FegnBF2ET+kU0jb/19QXNnDJ/97HJTIa7jpf
SQNeT4lmEihf87XLjHYWFznioazdRe26iM6ZJT3wrtJ+j1jdXU28hlRlA4pdsFyK
DwDDmSkZrrObSmm9n8QmU/TQvsrXyt8RQBcQ/UmbqTtT6lcFyV3PB31oRxVHDdOM
RPX3WdF1Ps9Ej1JmZa5gs42yPpSARZgYsTN+7vAIFvn+TQACHqSxPmuEb3EoscwD
j4vYkqHPK8yL19Hnj6QTWffYVMMafJwJRyH7EImG+mfyzm4UJvPhXnbAyV7gt0mG
U1/DNKgVm3F0kCUGzQSD9tVRZyCYMCSG6t6CmiVSF7NHmqkuXvrqSOQF22S0l4DK
LM6YJ79YalXCrjiXWWCvSvrKh7z4nIkTZZTnSt6Z+KOF9saw0M6dkcwBeAZOeOOn
Si3bgfHIuLxE19fQbbES+aamWkgO9D+vI1TEOkXG2RV3xtI5KkfL6yOBHbKF7XTs
btK/Hj0FBaKewjtxn3HkXaqH5yajhphqznXsy5Az2a8jl1PCzx9z7fjHucRd1anZ
IAY9sn6SnMI6HvDmDasW+2s0onzPDHWK4ItkowNz2m90tH1L/IR5c6u1bCrBzUHS
ImlDQucr/tc59apGp6MJbmnb56cgz+Mr+b+rIIx+JuvH66zUIEg2a6Hy8BVaqzsy
40tcNQh0L25Y6NNsbE7gvgBQyHp47odB3fqZUK0uCsYOjDEoZCycvn0LxuKSZja3
m7ks/MtgmsgKbQDp8/z7OYMK24pVFJAZQn1unyNYHhV2Osjsm96XmCxS0J0HtzOI
8zI7HNnPerA1y665qtUNFb/2LN6LJQ0G7q2UQAiYgtGL5iavu/BQxGvzjuxo6fK3
XCB/POUx5EJVZqjbNNcEysauqqrI/CZtteOc9qqnluP0e23i5LDAJ40ozqMp7Dgg
L60N8ZyCiNg4q3EEvUttQoYQxzGSl+yQ1n4b2vm/3KYX/UlmbCkG+YvSn+ROLHbW
v8J0mWYrCcEbvmZJ/1RJXca6eiWYzPd6iu4U2GfVac7frIpUA/21KKUiJfyMOwR7
HOW1Hl0ecoelGOy9R8FPg8tosH33brVVbVJojgYOWsbYedt94ge6pWt5KvI0j3jD
J3JmcUoU8u4Bv5P0g8oMJhViJxRcn/Mkf25nwZmWU51IV40vzY6+2/4LnJvm2Q4n
DNHWCG384UfD52ghPjYwX8g9XXMOiEsRSkUcczx//834wqaWgvQQRL+eAKVFs44i
MHgTgAOcZfLucgThXKZjmbEYjl6WQ3ST1jvFh95I0D0Xa00xoCKC5KqQpqYQR7p3
WRqAq5xrwNl/2XKPNKzQ4DDEDkhMWK2FG8y8StbBbx4TujH2PCTyuTbdke1fKlTJ
VaAJArgfpl6sa7H+z5d+uRqFP74pdwG/7iCFqPtNeWQPjUSQDfC/2+ZiK5zpyAa/
kTarcEk8BmY+75X8hR1E9efB0F/bCVVQBn5ESOJc40JWollVsuOdKaXEIGLX8QY2
5sZSVZPKIJdOUEgz6nTxDuZjPE5D9kDdVjXEzpiSVVHYorlP7/qF+dhFwZd5/M+M
A5dJP2ZGCzwmsOirfqg0Y/PBCiInIr02DBB2/8Si0alIQphepeV8a/B66JwghO1r
MccwSOfHLMlBkzZzVvrXm2PveOP+tW9rlwXzBkcWxHFi1mG+SM+XI2+IwkHGeAvq
jGBjFzV7NdM5akje6r/5/mqbuDGxKbOlb+PH2UxVzFlZxwF8Az3DdenhC5in5GXI
Hc3oa9reC603jBgoxW5bp3vxzpk8jnAxWWDjN5BUOvkz7NgsexulM0a5iEOZY0Y9
4R2lxASxR/Ngyxqc0LHCC2HAEtDk+uk6VTHjxkIhgo4lDUzksCOw7+7dWxN2l0mr
lwNqhFn9unM/4kNNH1/H7d7VSx3l1pWxlyeCRq1x5jiWinPHwGZ1LdkVjSJuof4x
KFBAFzJRBFMO1RY1YBuXKxKfdoCaK41tWoVNL09dHdzBLy++kVP6n0Mo/2JKLJXz
leRPiu/XKHiqL8lPtLd5EI0vcRb3KtKEHAeeukFfHBqZeL8u5G9emfKXQ01gEqep
QW1lfd9P5kf/tEoUXKkfO3UNXl8GMIQFRPMEi884wjY2kdWPdeDlHj0TpyibyGoQ
lcJ2iLLWP2gxmC86+d0FFboDPOSQK7hZaLQKAubJp/d89SlPKrjLgWGsx+LobFhL
f53cx9rudoinlI9fzrBF2W5TLoTQm9NjrqZAW372XQ3ZQuAp4raSG4Bw7a9RLH9G
2ZbaLloiRrCNnfF8sTtN/z7owUJGeFo034LJ6OoW4dClSu6gwXdpqPOBSqm0BWBp
ze7lDXtzNh6HuigoJQkaxl1M0iKkNcuu7OqdAZzu0a4pootGwwBAVOCu4kqpFpGf
SOXU3p8ye590zOnMUvgWlaZO3CigKEeprCqxhCK+jn2dj1oF1e5cgvErXHXT9/+/
zZokcEDNwCaA5k9PeyniagUMPyElP796NgsXQBqPmfwVMZLoYkvm7+Af0/y5Hv4E
lDL5hhssPZPFsEvFeNI36LpqKJi57vcSX/oONb4YlXr0c1aB9W9ouM4ZEApKhn8L
IK91gv10SeMBR+mpiHWBGYSEdvSu/Yg2nt7Ur69XyRyavsUeGKxiFp5XgcOVW58D
+bZda3nCMHnlSFZqs/MobjaOMwrDIBhfL+HFhO6DagHbXhG3a42Y2EyXuTQO8pFD
UQLkV9p74WELXdtuu2reK3q0F+ya7ZdnNUSO9hURlgEW4RGRY+WjlyXo6wnbWRf1
/20LHqO3wr0q8GDfdmoJRp5y6KLswe/3V5PWIEi/D/6yEowR/K4QY3xqLINUnWJc
zy18y76SjdrY1qQmZJKhgmrA21opxno5nTLfUyetJEcbdWFyZ7zu8fDPFjxLUhci
0DK+H+p6qMtxPgppTjsgvQM+qO7rmnyXe5e4SJ/dooFFP/g5Tu2Zv/DnxlOyFG5u
YHqtwhp1PyGb9WnMLuB43pa6NlE2R8ZbbagSTttVQxW+2WjXYMrjasicpuaMDZDv
1N8WAE9P6rMyxHIlmlCduYa8zQlIeITv/rbXbeeXdAq1pXTiOF98xhrd0xRlCptL
05h1JtzTJDIT9yZ/p/DFx55a7jbZteKqk2cdXfzSx5u5WdtCIgWfeMyG9QM3VVRi
mGF4avSNiNfc/uM1Wyhj/nsA5bsEKob/Q9Smai2m7SSXufGBvWzpr/HD33NLjX5D
QeBNK4mDU0kVI1pxm4U9ZVtpUvAF36JkgKLhuFTaDoV9r4z9ornhl20+crqwEWoe
6gka1r6Q1h7r0d2uxXih+Ux5rhA63c2846oVlvjy345IpyFd4BwkeTW4qhy1Oh9C
gUo85kyt/jHkHjx04XjRmFSC3R/u4bMYZ3ssAaS4xvXyKcORFq/Wr6SUQqsBdG5n
6p3gg+o+fpEJr34C7CuU5ltjw5YsUXz7L8ja3o6Fy7kKujP1yYN8ZRkn54R70Q+R
Wh8DOO4p6uz9QiW+sfqaMLyDSSvi+zKig09JCiguoLyjtlMNeIZfIeAoHLxC96FL
M0sD+cinDZgm25Jnp6yGsW10h2EFk/b+0ps855G6y4AyfAMW6WSIJWPpydmgCMHz
crzFblW6yzcarcVJ8doDXad/Jr+AJkauEHQulq3QRi6f2TIp9OSFGW6tNhaKy1c4
PS3JqijNAHVaN8JYM+FAwLazEdcAT6P7dtjfWcnm4ADvJMou+YvshwIZZDnXoOks
zpg65wiiPEKE6U/Nv28AnOR2Xri0x+QoJlR93+FPwcaz+hghLyHC2o0cp/DSZC4X
psLFJIZOlgDTV1/dOnBUMKlei34eeOFEKas3e9WoJsHbJuaVZJYF6JlAz0muRzvj
h8obhFmpJj/tZqBbJ4Pf2n1TjBv8Rc5l1XVdhKr+F6KBPtITCCNebPZo039SnvBN
butjkQSeGI/zVQu0jpflxPcRw4UD0oTRtYPrgQx/vQoaJ9n0AQbQyH2ybl5eldGx
4i36aXG1Se675BImd8wVgLRo2L2VgwH9+Ya62n4yvbjY1Dtlcz11HmkYeHTiLToS
+oElgEPuJq/gVzxxJung383PEY+XCJDPHLh8qGfyJdf4skjpTBxWMG9k7cD5XIdF
bI4ersIjsjhEprtM/OWSmUrESiq9esJSdlKou5FkKTJvAM65Wn6n1dlIZF4r7bve
CQGce4WlZvCJw+yAAm6cPq6rKA2NHAju04kigL4Hkc3YHFUwfOQl67IYAm5qVFYL
xQflBBBgTxoDdSIudgKzwSp4EQDjGUOXYSCN2l1eTpZAKkTMLTXMCaZINSW80tUo
s400OF5CFdWb2XefmSurNuR39FnWV7efPjcemZnbfoV/zxeiOR7WOvcx+QfrAl/0
023pChQE196DC2xDlWrKjOPtbrRceCAjC15Lmyn+ZKplTrTljYignKVbZGnoAy4P
L37QJqL5/6kGwOgn3cDP1gRd9qidgcxKNOK3BHvDtN4zxLXXRkWpXjiUvNu9q9Es
ZKWwap710VlBGXoCfPX2YqbvkImAdxBxPkS3F+JMIOb5xGkSm4af4v43zQRrzTgO
g8aI9iYHQ9PCPoMI+xQsNmhiAnFW7kzdwHf/IQETMh/l9os+1E/CpFea1jQgf5D/
uiAnxMyjFEdhzY+wpAwgQ1z2zbniIshsde9WBguu5CYcATx/CZom73ERDrk78Yfp
OAAxc4VWzuIPb1dec5Dhn8r3+Gw9jdQsJHhn7S2wCvXqUxNers7ojbuR+aXKy3TF
RAetTq2POyJ4aXnJM5v/LT4XgpDMJIC/YMdg/yjyaf0mYw12FnT+7PXspU0ELbxF
F0NjuW1LV8hwl06GV3KTKEuT3e2YG9zvtMSzO74QksEpLpYBTRGdFep2FRwLUuUv
za37uTMzafP67vA8rcWsOrSinCnx+3qeAjSwbzREvA84VdJkNzzT93FaIl6F9MBO
n0QvAEKic6DvOD7WMgaAyKLTXAN42PKXax25TBvUVQJkyA2mQ7rKEJbqzeUBn5/6
OYSXLtUTBaM84Oz3oDSvZ+N+7cWny7Yd4B2mCDjfRZB4SgJX15gwZ+u3Ow+pJMIA
WCMYi7+yffADXykckEe9khTvHPLFtO0fcfc7C7+LL/gSOydBM05Pid2wtDB3piIj
XIoibiFtUDUGnj+4UHqFXaRaHzTtNxOv1r9hEb7F++vcMxokPtqyzsJ/nTwjF9/p
TiN4XkRxHqBSGgLDvLK+xuD8m4/jFP1d9uxF/snyNKgkOMP2MSZe6ZXPxoSVKqPw
GsVXvRj2MZciHHx6ZX4E5MDKaoetBcVzsXl8J/vao7PU4Z1eVHMCqPpIPougRmag
qO3MSfBhNxsJNCGbVqv2SBOwMPqp5R+BE2k9nqDHpN7CtgnoNnbQMvjwdgtIo1U6
CMuIiKOFynhLd5ssRzGez5jtQgt4F5gvWyln7S9L2zk/4r1PsBdAYbSK/k438r9J
FQeiW0GXvBWeYfEQNS47H1S64x0JZw90DzoU6/lO7Sv3FoO7h9YW318zmRHMNiNp
td21+D4ueTbimU6GPj645G77pK7xZbZv9nOVb88XIaBjIt42I1+9iBk+2ak8m9mH
Wao5/hRuznuMqgS2S7q0fIyiiMqzipGLuaWFY9yf2/ZoQ5HFf/cUcyuum0bCljX3
tn8KjM/02dxw7j9HHEV6CxxyBgrSUxxKvJYUEf5zWSjeR6E37Fy0wjTZKKCsJ84n
WEvYv1WCoGql0wdpz9+lqSV5+DKGzgU6pSxXID8z+KxJUgwTFZYtQagLyy/uE4o2
lS6Zd4Fu3uKu7AC+xt+f0Lxtfp0G6Ha2bQsq7ClDRt/F65OtJY17vCXsMEjI/wDu
vgH8XEOMwQy7UY4N2tp2Rxbc21PIJYi6zArmvFsRq0k0LmCiQxKuIhXYmgoiNDkP
r32N8TmdvHt0KgIsX+9TQmj15cn/Ng2vOpY5xrUHYOOamDw45ZE0mJwtk/aPwXsT
1/Kxd4hlnz7Xw0OY+w0OO7TxUgC8OgRZo8tzDlawdgQpsS3NKxD8gVUxkNesWDpL
ZaDfBhRVQynh/1KBg7ObMNaHd2A/3WYno/Ff8ebb/yyLz/yqPiwNUJpDIVZjdKnt
5gEY1Wm8qgNwkWCc2n3/qZ5giC35rSfLwlp8cTR39A5VHeg18l4k8pZdBZ4IdyFH
rXYqQED+y3uf83nMOdWekiOoIsOmN5eV2L7DqdHSEpvVaxQH8nDx467WO6VCls8t
3vKH+OG+ykPmbiPQQWZwTm6BD5UbCeEUuEfNPV7UuP/ckNL5aS5PWuO3Bh0SjZG+
oUyGWwDQMVvwDsVA245zryNeNxYR300VLDzMB9nquuRqz/JsjIrrkR9fv2x7TLDF
7toVU8A+m/thDh8BKShu3gRyMm8+eH81EIJNcj7kkZHHge4Lnelgg/2g1fKjDxV7
FBBb8fYWDR/JcQYNPMLAxRhsq2r8eaMMwkL+lsyCnHPNyvd8suCPNylMH5lYIr55
kukrV9sS+2B4rc83hGe40Bq/K3FQpkI7+PWn3R9/I+xPjhLe8uc1ihWorEo13srb
kC4QM7xiwG4rB32gyW94k1Yo0hO9QPn3mxocPOdGY5CcIhtMa2p+olK6fqSGJpzV
Yto3hzdoVT6S5nIlZZuqz+mbmD0FHGeimFNk9xvCNhkPbSmm6VzMQxIe1Hr7DcXw
+nqYcJHu2xvVswdEdhYEoHXVjRvcFFNSAxYtIgE24CBH2b+m8hQvsCiMinvazt9p
Rq5pAyzpPfmNkWzPPBxQsbKJqk33ocG62uG3yzBqcTsVu/wQKPR9/6Xgx1Swe2hY
LQJ6Azcos5GmckkGALE5IDo6PotAs1og4r/JJi1M1KffNgFermrRE0aVLcbRBMRJ
U+JK4Ws22HoWo5ZpoAYXyhaNfg8mq0jXTOB99efdJXAPHbHMtLURV2iAy24sUHSe
twPgR8zXsEwTci/dUZKDnH4lgO0cqFi2rhgFT3zlsuima7CRLUNbjn+A2tm9lY2J
9IzBEz1SFmW6bbQZmQFtJGkeZiLJ+ZNRymM00zXFPEdgilQWpfONLbLLgPzLoue7
nXeRLFQJoNR4oU9xNwgTW9i1xwBwUFEnY7ly2xNZWQdnjAx6AVGoZhAGEM/TIEAE
rZuNOkcK7ZRNBa4OtgMizA9YqumCQlCPrlYmY7SQrZGOYFMEgDOEGpBjIJkbB5Gp
M67I6+cgMi1AvnCUYksVkRXavpJgjxZP6X4G5P8nOvImYrgZs9MnUibUkUdPWvK4
aUtfD3oaV8e9v7gs1Bq52KKr58NSPoto3NgrPEFo/oFl3mbs72+F31HvcyNpN8tb
MEZerXnqUdGpeHtsBmhCcPgHPvG+VdiwtqF1huz0bm6Ifaz2CtXhaGk3221UFCyB
PufZMd7k9YG1seXoFxrWGKZS8uYIKnxFXEAbojmSFFNsqJI7v0kkkgpu1hSsc6cd
rt0QlNTNQjXJGdGkePbiKepdpLaY3EeYE8XxnMePOpBb0b3MRhZfKZqkK65+mf5k
em4pMm6U97IIqUN9gMu7Rsyra1wxPe6NW5O/Tsfn6kkgydyEd3Epia/6x4/3ldTM
AE58e62/6v8MvLa1SnOb3ETqZxeFahU3uKxpC/oYGf18uGfjfDKeFS3sSdj7TqLJ
6caceWDk7QMupHlLFLcPqtExwK+zUSBEXua6NB17yITNl5w3kDSjBq4sF5GXrHZK
cWIGz8YG0xfkTJEE+0qR98VMi6P5jgKF2ZafjUvGgN5/9ha5Otlv/K7NtpTDT0VC
GYF26j55QRBKs3a4pMy1MwFn63l+TZ+MIsFTwyucDAhOdkTZJl3AO+skDAgUMGO3
hUBLNIKIiQpFm0NvAmeIMFX4SM1HHUYBp7tt5zsedaldGIuUDevmIs1jlfbcFm7H
16GN/wAaasV3cgVJ4qL09ry4qtpK/aZ780C1wZUZ1XriMV3lLbNgGeYu96uumqXK
V1r6CdKz4YYPHkfJcpbB7gp+zz9+uGoDlDUuwnA9KNlnVNN9Z1JKOE5IM8Mg2vdJ
1hlRWWG9Uzz/yV60XNt0GclSSv9v9FpGRMranZbmwSisCvx1ZdyxOa0ic5ANGzvc
+zwvv4E7vlf9cGcr17e6TxSswigYzdYFFOepkD8psm08fkGwaaQyFUqb12szqO70
i9zBRl1ZVGPgBI0p6ufPDXdct9cbRU7GXTDIro6A4Esx2zuJMopblPbjecT8aGpD
PZ+T+557SbDpzzumeyEERooWRN0AMP0YsdtSRNXfRkeMZQXH7MAhr177vWM6YtY8
niKyWt7hDOuwueUD9vgdzsOrDWN+s4SyxGeRfsSUFRoA2yimnoyS3Ukj5Tszk9Np
fnEF8rKq9NSuWQjJxvUK4HAyKHi1vGFa4HPqiHmVKK5Eww6ZDQvU+cXP5CNTUOYA
KQ6NIUbcrJDQqhmRC4LnaGTEbIi5zSGD9rX8ptYRkJtxjnhQVDnBGIFTJH34Z7ob
ZtNuewye1Fa7/5BNbpN9emhArO8yxeCw+zJy6GYisB58vrBfjHe95Lav8GGIZw7A
6ZIcY6VzGsPbzPi4iGD3fin+gRV+HDJyfxu5UAdFGh58FSzxDXgBtAhCmEPxCbMT
QhcTcV9Px8rTEinK2uNLlfq1ZrX26cQCBXvSOuNXOpHOBt44K74IuFS6dZC5qTNO
72GyNX9Y4jvQEl9d0Hgs4kpEuvyEEzZQShvR3trtCpIf8tP57ip/hosaMT4z4XEI
IhYcWyZB6sEHQvkYOzu/LP8E+ImU0yqt0j/j7JpdWtHAEtGliE4Vh/68lu2qCJkd
44xbCmjIbSDu9qs9bK/nvw2bjinnIOpgLUbr75fM0QhfnH4t5M3Xd33jrk8ywnf0
nmn369hqqjLTH3ofQQsdeZRkJ1s9/W1Vh7i0QrajB8INxXzEFHr5DgIJ1CkTlJGY
yaRB8ag4EygXCQggx+t85ECHASxWNt8xlyFhT/G/G23hEgrueBiMuEmN4o8UpmeC
SJuXiQKQTOmLcmeb0Bef9lOSjSDdDnTeF52ancwIKwd5ifFzw5LB4nfgUcKXiUiD
TCapa2WsHDd3KEEwwA6y5PB2R/IFutr+3vxITCtyZkXvtR2L6V/XeLzsxOzR5asV
TuvXgSfCtwwc3t86qJZcTmK4w9BqngLv+CZG+gnCVQl4vs9kET18UvPnVnTki/KD
sd7Bi+5luJgicuQXLqX85z6CY5Y8iff03KC7ncAENVod3K8DIzPKIUtkEhXXujZO
kyKn3Cw6YmoXKCM8ieBzAJzAIAO6Fawat2qnf9jVWFZNfmohd8WwtJOqFU7kWoX2
WOZEPYGx76W6YmINo8Fs3o5InVloEM4J5GvRkcD1TGr0YI0af+m6neDXcYKD7brQ
Up1PCvSa56Ty9/bGrMueMxxZKU4ikS+LWsyGM52AS9oaNjrFdMNxvZlCEEQq+p3W
eZCmlO0MSVcaUoWtBeNRh1gFd14fxpraTHYOsNcrimA4YLDqcyyG0bIITjo/f3fp
9e1P66boZBG39gKkF7dQHYUczyMS1E0lsZKINpCLMsJvDlRv7enPZVm255tp6Kmz
dAlElphEapsx7PV/6fhtfsG/hacXsJDS6byfLenis43BQyw8+Q5vxU+d3mMdO2LI
YOHc6/dJ2hmuY+wX0IINFW1VaV+Cq56fuTPyYLMWs1oSqf9GcSU0erOqOe9GIV0W
VHNYPjz0XU/KgLHbrhB/VM1fI5AmtKFX3qQ1ypujDiV77wG+VLA2NnI5VIvvN3+U
ulBL5xQD75Yzw60eAcYFxtrrKgHcMxO7F4qBU1e+vl7S2aHG9WGm6eReuliTSMeC
Z3OVBGJmeWX2nc+4aIfltUYsLfXad6T0DiLSskV1MrXDfEKHqpUsdJpY77muOCdo
Ig8Vq063SeDx8zlGDyzog902igJVQcY42+bMCAyifWonvWMllvzXgfo3yZIyNzHE
0xvhkkduV1Np60XUM3iJrxc19cZFtqTI17ReAk+Se2QrzVnDqzgMglpOGwIRyqG0
5QIyOoet+kqKfqNpk7V+2cwxSewfg1wKLE+HbFBnbpuaovVJ54n3hTbOf4UcEKWn
eJRVWIzpWAJMdBTapRnHG1M4FFMdtTnR2GFIxhy09OYES0sjl18NA39QhCGFxVyz
fPWO6UM6i5/TmcbZx2aIMloADZlRE73E7q4QKB2nr/Jegoala2H34yn6xA1DqPX+
394jBYFSiYB/50eEq/90yEvksrukd71YsZi8cTdmo4IMV9pdUuQr7z51lb9nxCqj
KhXdWrQ9rvt5Ht+VZEiUyIgf++Ztw65tNgZaeDBhTW8BGeUdY5sKh5bxV9EBliSN
6k9Gde19wj7holZETOk2fddCbCEyrEKuKc6jGJE3VY2Htwx+Q3IEi1/rNnJr8i63
lp9hc0MsxXf97bBK2+bTwEI5ZkMM0jOSY/h1yw3+5TrpDjb7FZA5ZHUFaAS2G+mX
SKmU8veZiDjouSJGzG5exfUscD/eDZN/KkRhF6whgLAgjzhA3dAe21wfMj38a/JO
4Qf7fZCdZ9T78q8yc6juZ39WfzM48iBApkpLWYmq0u5b+feD0yiO4L1XI+Pf4Je3
3HcH0BhrWC2MpsO9ImAoytVugKvL487bVznGmN7+7OA9UiUHYf5ImpFhAJQUTt1N
oWbgAuVHw9va+9YgBL5Ht7e2GKT2XQXxGKLc8cjc71wgPlXKhIumQDFTEg/hkrC/
PpVXfB1RF3Jlv4wJhV143eNaeLr+8AHVJ/kZN/vJxFN0qtUibQYI8W4XkWfTaJhg
AYssHoY2/x0b54m951Qcu4T9cQpz0gihZ0RrRF/DCo2rAPxgvHUJ/eNAGoI2f3jX
wFOr5gBmPoDxyvvHhN4pgl6u7BuRdBI+sD/4+JFalTNTjwhOxhv4dOxiIdSHPWBA
9fnpYWlTHbZuEdI3WXRcBkTniG6qgWab5y23VS5jPUZ/8Qzx0uolb+Ut/SxdwWtE
wT1HKr9R1SD9cov1dL35ItXzy6d0WMS3Jqyvl9YNp3J0RISxML+tco5CPjc98dli
d8W5kvDAcnNcNPPQBsGjZ17mAj5NY+PxsaQowChg/A3Fx4eHB4bsifo39BHRMOvU
d2aWQf//zI4wsisLaLMoohzDz7z/PozGpWER9qkFrNm2Cd2JEUwwYwWa7f8D7vdX
a0pAQ5UIWPwjRwPtnIrF0wbqSpLovXHxuPim8P2SeasQotTaTHsiYH9SITc2316c
qSsFldQaEvlcChg1byPdYUxOA/YExDoA5kzUZSBxz+Cx/Oq2QF6OUlAruB8dIzhH
fo6O+R95oiqBkTh5bkDBQATBVc6Guj1llNH+F5p+RToyuH2hW+p+0PKwR6zQ5yau
U99xLzfuDhC1Nq9ArGaOB+t0rtFGMGwis4qGInebeGCvPpbpjcTqEqgdQVqwJ8Rp
jAB4r75frDlE0tb/ulGw0+WSIUp64hzvA0fEJCe21+4lexWOeyHjNblXAQhJkhE+
KktDbVCQdXBNMIAGyrVlgSOCAMpO6CvTmGRiefIVwPFc4LsfPq0eT8FG0N5hyHWX
FN/A+3r1S4OUuepTVZ8qlJqnTP0jeaa6rY0yXgVZs8N2NaXYg6Nxmoe73m6U0tBU
NHQ+YsxQ+OxqxJUO4ag2ooIKY7nmptdloOAB8ZvA5toW/FKgTh/Us8VqU/xDIKtG
kN4C8Rh4kIw7H5E1qUg9RDwF9bWRKxqZcZwntqVGgZw8lnZV+PWDYlBjAMQU2h+v
OQBCab4U+QREr4L8naP1F81hq6tkS/UDoGt/RyWMlZifp0XpnecITk/HVi0oZ3WI
RfGVcQv1Pvhq7c3MCmQlRvLtfbyhKdU8H/3plp+jNL4rA7lBJfg3uA4PFNH91iTu
5UNvcRaWuPpxu1E6+ph/fC8GTiUbT64joJfL540EfIolIsVibiJoVuD3GYCyDQf8
/tYnyxFTdYXavJui+Ko7hfgqZYEDwMyajf6hVJ1+eWKsPwASlEBBmgtv7rGL3cIP
HmY8sdpo/ihxjhOOD/4MZ2J4qvE5TppjybJhpSbOAPlNODo+t5BoLviz5sFIexgw
m3+InXA+N3xgKcA8dErzk/C0Iqo8nC+JL92JxH3KCYbCfauuK1ma0t5e7/GBGwpN
BNacV6uI90ebNj+DXLkUabkr53H8RORgmaiHXEzfabinhnM0rcyUvvDYZZp+uxhP
V69BUeVZB0nZ3NpBtm705j3cVTrUxuSem5YR2lYXXsu2sjEfgBzGPy7hX51ofCyQ
XJdmod7BwLmTAQ7aPdrp3GU1fw8v3SDaTm73rvLN+Jt53gSMjAaDuXzfajdJ+ahf
GMpl3XtLDjfXhp/CrHiSI9HVIKzFdcD78Qp3XuPp64aB9baOUzYPfKXjd8sDhf7O
qiW/PE9zCqGLHUay/MHjlmOobu+Tf/qs5RJ75COQaAvsO+WFomtIzgEIHhtsBs0w
Gg7nFN93/iL7u525NPPlYxYCqIlpyuPxNXRe5ptPne5oVgvXDWm29c986As4DSpz
SVXEDf5gdSBtnxDFCFeGR3ullCVNmLoDb7sTmA8v8oRwtseiTSgC77uBXeva+Mxt
TDlLyRzNU+fqF67nfI+3sjghfE/WGQm/PmIXM3NW9n28PeCWrG0hz3l5aaYJcsEq
6V1GB0YlHgSVbqhaiQDNr6d+AbK9ADwF7QBTsw02Rxx3rTnT93xVq/Jh5qJjm4Aj
hAR813e5CZbS+tQEcRIqeAUi8eOK/KrfZ/Wq+jEymf83LtP7UMaIAEKlZsLYmgzG
ht7CgRS29LSKiwiBeetyDbNEY55JVYbzgqBpgD4n/6tEMUckb2DlaC+UyvZbBFAg
HT0ApiI4l5FB+srXdYCDI4b7sXhe4FqT9t4cdymo406VQew5idZvYrQUUNvrwI/v
tKjymjVJBPP27zR54JSCC4vDhRBrA/6bmuI74cSNC/o9+DBhWTXHVRKcbxIw5Vfc
NzdwArnh6bxkaTIEZWz25OmGpC2yP8sse3O3/ojCqe7InZoMaPmDK6jskLFrbqi6
kZFzd/EEifeq7kLvSHiZK7lHQk/X3Ln0FZewRmnDTACPk6CzVtLu7MC9c5piJFWz
AcMSSf+Q3R9m5f4/17qexT7gllvujTp7C4RK1VuBn9+WIExvKkEVs4o20UlWq41A
JY69LlHb7HR84tyBXZO0OpJ52GQWKN2dZnIs1pbCV8/rT8IEUWcxQzcbMJxq4/gl
XTwJg9VRMMBKPvlrCGpn7X/IS0eaED3NtB7r4AE162Ed8voSW7Ilx8+1EfKt83OZ
Zm599M72tNtEqQWJKmya9OKRlomIYEDfetv0lqNS8OcuBaV7bqYR3RcRn6nLcanJ
h0MPJwa0/mfx4B9NHmWKyplDUaUbs7f/5VxWiJfgBvQazajAgiwGwpglChAFT1C3
2E+Ag/ff1mfUFXXE73ye7QMU1gwU+DmpVSFxdk5Vhefxm84GZ/WVwwU33ww2Odr1
BFl83M9E6JU9I49PjT0hO5JQpNSIQPMkM/NrCIiLUrlvO65orDvhc5Y0SCXFyIO3
jzWaUYjx1ssBDWhQvGc8x8RVG7ECDXuDlGEWlfebSrmuUnFrUWl1bwRagGC/E3N4
T11S1xb9Ydj0fNEn88y4kK9F4GIgPcAI1hyFwThw+GVXZIK2Dya/rMFT8Mm3S1wC
VP48uDbtoQvTzec8wStHuMFScUPnVJYScq9tPJjWV+zvZIRkxeVfmnPp6B2IUP2+
6m3a7otbESO9O6iUxh3jbtuEODrdmawHKKottgdd8tjKNxMdO6vc5VSirN77TbXe
xbq6aPDw5ra1DFgp8zf0pT2Xv8PqV7AZfTr9KDhvjWRlGbB12mUCv2CPJWDt4Nx0
wztSviAsrO6dzKYNpiEtNkPj+zlGMX5V86/AWAYEvTRMq1w+zB67mMY85/mnELRw
Hb1V+48PlxXuBypID5+McgFCqnUedf7uuEscWhY5Lu1Zha+636GHxYcq+1iNZ7Us
w9IiTPTS/OFrT5weaBQKiq9ZD6A7Q+Y1aOlHbnNJmSLTFtWMugxHhk1/h4VQvn5i
eujUVFJeLy2hRZsQ1U2qEUm8i/MWfbC2E5GKzl2kzAvChiypFIWQE3x8xewlYvVK
vKcg+wsKkEokQBYHDfgaIvMfNdsyJ750RRw0+OWdZdY2glItD1FO2C5snGVAT++E
rVlxRjMSJY/4BkCkRUPTG9ALBLxmSvtUk+K/ffWtLulIlt2BKCaf5Q8Si2CiCeXn
Jm2bG2wh1G0ki2Vwz7W8Sl95SNG3r89ARF916U7nlROo5F8mdVb6GGxni9TpMoKD
08sSk5qFVxc+VRTzBrDj9O2AwaL8uKM9d5palPtviG2Ypb5vDVfk46G05H7X4n5N
8HC0ew7J/IAOEp9/GjwmuwkD2/EQ4+XfJ5cOWCM0ZP+upX4tqHUHx2+0bcyCwlDa
tn862U88DRbx8MtB+G2/JlhgBg4csFTlhKHflTKcSfNO3EG4KGhSmLz7jqF3dUJA
IMFsmqed23qeoBuTl1Lnq/3JInRTcLGqzmj1Z1thsz9WAluOlwnPmiq9a1cquXrP
SgW7Ocz46bnwU0TRTA0I67cw4g6vo6SqBRKRU1njKQrvS9+efEEqh5SnnuRwfnmV
VEL53gTdVOxBMg2VXlyCLsOmxy9QV1fr5e5CSV3WEPgqDFDz1UaN05FJWI0+zzeu
csAuCqYC2uRp5iu/l8x47fyx0XNKnkNj+slj7X+mDr0EgncWEoyYQE+NLOFxDzzo
q0vZwhzjJsXmyAxylJUEHnNRSnSFW35askJBM5r6lk8ekM849CE9dw9Dp4MBD7Vt
OalxHjL3OTmArtXiz6m08PmVOrQ2ZfP8WIThHtrMc+4Dh9aKueMRIRN0dLddvvz/
zOu6SYb73aZQJ0bxA7D1IMUGqXdtXIpksbl2grGyXGyqdKUGB7L1PimwyWxxLRDm
sivnN4R3jJSTJEKufqeqEFTNUfNMUDEmAMtr6ZriYSY9TG92seW4Jj7IYXqCKCvI
IBK1gTiPVp5QY2sO1+t/RKXLSk4NUXpMcbF0m1VYITzLOXdaB+PWn+ZBcjrRzHVB
wEQk2eJs+Rh70UzvMHedJ0nzJI5FQguKt2FmfjufMHw3e9bfrctGZ7z5weJwg2q5
C0uP6JY8ULU0jzLu3+E5WpOfnQHm1XLc4/JXyFUUfGnEWWJ/gFMbBB9rXKtGYUQj
leTgZHz0NcemdzvkxDlDwaSmwQtIHEVbxxj76+BMe8Zv98hPLhKbFAAypGV0CNCo
oZiGcCtvqSleceME9WnQ4WPAlDacTNYGKwop5cdoe0IlzNBRiV8zjYrlt6Jg3HNI
+pUhhpfmudysNqym//5sKWQQeUabYqeCyqn4+rqhid7/WdZ10RKgbrqWQpDSs7g9
7+iOy+0A8H3DB3zUs3sYmLR/5pMXRdEQCyhBw3iMgT2DACxzFIAp3d0Qw5j+QreI
WHnGdv7zSmJzzsmhGdDgSPGS3biJwchWELmdMPUFetnwAOWvdmnb2gQUb6k3LDoF
7OA/cH50YGyPZ2a9b0UAcg3RJkmsNpSCJIbn6u2m/vF1Zp3qfOFmPgEEqgv2HXwM
HS8xf1ZvCVvS11zXvTiVditDPyOxWYrYljXIezat7KKrad/CtbfIE6fEPyCLlzqA
r5pX9N70UgVPmYIT337xK5IDEArHJ20hhDbZ3v/NWG7I+sZiAQz5T3ADpeJNAShl
J3cQRjPxXeuJtDQcib2PZUKEWN0Ra38du5zWIwK6Wv+KPVhcVR+RzLNyhN2LCF3g
rnGi7ecsao0e6/Y2YLHO+8S11Hr+Y3x+y3CIZeeGjB3YKyuK7FENahx5e9HHERze
OPzIBpvyEGVBoN5dCRkLGUoMWSxdx2WRTrXcbyTaD+3f9W2sdWVRIlf9lRSROaMM
kXTTZoQmVyKMtxkTjyM8Xh6JacNd0uNTEwGNz6F8OSIObqDHpW9+TTSD79VZDl2/
kcumTxVzHN+9hV6fBu8/LrpXzwfhfRuujt9+MiU1PIwdWDkcMUPHmcje4NxqZpTe
YdS0ZlSWdcORsLzhRDV4vPEo3oFDXQjL1m7Gi/2bn6K2Jw1vC0bPQz9Cj+1ahFPS
ofaDzjUi6ldWBWaX8HZFpelreHw42NLw3rFwEBfQfVM4ECNy/ziehR3w7nkLxaEm
ITlliUnagGDBOnPDQkoT+imkZwP92eSbX7VfL4T83wC72B54EVB5qGdbpaM/CnH9
2QTdzWUcVgU4K5ZI2jj5PwiyRWIaP4zbZ8rZpvIcttJixDKLVTx/kd/q8wCEKCG6
5Xcg9gZaPVHvKkFH85I15B4QWU8CDsmQ5HxZSXrhZm7IevFadarnxQgq1ZhPYA+s
mqRoYp0Fn0IUayxjqvj15B+FOyU6I7wjNtKY81s3khh4t5BX1aI3zQHTbShdkWiy
OXzpzSmkxjkxTzf1NAzgMw54/gmGZHxLlJZVYlyYHoKrWN9BJwe4x/nViEdLmNnh
+Mpcef4l/QteKFknczOMUp8NcEai5JmjjVH2aTkL8jDjcu2rHILgRhjImCbocXTj
hKRtrFvlIL5nKrhEtHJ24gREipgxWoJYMSFgfMAWtEYgU9+GWJGUKSFvMVMZGGpb
ks5nVn8SXlIGKCHYNMEXMoYnNu6xdfTLcy9SlfVlJ7SpjiNKi51nUJ4Uq7IMBXaK
ikfG4rHoxzr/EP/WcD/IEA+nkbji6GKX0BcugbNT60eN5W0IMbjzIJz6Ys+H1a7y
IHQzpzXFg0Oam/X7l+qYuJmeeNQejSmunKJ3C79yvlSRj/8Ua0Qu1t2D9EYYJTWo
uxNTgQScbXE89HnrCuunIy0lsaIKzftr86159DjgM0YaR/mJzmKD+gXeheeuPxFL
yhrcPGaB4ntsv2ayEVO3vwXkDs31axoevMbtKWAI9EQoozE4bcL0e5qe6V54wBfn
t+r3/+SSBSKLrpYtQNTlVpemGZj5ungpIhfkPDPwo2nPnJyyfECNR82+RHhjeobx
nunUlCQFuiSVaoq56TbuTvDMN7ThR4lhxIcswYJOatN9K9qC0Hs0xr7oA5STrl0G
aP2v2STw/XYvgz+PEwd7EjgnS3LOmAvCTk5dlQpvZLTrRWA444DsMh5JLzu7Z0vU
7CwQmirQduar91hLTd/+SsG2wVoN4LPs3M/+Jk/1idgHe3xoLqrBZlbB7iaHQ4JA
y/2LUO0pSuqD+ABdm8nLuelkLzrdWZwJ4Shj006Tk3zI/Y/L2BvU4kau1KkygnDb
Neo3f7pf+ts3utJDoNVqnQ6KKeqO4/xcJkV4IxMN+tcHSZJEQ7jOL5j+36Z5kfZU
saKpurYaSldSVf17KhdSjY1OWYqsd12lmzAAcdt008DwBZBBIJlOWLGU6ExSZE5Z
Wp6bHAK+J41IiesFO5wfT5ido8xqd0CL5QmqC48EvGjYVJ20+bMCfNaWgCwnQ5fJ
TUCkeitrB7Bf5SJv386j731nVvmH1qlz3gh4IfPIPpo9oc078gmr70K+QKZP7y5b
Az7r8YJzpCeBYlwvQpA55JD/Y8UuNsl38O7T6r6oRSF8vjbrCQoAk9hGPX5QVVdY
frEn6zL2Dz1gNRVH8pdzw8l3M8sU8mu3hRTBf7s2PtcvMDrXq00D6p8zPG8oDWhp
kqFzxM2snBFzHK13oIQAsgQd0YtHtXkk262TgtAikGK3DsXFmCzMy5GHGPqAMsM7
7AAwZp0taU5/obRSp3svFyyRk4RaUDg/jY6DeKECYMusby05284YycusK33qrDHH
JwSlg1T7VBLXtD3PvHkPJgabOezMGGom9HasWVt/uDkoiHW2F2a2mK0RRmA5f5sY
YyoT/1/llUXmq01PuQfBRkyQndA1SY4zFSVB2IEr1ZEVg+sbN/Kcby3lVADI6zwI
o5VgZQjdFWDTEEDtgpTqA+ayGsy923D2OEIG5hJLhYjdFr44eWoa49SwyLDNUxDZ
Uimo212fKz9ATIceqf9JhNkzH42HCPdwVAqdDGuvznFOQrJhsYJRauwZIv04NA0I
8GG6GAj/uuQkfmkokqRlsDJsKS0dnKXaET9Q9fPL9+/kmNvWZrvpHXO8wc6F2APs
MnM6cBXDApke9diWJ4IVSEUFgL31u+lvioIqJmjGZCdvGWH74R+e4zKNyKu+Z5bx
CrCpvxIVQ1kHt4VnWLsuYCYd93eILO7OQlRFmKRwY+7H0BH+S36FXjb3mDKU9/tZ
v/TwCfa59GSf9iglwa95pnM1l7doFQkszcFRKgcBggNJrfcxkMwBX4j1moAQcUyB
7//NiZtvOU9YmrAgvj+A0Sw7UebvrsEj50O12Xx6i1GS25iGOtArUC9yIUBes85k
C8pkXhdmHEkecnuLz0V+RkuFkGXwTmic0DaIxhuRz9AjS6US+1U9aIe3yGym9g71
wVx2vh+eDWvrQzZYdvnDsDD003/JrI8wC8btdxbBIxKHVunXU+5NXOzk3UhOCZCb
74z0wxGUEp9osR9tFC4Lk28QJNgpPsw4+p30O9Mdbl85xp5YqbwXSCkdqLsPzHkc
q27IzlCumuGparaSb4nXEXfWZxC0QRXpNW6AU7HWmPG5muC+7DTsuhNa8/gK3v5n
5elyuVBwtXMTXsrCKzJRgVm0wwUxQB73ijX/cGuoxBhihrlLiin099lwRy3DF17d
UOMppwkJU9wI+I45eimr9jd6JrID+v8P+FZ13iWWCtCfyLiO5WITHUf7cVWfMAL9
pzl+TXOpAdtOYndischlFXzTeGRUzEAYuSqBkqwMfwAATwpl9fUvYq6QtOKfDsMa
9vzS+0mURvlmLdz3FPtMwhIS+rIr/784Z8nbYMVXQVF5FknM+iE8v3Sn8cwWk0RL
x4cIqBYL557hh2lZ1j71KFz8jvrmX9HY8SoMOMMozjcAQKbVzg2XkeK9k8FEX9LR
jcPJ+b27jsbVQPfqOIwt1dCNWJQ3e3TsG1nx1MSl5Aqct7HOlCsaz5whvFA2gLu4
sTYz6xIvg5g20vQtii0WuJtMiZ4B1kRcfhJ9L9QKOy2oSUghA2dkpBcqiSO2RgXK
NWiQPfFK6/ET/+06w4FFPH9hQ5EwB6tB3GJzaXo/Vt5RdH4ewM44fxqOw0S1xH9I
+FfTn/VNUcvuDRVXGGEfRyu9qGWRsRxJ5ZOZsiNjoC5135XKnf9l0iKh8iKjAjtf
f+LXxjxJ085tKdi4bKqi6wBIwBb6DkDvVcENTIm7OOa1ktW/8cEI9MbiRMGucs+g
7tiXiMFLR9ZntkoOzyKD3H26LW1w21vtLnUTM2+JEpVIZDCyJVvO6qw2tW1WGwX1
GisKA4rVoX6wPWYTVU19Fy1UmrXSgrK1MhhPyNqrzYJaNdq96wNnHOpqG2B+3uFj
vClde0pthEmr8bHZ03foOvLFrzCN++MdIzlg9AL7PojJcfnc0BXsYJ/wqzM0lOSE
1i2jZofudiO8Poxc2e7WobeVd/kABm7AKxw1+u2mPpV2DP7aYHJ2s/15BvXcGSI6
e/OYEKQzHZY8q8feEzVKCAOrGp1Jhr01ajeQzJVCwnxxhqw6/RodiKCUYcvvwMUO
59U+osC4pLnxKBxd6wgJamPTk1lOywzYM5UFt3tEHxMmtcLX8U6ZCvZqt0Hnse1Q
K7zy1IKs+f1XwwM1gGVPQOmF3AuatNonpiCB+lh/sfOCX2nHkA+aK7zUdBf85xTd
1TUGdGphNVVESO4bP0m8sx4ULAtT2j0nwLrSQXWEQQ/u6fPnOLKUPOz3rCYjRf/v
PDK0pnSOYD+4GZ0pFSaf5bp2DTPFLusD9uY/ppYP8MDRRVnLzEYb/RKRSzAvYQMl
7KDv0j67y/fCcSALPBLbdZOAU6yI6YPZd2QZujH2Xhz1F9LPnTdN90v/6QL2EfNC
W+IH+XvG5TdwENsEqUejeGfQ+tgTASGVf2cxgZae3Kuws0DPG4ovSzweapFECYdE
3xZkX5pd0yxH9DioZ/noiyGmR2WDRyViZAy8JcVnIeUIKTZv9ClXSlS1f4M0ES7J
dcUHap0O+XBL/mK0DAJAvRph04ZVKBcHX4S+xuYZSqzdDlYtT7SDX6G6LecwoBzD
qTODgKyc7/2H/g1Llg4NCa+Wwl2JTrRfLuzgM+f19DiKsTDW4EQxfFVkeRQ2qsVu
NrJWoJmiMXe9LtZp5d86bOB0CFeshvGkVkdfV32/xuxUO5YugPzZaavZblD8ZFM1
JQ9PsZXj72sbQdcV/fazg/n2owdN2i6wD51H/2D54s1dld6yYafgDt+TlHhYzlIV
h8e4wOWOdEF1lOmOCul2LluXY8wFvtRU3jKzdusD+rl0k9HOkbz9XgTGF8oFsKg1
hbr3AQnf3Vwka/DpG+nYvCXSpa0NjudZ4lMxElDjl+xdTX29+AVqlw5+Gy+H8Oti
pPqy2koTJGw4Luo4e8c+KKWYwEmRkDNLSYcAb0A0WMCB9Ryes6IeQmjes/3hB3JD
hgIrI0WX/kuxd+aO3+9GEa+IlD3rT5w0dEaeKGmVcKm4YkaQlPJw6MtjswXYt36J
GZ0LdyplHqM9QqpJA0OIebTxf2jy0ujE8CG+16KG8ZcxFTH6vdog9QBDVZBGOxHQ
/u7qcBKVspYCZe5NsFqyx0W+lIsS7rdUPJQMqNpR5e+Wp+56UFM1leaLXUKqSAOB
hx+3eqLm4oIyBtz4geyok4ioL+Ni2wqJGt4C0zskQ69G0oQimr5UO3wQOnHWnsfj
3pEW3VDVUZYWzjHI8+qDjSXUIq7uBiZfUGTh6ndfsnOWRcHd3Ts9t0Wl/Z7OYy44
rtOlT3JgqLp6knF+qKXP0zBMu0kruguQsNiR6EbFWxYknzvMqyAKuHomAtMKaK+R
wcFySL4P9Fsb27GD7x4D5pUAFIB6KCVshe7/1edgrreWAz3xlB737Ac2zjL+3xbX
Oewa2YICVoJ0SejY82tIJJCR96cNttBgR2FXHrfG/0WkN4Zzo836WimsYm+BbpK7
TcBeA4/Ba9910MYYf7eISyA42MZa32fbEN44OVd/9VlJzsQlaAYFLKu8k+9mifQQ
9OCMLfCSfOOB+46/JvpCVxcLrZ1lYrmIcXTnUKp+g1CtmCjLLimcX5Wajor5rt52
W52FRMuvBKIj5FaBhYqPi8K77/CS8EYCRTfCUQWjs0TNDzef02BmBxIF+nT7z8Ib
uaSerWrVD+Hck+qYkI2zAQgw1fsLVtf7nIjI/O784qmy2AQeqP31yc4+pFsl+ByG
tEymMQAAID1V7n/BpxCIyTnETTULZEzrWPLINzKNfnpsejm/ZvXntvAjZbq0sLiZ
pyzoEYdwGZNRy1Ge3HXoAOmtg+74hBuHQ5jRoawnECFssvwIduM4DfVjF1GJGizp
tvSgHn0P09JtzzhT0pCvpXeauaTtmHciFJTB8C26fAYKo6qZsZ72SxDW9InPGxD5
Xfqky7ycSvaTdffcAXrr8W9+0dfZIRDqYFmY19Kn3xKRLNkJvp4RNg/Sl9ELNc+Z
dLIAoh+TkhfoGtehWwMPlVxG7Ji4oTS5XP+D4nCk3xOUaYiS8bvmWgNcFnqyV4z1
X0u2KlUzAZTms30v0di+31kAqkuRlNIHcP40/V2tNHiNeaN3xbOWh120Rscgva2U
aUKEX0GSC0qrcEkz5TQN48MfVzyPkPY546NSO+Dhc8zNitGUjHKo/whD/X8a9yfj
UfjIptjKb4ZV62dT8u+8MhuIfQVP4J0R+CHhRzbGI6pAwf1UV/3666u39f7ZPtED
5Wh/DX2xZZU94h4g51SD3C7qQGifRQ9IzgjgQfHGKl+FU/OJQkPg3NNZFpkrm14e
SyQLeBmT/XBmHy8HtbxCyeuG+SbEnpDXodZPxPlEZI6QowWWcUhwVGQ7ZUW+yAQ/
g7FmGK3cX8dM9em/qIwWfY5ODFs5E0sKb/qpAVCRZxohGMT7lBv9VVxO4EVJznt+
aRnTB8Y/wzExNgDrpr+yxzhnw2/ZzQF32xLUe20f753ZF5iQKOWO3OPjf6PPThk8
omObFeULRyT99r8iF2GasXRiUyYo4CJjvlc1TwdP946F4UA5mcNv6CvwJmApqpt3
cBkOVQZvbUzCQGQTY+xXdLLIBWAr1t5AOvVVDl/sUI6E5iLpjogGD7kJLZ/c4C7j
pKGyuuMw1qrHTYdVntuhKoizaxwIi35C7Gko7cQv9+Gn6jurX+7cFEyA8uNZNxcK
HaBD2bQTO6gSzSv6ygxpAwHaXcb6cjwG54EPklhKo9Gexml9BfmMrK8a0vZlPFLg
jieyp9PMD//8Jwh8T87pTezOX4xl0IMCjDlNA7YEBYEmRIfygQXoXrDlKvQpqae2
Z72+aDpgemoh+Iu72CVwCr/3gJZ528dlwlLtSu6NFFJj/GptBmqBdNdT/ln6cFdt
8vR+auQDLk5kEicCbRexhMe4ZtnGRwny2UKs1Dltlc2LSMHK3lET1UEgDaAWzFr1
3AEUhpMN5XB4ej2PgnjpxJG4FVDZ2rI2ffnd6GF+Or+5pt3oGYblJDU93SsAkChR
0qr8FFZV1+CYy2JrBGJMfAfOfm47j5MqAXTMdsAvSKbxRcjfFTA7DWNzz2pWaYjt
ZrJ3ANEx3Qv+NEsikqDJidWQd2T+eH6J0dP3fSDNI/cxzccie5+C+l7jEY5KXTP6
LQEnlZGXTkyIV3deA9Cm/RDkE/9vfdjahe1lfMInXfB0I5SW5HW/4DMKmA6bOg2v
pitil+Mzt+C5kqhQOl23uSTDLyPRJ8esOhkBzEFFBjWlq5pF3KBOYdmEwZpOot4D
gW0bg6W2PGInKpyfi087fXa1zGc0DAcjKFQJAcvJBMkymfSqMipnCb9GwAE98Yb8
3FuE1wxaCDRPrDLlUfemDtTPp/MjfvZTfA1TRyCvj6ZOMw3abzVzzm6w+ZGF3uTR
RfhjJU4IkPHq1lj6S2qGPSzH8Dkzg4udrsPZsMmz7ztucCnh1Vmrx13+GWOGB70c
w83l6pq/cPhqvcKycwwT32z+DHVr7BxuCiVmJRYJ8RBOdGOO2GwBimDMc8WuuGqg
Q8gRb/Pno23IbaXrAea0hJPQTs+eodOC/NEtGGNcO+D5ZEPXI+9nWrsQfL8Fq1UW
kF/B0xNtMJ0WI7Wn6cOOuMPMelN9pQZWgZMofH5pSAk7MnX8AXq3BTN7jDxVDfws
TVHm3IVhHvNbNDmdvet4QYpuF2PbtLOvebsLGkq3w+5reqL8qMU007DxIo5GmOuS
3ArAbJ3BaRCiQMyMAkdytHteVRRFzauOzI40fgDFNm0ysvcTJDArTPfEKOvPjf0p
CcENG5TXO/Lu/5K4/+nAjDdAesu4entxMkEn74P40UhHBRlrrntNNey3gRCRU5xr
eqM/FB/rlhNBNTs8CbW3uqLBr8CM4QtGavzu8F9wsi0uv9WHX80wuC8zxUoqjd8m
1gUAtZypG6Dc/oQCcXveY/OSiRWeTYrCOthYO9Snu4PQRxJb42M6nVNGZ+FpCLpc
HI168+Cd98YheJxp/ehxZ/hCe0XazYCljV3/3SUkTr0cgVSeV38q9/Sf6SHNUMlv
kPDczDxQZ3RuPAmPnQpZvTMkUb52kzPjc8YPocPwARi4N7yHdgjK4uZSM0RL6Vxi
4eV3bIFk1OCb5sP2+/kUpBpHkMogB2wsOyoq4IKwhkSA97WrOcdN0wmo/casdAYZ
oe+kHiUC61vy5rm35ThMEzwhrjQf1xnRHtX4+3tDzlLKWOgTPG5ywlZHIiz0nbHt
Rb2lGrEcw48hk9cnQ8rehfx04LBsTK2kzGmfIkRtLO2e4ZMToc0qKSFskGoU0GsF
xWsHfJV+CWGCZ9m2WIDLQmYKoFq3rzEd6USgE5qhuQ2Hf0zaXdN3fJ5OIccu+XYR
ms7qrLcQthezHP4mfWqAHbbx6hcLJiCHeL54AdT2t+ficsLh3EHTCMnP5XJQ/4Iu
8ox8Ob7c1wxKVo5kWRmqNhw/RFgJ5emZaZgijeYT2hjQ0zS4MZxVbC2Su5oSIPi8
2vQGxbrzE4uYXwDmyeicKTw8nr5xprxDdy+4na0b9FsiNV0NvfwHNYymrlbgYNyj
0UxUEgM5K2xS11lrefsSxluFTZ80IsXo2FKTFjV4uq4Q7UYylwyxwsCKT2la9WAM
gOCdOVn3H+iNJwoI/UXoSkQSZ81U1xQ8IQlVNU5g5YuOE+kaj2cbjTEbwzw5Ksc6
iC1kQpbowbQ7KmDh/MUftT3R+BpnrFaKTSBUc/9F4h5JjC9T7RFe7Lq8sWRaB1ZX
H+YFdJtqFnka01vCabCftOkQ9DdpUIRG4xJyj/TJaUEIYwwIlIXsSTIdutYQRYdV
1bErbOQaNejRYQJVMstpTaT+KSldYUicAc7pnm43iokcyj26rT8kY1jmBtG4q5JH
FivXcI85M7XbZUz/wGE9xhUrGiFSFcXpH/g/DkuZjWbkXm9jUY6JmxYTrOzB6W22
Mg2f3lMNvcrRli+U8xJnBfvAa3FV8cpT+94xM0BKGb/jkcRuFOFFy8SPE4w7GTeR
QzU8KXcpcX4pkzL2n7kFPYr9jtxlz2dusPkHeImzPnGh1gwedguxO0gCP8HUO7k7
tbOT/48kfl5FSSerUpRe3DLqyLQOoXJarEAkB2/Pmqx8SxXUs1n46b4qekxuTIC1
LnGLu+14MkkBnCMhZZIxLvuM/EefuCPz/GjlqnMK+doxPsXMee1FloTeT5ZcYXE+
tNgCb/SwF+qFolEHeAR6HvsjMiIMDOIivPZonMSnCkUgjqpQG/AiNJeNKgB0pB1+
WkQnnX0QmOlOmHU8A6VTHuQxKMGPX1CF1jEIoQkQjqMVhJPqOFVQbLMA8PDH3Smo
TABEeYj8GhP/bfOCQqIGXV233Fj2GwzcrCMEDE3ipfDgUE6JC63Ei9vNFiIWj15G
33KItH6x4VPS7iXAu1WiPkhEs+iRZgTSdii9FXIAwSEiexIbI2rJwpmxFZrIKf4e
ZviGsMi2dDWybd9oHbhMmiAtsAs7CsUgKTePvqGE7EIhj+vdDQCDiNjHsJw4Ww+g
A+CEw+1ASZT6mWeEPBFXkrRaz0dGROvxlRfVAMP4fJvyUWs+s+JrfKRFKxOx3soB
CjtZGeg8f8DfrxRzL0qr1FubOpibcpAgftKZKcHqSGwCaIpmQ1OrjEKKe5tFNu68
ihuCpGtO8hNAeswLX8hlFMnoXSKN17Dj2NO7N6P0di+WUG3PBCUC1VeHglg15RBG
Ja6kEYPUnFWgVadGpvuDHKuZ7TVSu/iQlJIVEFjg71B7jvcx38J5HbR1gp4ar3JW
TP4kIExR3naA3VUxa7X7YtQ2gvGlDkXMNgQjMv3RT/Bi2VxVcdMkaY1BSjjMUmk3
2Cvtt+o0+OahqfwBo5aYyK12a87Ruvf+N9916Eaz3HZnB3hv4ZixrN9kaIZT3qqd
n5vYSti8E/zxIA12V4dctTqBnPfqu5yJDYRBDO2V97UkVKFZH382zVodk7jO3bty
dYn2XMDPEVaBtvHtD26oBlYQf58I8q9PKSIngcN1AjpaML2WbgHf8JzApxiOygC7
SSSWHDy2mRCbha3slxMdehudatNCa9eDdlQM+6djhIcgosOHhhTffC7cDtQKxiKb
fGJ6yPS+RjOKAkII7pnFV/E8D5wdqrG+CLj6rTPZHB6dE94Y2VkGQBPwNMp8QQ5U
Khv48FyVJJZG3Zcx8TueqAeaa2F4PmeSvtRQQKflT1DcrOyTfdSmb+MHGGtCv4fY
ESKhigpWMGgs+bU/HErfPdbuploLTwxQ2a0mFgdyNgyRtWPijQeMNOSjdCzU8Eu2
twSISlixqluehuVLZXtC5C42cg85tF1fwUBap0UNwxcRb9T1YfEzA+ROf7PDN1Tv
+xS03Qly+nDYdHe/B5YsTRGpa+q0n1y0OZnB1GMGa0Ngi8soZqDntsln/stuDPz1
/pTQw+H8vMGwXKF2HlOVHoHpmbZveBR+6wehqrmeJ5Zdq8F2XYKzgb/He9BpHaG+
BFn6r1xPQOWFVb0T2WcWqiPTwEFhNmpVPC0Jz07usf/vTUIMjcxmmhd0bsH0c22r
gog1rp46iOSKEvhnBKmeFttA4Rj0eQPuAggjFHI3VPH17p9kabyIGhn/zp5fBWN2
TWW/N9gGk78AnJwPon3aG7SFLgMt57Q9bymToQGc5D0otbbPtB9rsUhg4O2RjN0S
Aa4QpszRVDQjetbDXRLrXtzDn3WDsJOPR5IEy1zKecF8A7n/Jb2mWLUQGRd5Tjl7
32wbiJO6x1A1FtG0OKMaDjxhYDXvVkjhsmXCan3pmY1tHcE0l4qc3tIMtAIE1TZJ
YpCe0bwZTzyJyn/lQfk8XCO9TvYtF+kUBMYW/T3I5j9PRxu1G4q4sYar0pJlXpSk
KVkz5vpepuo56j3Q3fcoeETM1ALw9eQzY7ApIypzv2QshgpaOLY4oaeyEjFizMdr
oxVfQjEb9o4shRIjH4IzTa7yIAiWP7Dr4NfZTi4bAvj7sPYcKAXc74EzRHSM//fE
Ii/RDS5WA9XboVI1dMnk+lqxw3bkyUtNoR+G3hwBjcmCk40KjXg8wCUstvzUQwRK
MMACXu6+5vvV618jQprJWYIKO8flO6IFYMEmat2+kvZo10nqFSOCdKJ+XsdAu0Bv
hw5XoOL0tOhPANtCiGNw2SYcMycjvOKgYHNhNsU3cpwopeUvf9xwrRa7ub6U6KqH
YjZXCsqxvu78L67xEYfcDWuIk3Xiw7HVyia+WCq+81LIdWlwy2Gu9Vf3zfSorO4z
FFfuJ3UuAC6fHEX7O4Jtcw0332gdQ/j5F9PejG24AVz2U1X9EbPj6fwNQ0y6E4Nl
P1dQ/HSGqgnclrTRY4MM8y6bjGLELRIvaNBZIBXHY/sxGFCAFEMDmJUNOW3GonsH
K2Xz5lIOSTC2SMm7U9fATfIPVvgyleoJ5cyi8puupkYZbuFIRvULIrALSgXVi1/P
LRII/GbQOmpa2g0D/qOmdw7HqQ2eMfZrKY2bZPdy2zQhxs9wVMPCQLL1NVe/HaXI
KVsMglpxlZtdiugzvWpkJ3uo9+ayZqGPQXzu+JD50h8iVIJawy5gPvwNF0xUqTzf
Dn8hwSHoblGmqADPBAS+svPBhWD0p02IEWAmhYKuc8Rdyt7eu2ITrvD1y53MW2aJ
7D6PRbAAzEWm6FaLpWMhJ5YSqGQYJUaIsvv8ZL4t+e8E5/WX+jUOdaF0NMqctXvT
pV4AlVfmYr9xxbhNOTjuIieK0QSGVkQKNn46bsn48aaDQjB+fmdcpxdwRmOn7lkv
/Qb+ap5e8hZUlxgrWb0CpMZLmpqcroEA6Oj2GMIPIYANLMGGChjwDCdXkHFpChZx
TZmzX6fcZZ+49aUgbZMZqRE7CTGzJGNa8R6AspLEOI9NbohE1mnIipvjfWWnrtXS
7VbavLfBF8bR4H+dcMAYS5MKVcklRE7yQd+Jf+mNiyydvSw+bMyLf2u3/m12G2LJ
iPW86LW9d5YGBdMCRji1x5JUXfFEREBlrjgNuIpMXplx0d1sFSELx1hdvxJ8RLaX
3KV7yQtNBR0D5AIo9TLeyrKNqiGYMg+KlMHb0tu2I2IUqOESYLKkbzn0gpZjebN7
Cfj7eCwiaMvhGnDiRrEL7Op5bFj72QGuBE1suVyRxVpEj4lXodEWmdJplfBQLroP
r0zUfm2csN02G7ZH6F8seF4qlE5sU4gevfD4EllHOn4v0P31o/S43pDY/iHrjhPr
GE3sxJEroW4efbHhiZK1PiyzTb9t49CnOWKkQznMhFaRWNiUF1oqP8QHWeKoIL+p
onIZF1So+aNuLWhKbXBzMQOd9w92DjBB5F/WC58wdfPvOcfb5Ywnf54af/YT0jXB
CWNw4LBG1DfbsxVMvW5KYrbt63wW6bO6z1nqeTYUSD3qRP0WuyS8w5dD0cb+qyUo
Fpe/Rqy30gDgEFGJf32cP6SXAzXBGqBp71poJndjzMX4GJ87V8+MDob0+I03Zkqw
IfLl61/n/7WMAwdjbKb608sixR6YxbQJFz9jhXPZtv5qNlcgP04vfVQT4desxJaI
xA30/eyV7BuxG/AuzLP2KjyiT/M8nrpi/lHdM+t3tWmbYbijQ8cTz5Cla7S8v2y5
BV3Hok3eipCNztwKVHnNIH899sfHNmEm7vQ6Dz5wW4q2k1/XgxftFWJ1LERHTEfq
97iqclCLlxj2lYR5MDr/ARBgPMtw6WuOT6uwfJnnRfFxFoIrp6g382Ku8d4N60qW
KlcAnVOkomBQpUkfaqmx9kdlXex3ZbDv4Bd8ZdLuhQrbSP1uGnsZqftlCtxbvvqK
ud/uhSCBReF/Di1skE4P7jUfsjtsqdhqNco4KYrCEzwg0XwGVK8amxGs2Hs3G51j
+81ZWWoUSfPSsScaqerpr/UgDME+Eq5XSIEambJ8qw6EYZVegse6kIM4pnEdCAvR
MdWOYFLX5xrLj6POihoPnSHDqsbkZoT7tIupQGvJncUjEgHGxrMXF5xvNVwxhBBl
elY1tDtptm2vXtj+Y1l4Lx3CGGaMyaLNO5goY3q+DmFLds7ehhUvcbIXGKacTIev
pC0W7ewrVHKjEoG+AObbYfKq8aVm/9Ev9LHEwu1FxTpNyeYN4ux7v0U0oL5dZlwi
MyKbScjBKfmpoCH9T9/+HGC4sIMrZc4NkpcC/qtgNd7YYkYB0i+1Nww5U8hJKSiv
N1B7oZUs/OoJjqZhD11uJY+T+2lFEOYrNhPOxti6jQBECHVZSO/ZDoXHwV4FX96d
FR1G49yxRqC0jJ9c0SzYFjy6MBZenNKfTnO1Yi1a4v2LsueaCaVKGMxtyFqV2Slx
I0TI/6WgEZtV8lmn2BjM18Wq8BA25wVyiE4udjlcxgDhZh35aV5zaNjuwfKHQGnl
VeU4RgWekAJxQ/NTy8Uzu9LvagYuwcKtmbb61aII3eZXWORc0O+Dg0+ug/CkAn8n
mNhXxJCTh2qwWiFuA1o6jXdg9hpojxkODqUHkVVaLCowLW2etDiomab/K/rGEK4u
kHCj737Ol6S3auMKGpBmZs3Pc/USClrcRZCFFDJVbzjzejiNQj1K6JiiRRWOtB04
/hr5X6D3xZh09QcZobcHzJVZRWVNajO+/d/v5Q0gKkkLeXR1A+p2P+h9az2+WNF+
hz02EIN0hhmTKlLBzA4NsE8F5/cIXJJgJFDv5y0mNvN0+1SF7J0CHgrUQRL1GFqE
0or1EVdtM9+YthBnY4IHYR3wutRkazyXo5ftTfjsSuLDwTMZcFHPn2DSZTfyqe3h
3RWW5IcUqO4BZZhPd0zuQnXUQ87cdC2JQDrjJvpuYnl8Jie5rjwQTffwSgReVxSu
XlxF0vlmWGnq+jV/Amf05PTtvj97Pez5oAeoVM0SWNQTF9I8gfPlshPG7e8bqMOd
IKEKP9BoqTO05S2Yo8cmF1Ln3q8B8vu3rH1k3hG3hWJELq4lJL8AgW+dlOb1Ef1L
fYn1etmco+xkIm13Bg8rgeFD01OVo3K4TyovUcB5ghbXC+wwkHZEM6ITdT5N4/Ej
wxO6phopVWRUXQQufNFZW1Sx4IVG680uosgK78KVwvQZvPDJrZtH153p4eTDy/ib
amEwJoNKib6XRn8d3jYhR2jxs9tqJsLkLK9l7ij2Ncel7PgojDC7TXDbVYAMK8rk
gIH8sdiLuY2EKYD1WUyJHf6qczBc+Azw2mHZ4Yo8WQtevU2kIBJNVubVmhRWG3La
/1WZgI0RVmy/lak+0tPXg0wtbGVyDLebpV85Iwj67rgheReO0rWYa49vVpv+fLEP
Ulvc+618DLAJivrzbiIbBat/tuvFbJvGl0I2AVeW733rnXyVXunTsdv0JrrWJGxA
eNpYpDIhYoq6BnoSXobXRhWRrAdgroAOvWXCF0QM5XlCuiUvoAf5QgnMk87rd88N
mrPUyQkR8wx/KsDlyNN4aNiP4z2CjY//NDblOenFOQN8F+YvN2ycm3G+Ao/4u0kV
RJNNS2KO4cgm11TyHCpki9uwQBccGr6UlY44LGUGbpi+1yqIZSH28mnG0xaDrmH/
4ukoaG19Qb1D5Bf32aA0AeLLp+NeRZumoGXJJIsUy50FeK0DH46SW1ncP1wqeEhU
LzTueDXQt8lGFkrmHnd7fkXUTl1A6i6jrjsYsRCRa4PowQ6tftZyfXxyva8J+OX0
TNF9ikcFJ8FpaorqlVni1r0TMMr4xHOkmKsb+tyVjKXbWUfxnp7tCLWKY8aBhSNH
M8O6mWGRvh5yLVJ9oMm23Yn00WZqRf6zrqYYXH/yCl0TwdMhg8OWwGLK1j4L9fFU
x3MIfPMEtIQtHTI8WWoJ+UWrYhGPx2o444aRlOLsHLCpiKS0LzFhs+294oi4JlCF
CW8OtsvyHlUmm/q/0Zsbpwh7zKK7eHVAnKo+POcKuI8Zmr14xYDFm/8NAyh5S8wO
C1sczm+2j0cqlfqRbrWoZXmdExBbqKaaVqZmAXMJy5uwd8lqeVBTgm/qxhVhcam6
aNPkMZVB3lDin8VTgHJ9/ho8i2Sn0X93iZtEnnwxHdPwpjoBd6Vwj9riCyLB7PGY
tsHxKYdvU4KC+WZOlR5733O6SFcFXLJxFx3W9IJHsxr0Z7U4t6xQsDAK+SnBjUP3
87mr429MCPIg0kWnBsl/qvfoXkeaWGAq3aGa16saofR+RIkpDQdMvDp0l1+MzgDk
EsVXxrL61NWs0raaYFq3GVkcZMuSXmiR+RAHZYUsdQLGnWbZYFHip/t9xvTOs3H9
+8C00EcFvGDux8gfBfHUK/20pr0j1R6LoNEuAw5khQhWE2Ay/V84796ZZILDFIWD
6/kBRIQQpsH6LB+SV1EE8b0HKiF2RybMBJseWqQjJ+FO9fJ8/MGTm7lJbiDLUPOi
Yrv940n/Eb7KJA4I9u/lVoGyqvmsmCJP2eladytoExM/jfZMffdfwtdeXpeQMqZk
H0KPFCJ87vntPhqhUC8xRsiRoDEhRuJCT+6I6rn9TIZIzgsU8m5571BPijVUMIyd
mVh60YOzsEthSMrlRck3+SMf13FOUvQVZaSXOBC+bnYlVR4TWHXWshCMw/UNlUne
ij2ocmqF0+PF3El+AWWZcoy0CzGxib9q6pr63yZlvYGeRTll2VAidyMk3ZVXUk55
41zK9Odjf8wKn0DwqZVeblVD5Xp7xaP3ek1lq8eqyxCs/P3H73ZCdP3eVhkT4UDb
OugccDmEwTW3p2IJDrTue1QsscdjHA2Ejkmxqm7qzSFh87P0JS/FSgWE8EsWAbWk
OjQwxRLfhKXFoHUHj7zL3jMhtTmgxEnkHhiv0j4rwJ+ecigDX2xlu1ek+ti80CaJ
EP+/KvgUe0iN8zjAB4ei35Dqo9us3xNGTSz9PcWq6wtxY94IDFLrXZDlKGH6McOl
jqHJI12tUapf0VW7xhe70E4PswYGmpsO40jnBL0oQF0walB6BBMf8EFfFaWfv3de
f5R0hhuZiftzYaarAMS41ojBhnW7RQiox/AyQK6I9b6YP1OxYFtYJAzfpypZkSgJ
edrqVskzKHO/CHImZrWEBGz07X1kFIJhkeMGCquq2uySarN7rwchvqIQ/EfJaj8H
h2B+DonpPH5Cy2/IEWiHUZ9Or8jq62ElYCtc8M+loPa2/KyiEf4+bD4cKAnUd4RX
BPj2wBR5fV06ggeyQvWWQFbQHlKDadmk5x/my0hs85/w8eFmqysVOvcBV2a5foz1
DZX5M3sdXTg91YVBhIY+/dY20UMvSXBfnPtE7+F7b1UDTZIv2MM7tNJL0SUSUY5s
cyS5+ljWZUflBjtdc2Xr+iS3xkFblaBgBDYuwZO7V8GIpRK4ZEqrwfQbFnNaP9x7
YeXEWLm+2w6Aaj4X6uZY95157Th3oUuuJxJNs8KNhW5yeUqUBdnxheXG7MoulGB0
nWsjwpfvQ5TJk3Rh/GUGLT7z+wSmRf5P4hxkra5YUvtw564nQek2ZAFcYPeXX755
KrR8seF02uOINpuRUFsv/sCkKFlUY23XNlBvmjOFS4RY0GhLsOKWZdoHRdk+NJIc
RLE1ZqQMwPXFeKlF+zm5IPrn+Z65CCNOisetWHOnV8q6VvEfQjxYbOIBsLuOX/jA
ksJ4HAlMlrjK734uw7dnDv6Fr7syFEB+ubBP1eQdoiRgQmI3I6YVNnC3aII0DMm6
yrxwph+Uuw+rVrUUaQM5rt0emJWrGcBKrPXXlZ11mtyV+lROT2G2zq+DQloacevP
0DdknG4fnH8gUC7ivIT1iYhNojlmDEngEVSVmSo7nn24ONUW2T4TlsXaG1f+F4VJ
nVpYDlwqSdeIiex7nh4B/YNaAtthxOllm/kljHXD9kYOtYj8C3YNpJS73RL4Jufl
B1Q4StrUFZfomKVrRGi/PSuolQ53lyJyRJIlzXXoROBOWPefsEbkXEfaUm22QzWe
AegX4sijjslPiC5lfPAqCxx2g/BFTqDogMlrgosV+vRpYzJMsq2LV0Kz5RV2czdw
+PWbjPVtiGiHIE0Sl+Cp/AP8PEe1pd95h6bBx2kWN9HBhKQzTL9nM0zMlK6PUf+f
5zo2FYzsQTn9GGcuDjxIT58i5jvN4sdyjzVuwcQdQNbLsBPu68BS0fybENGO/vEn
7bkTpfniF+SSB/fQ4cfSqFv3te7Pezt9RGpQe5V7ME+6qCOXMPrxlQS7xD777c+q
WwipegD9kYS0VK2l7ofwc3seedlKQddL1yDIYvoamN1bPreLjSRTIQ4mc/9sRREa
EgW+MFsJx/NCl/8C1I81IJi8BSSUAEVOclYdts5NL5aAV8ontC4zYKIKtOsdWCOG
NldAqKrcbqfO7b4/ydY2KFGM4FuqJ7ntKHOhxXeXMUJmbNlM3vYn46VzHtZRHvAQ
uCVs5Z4m/08FMGwz4Mb28j6JSyuUPOb4JToIP/HxGdLf7soFudewkVwFHQ/q8fqt
MM2hYktqpA7DtE51sjdcinrWZhHmoDy61geWCxNHXBCSPvBvlUudnx3CH+Wf2r+4
ViPKdHaSFh/d/XUx3TJcP+90I9UaCt7aM6me5sGcDqtI72sIZyZDqaroepn1Z6Ln
An+BBAcv7+yVxUIYu5D0yZE0wqGknRTANUgezjXJwgMCST2ycX7n7ZoNCHVd75O4
Hcui8aPQK+ouFSrrcuXMj8ruiHsQKJQr+W6Ohpp4JmheMGZN00/oeN6X6ZDmgeWK
xEZk3LUFXKvxf/l61h0wLD5L3wips+EzbRw6+agD2t3dCwvkspsqDrFEbQ1XMsUJ
m4tt5pANBezUm3utbDFqiATagDNWYw3FZCAGMlzQNd7wqlobsffaUoXZiDacJ1Z2
qnAfXVEzmAmPy3ot11FyJjT9KTGbJnEW2fkc4MXPPDTpsz+ZPlyXDQ6hA5qachqq
QrnqwOb7C1cTtCSY5MW5GpVDBfkxahhJqBNPytfEMwZZmBmZPrapY1sjCPinrb/L
PcTNND59FTED6Usd13XlDFzwUeFb4S+aWTiQCb84Wp+Wu+0KOL1Hj5Z1WUK1h3Ow
pASI7QOkbJO877n+t4l9os5TsBKj1H+p80uPpY6fH0VUutBUkSFQr+CHgj5LAUuD
kdd90+8yydTGsLDLrvhY3rnH7i3HleD4C7GW7iwK0d6ZuHBhgaTM7UzXbtlAseLa
Y5QLiIj9PUwS+oahbzAklGGwhB6wQ+Zi9RkT0xGZ2duhNCtrpo8a+Enpiycj+xcA
KzjlkUyEhVv7jh2mpnLXeXZGbCPsBlfuIAtIY0PikvxviiCyocZ+yX72AnMcaLE1
IKVZJoKP+I3XiuFZ0fx538JnCObBTU4vyScK+e1VlVvl4JAM0OpNDnUdMmJ7EZD7
QmlUeqF5y9VYH8e1GMzFEY9e3c7hRp/n8uzp9ErYK7vmOvXUB56rGaJxgYgiOJGH
xJw6O/DfbPlSjbqaubnRq8BExlviU52qJIZ6w+7qWCInntjDYVcSkCkU1kDQJQ4C
eg/WH2D8Xjl1DJVBBG8i1tItwoTm1SDjypoFl2qnZqHmmDomAgP2vDLbU4oyATZV
2oXhU4gTdYEEw3ctwxZJFTikOsR295afAsJd8DYXlEQS/4BaukBKhYCVMGEYRfnE
SZZvAXhkwr+KhLhE3BjggUJ52LGdEYcdt7d3LIHltehgx5wpB+PBiD2Jm4nVAAPx
jwD4hjPCYTTdkNJyrxPNWoYUtkRYlBbYRxoRUbTGRtbdPj3tNxs6UqDnrcP5XNyL
mRh/aRQ0yvo2Ngmiehn9lQG4iJPgM0v69J8CVjJkZSdSRbTQttaMVByc8WEfDBtx
UgNUmeWR6pxys/z2sHoN9LyLESfY8Ojqn77JtERkBx/2qX7D/j702uGi0Cnr2zCr
9DBKGZOcK7EXKTm9y8ja24eLdgbiWxP2UslbUbh6zH1rPTOiqEK8ieoOYv8Y450x
uj06QWJgslpkGl2akiOgQJKKcuZ1S3OQqxQl10W1/sfpNGZbR8w9heZslnj1AWWM
rj76WlqLUi2/q+O0YxUd3Up+ecTn1G7GNjddue26GzgRaXPcXtAeAICRzs3uwyAY
z2lZav5OOvLamxUIEV0nUb54kzZ12EHP8dMCF0dzSCPX2xl+U45Y7KV7lybisOJj
0MyEZYMIo2RxgiUeCDAYmsUwNKLDjT6rgZOvz6KFF4iVT2TZWSf7XinIP3xo4j08
G2flZOQoXv2GrCs4FsEGNLGxVOeLtSiKmQJXI75NYIyCfnyavfL/QfvS7Z2Y6mby
4tna8FtbKKD8AcjRiedlprn530VRzw5hnRI1rj+AvX6QK6aC2LK/XWQmVGda1zXF
T7h/75eX6QxaWqyvWE3Nlu8rB8CJOnSsfY/J82HqWAxmisNuScvSCcje2QfL84R6
malYok+lcQrVvgLvD2zj68Tk1aNR4K1m0xJngV8bwRAwgrvLz/WZauZoExtG1T2i
EKkp2y4qF0QoA4UVwy1LQROS6qiMrlKzsheLZLJ1jcBJSw+WNNcoPraauO1Rv7eS
T6IPTh8utWXQtgFNicv9fhWxfrTCWddzuLpEL9eG7C/43UJ0U4HpELipbD0cHA+F
AL46bPnz+B+1XU86rja4zzlQHFM2SEsugHGDuyqPX0l1riOdEcMYFIjikQBCtBgq
WGL9grTXe5x4dfLUyHhj/hnLTO3pWlzrpYZZEQ43FVpGQEfgtd/Ecpa8uabybLNG
Z34x15Wnk0+oJw5X3qVlr/c7opuNjh3itBsQOc37mzZ5kh5cnxnFeDm5kiKEzLEk
gta+2ED4NaOeqdacILROMhLi9QYzmkn75d989NDAjdMGSK1emjG3TzobMbpNksi/
jRsdgjBg3TSIW5QG7ZNYXWQptb7CnHUreVg3X4OmmZSjEf/mYMJ9f2Qo3aIlClnr
mwfztXLnFwPBZhx+A93HhcuEk20dsfxL1D66R11NjginkDGNXBZEe4+KWz4ZOdJ1
evxX+7/f6EptOKRJdCcYPYtXu1owoGDk4S79g4MzQzKoVBnP5PgehCyXgz1UvLWC
wZFkB67Vmah73cncUc+A2Wp2M0yDd5v2S6K7BdjdSxnZZCbVGGcNjwq4ZOanXBIx
bNdJjzV+2sKRaL+2Ba85Qj1uFk5LRdKSjatRLmdPtVLAH4l7IrsqZ6iTfLlN+B3/
qfUjmR0trTNcTiq/Eypb4dcrJ9P3yTJsJG7PRl4SxuB9YyZLHD1JzVIX7158Rnje
IML5RHd94oAS5EvaFK4dLUutoCRivV733bF3oehVicPQcS5KMpKCabTF/ygBZo0o
MjZArDp2jJgzx43cSvDXJyBtevVr3Ncf3FNJYLAoe3Mt/h1jRRqQ5jVm5O7DRLPK
4HIBSa5ZHTm4k8mOuw3tvunfqMdSW0fh9YKPcn8nHRlwj48NRkRLxuPHQl/Xt2Pf
/Mz7AXlnVYkz0agdgwYhsKaQpT2voAGQveseP5woyf7iBnedXNNWqCUn6DKOhEPG
XR3bCjKH2E48GHgj1zIBqpPtZzv68C8RnoGW66hw700j3lxDOqXCO96HowKfglLz
xunUY5fBk/irpMtCN28eUdC5Ny6oz7xAg55V3SdsodUenHfBv3+jANOb4U7WNTTo
xwM8TN6TFezyjihEJuGQ1rX64VSFCH+Da2M5vS8FYlqDCwMYVmyNzBivw0IGkxOZ
F0TyJ7mogvYrv8geoLYQcW3yJkuX3cPKY5WebUYIWzLa2TP+Kx9PAeW88wNWJLIe
KherISEJYkGjweEaxJE8pa7huVZbeALd4YfDgbwUWLuz9XDpXrt8/pmPMWj/DgmC
Rpx9ypXYYUmTak4vkuuGjD9f8Qe1BZpLAk4cmYHurDwDEP4BRHHD0R/EigJXSXcB
DBwkP+z5tlRflYKpaDNOB5E1uLP482FOb/SZL2QtkvUQ0A3Wi5+8J/KnoWfZ8v0S
1Uhf4jBYAhw/k9sSb0USB4Z1b5GulPVTQiNILlRO5SaPXynriM/Ci5fL0sSxhgH2
bPvsjHwKW/8Hf2v6s7bLnhmN4OBpEKbWdS7ZO+isQEpqcB0Em3S68968+q9YkTDz
rXeqcSW6IfkzfqqA0Wx4iKJMzjn+tpWw8e1JUhb82/VuKu3kcL3BqRJM77apZ4Gm
xeFBT8JEHMrFN+N4tsvCWuk4rOPEBIPa7XtxEeRebsQwa/BnA4dQJQ2V83oiQ5O3
fq2kV1ycUoZrDmDOy7lWCygXFCvqbwYuPihvwc72BKSyDDKnbiPqtrHCvQmOdo29
SbXuw2gpYGkoBwTRs3iNbjllkGPRjJiVleAn5TeQLlfX5kUgOFn3bkbtkJHgptaW
zylrOFUS56yH1gdznul9PfzIvW39lWb20QLX+DkbodLAxWh6TrUG4d3LU+78gPnK
uicubJVrl5sXxMIoFBoIzOZptBAECbqt54E13qgSDDGOEYSgdCaZjCLI/Qwk6GhN
mQsnr/eZRqV30XH4cUKt5+AK04iB/LU231Oej+TB5xIPIm7WLFY4XRmAAzpNiQCh
eddU9umf7RDZoLn/ODAxHf0iAiAw5CNM6HuRsZbCL7oJG8FXAI4xa8jR9aN7CkKN
iXitsvY0jBMsHmbXGc321pN0DDgkVP1KkQU64wc3HcQPrf0wPXd1skVDfq3Kjcw6
/Kx3vUOnHMqVkYbp7Z7TZZKX8KHcau6YWaOqYv/jHTsLAX2BkJT5Xi30Z7Rw651M
CxRy/84gtJnnx4ETcHn3EBk6D99NrSQqKlUSbO0sLh4hJ1RaFoL5gmQn2L6Z0C1+
LV1HUSRQdaVpDQ5blkRITU0rc3L0wTPpfwJUmnzubLA8xqnS0J6Ug9IdDN0vxlCG
jbkrZ3eVZA6IGmPXtMvb5K9FFtfTTytJVqb2L+APfH2c6sHYAJ49T0kz/hIcX9zX
g/gdkZWfjMEcqX3YgbEzR12nVCgWNNzRTHieoq0ijAJ31hDwL+eC+7Otvq5ZRBvv
VMAux1827vwe6L6rNoYmFzgygibIaFrPLjYvYdZR88KwGaNKW81hykflSvZLsKKf
PMsVfG+Gwc5H4PXUq4qfOxMYtmZlg7KriI3g+wPcuFFLz3RF34N3KC/HxwjYB4FH
2lbAH7Y1JqBeMa/yssGrVjptRJKHZVnPgT9MZ4dbLR5nYCscKqDLvLIwj7UJRIzq
MqZNQoBQU8bhOVzIDXe2kTxk4Tda3VFBtUWh+28W7275TEXypjx5c6dm4TASYg25
5wh8IblYcujBGFwDFHm+n2B4dDnBKA2PQ+YxZuByRekOR4jykO06s+E9RBMsMbBW
ip6Sf5ItF60RSjmUtAWw4mEGL7h+ZxpBr0cxPY+1pcjnMpWMYrrKpWxm2ulfz7lx
w0zg/RofL1QZ9L4rsdeZjlRil7N6oD8Uxo1qxiqwT2GMVSK6maS4HnK8Z7CNdUH4
VrB2U5kFv4NATv5Rof1eS1bIYqUG6qpTxvTzj5JGjGzrveRhVLnM9or5vk76rfp6
ngj3fpOR+bARerraTbAuOuxhQqPSxU1VbVlL+a0HSKQW2lozDNKOpY+b5DtYBhcs
Vdn9Ifw/Prpb5K8kmVehE0n9enIggD5qoXydkD5vTY/tMltln3N3r9hJm+BkzyNo
Dx+4SWPf2mFR5PE/mRREwMN50w8Bz5/XJXuN3TmwzsmgYXdsC3eoQwE8tD5KbWKp
tV8S485zYLRNLBhzddKims2p3mAwwK1oI0eDCFBIrHTo2zw3mJvQOVvgMcz9dHWp
yQueh83EOOabVZT4kCDbKYr0PTQEw+m++PaBQtWXJmFxv9hK8b34HYCWqZkwtFhj
w+wC/N1lrnoy8mpmODY7hwhrzYeAUn0mDGr24ko2wGjBxcPzaXXqvclviKP4s5Ny
LmNZ37/+5q7qUjVI9BMhcuYUfizMPEF64HX+t3nP4+30bpJEkfygKtGU4rgzeyGz
pBm8bQBaoKbggLZ11dJg6ej9gGC11J/wXrjjduV0z3abUGW5bQSS2wPU62AjAu1W
oB/GrsBvFlx9UTsoSqgWB9P5OCkKg91xH3hEL2WbkqqpSJv5vA3Fpa3uA8PaX9Hj
qU6JaFYCGZrgtknJa/ht9+ge8WZtFS8CLvTb0vXEpRWXcFoMnhbl3M3bC4MYsJJH
FtvJtH4orw0ZBTPyvehKTveSudTfJYEwr6Uagl46sSzh2wqKmJ2WlX8DJPRqLlgy
i9FCd5k0OLlO+9oOZ6XAoRN9i6ZElII29dW90mc7YkpfLDrRSBnCWMijmk7fpiqV
gMsi/cswqTsJS/U/LNueh/kkLKdk95u+DR8wk54IExdk3Cg/oT45447iz1N8R4Y8
CC0OzJNIiUQXr8yLUvEDWNMtQQm73nFEWJP2XkQiWykSBldSOQTjNNAcWjMRM7BK
4C3to2sywkURSSx4CX76b3EN5ETfY9IO+C/LiTeelPVz7pEq59s2uMVl+3i03sIq
GLBwHyFLAmKbcYtHs/v6qSxfYHPOX+o+IV0V52DFXiTCYOpaYUqjfpXrCcmYzVoC
ZsL8fViANvQYPfdHIw0o6bcF4jxs2HcPF1PbFvdVx1j5ctmcrNwYushFZLFjDJ+K
L4SZFWY/+s9b8Oc573q11eybgolyJdh/aAzzHsIoHM1m+DriNyUoliUha1z4+LWh
fLz0z2fYrYMAVHfZewet+T8oTV444+1kFwXd1cRtACY2+HyVpSqYMCa0lfbK8bS3
8nFBHzJarZECaiWGFoGvoUFGVtNczYwdRofNCL/H6CfwukR+tXb1k3MhM1ICNRgm
hd4EkE6hqSM7EORJTJttIwWzebcqViPSdUp9VV7VQ+0d1nZG1SN9dXxhC6xSVDCk
jA6qr3zJNJmiiz6lCWOKX21exqCNmGmi0pdRzueuNlEtBwdmllibuidu+nju7t4Q
znZFLH4JP/SRfW5iQDWz2gQXWk1QDkLTFWwGCuik7NSdptoDI4LiN4nCULcNs4Ja
/yIGmFPIC17iqyiy1qoUS0UVk8i7JP/gvxOWxljCCbP4g6RJTwFnXXTg9+t5qBYt
2Ll1oXwi8g5CgCFtxpR2aLhSq9jCjx7aZUWEl0DYKTsDCHRWiXxJ8OD1GXVzk8li
T8YrIgNuPit/+cei3AkAlCpwRQ5A96ha3oLi71kiIgJ7aw7T+97UF+/V7AEJ/i89
Q6BpOlGFGXqSGEH1HQcwEBuFuXS1Xvi22L8asAt/z6vPUmEkxvP+Qb/QO3PSmYx8
TlPmeYghyktuh8MKCHhAXKmypcadgX+Tvx38eEPrjQkowmhONSvWm1NgEpgZ79ll
9QGWL9159bfAjscTAJ7onx/enFHlwN43x9w77wIQUkRe2BafI2Tm8HHrx2TGlC2v
4GLW4nFHTJ+TpQ2hvazFZQLEOVjQictcTGkKKpazL1WQNDRdbbCSbuuiws0WKRb2
pvH1oF4b5bCPTREMTEBc0op3bXxmMBSeWCMVAcs2ItKOlQZ7uFyNjaEHOcmvnOpA
/2Xy7UqxyWJ8RCSEm9l3IECwp99TtuYpUFp5o10oQFk21ER0gzngQNaSPVwH7vtL
dzjBCyNaaYXWynerrvhSKwjSlDlTK2lSY3qRE2bG9YT58PNYuDBYC6nljROx3BDU
mTtd9BPeUAdj56deYp+p36UhNzgtTma9Yz8P5k62kNfDrprK7uBZyg7oipPKDTQ2
Q6CkPt/mgzA4nMQeh7sHCvJPB06CJkMFa9w3CXcY5JRhSm7akua//FKveWINcd3p
8Zeie5GwKoNFVlLibk7dy8pjtccdKFWf2d4tV1N40oHw1/IZmL8Y9wVIn7P9H4MX
Hf/MKlmnd/DWx+v57K+pwtCsbZP5UeX5nknQBJk4Era3dSigSVnsE0R53pO8nW/1
5FgKSUXdreqQvLh0NKlOrD79o1uInXUaVgkr882ZQ+Z4t3scE5jylmxBn8pXxHUm
MJMeoQs5CeK58VFqb+tk9K4cVKM/9aY5oCeD3czhSdaGtsg3UUWWUWgnef0wzDLz
JkXu+AaNyGBbVabHPeB5wTAaRsKr9rA4Lr/6kTsUY1XosVQ/RHJWRcBD5XdFo6sM
ZRpyle7YpYdarzq2kfdW8EnJfbRANG687WXR/t6jvuyXCOX/2wb07m2q2lv8tXrR
ga0MDVz4Uuh9lnT+fHf9Wpr/rqjQXn1fcUC0KVNo8uTYOdYF5aLFQ0ukjTXElh5F
/GN5Hiug3ZP6BCcj/tBPYDgkMN+QwEHIu/+kn9YLquwzK/AxEU+TnkZM+x4hh+Ck
tE6OMdCST3unmqr32O1ODi2GAJGWKV8WcTJg0SJ7VMwMAwQ8dkazbrMiNnfHT+57
U1wF0KqZhPOL9QMeFd8QMah6PhhFmABVNJCaxrOO3azfHO5S2piTREI7fGVkA43m
2fU1742tSiIQj48FY3kN8M/qB61ovT5ThCHFKQunGsB0sV9neq8QDqdoe6jPhMqz
+bIiT0xdLctmzoS8nj/nl0e2yP6nmLvvbFdfT6h/0jDZ061EWlxOFAWl2b/VJMiJ
WZoqDY8ac6gMJxteQn/PUtN+Ov//J+iqlD6xnHQ8pAX6hMCYO6bjxdpuKBtSQVDs
cBP3jMPCXl7skpAWHHCclqOh38dx/C0FlYhdDdvDpGTDQE6nJ7kzLTlsAO9ViOg3
KBECPkla0/h/PJPE5AWYy2pTLCud28RtfZe2yepiGmnXPbiHLbN5i6gynZH7u3V7
Nm/HGDA8k/9B4aTLbJoP3GSPkch70WLlEu0CvCZCcWfsMMiUABw0k5nITU6Hoc9r
r8x8vfnJCZcY8Vu4at+THmgxUdJRmI0cPu95CVETmDeSc+UJ1BHjpzRAJTzpXU32
XvdZk9VNZlUh+xahP2lmmUQRms9PUxCq9DvnXTzvHp8FqLdeTGz2wrJP2DOjulhJ
d2R8FrToaKJL1BlQ1TO28SY7iGLEHXgxUNzEUQNkf8InogogsB27OyHBF772HpmK
o7mMynY6eoXvdtL8I5s6aLnLAjTwc+doNLUz42KPOBlzomia4mDYCxaj8h0y8cJw
MGCqXHMvaoTIcuJ8bmfVP+IRuoNVaA9X0h9weFiEN9/WvS40e9BW8A3cZiJyoIae
9djjnmwLHpDx8OrT2cPX3ov6zLakpbzTv00wqoEv+9osS8BKpzr0XoaMFL/wmhH8
oiU1h3kG7scL9+jAQ3KpCB+BRBVjwiCfuake9Ro5OqprUMJBfd2iW2nfb78OGO2W
LqNFX584B4TnPIxt230pMo3rW7VMwEpSzyplArw5qXdUw8YHkm5610XfmEkQN8wY
ndEy/fq3Gr35AlyItcqM6+HrGCNiIsV00uwuVZF2TtfEvdT8gwS90XdoJFjaslR0
28C1dcvBK+OAjsa2hFFG+TEtIwdMjaUiiU0dK3l0sdAHW1gkHCIqj3O2R+lnyLAr
AvBLkNkSIyYFMnzv0kv9PWyvubI196C9y8a1zv5RBblBsWFCQyLqJbZP6kd7H2qH
DigIa/qkqG5vRb0lL9d7bQ2TrqKoDlq7Cikv5I75SfGcJtRf2HuChrDfOrrJTf/r
hkSn7F0VYTEmxuf3HF/Y2+KLEL/zJu8azhGk+nEuZwRRzeJ9TZAWqlXh+pWBMDSa
V/92KbBcWMj58+5xkqEfCmedL7m4xlW6jq0GfKabwN2N+4YWcHnKx8UuA386XgqC
lcH9ajUKBC/G3LGEWHZCRDVfw2HW7d+2CITLO1GMSrv/jPZZ3uZGhmE17R5nIumf
bfngzRDiF+z1E/I/KXLWnGjn+Ye5M54prKnQK+HscJi3Fe1L+BX42DFaP+5sloYJ
t91/P5Xf0csgP24KGAYGSBpJsuGl/bEpG89qSnUuZYUlfMbcyb72QSrrp9ohT9a2
njCvemgfSfrLPG9UaOh9PzfD9qVA7N7oGmphA+Ybi0UtL1t7pHcfMWx7E2nWlY1i
awY3tW6m1L78tx14BnaZWjq5vlPo/aKopLqYLaFs4XOOKmCqKAIgYqfTm/E9qKz7
S7KNi7EJR5+gxX31k2tHSiPlYFxut3drArrxFXx5x/4N+x3BP2rrNlLdeqyqXpN7
8vZF69moiB+otRMVIu8NABeeFHHaLUjQE+XquV/4hUAjKE7ugx1+TnPEIGCUf+x4
/tZ1CtYoBzDijBJkzHNLPkiJeJFjQZH8Ora0E99HYQdgkdda0TW9uiargukReZo3
thvHznaFrMhpaBRqVqCwpHx0TOb2JGPbnyfMR7LwshyUKPNAV3I3bN+LMtCXSbbC
9CHhlfKX1QBQXii5oM9x6/fyKvTiwFKQPOu9WRWgvBvBejPjhF9XEBKxjGIRq7EP
0FUCPct7UQKjPUPF2tCKyEkva0oym5Eh2G8orlMz1203nrN11g6GtapidsPkaDgH
sm69f47Y4yB9eHouAigGXCqU0ZOm/Ks+pCEIv3F5LedlXmwumvk9fFS/MuNsNRjK
lVGgKG5UaQIu5J2CsiKb7HL1XanXVVl2/1oPO86h8qJ9fHvgFUIlKTGzx2dxkKXg
AEypR6sCsiLNLHI7xHG6Gi6Cd+xGlBc4YMTJ5HRWDaQ/c//GG0SyoCHnGReygd/N
dtH9V7ZKdsgrAhMRmdjV1gr40FjpmEjdOXCfHH+9dN8Q8yE4WzUZQ/CunVu3cxW5
adzHyZDLJF/eE5GnID/I3pRPmk86yg4ehp5c6AhYrRBxBbQZ9RMDvVd2g9vLx/fF
8msqChcTI6o41mqtYcMUZiR/cZABhlxDy6HwxrU9BWop0xSkxpuW4zR84stkq0QQ
vFjFz+1UVoUA8qnbs3q6GnaEV+mDDOD7ltNZK1yONllkBe+Sxe10Qm+0nzlybKyk
24JVNfzYHhoouoDDaIOBu01/pwvas8+2IMmE7RO7b9TvWzo1bxYqrLkVEBjj672z
zcZr6O6GJEAOT0gPhgD3YjLGnETriHkfqz97Cz6Fz1BBlPDv/x52AB2LUW1mNBOF
RbhBsqTUt9B+/nl3aLPsvXw8+JGz7uTc8pnw5uyXIiMH0eDlomgX9/Rwyt5AspGG
5p+XZd/XpDMtSfJr6G5ZvgC8QeJYDzQljGr4hPWC/Sj0VTzUN+YdDKzReXTMX8jj
Rl9GWvhB9xSuxwPfo3LB2AcLB7sGi880O4n4bRa0cc/no//67T5cf4hK7Qge7HcE
HRIHs79hTNEtRj3uhB5++wcVmnSkp+wTs6lpW9UcasO5GC/BozAydZ/MwgSNro7T
lQjjIhsdZ8xFr/U1gcCJkh6twEgW+DhGrGahSuO8W5gH6RgX1wIp/nun0rIGJmMc
Fi2OJ3sakW6g+fUzeW+eedFaznp5jKMbOlFxIJn/YVKRsrw/iDP+4ESXvzSOmWHZ
N6/HXb4+m0Hdd6xmkUNdsbrrMWZIX4EKTHV8vmjKxQofNl1ySksUjvrnATLKGf4D
FdlaZoOhPOE+GrrrfiEM25uX2T1Y7bNiEmyosqH8OQjft3qESauzZg7lWiXJLth/
7MkMEgXeN3akzX8rOO7rxe0jyPdUZskcdM06LpS0KTWMAEI27V3mHClD9O8BCxGv
OdR+ja8PzKkLwPU3YJDFVqpQN1r080IJwghjdWUVd8D40qjbMwS/D7FDSUqgU3VV
rfu5UAM6TnfEzP7o+XDD+ib41a38qnBRYatpUmW+Lwaw0AF1ERb2pzHGmwIvMWMD
VonG9YzkUH7xMYWC4mHHOzNibDGKPwJAfV3ooVPnF+4bsf2BhTkHA49raA+FcVq7
YlLJnKqRVkqY07hoh8HCICqzDLBtBAQKeaPe6jIbysXSrYhPUMnyOhyJg250xJFY
2FVPUN2v0ALK0x0rU5A5EZtevEzWhwcp6+pNUAoThMi9mkC4r08sSdx7gD/vrtDc
mHUydKyB691ZKeBd/aHY8hydEb4JVPpyKDevyHem52U8nz+X/ySConCMnUtSbij2
4Gi+2jBFwtwyGo8GgF/2ywGPXWzVqrM3qVrUH6mh3Ezj9ipq01/P94lAQETw9wE/
WcDeKjfTZyfQmSHfo7OitYDU2SRwrfTkV4NdRM42hanbdGP6hblNrOylZxpz+Upr
veT1q9WtI3PkUVuclK2W1eMh/sd2fa+/7kO5xJvhan8YjSxdA805BnjiJ44Bn1Jp
Qee1Jb12Ju7YKeHW3E8Tl4zD4cyQDRHhQ8vWSPEBSkEJlCxCB09pX0paT8+LcWq+
NQFRRUntRtqRdZTk2QBWNXvIZl2qly5enQV/KCaih16wd/G3VRDBB/dMrRiafpXn
XbFmtiCt0k7gaBJHyjP+OWNx01NUSwmV5CEpKBEifG79YAYyNguboDMpOnMyIDW3
w7Rr7un0D4LhBhYC3j3yRbVWuwsgM2yAsPeHFHCZx0bzqIMBOFsygFeDJvyHE1wN
brItk1Fzw4dM/jM3ndgwX20EZMGfkKrhc3S58XuPDW9RbZQQTAPfYyUgpeUa5jPz
xcq1xaJ+Wn0Z+aUe10nazoZspSKEg6W+Mw03EuGKJE6soGvf/kVoXjySlTn0rhrW
F4Gs8+BqrH1N+6E1pGmDPFHN+f0Y1Tm/t/dXFHWGoBF7/EMOhsL7zo8vnLFpgd3/
FrKhXV7eH01d8iVkpC8dCdC2ZDTLT+nmMiyOriCWCfHw/jJIONdN+aMogaUYt4ic
RpyaopWEiXdQ6mdqCvjuA1qS+2pyAE3xvTFnt90SDaAxCm/B6DljfRtElEzHWrxK
7sGc7flA3wdtL+7kas0fGy2nbl1/SCSc9F0lOfFg4tUnTmY304c/pDOZ+J3bMZNf
ouq1GWqfBkMHfOFzslqEp130/Z7+CEdIgIR0cVOm3pDSJ8gggcw+uxm0EJdNSq6U
GeYqtNZTTRsMGut6v1K+P7X6T/9MdnJYBqGH/cQTFRJRZzDgvXhBlQmstCu5vXC0
Z7diV3/yFKtRgAofI54Bm3tYWcoD75ZJ4W1G2YiBbM5r681zJYkPA4fmp4J8srIr
V1IAWtF66lMSiqPvNwpo4f58HasLc/DXQfupxcHXakS37SqUAvlIYZXOKtYljRXz
cex/vMSNUGBZJ5YKMf0m6yHQF2plkY0GU0+JhOnO8CSSVMPbI/BEx9jLzdYcw/wi
uZykS6mrcry5wh63HFGP9hQOFHJZkaTxuoYcbzTOgeyWLMxNHmcV9r24TB4MsBps
hidlo3D5StiroOK6uS8hK/eO0DqnaLRDwS4nO4FR5Rb5T/HLb82vsHnSluFVb/5v
zH/UEvcxtbp2Zg8RGoJbd7T75+Q9urUuGVHLnugTtwfMlWrVi52efUQbDTDcL/CL
9TOhK0Ih1RiyKM9K1t5xnjjQx4NauaVBVLJTE7t3EwTXrfjxft9F6DfsmN6NGaeY
K0rmUysNxUxWC3X3utLixQ1P9KbwIHu70qIalk1UhPf6yhDdayVhbzcZpu/Qgq3m
Os+xXZKyCNC+QhowM+xmYIKWt2myhO38yNkh2buc9vZr32PvcKBEaOJrf9ZzZIab
yGaVznVcqUXbUisY77/g2zvTXXsxTBpaPtT3MvcwPSke3N6HRUq5ZDOSFQoRwHAv
L3CmGlsQrkVkecSNwA7Y2X4a9ry+3Vb78IWVFln3OkTO0YcoMlxjrb0wYtnjfWR5
ZKD3PzjY4oJgTOWZJDyOpfyyhePreZYmDnPT1IVGDnvsLJioB/fZOfOriZV70RCB
cPdEFeIeaXRIftJheiOdjQ93ewcW6kyNbZnyMh/LzygXqa3zC5SHBXESADOnbWAQ
tUXUyJOd3Q57QqFqivRe6AZRZvDHmxQPDkBFKjNZkCVPzUmtAtA+/BaWoByf4wAn
5UdtHYzxl4RCRsQegY0TuvVI1GOmW6F0TktudwhhyZeBunrhBfXtRcn8I7w3ZeEu
mF1wNbgv8IRcJiyNsl1ZVzbMTpqATPWQDJKz5C44Fjvn2j44ZYkIZJQd9OZyi2y5
5rfDREPDdD739qq4fjjMDrMxJSjDcTd6y4e7b/P5Kd8Qb0eGHgbnkhC6dojOxQ61
RZFH5/3UPRWz87Q0k2+RiZAwZ/uu5j1U/diXRqONY6u82oD6izhB2lq02AC3zfnx
pUyrsqEHfDUgeelhoyyb7H8jF+hj4HvhmWiXs7cYnHelVzIRa3WdpUwRCvec7Tdx
B9JrG1KUZHAU23fizR4cOsKe7Je/9Vldyi+XSKTcgHLObTEVPg/JvB/SNVULlpyv
1n6/0h5LaykKGxwDyk6LIjAzr8ACxnmaTgDa1vaWCUL8sOV+03qm7yhpiJq6Oy/u
h8gXWAKGU/k+2HTRfttAtwjluDwatTKRXjbLY+oobyLnov9gC5rLGi7Kjp5tn/Ad
SDgrbK8hU630PHQkwnDM13Y8QBLVa58xevuQOqBzztZL3u/CFUbgpv6rJc8MRUYU
CI/J2ffy2mxZ6zala9g/uv6iBoiqT3gA3ett6lkOw5lgPsInlHiAlhWIA0C/yrUC
9IcCD6UDz2rUbpNMH30OreKKA7Mf0ETwPgx5dWT/0w3rgf2DKx50X2yQsIQpUSbA
OI+tY1iGoiYbLVwWNtz/YHcng7axaAe7wPNHCYoWkMwxk5DraRb29BG7811+R1+m
N0dhh1K5r5wDl7H8YQX9QgxGiUfpfi3/VXrR/glkYCttpsfjrgst6ViV1ZkSIDWk
BlHL0eTu75Cf8DG52e8Cr33AFjjWz7MXtUnPMZI9f0EiPUfnFJBj+4GFbM0cUqcx
9doKKC2+XMJKR87DS2wOnfuOs8DzL9cZWzhNWvaTRAv5JnFxG5WfjP29CtbmemOT
oopWWuaVhVFuOhyVK0V/AHhvlKfAN7ob1TUKt6N6cGqWYsZUMhuKjq78YOk161tm
wQGGS9T+MZaAQQxG7PdGJFT89gYHiY0QO5bSI07tr2zHc9vP8x/BMkWZpDgKoaDA
Ja/5caEuegUSPrSdBlD9laQl3EN9cS2KZCdu3jYL/vuWNRyIgHQK+iuyLlBl1aCD
nHU204FwCZmY2h2kcXtOxR5n2VJaJFmbl1Skx+LGRRMRiGoNVNfgl4zn7jAW9d7N
/o53vqElEBvR84Von2kKU4wa0BgkKb3GANM1nHpbrS1KameKYl652ZMegRG+o7zi
mw6N0HAknQm0o2OwqZRNPi39h6vbLpjKoEKXB2JdC8wiIttdgYHYXgpvJWHcyBeD
ynWOy4j8JhXPRaHiF9AVRwRVp6Sz2/CPcZ0uymkld45+xuK+cNCCg4dWfwXE/ink
BEfifEe/x8sv/mMumP1uidNlIPOjScxjS/tyXBk7FD+di/xh9KFruHfcRAVMt8sy
uWXXXdnZGHwJpHdukhcNydtwnYuf9JyNHbRNQ3Rhz/nBuH7u4xu9HANmEN9ygxu8
MGp3ZaB+q76uwTrsbOxRpgAZ+zXZKqnTMbi6Q2vWAZ/ZzJwM+oHkkD94+CMX5zeg
nVY/KLqiG8HjB4p4Dyrj6Ap8oWe8vSdG5H4WhBHla/En7SsLn6ayyRGjFLdxVVTr
FM46Gv1kC1EkmdMpFb5OK06A/HHXSA/TuAXQIyolkuwI1hWRI5M5P1QmPAMZ79XH
woyrQmvY+Lr1vIUd7+gjHRbWoISfBFGPwnJ6RZaVPiy22zkDtSFj/vqeZKo3qglD
2ReQVxQNmG4zjR3x25Qkrr10VkVXGC/MNycB5l0tYSoLotLQR1kk8oPsPyyAu1bU
HetvrobplKvThsDW2umd67M0ZSgfeRqo2njUpDW/8HeIWa8IP6vtmpMgRmrk/ZqK
/ySiS5uhkM94aZFs7uyjuEbL3f8XW53xov09bZMr89u/juOVJTkF7guf4Fy+rUO5
kUTxknPCg08NGWkuf9sE4Wy1NTN1b6iiTkC6MNGYUC8lBvc8jJmwEZu5r9lbT40q
wo56bjRrsr7dDh4KzOn38KcLSRyCZlRsdIS+jw/zFfKP4iQDb5/v8c1BSZA42Yl4
NvKGIkihbeDrvEknoch2aF0zeqFAIUWBGxBjhKHE7yKZ1nwccJxeOlxJP2QJ/1Ne
MEacpPu4iAjfc0PQlINn+WEh0ITZK6LUaGpESdLRq7CHKrmw3D72PIJGq/hmHMuZ
P36LZ2AzmGGXdMDCA3gz0dnwhO7Xqdd3uB+CHrHggX6hkea7iXXg6HEdqmTNjRKq
3Lp5vQ9IMtLVAdryk+OcTaSgyXBPUUxGx5rxpVB6R02sj51kyGxFNkHUZJUgIUNh
bGiS0Z/glCcSWi4urUACVhldyzNk/LkaHVVVoVyfICyleyB0+MkwBZWZIIrhyx27
G76C0+E13UkqZ/hl4w/gCbEuOXmffUxMpkMZfr1QVCNB0voESlTYEn5PL7n0GpQz
RV1QPuccXt9uJU56U7PNlrOji+eKgWpZa+62JRzpxCD+evKxZyjk9cbbwtU89QEt
6EXuLoU6PbULy8j4HjQbZDvRT85KXuTINUJwXcEK8+I5CI/S88d/VgpFo3yWFj+T
VTmkfQpe1p9zkZ/3ltbs9nAFqThEYJIbOMj6lpsvDmTWzfVl7cKuibYbY20BvAxw
+S/zovSvqbTHFBLdeSq4rOyARAE5Ffmd+g5FmznKbSyqvVnrxZRv8L8UHLz9yieT
kXrT2CkT5C0YHWwT5oXgGWLx0qY1DIgTCfFVTOmXlV/yV7BoQq/ySgnNy0Gozkad
j7i7BQX/cHTwtAyehZOcQTjz5374+9u4hwB0qE3MBBUoiY+VSYkE+ppIirXX8W1P
E330Zpfz/UzINi+gS0iGypNwmkepxqaKbPlsG/8xkQW4orYCl+N2AyyraP/LHPlY
iAOfEkGB3gLWxkFcYufOjGybfpH3Vs2GpLklY7TQH5fgM+s0Zv2vDpKwn5bZMfoW
hjc8kfN5yTSMvSlrqzyCn6Pjk7fX+bHYi2p72yddzlaLOGx09fs+V/gGBSvjM6UY
/uW+hDEBbCWZSU69SmBI3ShhGUtqo4VSY4g7Yva5eQ6g8qEKpGzzatSy67rvdscD
3vapUroZlesy9R6p0LRBcSJ00iu+y65TwfwWVRh7803jQg0tqWBCnIXh+JWTJ8of
hvUz0mE/oNUvcYqqHlJr1exZnMNe5Li/2ZlMeCjXGBxbVBe4APJpYSSmqfP0ZA/k
z7zX6C7eDifZ94+iouV0iOfQkkkr0rSES/m4GlyNP4ceAA+dQ7fBziVQ2at0R6ph
WBU5tP39cr2fizSvL8bvZjEUKa3cie9Nk7BkHTdR3Z5z3cdCOHb9soBVvD6mFrh/
JtmElU6CI9yqFkgcM4SgXGajCfmDTK0TG1TZF+2ecNC+DyC9WKjvniO8B8NbrRaQ
na214/raGdWmAK7VywkAF8CZFVdpwubdUyKm7IDo8MX0MzH870zX6LasCNsbhlxG
cfya0kwRwDRzHUQ5Dj25ddJQGvu8oaeOFofbwMXos5XberVlFq2RbjhZtgaf6PAd
/ZVnq6CZdGykkd7Mi4sugREAjFs7qH35dqxmVMRFhGWO2KO6bLIay/fa3I6O5crX
TK5+VMcQZBv+l2yJ+0Qe0ZKhTM4YZ5Dn7LAogEXoxNDL/sWqdFfqxRs5vLT3uMO4
S/vv6FJkcOSTegSHVBMUu+N7SXriZMARdMHVs1cZDwbq+3pIRVJL2Qk2Zqe/yBUm
CzV9qzRtX/z1HvgXb/p9mubwfFjf8pcxMeJo9vAtGsPZba3JdVWfdbWiUuN7xCpj
zg5PzxqnYwcmsyd2HvjvXi4bJjK3c+EMBeeHeH/7SI5o+rLkSPhYSsO9BdOrMN7E
fqKjvdRZxxwj6lmvdKKCxbL4hqV3WRDpQRRYFRXJeLdwQMqMpEu1ZuQQ6SIGWmKT
+yFCnSEJZqz+BDSbUCQEnqAFJpMN6xqs3IJ6SlhIbKVz2DXUyxgS8h7RtTCyozKS
xjgBKQS/wCrFNStUBTsATvlcWRzKvgP+iD0fbe0CNGvNRwR/zN6/4AfDGmkSicL2
XoTBeBwLTeYMhx4NC8/sTrDoQa0iZFU91fLnpf84Djjv0wZq1o9cUr6iDQ5Pc7mV
QvPJDnuy/BotOPce56vbi19lFSuMYun+W3jAMSVV1+REVxyKrWkTKwwqSZaANWa/
Om2+/XGqJMxYdcXO3cp7ZG8ydDNXkpUGJqGopITL2hiLFENMzcAus1xT4d0Et+AQ
aRgOvKQBxnLfEGoV8GfxPK9rrEkapYUx2WWqYQ4c06q6yTjRIgqjKlWk0r36j942
kcI+l0NZ9mNyQhWawmVYB9eJplyi1zoj9ir5MsSp3ENrwuCsPoFLKX01aZdvizg7
Bloi1JbJ68TzbulNNWjYkUj4v65hiGm3nyF5TOGDVSFkVgDYTmxH5/wxAtlWvNgE
bvHYApDaXRz5Zx8etONbp2M/9ErOqK2QdoVPJIcEGR0mm1y5xDQrg1O/AQPuNhnS
K+IC0V0lYTVe4t71823v0lhpnOPOKHT89QQeK6fReZCKjoYak+HyUKa+Vi7osX0J
bZtp18IIyqTYA4EMAIT6Ge6skoUu6DwtfAckDM8FILTHaPpOV3I655sckAzlYdjb
6BBHBOEJFd/BDBbdERdntGLPoxHbK/KQB2DYPRZ9Fgle87+d3+1CzFRamRW0Pl0O
CbRYSBHrHj0lVNm6styldqgRTodJ0w0p6rwGCuI1XgDOJXVE4VIqtKRHdkZSUrGZ
7OyoRJhKRVH8l7unkhujXjZTDk3XYMIho5n+7j3/7ZS4q/gpKMyAQQeZeKIs8RTS
fHDUTDyZYeXgNKtKV2LKtxINp0BBgA3/konS4ynsN7CSn0A9iclXBXdXPYeXqVBz
ba0YT/CGJt3Z0DLdbcV+mXMK8hnSvqhLCknw22fw/6Jx9PjLol9xotPwVXr3Rpqh
8e9msW3ppDJ8kGKoX+BHTQhjFTP051DuJPGKsMjxtEq1u9R28oEKn4shbiEus62h
U3zGIUW9GQ0F6mcaY3VLQGuHS1ptu0eWnAaGDQpyfCoqU/0iKSCQ16i+nteOtBjm
A4qUYZ3Fn+KBKaDrfASGwLsW+LNlFbckJbKBN59/ZYHzh8BUgNX8bDfGR+xftvVn
wOuv8/BTCFFcCvar4vs2ZGsSSiwVRVsn9rsJhoOskz9oUAhjunYiyI1r+54bEFHk
VHGb6vl6dqjEUECKOBCDxOZMx5tK3RjDa0RO2JCFSlh3WQmrkxbRqw/BG56E/HPN
3mtz4NsYozSO0ia3KGdtPtILqn7PNLetWeok4aq2awxMh6ZBOrTNcPO4iZbK79jN
k7ZTYUy99o868fq19AYffbAoJ1D7G+g/9u0r5tCEVy4Spkg0NIpzWfrWx7uVmPnE
mQ9KE8m5PHlN7OCT2abiMYxk7u1u9BakaGO8B5qWkugQ9pPea7ECZsJ4cMKnhrq2
L0eQSJsBl/7wz5p/ibB1SQQva6GwXUfqSjDdtQNxy/pO0D+7RZDyIeXLeage3WZY
sUFWJGMCJuHwqHjL9aMtY1PSqDPaCYjsJUSiP6JnlvaNrXO4Eud5LnlTkTJa8Tv9
zyHmxXHCQbp7dQgeXeLX5WsPv6VL07YALesZj8kkWMaaq7U3vHjzvNJ2y/Q4hYdp
FvSZkcbOjG+DH3vfVrC7Z/ldEUaPj+jP0ppKZG9JNpK5kCttbOzhHGhPc0WG+bGe
qjUHNv5ylOejL45RnuCVaarJ176fQa4U9wIjKacfq2WqxZYLTWDvCz76N6QPbN8h
mkpgCcO4HX7pu8fYLEqyPFdVBvjMjUWdLX5NCeKb08r1IbJ+VsnZ36M11E7igaMw
gBQLhCvHN0enQfbG/Cdg1ZIV1pWlLBzun3WjTPvhMt/TDPYvcIu/BnJ4gUcSQUk8
w/pGrF8bahIARvb3eMUYkb9D0crKWak3DzTeenWrMZbxl7TKy+VPTi3MK+YDKll7
VAInzAM86MtcJEYmfLhwpW4jc5NyOfA5ZshCbCiEeizKsqEU8xlg9ivOk2piXapM
ziC+a0TwhjyklkvWYB+gMv+IFyFap8qAmF0gbmyLpQgr/HbsWSMDTNZ2HEl7HBDX
HBJtYtOETxKnkfaSqfWjQ5HUNom0KEcseUVgzMJ9mbiDUvcLnBeZ2aStyQzGN7rR
Y5PfT9T1/WMRwtFB7u9Fm2Q4RjPc9sfpTPIo96VCm7oAKGjV1mncsOmVzwjImF7K
JN7c5roCv+PcE6MdF7rayXe6M7Qe1FSTL8JZ5NLkGIMQz3bfrwGL9pQK8HyQ+beD
VRlnjx7AQahqGnMDiC9QVVKXBkePsHLLsyL4qiC1Ktam9UXw9mdKM56Gs+A7zgfN
0QvTuYsj5qqWaqRl44DRIjqmUurjbxJc4YoIhWWFNmhgihEmmgVl9WtzJiJiGBZR
YvlACN5KW8jOh1Ag7JO3BhRK9/I/P4/dK9gAfTsmaCuwYVoDwDfXQh2U7T+w049u
zzz+Gx0lozR4RD7iUzkVkwId3uckrvy5FiZTOPe9XYO8tXz9ftJMvywUq1CElRxR
atj7pQasU4lueg4gxMO0YXML9LY9lpyRIQSEJFruDZaFdrkHaoMAfsly23rOZ0Ex
x73ezjOWqEo8prH+NkNFPY2cceTgWQNtvHm+3PDCgg91Ctkv1B7U0Lm8L1QFDG1a
ZxsIHvTN03FD4T/tPj1asko6oRZqbOhlF1JcWnKn+BblIvfeb+ZSXQ30YhSmNGAd
4vNLlg+tJkJ3prMeh50MvQ4dV0xz9Pp7aNfJ//eHG0I4qvUhvVjuHzZEVIAiEMoB
dlWo1ZqzGTHDDOY7PP6L5DuihrPgPz7mGqllcTQXPFJ/gMb00apQdmxfl5U/NSr5
kg9/qZ60YtOsJq7SFr3YYNIQffcjkWd7RfIyV32wGUKebTo368EpuCUU6TjVfkkv
ozf2Yz45+WgwpmsjlKiP6Isvod9HrKZDziYRBbt+dQqz75dlP1/+GqQUjNh+VcHC
XJ9Ndim9MgU88ysKhX+HdH/4lkuk6JMbKngoXK3TNkwD/6JO/f8GnY8w3qKpmQDp
D4T2YHjUq2rC5goTQbw1klvE4RrX/D5xGwHXhzXnmf3woYBQieTQ5z86Tu6ZfKtH
YkXvAC33FVboXzwIaBdLo6pK/Rwfxa8hgBB1C4nAG/x8GG1dVhgzZtSYP/IOU9IF
PZGLMXFvzhvTuS69sNCO+qzkp8kf7tOVguH4wMxwiAoCDllMvX8VjUp3Z+/dAvFN
ZHhC7FhJD+tt/GGy18p1EkDdr3zyksdIsGeSSyvUEbMPF/wN1YSZCoT0JffQ/dSm
nHpM1UM/ICZOVil2s4oYNS1Tg8IQ00pYy0/XWEF10SKwgPqf2Dp+MzDdyKx76vzy
oHpCNA/AEBt5BFOdOBwLd1o7gXVSZ6yUHBlzHrtmtc8339zJOSEef+QCqA+KSKCN
ebL5nFDLP0Ye3XhxWusSnzoiK4UcphrN7aeKuLT5M/3BlzG3fGWOW9GmG7OTA5n8
HggPYvUL51bhM78xphEaZNFQ0uyPPqGRzsoHR1m5c7z47yqzNmUGTSQmqT5/jRcq
Ymlc10RyU57bs7FlhBjKGQEhKUXk5tPy7/Z8X7T7Iq8GOxz0O4uhvG5cYhQddC+e
sJhTBy9Rc+f8t/MrbzoQLTWV5TF1o8rFX7G1rFMiaWujDBevRIzYqzMAJS0w47cq
d5edNBE67BX9MOCSiYB2+JVxtAVp5VGJxKSrmZY76/KwguembTcvTC09XypVnn9i
8EpSjuaSXMCVj3Pm9cPw8gQai+7gm5V311LJcT/4v8vKYpZjKxIR8M5VjwuFuMU9
F5CkgB/xNqJ+YJ8nHCUT1KPBdMfCNKycei2ICPBPSoGC/1NPt/73K/NP34WH3o2U
cI6PhlMM4vFQxNjIQCTMEEOKsHPiozD6BJmaZoPz0q2R98BzTJPB33pDDUkZEGea
My++MtmF5JVsU/z4LFHqgMcIPbwkgGeSnlPOI4+kaVYp4xOMFvfS5gUpCHIbJzzo
cW/qxjKiMLw3SyUVXyuft7aLEEFuHoxSi/KgUM3VUhrReFEwSMWjeX+e5unmsM3q
dH8Rf2l/Wx7cBgD9QGIkffV9acDy7vBL3Yvcd4UVFlx0I9yghHoyvKHlmdKePplT
Aw+Pt0ft4LryUtrhLq+OxlgLW6W7c9wV+Cigm/9Q7hJF72wsXZjnu71KdmU/yvqn
NbGn3azVgF5PxD4Qai32BFukTRpOMQJkqIu86/7XV+XJ/YtDCFhmgqDnn97rXIbD
1JkZ6lRrzgWYWt6V3TSno8SL26BUimb384O1V28PBiCic5T/UO8meZ8hvQ9ORjWh
AqLJwNuw9rn5EuqJRMMha8z6yDbcUW6uWCS9I4IdY0TeuF4ECLGH2vH1ITyNuujX
mO/jDHR2kGpK9RsTdNQ3XMpFOFewhOM9dZ7CILfehPZi1qFs0AmXT7OFR3NoU4L7
uyZ+rxAbTXtAZXhA+3Yu0N5bHkp0oW+qZfTOE640JWzE0xhpwMMzSSp0zhxwTzEa
KmQNzKvYCI5MjA5KGVc3W/BEA9atCA8ZieuqzyTuD6y5MzUwZQf7AZn2RVWUd7WJ
1RX4ZcpKg/ElYx2/E5gy3orhuIiLqHGvTaz3DJfS+oqtpSKsyQTm0YQ6EEYYu3wS
XNPUTRp0bN4qreTxZqpF10Ebvq1mvBJi1/XJxd5EMHz5TOSeVKWEpxaGn5vaDfB+
keR0RLU7PV2/ANVeVcnlcvEjNg6scMdrWq0mt38ZAZshCk8fWThAy0nTT3OPo2qM
CfivbRrAqRHFYyG5amZsemeZPsqD8C24g+pRfAHyeRRC41L0OYz35g3b8t7n3IOy
DU0WBnbIQz62yr7mn4Hp863l/njPlQ6QnV94+EwCs1M9PZy2mPuLCi97/2WJ5wW3
RI2hEvfCR/N9wFwmhqPSGqntlg4mrKKfmA0Ub3jLgC/8vbfhzOXzKrPwbOAQQ+QF
8eb46/ofcqSw687SkBtGSezkaRF7eVDjZKu+ydvds1n/12YPPfVCWZAGUuklrVLf
3BIy/ewEEAXfmHkhpcCNJxavlhAWn4L+BvvtAc9fN24Z9CVkLxE64hschUFo3vJE
OU4NrDMu/HHW/izuDmDfE8NlOIxonO7c8uFZYvQCmXqVPZCUN3AmesjXqQYar8qy
gFaOgVWsMFyDTzEMOvUXWHmxuS6EGr/d8AshHIw37reGhPXjNgT/xeG6Yder0GBF
owX0cavgug3G34CnDx2ASC4yQkEFPmqtOkK2OOW/4y+dgMohSGy5UJSI0eN9ztf4
ctoyY6Iaand+7NRTBCwzbiBH01/vcebWA4diO8+DaETg0CPC+oLJ4UyQevuHGhHk
TRjZCckSV0qas5iy7HSHesA16TWFq2tHeiWmPTmlOvYDXVxzggBJxx89TAV7byTx
CwSBm4cC+QNCyZOvIWSTIsW7tOau/jZ9BLVOJEp/rIE++bBohciJ3TqZthSdWUPE
y7Hw0j4dl9uxnxv+jwvbqrb+u2AbKrcET1OGyoLDkZXY0sqgD7Kbxu0YeDx/OWrq
uriq4fM8G7DVPVjGc/VflgfUL4aBILWDCekIWlf2TLzCV068OYpWZDuUKN+dXK0M
UitGJVlhI1rP6Dperup520AhzBdku/uumU3q803EfjODqVrGUHo3VDCFMOGLsEs/
Ki0X+iKtZziCsbjW/F2AfKu2bBVlmAdf6wCV1ljr4MFvNF+X/++IbwBJqAEgmukP
Samx08gQTTO/Bn9NlpqRCrL+itSdun3qOP6BOp9XUV9FkG+GT0PSw+ixiG7EAkjf
YOkBx4XW5Fn6OOAlWgWPhJ+wbMTmRZMzZbStmqqTDl/F6Yh7WvSSkLNabedxOCGo
11bY3m4OoLgn51OqIjZ5wXfVrOJksKzIayvOMGvxlwG4a4la8qPdtK+nP66WG6EN
a5DmFjdVzPYBciWcdicks4QaI32kpDNNQyjWiB+SL4JIGvQLozTtaH8bSeSWVCny
GNwUv3ENIRIBe9v8KKME8N2rCHTx9sqLuPzFKME7GeiSZift60pmt3jHrxgLKBP/
025vLPZRA6WJCfCh4dFMXlwK+63Ziey88oJHJGH35XKFjFKB6BnM8Hp9Ix7Ph2jN
BpjTytX2pnGTaYbhvNGn2A0t9nV4hi77lukDkH7/ke1IFdz1UhSAx0pN0C9ZOsJf
ur2h8pCLHxG35IDyq3sRjZ4MRlKPCNVTV8R56ffAo/7k6YU5die6oGT/FjrFaNr+
0I76gr0V2ZlPXDkDXXgEvU8vF+kbJw2HaYWWGcbzAv/gYJqCgY+Te3iQrXs6EtRg
HqEAt1s7bscEbH3LVPpZ1jnONLlpUmwhW9uvAgFcOoyfbJliXZa6GkwOH4ENX2xv
XpU5i2DLaRHjzqihv+j7hCBCbBRPsrDNP08csTFxEX490Mar3qb0BRM4XtW/L7FD
vDARtH/e9c555xOAb5KFivSk8kO+jS+kL25R9uzAZtQGP4+JSGe6173koBv5ukBW
vADNTq+YJAX4IyG5erCPuS10pxWilCcOA5Ss38FhJdUpQ2d4wPUDzOQvCbq+l9Pb
pBkeS2Rdxl5N/pAYmoHTYJcfOuG+gRuy12qP8CcnuTQcmLU9oqdoccaQoCOLmLfS
xNeRmA2aDcVhPW1enYLwkZ3yKBNU+c3VhMjbQs2EoXhqjkoXktJciVF48SUbkr+f
P/fVBMIXSTp/P6OpCufQPyUQWcPXY+5zDTlvEgAM0FVvanspmoho1hgFvb/chtvj
45x+kEaCEUtosYHQEeSAU3HSwPSAXVIUYyn1b9mP9HH7t6tZeKJW1dfT0RIJO7DS
QwZiWLY0hQkOwQ7J+/eQGy9X4JjhLbGLnv2iA9oeIWD03eejU8wKfMCsE2NvWpJ4
IjS+Msd8GSri40vrQ38SW2YqE3JdOcmilhH0lNo0/rnW+SmhlK0s0wPpxOSJEK+m
3kyiIDLsq4oSfwZKZGGWk38qQg6or+0jxZ65s98lauQ6p1KREdNqKblWQiaMUiZs
YkuXhZKo0gyYFlsTptZPb4LN775lBgd9a5cACnVa5voBdwYM+CIGbVnCZlTLVk0k
uZm7mC7+l8Fd9qGe65tDppqUIO12iZU0Tv9pY83+H6t/V63Y9ObHFniRcurD74WR
t2fZjcM+wh3CbsIbSMTHyRQrpG31KQctDm7CZFbP9tI7lXrXA7v88LBisqYFeevV
+wMJV4xylhqeWxIOsnX0j/aec+0majUvYohsJLh0qYWZI6HlqTjejfI+AtuSXJf3
k/RoDW2Kw9qJf7O+T9TBKV0wtdDjO6T7ewODjccsgwfTE27Tf9bZTNUYNw25shIM
O05s96zJtX59pZW6NanYQ4roQe8NS6zGv7aadyx/IcUaTgDLOjw0MrbJya9HoSWu
me6lCjfWMYFD24HW3ZGQLjeFNSnouhCAcEKX4M9Zo3wnBRemM1T+C3YjAQhVIl8o
mSstHtXil1lsWrKygmO6f/HobU1vDI/jOdKwDf1VLu2+klT5ZRvoKOKrN/EeMoe5
jOZSmipxDs0xWm7RYfJTMSyv/QVcxuyzNFEE6sEySAC1mO8fhzgcQgXyFKZNB0yj
QeFsGdDGVSzE6/QZj4en1YNAJyXGS4I3pamgHR58qnpbf6fFx7eF9KHQ1LMMJzpX
4hb8Ds1HjCJetBtzwEj/0AI9VqmkRLEJFaGAvcmw53r+eBrLXOSsAqUxmSYulLjW
lBWjEK/LgOZOHxg6C1ceS1iexaFc3/cx1TSe4Q6WUNFhQ01XGpre7D5MRUyLXPbL
Bg2LJXhwash8Pzl+Cl8p0uuR8IB8ZO10QRpWACUsYBtWptxTcgK3p9cWAi0Uatbz
bK1xLs5yfN2HSIoPlIS5obHo+RgVopDutQAT4ojWqiHFstyIJXAgb4UD1G3kYJXv
W82mPFocGBZ/2jYHBodh1gfHkNnH/CrXwzaPrfF0JNGRF404LRmCy9Z0SKJ/JU4/
qZvJU3/zs1WB5sd4N8jikuIBz3mxsLNRCpW2WjjxyzFzI8ggk9Td5HQNEG6GMdk1
BYBDLKSXEfji9wtHolddSKU02YFqu/8e4bX+v0oa3fFJc3Uu4c8ehW8pLfNrz8A5
FDgAJde/vDWeZenA2KbRXlil0QQcH2D0cnG/eIbV1I8jJJXmMGkNUPwVMPVk+RFI
RmZyGZWQRCUT0hkUeHPXwNt1ZMNnrnMTuQ0r+MzgrnDWXjlbEGpb/ygxsoMyrXTA
9uKW0gClqTg9TyjLS5hhv8W7ldRxFNBm43vKOfCqoqjNB61C+hOzaiJ7hbNtLy+O
EYEI/Cbpq+DXAPxknv7SLCAaX/Y5dYqaJGmsqQ7e1d7cwyEES5fYmkCTpLnj16Jt
GMjwmxTDMTDXw9WQPkC2B9V3C8gn4VO7GT6HQEuwKkNOdhkM/feCdYa1IRHj7XwN
9A/M/rOFH3wI1cRSWq9nmz2+yHBjHkxY58AYM78UtVs7COn4N7ikYFI90aMXsnEk
vkmVIyTYEZE1UnvDqGAZU1Q7ssxxJyild7aTHpN9c1Utb7/gLOK0DqdAaRmWHomy
+GPPa9QpXllBemQadvaMm+O+kZ0lo87J4e2vDn3nnztVsytM46kd3RADQrQ4b51v
y3NsnVohtu9V7Y1mI+HSkUEGlhpZGPvAJhft8bENakCcH1QQ34qOApKcEJQO2EiZ
dkJQeugTCTu6gHAZFd7mLJ8Mfi+P7cXFQQAmoibgr3/2Dkq+PE/DpaH0YzKXgMXI
7Ez+6cPl0ehydUMKZ+nzWwhTvHt1/rIvIWwa1hz3athyXxH2k2P4lNRjbRaOXWHX
/WU74GShbAZmhASSrS/7trr8KhsoRdWoNTq4ZhUDm7XXRhU9WpWbTr40OSuyLCI0
a+FvI/8PxNIiDoVlwTEw6Na4Wnnkb5/dH7ojtWuH1oZbrW/bJO/9vh/a9Awwa+PL
n6G1ujJ4MQzD/hlfTkxjJ5v6aYktzuXe9PSSeVBHLUbxbQE2qwKs58i+uDIDMpH4
6mfaW3E8Zy63hp8eEAB21Lc49M3HlwnbQTHt9BlBFkSMWSpV72GheOpYRFgHz55P
0WzNHIDEyAJuxRqk9iT1Yl126BGztVEJfS/NeR2ki2Ukvfh1EB0AnMzB4SzFwMOt
1wp0PJGD1m6GH26JuKzDM5c1sghwm6W4tudKrQLfqqG44+e4nXVhIXidii7B4Atl
ibE2uQ8iLb4Fp/Ol/73fjpgBRkflAqi8a2xPTcH47nxFEWmiHWCZwDoH+j0p2MR9
RCi2h8dbgsTk7btwKmT5qN/JAixcKvstfNFs9MvY0Qiejh5zaRFqvCCTEOVsbfyP
Nn+H50cTxLW5D+zRkcGuPH1QrpoE9taWXifI7BX1aWgUs63jp3ihs1KefBQbvakk
/jgVRisqdlrO2whJbd60gyOXsDNBXLAp4PXtqkLjzD/ez8IolW9OB8zqoaL1qXw0
Dz5KTiuGOQrsKaRSehbLVmJO988tq4i3iddzvtS33wJjsjiwTJbCdVkm1fKtSt1N
ZDf0wSo78ymiQyY9VvZMqiMvLRAax54mO7Dzf5KNTcG1t0z5DYDW7lK40SW2mSQ6
MoMFdcVC78DQ4oqPnmgW4f3qpPIZMn35TddqTSJWclFJ3Jty7hiRZdPYSo8n4TyI
qR1iU5xzB8WljeDzAWWwrpBizqpACkbkNXuWVw8Rd3j8z98fdSues+lhBDfd1sSj
mXw79NW9YBV5qtmHffsYEol8Cyknc5CwElCXBqWla0pyzlQd2EkCOHwgP7TE/TZJ
w9s9K8KK633MrJaZpFwyBe/mbCaOFVUz+ZJxuemV/uhmstDDJraGXUcvnp2rcOmz
NtmGFfB5yKdYBQbA18003/6HPJoIzuI5SS3Hc/yP+IrgY3t8QRpKCrI+hs/GLd7X
OtO8jIXOe6MXaep9p9VII0azvz/UpjofXf4wK5RdnNsJJ0vxM/R/P9WvYuTYaStc
cKJnmXmWv3G94XA6ShM9VA3YAxtfvUCqJrRy/N0zj4+1tj7rNn3o4auLjsQE8+qN
ZQC5zFnINrDFbzOx5SPrNfR3C3vylbmPUIRDzhMWzHJfyYcmyjVGSxFkp2jUerPs
M6GVPBOWOYaJc8gftNsF2IuLaexNeh8V7nZE8cBAxJlzZG62IYM6J2boWoPsmwEh
H9kaMM6Y8DusQD95HHyENNitvmT4h5PlD3sEAlG4Qxogn1o68FS5I0m2KZcF6FTV
JEfaTH49yXg12MR6Pvj0RxPiHTs1lcjOfz+DeGWlFeRWFbZmhlIhj6YB/NbYWq9P
U0pblDj2sgLNRwCRxPJjgj3axzJxkg1KG53DKiEIkelwb9ks8hexCTrDtu7MKbgi
Jc9fctRmeXW+WzN8O5T2c5rWQZ6siwB87NYxHsctlYhS5+25jf8ofhBu315mNVHQ
ojmN+j3V/4OqfuNaA0+0ugXsdibuvu/yoDiLh7/ZkAjbOrKwS5VEcuOZFp85zOui
myPNGi6LR6jb2ko/NtkhqKak+3w+7bkzqwkCTeOCENE+A4IlhX95T+4v9epzwZaP
gbGIE1BL1Di0m2+f8NAhLfyXwxDgXSEyDClH5n2r7cGsbx8LzMHZUVhIDBEzDKvw
G28/b0ssnPr+OdZFk6lRYb/CvoMgIMhDZicW1S9JajXsNPwObB/aBZoglkKpaJxL
WwdpmDQkAwX7yWbrdOoDDt+vxfVJg5HUbypjRqtAvJQ93Qzw+cygKLJ0ns31Vsku
BRQ3d5hrAmOKfUTDjk2OlSmmeVv+OG/Itxb09rR0yIBhj4QHzFs+i6sAnXqstsqi
zBKL08c0HBoFteRQyGwK1F0r2jqYXoXvC923xDrplPr2CcT7WykCI3LQKuhB/kp4
KjwARTozVNGNuWKt7dFBYU8L6IYftSZyz0Av7mLFYsAqcL1os2XHxdL04HNc6Bb+
hGGabhiVtzJsX8s/fVHWoS64n3VXAFdvs0lQDGyNZWyuC2mXBoSwzN6EDGrfpY6S
YlUEP3TRGSfz/jPmkrK+u/voMmsdDXlgLUhvNnGa4ugTHHw5ckl+hNECmxr27nG6
TCpRrKlTjXsq29GHVwl1zhkDDsCX4VuKe+4eyqKqRGVPMUmOgEED02CL5BBKOPkJ
XA+Q+9H6y9ZHj98GIvTOXhpYcQtvr+FXjH9gm1PQuEK7T9PvMIacBYd6YXuGYXvn
PWz53K8yhfhF7rWeR0c17iMSOaV9zQ6LcL/SgJlF2qHHxbj22iMVf6GGoZlVC+Ln
aIvb2N9yugVi/hszDLLWl6y4yoOFQdD4N9pYJmpazgWs+27M02BpU5Hh/8J5oESZ
WE3zX8tm5vE+lwDNxUbkheGQe0z1ASCqrILdnLWDBTHN7dMQ3m/+H0I80BRrzQdO
DeBhUJegmmUN08+aKAWvme0a4m7nLNJYNqjqsE4750RDra90xVuVM0Ih7Cy39dSZ
m2bz0uFDITTGK8LNhxN7PSOM0yLV2hgJO7SUY5lezs5PKqswVxXUk00yAfUDBBqm
JJc3FtxwtnkAEgUWoea5pFOnCQ8/wFC+VwORNQ0HCzsiyzH4NNJ68dUcaVFy2MGe
YVzUf4IltEiY+19e9mrLLn7dkDqWNd9Y06tDKOZT+3fvhFUC3AN5LYzTMb1j2NbM
2Zy5ISRvaLLfafH+Mke0pjB2AJRMF3KI8kCQiKOn++npUu07xL7+kclza+IJ7OlO
hBW9qYi3FJPrL+adf0jmU6aXT7Ychgy97XG5/eLrDl+ot2g4746SSvigB1xnplOD
+NfyB2bngP9S9higL1FJc8ZV7Jy+kCprOp2W4b+HrJPwJkGU0yf2h4H2//1pynHE
zWeFd0FpBlbeYb6fcFpCzMWDGu7mAnlg9bOFVJbZNN5c/js0Fw+zRz2G6coqE+Gb
F6/Y3XcyQ7cjM5EbDZEGxCTqx8xk/bNer2yPIzWYTZzplM1dxfjcjX5C82BPSE+8
fLA6QPXviiBJZm2AuK0BngUg4KY1qG9Svo1rjsq/ndDtubIa72OyjjXR4KfDdktm
6BKd7qw1AJISnLyhIJSq5J2BGLHV6wCTzovGqEa0a+9CD92NDr2h9NM6EYGLRP9L
PPt+7ptEFeT/E2zrldlPn6KLcEjtORNdLLRvjT5waWDpkjn+q09hDeEs8HulOrUi
sC40REc6DVgHXFGSIF2e28hz8jWf4YBLYQYbxCTeQQ+26Ptm2D9FJZQh7y6gyEsG
i8qoXQUvyNkkN5jatnRGCvT6b5msQMWs0mq3RRClA6+ESFT4L8xrw1hx4LBkclrm
e7IIpzcTPMWnRUxrzg5d/KExih33kkyks2BBS5MX8dsoxqWD+sWkaWMjEN6W8PZk
ZHZD60dY/4/BYnO5JNffJgZc+E0494gww4MQMcq2ZML0j1Fx5l3VatYGkQBKfmXR
xa0Wl0C43wAxQFoI3qmhdWnPaoDcaxq3DfWPacvnQaS2SjM2B35oS9LJ0NhOS0R0
teAxLZqWJHajW5bwDw/8k6abH8MiWbUz+oPJhTZuKZsDBxYp6VnBM3DPHARGnzvj
xc+Aa8fvVTdMdnBlUsx6vIoSY1n++lRXcahhJcWS37wbqF9NMhJiqPhmU5PhlXVt
EOqZeibDrgf3TuuPPrz54pRc/ex1jMmYaE+2gqS/Q5ksjbgxE1alFUDHqZ3tijVJ
wboQf9P8OgK4PCS0D5i7Qktz238z6U9kl5hBOQx0xYb6EOV6/BQOi/UHAv8s/jjc
9o52Q+whxgpgGjYDqIebq/QqqiUY57Mdvf9nJIymztFDWKRdp5OMntMt78TQ6FW8
KAW7gW0mbg9PGNKtOUrzLp6q5eIqGuyXMW7AajxwVyvw5s03ltiGRIkv3OJZy5dw
9WtsOvomQVapM8mE6i5Z5Ag/AjgQPMzrRoevKmHCnzkp4SgsZE9EnvwXjggBUFTz
kEUxDyhBkSXDRvwjII7QFQcGLKNt1OaouAnS0bpBSiXh+knfuejsO0uOnPlOoGA/
wbqO9UDvQeCuQudqBXGEQ5X2LjUJdWdPksubEO/DltTQA+2vEhMdlbMNFwNDC5tU
1S+LZxeEmEc2mozg3EzD5qwJdAgGDjuyD31v71RJof/rrNpcMMdWFdoCbxDM4DoD
HJn5WksYJNwa+KyQQ1I+x2wNVXuHrP3yzdQLQtnLDcbV4T3rZbHTlmu+hV9Mn17U
it0NcOwIIVhK2SkBimz7i4tlpSzvO+Zv/x+3sJfU3SdP2N9eVKREofN/E+61o1gy
6Pq0TByorodVH/QNCDIJ7qgYXCrRQ7YvLu72V2UeNgg2zuU6WzdBridsiOO5svIm
KgFAvzHCn0Ff5rpX+Sl7S+thRulfZRkC0gYnjmADkxwxco9Zbz7AcwDZFoI4z/zx
WHOltElQSDd0sl3diWe3SmWcQkTcF7DwNdja3X5upMKtM1Qhb9R9LmS+ko5HDnLi
wX7RTvCifKjQqgS0NR1Jp/Su0BsrTZ1JwFfQN9Mvwar5K68NncDAbjU5D9+yV+Fa
zb6ST/S0bOIhkCQTcn4qiJRTRJB863tbuJI8w5BtkXbpwXnc5k/DHq9vGBKr02Lm
xdNQv4Xq0XbQ2TpVVjjcNma4U497DRhWO9QP2rxRJtfdVkdL2R+L+oUwQ1c8UYUl
jt47V1ufZsKCri/T6yFdgNQnh8iu6yPwsqc5SzAF/McyaB66OJ6T4s1x8pwEOXeM
rGQUSMV8Skoj6E/IlahBZ0atOcTVVRxGwfhak7Uek2r/aaUTAdCTK7Ci3WDLn53m
00sDhO+KjAJWtmfvX8mm8Vt8gjV++kFsT4notB53PxMRAvaYiUDqyXU1HOKnsQ4A
OUrzB8T9iltvD8fgSBu6CP9/9C1IBjgwLXGv94Ew424TMSu8Ksl2fpwaQFkR694Q
bGQFSfBHYbL8M3EzQlkMghQAC4bnnJhz/ClIZLnZ63Ryh4XOt1F6lTtWZ/x0OfYP
hLtuNcRwG7zwACXU6gPvZUz1KCMGdB15iWW8UBn1XJM8fJKP6+kQ0p/31uTgUAXE
aLiu918OgCmkfRrmbhCHUfW5TS+vDAtx3ZBbTX5aJKvR9sRvZUxwAT/wDspv3U29
SW8OQ/WKiBMGpWCeoRD2GQ13Cv6o7ld5BwCMTlX4d2SCZFs9LyPLmV3CErN7aUWx
0Ei2yp1NkJXVxg9s1tEGe+eYRWk1ADbMwKZDb5Iok5dEbneGQKfT/yNGwdqd7109
OdXyE33xzyTdcMl+Kt30Vxu/RNItm8ScLPkt/98LPUg+XKAOoCRGiFG3G05UM46W
+pUr44JRyFYOL22D1XFD4hsfvswVziW4TCttipJXHvyPYxgUg+3ZZbBcXGIEpWbi
jjuYKHS1k74G1avwnqOf3hFTsFoQR7y1AxhQwGmycqfEfNifCI54jQksoSeJVf0C
gUU8n9Pg2TxHTxImI3btyd375SH7sI4pRLKn/b8gFhf45cKDUvrIuMDeXj888tSk
UBaUVeOG5Y6PWcVJAtrriVxF/Y1MAAwoyrxOnH4hOG34L8f51XBAbqTT3AXdAaF6
3QHhRXJr2mrmo6MoygjqbG2TtekGbVdmGsnk35+kbS4kdYGBZ1Hk9ElMAahpN+li
3yGoGY4Zhag7QInhCaOsGuE30tjFb9JrPoCRqTR+F4zlVOxzEqneWwuHsB9yIyUQ
34gVy0YIdGQP4gq+xw15VYjLIubFw3gkTpbKa8tfPXbGNMSvw/XkTsXdTw8qjpuY
k6yASaeQl4rckKaSwTEI9xjMi+nke0ih3etD2ZbJ+LSwaDBBYhNTosW2wvDZLYum
q26uxuJa8GeX1t+0H86aqg8+qT5fq7YevPdeSxAFLcPmUDPGx0pP5Cd/+DibiLC7
2GoEh0jC1pZcaNYn9Ybr5REHRUKjMq3/AFnbNuY7xVMFO57qzXZb+o5Q2E1qudfw
cO6fczYgfDZoMmE/pAs4Xo10R5R1WBRPWgRaloIeITPeMclW67Aq1QG1R9CZXB+t
WVkFXJUS7JfAHri2kqaH8wXJoBEsjOBDBk7/R0FWIVDntsf2FJw8CtWP8AfXNhAu
/0InXvlSC+MfT0FHBV6QwP9NdL8P2gW20R6jFl+qAJklBMMcKiKk+FQQj/l8qYPh
KaCzT5qq8pdWU8qK33DXOSpinubGuVVgtq/SqKLPwwyDZVBNRrhbI6vCbqUyK/QB
Z+DTnVjOL5tjNCaeseCnQDdfjyQr73fK7NRy94CBLdM204s635nZa037zd+LfB0e
vp8xxQzYUiyk1WWST9yUyLZUAuWPKaz8CKHjsS5fUqG3UL0LPCBBYCdjZUfem/2G
R6uTBGl9Mz9/lG0EJYPuz3eiOrBMaiFT47FLDyGYk3hIx5mYF0OMEN349NlKdsCL
K85RsPcMMhD2gyffp+Xp9u1HJggFJvXHm8r7ngg89gknMtjlb4+mkaZXbNvHLpfl
+BACaM6ewgmm1R1KupRcq5Fsi35CpMtJTLmmXqteV6ejlgLbLXA1YmAWuhllLwj6
hlJXMgdgefxxDt6MYE2nix5SAO8i1/PVm9rI+axQXAX9BmTOdc/6SkoxgNaLyST+
CDTqGkrIVHzi4mk4aDKucLlE4ludXxHYLQbm53EJQlFHubL6bqussSYzY7T2tuUn
a0CmzzWtdNA8VHO3Zj8BjGnK6lqu6fxIK2PA98+g06zYa9ov1T5wK3BQKNWGl4BC
qF8Nxf3nyePFvfGnHomSlwBCznlcO6el2cBXRMINzH7w0sWbdPKBYs6y1qw8rNjJ
7MtCsauMJ+jlqb5WTQSmKhiZM+warTPfiQuOsCAIa+ehgtlGfxQDR5pyo+5HTaqp
qwwYdW1ezoLB/eKGY9HAw3z3kVujfjZvTo24DkIxTQT9ZlWEzkkouwN0nCg41qAC
GCzpzhdymVGQG+/4fJo8MjPkdV67gPU6VGDxTSnalEfZIA0oIKRdMvJAa32Dvkis
ewcNHwDrwMRh4RPjPtRwJtDWm5oRO0MVkLpPRq6UvnXC5Mz/nai/5DMJqwD08cTT
OUuC/811dxNjLpeyLgiYTgeeoxniQSMgsfpzryxhhGbddRk43sxWXkwOnfbYYiw4
Jii8V9wSdwpnrIbS0fFZCgfSu1E+nDazW4IFsTGqq2HqfuB9xng3l4pSmLkfy/RF
GazdJu1LrIopsi9sDFU+311eiXxXNqZk7LkwDLgmUtCAaYbvBvAzV5eTc8P6TXmG
Y4G2p0y06v+8wBs/OzHp2BQXM+0xKv1KoCf/gV0db/sNlA/w4qfT/IlTeoZ9Tlti
pE4iXTfEzX4e5FvFyQMBRVEn67TIE+QSYPzCyFVGdZr16gdPFCRc1drkaa3ECGgF
CaJqNxTOdHHGrhWmS7hPr4ELuQZuFcGVRm8svfW6DdLJZkuyhSZB5Y3NWs7yxQLa
sbSQi7CvL9xGzzT+qkCpN9RmlRm5M2Y8O4FKyAOGnmORv/yD5XeCxty0k8F/8Bxh
GiDysdfec5pJlUInVUL7vLuKa8CrMcf4xvJj1Xn/kkrW/76pJmEpjVGGaPhO6RjO
7aa80uTkH2VC/QX1UP/futu1KlzKUl1oSscOZ8UfY9Utsc/7RGOIEhNgulRF9eEy
KFWOepVfg9IocST2DvfeRp/32RI18txxCnVHtc+Gw9jNXwxo5ddsZj1uBQpZKXED
9baEAlt4leqNfw7QAZAuujpyBuO9sa64PS0AomwxU8ldJPVM+8qrmTL7jXMtVw4f
4GafLeDTqHruAivEnoeUbKWRhIokSQf7MOjNwVseLTNed9busnI1/JPRQCkDkzvD
iesmXu2XlxAdTAA2QAfnpXZW9LnSCCDhMYbHY++hgz/XJaYfMRFIhTKCmMoucsed
/GmK3vgQQ/ldN3vq9uH/NprHs/sDv1VxmsPAdG5p/r7mpcnUhTEdUXBIA6LZUrt4
NtdBm/aolK+wdTV50+Y0k0dpFTqbb6XecLP8KZW4EolGmjZoWnE1Ho3Fo/4KbzyN
ILnu5vKy2lNl17QU/eq44wk093j2kw5mbRvNMzHBGNf0YtdbnmpBgXBM2potYTij
VBwebf3LkWMC0CCaIl0HSupCWWeFeFpOSCH6GF/OfHjJnaLrSoANYkXuu0hu3cit
gWiPO9nJ4+A66yCzAP6IWTgZlZ10hzK8E02t8xKj16kAxK8iXJL6ngzspwOfkV1q
KX2Pz5v+tDwPriqUquveNsDPprbvmV2/69zhKzI8l40M+puFiRvOjarEVJopThiP
L3VsLN3CDc5ou2ti175MaBQoOZ7Hzc2v+EOP4gTAHRLRBTRp4RL1e99JF52z5nuF
AYMiEGA6Srlv7cPDINc0ZntZVEZXVMZ1SwZZUbwByelkI6SjcSGHoZsn8lrW0LCb
3WnrCD2o1JjscNJ2kIf8/Z+e5qoGus59+CDiLzbv4H249mSe1tJj+Nahs4DG4sIZ
dAYvXy7k1Ml8H5FAasZTf6ruJImc6kzcmpBMGU6ov+L6jxT4gQQiI8DMLYcslWUi
wLfo+imeMLh9f3ZcFgkUPPSOfygRjLNbVblX/GKiHza1wV3isUP8Iku+H82e57o5
2mP1VzRqx7yxigZeRE8NwhFMKhas6TuO/ix4b2D2lHJvDGyBNx7604dYeLWII+Yy
Y4GZFMREFHa8aXBxvROo6+weIlAanTSEL/8+PG3N7WF1L3f5x6ZB4IknxdW0sLJM
5tTApbZgl2IWa4+2zCR4h9gPZMC0+7agB/e0HTzELRz2qnsIKqdJaSyq9rySdbTK
ReToI323FjKrpqXk/JzSBiBMqLvtnWx8fq0/liOnES68menkf2wVLSeUBRQ2XyLJ
uYGQdH5LsJCK9vH+bk0f4UqLXQDGBecwvGVKltOE7SuZPu46EjM1Gug6eOxATL2K
f5kymQNeQjC8vlD28fxJhkJIPqggAcPtZ71Ndh/Oq1UpocNiaesvsxxf6dB02ESN
uLWPZrUcI1MXL+l/LEkBLkAFsZSRRnuWW1wxTDJbq311bCD8b6tGaukuFPTf0z8a
n8qf6LWTdjJoMtPkvXBUvXwXlXTVzFHaMsYhE4QEUqSZFU/icBelzjEFwM0GWap1
dxWOmHkBHUbrSvz7M71Or+bWbcbtlOzKgtpWca8cLXkwCFtDJl6bNrQfUCduedl9
Db+bDgbfHZTRXctZE6xAm62M+Z2qA/oEtArMUHsbcjh5gw/ppH/2Oap3C9ijc1jI
TArJUC53TKYpqTlOysumVV11RlmvP0/u4qP+v2Q4K5siS61BOVyaOSTBZImfNYpS
6FosfJbIGnbcInrtlL/LfPtx4gqzBgZpBARHIl8KC4nDieBzA89QcDsi9jrjrC7z
JuBOyCS9jKoNiEBb3zX2QL3wODLzVoWWvEjP01CAGcm7s76bK+RCBz2UeCaILf63
R126maxLQ8roT+jFuNLwF22NvOWVsn8t21TkX10OeZdCuMus5MDHjuhhdwm3q5Qe
Y8RaqASV1WYaT2IhlJRoXB7JIJyR35HIE5PuS0Mbr57V22u7ZpFEB/AHwWFhtDG8
RDsMMAtPbs700bFiTsX328Factc0bPvtDdj0Ap5e/zBT7N5Y6DWqw80P6PmNOxYi
VwoH+2nKEX5uJ2AyIHapJbm8PbS0YeLJI0rOtzxelFNQ7D0rY85TwV5feDrh82/x
YndsQgLkZymP8U+sfknouIoDItienX89Lax2s5BcxdaI5MXpQ1RJ+xoRLAeFo+P3
nSJyrhxspPLCPhEMzpVk2lSx5iyoHU6dFevC9nOYtgZJ9aI/iGD/nT+FYxEuq4K0
WY96pFF/k1tMkTxtIbaDE1Xucf6gEiKooOkZyI3lUVBvJYMMZMC9tbteqU4I6/TI
n3FIC6lmV4k15QDtpPXxZ7ULTcZ0u2KwuSLJEfYl+GS/2x5TlR1jidU/MJcucEv4
mlo7uYlam1MlvJKzt/K/xgtw6DETvakzwNjbLmbvwtt6+RSOzSJLi4fcaqICuq21
hGwT1onbi3iZeq2p8A3CYjC9gBeGFe9+KCOYke3R9pUt56PQyS5CCnwC2GiSaK9E
cLvw501DA1qTVVVsdj0lDtbJ5MctAGSWsum1AyKl391062nSimbT72ohuEQUk+yp
a50R79McFfBi5QfOZyfvOvFxX6OWCJCYpRjtZGyvBJBCCH2N1bpntFwDllyn0mKx
GbiNCFHAr6YErvnATcb5D6jbnod/APVfa0QiotOkg5+BsfjC9gIYN5UqIJaNof1s
jSPY4bheAnT6iW+0yjqBuzScpozUiHdxHPSCtr1KnDIIKrHqW9mUFtFOpJQloG0e
32vszsI6K+D4JS48TSSct48UFzkWV12FyvTUNPbBzIK1MtAzUy9yf4l5UuK88L4i
raNK2f0VVgHi1BUxvEO/isOnrwjIfseJqkt7EMFyieYgqok8z/m3D4RS+s/EXPwo
MPIz0FPcKilFf8WTGDQqzXcJEXxmWFuYGmoh0zQYYpQ4lMLAZs1BtMTt3JQXKk6G
eo5NWPi4RmI6NY7hsccXHuWsJrssteTv+RQuKHoLmVj8TL/mkq/mYLuIzb6hpEtY
6Uh0FhB+Hrh3ibLgcDPu5Wjnrzc1YtDf6hip/FP+FjAGc1Dp3+oezCxGOTh9PtvE
9gMvbUnISfFrn6onbQ3TwgyK3gR6DGlAdas5rOu3KqVAROkbM9nCXaScLKvkArPh
JqZ86scxM9DflxYG+vLRhMGI3wEViKIPSgfH/x15x4ek0HMA+9USORK/DoL5r+Rg
rEwRoMWlal7Ncqy1kEkfsEFo2tWV631H+JOT/SJiD71cApGBHL1Zd32OMGV63Uys
E2x3iMPiLx9Yg3zDtqhO+V14N9I/JCfrIF+0RwTTqz9QbzErbThVxW+HT+4uTq7p
WgxsjAtZCKhpkvsq781Ij6c5T3euMQpMRCttvZkGFs4Fk5TNtoru/bvdGqAtyVGH
/MMxP2zbcGVxSevbjo4HuVKQ3FM5qMfulR7G8b5SLsamz7Utp3Iwms4FkOuWiKmi
/D8RWPQZT5I4Qh69o12iXQ6U8PuOx65fHEWh4OaOWuqE1uKIzE4oAvedy34gSYeW
2o2xQMElJNJZ/5cabUre3OcP64avL95M0hjUG2XoXdpllv2S8bcTHgoTFBBtTzKD
emrpXfrsRivSV+0x+HIlLFx5O4a+Z+vsFvUs7Iko+tE4Mn9tiU0ELnMboOev6mIu
SB4w54OamTvz2RlZjP0Q3ViHN5LjMpa4SRivFn44l1brO32m1VyOW9UgEmxq7HjX
uO5WZJo6jc+v8RA20S2SaKyiCkYli32QDtH3G1E9MKpqVxRK8re9xDAV8+MM7FVq
vaS9evYYzEr2CobX3PhyA5p11Nmr8tglYV9/Yl5rZ0z18iOEhX/x7EU12Z9JCw//
TX4lEpUovTltzYfuRzoienWWQu1WK4N/bZg8sNq6gpHr2O1Oh/WTn0tr/9OTUAcd
qdBG+seh9OMFzoM+9FnH80UMaqYYh33v4Tt/XTx6Is6knS4q9yFEnuTFIWsVaS2W
MNUEoqreumv2Ft90GMtjOTYGK/eLgYSkJTK6SaumPS76A4fq5Xf4sJQWBAuompB+
alETL7batef3OcEZxzuaYbBTOb6ZkImM6oOWALXtCOld6k1tzfL/gDp+m+B2E/7T
tum8Cu5W8Jism2epbg2/vsSycdro87r6Co2dOKDsUZErYXQgzdjrWSfwqAnj3oUd
6gLBm3Oon49YY90HfVq7tlwwVKFEyZ12ej0L13cCJfGhX7C1WfVE6g6UPwQZ5ti9
gWN/TmfWc1BXxYd1pEdOl+HLYs+tgD08gTlqygZzIZQZd56SJqI2Q22yl3qhlEFj
yjxYfA9spoXYse73hibULXVuf0seMZ1RLqNeYQFqI3UR2DlvQCs0MUFsHWS1eyyY
O3gtZmHBU5Pi4166mZ+zbmTlVCLIvXHAJ3QvX5fAQLyZAUoQZO5wcouPTISdo7eo
Zhj1VvIeVm4dZf612s2/CSH7XzG68NDeFWlbt8iCLWo13PMTykrH0T/ceKhwuyWh
h7TVdNitRPJ/vo3hYmPJzl/ngJMiAQgLsT0FLsenp37wTtHShgctaech5mOJx8aY
Tn5hQIe0Mv0HpgZqhAVtIZMQSslmcOL6f3pSH0UtRCG82AGneSpgc7Fn3fCVlryl
QP2bOd3eXvAeS7ItYS0R6mV4BMsWlSUZM6FmJLA7+05+oaZolMbAhZlEzm6vknXh
tXsks/LbTaTRGD/wWVWwmXVD6b4OsiCogcgECIWL+Iz8sz6+8mrr3nrOVfyPN/Ov
vQ+qeYtCOcZ6MOE3gdUMrxGERvc2kILNKYaeRdbFJ1wSLku0VfDYKlObsUN4FFxo
toW5765pongM7p8tz0ShjaEkGWgWVu3I58pI3zDDbJI/Rk4sq40q79DXT9RkD+uK
O//V3G6FPZ222UeJksx4jlas/9ubo7iXdUIZCVznksUpmHixuLC20SActFQDtNya
r7wRHOpHcu5HmHZat2/MrLXACNpMwBPsWT/oyrmsxfImM4hNQbXNlh065TR84HM3
XOgIKHSiPEo97eByo6QevWsDncfpn42fPX9skAQglwH2NF5WNRsMQnoK/d0Gz1IO
/P4I/Owf5XOucwKXlaadD9Q1X/7x4IwWewFnG366tNpCyiTsZqGP5tK81tgJp2KD
8AUS8b/ouWQnKMuxSHs4VQ6BapgANlDictP3Kp5vzQSFgt8BMAoJBYFp2/PV27FV
fNJ6IA2UpX1SqkZk5hy4EwsfEn2VRdtIPxfZt0FbZ/YoNGxZPFxzRrw+uCyJJotJ
wo8LgiqjPCklpurEC9nPdxP7PbWJ+jJsUOTnFz3eSDzngITH7MQxWz6bDoWaUQv+
FAm3qrBqDKuVAnedPx5aDSVxdS9QG5B8rd2ltQALup2ki1OnxYz076VFehnjiepE
/Xs3xnY5F1+LBkFygWFfRWRDQ8fx3Kzr0v4uiRqKTpTpZfY2V3o/UWjKOWE9hQma
NGSRKI3/lyjVAoOgNWKTu1Pw5B9yx9qzEN6PcEZ4M2LD/ZzVsVwyODnmcW/ikMny
cqY0KgPU7b2CvUxer84KpTeoeMEB9L003bdvTJ1rwapt9sDXb0mUhWCtmTSY0+9x
oA9xZZdHEr9MiDtwuvapC10T9sQ4NFoziREtot893dghhNylKK7I3T+ADM0o2yiA
gzVggM+LY2zlfdiHAQieYh3cFC4GCk42zl1V40koh/YRo2sp8BtQ1gjCPZ7upXBw
xzCU9JECsbwaffOCQJs9jIYDcjDapV/mxRiB4Zm7WMaQoL0Mi9qJFij+U/FlrmqI
gRwcckiNJvfAYx9SpqOewWYaiWBHN6leh4HGcLbta7WYi1sVbSrlJsobcQWWy43O
xL4XJ85YsfGDKsOwELpXBGeRjkV64X5/SVlrckfs6eebeeNVTTSTdHY7V+7e0CJ9
eeeD4tEyyg9iwXB3TYa939r9Biqxvzy6yCzfMYZ1ingplHNvVGtY8srZrd52hn1m
+7i0H9gxtFxLp2oCUYLNSO3rvnI6WT9FocAA3wSPnA6nW7LrQLA8lKQccd0yb06y
934iAvH6YyDqIg6x4iKTDWlkbE8Np0gRvQj2AwCjKcYXebb4hByv2u6zH4XQjk94
MpcRdQTXyHOx0yXhhAVeu8fqKgElJalK5pqixGx45WoA9SBNgXkjPwa7C/lhK3SJ
X/im4H/hHgGvt9/iJ2JvOqjbseuI+F7DVjPpg00kwBJPCBW0spRZ+8ymFBA+fUwe
h4G6KQf6AIMgw1ksWR1uNHurRIh9H8XyGzRD2KkgJI4X447h0SPEluE3BNE4epIx
eYY3kJHA0QBY8nzTnr6gYyN1vPABU4hdnR7woaIW22btLnjRu/OOAB8d0t+McIhG
0Xc2h7but4syOa5A2wRonvccIOARx28IBp2JkmhXtMdyH+cIIOeWVcwiPPqXaSAg
8isP9lb80g0OrRsA9PA/q/buFAGqZWYntWKTKy00cRtIYsEWObr2HxTH7eKDqJUk
o/qMeKuq6GkoZ0oLW76UPRkR/G3xhOBjKwqltItBrYFi8SDWC4AMs3HBRfZwrhTe
13rfc/JndG3AZWKAQ5UTRfDBw+LWoF3mKJisDKKdS2XuNvwhioTNpYpcaE+gcFZf
zyDCGMI3Iq/6fXDxidg49Rz3lQ1z7mBBKW3UKzdb6OwV7OzOxw+2v+BgE099DWwR
LJcksFUYWdSHj2qYnTA4uqxAFLHW8oK/etfcWndyYO9tAjzRtDSL4ftEO2zJox7L
26kGmWhTxQN9Cizzc1hwVHYr/Jt6midUYliHVR91TUoFWjsR+JKOm8bDzZDQrF04
Pff7IR0bdcZM04+GhG7cO2g2wAPjGTMb91fETYVyjuvd7dqnPO7ZrUp25ZlUGP6/
6EWREeQ+27tWJN+In2Cry8psdLY8y+DMW9ulUeoLSl3gsWXqtH8h09H1NoKL72Yq
o4nWTPUsZsiesEydGy84/31+2LWYNBObXiMXQSFqkSZH94O3u+o8PkouGcZuY6cC
idW13LZi4c4ZYHXgkryK698U0CZvaTRV9SbvE63jcAbWSVjqy+uksZbTTmFbDIcg
TwJu+pXseDWhVCs+jGiuUwtfXGPxkkLMzWrdeGwwtJWovTvWpexPXSVWaP27ED6Q
72XSJ+GZm3K1fpIhMw81aTXC2HK0YDWSLmKAgVlApKPzD0V0ceQetwZseu2CsfGE
hhqtzDRfDj2I+pwVA/3YH+SHvvdTBNp+IExTrhm1d/Ua434OumY8Z2mlfD4yxJhn
cOopyyjxOEG5Rc39kNZTfBwc5h2cBcQodXSfnI9mkHSMjMiZzz+Xz/bm5ipvzu8i
kj2+JOEJvsjccr/MofwSia3jrsSwMMppkpbpjzc2x7ub8sDzASi0KJ8uGr9DefL6
VbeQ22rPd2wxRxkt5ypKoziGwnBt3Ys0NERZI1+NLTYF1SE2538FFpY/B7ukmyLl
vH0uUq9z4xQJpVzBChg+1wY8QqkBf4XhdnG6X1f+W8XmP54fNengpBQp08x2rLyr
QclljeWzy55mW/lcvhEercDEmCnwlHjgFEvlJkW8WhgElDcZ1NPhNI+2yUN2keP1
5dKFtTprw0/5ATsOZ2QUyM6BL8RrpUeCaLggTHtQOlCPSSUqy3LhV8CIpwwBqmu8
61Xo6EWP6lxGFFbDngrz286FrRjuKTYB59XDcSMDhRFrGrRgvlok89N4Os8l3285
f8hrQ2zTydcbG+PJM8LWpOdaBiEXjwuGoVCTcB43OYEc+e5Qb3shJVWkgN1iNlzL
HzLcDLkvfhml9f3IF2Wj+BUAraNH090kMW9AlIS2GhdbM+aKvW/0h0qSOVtSmzom
4tx4lJksZq0HZ/eTyH+xHzkb5NoB4FKrm8DRRRuukdDu61XP2wtQ1dgmiS1lOWDX
KzPhwhwX0zWqPKEgyCZGAbaa6ti0sByzg8g0YU+zxNLNz2A1oUHWMkR5tE0sGbce
u+0svHY0D4dbCl+YYjL1uGx1cY+NhA17jRDLiCkFKfFT4vsouPzxhbxRHnRbiJ11
/YvigrRq4pJlU0bt2BWw+FT2WN0M+g40ris7pdgtricmq/3rvHMZmD/XrACzB2w6
aHUrc+nA7B27B9KPvFVUOI6mkkQeFbqdNLhiVZ/7R6Tm61wlflqNJMlx3NM720TS
VlOtdKgXO9P2jhOBJqUfNr+jEHlCJaWRoxlZSigBSvb06++cPPBXOojspOV9+PFI
qJj2zTmPyOHGhAzF1fXAMY+iGKKEURfmeze2BU6FEHFcT6AyBSRrYJsYYygxMbmP
Lng6lVhU1Z69ceOC+2XZakFYZNClzL21MaaXe2t/gAXw2OmuMmaWCy42YIg82pv3
zfe6/elB70szc+PPnCY0itMq/h58rwbE1mSzbF40WB73d/kstIvvXopqYAMwqZAb
Dg7CZBvSkc0wgLigH/bet2evVWsJV1QSjB9iTKmgiA8bp82AHj8QvMLGfJu2D6ie
bWzTAvytzNHA1C3qbQUSzniIVaLt8beNR9zQaIPy/Fe9oVaazP8NuH5a8CG3I9p4
5Vmm8Isj+MqDu+1f3NFt+pzwiQ6nPsQtQ5mBFjMO/vuFEjIECEb8v3sSQDL1L5pY
xGiOgVPZG1XVL5Jse0H/eBImdpIbGLjhUktwoHO5QSrGaq6IHeYmf0UJweN99Roc
wrLhoJPue8Lw5AyDctXj9wmaOUGwmfh6Igh+D1s2SwYZ+LvDcUs3xmdQgPCnUmKU
GfEDgeqmtyr2IvF+jo0+xdKp1k+UL+hC6XjCiRTE2NCJTZmGUDV1E0JFTYM1Bfkb
JkEHLvykvJX4XmzauGT+vwpMzzS21poh+OddVGt5kqC7xyxlZiAzs2R3xuK0lgfZ
qBAiI+MVeRFSZFuLBevVMDe627xtFHsIEfmxnJ8c2snbYeoV9tlTUQS5jUmWEqxe
8o47WorncVVk0s7st2ljeL3QhwyELMKiLcl629+Jzd5fLk4kH5heQ9XmRgbgh32x
YvS2dtYIe2OH5ZD1l5KTnF/It/+mgmlf8BrffCTXCyBZiEtS70DdAZhhEbowiXld
gea+IdYmwkVtDI5ttumY/Te88w+3+h7yD7LouWGBANVaWJAfvi4sahhgzMB+S1rb
kwHzHpm6JNykA2IfNv7kncejSlYtSypLvLiD5v/s0QDLxsFBg/01wVO001RXnUiS
+KobfkyJfPhuPswsWvYK/aCGeFDIWnRtCD2yZOse+DvLnvKwYo6u1/VzCEdWgvBf
TELs/GWk8PAH6OtSJBtKgJnbIB2Sn2tn+pqcs5/y+NYHNW41OLOYqpURkIAT9TX+
F04LmROhSydXa6CF/M5jpjlzWFE57Rzy7VtGy4MUL7eHPvnrtSlqjt0AAZ1VufC+
BsJktMIdwEGl7CfaGszUZXY/YiSQkRgvnO5ZiWo8to0G1YyELBqpkiWCSL6cBjC5
fIl37+2klWuMUNEqjeOJ907ZY4cO5rfYhebJDcF0h7JBlFQYmHi//0iNcIUiLHcz
YOYh4K2go5IWY4pNgHugC5ZXJC08C1j1kHgy1H0/xt3nnk3awabVugOq6scgE7j0
nbk1NyBv0nK35NbMHiHxP0KkaV9NE8qOFqjjCqnBh+vFmJrJvy+3tCyCqE1q0wiA
paPilOegyq0ZxboGz5kB8XhRuQoX4unq7S4zEBgE0VyYfFc1RyXX2OszN3s894vm
4hd+QYFkKVxkW4r7PFgIdFevSsljd01TsJf8nShU5AdjwHCANb/toFYH/v9sIUAj
zVVLRVp7xzyUGsN4Upm40Tkart5TqyzGV5MXUk7/xv3mzspFZ7o7DHF1WgR7K+pD
R4aSk0JeFZEmOW9Fm6DybwfVWGynsm3Ytz62duSFn3zHwlwR2R+llCaUm+sI0wHA
xehGjP2M5SrIBRAel00O/8aqklM0D6dIQjZsCspaBub3j+mAWjlk/wV3IpzHPy8d
uX73AKHdJiYCVjKOpiWTmOiuCbOoZsSWqQuRIZFi1+8xXTWwj85/FpF1ZPNXCV+y
Z1On5TBynlNq234nc1yr0Ei6pem44Qi4t5epOHW60wWkaJvCpXdDa6jIzLJcftMX
n06q9sqW/V8BZuVGd4jvENmUmhdGtnShYjReRLgeFbainxDC/8O5s/u/2MoNTOPY
W5L8Mic03I6gdbudfM07LaV87LbN3IG/6ZVkI0SwSLRFRghjFOSjCSJAbx8KnaoC
u/Cuu7vdkQ9f+WRxkYpuCEFN+a/rw9sPW7ZltqpbPgST3B7FJsIh5r9jMxedxfIy
UuM6afIg5CgvCQAXasrKDVsCQm+0fL/sMwYv1mrEHRI9jdJwKO+ncZ7bjWjPVLnr
bDD97C9YMM4Q/m+maJ1EzO6w+U0hyAQNOAu0egvdOPih1FWG5QyD6FRyVbs8ZRIl
IvpCsG4dpnM4z8k1O/uGGiyYilDfHcMlHAdODpPz7NDDDNRD9RA6YpIGKpQmP2V8
4zHpift0wDv5/BRUL8y5fR5X6irqTKIN4338TtDgo8jW0wEhfuQMT/4Hop1PoQKf
vkoQFHB5xun8K9hTGyRqSV0THUyOSXGoqziJoAo9URsyq5m8zQThbpKfTii8Wjx0
1tQAOoD+W97klKNtG7+m6A28AhWmO4aIkeJJtCjpG8Bc2ARr4C6iv4xnUs2wTnaD
auyBbJdkk2NziBwlveEZvr6Tiksxtu5eV1bPve/p2VpgVB2ZjhG6Snn+jTGQapnc
P+FMqd7QLEiae4s036dxpW2951Y/TMIS/v7aZh9Mn4jHo6XxvwQ8+mGOTSx7dXVA
9mEdLdWwnGAsw7g/wMH7bEafRYhP5b3j+lucXgSrVSX/lXuYQgiQXtrAAmP0UJ/V
86SrNiflESNV+uTM32CCb9rTjQr2W4k5OKZz+z+A1CJdY/9thnGIOH41QxKa03Cb
UHDArfZbE7OmJe/skd+i+OidtTtYfHpmfM5lvjS69Vzr4O1kG11+bS2WAQzqxvRv
ovLXZz+sNEYg2+nv0Pmh92HR+1q8mhG2uBnxURQPvvTpSHtMjjM7fUI/XSrFQ9zs
beVuQkLq9Q3Gb2cgAtQhFsVEkbrmNT8hg72FUaN3S20ap187msro/DqWWY9YhBcX
xMtKxCeXvtypxDMjR5FLjtBODVJyzA/ZloPd/suwkOHUz9A9/CXWwd/k0SDT4mBN
EOK1MXJFKEf/7lO+2GN8JxJV8SwxXBhJcZ6NMDU5QWypQfK8PtGizWb57JapVTEO
qItaQhi1BEX0EsklWa6l8HfhgbqQpNbZRhKuzUYFzbLLIhFRWFbv3sKNAgGbRu6G
Q6jEzF9RTN3ajoXKIatmTgP0Wu9aYWH3xcW5sk1aKtk8eoplXWSPHiRiNi3fXM8a
Hja070lbnExBKrTJJHdZ2vU++y0wOHgVzv+IXNl8K0Rm7nI9oAzHZSAV+sdNvG1+
vxcP5NFEO7iIYzl7GLLBTZwxifjHyyfNbaf5akUcOoz53vsI0ABHSluJM6/9l1Jz
no01fIDiY9ZlK8x8ZwMV++vRGmiyoKhHgqB2Xc6rWCAMEGlQxtrHn5QaOsHs3Twg
CfkiBkoQLWqwsB1spW1yI2i4yP8Q3DdTbQT1NuQ4Z2DeEHjfo8JEr7V/eMne19zm
DO6ZmlJI+U2BkmuC8hIxxaJIjw+9Kn+G6Cj/i5iY1W4sRuM7lUFaNeKb2vLhZnAD
eR8dCUPiXPAvtrKrIWjQcM3UkhGbI5OL/iuW5yp1gpNdmsY3AslDCW/WdSGRmb+F
whCQ1FMxiXoD5vE8hUzJ/IzFpuvkISrtuQ+bB3DiXZeaGrU8UPGjs+Ios6HefRhx
2eLzQr9R5hDHq/S4NugCCe2Waf9cwxasSVk7wjsWp5e7IYULTESMTGemH63vOiO4
coXyARDExIZnwE43ykfF/kTfBTwk41R/iokMC63A0d2oXRWabP3oK2cfVsws8Pz8
SMSDd27hZQonxM9f52Zy0hUUg1VaTzD1m2fHvuG4uJ27F0b8uS3aj3ihRf+oO9jy
+rVNpJeJNlnvbuv6ti8UGyxXl7h8945bZpxGlxJrUzUJZJv/T5wNZkBa1LPvriCd
p2od3a8z2/0jaB9I5rFkbX6LuiZ0F40lZ/d9zBjyw2EAh/W0znBJCYdRlcaW1Sc8
BUz/FZtCfOX2tlYAQxuNXJ1TEv8nDs0DLZXoFu4jF2/ET4aaPlwf8yB4Dhvy85oO
g+uzki63nFQ5Iy4aVwdI6DmVv4i1oOlqQJZGEn3BoVJpRqa+81zNgiMM/HgdIb7a
VEdWrs8cWL3iVmq2mgqsDHlshJ1QS1e8T9Nx2Rgdc/3axCXq81iHwSwyb1zoXv86
CZxgoMoI1BlrLjWacmRU0VPEoONNSoCfvhZwMt5N8G10TGLbhk7eUgHgurJ3fhlU
4OnUplMx5CCJsnLml0xU3orGjir24o5yuG6PXc9SDTX+Wh0MQ34e/n/qiepQmWE6
IjxgWQMFgeOrAazsluUOmfwJfENsSPXvdO0kxB/F9FWiQ/XDoeSb25FSAHycnBbn
0pXzL2Ln7kJFh4gDgdQU/JHEYf1YzRs4EH+3nCvft+MUC2Mu9xGVebDUyv12EyAq
IExh6KFBSWrYz+A5UE285HKBIK1gwABfAEAFzo3r1zW9RqBKszxR9lbJeF67EwwB
9KeJa65haLF9/0Y19ua+JGRRiU7zVoKMRVwY6agH4c7jpG0Ad0EqaXWe1V4gfURS
vx1I3JS/QvB+rpASHQSTBAhDdLRIP05cyWB1eUQcMUDF6Vfech7Dk5K5SEzTpAwE
TiyZNV+ysRUE6z43cKZRyz08gdT0AmAhmtkAOjljF9I9JN4NkV64Gymctmse7FMr
wQbXGX40leXoabgcQD8MxzxbmJxqO05jUI3bX8jRuQ48XMAzfbzOVaJ0XFp0X+HB
VskMsitwlKxNPFCpQR8ksxE5xmol5/RWr9Nq09G8/s4oo6dTZGlum4Vf3OU3sWtE
k+wVIeA1eAs7HcgiMJ5CzGX0sqi02ovOlakh8Dwl27QOmgc0QeOgPp3MDqvTucEy
tFsjYG/zSka80czWR//4Kxn/OdpFV/KQEZN1IMLcfL/FvwHvQ6L5naclLo1j9ZPL
AgYTdSSiQ17MzmKYdvO6Lr03KJkg0bHr+eq8wpEo76I1L4qe9c7UNxeQfJqtbRps
qc8aFLxwHrD16waVqGQfgVRZRiszt8zVi57zjQDaSQzbISPzT6fWph/RP+FsoVzx
SWcfu7HFnb8QkejC3fHZ/nNICzh2kuibgYjyfr4v/r8DB3LUKNpDxoslD40N35nD
REjsiOKR+nqx7NUTlyE+klpKbpP3OXQcoeIHyHSdF4iuufjsrRc5sSsh17CNJwl7
V4/3hdLUNWmVXHd2PBpVDXTTVnq1ArIucauAXbgpz33vXj6Imwjw95miy8nOqDhT
eHAiXgfangFLPdRWuf2MNGv/VbSA9d0s2lWJLiOO/6D+Gu/jMfpCGldOipU0Ev6C
+QZbtvAK6ISxjs+HkEFY3x9X7miALELirrRZqWFV0DZhXZ3jJhGy9XQJxKVm9F6L
zGnZXOV/A0lobASc/t+bOtBI2a+dO9RQMCzzYkv3j6h1l/y01WU19lvJkSOY8Ni5
gkAOpCmsGNxIoOo+Wn93H4n0ovspKPsAUXcdZaHO+dzuBM2G3MhmnAM1myGaAhpp
mqriWldKIKM7QqAK9P/QB3SLEiEg+/GMhuAvCXLkbsuuBP//nfn/WchJkXHXlt3T
CkBYpe+Buq25Jr75rsPb9V3Cc2/AbDid9ziUV5f406tj/lqEDKAqD1+dRCBXR8u2
TglrrsYpyTvoZlxnJry5xBzYA/ET4ucz3AhRyHJb2X5nB8lO8yV7q5fK7nE5CWu6
ZhB7hEpU0IT14ldYFl9vNcbevYfUAFN+z3heFmK+tu+rGTdnf5zPDBcqwMVzhtr+
TkJSBV/8h96BQbGbW1YivG32YrxfUZ1JlVyk+fC12LAKuCR4e+DoSGbbecq+0POh
/h0CcPgYvQLy8ZRQXwm7A51knqEV9S0GQIV8/0Llr6IAJLY9yjFJfLraBiWIo1tn
x4ojRr/R82XbJseUkbt0U+k/Ok2RBchY0G62o9pjS7rE8DfTiNtUIUuZBODxy+Ek
DBPu9ZV1Wdg2+2Jzsf7FIwXr1yb13Ux5Pvulh0SdAUqu0xg/jlqfpidmVEklPrH2
KJKtPDjiY6NE2nE7k5fYY23mX4PV/RZn1nsXIsPUomO9gr1BvAxhQAiQn/ULtaRt
oelKGFV8b7DsPWgSHJPQD8MowjaNYemBhpP+TdLCpE/FIAU9bdigtzp7l6jvjk04
7oT0PN5HfIrJQI9jz9W+xWsxh55JDT+87SSX5LbkSQc5OPjfoAOMqJ5/yeHs2HyM
VfZu3dEp/ANH0MmnJGBrfVG11sB1SvOcju4T1bHEl2wXymAuvmac5IcD3cuJ2SVE
iGbbeEXawYSMdorPTmh9zES3J29Zhchohh7k17cGEbUywXNTsJ5Yh+iCDNJRUbu4
YYcq93naZOUA6WTKrQpToAZcEpz1cshXqMGHkfweyELb7yYHS7w/tcZxdXPfTdZ8
6ply5XQ1+UHW4GwdPdPwFr1CMBcchpzSM3PaR7Pi2damM9z8PMa6jE0CUrH1WJoY
TCJItkJ10QD/+akDn1We2Z7oqJ3Vn6yhJ3veHIQiXiEImNZyxiqkzVyOA3BOtuQa
/vj0X9q2a9+83Q6wMOIgpyWVBkLW/1gRA7X0E5V26ocw/52vh84+0FSzN7bO1JPO
uqMqU0KXqTrFQ8achYW6sWb65mgJxj46D5YohMNZcrHAehLowLaE0MSFjPIbdK9O
FnVbYM03V/fZuQFA5f1n2nLoIAp29maqjXILwSqQwBl+FDw+KRzl633xf6AB4ZQ7
iAYmECbOnexxfCHIYOT6g94tC/eaySil8IdaWoAgDOjvjlosOOYKaloEvnZ+K3JX
lZYUJyNEcf77xUmSmJqFKxyQC6gEaYLm4w6Qa47TQsIspKne6XWHe1oMQGoxTqkD
S3dAeBGBFMF7oIn/OfQ6GqpFRJfYpZHMIWsQZ2en2AOv5TSBWcZFVeyHtzqgeSJj
jsCyGP74TTTn8ckDmBLvDcysmpV1oCKbp4GnkrkKZ1xB3Bzi+8tYgXXYKfpWGCUy
Pw/qSp8+hPH2JdyX76DDvy8zRTP24vNQSl4dCZSQFRjozc1Is3nQ10uDTanO4FEB
lz3YBjtLfQEMlBN6HyiWyN77PD/X49T9a0LkRNRY2C2LMxiYiShT4JwU3gVyHbmn
duDUQ9I+uH+caFerxVKSuahjOVDnL8tnVU2Qmaf4hXMPcg83/raENA+dFYaQBU1T
xiOSfgf4pHgsJBssMvG5ztsheVaC+b4IOZmqopOWNqMIpl+RFNYI+yWobmiPOhjE
JgJqpxW2nFXs0o1cDcaeLH6ZkkPi9a08FpdUXVcE94gOvgwa45kiX4kJDEH9jDsi
pfE2V4IImqrdMva31L10rQXkmEqq2w9ninnThzg6rKDHA8DbnacIdF+0Yy197gos
AgpvR7XG1SHUx4m7NS/zB2qZD1VhbpWkybpa5LbIpy8WtX8MdnjvjkCNTb/mUIfE
T3lMDiIm1V+ddSwjSKp3tY04pm/s1I2LXg+f6hX6drjlUObFKkSJdAyBrZzVaA6A
3U1wfH9AimwgR7khG3N6/Ni9TojGLN0rjlqlipRg+0sPKGPxUvUmrM/JG+R0EzKB
aQYxfsx0ap8meDqeZY6MoVZKHetgdOR50nILsgLzw2yQMI1EY+OHoNJha2ktqDGS
c3Zmh+3fIne5qhYM45WqjAtLswx1tXuVB0agJLGAcR48J8b1Y8qoLSwINfTfc8wv
p2HBH4QipuRZQMrAV5cKyvpQYy6rfPyeDUdtudKZ8y/kCx5YDoHMm6K/a9ByHpHs
mrvgoUDcYdiWzvV59O2dv5D8oYjDv2f/sPbBFx8h8Ieeh6VHZiNuVat2jWNNx81W
sjZqKn0Mogah0hSOd7wqGCpiHa7Xr+qKKPJt1GpVLPgHjLoFEL2D4JX9WQxCP8YP
RxrWjaknqg/QqJEe4iXn9i1GtDIU1SF1BHcp0XYeMdpgZRH13OcsUtVgHLgIqLNT
3oPo0cGXOL3ZhsJmJIfAv8cb9EK/h1BvuYm+mnPxnLKW6puEicEOf0Mg+3GGudi5
kXMx0ydtLmUHuGSDKxXjrsT9+v9DfLW8kkcDGGH9OvsCIDnan/D2ECkp6lj6ut6F
4QUAJcc6JBvk2m2YfX1i+8FGmiUcIOPj1eTkGywiiMWcG4qtUnt7nYP/tRGPPjyI
Wj5/gj2gGys5RXectlFILsXYyObI7ygK6zBTaK+RMzlp9m1JDvjZYx3Ry+T2mTPF
c6NWfbOfIMilksz/dWsYDp7yKwY3ZIqPjvaoyxU2z9KoeoGzq4owLB+EcIPCNux2
Hn5DNhHMDRE9g8P7UQlyEMYjUYFu3doT5PuRdIbL6/1JMqiuIrGt3zwrYaI9y3Vv
R/IBag3JyEreypk6oeVriXfgX/RRXL1rGjiH5XOtCX4HGPA9+ExNScmVyjtb13ei
0OI6GEeMP+gFsOHRVUsmGSFoLr8Z2aSFKTNDsvAErAz0/QYF62ibi1fYOqhNufkK
e9omOeEMgU3pzmWYkWZTV2iukIorzmX4JRsr+JuBm3vZ12BoHxm2nK/LyRRehjRo
hfAKsG6KGXr5LQNM1ZDZBepgqBUvBuBAUyp0DvMf5H3d7m/yejGaNegNjzrUcqF8
BPlf+SlINy/JnnZ9cjQnx2HQsBgC5/6OoBxQag+ZKnRu4h5xnjDH0dERmwFxMaOR
k5PXoi4Wp4dslbW9uqaO5tRS2c/eL8CGyysW9DhK2i4oYdJDzH5yzMY63a5hVBme
e5U+pt1BDuLStwLka/XugftZ+ZjUnRqyC63pMB0xXD3NE2fESwugy9yD8TGkSCMW
MIl3+F2iqq9zxgtmX50GFF3MMyFNIeoimUVqvTZB+Jf77SWNmkK1duFWZr+cAVlS
CuIZh+c9nt8ZNi8phF0KWbH/Pm1IZaBX6hLKiMoe/XHTggtXw1SOzG1B3Gou0Vu5
NrHcOw4Be4/yr/mN1IUWnhNdaWPw01y9txHP75Sw+ssRgM9mJIdW06qc+AM/6tCm
BJZBD0YWJ+Tl84qhr9+27a2M55xVbIUXcBQxoCes7SaE/P62dMZNdLVTvxJMNCKY
1ReWZe3M8yl+m6xT4JOszwsPUftsif+U1E+x/6rvRCWt2izOiprGJSQhJczTacJW
qXTSjZH3DuFm0aRfhx8oT28YUiLqg2QYzpV2cEoktD3x7SrEJo5gFDVZQPuqk8UO
8HGB+otc+9UfG100eg0pxq1HER/nS9fQC0sXRaeS8vuCGckyMOt1LWqC4uIOU/2o
MUeqDzZXXakS2kQ2+74aUc8rUOHyXElmxjGv+TLpFMOtwSd8Sfq3ZoCC4/PNi4ZK
fmK3hiNuXGDSBdBQXoKOWPCg2dClvRetNvdjdCmdtqvloNfuk5oVF4eN0/kAzJ9G
DMbP4oGuS9SBPZeYq9q5xL9UiFZlqfYcrrWlJVHU9D/npXC4GOJCg88STG+o5RtG
UIEvDSeed4u1q3EmA0cyHneN1szdpgc9haKulokoD+dg9wB96quPHtsjpXFPCnUB
aQY3KO1i/L4Mh8h80d7ITjYfU7AJ02PGJ/rPVZOLx/gHBgXnSbpd6A055H47A4UC
zkyQzPCwYhTPcGWZ7Pa27VWoKmEBOgpwOsAngU1P2cdt+9Fh5cAteJseF4FL9HY3
RAggdoZHPyPgPoXI6Pj4Up8X5jbrpGiuD1xNNeFQj6elfxE0sYzdN/F3BzbZZc2s
jbOom5xABuQBnGNVt21w3Mc4my59QGjYKgyGRQ8W30bK0v0lqh4RZMRK2g6xkEnu
Qv7/PacfKjUnPO2LuHh2O7mItJinM3QJgjIYNE00PGtIqzOEPIJCmZLsbp06oPkW
7Hljs/LMJV2JuiLwTrPlbWN8Ypx+TmsLi1aSEAi+7Kh5kEDhRm8KiU5wWj+NhHj0
QGE/qIUmj39+yJhfJCJ8SUuiougE3Mo17Mz9DOlVDTTdpQb+dcFi96H4zEqNS1S4
g/Cx8L2reY/IrRyxLomaNxztasO/0Jl178PAUeqCAvFIv/pEs6qwy9xAeh0UDZeD
1YIHTLGBAGMFPFu8Nw81WQO6HZpa7yf3n0fpEqbuwsWz4YS2yJKInu9pTn5fgMcT
ncTGdHdOg3t12nxWzeKGsOaizEOMM4E8GvluzVliNw4lc85aBAU6mwU2CzIWKy9t
aAGLFv2oC9iZKeRMv5GMjcG6L1OTTLmjBsw7miXcVREwFirTTvUMMkdtfPXOtJ+q
vRcGQlTAThctPD4ktMCIB45Fj6tuDnPvOqNhOwfJ9pvY1GjogxkOMvVvs2hO7TE9
oOVty6WE/eXFbBjSWsv9dHhEMSx9datq9tZ9/SsqwV94rywWFuhj38IydON6iFAD
3c7WrUbm8RQm3q2foQJpWm/b/v99uVZuVRM5Cry/pzh9ZxktQKd8c9usjyAMgF6k
/GdGo27CC8ShWJE+BfPgKfSAi+bAdGW9W4B8Pi23Q3rMBJlnCOSoP4q1yt5VLgOa
xNcnv7ZYSjco3kLOZU22Md11yqFVxAfLgUcElc9fhroTnu83b8tf9xTY3+N/9CNn
Y6VjGrmTdC6PQiRNrrzGal4fc/rr2E9kZYKf7JI0DeU19SoDkYRXO9TmTVez8O1q
oFykLZ/dI2KE7hZnDtLEra28oZQzy/5mbEgnvVkCrzQd+c9cYIb7jy9H434hOA34
RcLKP64+kdeRnk/smRIvAMzDXTzkQrSo5QgfRQfybTrF3IOO65iknVBeLnbFb1SX
eyXXggCnswnA+5bNSLUJuQRaF6gsdKF2tU9KQgCGlk3Vy3ySQfuKKqx2OS0G3srn
E+rm0bpTF2OGqlqVgIExaO+RqtMCS1W2Qee2XPHeMVGqdf4KUBS2Ij+rpJuCxbJT
5VebTyOLvRVeQgWmD7m+tKq84ac2MkteGt3i8yYsTzJldLX1u7M7Ok5H6yiaEs81
DMioL+aOs6IP5+HcHWx7tsJWKD+IQ4Nt41mxTjJG1uV11yAb4QhGtFUqpJZ9OWwD
yaUwHguROpDycGODPQBPTiCSJqZsnPDDNECnm1tYkYCd+hoe48TJSuLLXhQBCQl2
2NES6i4gi0tro7e593Sjxdijeudm8/Fuw1FvGa24/IOfYnjv3nvXuKWZVhus5g4i
uZePsCQoqclODLH+HJUFEF1R86tm8HoK+tjpgfsW7dJZ4qWczHsmyAwrooWK6b/G
eVBrLteQDl1uJHjN9Wdw14OxCzPF140TxtRRWgHNldfk9Awoa6xtphbqX7U+B+0f
GMUQjiOdjV+tLLlWaVCvlQRotq/TDz5lByufGKGlR0RrnP+JrcXYkuvHLbUERWGI
BwiMXv4xPfA89tvEQKkCUqdJNzjQxvUmN3Up3cIQcwOMatFsUlIJOpBowgdHMPeM
MQn8mx/9MjL/eZEi+XA6DmK9xfRR1vStBdgPlTIMTrvyRCAnss3pJTG007hoq1kX
l+JR507naMn+eG63wpp297C5zr0C+fvhwhnkwIxI25sn3lXy0eCwqzSkoCjvvC1t
Gbv7yHWiSM9RxUIOfwxQax4+9eBRFrvXmj5JVzeb9FP83xAb65m599qvtKpcn/NB
CDX+4C7s4unLrmzLy/Quo6RryNLt2PFFiZBp5dI8T3exEnLrMbzIgHEXRVQAwUIs
HRLrycVf19j91AghVODWJagfFvwUEPVkR+5eIUXRBVC2XTIkDSACDvf+XXcTnU+t
lfLQEmGwy6CgpktTtFNvbsKQ26YqWG5qFaDH3Jt792+9qR1a9XGejrR5s1dinXoC
QKG3dS+AaWjnUFh59vDdWkw9h48j7J/TYknrlP5/TL9hpah3Afo/Nzlg1YFBTIYu
fISxXtBPwZ+gPxpY9tT+Y2/GkFWszyI2yNXpf8+iOCdBIeCvcu2qH2g06pwQcWz2
86JUnGuiPvt2KgE7mcU2jYLZrEyHrkup/PxVZ4armcueSNDedOkYCgvCFs+GZABX
isLruYXSRXtmfpapqZM8SWhfGpIhF00Q0kAA8dvWugA7uX0gx0TW/IA4ITCmE7h2
KyODGLD7cKQdRsgF3Wzbt8/K4E9gLLwFfsAfonTA00SiWjVPSovyK4tmsGn/9yRN
cIFrUIJI939jiXyaJAMvluStEEGadsfqLYBNcbjIxzxu9ZaTu7N6/Pne9aYuGSvr
NenZrc0UNCDUIS5b5DGNYYWUYehVBetQSp9CCzwcHbbtMdDBmBdePjPnsR7pzrdU
tBmVbUR1Fz69JEF5PYjT2QanHW/8Zd1ocBmew/qUJEeVVxUOml3OrgzQbITpRfda
Ppc3Q/WS+4X1kOBVIZCMxeY+SJaOmuMK7KdfEokyQnZ1WUiZJ0JgQaQMiJDEb4xB
l5UHhEWuSgoEdpZJNSJ3jPY/vt/e4QnrAsg3kX4bRNIaoZYZUR+kDzMpilS3uILg
XZy3aFj67KDJFZ5a5EAWU4tYJTGJlmDJO7qCuJFje0TkTU/wjXEAJoUI1m1styqO
j6/+v9kf34jBnq7v5I43QCx1tXdhwBIcZJwe/u+P/XqVVv+v69yQY85XmMrA1UdN
hJmOIN9z+PzYNhcAhIDrQccsfaOvyf8ZAi3pGho3bus0MPXw8JcBB1iludeZ7Jvj
Qu0izEZlpcEEMZPrHiX3cVA1uYymtd9GseZeftGVDkC+zggav3kjWeaFv4v72Zly
BQaJb64pDVicXAYZv6pux4N/S5QBXsHT6JQ5SQhTYJQkOFokNxKcskrWNxTVXaE/
q5EoHpdnQ0Ajjz11TAD0/zqllWYOwqaUKIUT3Unp/iqyRlzKK7UQV1zvDDsma3WK
wg4TNbRvSeHH79AsE7K5xGOazBBbKDspNJTOBV63c27qZ4YyHPrY7oT9ebn8rg1w
bx4bi2aBtMPuZkLggHZVpg7u7CZ6Sdn0HFpXU0OGx9Y8iLSokN2EsGQlR9MwCFpk
+u5z5rnlfHIYEe8P9xzvaex4xM4GN6djoN16JqQFO4gZiOjLHVRxwp69wZfkc3uF
OLEzgS10hD6GF2h6kYa+8y/U1rw3qqelIAFNebJqjc3lv1DwUJRl17KX5n/lr1cZ
4Q+7nVKBzcGCEfFQ2lOeHRJDwCd3wBmsk+sKyhzwj+RIcLJ3rl80OmDs47eb+pku
0oMCZTArDD6x/PSjiJ41kRQMVyuBZJT+tIx3x40W85//EOag+dT7K48Or4krZLXg
KqgZtj3pR834nk2iLowR9TTXCEvvf4wFDz30SysiVo420jJo5d5QNBQqg5WtnWeu
BWs41f5R/L2My/uetaywElnnXoH/AvswcALY6T/56hZmcA6cJjlI4yOjsq8bM+Qx
UJHi474aEmimzBucDt9FnHKCWiM1zWtLcSRT6KppflwEr6fjvigYRIUrmBrUsp1e
yACRCYNuDTHsCoVlIGdHi8exhCfqvoQFiLvOu2/7yk0M+2swppptQ5+xORU7r2SQ
zlqBhEmnkCcNTBLDUN3emhpDFiWwqtQf18gWI/TGXWaW9qcnn3Sv2OaBsk9nrIA0
GeR5twv8Xa+TLBjmv6/S/SF1CQ6Rn//enplRpfBmLlvJPBQ1xDDIUmASluCuTgAx
RX0riZRtXq+VY9tUDVcxIzDcAgc3/ieA+BAGWzCMyWWgqt62QUqGIgYgQT00etMt
N+JS+OK0H+uCstuQHFUux+aR4lZtZT+SrESL7fgM3GfRJV2LUYvY8t6yL1HhCr6G
YxfBz2flukIqLTHCUsJMJj/T/9IhyK+rZiUoGgflM8I/vw0xU3V75t5hm/M5EnXb
o9aNVDEmUE89/ZT6AWvx/F3oSKgwGGOW+wh+JRGuD6KXmjuFaJlG694cly390cC6
C9/CN65Zje83AmiJcBkXwqDyjiBvvoDG1Y7QMOWmy9uPcMrfKbIabykJEd2bDeq/
DO0BpHo83lWvQDdOYskrQW+X849FFGp8//SMNaWPYRPXuoF5x+NCiZgLihx0RdYi
6pcVUELA/afY95fEH02Qkmwjq2RMmtXjmvEMLZ1nlVZBkmzEJxyZwrHIGmY98wet
hvJxOdROU1Sxb+QCIRPunhiqPToqPZ9aDTsqK2xTBh+eGUM35w8DxKByi0QINNal
me0KAHoJpr5hJ9vb4l+YSLWJgOKPRQIktfmhV/y/KFcx903lzCEz5mJKVlMc7cDR
FwL0SERL5lZbdO7KbiJPIQA2lIzF2E5Ip8Nwpgbtkf4EPGl8dxWpyRWHnA77QP2x
zhz1JTix3YXbEQA3T+NpJK2/nOhUuwaD/31tpAQhgVQCNBsFEKMW+Q42554EmPSR
IIoP89ij0WO5eYx67L73ZflTLvTJjO2xboRkQqk9iiUcaFLRAghPRlWNlN3SRXU9
ndMa8kFc60n3JwXxNrVDD+D3F1tyw+FZ+UCbTrJKZivFJoQxQkxQAd+WGdDKSyx/
f+1bpzB2ApsNunXlr1UBrAzoxdeLEVNWrMxI4qQBVdca6f1rjDMcsdD6ozD+c5UJ
IU+zB2gkV4UVA6bW1ZNcGcHWz5D58ZN/w3s+FA9wP1KOi4iEkFxE2ekKrAW85tfZ
2WI5N46eIWT0H8boAQ7OOMiRDnr2oUYho79o9JKqbYJMfkiOJvSP1+pzsxL0JcHj
m7+eOlTpIG/GdlMcqt687BXQrJKZOckk3jgcdMcTU7NpSaHiNVFG+pq2EYxRvF8W
IdIxOC2CvFlXP0pkx2I/VYIXGgEWtKsiobhbYNV6m3khB5Imi/AkmLOLQnfUYu0z
Ucl6IRfxgQHJPTg/aBKldkScpPpDNdEW4jv+o09Q+MtL3kr2roCQeabPIaf40Isx
s7zpvryfPM++GHa5ACAGHTyS7hPWId5VYFmmW+2S/gIYY84fJhSWQWEIHpZRDf0D
6OfFJb9+gSgJuntwPk8VbTX6PELyYyAcWIzjWPFOEs7yhlT/o1v8WXU3jJtrhSSn
/9OmKL2hgp3EV8T01XY1/fxbra9pGffkjN4CCXUJLj99RKGfZ7g+g2mGR0PLLoq8
bqtpbG7Em1ak0/L3nv+h33AxpRGjrJ3FvQIW2ueOTtY5/TeEXm/9cXA2L+72cr3A
XGL0innLpKTP03Q4TCqznnIVSyocqusvi6jBeWDCi7Tw8NCJa57SS4gwByqERvnc
qkAKX14220DvJ5pjkpSeMfmnz7he6a5iOHnWFEGiX4dSM9V4/6EjiFCuG23HN96h
3bmkoUlGmsYylECzB2d9aKLVQbF76m8OqWOlj2fJslAEGtSXzUFaIiDcdXHPWS05
rJ3MCvd+zGY0wTUfbyCvQuN6nmMSbKzY1Qo+hiWy5n0LDfbnFM6HNqW7ifd5pYKI
vM1+uq55tcaPgV/F+ergVM/x/MRjIxlKPGjHog1TwGD1fgUPJ2Q5uLXHyul0/9xL
mt1yLHBaNT8UIIAaINoiSAQ9ru4qVDt1euc7FXISL5CIPQYP/68b2UE24gLtlMI7
+IFe1DF7cNL+yBv0pg81s8jRi+duMBCeUXhxg4t8yamSFZNMRrjzGz/noyE4SkFm
50ynCr9dOhJbr6UTJ0ZbSviaV6aCNUOT2+Q6Befq1cc8AqNdhkEw8uqMZO8PgZC0
v1Ky8zJFO7spPYcHhu/KIy+WTffO3iRA6rmMxDrdWXdjqWkS+NVamJz4hL7rLn/R
ku5VKTlRHupgiuVcRF1T7fophaYidsVA0F37ZDj+tdo5dttwW2jCnzDGSFvloQOq
65qL7yErVVGhFIxsL6RVvjO+av9GLLWKNfiKzwZcSGEla0MQG9/vJpuUYxNuoMQ6
12l5Z+d+F5zbXZaVs0TOStBGovsBsFaj82zBpEKGeCxfus5nTUL2dvGaPyZ5/R6Y
FWlV12Aw7gerzdate5h6l1Oxw+gvWBpwmcGNxb0IRjD+Ba6TtwW1qcmJkip48Oie
5zR8fTnhQ/SbxynQGyiZbFs5mqb/byRzI4LuUm+AHTq4Srqd7R5CKlLegu9ejG1J
hYaZSlzhzPQx2RNh1cPJ4o2rxKdGB+LyrG3UmtEmYal93h86TB7kzZ37CjzLYKXt
UBsKevf5PCZe9j1d7VIVuS/0p6CL0iId+TP3YUWSTb0JCSfcNnxXA6Moig85hSUl
FygSHtPfBDYKCxSSs4kqluJbpjz07HUcULu+a9Bi5RBuEdRW0wazSv+cIj95D/HT
X8EuL/SKJFs4JYCWmb7Dii6CUSVrBvS/Adls6H/4prl301R4KJawSQUofR2si9oL
52jwd8FcFlfJnf4oVNwB/RW3xVyzZrtpxDqjy6WqA+WzAylj7aHrOj59AZHbsKTq
YjQkw7yBoDtpf1CCUiURtHp/mRrF2cxs6BrG7B4fgHUSj2NNk0lMRx5qQ86HwnNg
QBdNBkgjGlFt5k7kRzCMO5iadEO1KYboXM1W6l41QYcuEUpsXhAs0zWZpsGkyy0H
LmvISxuhSOR6dFWu0qNYGG6lsix1et9wSLmGq3/YgHL7N7BJcef7UZ2SYql3vBtt
4sf061o5bHHVCepPdiqCmLNTHFXK1sNoX5+S2mJ3PXUiUduf+1kPZowg+/2/rF/a
P5tvDDMOADGr0OmsA5Wc2o2fxtxsitUEKzVNgwHVhhbXyO/LdsPWe4vDLmEznZgQ
Dd6Gvj6iPn7SaMq9Q7TjWNZ3yxqrTxrUOHuXiSJgmS8QxRLDG1ggauJGIgG3VNIS
bkSyYRgGg0UNsKLs08Wb8lv7wtkYHXDthnDUwwhhqezoBuXkl7C9NBSgR5IOqlvY
DAGiaFJT/ZsVEdrcg19cKiWM4ZMQemyG76SvlhRx04YSWZEVqloq9p5UmjoBzboc
SLin93eOCVPWAjeys8mDbC/pp/C48/LVDE/4esVPMUE2lcuNoZjaqZCN6EaEOixU
E7oaPPZQeEOBQ8XKhjLpIlgGvMWWEKB+S6zdJgeqrcD3GxJFFwxuciOooK1UXPqN
rslPLM/NGMGcxCEny6DlFftc2Ezi9TBRLojjU18b5F+xX+Zz0dHuzBy192NS7BXv
AfNRn+bZ/WOdvKR1dCeWYr9FTQoDRVaozocBGuq70oDt6vPOxzT3psF1FnRsD6cn
uBAhNlIKRhzUUZJzrSFuJTqdsjSsCm86t3N0yteq6cYupKxdisbtUPtobFeI0b+5
FhDPhAUts9ZVDwVk3gWAt804NDiqFfMZe7MMQ10URzeE3hwfc/sizyRCdVVmWlpr
m9Luty0EbXSJPqRcyI6ahADhQGY579jAc4TgqqmM/B0d8M30lUpfu15KP6sQ+sUq
RVXGAg1NL43QDAriwubl+sCntj+0AVRPRSO3lrY2KEcFeom+ieG9nPHlKCKTf4oL
tRyPCZhaC/7A5XOVF94TEt3a+Tt9RNFlTuo40gnDi7pE7UM5yJuGYnb2J64Rbucj
gDVRE68lqWL8+kq9sSc6H/qbtEZKc16N/BdsHEgLU0amGcQd2cR4mjnRcpf6Gyl2
4bnxvCo2qLMHzv1DYg/U+E1g2gJCioGt5vL7IRAaoI8geWqf29XrvgkJ+irgFBFC
gNy+zkCrX2kgYlxBe1Ew16oijjeQJyo4/GT/qguqg9OaElwJkp3hVXwSr4iE6248
IUeAV3vHU6ujxPl/dyOoGit7gq00FvQBpbtlYUJ9rr8nOpKrgxvF9+ZhfqZMxO9x
NEA1fzkYSQ0i1J3tLUGaHafnS2HR2HprcihDOofirmQwsibz+MXzGY2GbTI/JPWD
Dpm2EQXRnKiIZPHyNJLsOnMf/ncwMsqffPKvvYZ88oRzghya7hqdo9fi1qq4PclC
l+RcEFyn/04eD3fLjHUWm27rH4pMJAxYZVZCbEL4wKaQVc5mRPwn+cgBeTtLM0nP
SGAmf2WwjTw3sqCh/qYoBkL7xr4FcbA8AaJ6LINxzrSAzLMQz4IRy3sGgoaEkgcy
Hh//2IPF+9Icu1M3d0AXkwhpkNv0EdynA1HBjcN/erjAFAg5MugmyKjUJcSdDO48
wzqTTJ6q5YGdS+iu7uzxoRqM+O60oV1sa2+N+EQ1aiKwO9h3lyjrMMWO/zhMa9Vm
yKKFpFH13ofzZHzBZ9sp3tN4wXOr5zsEnK5c+ptZCY0vbeU2GpPYfwhSO02Fb5mO
pmW973wtxfdsbvbOv4G/xrY+CErD3tVv/FGtT25WAFnn9X731RGQyle51NaoP8xs
ab9PLWwbXhIOknM9iokzkRB7Ji8+pgrPCsWiX1Mhz/HavUshqx/Igfhe5V7BvzG+
mPX9I6qKLWzy59UQO2uI/v7rhUiwvQdRZOdOKfWRmABFobTyrSLrGQUezyWEoQIL
pxwDBDpBeGmFwEDkwIakzTzpwBKpYTYgsmWmJbXzey78cYD9g1WF8b6mL1KYiouK
p42VjPsfQNn73Z1jFLZyM1+JblAvpX7SLTDecroGdkN1gzWy+rZp0FT6aP/Yh2VY
tN6n6Vdr8VCWhF8ne9N3tjgPkd7jvdqieIC49CpWgeErjUF2Qm3Kzloje7psbPJQ
dqEGyG0BpizVf1MlIVNBGW6mSJv5BWBlPe/6NmT7jhKfUaxSWIXw8svGyDkMnKkh
0VCmlXFL0ZJoA8ZMDnwzLywFacC4XNVL4HBn6OobWvF7fhsbKQoetv2ieO36Dhvm
cFoDyPOYM4T8VYqRoBbOzSCKezbVVrzPzyfakqbTUj3+MBEeDmbGsaQG4/SWgXQa
66qLKE7/YycL/ol20W4OcRXhPdOe7Arplz4Z2eMoZB+2vpJ3PXBYUwNL4xt9iS3m
Ntu+NowwJv9xBmHjTiCW5QNssHveixHkgwKk7TYGZPHdmhQubbS1GX4KFhpPahhC
Wt75YtZHovhefL6zWQEUqeEK+QLC6ynixqTXiJKVdxOYDiVKEVE8IuP0Mvgh6WAA
ey8L1OX1oYVMHfm0Gqfm8RUk0YYOTc4w5fHPWdrXKWHub1usDwwPLkTXEemPrjw7
LJoGMiuhsXWtA+Gz4xWw5tKuPHQdM2uT6yYxVh9pnRqda7bof3mymjL6aFWw7jNd
0IwRIeY+AdEld7q1X+iZYQaTmJB/qQFju7eZ2QFF2K2Q/vwOCQ+PyatXcMlzWicd
A5A3ziKF0oYKVG3lyaxnxuJzgBvgzrEWVug8vgmd0Xe1+EUXRn6yIDLT/WiqvXcf
5stZCQ9i9dhzHgmv8ch1OCa/6Kv+yGpEp415Zqp1fnCLJLhTVbx66dEQIHUMqK1M
y7+QSDOKI2Q3BI5ySB7hBfeMAFPadWACmgLZ969dMawrAlmOvkIwgvnRQo3jYKBA
FIn2/Ub00yLM+ip40oSNJrEurEUxMb/eVh7BPnAapUncz8GIhk6mrLNdc/E7hINe
FFUC2l+TLfLYQ8AOHzG8XhHyKgmg638egNKfEJQcozI1dYv8TYZXXmf0U5UllkF2
Z6qL3Xz+4Nz/mWLV+PkmcG1PA2NoptDREaiIQS1unxW3VTqT9ItlHLRGFCyhJQ3N
75eJSfli5rmgOugfaD0kM/sqQC2u1y6x5j34ZVwTPz2Cmvq6Ns9GI/+WZyxHh0jk
ZP6QThS76P00D6Z4da6l2yojpWf1pqvH2ZlUsB0K30SrkZ3tuGkSb1osbpErBo+W
pX000ZcyTfIp3u7Rs3MDJxq9sqnwM/yYrqvYQH6ES1ZtSYUIccjw1VKyfC8KYtT+
zfDhxRS8SMaB6kYKnkL0blwdWVsqllYQA5X2956HuTGi/R3a7sLa/ewDClBZqmxK
l9j4JABRro5Lh/LVtSnzVNVhbCb4IHYQwGhb6iG+RtUNEfGVOpDs7H9dqwO5bSjV
Zf/7fvCo860OaDBXZOq+pJC3+90R6gYZWg3Kh8uphR578OcfcF61CBSD42BxALl/
L51g3GxGlfsn46ujgNYLKEj6j45RXCWzTuSNuMZH73qBZjL90smlhB6MqkuaztxB
b6fW/Nxw/Z63mtCt9kLVWb0iHz7KbIztzpvQP6J+FQpw3AdVR9+NA/cX7SXRR4C+
GUAc9L+ItOUdF3jau0M6PCVgM1QcROG69l67gCe2h4rqYEFOF18d/aLiDJ7fAGgI
/YDXd4HFl4j2F9zC4pPOzQ5GItpzHvz7NApvNjwTNyeVxf3uFJoCr05pMebCLQQY
/S0mv/vFl1uyoIuyUeU+1RPx3amsOszsuJe+4EuzJH+3HMo2SFim5POkusKhBg41
5zgFa/jTzjdOeOY0zas5YvXkitAtqP+wROdGeCaNr4EoUaVssnSfg5F5sTmt+/TX
yShFNZpleM49UbB8UMmXpf6PdVWNlkmyITKrz7YyrzmiKQdy7yOKp+enU4m4ilLv
bDKclo8sUqkXD5X2js1WxwRCn/vnw4/TqK6zEPWrFX3Z/+7gAJ0JvkJexWjbIZXv
jZe6HcjU091tDb6n4HyG5IOcIMm6N5+E0qZ6VMT10isnoocH16axQrK+hUPNqcO5
hsbTWdlr0kZgGrp7Oq/EBHA76/6q9m9UoEt0XbSwu3EtkOQSZWGcXD+woKdsl6yq
aWgc+5ykLpJGKekOBRLUzS2B5a6whHk+lJbhlF1wd8sbporFIeUpOR6mkSPvSHI1
DMKa2RX4TJSQrRhVGUBvqhORikXYCyJQKrQwAndMTv5qnmvOLC6VggxH+doyPg+E
gU7UXhffedlDVyHIhuf7knsfPKlvg8AOjtnGcRysovdqIk/sun8k1Iz0XqwIh66X
akgz+c+qwPdEng29zlFuH4aCSzEBS0vH8757HnpfNMzgmHB3/fsyqkacwwagOkk5
AfNQolyj5tJhoFUFqbHbnqZa3VoL4pVLc96IgUmYJvfO+oHyA9Lo6c3EDJX/L0SD
51ZAmoCp1zfMlznMByiXEi57SVD24UbqQYS4uBQEvhmZZ/5CU2NtzVa6VeARAzRv
VTfG+NjibuOmng16Pz9qwdtgyTkpfbLdmo4+4Ax5EXEsBA32MvxRG4kbMVwuTCHL
G9SDjY3qJR6Ihx9RHUD4xsZRKkRGiXOmXlH8Pj+7ROJifHq0BDszs7RUYZHTYuOA
YwM0ZWC1iqzZjoDg1MSzmwDAGqJsqc3X7YB0N6bv41bk2m1G+kfSXYkSxaLCUwiX
jrDtBWk5a66dT41yng9OhVF8ENSRcGG4LBkq2EzSGBSsfxRHpuMLNHWUH7udLBzq
H/eG8VzLXioKi/KdEm/jqUqSRR0OQWo0xBj3yH7e5bh89OGsPcZSJFLDpqXlAN8n
JTBxT8891nRPhZkP0F4MfdJbz6TlCrBpKaMoJDqu1SsiRytctE2B4+K6zZjt36Rn
dwl/VGe0pFE3olud1MJqbFuNPWHPp74jaC/FwMMTxE3G33RhgoW9hK7AkXdG8s/1
hqklvghsEruuogRGuTdHe3QFEZPah3LBONVenJ6cGUBkZ1LpgMc4AN0bQHLZOXqH
Cfoma+sOjN8lki047k3DNcgh0KHQyAwwAAMp324zTVCSXAQDhX+YzaFaVfaqYDJX
iZ2zCWoThvkqT/aX2ySf14p7Y1hUgHeUAOdbTT9hs3R7ygH4wBxhTw+N4tIqYX+l
zBNrKHG753OjlAbU+zHneAFvocQOwULjB6gnbe/E9PeU4knUlSfqaT0cOof+1pWm
rwzEslPFUdTt0eGVHqv63nD/jNIz4WrT/3GipEEB+RQtHZtZPM5tjDMws/ddGwrG
mTYjETBA3z3lPS8l6PryGk9zY8UAEaI4OABc45AW11xRQN5/KjPknLP4Rl69aYff
nDBoupakDTpzdQJscV7Qdt9OUOJVqMIoC3p8DS25Siin7Wq72aK2mncjoSSREA9A
2n9LBDowuTZTVPnUk0+9X3dW1Z2ZRreyg7Tx1b6KDIkzLjvbJcBjW8Ut3Rn0YvH/
Nsy3Q+l7tM0/N51wphR9dOvKv4gL+Vi1yxmr9T5BW4arbVo1Ebd7jCBUcV3hXAeN
/0SBIsKmCf7/1AOOCTQ7fj6Sd+kx2UKTs2lTXO/+Qn2C8pUnqZ4L6jSLym83x7sq
vSaZxpVk2x4wodiOUCMu39EwIwsY58WStAa9/pYdjOmUHK7BmBho+Gd3DUDpPG15
eSqRLEOiR+ZY0WqJur9UkoP99tvpOEvbquhdO0FNQnFrT1jDkkJV8iAOi9lo0f/C
iBaklEi7G/zCmeUSXvA03+lGqLeckkeSABXWXwUPkBICy2KGC4e3h8WgLAu9KQwA
HIuKqkNJBm3ORzyuRtIbRyysqjUfnSwWDoTyRGfIhkWASyclAsTyTbqxXTfS/jyw
zWTTZTLsep4EhWlxNI80dBur4mWpZwt+NPVoNYp2tpPteCKF1oyLRZ+/CbKALbLc
wMzdjtGVx+vbno6UVK8TkvVw8ndaRD9Da3TZGtmLLY5bA2Vs5EhSzZFFiGOhVCWf
SeJU//62wLJhf2EpkCaWQIgl3RfJQ4DcJ4lWI/chuZxoaFIsMWRgPYoA1t6raJ46
r85d1iqk09Zb9ZRNd/lykAsRro5FwIaF3tI4pxoNTW0eEdibWLRroGT+s9QTfRUX
W03mmGI+Pno5AHbTI4mUETPPiIc86ghFOsIJDTZdI5WN7NKratyeMSH58R80VRuB
Jxy/nrCnu76yz8zy92q/AkNsRf0CYiFGXZzxOXPAdGmoJKo+t7qcH6y7uSIqyA8e
559SqNXddWQP5IlY9XV4eMFo8UIYY/khLTpd0Y9zLKpBFctsArtoyoyIC/rZCGoF
xGWjBntUvAQl5Byz6+LKY9NO3MFdGVRtvMuZNlNmFaKXsOfBHtJx/cxI/uJOJ1rK
B8Mbdt14/vZ+cPPQSUUAa9SLteJg7DNg3RKii19AtVCk157cOSxBczlKzhKnETzc
+0QiAkYhhNbBCj0JOEdsfGkDe6SzIjoX3koBJYQQJKIBtFMSOmHikVbayPEqHQA/
GCzxlLCxY7Xiioy71F96qk3P7ni0I+Gx753SAwqFm6ord9HnWooUETGrPyR1fwr0
ElWqjCWfyKiaZjmX/LNRPeIK0qgmVBKJ8LWxTqmzJ6aEbI0TYSSDoEyWO1ZnDdbo
qxb8dK15Bfre2bK4fR+NjAq40A1EL+mEl6IcRJXUQq0ycE4t3ipURlU876cCYW22
8iB6wyx1aJJEIz5+unQzCrJPcXxxCkVQY/WE1+4Jpz5S8ojnWlmV1OblseY00d80
ovs8ZiJnCvVlHt/m8aSin6GZh+eG28VydDQNBPDH5JAFA763YZSr30GkNR0HSV72
hHpFYmoVNF4pgmM7jXwBRJc4xjxZihgfUXNgf5xVLuJtinIZs9M076nSWXILb78Q
Xbt/x6f409Uo2ES2Yn54WYdGzCuEkok/a3bQqc22R4nLWo8R2aUnwIFMxMc5qXwa
ReNKfIzbJbGfd8wqfy9ar74RGL6dkNG2a4GpuPN1k6UgIkXKNna6Er4UxDYkCmTS
A+5alFuqsLgpNLsLhs/vjsGNXyvNnIptVUWZGIX37hAQMbWa6EhBgACl0rbnn2ws
M6B6zfIsWfXkCyW13Y+dC4CX83AL3qiF5W5/01wRvgTCzYJjPUpX+hZelV8/+i3U
vx4aL6gNX8IjWHeMYqwnfNTP0EBPszSYJgzlsWB/dqNXccDZgLiOwwGM5XXkCkRu
lmxnXTowQaJjZNXeORHuBww/J3v0dd4StAWo6iVNb1dIbUFO9Qw1BUxmdDZpFpKE
BtcyjitlZnzyVq0ODGVdaPNXUrPU7sdyX6ukySQQ1FJBXdUw+sEa8p72XlVCBHAN
08FUEpknD32JJa4vKaNiUNO8bF+TtW93ObuB0ODkpKvjhUVtxXsJ4wzMdSqpab65
qdAW5aQIiArmvemztVlQF+y9/jdlNkBje8/fG7iEmsBKhDQ4jIsqXKcmvj4UUEto
8vk0+O+BlHI72Epf+BEKEkH/fp4xHcQ4iz04Ue/j5rA3OEKqw6rr5qMaN00PP7v0
GOMl06kaw7kQkCIIHYMlagzco2OORAtGP4jCR3nOgt+/YWkQQ1E7/ZXKeI2Qbk0T
4AWGJBF5ICNGac8k6YkgeeLS8je4E7D21sXuHe1U/Omrd//kDAYZR9xznELwEGUA
lK5iLxzsW2r2rSDKFS/wAnCd2l8GrKDdD+/0cX4qb9cWt7cKSV1kpc1R3bBOrj9f
W6Dc3/60Lkp0ie2zvsAfi8EBR3EGHPoU1TmiKOXzsaqio2kGLsxjUq37sCJzWB3r
M8wSLjxsQmERAGY4llUjgRKgNvRYVLh7KqSgbeVB9EKCH566OP1dCBiB/o4whg/U
+CLpr0tIL3haAUkKQD63ZOi2rgN4PgjPJnOcxsYxVTw6T6sv3kTR8jEeREGGQLA3
fyK2xEWUdITorxSx6BOAFR3LxhYdRhytmjhvBTQt85QyBAcqmxjNn7vF/uFLi0eb
LoFDBnpiQLkgZtta8oh74eO0ow+GbaCeK/LEsLalFuvmLG/oQgJobyyaIllSAzpk
lW9YYelWgaNEOKLupNH+7mzz3GBRpzVMKE9TaBX0UwaKnpNzcQ/SXmE9SZUyOIJL
y84Y1epbYMR9TgIxEvOaWsyHhRFxbFDHocUvN0qfc7uuiYymu0iZ04TsetHOldTT
bq9p6UZR/3I1nHpyqeSX2+GKKT9zeBkxegkR/Jr/rX8/+b0nif4oT/7h80GZrZdC
OLYVt+khhuEpFF70JlQz2SX4FfczHTK4FEJjbh8ldCzcBW76Bnxljt+N/XDLP3F+
WKyrPHilUJGxtjIl9dnZz1DZYD98co8Smjdp3BvunZDtXSDP/htgK9NOitdAqQNY
Iop7RVu6gFvpvliUtEwHljalwMdmRGPupVOInCFurmfv5PJ5Q/XQo1Bpawz3NrpA
MW/bLsduz2hbAL+1YRjrroYZjnJANfh+zyOspHGAvsoqasHrmUPF491LnOobAWHN
qxlwUlaplcAgwttz5SeMRhkcGI2Bh/XJSv5s4qT+alUtIxL+q47mAYU9ZzXWOkvW
hplVJjhXZvEqLOfDTlJuBm1GQP2pOjZENucEldQP2LCQOsyhPRqD047I5vZvpbOP
Djc92E+nnWzKTWd6YUGWB1HLegVi6qBHQ3ACq9mJ5MvH5cVFbC8f8y+5jk1Pq2B/
QLSM2g1BLjd6b1332/FbOysBljzKI3GqV7TeIHbrEt5AJ5soK8YQ8gBOthUoej8Q
ce2qPjo8JtHXqU57Sb/OA7KcO4fSi2XJyw64RJ2NI03uPkMrpp1+VHRmjFgthr47
TV7oruCXIG+HROoU9tvS4SLBpDaDZA/Owj6iHRnK+eBdjfgwEm7Nes/1XoI2gsAB
xGbLmtJjf2PBA6DxnlXoasdZMv6HMmQ+T/suTQiBOXmN/IEn2+j2GfEdrhUZWyEt
188WsO93Fy/WA9+ZZFR408DnF9dezKTW/wpt+4uACxFTAN33on969gpV4ioSR7Ps
wdXpeiXWy4J1x24FvQwwoYTWRW1mj3zsytxGGxKTPET92I2oJ1pS2aZwCqlm3z4X
PtmCq6JqEuB6V9Bt0ydDqn3pXy59IJ6vyfU9VPN5CsSUELz0/2cwFqIOBaXjzdJ9
UT+EVB0l7vJtbcvQDVASXttVOZBkW0gRqwogVHmhu43p5hiDSwft6dAarjaJF6c6
SiwBa276e7iYFU3cjXe3eESISxTERh2g8SsaZKlRkcUJ3r1nfncNgE0NqaXUAyu5
sFwJLYNtjFwHkIImzUN2cwcyWMpO2UKDFmGcFgGoLHieK2VCrbD7dt4S0YAMR+cp
EHCACqLrgV/eyQ+CEYGUgrK9ke3CwaFKBtfGyeppNO0PXBfWK4LuFXJtL/5pXqew
Zbb4WOO1/Yg+D563/nkeDxDNRW94uu8RtR2pdfTaTU63gyqnzNbay8zo89j4PFbN
yWN8LphCvhnJm9JIXtmady9uDzpRRf1LlfyLLM5B+/550bzy2JW0T3h335RC9xzO
67R+WO3Wa4XPA3MjiGiYxzbIr2Px0IprgIFmgLdm85P7buNm6BeUcKWfETJcXkZO
kfIvtNyjHnFPSdT7OwQ8+U+D1StdS1e9eHu3wSQ0GXXScbXfPRbkFYa6K+MFp5sN
mKGc1067bZzqFnP7B/oGeHpC56NLyv8/8Kd6b+JkXiviSpXhNvhbvZpGPyLLRLQW
mjf+h6I7avA+IxPI9WSI/9s5SVTnr1+ptOUrYwY+j5GMZgU4DeKqIHi+TZ+MdT2/
xeXaFI1jUJSsMO0UIB33U05RTTtyKxRHTBh8Eip9fDZ5ftkHq3nALFhDbwMQNSp/
0obftLUQUstqYnL28YoKvy/GSPvo9V+swYgEj6Z5B8lKNPqITPSFRrrSS1hh/+9e
KTFIVjnoUEVcMROYe3RYvfSqB27tzPFUJlbrOpBklYgKg34NLU131awt20hRmRCJ
Jcu4yXUxSrNrVefAmHp+wjhtpuHkmNtQPDrjpr9xqzeHH8zaa9lHySKlQJRzouJU
UVD1wbh+0E2qOL/VBV1DSlQMp6wavpe2bfTIeZ/0sxr8UFv3aY86CuEjeLZwzhEf
mIrpGr4+TVF4KE+PO+7d/6DgMhHiXP/KOFTcuYbplNsI1A4Ea92MEJq0VDuQx6rg
JBWHJZLDraUpUaPqLHowBwwz2t7xcJqo+mfW+GGf3XEC9WNsVcd/RMaNC/MiWcsz
2/I5/6dJIlmAzqXPpYHO2Y5+kwKJOrTMpnokJIlNwPTQRG2V/VJmtwzYKtT3HYkU
DcgSRkp6YNm1LyGfvkrTpC0WUOJ+Yl8HCptzrs45wR4R/6MWEBCuLlISdzdHukp3
OFr7LVla+BsmFjKH9J4FsUWkMYLF7Til0fBylxNa/WcokkFXfixik9U1yShGQ0ry
wrXFKiUTNvyDnq8yfn67JHnJFRibuUkWOg23cU35idXIhggu7XIHX3i63TyKiJ+b
/kIOwO57MG9K4xzCi/5CGJJRXs0fk2bnFDN019tudl2Kd9lib6DudbEcaRIAShmw
g6GCHILB4E1whiTMLl8Y27T8h4VKvdgHDqYBiaLSJUuH3hDmIFKBPMPFZ3r0S4yF
TqXM4pHELTLmBvSd0klLUq30tde3oZmE42O1lXqtiX81AJ2O2MXuuEnEyEQJk3Q0
oC3nKmmBxOvrAovCzFGNrg2g4QOyoiTxfGsqgDzkGyYjwHFbChRycCd65f+Dodgw
+/5nHFV4uyggNmYCRonGgf6gdoTcrvUa8fjRTM4yZPZjHcFhA8ZhJIqBypUzmNyG
jmPeMqK4VboEc6/JdLkPVf4TjJ217ae+jxdBFUsHXcHHFrcFyYzQ/0t/xAhhViK0
ESCh2tSu047BVeBXmyDBRzKA55tMAjLaaDx6OOlbOT4xIvUjN2yyjRnhZEJfHnTC
xwL2XszrO/OcMb2J/jr4/uPJ+kH5ZPYoi3hhg2Wz6hTcAqgISnW+4Y3IZgRaG9Ay
JhVFS4opU+ys6bS874F7F/wHis7ZX4fVnqMe9EGAqk3xieNV3Hhch/UGIh/rruvq
DYoDAkZCdhqMpK7lpFg4y9uWwfiXq1Gy6a93DFogHv1uFSWBJ/xOB+4WnpOFP/Se
wCdYDTmzhIr8oUpG8vZ8nxkTplh8xZ7Bum3ePrQZiCDDtz47wRfef4PsvFadOJVw
olPn+4uZjY5/3JTeEu+hHi0qOPSUzmGMvj2uG1PpxKI0KR2xxwzi9ZG+aetbCx9Y
ztJ4LHqQW4xeb847djMmOIL9yIE8FnJtkEVemM+pkJlwXkLlc+kKtzmf3d56VDat
o68cefzsCtxKB5u2OoLzQE5UKCOntDJgzbrRNyZoyC3kIqr1bpr/PVRed+/wj58i
dzXym3sX6zoEZhRuGj6EHYeGP9283eUG0KG+mQdG6Mcc4KQbSA6bPkJku5KhCksG
pGom2rW1pfjOW0OFLquS8/d/Pt3p0tPJi9b42ONfxREvZwdrg2bYRWKjZnrTUSzN
B4ighJhNoZLfkvrfiADfuN9NZoaET8p1ishWxv3ZHfLwa3jSuSKe9X5+L4DgWs2z
wftTPDU0uSnI1+FMYlk066JpbwXxhJXMYPJvJsRL/YAhuV3B/Z+/WgHxcyv7rJ4r
DFk/XmcboCYTIdR5G4Bobyl0i4zjB9ap0pexi8pZ4g4nRIoExdtVB0B1zE5B3Uoy
Clh251+ZQhGhYdUvCzzRUsN6cVh9xCKt3HszceLN0OMrr3dKF/y0zqfar9adCj6g
wGjGSa/VvGz25ENXrSycR9MXwcDNy473kxq4I1/+YYgUzdVhUON1VI029abtY3SG
nWALS4aBhOtGOuAM0ex765xH+gEn3qJrSQD8UG7UwbDtfzQb50899YFT7qtQcN27
+7KlmkAI1j2SM2CyQA49jvIPphlsP0kCRxUXL/mbcrI+KZ7icM+01pkWLWRtMQ5T
PPbJjxo3Q+bAMoGlGbkJ9JTq5+QtQ5rA7myTTIAhXi4QY+9a2j2fpnhIeGlpGxjn
33+fQDGuUFsElXIl7leV5zZt3DZARgJ7L2Kq1QIWA2rl64z6xOrcnFe0mDWI3xXB
/EORNLRi9YfN2Vf7RwuxtvARLfU+PWPvlsWYdMEZxk9DLu9BRsDMeNol71haDcdi
ymYty+WPN+cVrA3aisC7d0lo3tOo7qMDi8DYNf5bx4LqpHR114wfqiC0UYi64nIk
zjalMABthAcsMsMCYlaLEXMPIWnfjFDL+4yHn7p/QqJWQsxC9f5YLbu/cU4ae0YI
84+wwVBd8j1YSM5QEVj0RGE/gRFlF8QKRYAotGeO0ga1IwOPmn4CaugxC9oAlUUK
wviWBNs8jDXCYIu8mDRQcX3fTFMdlIb7XPG/Bl89mGA36KrxwPEpaLhTLhOQbOzu
2coiDGmUflT6EHJFpLH1cgm/u9f4Q590rgtXynLD3naLxo/yov/tiO8VwwO/6AjF
nIJ/amhyx8qQB41AySTPIzpxmZ26iUIadZvmbZfHvdtCIK9N8y/UYmt3kmvpJeMg
dyz87UV7N9CLwTPCYFXAyCXFEdVwnSYKmdcQak250n+22EMznpMsGeBF5Fk47NW4
V0MMnRAV5s2FYQtIRPi+P1zFt/vcTSXlgoPbTo/i2Y8sSbAf+KcuRizxt7dZlw7X
/4xnaN0fVnA29vUtNhXRJ4Kid41asV7DYs/OlH2Tbij908VeN6WpimBXj330YuH7
gdOycyAXOQlA0q6NLwC9P0TdSyFgSUbj1HCVGLsEMHOnS0jke8KsqiKH7RSzStfz
vWwDNYXRTiSuPK+9kxeVrgi3VqM7+uew4uRSyw1A7q4vD5/rmoO1oIkMFojrkH20
uaDSIecFhVGkeSfBbEajfcS1uiVlase8nYAoM+8+X7U17Hf9H6mVG/Dbv/0fasyZ
PGp3ItDtTGxk+cNhWYx3u5DUUw/zE2x9pOH5L4FOqzF7ExUxfWb64dWjzEmZKjE+
Cefke/vFgH31+0IugQZG51S7i+W0KQMq0CX+z/JmbxuuGeLS0E1XNTbbq1cBkFO3
FiBD6SMIUutU7N2TNj0jGRuNXaBZc6Evw1JhkJ5bdu0KFmgIcaNue2Gg1rDo2tc2
PLerthH11vOy79tHGkzgi3jR4CWaZsGDdhEHEtcHCrWb63e3xaiUTujZ7VYZhGCE
XWzfXss19ObfctCd8FEbJFYzeG/3fZOn/W2u7+qgXgUcXBScm6ZzXQ7HqbXwUwiJ
DWIOVCS1M0oZOaM9oEwGKQ+UFw4J9w7yu1GIs1y/qORcfCKCVCUXxKu8hOJ/5wzy
rkCb57FBMJrhxcTd+tBwhSPFMb9sOv4XXzN8NDPvN2WO4Bvl9Ud7xyTu6VlZuejj
8x9jk3kZBoXuUPJOTpGzeTWTk48d0yXu62mMmwc3+cXkLTbnRN0kT0PcFpmSN6wJ
cWJuiv8y2Z9ndPXls1wSHfzMp0mlgIaFw3M7vAZuzgDVPZtsXRjX02BGvucPhVTD
x2naQ637QOPK15icSblbgRkHr2iGtKmIAgEiXVjSB5kBWKWhU2dIBZhNlCcQHZmY
yzkUBw7j6Jt66433rf81fguXmrsCQxA0ZLkQwDrtA2SqD8s0M/8JSOl3NWh1eRqz
0Uwr5HDHEEyrJj8P2Hs6UzMHmU02WUzEX+ryL4M8LDOTUlTrPFXMvn1/hI243aPc
XZUMew71ZmIC/BIxZgE9fAT/R/hOxtnkFpVEZb38XL5aZ0JiGIefIO56lTxw7Xs7
JEn7uf6HZ3E/ywz1Wr3Fz0ZpqOfSAajHX78pyUCVlX0ghEcvY9T26NsdzIMz2VnY
Yn+B3OSslZHsA1tQ70d4IJx/aMLdut4PUyZ/I8zXQFTlGAA6P3VVNuaftCblgght
HewwdbgHG3uE30IvnIUGH4RKRv2V8rgWIFoqZq7gypszAtmLDz58A2BnZvzgahc6
VxWAAnR3CAQOjV3lpOwVxcJYGjayVMAjKU4V0rIK1cYzomgiPQ2EyJyGFXeL22Ub
+rt68S5FgvnzYuAmYTsJ80pThxx1SFxP9kSRs1YteEDwIvh/a6DUxMauvnImjpQu
nH/AxFdc2Cn9Bw4SpXRsOhU5Dfhwtr/GNNN5xKRgNIxGIjYNIqDmH6NdyDDM4yFr
nyvUDZhel20xrAxzjap3PllFlSdI91LKMs50PxgVSqzG35HHF+BjIl8KyHvUDrJS
ivD9az/cJ4HXTECkJFKBFpY/P8Q613Go94QV9I5ZPjmTXO2LT+hWXAspMn2qVcIJ
bbdVp1PnZ8AZ82E6oke43ONOpnVNNOJNATxA0Y8Qdu0umSA9Jn5VPjUjOpypcDdp
RVU48Qso8QD7hzR65MxvWMnm2royfriWtWfz+eNFvjDna1CUEDiglug3y4uC3nJI
wXgy54/WNprKfYnL/ilSOF11gqoSTsV6go+6iXg5lE0BRgnSvKrNIeYsFjgFarGb
fimrY3vL/+QIL9bonL5Eh+0/6I14Euqt6xhIK1sYxDSn56UieWOi3A80qLgQKVsR
ns98CgRLMf76eCLM78lXrrccA3pBh5SiGhQkKxj7mroOPNspFtvndsEiLZ8M6n94
ghVIMSsoTnm+6Wy+6tk5v1NapO3sU742p0GsfQU5uVbteV04WSeEWinXihOM0fTq
iS78UdAp5MXL7zqu3a/RJNL2oxK8lo9JMmm1zQlwMBF3KCGZGny7mWcm3ejat+89
i/quqdndEtRynU6fgVWnROQYpapDvXbixgzIA/Z2DPjlkxQDO0Rethy/0j4cLCqq
ONrzC79ThnKbKzbOIEwsmFQv0UX9ai7ae53qqSUBkUJI12tNbLaVrbTdHZQYaOHJ
QgIQi2zugXHMMeb3oYhqwHm4A7kvyCB/boGbbud03c3TEF8ZXpa9hAnMbMj5dTw7
vF/WfCT0muuugIGBouXr9t0hYJXXpkbJslOfCZ4cuB+xAFLhwtdxIlMJMJEs2Kac
6ZFJmJ+u+yP60mVy3atqjFVcyNRrAZhn/4meOPvvYp1rnHK+bQ1hYD8vcnpPmiZc
dJtJbhbkypEUnn5nT8NEIsypO7iV6utz3ZgmUiWKJ6g5/TA9feF6anmVTrqGHecm
tZf/EfKIUrKzZFZ6J/Tbyc7quRnLDtCEPDJVkIbcVHiQV40gByhmIxajRLgyqQag
rgkrJ8s7lvGDRtn6MiNzQQNl1w4m5MY6CLaLL53v5mmOY6Vu1R/HmaIBmVSR3Cyi
A/y/XEf7D+Qlq2IMqSiS8QlBvBV903BMF9WI97IORKB7Q1ESL9fDdxUsAu+5Ypjw
Jcg8cQI01aQO/PfY3rVq4Oqw7wrFPNUybO+amdteYIOl2ckcE8CvHNca8+CHnXEn
YwrYAbCX6Jkv32k9w5d3IvMW1jU4ujwb4RqGq5A30+LxXuiDMqKxRfl6DdErtkmv
NpTEzvVezP8tKd9YDkKq0W1h2FnJgC8famR3LJ38PcYMwc61zo6q9uPsMM0U4UP1
D4MvjYmI/3jKnZujjfAciAgUIskp/cmwEkOKBHyS+cUKv3JmsaoZo7w7OcO8t1lU
5wmrv4yRZnrS5oOxWEMl9dMGuxLlxbpuOGjRX1iRAXjDXxzpaE10xKLYUyvOBugs
Y1AdFc7UMqCJUwUhYbXl8ymTfyZR0lidNjOlj3ITmcedf/BInmF94M1bxDfAScXK
JJVnswjndOa/YlrJHT3TEhaye0EQF8HiQ39LKOk0IBCsxMkTYidB70YZj3JxiW7E
zeKekSds+17L/ggWYPxcBijq+uTy2HJSH8gtnkddSgJXMp619FIrAm6gXyFt/y1l
5bvPk1SqEfpBSSuSzglxhEdkBoOoS7q+KgWEFLG20YwDuNGWFc7s4QW3AkR51anS
OfR3JcRb0aGZWSKTVBqHojZPAhRNqW1LX7wIGHQX5IpXTAtqcp1r0tW1AgtagQUL
ufpyfXlmceXc6U7oqPP4KM9h/Aqf/3hvM63F+BvEMqdOeM8xetQjZ7m9lO0Mm5cp
fLgeSPTQd+hI1oixZRWfKPFYB5HRDWqFOEmhkLDNdQNbFdrijN3jMZYpkTDrYALb
iXybXQEesufZGbq59FexbAw8ONdTFC03RTdKgSg1hN2BVu3v98Cz8IoKvA/9+5zl
KSxjnGM57d+Z9ZwJalptm9H5qC3bnrkT8bLRMU/N5QcbCkeyfi9mKiErBumepQIA
Qae1Ld1H9u8eikGmldEiuYRWYZKc9sZIjArsSy8iTFurr7QYW5klDPE+kWyJhS0h
/sB2wqrHxW2qtkycAybLzyywPXunLPvVE3ynjpbjvNJaFv8w55mPAMAVEmXJWj0/
3paAth+wIiqeWqQgJ4ZQk0aCQf7o29zUR+3jOarui/A6UVm6k3DqKET7+5MuO/rL
4KUCYt4yZm2ZsmytdjKuk3/fOxj1T3/7GFIdSa8fDuta6qc8E+r4wlNqnqJMCAyN
AwMSI7s/LEy/RSgZIszTEr79ZSEfRUWA4xyQ2HP2a8jPWFQC1Y0Cgk1efFi+W/Vr
8kiK4InMTaPdl1TlGZ567q4OUR1NyYJPxFWmqx8BPo0H4jbFZfZfPMWPxuQ083kE
yyoWvlO4JSKjwD8JrMowRXnUpawb3k3oRhK7itB7Wm4AnYq3tqnrpUQ543bh8PLc
E+3hWmWXG8YLbpPhp8h85H4U0A5Vxn63OmFrc3UD3DrkwBaLIMwvd0da0GhoPWgV
lixYaZXKizol7949EosDqmDz6KCvo5lfuH2dCgRnV57RW5N1jxH8piTit1VVx6/L
RLbGy6EN4IQKiVd8TJI9r+VfKqYU9qwKZzcXHUUAhHvt4tTarNbAe20fhUYATok4
8Mg/qtnqIeR5xOA0OA7H4tFhjKFLDu2LTIzWQft7WsTZweH2BBQbN+lzb7N171Ap
i5mKVzbzhpNwhNWyES5d9dMu5BwTm0gh4O/uCtFR+q4LndEglvfUuHAng5qCj/3u
dD+S/vEJGqP+5ty0jd+1ql5Tyi3jO+tf9Wc2/7O60VKz8aSsPJfIe67rCg7sdAP6
yavm/10elJlZfazPU3Rbb1sw4HtPzjsXf6nXjcsAo8ekgs0XJa1DkMTVmHY27adV
bdtXePe/VnWGxDsk52ZqWRf4XrJ++8eni9Be3Xz5206TN9KDymgHWv0CUtJPhN9X
EdTxsZH6EptR2/pnUc796fmn/P8Tv2e+ci+cOqEUOOYJZB3TJC40VGAKKNCHEjAV
xP1ML7JG/qmlkPUy3MluUhEkXXxXfhSldtFLtKQY5zQfNbUUxT5aiOO7/Yvzgux9
ZG9kj+9TPXoIEWilzRHrG2khBvnzmsr6UPS7ins3CNm3iUIfYCCyr4vOf6Nm+KYf
yJTVwJTMNwtEJxPF0/1p5esgTi3wbrT3Vyc3QZctRQTCSQOaqzCzMKpk2biVkOuR
GesHGeNbsdXHdb0RR4XFHKxW5FBSz+p1psboRoV4hnZvxx96D/DCZ2ifS7DOnp/I
gOORs2lkeFP5EUcuruushPnycxEayvWKrnizczABQFDZC3+bF92lunmxJwjpD3b1
S9aJyearPF88WgXotRqqmxe0cMz91Mveq6D1tfRLqLUx9efMVdr7WiBHM1NJVXpd
SoaPm70vMLCicxaM7y5zIQ3BIKIlY4new6dismmd2oI3TF8lerCqEUYRoMZlChUv
36E4pOMV/zwUvOObiTcDDY2k+KFHGfKZh7oOTXQQvoou8/QXnX4MdG/MmHCYjmR2
voeb6oTtrowKPmsqwfYqdG5mYvQ4kJ46YUkK34SoSJ0xj3xiDB2CYBQd3A1Wd0c4
mUa68s5tK5xv+tgIGF9TteTIrbo3CWvMrKfripUou01btEFqp6NBXJtBD3UWtKCQ
uf+2NcYbVD3obDb5AYsh40hc/J6A1OAW9tS9xmIOaWoY5r4wqsQbCAxX/jYJ0Kvc
uodL1FZMqNqLY8p9pI8DLIRCt267Fbu7uSp2PvN+IHLe27dWHrP6fAY63Z1UXQ9o
cXUaI5JLdKo45nF1PpODtIno6ebqa7BtbHU/RB9tssmS1wRbbava9X/siGtHAO4Y
oWPvfMPxR5N62Xc9H9qxw4RdeSCetJLtuGocf5gqBhv0bCDrBW9VjXhHxxViMYF/
vK7iyp9J5fN2J2mM71n36PcJrppOrjfNtT7eL/AjR8UqDvvt3JjbjgOvUqUX6/3+
jyka2UVw9h6E2h8cpwV4cuxOeCAWZo8ySQbGiU564qt0g/5RiV8AjePsWeCkDHsI
dfHXAs+75T+Eysme8fkdqf7wN75UlWBk1iJMx/tOvnMGCyT/KPouaxN4EvoVmfQn
RA/CuI2Lwr9VsRrdtLo81TgMddpu/0K6wl89UDiD78iziLflagpy+t2adJUD6t4f
hFfaWJSzwAxVk2dr8iCnDw76e6P4aWl24SoGzWI0FEuKRdfwTYNtsQHG+4p62IeK
XWwlvJdEw0BZ6lwGFNEIByjRQ0az/fyHDMqSGqlUAIOb65J3qRp2m36q21FD4rNx
p8JLzd1h7+5OcUfTZSyRR9fmBkICPbf2QcJxS/o86zHdbnAJenPCK9JnuLEhane0
67Ryj9a1vRvNzWfdDhc/Y/ERsbNLKmQd4pBbzviNtID3x3thL4oV+P0u2ENyLQZh
VNkvvy/hy1S4g+FOPIM8e72GVIGQjQuPuWoGFayNXctkUiQaD0tuzfTS1rYQrE66
OAy31aXo9o/UPFLw2YU7VJgv8GPi1gMdmGn9eSDBiMj6bvBJlJZ6R40kmhtaVW8n
qZaCbvvDdJib/cIaD5GGXrDZIvizaEGNoQEqqh/GpIDofDpOrlY1gHNWcgp+LOiI
uKSXsNpcwQBBXj2eDVKiKqyYcP14A7b1/e9MOOLmX/V/ZbMsOnqjTwmU3UBDNvfm
OjWWJ/e/kNSyvPHRcRgWgfo+hG8AzrgKAk4mDUL5jR3jXQgPFuiKY2kl9YHprUHA
j7AKlKCcCJQGLpk+FsLaMr+9/kuNYq9gGQuKYtJ2XImCs2fZb9hCu02o5/e8V9Zp
F1Qz8MYkQyFUz/j1viKfkjEd8c6tBE4op13ANPw57SitCuH4QdI5D5Y35TBdomDr
RH8+5BHrmIiE9Hjsw0V2p95X5XHZJ/AmcKO6awOayP/gXQLJtWsinpFGjQCu6yI4
EXt3WXIAgzpDAv7kc16INq6DQKQx5sEBjaB1o9HGnJXCgeG4IsVLY/dBFxanJAp+
FHNbpFY4qXPgGJl/Wx5WheGZ2D73grWQnWTWVows4EAhXBS4tSWD4hSCFApW+EMZ
NMDOYWLOdCi4xVQASezlPe+XIEign2e2c1gqTbQa7DKpDv08FaT039IiiWoaF5JV
JZ/MnC1um+e/t3CZ7sZisJiCeVEpZsz+ZOFGesDqdnH2eWZVK5YIepKotHQYO4OJ
vz9Ttta6Cz3F3RY/RslmGNs3Sqa12aRHFfPWVqbJ+Cf8gOqEg9HdsdmMuisby4PH
+GkGBdNtIXctBCKfmriSKkwnWbh4V6zJg2LeVMDbWGkVyPZ28HXY/M2Ug7BDk9o+
wyDuzY2S302GumFH9iZUhNLlVMSbJKORhJtDvqKjIWRvqXWaGq1MQZpoNcM+e4jO
0NzKo3ztDSnjCU99uGx6J2e95sYiPtvAicZrOaB7INXxDFYuvyXIBZNhpBCnq13z
s/3+/QXi4CAwdDdgqVKJjRzmcPoSQ4W4D5kRIZq4kGywBe9Rwkn8hE8/DoGp6fWh
rL5IAUxQplrfwjjGQICbct/atopebIJCKAGEVQCVrjjlUoJ8Eajhu5F8xk9qnhPx
8ndK/PrFbfFjLTxOenfA3ZQbBKhFk1yrwHNs4Ilz8RCpfi6FqMOL0a48E6A5KBkL
RdoR5NfrYidNz7G+baFLA8lTMEZXgTpP7mBcbBZS6emIFCyR40xt2VgFrS9H5Pdr
tLV3rogj9k3ostIVg3WdnA4hGQo0+DaLHvp0aaX03+lbNb4WQgQT1svQZDDqA88A
KfU3g8lVcE5/MWeV3CtBYjl9ddhOy9vILz/fipm682dbIH8JsTfPAauSxNSB2lNj
L5qazU911pLv1OG06Iodym/zhh5A0MNE30+AP8Zxo/8UZoeCA29ZAKsopmIaYO13
E2jmI2gahTncvpcPKzX0oFYtuZkgSpdTRTpUaz9A0nRRchLI0trh/jpJop/e6Rjo
H2etNGV7KL9lMHbVBTkSc5bK7MTPVu7CeWVHeGBVs+hjyqogIQMuzZFARaKCG5KL
r6eErH8fW82A2b+5vnCD97ezS+l1+qe1m7fsk2lbVFuhnx8z8llVS/eBwNcoZnqb
MwkaLv5WPPxkp/8Eo20NFfTUiFqRMhgX8MNMaYkqm2hRveo8i3KTVm0+mg/EO4SO
fDZx599X4fBFc/LiBwVHDoFSB4WKKDHXOa7TlrJT3KMV7iN2LEia7fPzNW0L7pZW
qNcvpkhhCCBKgDeFmI9b2A917hLRKswomrXfoeVpd8oFh/EBIilxovrccibO3sJQ
XqrTYcP5Pfu5DJ5cZJ/1us5tuLTxQb5cTmuysE5OYCtHZ+rqM7iZoCP2xCRLlOiQ
t73yHBmQlCWViOdvKdWuxSO5MJVOzOn2doKoxKp/sysgQcIYu5igAreOVZrHLCNm
jyCpV6T3428pybSI9dRJCHF1h9ecjFsZxo5+QJlrPYxccaLLu15DK3l41qRoOmP3
nLm2PtDJ0kCFSZitVA8LEF4r8mTWzxgdJ9OfGQLJm8tQYVzk9qurDXMsY/4HAUbm
281z3za1AY4//liIWEybjKbZxL1QqvOl1Cyd6qL+EihDvOoznAYI42f/7NhNEfOJ
wX8dgd1hifgBpWkDQuZ4Td3OcMenHti6WDXaVVOuzKwujwtHELP3JaErn1Mj3tdd
cxUo5MYVEcrjPG83tu49c4KBl8JxWaGNZbQRTBdNZa1ryh6bpqVpPjxiYE2PX99C
Gk8C4/jNMjoqusgkCs4jOvP6DCsFj5M2iVKg1x8VMpwvNxdz5IqJlz92JdjxGuY0
8gmk2kjK4TqSqka1mnaTUGatmBMbL/u9fr223GzcPwnl3cERW2CB6A0BWGixfhxM
5taKJ9evSYerSJNA7OnMVwtTg2dX2OkNMG8DlrkU4bHfxOf0pMEq4vMHo/RXWNOr
tiIGE6QlmszdXrj2lQe8ntMtUAVi4bPtIez8YMFS8wYdR7VbRfDAzSAGh//EfcXu
6t27+LPz3Z52fRiOzKg0PiWEYEcOEKvCzhisVZUefhxcxNvx/m3oKoPQDWTmsTPJ
S6o4aN4rlxTIFd001cEUg0c0PhJXIbGWsxfj/1vwAYXkjMrSpaagBM5KvoFiOPcq
l/f4lylyTPdVAen1RSMfwkDCE0gWUcABjNCQeWUhj7Y3XldPn1elmqSKDc5noeX4
I4GIdgX5QW0bx8UH4bBfVBf/5slLJOWPmwfn/wcd2sILA08a7ZNEYL/yhA81ySzB
4hcrkJum9laAJh8HXy6ylByA4V/zsG3619FSQlwGJCm/UeYMIUZKkMS+mAn+On4z
1JaLITB58m6e34ochoV3mw+80mSOeIMK0QxS3DuLb5qgUWIQOjQ2w3nrIXNCgcxz
uKxey1+0xDQMl/ODI9JhFx3V4PmUChq5XLOjDa0M0iuLMZqMnqK42mORDXG/YarI
iSVgV72jHRL2erDBOk8dguRFvYo8wbUpmrhjSJaV7VjsyZTGDRrK8Cp6w0zd3YWD
vGcyslyKpXPCeOc3PujySZVzUx87Q704hbSbzRRu7xQTii1q7gBiqcjM4/uiciGq
hOiCE5oeYNiH6mYOa1e+q7ZqS6FEwWv5J4jT8n3FLahrEgUndGhWFPjcduaUmjRS
3V+LI2lnaUKNraQ7dlWQLkP6aArqEaKzdpm7bkvx84/WUVWVn9OkvayEbo22cIYh
LAVpZREr3R/VCZasiZmxJgz4A0CoiWUlyBGEi+pQC6vvdBF1NMjxlDcUp1BkuEYk
K6B7qzvqUwZ5tqCyz3jLM8NeJw9prqdIf2v2UylKNRjodnGzsOTBKO6W5Ovpxz+C
OKU9iDRxm//sXS4inO5z39Frq2ad9oHmnMn7PR/Iq9w5ljc7APiLJXeqFbtrkANA
lO31f0mARgJT1ycLokEwG6DfV5dR0FavN9XuWxbZclfH3uTgtHhLVEVS1kp+wcON
s3tlfLAaqrPBoTUr/Q/IQoRyqICSW1ywj6mFmlLFaAF1DB5b+xRMbYNJbdl42S/V
EW3ybSwS9Aq4AIBky+8vuwqM9Q1l70bwvqgBw1ZmX6eTSOLhDTQfMPpmUXjBw+0f
m7GRzk3eLteQGBAFsnGnlEsURw+EEt5rGP5FcWzUB7dnJPhK8QrYmsBT7VzRq4Kv
wKs455KYInyeFsWJ9ovjWTprP9gR1NwRUUqyQU77g7ry0Lxh2Udloi3Fxi4LiGXu
F1yAXwfMS6y6FdBZVirZ//s9ICSy7d0uDO5J9z00MDCOmc+uXn0GfeCLsWgL7mrk
/O1Zz59lmMGEOnpNZVwzWHB9bqdaOafsVghJinGyniBfXynd5/lakOh99LQkn5v+
5sjSbnbMfDOzYPSGaQXsA+b6dGCAOmD2Bg6Duint7J7GxGkTpnzxn5UtQQHxyCUZ
QeaoxAifqXEbBf/OOiE5KxRe3bRJ0FRB2Zf0RXg/WxWTO3+y3I8EQxRRcd9BGNvI
pV2b3pTb+XUDAY3J0r58Drd0/p3cjdRIbL/ZEdgc8Zkr4TD2Zlka0jiIzIBJslVN
HkzpwKbpftbD7+paN/gD6pN8tvhDvNedPOFwtzeW045Qup5qpPeHvGNse++tBJ0H
/x01POyBAPAzz6dpLoLtgDpwB0RjbBOeqGIzjQ8lEI1Uc0vFRgtPxt2ZGd3n6r22
F8qECwpdqgnLTvFdmwZIOV2XSCoACClBw2dorLFHVDCdYqOzldVlSgw25WSTqN9f
QIIZyOzfzjIHC61sEc6CrosSZxRiHArLGi5K9gmcZsu7KKxiWbe3jbyDFZPaBTjk
hYP9UiZvOgVAa3Aid7Yhr4799hoDDsoy8u8QcZ8wiUSIfqsMy442lGskGffM0tqi
Yi9DHcOxTTfzsVQc108SLo+9FTfYUgItmwiaRoAyIrGfLo6fo5MB2d5cIu5Vt5kB
I4ZVdkfsEUHnL9zeZlSf1m/PinQlaxq+Yef096xf1rXqfIwBL6eRlMM6SsqgTe2c
W3OLWiufZysBCpTJTtbKTYF6O6Zhu6hyyl0KqD0NfFlyy6AG50bGDb8KUwOr+hDX
6R/gfeItJvpKfR7G+7TPsVhsjTRr4vGi2zTC9xWALb6YEJfQObk5O3n0oZwdmPDt
MdwJfaw7jI2DCV2P+7mBPj55x86AdesNtkwxF4LYZf0/5oUWsAsu4d07RHPj7Avu
IkgGbWrPX1vt43cjOvhn62UC+n9meMePUleAp++pO3uDm9Q3CY+TtTUIX1z/EM07
JYjMxM7BE73EQ2py0uj//JWqwsCxRzQPQy9U9F9aJXYQix9JUlfKw87bvHwngAsI
CgtJjzgLYNEAzfoZm3jBZCDgSsu8aIE09F/zWoGueqeLWPC1C7y38qJS+3KqZ33n
y6hnQTuIdDl2gVmasKpPQKfllg/KAffYaTr4yLkBjn+FQjLXfhIIffkmrhbamRv8
mgI1352YoxA9wA2FltpBl407j16iv64fAYfZEl+kqYKy0QHOQgr/qUP27IDzlQKy
AZbKrvwBmx1Z7nfwDSSxRTs9H1O2eIwH8TjIlLOpBkH2HmmEKZSmi7fMV3SGqsVe
t5cEYxEfwrAPE7d8AJeo2J+FWJhktC352xSl4NL+rh2QTr6evIDF9xD016VjS4kw
teeLhWxsmGiqwKAgSaut49ur9OTwyE0IF/dcBxOfRls14gN0L+xvScR4F8iXhjMM
aeQI5uKsL7+1LuLpm3FNRmwWckctto+VKyWL5PVhDWGIRbjXFFxPDqC4w/xAgu2R
eSjZ6Em4RTjLAtSJP9n5xHcGo5Upf3gyFuXST9xkIlynDSQXllolxhDHG65xwJUA
xbvLzp9kbNglbuOklhMNJ9/VmFCoB6VftqoL1RY/R9y0rxzQbXlKWjVyk3UIKNTZ
7YEIyPVA2fsIosg8WnxHFFivX+cPztWHwFVIYbbcLopWAApg+NragJ6L901yEKiF
vEBXX3IHAQgEHSph/HAx3OD/ZG6K+NpHobfWowUIpPTxQQHAKI5fPAWOYdwoEniF
/1fxRSmCy1tPA/bsVrLYwpfKn8hBovcHizc4AkShKL5r5DShl+Uoiyed3qcJYlxG
r2OYSlAau1DoTJy3sA9XOa8m6znKHO3/WEckpijBQDeQ/ALtsCGz0T+8qlcdAZ0s
qPS4PuZHOXUD5rCBRRr8zF1F3zYWLe/IBX60VcYQf3SGMPGvBbiDbVNQrWh9gGpg
y7aZnAwgwto01hsnCVQFyyysT5SVffVQU8AnAz+fDLbZ/rxoSKVoU7LGOnzL4Tcr
wkR1q2Uc+KuA9ZvHa3ODYtpqVXB/JX+nUhaNNkoLhJIOfNkQX0P0RGDxIsCWq5Kt
Yqd3bsk/hA9V5C+sOq9NjETcAflMsNGku2V+wwozEBPEIdxZ0arAwH/ECJSnBUoV
7Ah8ZnPZrZUQjuWNJeERq7AgOE7H1UD1lZBM0ZuMKEJE+NaCO3f+EYTvc7L0QIGq
asNPSUxO/swiKdGM+pvTHxL/RMwAb19Yq0RFyDNOF+xkwM6+P1GjpO8PQkJFCZyi
6ORcwGZgrggjA9tfia49HlJpYZhG7tZ5556G5porpwapHj5tQ2vPplgrPxJs+HyM
nbG3ZQeLXBObJrL8aCcUdhiU5XPbCY13ciPZoO9vKEy5RwQ4Wr5zbkLO5GyGDu+f
QXRMsO8cG1a/wM+DmvvaFA4dxKCg8xapvBseihPpBP7Z7m91oBJ8MHN6uggsWfKn
mqnwyfmA1N5K/XFj9fbnEBh1VEHiGdUoqVpoNGtK8a5WHgTdDok7OZaUVwyWROjq
5Pyd1E4h/FjVFsMMBbW8RkhU7Fv9oBSLv2i3lUcKmFe9HLoP+6eIfNsvUNqxC4Tl
YPhN6hoyJG77PsrQRfsxNfI/4ReRqFzftwRzlShxrC6mwET6B14TfJhBjNlA29bc
s9ndsEgZ794TVDXnXW8GYDTpXlC4B7LK7kD5g/436PXshB6Y3vApYpHcUeMB332A
xBAGnSVtVzogkEUnvAWbFHgyKAY92ga8b+bKJr9jYDCOoodcebWrCojWT72/1CAw
i2MsLG1VlK75A8NMdHAbb3qyLMasHtoxXq5tL+jG7GgX5E1xklh11UWyL4kbDih6
Jli515vl1kVXedydxSLIg3i8/wB62+riHFZsIgq5FMKiGVuY3TaYaGjXMS/zUpMQ
QD0AWTXHISzSN2KvWBhGi9cUVIC0Jc/0wjqD3z+kuAsP9vGfTTSfgk8GiEYBHOlg
P13a3X8V5oBob+FplHoI8mFGdxKvqWPvULxcb3Nf2ddPuhx9RcHBhfkUKz85RDcE
EgPeoSU4R5FgcA3rHiJvM7ey+wwp+kxuAYGKfIu1CvsRl2XluKBP00qfo7HFhuww
FpO/9AbwYIqErue5tWEfnDPfHp3WiV3qQYaqDtwlkPRwFBbEi1S7ZlkJJ112CR6Q
vAgraplrb3TxHnO5Rk9SIItLwk/2fed3ipC7e/LCJfLGt20uN0yN3JRLQ4qYkTEg
sE+X5AFC1cb6HjlRl6aatsN/fxyg2hOTd64gvWNHSmtUUW1rL6YHo55D2+BEDOen
of5BcMY9KPCD9h6LriSM/fX6KmihNh4l6pJefIOk+2K8GCiJmIRPnoznhOW5ADem
9NDVX8j86nIGi7AVv5/+ed7doFqzMsTkcITN78PJIBHcSpepKeckAlnN9PgIh7/t
3Bhc4WKixujfAo8PZAvZOcOWoMtSbvvhsshYKtpauqhtqCoFW5YoXiQG0QWqLwwa
GUe0eh8gzLdo6OrETMFPvdjK7E3bCqKmuNVniJ0i34PTmjKlWZc7Cga7p5Qp5nw0
1QOgF+A+oi8PK8qZ4tvTNzmc3cdvwbA1tu6e2/bA4XRr04O/5t+i2PxkW98FUGek
RcsuYMgBgaGeRI/2lIn0sGA1X5nXOS1ch/t2xcPTwRNMvJ60sRHRagfnLD+T8/od
keeE+f79D9bBDxRU9MLc7FuW4uayck09AErNFmArJ0n+S24Qwf7QXLHf9S9Yq3G9
yLfruMrzQhrNf7jlXEQPYaNEyRVW7uFJsVrhXSHBn1Yc3SyxCl+/JptYfYhC1yHJ
rC8PKRsG0DvgJ0RY0AyiqXxS8TR8U3psf3/EnixIRlchdSmpV09xKvSL20AzwFyZ
Vk625JaTmoJh092kIvDYNQlmdZvzSwhY3z7kehNHXzI8bKKA44R9FejQh8idZfWY
QT6X1wuVfuUedxRl66fvupecqDpKUq1/20xQsSJRFOz1mtoBjSI3v3clPIKUK8L+
UzvCqr1v0/c1yhhSB4n6+r9UjzL9aikEvYaeHjZBPUbF7vISl9AVkecu4bPovOV7
liR3nwMe3akDZL+PFoGwT4WxCl+cfWlz/TqNpqGFO0zi6jy8XJD2gNTkrNhlumWu
VSMa68tk4wDDCdzlItMqxG6UyWQf9s05Tl9drN519ZBNL9KQ6LUq/8QCtPnLPO9n
N/7ElLJkfPbMcNWlAmbeOCODM4ishfi27Rx1QAuYxRZkFrp5tVybFrtcIKaOrw12
xgp5/IqF4TMf2CIdg88hEH87Dok2bNjlK3jgn6tA8oFvmBJ50301PwULVmY8WVAT
CsFgTfhMvyMRnvxiotwHf69miIzf37vnRh73mJ+HD3m/9Cz0opMQ5OxsYorqLYcr
GutYXR40cWoCKhCUCMaIIUdNqrk67tzNcHNmbesy3uoHSq7UHr6ue65/Q+Nu60gr
vaZ1jOby5FIGJlSTYD8uokMAfLBdOUHAz2TFn9iggdZfkSB+PAMJ+UUSMABfFm+h
uLc22EwiwIVrj3tMHyrTBBJWR5JgX1k5Dn+J9A52Q6P3VNud93wwYLhXPcBrEFBd
qY923NiZ3rCeW1t/n0fUQjaqRrqOX84IiWN2gHROsg2zyYO1ZqGBctyAc/17P1Hx
Pa6r+Lr5LXK+gJnHdsj3o78SG6TGeRN6eEeVTSsWib8yZE6RlITRIdTObWBr+us6
UvQVh6JbBsrwb12p42D4EyrAEZapLXqSt7dYqoSR9wSYCWDN3vbQZRMxg3KVXfQA
rAbyJ8Bg0YyH0l6zzsC1vZsTE5jT7rcKqWv5dkmogTttLMLRecDVGDX6ePYtPCDN
x2zxSMqWdXilSDb6kIE5M6aQkvjJ2NTg775+wLizwc8lumpyklmCMqG7eFxyniBM
X9rERn0zRwZHjGWO4kIArkpIqINMAq4umbR9YiROUK5QH9NNXzOPlbTSnPdf9wu/
uAhuwVYDSGxxQJXV3lPyJWbgRhAAml6c0qHxgSVYekFxcFwTz495P8CreZ81OgTO
x0sOsBkwg7VWaQsuS+aEgeKA3Jk2ronXNfI0T8+ZHCc9pDl/5qzPJ67IV210qv5B
izYVI8NKlHeqYmq7xwJed9dOk/Fug5+D8jokB+S9MKOMHu2T1VPe2PVKHg/98BS7
sVRxn0zq1mfYiOd9ufuFguI1uuSuvOlTaID0McbgJhO3xEVU/I7RxqVitvmDDhiG
uojqum1fL9i6RHnNp9iapAp0EUh5U/vRc+F1CsFIaOiaVWZQYjBC62dUbkEgiuZI
35Hb1kTeJsHOuY4JQoBT+2aUZhZALhLQDBJEjj5DXseBzlq1aOCptd+L8/3NRqRR
4gcMvZThBxmUh2v2xzR+yts3IUsvFf/7Qp+t4rpa9RURDfqBh46VZltHCV/tWBsu
OPvRSekYHlhfjrwmstiN4G3Rt0iBr68UETDX9FJfTHjRU0i9jrXpiC1m1s3unyds
fLifHnArK3nVUY/daUUXO0A5YqFgw755RDfwIImKEJPQ6BdxUncIIqPAQLJyZj+/
QGMZS+TcXYX9p5I8ElcywXcm8XBhmiQjBIHXEZqLNZ8cB4l9FiCbG6erhgMtThse
CR7/rRaHkzxmDhqiOKlI/VPFvqVtVCuIPd2vY/EtdMEtASnOf2hNdB8QZTtdv7XM
LXa11a2ck+UnMCGAhO/b2fr+cCTmZ/AqlwoTYgM/t/pWsob6WfO0iemKUuL07XJq
Mt3t4EPwIoPIKsVAOPrMLzcIVX5D2jfGvUlvnh5IDOQJh7M0SNweoQVBxeVrGWrx
Ujaqw+SeDfkZlRMfwhNpxXN7kCuy2vRDDgDwLDpZfSrnZnJZRK9xJmLYSDyS6gH1
lar8Z9trxehN+rpSDE+8PgF11PmoGVM43fV9Z1ARrVMaZfT1TCdcKz5WYaY9EmfG
a658lND28lF7anJUxiHe+anIKuSAXE+YNYVQpjd74IrW8vkXKt8HsnH0RgKm6Jog
pADIa2C1dp2a9qePJI5Hcc8RCk1SsUuhQPmgOjd0kCqodAjIY9D1Km0ziGVHivzc
KVo0NBmVzrq82iuDB8fiPKSl4J8VNjtsypi07JRo8zE2rZo0z2HghWQaeGeoJLqc
hYxd0K4Lwh8i/YOoX37ekxXXvfKAHR5MjMQJxgnUO0ktTvWXv535KhiudCP5JAJl
dID+6NHOoxDalCiP7MsKtB+3s7hO9HBXaXG+Jni+J8ezK9NFa4GaHqY7U9PoWMoI
9pg7usdNS3dCpEBr0yOKvrC5Glt3053snjJVvdlx/kD3rE48pU4J9HRPZ4M0UZT5
0PJIi+H7tnx90+5i4ddw1XA2kJ7AIL90iwtQDYQY8peuIZWOpYQxBFyTriN3RSWN
qj/0L+wQhLdIsqGTVnC51+4JbfqxVG1hSPba0DhT0wNbwMneC/jl2yp9zag6hwBy
C77eKTl1ai2fL+wtakfuQhjHRs6oNqGVhtdpyq3asQhoDKgPhu5hQoL0XRJXeIFN
dupGlOAMk7WTMmh6u2QRHf5Lr6buAebQ1qiGkUUGsgP8elsIe619vVwkOVIWLOkv
kgLfgf+/fEqGrMaF2ihDP3KVJ63g7pOhy1ka4uctTasEY4skKOxPjpYAJqh61atw
w05iP23yUxfWTk2I6H/WnTOvmrCdP/JFVIV7Y9MEUoaoVbbmjLL4Y1ROrchJW0Pb
6RGfMPOiyxcQ23trwVgGvPaE8sutlqXX8nqQEVLBhIxE7/YtGXAijgtNxdhrlr/e
zBXIuxz64ufJ5TkGYOwiUQhBtvHpcH5ki6vrZ+ey+09GzBpud/bNAWP3eW/P+Btg
xChVcQIho3CPX+bgh4/apI0R9OedpcV3HyauA8k4RiSDZ/9FE2t4PyLaaUjRXIF+
FqnyfwXSo5g29OQf4mtnzNKwjA/0T/xkKiwGVuQ3NyzEf1MjTvWgw+ae4BXeaevS
6/yE7sTjCUYu7nVivpJMsruQ+tpOhU6jLSdEdCfz6nWRJojkPShx6lHvWll23+Nd
EUhzHEWgGPI3tRfrgem5zL4TnPz+mdDf6Jt3q6H7/iVt6l70TfHAAaxFILRaObqz
mWvoRFcHA+s3j1+K0bduaFRYQ+FjzX4d2FbZS4zo483jW4Dn/Tyx1bmvNA4U+3Bk
1XSdbneBfZ0FtunK9yCceRpGLmTPQQtZyHqca/LBF69rxqacYDB4AIXe4/5/48+4
Wyc7SV6LGeo93vz0SaZGWEuavPhxsGjKnCxuaJ5ks6Kz3vFHtVbAOA2yxsxYX53p
T1pcd+oVB31ApJVHV1ube0ZpEdRNv6DvqnJUHVchShvymWiob3fF/YAKrHAgxo5d
qKAQ1e44XsCgzwD/wzuhFUD9wqmExOyvx+sVEvSKT9WcXL4W/63mxYGhfkupn6bD
IUnosSiuhLmxUfxDG6dwFt/jnT259Ad2hbVE9qTWHQaXcZj2KuV3De/2r52C8J8j
NdQtv77/KCpOhLGcJm+4j0nbBzAeQhHPDjCxeA5whbFxE3l5A0CXP4cs7+TosIQb
9on7BxY4nFqTIZSVpAkVVCd6IE6DeWPgpjq9OErcvnqQGSdAZP2zv3w3yLQH11P9
muqht7B2DOu75/1HH2yQaABNHgTqnlSblbpMlonoQrxUx23W3Wb1/KUr2ChQuPKD
dI+Xp2Eum5tVZ63/DCVBxqGAT4LSsf9+YUYjloTgfQzJo1Eluw0KwkR2zoEvC3QV
Y5mgM8uHSD98ND+g/zXxZMtxEFPD+rUETyBk0y16uk9zzQ5pbnSG4PNNMdtEz6Q8
IF5aq/ZqzjdBdZGf+/j1PA1gkMCaiugJ523RfLSqkux5679uZXjE5IBbcng23n24
R/wKrRLBNGTcr5KTJ3jwm9hBM7N753w6PSru+cAO+oVoMp1ZlM0JZ7UE1GT6a71X
nxE9n8wsL981xaH4eAXy/cftTorCA96v+gEGs5Ee1Ge4fbYQCF3vo62ABZ5pAUuG
EmWqmIHEjo0xZasvq1aX0XG9yCwdMxl7fpDbCwO/fuRX1TkA70tNGxbcviVfqdYs
zh2oN3fvD+wn1yCQk9vcP6Mq9eBwCLAZ6n8V4g/l06NyFkUYumWEtn91vcTQ0WQF
fDDZkfswT/+u+smkAeszS4kirgfZEadVtLHGy4h9ybIquts88PPiPM8lMg7qt8lN
fcLkQeSNmy9mO/hmbRHEV1jxadwMTMlgoB8Fh9gmWnRC5x2g+Fp0Gy5bbCSWdj4J
RYKPsYJibHDCsFSFyLEC5dNIeo/ECOaklpZQcWdDH0bg/fk0ObOKZxfGyh7B73ne
EoxzGDYj33JGecJS5ZpPu6ceAyCphUSsORjL9pxqhyRWmdHILLANGAqXtTHcCf0X
KvHDrHV/SU4HgU7pRP2jD9Aogjq58UulsYqxDJRSWdN6MD12sWyvKfTuZeI/T/ve
R52QsWV6WG1e5ZZMMQCy2eTSLInxxItbXavWge8rVA95s47imCJY1CADb/QX9iYl
AYh+8PlXnR2ZaFv0QF8KnwggZu6O7z6yJtSR9caDZ4uWsCysivGrkAmxSaUYQR2g
xS1X5ncE3dXdvQcGjiTqNVjszFMUTWlSJkrJ9cpicQKpDNNdPYdoTeAoq7p4+HBj
zi1zqSDteV0/bluupnJh8C/USWM3HAr9+YiZAbjJCII+5L7cKpGPvN+Tgz+hJc8d
K4x84rs1gnRO9Ewaif/PJ8yrGDCpwTfMVON28ccivf79CBWU6tJptqEv3WFYeckK
yqE2pcp4gdaIoDEhJPJIzGfGhact7cZ9BwRsnG+RkiXwBt6yRBy7tU/YQAbjFjps
qPsetyAtX743HGiqu8cxho6sEGgdRP282e7OtGp6jHTypzL4oqPvgXiWt5DKysJD
WmT6r/luIC+Ty3wefBJqNWLrOxx81QKsDawgViIKhb7a5k8ch4jawopIpDQIEohs
O7k3CxQ//bH42HJgp9+Xlr2o9j0ChRzluLV5BNfhlDvxTQAYyfSHv7FUFMI3+YDP
Twqmj4Vj5Lz2HxKFg7x5xQsXxSLbfQr8rgjNtUSd+sRZKXkJQcp8hxrp6TQ8iDcW
zPgbTNoAiIkZuJOi2mBMsECfvzT5I4HdnTX/GtHZEfthPf32DpozasjQ+FdLSBfi
uMNYXbAiw1fmXDDoHPCakwreOv3ckH9O+JmtGgo+/21PSbykMVRAP6gQRmeS40zT
51yTB8Yvg6uta4q0MBPN7lpEZc/UwYsopW2tkyh1olA7u/l4vzfNhhzCIBW8oQq4
Hl58ewXT/I6xkhScxq1lg6AdGQVqASKYLDbAuHXyETP6BfsjoPVa4S5OgRrOK8bq
bYfBJjORdwjvCKd5/qAkKe4nritHnsBYwAytxJWoIr5jYBEoq+OvB9gMzkt6WlDf
ystWyu+c44KtBcXQdmU56hZTZPenenT53SjoWFjGc+st6ONo1AUnN7ZRHfvqh3Un
GI79GjBlebHyVhkLMXObnGOo1y2RI4+s47aHROWcTh+wBYJ/9JAnjkSsauH9ZBr4
bAaFMhz/RlRlwDQety6CHvYeM/y22vvfFeUhxWkWBRiHbZk4svm3zCdCkqfw9OW3
KzR/j07zHu7LmDLHENDxF2CTjKRWfNDpw0tGVmpdhQL6oBqTDBxxaiEdVUb7fip+
prz4vmE5S7p/STnYjSrwinxt5k9hy1BGR3XUjLWg/Y4ZRHhGATm7LDpjLy0giI7s
jDmcrtcjf8/WZfOoJlXge6WHs52g8+NViqxtXlrCXEBZGTWIFHF2dboehNpaSK8V
TXJoYkep1HBnvD/7US/sy7llOSpFQGmhvUEaWC4d6TCNuwWGkyah+IJad9CSnWwX
A/pWNx8P3mdj28KtHf05YUk7DYoAlHfFKEi/+tCIErloQOjZMn7NuElNiEKI1MTd
uCzG9jraa3mC+gos/9lrcYNXsaWvGwSLn4jgghwA2wIt9F5aAHqVWI2gLXA5hB1S
yrzDzJXiFCL/hPgzlm8ohxsSwW0lgvuIBKOrmHNtgWv6AsuwvpXWxIcJxnD7b8xh
C+dk6k4FdU+atezMQAXzVygrw7PTgeOM8Fb5LX1DJM62g6co7UIt6Tp9nb1VECXO
2tX+y2g1TBj4ENWpLRgHzUl+RIF4joW5ARmGTMbMQhLKfGpAlrU30go44x887FW8
xreYBKxjy6iHZf9p5ss5Ulvo4o0bDEKlzXwNicZHEwSt70AEj56mnoIgrfmIZfx6
qhL9OYH3d2mpP2soyd5d3tFP8ga7KFA7MEVzpxkV/fsjt+7vGnwsFF8rQu17UV7C
41zxOFvUwykFugl6EvPl5pCjr/BuuEdpsh0x/eqIzscGNd8EfCQVvRwVVC+9ZHwH
JhATeug/TrhuDEHQz8o55LSUDGpTvzLf2ufcljuQX1g+87xjKPIOFFPSHA2I9hPK
nwX10dmLCr6VMCcQMo6SAB+dAp411qQHFc/D0HaIwjEyxEa/kyaLOXH/bDjfQ7Vs
HrwFoaEDbgLvg2Ps6+iqdrygOD2WZSILdYNmAxEs/6Z0E+JjFJxjkUIapRuKmWp1
lemrRVS2PzbnHo+YgMP94Iu4DdaAM0x34oWUFK0ZuHOyHfasP4ce+rlV/eWhMH8X
b9PwwZybuSEd0Ej2UpnwI3uCs/Fx49cJYDQmNexSJ7btLJDHGBCRPf+D2xHO9Zgd
yt2PLhxBP4eA7k1uNFYqct3WtccU8moXyk+bkoo1acz9lfqVT4Wp8VAuFXaLSCkv
JhNk/aRzhl3XEnb5UKHH/H/HqCGekZ/Fg50GX0DDa1m7NxNDX7vutSb8hVlbAU+g
/iKpv3yOjW5GY8q3EsqRO+VmSckQ1EYB+QfUx9t4kFwJqFFPsBoPC+04Fbpsz3U7
3qE9nd0KqqwPk6SlszIX1fG+TyAZy71lPMpe8VoOnsHZUnHWD6l/cXOHRmMlCrxZ
1Ce0QhaDCQ60WRiQv2a8HScagysRGOnbPBzj0mPYqU1MReDjvs94yKuTnKcUPSt+
2XGMUgAJFAJ7hjwm9kFJ4/pnCIb9wodstoTbmRFCx9PXVwHtPPJCmBToa9wvoF6v
6nNLZrwENzbECYYiTXIOhrAPLnqVUV48LsOaTbrKuJXqosT+4GQ6O8C2/F61EeGL
ishcXaZkQChlhBperK5Rm9sItYlbH14qqF34GsRA1xiHfQxKNLNiDVvT3ciHky/h
4UCYqIO7bP3U6XU0C3epvBfL+5GtxS+QM2Mk1ZR7RlnFMjJtFp4CqEKuy39EmCPM
X2Ar5XsxOYYSCovap0VBqFDQy4/zr/Z265Yw3hmZrYTLKm+3Kz0ZycAn7f/VA2jj
Qcnp43eopreddvEUcOMZqF3A5q7bF4GfO8ri8UidhfJywvprUELwsJ53XBlvC/l9
UVhDjkLQlrYM9Enz9xqpdERAtaoaiNAqwDpEPqK23Ri1X8lnUV5mlNwCEY3CTsBQ
W9ipARAA/S5VtmORcqP6rzCL2jfI9LMjli9PoSUg0JecMvvfWSwAaxaFWA3d45y1
+YUC0AxZmIiP4lodb+W0TQwW5IY2bAacSZdrHWm1o2zzCxYBGV3rrQSBdWoz4PA4
M5w+oygxPDHhxBhdujF8oQQtVTiA4ywUVIXxqi3nMFuGedvMnwLSqWLnFfKu0F4P
MclVRAm47t6q5A9O1zsHT1zJR6D2vzEG2Mst8awdw21tuKQZL9p9+Z/mE4v/+jZ8
F4ZNnqWQR/K3RZ3xiVn7QMjozh2XNp/4tT7xEHDgvtmeSaj12AyZRAUzcria5hSm
r1XFokVQALDNBUgQZ5qtfKdEt+lFadtG+rtosWtBoPxq11T77MT+Gk8HDNBVx5Y3
fu9FxMVczYNAqn4A4gtoS18CBu1x0QJ4Jho505jWYLr/2vIOaSzroUBLFP4Hio/N
Fxnb1nOzsAoMiRg2IhRqFQY+1Y0Tsy6bqP2gD5lsCmKad+4x9dBEvEx5sMrRe+LZ
giv8UQKn5w4cwEW7Zhc4aknjj0izYckiPsxhD1tlj3zGNI2WD0Gz5bGwhBsoIXGu
Ft1qNszi2RW8Z+mZgWRZc3OefY+1wO4F1pBxv7CxJWm5uKsAZEdnm7RwoemVdxkX
8BT59MJrl/L7VTqr0EYjHepYpGoCtLdKv1830JBAQ12fGPgLcFVf7a06Gnp7Hf0p
aCoRu/NzE6gz7icrbgWo5zNIuuBBxToU2S2gpB/qxxBS27mG2o/qAwGRQBSlCOzk
QO44L9wWpxCp0dN30Ht/PsXtv34G7XwIj74ohve7Pa6k8o0sczBmmpLwlTgNuJSL
kEP1pJ96Mr7V2VnidPGRaUGQDJgHJUr+wjwpcIkeqkkr1fdYJH0a2CqnAGa7utsc
WyhVevNSH0HcZeCY3uWR0HT513HGMq3E9gObgfGXI6oeBKXeFsXi75WUAOLf4SAp
h222tXoV7Sqd9bODCJqN3YJm1HtKnZ/DtBdih4vQxFKzeGrOg0SOvHX8JM+cIye9
/OX8HquLWd8Qv3xAr9QCrIqvQeFIKOCRondKyz3VFGJHGctihOr60c5u1KSko6Mb
ynVqNpKSwahpkGHd8SCPpZ5iZ71D3osZUlJmSfd9AKPttcpUTyH5oGNrrjWajFzL
qOackwdIlT/Gm3nUD/XiC7RzqvZinT9ASScDa1MS4ZQ9/kD1QCrPnn6HXgk0J8Af
PNbciJwhqyHpBKL4bpH1CfpiSc5fftXG5d7DjSdV0XcczE8krYbNr9Qsp4e0BzSt
M6YEZRB23qe4cSYiGoOfiysMbpu2l+xzwdrl9uLMkQe6/dZw6YiwXnORqflfu+hG
uumZvTalwWTTnlPfjJnM0lY+3dpdmEXHRgPpfSQvmTWAnvfibUVfBSsjxK+zLH8D
BP0Pw1YxeCZFNIdrHDmjYAZb8SZR7XfpInciCUYtdJg8HtYHTCaWURGv29bUTXDK
mRKuDKeuPtXo/HxB4y33p68hDGMjv8K+IAs9sU3cZYDIghBjQ0cX5iexdZzppdjG
UckLuVwWDO32ndhd6QTjb7HQmbpGCsDo6wkEppc53oEIJwxOz9OqZtqlUOGo/cAL
cjMXGunRpYEsznACJp+UD5WKEbiWJ/oY6p+VUH8X2q0PAMr4bhn6NI+Vskkh/aaZ
4yXjIxj/C+EegQtLD3hLfgQ9k6Bi1z/p1bAC3WWwECkr0Otjghg1UtwnFjU9WTRz
fKQJSBJhkkM5jQasUHuI2KCP7CqrOyvOR91wubLdjoZM5mjEOiGwMplixh9KTZsU
SzyS0vgIJqnJKjwwfmZqi54GGreK4skGz1FiECJ8Ks2pYzCi3E3WWpJmKXmfVZnH
+XhBOr+OGyh1MBYOBHlEon3ySQP6D0BwA1j4pencrQstskwra+ujN+sXW6VuKGGA
5/pxCD4yIN0GRm3LbceJ7Nqd1pLk/dyiq9F8LAUDXiNPnZS2MIM3Lir4nNgPBwQ+
7Jk7EpfQgZGGyvltPvKKX3+cfycXw8Gzhxpj0u/KzcuslnAV+L0+Ob6t2MEqdsk8
AvMTfg4zxzEFl+kbtoj566tyypukD+lHEFiAKeb0Qk/B0/vBjs3Gi7HYRgoA/tdq
f1+ukt16cpDLICw43GlzgKail25U+Rf5y53UKaF7TjqD8mtQtLOYPCYzAtcMoPaW
FuILd0cjB7OwneECInIWVOw2ozZd0XN9LlhG2fUPQp3ClOz+4HGuKfOeC8czARbb
m7CnGRvrxOTvBD0CheQtCP2kWBoRD4bx5akXZpucJoaaWtovsfU6Mofnk9KHHdHz
bpHlAHsM5HV1ztOB6q/Q7jWYuPwqm0lqnD1SlAugPunM4V9qvjchqI8gbOn1vz1/
TwB9+PWqCnI/70baO2wrkYaYC7x9GZp4CsqSOPM5Ko0yFUZbldH05NwX+bMXAkUs
27BmE2j2drAS7FAHiW45SfnIWmsqu5eZpQkNt59UygzUW6/WbbPgXzjRufq9bSfp
ZmvfpTgaIA1RVtYhsRrFAWaz5/1/qR3feUhASgHESGYzsaVoMsnkUSzyMmUZ5gNt
qRArPA+Nqd8RU4XzijqOa0STnEvf7f/nf7JtBrkiOCgCCElFyIAYsHXej4U+E8XQ
dbutA0bYniKa5LmCj7BIDKX1XxJeLlGxm9XBlfeCGdGaz5uGkveMQ6m/blkGLIOm
LAM4F5BkNP+qVMeCoC9jqJFuOr0j4ruM+f1Ym5z1iXWqiclSoVaEaRsmY1G6bfwM
/XDhjZaHdZ6EC+95oqJHrQybxP4s+bDvPBepVtraWGsJ41+YXdbfFhlrppb3hQ3S
uQ9KITvAhnrZunACwvwZvG+JhGQEN6MTj7cGx1YtETq30S8FWwRGP4JAg/F4zayM
QECxgTeQnn4F4wcnrNuJfaCCJ10okR0t/ZqZYY7IL2nGSlKm7XKPMDJ7GPf8p/s7
o1kDwQQxcwpp2sS072d2aBOJEgP/dniQeXsfcPiGUu28u2/iWBFzMIq9mjYYTpPi
4hmsxAAXbx5N1bfFg9d6SvIgebJVcmwtY4z7nb0ob9/6DNkfneKl4bi4BETMNhQN
/NPfrIZOa2NxLmwodHvYDaBx+90csTIjPOpdUqxfYeFYY4tbsHP5+Wowzpz6/zMN
bVNvsMykgtB+6h8MQXZcM87bL+gZQze3OugGnIpacAdfzelubvX5hNfY5UBeCNnM
SC+hglLq3x0l3uao4woYkfvvbmUJr7/e0OWQOKLgrSZqhGUDpmXFX0QuMwNWxr3r
617NTnr2C8s0CpE3lQQxLtt/FyqgvvIQDsmFFrwWl2UjMt70MT9l7rb7vWKdkJ06
Qu3/r22w522eJoY15XD46N6meU+i3rVPq8tOaKk+UvOjoZ4aZ2lm6WYJ56Wl6Djn
BUidjZLkkD+UTqvIhTaYhrt9CdC1KVWKpjRCGGGYSdRiZbITdWghVA0IywCe8w2n
NEHAJwaOispi9m7638ytH+3K45U3/nJ+tgm/agx1GUob533ZMPK02Ezd6vRmXzwB
Yzzlz9cUG9EAxaChD1H0kl5jwfHu8cu6kCJsqv+mjkgi3Jl07R5OilOuECbXKiM0
0GPQ8Pp7witQp3t6L3HqjOqY42ielUbIegxZ3hf/hnX7tYJBMicOSo/xpLkJWu+D
24yUKH1+X9NptMqXMUDwKey6KgZ0C5JjOlqg91GtR9fSyNgj34HIaxI67Xdy+JEN
MX8zhf4FmeMXg/qUqRKuuWtcWEpIDZZl8YlJ+UswgWGjBb9TAB2H9ZDxx/7j0P53
TUFq2yiESNz1rvf4G2bDS//9KpGKkvaQtLpC4SkvBixW1WGUuv9WKqmAKojwtbgN
eCNXVKlqmBouLJH7uJyMCWaPdIAh67e1P93gn1QhSeZPJCHNUG9AwgIB06OKjdjz
KJdcIGtjx5LjN5Xr8q3gFscmLcaB2xXxl9NgVVBxhHIS1zacI//TbIBGKAb9hT6Q
jYtYymaTMlmxYwcDugyZg+IN/TUUFHja3XLmt+njIFdmkH8ZC3sDBc4dSjwdvQvw
tdmGE4Th8bj+zHEDq75w7jbOdOtHqWMfFAFxyDGy4kosvSM/0RlFJPx1ksKubxco
iVLcl7kESPPS12pV4CXd6D9CX6rb7RntMGK9WfXLZ4yIEv43Ex5eGnVfL4IPlKdn
meodTZSzq6+EDofEfr4QVmeMVgAlPp24Xj8kPUaLTJRRMeWTwNEHIArkYuU0auFX
1NHipRdXD1m0gTfj+Ums0YkKmXEi6/4dtE8mfR/HrRunMpEo/Vto+aZJ3TcgulCB
HcEmL+8uSyfOGxwBryNxyVTYBTci4S6H8ZSiTM3yRZI/NOdcCPsiruWwhb5Z3P90
QRU5/n9tYEejDwVS8418kfcRhzxMI1iJ+Y5g5kWD9JsiAaiZjg0+tbs6SJ4m+eM+
ceXZi0wFpE4myV7jrjiVBqZ4Qnf5e9DXqvy6pdzJrEyQjrEGzUpWOzQDZNo9DROM
92OqF3QswQpr5CTB6B/mCaaDssWgCQKKaJB+ekVSI6BLCzKCqjqrj1o/aEDezR6a
0l5YtlkG4e+04HRZsf9cqppkx2vPqsQKpi9W/6vuUT3JDUuVFyqW3TBqUOSrXr7J
528tUeKJ2WN/qHP2VylB/j6OjPjtWdqsVNICH+IWvAEVQpavYuEpAHTyFRgQAbWS
TYvXzBmuPYZfTVGX9b3Bvz0w16wGW7nM2uW9nY+79KpqhzxVpOK7O8fWO2aUsXFh
etb+9U5mUmqOpqgqyZnKIHHKVlYSIOQRghZm4z8teGVehlcRvChb/nHj/tWueK2c
8QJAm+Sw3dZIEDqFPzj8SEPCMrduML40sQdDoEpC8zRXhqENj7i+XF37TchZVrB5
Fem8p6WEuS+UUl6ypHFjqrG9kbUNl5fiBrOQmMQGff2h/65toXnVhyTTd96P42+c
fSsm7Rf04LzYbCv1NrvbMmV9qHXuyELvr0HEc6tAh3/ko2Tf2eF242mDOvOEyeg4
YImoSL8g2rVn73LJY5yhwkQr9JFf7Sb3AfIlv4Lv3aoYVcAukbim2x7SFYb5APVN
qhf/zi5b9evvaJVanjIJ28otp0lbOT/pS+fcuQfWc5csMwfmXPvdKLUBJwzz2PDT
KuyYtOeVZPFwuxXhI+nTosnHr9i0APrsdvbcyuqg4stlS+ocmHiwifyEE1abuh9C
3QYUyt2nXVNoZraQD0NdCg+dKDKZ+bON+8fWFkSZsw1Fs5JWJDzE0erB/x/Gth62
Cxwu6M6SfIo6NjbW9L1rxVBQcWmCtDUpovFWsDO0qxU6MVrhF0so0KzgKy2T58mv
JtWaUUQsKnsRfT+HUY7vGu1CeiCxST3XdQ8k5qojBWwlpMEHPiz7O7ULTY60gi/e
qiBRB4FndR9ub9n+BpZ5lpEru0czC2dnAe2bB/0sg121VqnLa6cHoc+YaXDiS0WJ
MHJW8MY6m4DIqAo5D1YJ+vGmo5s1JIgslPKeBCzOheSNqwy1Bcv8wLVUSD+vfpUG
L1Ub//5qdjArauIekohPIfCDSA8YZDrp88127hQNFU5tc3gY68pCYtBgGKxn1xy/
z8bhh/eHN4jw7qdMu25/7zUu0zCSSeyUcUhrzosD4E49e0mbviQclfAQX7EVOguW
cwfrFY79Mav+IDQZk1wdu19ZDPbgoTpslCxeVdGkMeseXndF95ZePxK9onurolg1
+7VqMAC9itf0vnh4XuK8BG38ZNakj9en/uRNLnbid8umXsMt3UGgIZAmlaY2jjzm
TTtdZqGV6L9VUZjSqIcoZb8ZPInmREv6zccYdg03sYg6B3W7USXEKBCK+65Ar8A6
+0ew+0enDmPuAsWHhTWJNCwoqV63cF/qX8yCLWSvXdru8Bai4Dxn90bxDqob6jC4
4Cxg2SA2K/8oWFi3a3zGnk2IEhmdam7mv07QBWOPzPLH68zCW17CsGCiWf8WziGF
f/hIZRogQjHpGEt1zFNNWMJLUm3pNK5BWm5rTIur2JyES3DDVzvOs4eE8XS8bEx5
wtzRz3Y9GSA1iDGy1oCNC0/7FUMrcG48DokR/Rc6h1f+ItuK8eT+33wNDRveWmSV
c7ErVgn0ifA9ED9L41iP3RkviUAKjbiLxrPyNCQ7p1pC0EOYfb80OBFiZ4is+ynV
LAM0qE03vqfpD8CaIWwn0NVU5zoOnNyE/5LFswEqFHATIHDVC9cFE62dJ/peBg4e
ztRA87/uAX+uuyqY8V7Q2h/y2Qux6hgX49XFki0nVp/AQerGE9RmjGbV3uZugDSk
n+IOlI9NiknnQbFYFjaHAkCDpcEFTprKWKCp3LOvWzJcL020DNtIaQD5FGu3Gcoa
i3X7HRiaDmxK/kHkYr0eXGogmfYQA7JNQMXMK2HuGk+cJHJI9yCdOEO5jMkE+/2x
2kwfW++8Dhv2x2QDRvLztsmc1BV1QYSWPX8f0IqtYoFDv9kfW3Zd6l8AodGaAiBS
Yc0MWgf4JNKbJ/p7pcJvy9yX8hzPZF3QlUgiGZC8URSu+P3/RxJ997eSBJm75oqq
qWNRYN8WrC26UqRjvml/25zlb/C2brCLTvj2tJnAcsl4tfnRO8Vf+s6vj9SR4di1
/+8LpBaWtf+WvBpHuan/GFE/Ln8lRuZHo3JwL7Tet2GUKrmh2arWQhrFGPj9A4+6
wgoO4kd6phRY2F9F4RJJH6fznljDRwUw6KpahhsF4QSvPwCauWcnahv9QKVUYSft
0tzpvxGsNq+cLYV6Mw/qDN6nux8cvZEDkMPffRCB2qy58vYy7cRziv1bvje4ckW+
Ttb5Nfdp0rCHqez3NWO8Z5Wj4jKtgWuNZ77ddVIULsb1uoh7112YD6GMy2B8XDo5
e5VPZ3fT2sXH5Yl2hKbN9KiXC6D3z8+DPzOPC6mli9Chc1u5YNO22k2puU829IC/
u/SoE2DAWYa9AnZDMAYKvwle6N2RBmYqBFe/n1W38fd+G3/Stljv+rVoqcNISvI9
wFGQ+X8sUxQ4xGnVKGuZdcKpX9EuReGTF/gL67fQ9+KtBhjELPNI/N62vt8x84Q3
C5+a3sjS8/MUjmatvadW2bvM65MSxRM9qD8050ZWJXJs2dbPDoy1FZz3A1AZXKu1
HHY9VajTyKajJS4Gr988qeZsRX5UUWXpJFIEwCd9+7mxp5UVdno+INjrzP5p9VVu
uDBTABS5+WuJ8Rs7OS50exGkeyAf7Exe+OUtxH1c8R1xuyX5bH+T85MTE0g5On2P
cUV15Id/KInZ8MYf2gu7ms8UsNX6SiWHlcVZo5IeERulPQjwLWkPZAVk4fidd9a8
/tYUKg0CdDQUmyyx7lFoZf7/GAHs+Nalm6t3tej7nTOXlSha9zBx+M7wTtESBLR8
zSW4YFPkM82ohGwfCa+6A23305K3RxNGvhq0hGv5BuUglAUjYK8LXC2irsP+TETL
lnbGQGL8d+s0aF5dwLpNinaNZofeAVwJbo0JGYsmXVDtCbN5Bdg2I+W2J33ZOkr4
utxu6DosgB68zamWuuW9njWE0pqZP9r6xjhqwyt+/dJLC9myBoeheW5/s4c7gU5p
yjmbiPcnEOiPWGYVnqNBN44ACQ/bpeoGI9Kc95vqgzQVusQZL9IXZLQlypzNt41u
drLmw7Mh5ALsTIK6688/NLTXWOiI4Wq9TlxsyqMMA5wKzgyXbjr0HDp0MYx0F2Ij
r6EDhkLcLMtds/JhaTiym/d6e8QcyMyEQ99d57tOWuKuDriIWbHXboGjdwQRhAgJ
UQvmPztnyeFbabaScoih48npRq9qHp/TrS/usyPpNzgCmb5iRg8AqnaL5amPpp2n
X8HH8HRdEPpjxQT1C5C5BLuQkBzKy2vX83isy/kkmUu7TeDvwkpY4ZoL/9qB9pRB
beVQbVaU1BubtH73x6OR2I6+fkxT89RUNApL6W2U8nUo055JkeVOJ1jiAtbNECDe
2eu8Y4+vfX4o7C+Tjr5ZtIYrWsoFtgXYHERulqzCw7HF3gUWbjQ8lY9D5SMTLsl/
AXZzWsfsODmQ5Sq/7M4SNq+HUcHQIoEFHQRyg4fHCtCWTR9Dj8cWwLpBWpGJrB12
fx/13TIsNPHFu5YB6bzQz3QEyGRrd0/tFiwyA9NRTI1LEbJNEiv5+4kMkvLJsOOC
I1bos+LvQ5h4oTVe8L56hYKaQV3HlBY0Ny56jlqCZFroOvgW2mDok8kMmQk3fEs+
aDIzwOvLD/3ewCjz+E2OnKRJ2ID9yKff88bm99SbCae3H86IXn5fvgIGaL5QsoGu
U5pV0htAwNWmcMu3kB7bCbkrzMCXPWGvWVkKORIu30AlXaqdfgLspFodJJE1HHbk
GcEiUg/KZvAOYT6mua2tAf4W/Qb4JzJ3bOTVGjRpRYyF1oG1IgpLYTVXWe5gSD6y
KE8/zCxHDQ9tymnnRp8SyXI+QwDp2zdPf6KgMqMIxKGUrgqfJNTaomQbqgspk4My
TdVj4TIXnsy2fF0rt9vgDzLyPrSX/y2zzcigsbiuJ5dGxVWYIzg/3JST2vGlPZFx
hKq1TfN9t89ZXxQr3tIbpapg6rxFhCZwDr1TeUU8WFd59EAl8Yw/EtSRTrBdeKtU
Io9uQOZIYgMIypHStUKQO72nN88syCy2logGl+P1frss+cB7To4UTa5i5ydkXI9k
edGZ3YlTnA2OPfTckD1pwg5HKFxHtKTIelJ1cvSCrXmWSMYPZKPxTnU5KIVoRgTr
nlxu8cHuZkDYfqvvis0Jnn+N2T7EoJib5dC4lx2m1llfyupdflszFK+4IOSWbUHh
/jtZah7UPTiIJj6ziJurBgamEih0Sgs32B4SscwlL+RiB0MhU/2kWJNIdxPUfMgF
G3zzlBSTkQb8V7w0SeaOFgfka/leqnPbTBAo6fXdxbHCagpBS3bd72goHAgjqFEv
gaaYv6u8Qr9hCcvGFK2U7YZhhhUi2ZEj04/caLYLbNUFQmrUvYSlLyOkH8XaGPcy
A4UjGsASlgYkxthM4mi8U1qp+cPiIkTX/aEOHcO3eQc8YRI+BmcGmYLNDdjaSO2m
RL1HXXgBgZJnJ3Rohuv+39X4xAVFfJtMTiVIHCIY1LjvIfE8MXEnSHtHsrfu8ega
YCxx5jIwZsCS13sKeGZPDGfDPdFlVVBFMPJ5ulJqemmcevXIlFTVdp+s90dzAlia
tgWSgR6AzCytDaulLE+Hdb+yk+Y6tHaHOB/5/N9HgKhLVPUWKxCEaE7PkLBIEGdw
82Wl11UtdkAFsVVKeUuZ+2xCqxcvTC3U0uPHsbWWLEKOD7DBayQi2k7XX6eB54RS
0l/3PeIiaH+rpc36GKSB70tDQSOqbL/5o7xtf4ZdhLzQX9xQNrxDF7Zd5ePHErmS
wiK2+PdTBgIS218hM5J91iW+7zZNW54lXkyErqaaYXOHrmW5VXb1CNyNf6rTs6IC
dLdfUkP9/Sy1WmVj720PYwgH/OgSE2JNZBwytdzdrIEEpwTj3B4OnQ2PQ25knoXF
4DriiAeeG2tRGNoLSpvhOsYyYsSgyv7HmbPLaTUsYnpwnJkRyyUf0UHq3c01JP6u
niCS6OcVpdETrovn3cX9X2SEFGyADqNbFK7AMTXW/uy6xOlhtCkHRGlJFjJtJbxZ
DTGR6fHSso0x8PMm6G2k6t68yD6raC8FgG1ZAoDbJyqJ66oym4OPyPB723FCDd/O
N8Wa8MXz46YdTxbHR2xzlqvTzZ1IXzew0BpIE5kpXs6YBT3VZolYF/PiKlXefuSU
HuNNx3gVL8XPKLstJ0Vk77jW8krHV7VlBVRJcfo/PGLBMoZ8Xfyw0G2CBP2YAXL9
LUDLZurNeL7r72mL5B93dByeJSzIjRD9WkFqaa+OUJgLqoHrEUYmvwX9eJK5LmiX
WsQeOawAT5E8tqfU1edn50AkV9icsA0NPihEsxPdNGpyokoxovG51SUxm9ofor7W
SHl0Qus72iCT4ebJ01uFe6FWGT7YwN3QdbOl9DDlWKmpJWhAv1ngM+AUW0UQ1gop
wWEyol1MrKko/ux2B6NytOMmW8T9stNJEZCMPioh7MgcXeV84bekrlU6XSGV73DS
iMYsiLQsFb/xQHKBShLROOjaCPonvj9OQqh8K0eb2QoDXCl91ff2OiecfkUBpmbt
8VweP/rDVfhRSVozLNbeni4WyuolFygRkZ1LhCquJUhfrdPotd8/sZt/J2F0gFiY
ovtdWT7cgrJfz0OkS5iFwuGAny8F1K4YpAXhlRQTuxS6+EN8JCidMcNH3grGRmz4
tkyjhBI3Bt5WbGwTyRbMPJHPuehLUZ9zCTxqdGLKLZCxi8Z9ECjxh1GlfzCzBhUg
xZVtdLL1T6eUH8t7acqXM7DpfFRWOkYyI+e6ogmnkmTMsf2KHdIeRzD0kTZf5oOd
rhZtZ9qzrcL9v2KEFtf1gHM2QkkP5/Tvl1XkFR6GMXxNLlnM9WRaVoDQEAVoRHEf
VXNG6l5mEtCg5mM4PeoqBU32M0v1elMM5k72Pg8TlL5B9vv+43a6UeqK5boUd8B8
+YMI2aZnQcRvdAHxOO4ZIvF6HmV9YX52Hp/CASPVcD6JsS8A/xu4Rb9AkWoA7Aou
OdNlgr8MkNWIdkI+HdbgXjvoqrr6Em2f4jvkNdkdtPnC0WE/j+2PMjX/Cx3KKVrN
6qeLTFc/OLrvFTl5TVg9zkyif7CNvBYQqQj4Zq2elCCjP2ShfGpERFqBgkisFD1j
DqbV6hAF3cWvUWtj3U3GJgAbGi34wmfXvHXhYUxhkR3yH/ne5hKdv3H46xpSUIe4
lu9f8ztEYIi+AC2zi8ogB0N5yoTAe8ItNJepn8H3J3JJhQPw8Fm4mK5TafR/6NbM
SAxQRSMIeJ7opJ936eVeBPWMhm93qJgtQSybYOAuM7+zJbP/Crx+YsEZVX+S3pdl
C5bnI0saL8tiHAkRsTuMCTBh6IPU0em6bCWOlguKPfBBe0wrie5+PphIRAB6Nwhc
5nwDS9tbCaouSzMvXbAnRq8ouD6ZN7DADsKk4UwWIFf6RiRJOgXftoGq+z1gQ0oq
nAYLaC37LQSdHRYs1zB2I97pnOntsE1mfiMUjrH0wv9CeZstW61E26AqVprbkg8o
zZdScDSNhzEoW69/QK4wDHFxemuRTPEMYrodw6FF4nNPYnvY4o4LLQZBM7PW/mpT
Zbe/fwut2jYlWGicXQ5mPWvGwg+BUe8vC5gsRCGyU+5iTrD98m7bKCk1/ay4iNVs
7aIkkXeti/ziXpJRx7agULVCTcQQtkUnJdv0NJiJZvDn7TE70SXZiamwZcMtqekF
9wqf2kjLDw3BGlFE3M7U3PTjRAaBbKJMyYcA+Qi/PM6mybPSwYRHet+iXXTZsUTz
ZRAXGifpPCZiG8SYVO6TmNx2GqW2su20T6jEFgBexSDZueiCZuDqEpoMoc7Vfx9C
2wsKy2ptY+bI6jLSJGC6BP7osGi9YqT35fqt25h+Rrb1UCT+nEb61L8rCiQuFcXE
EDgPgcHKYzuiwdKyDTOYTZZf3YTBbynOjkEBwftV0OWWo4+v2m0vTroUsUIpJJ22
rhA/1q+1q8hd1X3weVgpfsvmAf1Dtq/qCK+97OA0UtWsRH/tHKFeUz11lqKmqvde
itvA/UWFG7dyylo14Rzerx8usojkLaYf2ViFEt+v5JAbloGFeIqcPy3wQ9h/Pdql
2Sj3LG4mtA2RPVM9owl2XOxyRw0merUMYK4l3zK4cQYlLKIAmhkofTMA3kkJITSu
O7KgHHkzke1Kcj6SdXEGYnYPV2g5xL5XHk2eZjxxI3/EV01+Ui4bQeQFIUfGGhyU
hu4U0jvFbXioqMAWCAYNRHpjZPc2MC/rCHJcIO741juMimpXuKOy8h1pZQQP2IID
L7rR/hbAwT9n6ml/0+Njx+LE+M4MICdL1pXLklx+hoE7fIi+f6/xypt4NB6U8wfG
B17tEuH8HRdJWhtxWXXjcnNlzImUIsmE+RGNkJ36S14zb1SZvE6AizW1rsluPmzU
oGBvuaupZBjuO1rzZBboKbHfNODmTXJ5TZdEahCSNt61GCAW8HPLba0LCQc+jwnE
/65j4M1lksvLaWjnIjpwHmVq1RwjN8EFr2BKwQWYQLi8tzS7KroDh4p5wS5y8zAB
wLrvx4wMRji1+wosCDeEKccIzJU1GeB9EH987dq3pigWXMqEXUQJbfKIX3QmF4Bw
9hjDPYih+2tHU/pD8PK+yA8oTH9hiCdIO5h4uCjOndjKqQ9rnljCIU9o6Z+Juigl
/QKt46mAPfsSSL58hrp049sn1I3gmri2QOTZMkklVvmkUXRoZVou4nPALK+/tQxA
ZS6AbWl1gENogFIIB3hEYt0CCb5sc4x5iIQf0qKpqMURj6r7ZMStTWuBET349SXo
L+yYpvQXZKdxN4zm1q8+NvSNppEQgRu/gc0RXe9KiGz969bHqmUDd8ctfZIqz7Hy
3ERhQrGQXJCycfKTuoRVt64tny94anzCb3RJpjgiGvmKJr2VyfGKIntx0z0GcP1P
5KQMqmXZE+9S/WGtZMPuDsCYOAbt5AJIiv2EpoFa0xlFlLP2tqSr6jp8kpDikSdK
5oWTRGqGxJDWHDaEIuu7hHUjNQCCRztJF73avbH9dfISmjlpQxsiqloiC7W6mahJ
HQ2IzzXWhPMQTISewf+1yyCEmSrrEmezpcf24GREq+q1PoG0ryQlSD4+qqT2hbnW
tbChhmNj9GFznBfR+c/eL5KxCI6UCCMK8mXdsueXpVrUkgbctsPa2wS/B5PZNVN2
rbUGod0YQAOGVgvkk7cK6BLVlbkam/zRTvBc2eTFV3Fkj13LHGMSnBaRL98pjOwS
xtGEa1PSh+czBy6W9P0HE4Jaxx0qHKOFgU+hoCRiDGUE/wKrFgNAgUckAiPs/MOR
JeqWI4WUy0EsaMkGNF7ika4cczB96VYJV79NTbQiR15NhGsHjHXPrTBBCH7xD5wD
oYIB1fMTNdAlZoZ4Acblehpve+ZqCecve68Vp+DTuU+lth4WK10PWB6YDTAFlVEX
rimb0dT1PA3UiqXkojWuAOub7osUjjMd/3jKEeT3GJtFbKBz3Cq/TvT9N2AZlTRF
3ypn8a/ZQpgZZH7H20RqSkNLN2vZb2dvHrpXNPGiVrYoeJDgVXkYl3HfI5mI1tne
Auy8JUDEA+PPLDSDwF+xPyHhhmCVfasSVRPm8/C92IJZu0csNT6DL1+ISdbNoUce
cZ8XghKiGpSJYTy1lZxYYE7XvRHyjJI6qGaFwvySMjXvAkiqXOfVoUlWybkiFEd1
D46X9suFooETTBYPnTzrUFgKJmkLPRZhRW258yIgCjJZ7k4/jEcqQP68It/rVFiL
GuUWDwLD/xZKcUPOSF08y6DdIeiajKKyDVoQOuRYhDT0IygArWTPSbKsJm2tGCCD
AibDvCBqgpYf/yIRLV8fQe6PbsTQNWgroCB3cK4gRxA5hdNJtgT5cNCosK9tapM7
MdbI6dGuYp1GuY6gPQ5faDXsXBl+U8h9L3Y6JALJBju+g9aFk/6L59CdQExlCqG8
Q/wWaz2Krhnjk0FUy29Wvy0gXrjidmI53Mft4L5rFQ9I4/Zd7pZMgBC50DpseE9K
ARw5JPhjhN6nZZkrAHia1I8PHeQbIJP7Ru6qv/nkBXLxD7Baz0Q58sB4/bEnJISs
6J8BZ84tjEk+sbILHXbcDWJP818zOcfmC9b1kqQUAAOe10Orbs9Qm1MhAM3pXEtX
BJh7ggmV2rNXIJLujpKaurV6jopPBRTjwmkmLqVVDh151mG7PeMvT3K5jNdViT9/
8RqB0WSAH1/Ph79cp6i8o6L37TbyBVTtzqbIyZDq0VndKD3cqMgR2GdUUcts/L0L
D/C/SRpI+UD3dEeQglLmp0qTfcjPa+unLydXJ0B7OVKBtWA/Z4isX1wudzQ7LZP8
Aa0eGHUx3TDXRjYTpxgHoslbMKbq9Fqkx41c8KMiFUGe9SbevY6htKAow0yONSK0
fyLKVmvrNSli6654NTVBvXuRgM4XpIXU3pzoDSkZN6DumL6cRirG+iQLcXyXn9TM
N17D5vrx4V5FzfSXjZndN26SKVHzV/0Ss0YYoK1Lu59HxToVNWCK09j7deCwib5F
vYt7lgagdpbZ1nLcykruLTqoCavQX18S1FiB9tF0swVY8Rx0c5MrQCXVLyJIoFy+
cXu8qsilvO1qcM1iDYNOktVmYS4mLZjXjEc84sndAGnA5nhqurbpn4/sx8Gorj2G
zWuYvZ4aBxzlhprVePeh3e+F1maHwzbuoxt4yzu9lD8F+oc/wJl2kubyPbQJfS68
LZNyU2zYCAoc4RdWRMQTyLVKEXKM8/mmlRyQ1Wx5YdRq0WeLgbsjEDAmyZRjyvC5
UlGjbfVpwzKkNvRc5IGillSsRIuMGjyMbZ2GPNWAXkZUhdIMxP+5MGqjbmywxdRm
aSI2kmYk2mZQEGbj6JWzuT+RetmSCXBOh3ZVYVUxVnuMbMwoYPa6gobqG8g137GE
AMjISGylOFAA5Z2IHkxwfx7iAam096HBbJEfkK2XhUDBNjSO05D4M34vfWUvBrx6
5nwyZIUxCzIT7E/MBRs1LWfI3CUi2Ex2+g1Yape5xlnXMNuVpywVLBV7PI2FEa9N
pvtBR4kjFg4Y9kTbrCyMI5O7ByGkSdOY4VX0TY6PGLZr0Od8hUXFsMOtLoB2WP9O
ih6VXUYFfQDNAPMNxFB8l0vsdeQU4mJi8RdfIlrMJRSSsJcWAvxzhzUo/89paTJW
vy8ByITtsUAOKPkK0U5aec2pfImCcRkurryA8pM+LirltnKB5sli+po8PV2wb1ny
5hK6MR5etEMEZfOw3m5vQZiWJo1287HmAHTpQJqmyCMlarAZK21vXMZORztZ1zEB
cOrvsjoHJq0qCzCOLveMobV7UFQEmuhiirkNGjgymRMG2+L8M28eCfI7xoc4GDS0
jxInjQ1HAben/ZPgPXijOJsXHcGVeJ5B6vhuqOOOfhAaY9ALFOTvTgkWnpwZondq
iHIfukrpmams8yvOAcs6y2HO9i/0V5JhaBfmb/3nfOFahfNngoWj1/GpSY24kC76
sAeggMuRHt5oM8i2OzBjg5gg79tjyjmyj5WDb5tcVvx8DiyJ49vinboM3P/HvZR1
Tj6ZQbtNT1cqIoNKJn2FhnJ1RQcDZWg8xVvr/fI4+9fh9t7sfo0Nr0n6NMalhzUf
+3RCIEu8RoGbogoPqE/uk+7wqxOMCluuseJciV9H522PdT4VTBBWPXVvCUjHukOo
a2I7GBDIfFU73TBoftWUXm+XnWNey1sIlJ6BIsDrX2feyzrcROURajx79Qs+GO7O
IFT3X0/faJ02KvbGGIdxjIAO23LJXlYYNdAG0vfVoMWD+OdPD+8bEtyJ/SS/dV9f
7hD0p5qYk0hBN4vuRjaIpvPcnznLlO4xYbrrxbjDBJW2Fuw3uisNa3zX1pnvtkuy
AYAGTROAmBiKtU7YTxR40bqCaDcLeNSb4Otg39rBxDgywI+MojJajfQEgjmeg2eW
sEWygwTuvMbhxZaDE72VGEkv9/Nb2btPtGY5PQySVyHH2A5Sq14EgQ77ha3f68G4
NEIygUKNaZ0PAAeUpLxToK9vL1B5nM/hwOTU3uGkdMS3mMj1qeXwPven4v9AoBPv
tGbMlZwIJC1N7XBnyBMlrFttxDb+RFiRJGJOOjpBET9S1NUdAQlfCVDORjmHVZgK
JUfGK5z4dT1bxikUamv65WktcljOG5ANkKN3LS3eOUSiBwvx1aV+3AHYNqlVy0KH
XoTgWL+l6L2QhBpQ0uBuijBI8+Vym0NYdN9AZMIMpcWXo/OjFmggltJ/pkZeg7hV
O28o/fXA7MpoKKwaGS6WWUGoGwCFgSzhPOfWfU9TQ2URjaR/Hyy/gUvgMx6DSUzd
4qSq5mrHb+fGi5bNEs/CFqmoV/6EDYq/NYf6vQcUAmxx1GMw/dZ81q5WiJjxgQNz
EYxghC0A/eBUrfZkS1j4ghIGqa1OCcZBoD8CtUQM0FbqjID3NOB6pcZSpC8lhLwY
neNkv9j+VypI/QxhxGfuyx7oqwiTRFRQXGhINxWs5Y9bbzux9xxXD2Z4t9YfriC5
Mb1rEaOX+4N6yh8tMpAXafQ9Sgj+EvB7gBUC4gCki0ilgaXoA/pbWmvwUkAjh7wS
fyWZzOIP7LmHsfaYn21MDaAiMCc06OFAe/WqhsZKGOJx1+PvDnyxuoU1p9XSh08D
a7MJ6aRmaHBL45kuQrYmlwi8P/lk7QZkvxqhDza+/+dOgEmdkaQgr8xMKs2ZdC1Y
puRt+hfNeYjcRhMf2CFkB3V08y0qPD7slC8BYtynk3XTN103JJQ86UYGlXbApHdJ
42Ls7f5D3hBKNSWJTqNct5JPBO2Bmc/baQOGdBN6klxLtTqjFvI/nWSil5zt2uzA
ZybPVrGYsECkfK3pKNJq35lnFaTkcIGC/aNwqkdrI05qonPKmXLnlh7BvhQJOP6I
vunUG3BomG6AFISES6MAlm2WcDdwdEZZtkLLTefg2ZPOCakQuRgYLA/E8aTcoL8G
kh+GMRhmgnuSuLpMAw8SXwsajwc3218+4uF8v9RF0b3VpCNhhaVuUuRWEzodde5y
m58CUr6/k7ebqtlejikfsnczGhFgAq/sEBtHAci7QAHy3X7ZIuv5dGyLtfh+KGW2
ivEG80MA7nMUNW/Yvk/EZ1CmoPbeFVTi1vk5atLuB+T7c4hY0LLtlnlJ171zhFZq
eWIZczyiyyH2U9yhmTIfrh2lcPPQIRc3tt614W2HQLItjer92YxpgQAD1JzQLCqN
u/snlMwxyzOTAODrr/yKqPLOWaLV9npaGklO+leCnkrX30Q4aUiYuDm2LTYVqrcd
2ABibfbJsLpytgLYltQdefRoh7UstPk0miNrTEwuHBqHeS/IJ24yvQ0+ajU9o4Da
bZNu1sSIQDsjuucU1tEbiWUEVK3lKXdySlw/lI+RaZqMxD4fyS9a/vGX62HHTD5B
9vNZgNwyGfq3YR7fuXQ/LrqiK2kiOD4C87mYS433wN7J7SU3xfUJctPlk0AWQzjI
tn7ewXou+okuTRhTnk8fn2kJTOCqzZrUDvx+sBDQ1cGK5w/U7EcMDi3lgY99SP58
B0KYX+WWsrdSEcofgPSNE44E5z7WFydIwddnDpJm2cLDCPoUNL53kcW6+Haj+qHm
R2qC3KyyAa3BBVBR0tjX9alNJYQki2QABwK4Xrwb2BPKJcdiATtBr5PHl+eofJtm
s1m51nWXdRlG2cWEoWVB6BG9BCtMQN3PZKbdXxaDZxMOCSV0Dpqu5q+MY9K1wvrE
noa8eroKqJy4nYCJVRs6Ir+vb9bA4QVcM7YnXJAZLgvj/L7+WwclFRBRz4e3F/6j
fpLreUECu5kFD7wzTu3Cly5gIF5qgfWL1wzz1F1Jc9JlqMGSIsQrZuxjVjFd33Yi
qpr/m7EVX1crBduvXXCPrq55t7wSiq6tecN3iObwW7HyeLc2MQd6OFrZu9RG/deB
xnHAU8xgT+v97Ws9HuvIfKgF6Aghtp34O1b9gHvpIkuzgFyXVsbZ3jcz5Tp8iwzG
WIlLJ2G9YrcYpCCM6eMqUlSTds1pWJ1qPsLrrLlnnWtY7VYjGnpFK4eIYpmqPjDS
Ej5B3ubrM0VNOkR3EMviQAGTrOJ5gH++U/WWE4FzmU7TkCm2oFlepeCQwwVO5oLr
DnCFehDcHsQfAgJ5uzXzBk6o3pC+nxLhqiKG+Yo2hvrpWhxZDO/MDbG1rLuKnYWD
SkpgiEo1m/UXMyy6rgxo5HLoeqaTX2xepjymkYdBDJ3kjiDFeCFvCIgCwfatxlBw
kVYWBSR9KjXf0AyQIZybG/sMsiXcejCwO3DufAWp5cWNwhOiO7Qf7QSHUkEEAJ5O
NGvx41myuwi/TAWoy/5LrUSB9YPpUdZD3arIEaqwGJRikgTshVlqVkPPJb82SdyO
/GCLdW9FkqLLrIjBhF6ywoenfT6UPXY6pTFuZD274hnktktkp2jPNXndZJPXmH52
12KFHE/NvynexJIUXY164AMmllb6oiSwnK9hn/mLTFZJnnfZlE3Gpu6etO1k6eqc
6ejBzEra8vA6kQy8xVX85qeJ3jxdgJP51e4KmMXjBWoe4W/ZNKCHzPJMcgtQ/izY
8aqy5CCkO4/+ovhl4eKRuUW2BaDU6YmNNt33KfugamBCfQqQR1A/P/c5aNNMK0KG
fCuuIcdjDctTfTEQyjwA2hufj2HUtfJELrzWzn5K+krdfr+w5gmmE8AYtnwqWZb5
FlPHOPPNsnoFKo77dYczT3+6ryiIk4N5jk294RNcGpaNcUqsSZmwOBnwqhTsNb21
7xJHVvHzf+uB7onqkBEVbalS4cZFdjv6KZxdPD4qxQb3v5fO52QEa7KyXbWBjbDi
WjER57n6wVvQnvsrA5WK5MZROk5WD4QouEDERlxr/QdsjCGWWlKqe3rhGzzSTWQu
9020I5VNLcpjrmIOxSJJ4ntiN/y9Fza3ImwXz/ZVv03XlQqNAvVScKu6dBy16UNq
1vbhlnLcXxf0nayHNLXPHshHPH40h+w/67ecGHJCP89cCmVnsbjXpRZd5lMSBLtw
PUITXoGeDuBqgTT+GM8Y/MRhMesluR904LX3ZeFkPHlNx+Xj1ZU2nMn3kaJOowe8
OjU/tgEe8X7or6uttyQ8Jg8lOuBflGnvnkCV4LD/V40KXNKkjR8WvAv6cLmsv+p/
PIJcWV5fawx58DZGDOV+WduDqWeO/YHSlMkxx3E4yLBP05xORzRLFQ2YSAp8/3A8
Ay6xRc92SwaKXdTQiDdI1/G39KIB7DfmE7+HINGljwa+/YG9TI7Ub2ZeWEu694n0
Mxn4qWZEo812KUDVLpe9W8RNJsQZp9ga1MdvnJpPc2sGAIqDj2DWjE/k41ej2QIV
CREt6bKxI/0K+IvwwfWfkJusw2hNjpLBrijbbGrCZl/lbXO5ex04s1neC/e8V9n6
Rxxhxvq81+TBrOqpwW8a5sCl/a/1EamxX/KVYPRiQ7QszpN/JZR82XwPew4Avq6a
8SQkcjILM92IYgQrzYtbEKMGz2LnmWclO6Zv77Y2vK1eed+eOuHuu3ZYrDSVNTFr
ceGmNy0cuim8OeGLqqVQLSkPngle6ak3+KONcjg6+mJQZtUvgIG2tdbBzZmeEO8i
foL1+xna19owXHdEAShxq/avEadTTqocy65rG7yauSkK2b3Q6U3IoK8LVFlCqDMq
oyivXU7pXJEWeX49dh1wdBKb6hi6CF4CdSTeHhJGm70npnAPu6jYEdHV35jVEMc9
b1qdJvF9sh1jME65X9KP8VcAG+80U5WHLZw8l3MSmUA+R9bjHN8Sykk4dFv4vmPW
hu9cvN242qBlTsWo49/uPQ+GxKGBwjo1I2wj1fK35/az23Ywoh5A9/jm0FpMKFtq
+u/T76WmkrRsitkFxZSULpyQy+5FORCekNz+PrnqGvugHwLfXB4kmCSEVPcRtBKC
C2YDDtGLdvhhN1tZCyzkosqfLxwxHi3d92LCb71qKlibuF7M9iiDpkXKHTYZZytd
dkgsn4R9H4EzXgaBpkN008b4O21D/Pb2vgvlKDq5vZLuT2nPrM9JRPjEi0/iHQZf
AQrc2Khs86J+9DUfTuyaErhLz21zOXZL6x6rH7R3eht4G5bDVVhcVKOkAEOU8BPx
gSw5j1rT8hQGkWcv2SKpkvFNwQaAaYQBBROBF08XxPjZ4BKUyLt/DGiO0BcftzTR
G4p03l44uhjScuVLFmdC2SNEWeqQPWAckIrk+hldjSv/CT+m8KpVU+bTE1KphkGi
iEzaM658CsA+cVsSb4UAW3VN5SHnxBjT2XOAh+mv+y7AVQsEOuh+U3ZATNKLxoe5
kAuOcfpbGe1V+atTI/4f+T9xy4D8xb1rJRcAtA2s/8EHM3j9cp6eHq0jUV3eEK6U
kgN9Uciqla520Io2NTi4CH/FuU18HDxFH9nLxZnw/3K59nnnbDI8pQ1kcLe3YGll
c192drmkliajGw7AbP8O2904kRsrngJ/d2kXH7fGXfxg7QsuqMrDM4NuJ6Kfy5B6
LqAqTuUyDp3gSYU2CS/S1bQOR1otX/DmFYSZxbVhBPaJXmp9EoI6GDuUtljbtrW1
kVgHwI+gzl93zyqoavUbSG2R36uo39IhN62q8WGIFkTRVKHF8qUh4+gqsZVe7w7p
yY53mS6ZaiSICAIXaAjn5/4PWb/rHpIXDIqeI/Lb4l0ADopkdEp+U/wq/SESLYJF
vbVFG8i8u3SieqR5lMCeuXfOsL5QOryNZ22uQji9glmaErJKkkSKj/9Wr27h+Gh5
nZIHNZ0vET7BYoU6AcKVQ6Qlvl734VOHXjrspt0QemCy/xDPCf6+7x8XiaQgoaQ2
/vbOb95rVOoRONpMc+UeoxPzV+9TrJUcxCLPqpQxRKrBqdlx7FwAvyFwLLF3ChBK
6uO536zGfIhjyU/aWw0I13zDRnVF1/ydm3Jeboh8UeApp+2Gg5Pg78pqdYTbL99s
pklG3Jt1wJmJJiPCVzvQ0MGYIES1k62OYs+8F/EAPUYew7DV+mWP3MUASaVS2211
4zfMkA77Fi3Qd3LbS0qvfnR9zVjizRfxuivXbQRTGS41i34wmIzZfU5NpX5OUwSP
8R/eE+hASHcPjOH8x168l4B0YXoh3wuNL2YTnpjzGu0WpO49OzwF1k8JuzvzPz6A
rntNNZrNBKu2YBQCH7ziHKtHUuoffVu44+1Rq7RaQ/not6ta17jVDqi/97XvUARp
oV52WIT78H7ij8swRMYiSOoVnOJSACQAmZ2EJFPgVTMUWJ7kQVV33kJy0skddnsI
S7TP+ms/jUzlbMD76siiiI7IqVnwjfCz5I8qvt8dncYljIl9iLwqVVYwZpeF3Nyf
UFZt+5LX29ahnSthErbcOCtc7nolHU4ks0mhbHjAPVG0mlvvJ54W1rfF+teADpeJ
KQV95NTE3gBX0pToMrjeDmT04PGJIth6akX1D++GJXKz3yWy4CH3JJkbRLqIG17Y
Ro0FdRMvLc7sDrYyN51P+fjLDO/Rq6NedmNRrFP9lWgPDcfbbEZ6T620oNBS2Mre
9/ovwcbUn/tSYs4WKghmvZbE3YFg7B/2uiYJd0A/6nhCVRDjT/QUM5TXcW2h8CBq
1h+fGFNB3MQcQShH/H5sxxtb6wAItF/O851fzVpYoHS4Cs5g6KT2gj6FfAr3wSnz
1Spm+7oUXApY0J2/VoMupP1V3MGHik9oRLdwTGSYArzGg3w60nsdn31avE5/iR+D
aofSH5QnO9a3biPPelNVbEzB0R6gDoOI8WLazY6TZmQNtmQDVADqZ48+zUTn9/Na
tdsBcXHO+SfuGQ6goPUs0Gg1OfpXd0H167ec9Pofh3gO2QOVd7jN5O5m0VICq66p
b4CSAXUE518c63Fc7isCx0Rq0tw3KdYqAuJSZ/S5c3HT6JJzhXoGbdDmqHoTh4LI
YXlywQ4jpNLDjzNbjIkhv8gZ+KiW9BB8lND8RejyQGJ2R/L2+nXo3JOHAi893TY2
rozNUdmtviZdQBk64GBdNz/NJTc0caWSQMvthiaaqS2PCdeB1+N6wepEnagrR3LE
zV0NjMFqqFFB1DNTzjSY586RGQo1UkbV0OyucjthVerkTzmU8rl5N9DFGLpz2EW1
fApAU3IR0ZE7M3dfUZnZtR0CdL4JixjddpE4or3fqCYK3ZM/saYzuyBYdWsMaw5N
u17XmTUsfvy3ldvuk+ipaHl5bTghnwulEqrRyxw+h+2wZOWVkxEutfpmKV3HRpA7
CyvMYYtf4GteGo1KKe4NjugLjRwqjXudhwiFw5E7tzhT0zpueprPMsEdxCSOftQq
5Q3wcCx55r8s/coF9xPqA1G4iSHW38DNj/9+zvN7W7VEHFFIvURysJ/NvZLQwxhL
zDZGraOVcNltSlhv3L75E8N7fn3/NdshjyMjx1O0JAxE8FDWrGp/126ZgdRJ6nSH
Y1EQ0VpDZNSZrbbcoBTrHkjl0mti8ovcNJZLqjl0xjnJi+jKEzbNIwdWpWoh7KYW
S0JpMJgc8Upol8HDZG9J3nK+cdgv8Vk+fi5bDCBk4CWixBGSFzQ84D+L7ndext7H
BiK0W/VIOMApMcejW1gMdr3R65YFQLJOQ8nlnO9Ikt91QrdMoPqKcd/mcYwNd7/Q
Ir1+6yqpBEknRTvJ6eONefCTH9RNZemRjksiXh4SJC0NEZKYOdnr9DRfHdHd3Z9s
leyxc6/mWXwo3zNaTByxA6QjWMjBPpa5ocmEIaWZpr8Uh7RiLL0D1kaHCwyxUAj5
kUqlHgV4jDt9QfxCNFfnMTnzO2wx2uu2ltu7Y1mgHcybhv8YBsoJ0AaABX8wSTsz
rOC/YDNegOiwTuSVeDHJm37cFpyqTOz1HRG1iv6bJQhDF3bgxaoaDyCGprnnvDYo
zfbzh5Knjz/yOnN/LwQp2Aakwd6z0BkvnHRJG5f2VncHSl8NAspNOp59dHX6ctbE
rPEzkCEjB7QnuVursq9vgy9qLSBtYdSKUqB/7Fty5uHYb2rExMmHVRe2V9WCQbjQ
rbUceO5KcazbrMQnCth9+984P4pbb2OyaJBE7JTIQ5EtCT8Al8OF/sqcms6nYwHE
wO6Inoyl2yzDcNKm0Ko22D3n/VaRe0kD/mNkzKPtcKrHyGbzVbH5twLiJznMNDch
wTZwyNLIgEAHSrjYbWCkz2auykw9fp4FkEDd9rcqMKEyPEfuIljGF3ni2EpS7z5F
EGiZiOMkFVEkeBqpxXpn2FD5pNyGqxXYaK53ycwDSy6AOjFWIe5ty3c4ZV+0JF0i
O2I0ZrRdQDku0menN4+YCS+lRuN9sp+LLyaCMoKY5kRERL+A+X0qmNwHK9EE4SQ+
wEu1MFXF9qX8Lqnu447rM+iBTbx9Yzlu/Q/8WA+SqGMomkTV9tCvU68JkTV/S5iE
4Vl1W3jc2L6EAsw0BCJkrbmZWO4LnWEHzpAS2CpoPzrEsmF2jKnYYy4q98F+1yS7
ht1WQFRFlKgLOLq2TWuQYtFM9hbAUgR3p9UgK7Luqlmq2L0+HPLIrA08yURZCj7I
VDV2SIIe2tJUWq2t//6og4wFH3R3z7iBkOUE4v/yZJ4kKBMz09iXKfPD7TUf1SJm
AHTezdYQJ+FPnMJGcRUn9UTtHiOv8iYFor6GRGujjFw5REzqzg4e2EUCyCx9gTJi
RZ3Mi2Ddy8cFWhr8RxA5dMiioGAxCcuzoCLDQH0yogEU2YyG6WcOGP/kNmXw1AYI
acClzFoi3YgToxXW+BQdAdHWl0l4dOVAwRFrolUbBiDoTPvn9OAH7EgETqcecgrD
96X2KTs0GwzKoafogtLMR9IJaB0TUOVrm7RARMNxAPJgtbeea+gQ9z4Sn2X9c9pK
1qha7AzBTkKjPNrw9WJg1ypHoAjZKgwNxuqR3i8eHNXPsJyzqTvXDUx/eLhDYtkv
5jQZeJvShXtXVmm7pr0EYqBNMP1AZsjRsCCz65HNbEB+rylzM05+iG4ZggwgO8XQ
CXjmgszyZ19nrtNYpMQUCwYga3qN9LbuEsv65mUqbB+HGBO+GU0n71Vxn69e/GxH
fHlwCci6mRekLbZpig5SvMQ5F52YdgJr0AWoDFxqpgCqyNlyrl1x/XbvIl0qSKVd
N6YXAFc0qapsZPr1hsEyL9hnuP0K1yuQYHVWNoHi09ynQVA9hM1n6VFwMch5upK4
LP4uFOhRsQo2ztoZmTVPPA9l2Z/D8mERhfkg/smvhUSscjEie1qrjkgFrCS5X7lI
Cn+Bs9R96qhfTXoAWfiC/dBnv5tNDGFbRswAQELPmYYB/VIlt6X3Q3gohBjgnSz+
/i1nNkNV1na1woH3MwvwTvEkDHFCUm+3eCXp0FzVStoFFpTrdLsbDISf2bokU0Sp
uKS5BVQksJtYL3NsZjNyPndcT6VU2Civ/IDNBeHumX68xeYDII5QCPpd5ErvZUwx
PvOnwb+FSevK+YS+Qr0A+HJ243r3PKi2HF6su151lLvSbE+wTWyMeYCJ9LiGveSa
B6LF7mJS+Z6bCpF7P44CtN5LfauWowxpMO6uyJX5Tfk6h4zf3MCneibD/jXyqpie
DQkRHKSqOSBnHg6myND999iDVqyjHGmFIoYnsB9nA5Z2FaGHnW9TH2ZFOgFEEi4H
QmQpaYH48lqd1yp0C2Q+8CgYnMc7M+4nEexiBOkjePErvYbIpRDGXsYNW72mP1OP
oqVaufe+L5aGg+mCeFO/NLEokAItdmNm4ZQi0fBDAYq/R1HwgsC6TBKb9N4HC22y
DqZGZcoPi1ffc3WuPNJgAAolPbGb+y/4pSac55oyAOcfobt9hBg1VJoOgfjV5CM6
+9MbrA03LQvcjQuFvsWvT6AKcmybfwruGHCl06KY6mSO8nPry6rcOebnFIMvwfkN
dy+1WQYNKofIZe7PagPDde+XAEIFYzaXnlh8PocUYaXzXYer6Ns3TFSQDRpIaobb
jUAJWRaEx7AJyoGAAtSHw5KSODSb2khw3J2vfafWMyreueyRAUbxb+itrw03bCM7
K9A4+ktXic/GdHoG86x0cnr3n0FDLXNZhJobR326WKLqFYLb7VLlZqSxuEWsH6x3
rljKE4OtlUltLq7q+g/WKysyKFy+2mSaE8YWDApoGXRN2/loWc6oCiFMjwccEnE4
+KigVhvVZuz4/QIPQ+aZwp8boOUSGhhJOQvrfxuaNxLes2/VjpccRF0w0Ge9rK1C
zMzT7EeXIUXGf2caYnLtDtVe++/l28BW7qNmLN5+aVm7rAhsgTODFYAMErl6JUmq
6oRdtdSOrAnn7dKjV6SOulJ1/pcMDUxDo8pJMQSIUS94pX4Q8N1ZYpSTANlVpH08
AOtSd8A2Tt3rbAC27uSsTHHnyv6HToukVammKeyJSkxH7C8WyLqNviTw/ylxtMnE
V71+moStyYswnpvhNaXb489US0bKVsZFTriYop+gmkTiwyutC2aNO0RjNxv83swx
zYocBRTH//YWPN+7waO0qE+fStY1Cwv/AatuKTrt6PJwMOIBiOe5i8+nGzEgy5q9
6utszVyfwfNuMmGnulXC0SdXKgdfhFg6232yaZ7oIy5LK+dqNpZD7ZEN4t99Y9AQ
SsmJIacFyqtkcQ+22eVUI/L4fvuTGV4dowl8BJbs2iErc1bBKEQxitJuWySemEPk
vdTGlOjrsWA5Odl8Sol72eKjHTpct2mfmHCT3vrUnk305LaEmVobb9A+qYT8jbxl
nUj/SB5cfmw/rpOT/44aP5asp7MFoq2IdMZ1JBypXZfgE9p5Bt6evO9pOtrUfD0m
QBOzNlsJUzx7cAOCsLWZIJ6b76xD64KrtpStkOJYBOLWlFl5V0ugZue0XykgZzxA
vVldNi3AZvUH5Q3qlHOPCNJdvB5A7SKxvvTaVsGzzxuznKemuOt6LUr52GosnzKe
xUy2Pc70GOJkfBBZWwnDn48tVqikZNdJWB3qgRlWehLWrtfLCuHcUAh9CjG1taiL
cmknGE381I1bKfPxNrYw0kOAYsA/1OJJ+Bk4gdvP3nk+1dOhCc47CBD0Q+x9ZcAZ
OpRm85nVBhZqVYjeSIjE668F7bJ4fSh+vBg6Ng72opZFmPGH1oyQDKRDWmD8MgDC
/tEcSqQ6Bi7Lor6Vdb2yEAdpxqF1MGDPNvv0D6Z1YeW6u6JwJvt9dt9S5/3/NaYc
LhKcG4wYKAyQ+uuo2iUt4fey1pIsQCbrUBYlQV9ZZ4m9wXvhtYZpVNYkcKtHe+2i
LapH1iNNQFKRXQ9ya45wVjRV7TY7qlSzV3h+PIONkriIojw8NUUyq60yUFqRQuhM
ty4lkW2RdT1//rH8y9DcBcE6qdDaRiD6mh2T7nGaw3GeDf5o7tGtoK3NxzLwLYiF
tu8BSg/ADFCzFzmkxgkWCec4lp+WT6GuR9+Z6HZdoVaLHcdItRpUX+4FOcBSyjKb
MFKS3TAvF5yMSg4hHnf2CvbXyiDhTp6doNL0SjIbeYwPHbKCKyK0b/KnK8U3bSJV
BNIMPmBUeyi3o0ggvOJQm/7+wJkdQJHo1phaNwFGhlVrXL7xYetV+irIrRjGN3yG
ht5D19w6vw0hTnxp0P+FjvR+mpqcs4zEYphxzx2l+lzWx+wJcBlikIs+WRyWv4TF
NwCKTXTQe+vq+dd7KOjifMm5vOQnHfCsVZwRutYdjTUzePE9ZSUPZfDZMnQp94zl
temcby0psPTboQ0JGeXdbvt65FPRY3QOnlZ/L3clAWRyPb2pqBMRFRgLquOVQRF9
6ftJCpTGDK+dnAIY8x9tH4RLiWEjNM4q/G659XmuWL+AFAw3qCb9qRqAr5nEG8AE
dgBCP9irUZ2zUJ7OIMTQ3rKVzlDVni+cwzklkTqe6jrO42qUTJM4/AxyRadWbMyR
rWzJYwSuSln+rX02IGcYzpwKorucILz1Zx5OXce7mLkvSRMD3L8FVO64V08JT4YN
9i4qgE91o1TfcMpsawGpMwTewSUWHO3Vi7JSE5OShf8JnVnLvEXk4squi9nBSYVu
915J4jQwEOdMcgTl6TfJsu8WLQ/Dz4X4v6KuSabGqVB8MsIzwIUdX4DMkmaRQQVK
2K2GXyrWa2m8BjxxjS8hDZsJGkg3jEiMH0DZTy471R8PYK6OAyxG4d9mbqAa6iju
7R0CYwAnSXv5XW3lXRWnkAeSTe41aIAJtNIl+2fXIN1wnqKyRp0Y/AhuU+GnxnkC
o9is5myLHiNhLEITyavhiqOzkpK1yr/DENFT8NxBWpzgnxXZLJ4IFv8wRkwLshUu
FBDDSnQBd4syepUFlNgzlqg/zvS3hsMYzQgqW6figEPpEwQ1LkuhwP72dfb6ZRGV
WApvG5HukAiDwHZnhqInnlHhBFEGtsEzNqF8FhLmX1G3LzBvwbPbxpUU+afS9BNM
9fYQLHop+xklulf+9j4auTkdpCRkBrfJkiVJRwACbQo2SPSqzLiV1Yf/SCB+3zjr
5Wb7DjJ/7rsd8LAT6DZiVcgmk6Sws9cjjrEByc48xsO3YcUGMl4ZNmtAsXNJeJ1w
j+qgxzPdrCgCYLuYngeQPcNwDtfoo856LxEZocj9hdn6ienjoQhXtJHxBTxKGS12
IQeRvmvvIraLRM+xTvbMQTrZbI3v9t7OYuWDo3mRCr1u6us9RQozvR/Gq0Q5K7vp
VJGLFlpPX3CiCzHvOy6DhdDN2pL2bUnUBTWZVadFxroMAZiUTnliFIRBqLofY5pJ
K71FDyy4TfUCr+JMB/hCPasttqZ5VMAXV6K8Ctx8Iq+boHNNAh4H54h7Pj2QdP9N
bapaKJhcEEW4yVKazI50J18Vl93Gr0Cc30lshKNBtS/ayIdIQ9E6XrgC+YRLuJ0E
lzhRXf1S65tpUn9zH2vbaUSLCo9LWnh87+8opK3okGAunjpDsbvKk7JXPIMVzn72
L8eK1hps0SvKw7/Rp+ukX6db1hTqVo+4Q/pDHSrclGHXAcV9YdhEkNlM9FD3ioWK
KlGUhNWVa2K37TO34c/cD/X5j1MjaerLjyEI+NmOM3ypKBqrhd1B2zmUIRE2HjMP
GjpMuf8kdIv/yod4zUmySxnu42mR7UUGQjZZpmYULq9rD9eGFvrSHGChOMmbz4Ns
suZky/ah457ko4UiXbnk9kPfVHzZds2KKFG/VS4s5rHxesYK8pJyrkBOzDdhIZkX
Ql8lORFYLR05+Tij2d3wMLCMA/znOlZhO9qU+kJjElScyrfeBMs+TjImTUk87shr
A1rskO/4iFgDXBOVKCDz3Hvp8UPaX069xL/ZeoJMdVVio+vNiPeAYNK3k4BoKFsE
iXO2Z362RzXvwC7MAqEOf+cEO22UE6eXbfBzorKNGG2uE9EgJtBEQ103bS49vZM1
TqnfI+e0K+y1Wt+0NyQJ2zT7h3PQRr3FAsvcnRg8XZa5m0yRrSZKv1Z1kh5ctOKo
CBD7wqR0p7JPa65dHGvmdQPpnExCi2JMkzdv3+xDGzWuPql41ZEJHmfFp4PKeGkl
TY1vD9/x/u27EAouCkYDprtNpAC7+67uXOpns8IdoV9xqmUgWWnRnbX9b6WgpGDE
a4FTZAERF+t2GKJSa1XtaXj/5SBaOzJre0msg9w5MiLpvB8fJ7+bdnvwXEu+R7zO
O7oVg1VGZohnBsPoNucgVtB7pLkHNuhy5IAVU2yNArRrC1R7Apxboos2KKTnQx11
n7S3i5IAVFQYmRVxO43wpv5eLB9pcfRQaeDNwbAOtVaPiORyQPyFd+uCWQ6vGGxq
LTdsy81QMw8aeQ7CXUD4u99+7v+zcK7woFnjw8FXnsIyPw0dVkbxSF7WOJXyW8mX
E6wUVmxGMFledDL7FQ67yiaLBq5Iajic8utKE33vxhqN1EvoQfgYMZsYADtOjdfQ
vbzAYViywVcsixUHtCI0m/p5Hbufxthmg5aZzjhLGkTeqEeCwhGj/kJDHRQuQ8sR
+MxOOJKBWsQdmlTbmojyKEbMPum1dGhW5ql8/gCflXHW5/re0Lz7T5ZMbbTBOlqg
OE7omxhDbxDlo5fPEEnv18AwFsLvt/dFWODns1jqoXZfLIcHPGkdKhtq732GMYAK
FFfTThapLFelSQeqAkvVtkgmRo6pdMOaf6Q86HX8gV1sndRMah6PQV4RTMqDSipI
E7MUy0MU7PI2vOiZuZ+JtaS8o5fAU/XXQ01pO9bG4hlnZpjhRBLwWmqPIaJzhTCW
Wuu9eH3/UPNu6FmwItPBx6AS9mAG9zziOx2r8XaVR5qnuB5Saa4NipP6g5wMC2sq
rSZam6e9JG1aNsMUqPdtpKfWdYXrX+D+IbO4NmbDNN+qwVW06MypLFm2V1sCUsnK
k545fza0vOO5mNPMFgjboeRAOW1ZwRH2mFaImEdhSq8pXys/f4C7o70xHEkXNV7y
hvE3gcopUKUQ3j09T66544AZPErtlfnwTgN7iC5DMv2rgqZY9lZm3pUH8XVq5wJc
88QtiozAR+G0JZKjMzptwhUjt0+Na8U9cRVp5EGS6SgzweZdKaveH5RrZYRzzJeN
jpDjt0utWT72SXMwUMnWQ2Y0qMk6ITVsSRXIMJj5q82J4zvzOUbrJtVFfJkAb9PB
/dJ9qP/Dt/GSKyHIuTUBbojbUC92BnXFbykxnbaiJPDUNFfRmzyVW2pS8FjtfGKb
F+N2N9uJ3MWzK4BZhf3GR9lRv6E5NSFR4S2ZHv68dHsohqOmyzbmLRiccRRrFjtg
EJpG4Olx92W+cNhbg4UgHCajqR3ntAWvX1DO8H8W8YoYa+/XNFzkwoIWshpZ80u0
NW7jra2edW5SwxvhMybOj4N5bD6WuAxlGm08ra8PH0ffuYP2txd9jKVKkco8GJ1S
mGpfFZvS43dsrX6G7H51vFWBY3MMLMVZ/yTlqE4E5ILCcUt9vIHKcIOgF04anSok
Qk59MrCPxsyi1K6PxHkTOwSa07BNomciyG10x+0SVs7KwB4Kf0y6a2Cvqwbq3/v8
IaTFWSCQjlJsDMb9a247CEPbVP5BS2WPoC7YPAAT6bWDTWKDgO8IZ6e9RAdx4ojq
8H9qEDCwJchPvT6wdPN3iab7RYrk4p6bzdapy1uwFs3zddrW6JDgisCvlfjf4O19
dtLyouq4PWyGiV4mwYtpfmH8Fhz7mC5R/g501Kc2PIBp+eHWK75niVs0eS7QenLq
8c8IHHlFTUU5hHxjIIJKwxl0EjdfqJCex8AuT3K+AFioVdsvVeyzehkmq9SylKrj
lZ9cBLQEFrR9M44sfP6iXGjdv54Yu3dUKIQSPkyPHg1ovn5raWgI0EnETTyY9Py4
t0cjkiSROyR/+mVJjVXY635X+zIeEHqnXgcpRsLHq/fBGTbrLaOan5m7/F+8L9ne
xPvAhc11ySpBMKCBAKrGx4Sr0xk1Q4dF4s4YZfgxV4zpCxeewbzB+ExN3+uT3MeX
l766NCL9bupnYr7JkEOtqG5psaolrtLtYIIhurvlM3sPGqtseYV4yE7GfXPoiQOK
LtY7xwVM5bicsFoWs64za0/+PaPDTQ8tBM2ZXvkAF6D990iaMQgUTP84m7xNxXeX
b6ZuEicK0zH2Ku2pNewS7aBf+yXjTpvm4AkjGfjryzVBQ2EnXEKco0Esh+n1NTdz
4T57gSGKk9BpRZrtt5//Xr50lsGIYuZ6YMMx5VENS6iLwzrSa3Cul09ctTJqHru7
eHEe4Y4sR186/F5xYfBcXExvxV8TI28UhSHgb25HtZr6TYJF00LUmEUjkOa8boDE
kaN+/zs0UXvWzuRl5Bz9PC65V2M2wScmxKwAADwXIIAaJOkI0xUBcTt6LdGtJZ4/
17IrI4+OUuD0OXfpf0VgU5bYaPUFmsS7scqS+uP3J/EIoLpYytpr7VyesKzE9deD
US0zN5gLKqKGp38PE1hMKkfQa7XBtkJgURk+hC03kwe4YnRBf/IKBOQK7zVfpKnE
VVxDdMnnFXew2ebelbf8hwPnYAUJFchzpkAPDpfSdvBVxSEuE0SdCbVzhen9jlDx
6yYC7r87b7oLuvdaewV67HS+AF1y+pqi7BAMLj9V5gTlwoNzLipteBHVs5ekFJdl
qQtDZtzAdpz6xkhEJTUAzW3YWGNRnXIezS75W0V1uthmWcqkcmaUkWL4g1f1ksu8
uIKVY39wXU/ssPdTKBZblv7NdPHLjB4prxVi1TR+rmwbEkqmFCu2RdKpI2yzIY6B
y/muZ6IqyCPpmrQzDX3j/Ua3AU1rA0hRw8OahnK4lT+HEmp5zEQNnXrTE+MhikAq
CEb9c7A48dYHZZPLvYuJbo4BPU82/tIIv4VdQSlFd47sBhjwoCW7YBOXS1F5mtcu
1ABL1FoXIjAjwwBO8pCLCcs3i2zDwX9Zti0D/GCuN0OiChvrWXRJvpuvGdScv7Li
f6tc/+rzzKeBZ8GIovVpACZ+Hm0fAZQuESX6qJp2sdCDUSS+ZcjsEd4VRPRQiBjL
o6WKilEu8GGZm0KuFWv1KPqlov6QigpYuKK7qhZIVLE5RIs+I92PlU5D6/36Re/x
C/cZeWDHcrwIiYnzWO3HMphIYjNCGdjY5N85mq7PGCk4OMYFV/lPZa9aOBMr48Ea
8DaShpOkzIv2fjkBjsrFAPEaVRfu2TD1secTMg1hlXgBcAWZnO3JJVUqwWO7rBiA
tK4bjE3dDZlJWXIF51auA/Vny5qZ1V1KYEO0gDPzxYZsii4GZqo4eJDjqvqVSDoi
qSaKrtBOyBrgKOzTYocMjQHCU3b4BIadaJYij0tvivlUnKM+WYSwvE9FuWRy/gLq
LEzb7FQgjK+ABL0N7rpg8RER5gd+AORaRwwIUbzu7jdan3fhvMMWkhSUq23yUZAW
+J9Ptyfp3PpdrZO6Tt7OTeE/87bHdRyWMD+bhgOFh76aUs67+BoFcYfReTLvcOvU
XApWbYwocyqtM0U20IYK7MWUh1KO9X8QLk7gkbjW4E9fATwsnZj+sGVGB4avLLnY
IL3Y3TcRiUV5Wutfrv2OSxQSNS7RQk6UotbjLVZ2BWrv1SGVwly8yMh81g1/5eIV
/KUlpemhbTdv+JfvDxfxmad7352QdqqFOVgPMBOBYo/QaZSelumFlp/SfGMfZH15
KG5dkIfwE3owqym2/AyQgEmJagomp7pXtdJ5/lRIhImly4T7w2uGMrUaYlmTCf2c
MczPV+FpIKrc+XpT3CKDHvRXakE3BAmZCz3BHDsODbihLgf7u0a/CkQYOpu5uG6s
LHfPoESExj8ATiq+F2OOEbsPGCBdGiXMQZk3r3nXkeFcqcZXQ6TKnZyASiGWKzv6
zT/5X0EOIt9o+CxS4jlR/G7ubZ8AAPZQoM2MmLRt/XZyz9eh9ZyHfyarjCzKi2zj
qSNby4DTOkxcBNHck+cJsrDFeI5dmjkEBYgj6j6V3G5WfBlbH0uhU5h0NJ0okjS4
bAl2nTHKZgAQTOK9GjGb2gt5SrEiguEchgi1WcvImi5uIqM+sew9tQI4KQE10rKS
JMGEKZk0QgMCK8A1YPl4teukAm9nCFaA0mUPynoC2bp/i2uX7BnLjA9nggkNp4t0
f4ESj7itccmKKmmH422FbAilBihofeuZPovpp4sFT4+yZlJSmIGiMKZApfCiXUO6
yvq+9axr+4PzcAHKk8uikhR4iJd9Gbvt8hq5CFFnCADdFnNywWGAhzjTB8fTRmre
cth9+KKYfolUQuNked/sGPbiVMKulhEkTkRJC2pWNdULUL7SJol8FCDtH5a6peVY
Q1r7FTJ5ean1G5KQ3NyCpIjuy2QAvJNf0stV/denm7phJdf4VsUlcQiGTRxeI7OX
HC3Z42bEx4VKd4nYRnjIbQnX79LbMlWd8Hd4oXKlzsGWBRBuWwVoNKtzkSBseOdI
hS57Lc/4jba2lcrLUkXTxsU4wMkXNxYUqr3TeyqWKm5ae32m7LtTmnvjQbC98YAH
Ut5agiPTV7y3WHofAgMnpxvzW2y3HHiSdBhpu611Z6+W6gE0HvrCunzK2PCZ3mjL
oF/76Fm7ioZ5eaLb7s5+JfYt4b0MCIjqZPjKY35pJI436PGjUPXz4eeWqy70MtyD
fU6vcYnHxejXw479FG7jbDcGm1tScLv2vmWiJMr9wM58YhS8vwwin0z7KsuxaJwH
lvV7ad3oULLqqRxc0S4vacA9kP+l+0IzWxSDOuR3ecVXISMPkZuBYRA1Tj6MjPzf
bysdXZihtDCrsqJGZRwD/CmA8Fsh8XqNPwCaaZkjvp8ar+bjgPcfblPM4509EDWH
dnuB2dfA24Pm0RFhGt7gdXt/AH3jb/XGzPrDhRIVLXdb5aNeFRH7mT2EF8MmCg2N
aWmeOxeTBCqD3knXPFBngmGjG14KOM537IBMS99DahlG4QswaiXyq+arJumiy1RX
m9E0PwszOfuk6xlC2qEg4TzXXAllVT3LXev6SdUgFW5mJ7+MJx15J3EY0RpoVCzZ
vjUtJC81gq2ZBA7yaoyOkzAZJvcOZPl0HpKuPNx9Bn/8O2LQRVLITIGNnL//B4YR
k2jTcSC++zBC4vK8KBjlqa6xjSP9jBarO01q3f1VSuq4bExJiDfVnqC4FhzqZTY3
SNkpKeRNSzGAni7fjfp1+QoGl+noGwSWZupVwas7aXlcRZKpntuidBaDbhFA9e8L
d62c2Y8Rivo8ssnG1Ei/xHB4lkC9yWFrELq4G9AQryJ7cNNvRRYVnLzT8oFpb1N8
KBon/Ki9thmOULz6tc+/REAsD4o6eZe44zE0YLkj89HThdm2pUGg2wxNHe1EaV7j
RKyQqCukXWd8xYFPiJc0+ozeKNqpNefGkk4zvyMszcZbF6hDf54RMi4Go52RDTYy
NodChn580K1Glw5qcDWPhad8R25Fg4PNusytLiN/3TGVHDFiG2FIgnagcgVgjdcH
QaZRkdngcHKjx2pCQ6zTTy/gWILFiIfztX7JzZNpEWhTk5o97nCipeSYEi3Tj55G
ARw9Tl9tuxqAMYGr8eGD2sGke3CSzwTMmkGvLtk1MT28ytEnKyFP7LJPMddTp9CA
CLmeeHtcEU17aM6mhvNI6tYPI+x4fzzLpUn2WBWondwVcMqaxWAEDx6j8FRHWBf6
eipnClPo9Y94DclLq6PFFj4Me/LOQ9uh4rBBrPgkgIGYWfnb2wl1o6dGsQzMbZYI
BCgNPpFBeBKRZWx2Z/23Y2KNJ5Gzz16hJERu5W1oMiMx/g/u3+5KV3+Hrhdbm1AN
cLP3Aa6EjZgS6dJXV4FPaAnd5dvVKA05xcA+PmIdVEyQPXSPWvSlX8mYZxZGmukA
fUVEyTLrqCBlmINgB3fFHubhI/giHK4DqGmi/+k95N0BCZskB/DgmFltqKa5oy01
fOWeXfk2hHtrdrlBqP072HZ289JBcpEGETTn6XGFXw7VhV+R8h9UJFaI8H+5H9W2
d0u4/pzTtxWtYaSo0J5MX5QxHsdOaBFrWAaYR/5dUqGC5M7HHOTlflMJDCE0CkTn
1Eq6WXNXb1J4YjKojUB3gYamiT0xh1ZS0fSXHx5aX0fYUOYojof+e3tPJUiG/m8m
tb1D0GecxTRlzup2DQmoP20nTWzndNz7iupUBZd9grBZ6GHmkIGbwz00uXgng2FO
a9qKNOU8ZaBMLHMiHgLeiEqPTNoI9m91fEf3c3XOoEtfc2V+aoeBw8+xpdaEgkw4
bPkFrGahM0P9sZJ3W0n0mwJgQo8npQEWQ1Z4FXU4GWByDFSeZgyMm4Q/AtrNQo0i
kBO2VT+WQg8H8tyVeOJzv8gRn7dqrsFPpcwRTOi56F0Ai5mpbc2WX9tLnY6GYIGh
PsPCdDn07vlfPalYIjlgDA46gxpkRVPut0nm15tJDDkVAoXpXX5lgUWaYTyfwVZo
Y7XoWlp29+4TItb/Qbkquwq8ZyGQ+Wl6RguHWsQRDh4GEzjFmQkGZCHObM7W8/2Q
c8IB7+AnNYeKd5D0sSVwzmpLP/vLk0Hkfea2gCvnCZzJL+Iz4BEMWU+EHCuudrmE
GO7W5Lj+FjGdn19rXREWkdctKvebb4ipaVw03HQASiDMRmikrvg1xnOfeDZ5p+Nf
N8+9qjUNv9E3yaSGD2vvL4Xekz380p7iAUUsx3AT24Zzkiia/u2ySLCAoVHGXqCL
gQ7ujdLui2wcGt1RrcX3h7OZyjGL1nQZOUAHKLlnNErksYjCnsAtcmtZdKDUBXDf
c5CZCPg/7oWfdwXPpnoSXGaPvQVIoVCsxRs/X1HHa0FJ3RiH1j4eN06dv6XrFiBB
juc49lDX+DVkeJwrBy46SWw0dVAyWNMhulKwHN3A8x8wlGf7zwqO6PKqFiRxzn/x
gpen97YVYDK+I3yxEYBg9ThbBrUFT+24jvm8AWC7pJgImH4+TFwELfS0JDD3FJee
FbIf/8kxvdeEZTjMvTbwCdeFztoIGaxzJkL7CmtielcBrRN9eLXG/1g1GYCNAFcI
H/Pd9gNhSVv2S1Jap+HKxb6wUB+pdt8nBrB36A4sUgh5PuFiIhQAcedV9oGUH+dc
QjfQ96JERpvamwbI6VWSBr94Av1o4QohtNNxHghjc+4M5aVM7y/TV11NTprp+xCT
SaAwzlEV0RYz/u4Qs2FE6Lqc3wZUsCmMLBO7y4AuXgGJEusSABa72IltsEZn/HLQ
HJM6y26iyrV5qodFij7OLcxPQTedITNcXrjqEQN1Sp1XyZHqNlZUSCgwpjHIiPWw
qEOQcVTnU+mdH8wkCisCbXq1E5cg8j/cwtsuHv5hYMEfvtTOXnG+8bEj9bUVEHCr
QLVspY03jG2frEHbyqcdxo6D70pXToTWvu69K4LDfT+N+/l0vOFVa4mY7HHttRgm
sEKazrS+ZQH89lPW7XfXMDtT9zLNkv+WVVpAV8GUkp2XoV6LO9f8o0AeoheloEXT
CkgpeLxiqWjt8d8qm1+i1oTs4IRg3Y6hafSCVEv8cKoSFAYsd5Q9br03f6ve7I3s
RisCRi81GgtGXpjJGflLfJJLRBnzA1SjZKorPh7BImIQUrJJ6khypKn+ZRxsLgXV
BYvI+TFjIz1p2RMelW3iDsITaZjtctLTQXG3dI4oplbtDi8hZiO1qk53QKTeCOpb
KU90ZASPYdzoV0/YSd5T29zBTaPGkvx6zK52m3+3wxuq/MKeMA0Q4sT7QRX2q6fT
DyJVveC+f4jQazPDy8egmRhIm7Bfc+INgAug7qJItldbyUllBBqupWinU57GXLc9
BNviBHplPd4poWSWWP2J8JWOlpa1LfnSjkyalBggGWVkIF97ZMY5wWmC9dOb3nQl
vBMNmRFcB+wDHMWWXaKgicEGYaXKPAdMa0AVcGqgilcUo+V1HXVgJUuZav6evFr0
eLf7VaChdz131OOvHPtSNwaU7ssWL+DvDu2I+ot4Xw+wPii8XY/NUNo8DsEpGXSR
df0RFkUGlXohAnysRzhDp9fo7blP6LzvVlzuqmnRQp5lkhVvsexhR6BzCMgnPvvS
WvGQMWKuMgTmdx0cnAVFoKTWTt6Oyc8YCIL40ACUQ91LIVsKf/9BYBK2rycvYhec
Kc3dUe/ZZNaxjokJwShYPdB5s4gvyAKKSEmpGERFogqUw0l5RG+cnulN+lSamMTx
Hwk8S85ocxzEKcULEcH7Bn6DkYKJpLGl5xA30xkYfIjigIMDdm8W/5WAKJS2+CcY
UMASOfPEUGwHBvFfw17wos7Ydd9GqknNncNUNB9r+7kaj00uEDKwrufbvTD47GYo
US1zCF6cAr45CCjaZreQvzUwfAZXcZmgJYxTP7iHOhZnhpss7yP/vwEqzfvk7VtJ
orMqk3fvYfztaLBK3ZjrNWmVdTDRgoRCbldyItlycX9Y/Asy32UbJp/EwOSjaLPW
PWLL9m/+8xnoVxw4XswZtxLUd94qqVTmGBMnFGi99+ECYgSH/HFfpP1UTVciJb07
o5Bb449PsF9q5vT6jiaNVryPqVQkgNn1DzvMlhQxhMT8hf1rq+u9VgIvGXoqtXH1
I3HSO9CXrlsNhjxn7hZlwFUUOzCaGNqk3o+KvHC1xzUHlzw6KJwvwq15jsBr3HGq
olLDlN2FEGimnm91IJFWFuaesiPrujGih7+MTzxl8DSHpb1+bwCj167nIl51n8xd
qIAA4r6T7hM7FHPBpMgetxTUDo/QUt9EXRha4rZSGz1rRTPpQuUFNwecRFIfl1bw
GIYbm977r5EFVQ2pRCk7kjOJu+qHwBeGcPSedDQiIaBAm4M7kUxKKaNfyTtwEwGV
pjGSoo1q0Iz+p3dinnV+nS7woZmKZ9onLtF+4rDsKZfYh76xGJPghI2KipsYmHpN
wDToxigPBajrQUBuA3Y9mfcrFOto+KTsZZVyX8sOcnH2PGE13BpV4Wh4dwgQ5Kza
IxSro7vt/FU2P0HESYmtz33AVQQ8g1S6LMTx0XMR1UF8WzxUJs1pw+jC259JNAIb
Rak21Xekj14DkV2jQP2wtCv7DMUA9pKl6LsXLjBFhEQlSVQG8RlgNZJDTTL0J9HY
R7B3eACrMNjKmzWXJja03yRok14QDutyRveYq7888xktMoenCT8i0gUHeqe7oipB
2ecynptKe/QhMQgxw1WRZaYMSqHckr9HpDSQlMm51kl99c0R5WINgRCYJAEz4ACz
w7ivTtAZKnRFLZr+5v191wowLuXv0wZWQhlpdRRCLLcpv9Y3GSqzqwL/EEk/80rw
wR+mS6qegpxQpo4TfR77p/QbaiJrpphvNoNKNQmUyTdZ6AzUD1oBMvhmtx0yoELE
W02fz8upXjmnk0HI83Fs0mRdHiBCNinuqZOY4vc1tTEREKV1pEa6axu2kbxoPuy7
qgQHj4sAjSMzb/ATqDUb2umPfWrhZf9A5jswZRmCZ4vlMaqbEQ+kxv6uKiH/i8mT
gBd6ZM7DNfqC2wBoH6m/oSMzi4+O9Amj/rUCaMF8IN/5Bz9y+3LM+3+j1UckZnLC
scF71aNWlcCZgUNKyzuwGiD8ZwmOZxsAB63zLpR2x8d5x1hOHhq09Eaj1FAGzkZ5
TlUYS4f3FA1CJzyTwUFETo9Z5pBhcd6kOdGDT3Jvcs4GlYKxYKF9h8N9+jjbZP7h
O1wg2fo5ySShmzJFwRuxYliWFFwjrJ5dbSdPFrsmsooKhSnJyQSdx5QJKbxt0Uqd
v56uPGg5iWm9yqHFTCN4QBm9WFJtJARq5zoyL+uXO5rdzwU4KgCeegiNMDw400li
CuFSSGeQD8WYeFGJAksH+rkX4mqJ/NUVjhukcp6tYZ0LPTCCWdwlC2ofMuaoJopo
RkRrmfOj1sqpZYL1s4I4cvzJOHx8pNWM/qC5H+KuJqEDF4ttXKUhjX4+BCPGnwnx
/c+qlbSuH+0TP5NUjvcMBVfrhgATFWEmRKxgITD2+WBHK0s7pGK9YDH/dM1kOh3X
ipFm2H6cwut3YnGPdGEsb1TzwjF6NESYSSTB85qFu3Zg/yBJ+Jyrie1J53YD1dJ/
C5gEEb9tmU2B+KU0mC33QTlrYueyh7YQxu6kGoaZOkrPdeCDmbTvWyzI5V5zxfFG
uEgjs29nDQKVVh6M4NmYAWtycEWlXBIgXo8ZBtn4y4DErUhBT3zryN9jRMebsc5R
Go52i41zdLiF7a6Q6CTyciN3z/O3gGRY7JzI6S9rlh4HIZ10s1ZAIf+gJxkVOY67
yUAtmx9LByJcbbEpg/xdy207TRRHnZKpEewtTXufU02ZDGgoSquxOBkl4+6bfJTw
5Zj7Y0s6WrKB9wtKl51E73raXnmSk72ma24KzmMmVXhsIkYHdRnmqWnnxuIZrwre
YKJKoV3PO6CIolLOmR8KLmD/7f2p4wFOxvMeeYZu4PdXK/NVhn1RiNrUbuGALpfV
J7pTxdC1kWwbZWlxj1lDk7P8kKxGcmL+tCsvJ1RgQ2JSdS8KpN86VHI2fezrc8DZ
ZZTlQT4oJlKQOAxI021KLvFoDYk5yk4ouVUkXM2qO6PKI4ahbqR5jlE98nOAQ/+Q
3SjZYZYAfT2TRRbm3jU1/2OCOPfRYhJ5AaCAXQG4yWCMpTc//3+TBJgYdw92Fj6X
Rw9P/ePcbgUvH4jLprgGdEdMWtb+3TEY/uJPkWmFT3g1YPCENSOh49UIB1HzzNuQ
YABiKOyHUhyWfBXKYnSlFYF9f4R9wu/Tl1rlD2Neb1Zw/FJEqdggPWHYYSbPSLke
VxkEcroTFt8II7Bl+w5/gjLZu37hunHOGW7LEdXzMfMjfXcdtySWsOArCUcvZi2a
OBSh0WWb+U3WC4C0w7/+XEVnlTOpWCEcrGT2f/W/JcDVPmr7UbaXmD/ZNVeKPOaV
Gh7FWrFWEc/3nGmw6lQPqbQcoc1LLoRbcOHjcu/I0GaWkbdJ2+O6018hBvCowJns
ZEcspRj5tvB7zvVGcQncbNNsqA4Cq4YFNne3wyOrogQ5ymayMSwx5NrDDxyoNBOF
d+/wzO9LFsxKJmkjMfEeOumf9wyNEZGrwx4dPFOhXqrt1f7yK6eDYdpC9a7ezKwY
pXAd5WbGJQ5DYkUkxLHB1VerPVcPW92/HtIjF9fntSCSvRI7oF/KsQ+M1OrV2CQE
lFu3/xwIwXuKvyDHCaRx4DTGKQu9qteKWOOFEqBhygO+3GeSSWnjaMkgWMklwEG6
KWyq4K3D3vMpqiu8yFK4X4S3ZZw+TCTlVisCjLee47T7bhpDv/OP5512TrESeIDW
Rg7VSwZe+uNj+1Uk9/zG//7roigdda+S5xw1qAKIDjDESpypYtOibPYRlAzRJ2KG
UEE5opg3c3AHxwHmE3cvyu+rptwv77lwWfSyZDDXmgqlNeWa7DnRF70JqJYxIWS1
ZdUdCk5IKonmQoGKtsPW3sYWGtRIObUclHf9HGvncGWAQZ9TNYj7X8KlNNU4mRSn
eUn9h/3oYhtaHbmraXn9UvrG3OFjWyOGvQRc44meobV8ERXeddX9h5MJVMEyIGtz
HKjKTiz83U8Y5CuIRrqXWYs0RA4mR/RfQ2ySmc6qwesGP5TmFNiLbw3MvNsDVXOP
EDeP+pwZsfG68YsvqBOUBoscNc35QlTBOm+GiAqrIFFMARbn+W+AqmZ95pxgvo0W
OFNr/dKawRTLL1I1Uj5Ph4yLzjxpqs5LR458BuNrmjmye8iZsMPSNvbyzI9/5NVQ
lyRh6Y/G3roOo4OttSNBdx2RGn8lFeBIOMUMS3g7ws3kAsKB/wkny7B1xDTcY549
StHtWQRjeJTC/RDammtxLyi7OKje5tfDV4iE0nJJacUpj4uZjm9xNl0f2T2oWabx
/cpDbHwKzRkswsTqxGcp2UBakalfIoDj1NwBJrvW8MMSyDPFI1vzwANCRZRhMXsu
/2aD9dSq6d4UowG8oe6Kec5qRaDR6UTHw1yZNW0Vq5u4KqNarIY6exHkff+zF/7Y
MSdNaTkY4xNnzRdDJkH8JXsMlpOoHPCZnViM4kD38bZZOYu7z7JPeSQOQjAgbne/
HogoyhpdJSVX4DMO6D20U1fjmJhpdy8eGyHHTPmkERB6uYfwkb733BiRc9gjPVer
zOLKwreX8gQTMKj8lL7T0oVTbcn5bOsac7KDESSHeM0dyw9ss3b7vlmibFRChrsS
fnHcJChq2+8iYdV2OO9oYUyoxvqFYPR+4nFLRspOcw6UqYBnQt4Xe95vFGqhG20C
3GF52Zz7wrwXICFYj4VaroNb5FTTrv9Gk/CWYw3qDLfW0aWg7hCkgjlHxaHGOCq3
Cky2ky9A7cmEeM0jlZ4IzHkoFT7OpbS9rRH5q7VV7oG1RulypB9BBUZZvnY+gYvp
7reya5M7uRRUzZezK1646vrrXpkm8qmwcka1qSamdKiP1JzD23e9gdJapdDBrDhU
LNBH1+gHDZQRBn8uDcCU3ZtJ4Pw7pzaELtDLFe9mewZ/CfjKLmwAK1NPQz1HAsdo
7YGQh7697il77PEAunKLZRy3HqBg5E4eQoxGVsI6v85LB3ApqWKVFlw/uEsUZdPU
KmO8vhFGbum42iPlL5tdI3CkwYyl4FynP6zYInUWzdSXJDgJTlJsjXhwkvgPUnQJ
ds4phhVMWIUPa71UJSfR31OU9VdxUsLFVSKuaxeJ7EkiMkJ/Ju7CnOkxpYFntukY
2+GaCnkxi1Hw3sTQ/oeYrE6znJa2INebWGYuojM6Gmotjeqx6psAL5hLnfxdcIXK
5Io84hRO3vGvlQYZAX02Z27usCJ94huef5OthUrtVyuFz43w25sDTYSliV/LQpHi
A+7TsngC8CrNk9IyM9Za9zfX6/yg5uSlhe3ptRwnSlLCzj/2d1EfK6t+gRBEoNnd
+yHzC64U1WRm65jToLtgvY+g8vyobyqenJyFM0gw30bM4JzJ/Hc+8VTpQ51b94W1
mxA42p9MAjDZJolkbml2+L2mlU6nbQO4dXblbGyiczAoCvgbiJvElrcFSaeLtSON
Lzq5iOqyrurRqtuFWCcHFi2BtuPFAjtY4jR+DzdCjkK/pU1pZ5tSTHJiIxbtd20y
1IRQ23bJL6cI4zGY2kUFSpzczgVtMBNAlT+ZFx/2kNXARZcNwzHpe4n4ROkIVYOZ
qarEX+mZJxyQfn4ijNJ04ZavFxG754nwMCbTcfccN0230oG4dukA+yApQ5P0sVjs
eIS+9MxSHOWB+OY2fxw13CTsohT3ePXREF2fWITMM4XhobXgX+ijXwIwCSfa5U0L
dXOF1NsvFRIjzcgMshZ0S37hm0Fk0akhwvI1YbiXU4E6goi6IHz2R+FV65z0qzWI
fEShNQXXaebM7SGG6XLEcfcTEIb/WnEnMg0dtvJ9sJGYBIR6OxQCWBUWFujvDoU+
Gou8zUTA3ZSGEvSL2BLWAbZAWQmcmOlr+GhojfzGqwTKXKxd3kEvN9tzzeSsU/WD
FzHzlNISUblYTPK7wRcaOIh7rW4g3mRLTPBCmggxksorlfgqwzK68krZw8OAcJn9
GrZhVobHnM3isk8kgUHrJTqb5fxypqY8j6A9G2RxKKZNdTdUcg5PqMxV6c9s+tTN
CgzMfyWFyIfgsjXAz8vx5ZVWUrfEPhgIDzyA4VdNM2rLOlVLjP/FYWNr/egzD4mQ
jtBQtX47xgPXE2awz7cVfFHmXgSSIagebkB03QGHGnqm6CD+RkNOIxsFmm66nyQF
V1ruaMB+M/ERxO/JjyHhrqBLsJ7Z4uDV+91zHhEFgfnnNBYK3H4BV4AS1+0tPxxl
9gH8I5bkQmHtClqG/RIgV8aNH/8CoB1eCC6p3fZBWnifSyU8RTjvSh8WjwgUI42s
V+80UDAJF8HGoVUmZEtQzQj0AUvqmuY4yY6hd0GTuszRRqB2l5C5ihGYhfcmVLo8
67dmtuX1Msj1q6VAwXBm1GJyKlvvUlVHjsdQ0Han0lAcUhYRB05IYnAQsWzIKNBP
rLhGoYw16hF/REHvrExspQ4KbXJmu9llxRzOlZou9W2PA3BgR84Pa691GdxOXwwy
rKdihga+2bUwFwa3w7h4vKUl+cbwkJZ0Dq6wyT+d5Ytn+jFK9aulPyJ0ukoa80FQ
8nReQnMePZqKcZ6zD65zKsKXIYLy0qwwEhmJ5xpAhEv70J18K23YVfSYwvJFNtGz
UyVBEb+VPlle7LLgpYG3lb3Sfo2whPUpwji2R94SP8zcyLj2AjXmz8sTTqhViRZ7
q6wYPMyPoiIafxvRkgZjzRnDwjE7bT/nzW/fId+kZAlWoWXaCwIChbprhUQ9i+n8
IbjUOupL7ruCfJzlAFIIFlgLDJ0ZFHX4afJMizYy9HnlRXMjiOTiyUdCjA5S4yo4
uJ3u6Y1OCT7OQdCPfpkqIVsAQfAx8k9wvjC0XDhZu4xYVWJrhJrDK8f+awfpHNFk
LJhix7zru+OFZ9gsUZN84ouSryACBTXdvZM7bsYX+W4w4fYQUr+WCxsz7m5/AdOH
o61WLAJtKScBBYKuQhG52EINWcdavw+mpNVcaLJskjlgbTo0+/c7KkaHfcYA31fH
+vQsA00vkHEDEpUVwk0QDhsmuW2ytWw6mirXXQ6yhVi8+1TjvIqUjkJAtPJzYfO3
0U31J/F9AZ8nBFRALWRcza9a2MIUpMFHpSMXwgRDlNzeMbBiN7ksI/1tluZK9oFt
fESvYGvl4In8i17EpzQAckIcQ6Ftm33IUBrqz3iAI8x0erZpIz8J9GLfLoCIZSIq
lrv5OVs+ORBupdf5KBLnqJ0Jt/WupcpZgpNN/JCW3jVGrPVtBgUSsBBLR4K9/VnX
j2fvTiQjd8MGHuvmmfPrhqBpfC+SFlW3schnOOwsRKs3ZVIPJOZ03qsj6uFGfvW6
ubb+7+WbogHKpBDR96RJn3fTJ/DW06P3kzx8H9eHpnAbZegZhnotht3HwMMuz+5o
Ghl7eLZqIWlpPlqoszNl96FRQY0wc3nMsBKy8r+xap2KLjTJfzx2voK0lde7qd3w
GMBSMir3OqWt7acIGjnl6C4jq91x8ZvtKIL8zoarsY29rjFJUJqKYOIeQXOpKfcv
fbJjiFv8UkXiWTWFlmIBBmifOK6SeQ14bPQQPro8QZCkTv4NOlNsfYSrqdfx/n9B
nQOgSwlfp+tj/BBHnW4GPf/vWZxFkwXdq3xKpWOcf5JX4ltFXOrEBgb/dk2p+mrH
BanlgG74OBP91x4rAC2kVePJqw9aFhzW5v7sxpX0O/rzy0MtzOB36kqaXWST60qn
P1kjq8LrjAXBZAjMiJBVQ8luG733QuBqdpBBgIz3nB4IjSH9hp50hW8reW+ltiSP
YPGLtbfiB/wxNtv5lGM5rFs7jhViVnH4r958ZwME8X1qDblk6OVmp5IiHlhTiyuB
QgrtcYEMmLFYOshrsXmzsEwDb9Xhq96sq0cNvGHA5oyloPrhJq6U4K3hFGW3lM+N
FE5IzQBm+cCiGnVTmLx9h5jO16tzpBiRhwmlKuKu5QBRCllwC84MkDXBiIsfoczp
gAUWl422isp4ZQJcv8JFVy5g1lQlLkeDKKAC+CLKiQkfQf6ioYo4hD7s1D8nCZrB
ZeXZL4GPZO51ZUeYhfL/PZeoPIrWtpL/TC10r0WtAmfMZnRqepx8JUSG/2aikouv
D4tzg3jLr5npToFPPnoLlbD8tR88wsVnCPshIWo932jac+bMI+VN+U+GeWHjvaLk
XeRih+fx6WzcN746vqSkMkyzPSNcTwACIqqjIs4tTdcmbCRPaqHFv5YbcvBqRbBu
KitnpbekATIvBepaJQkiDkFsIvjEZgVaduWoh+/Fz5RjCHpYKs1+VefY6LhPmP3i
i4M2N0QM2U8gWTtlfHWRHw/z7nO/IK4UV7kBiLBD5gNJrFYczd6DVntUB24X/zcE
e8eMRo8PFgUgMxIembX6yRpwxM+/Tm0bYdEJIfjnoM/UAQyugQaKGj/99wXgq5Ng
oehG0luVkLSLMs9y//j5rFIZfXxe0k32IPBJETtqD1pTocrcIuGQEBC5jc4jsDu+
pGERovHx/imVpFttE/QLhl6e1yg5T3vGP88TbHQ4ui69RjHSrOYIyrvkkGS7mVPm
Qca8HSclZVERNKYgjSCAeOQhzUP0mtYKTZ+fpsKexyw1GUBHmLgDzK8jSnkxN6I4
Imfn0pp2MzEJgu5WsU1fux4w/N3ih1NA6JPKtMtGXWOXRDdptuJHEcRqCByVQ7aV
5nOVx6tEXMVHi96Ac89kdwXuMrbKlXPQZiK9qkyfzSEfIv2HYMp+2Qhqfz5AILp5
ztnmP6+HgL2Svt0gwMPAcZnlL4uldHTUL4AnA24/Mk7EO+fGsLinnLEPPTL3qLTQ
hejxyYI4lmzHnP0b/yOXSLEwP5t01rRjzqscqAvieUmZVTutXKUVckI1vNNEDE1t
zFZUaFfQOpkNmZyGEZYbY0p6RP+Rdj1xJXmeGYw6gjOQNjGHoPkjPKohaxlKvScN
HEDAkE9exBgbs1YozUcmAMPgRHnqFQhIkzi6KxgOE4dHMZchulWuyMmN9O/aIBhC
+AaMDxD7L4bPGHVzCP12QuemMRPyLxW7i7CvrwynUQrZGN7ZJIbobefzDGWB0hWa
VdUWa6pmcgo/miwxLFNwHt45MaZuGRMn1ZV4y27ZI/b4rcpBdVh8NW9DwgtTWSrK
bVXCVARw4SzaHJhpv3EJUw4alpGiQhTlaD4ZoZIhmJ2qZT0Svv03HdxX/cPbWfr0
dRg9i9AOdOBGEcInbL05G4YvgQXx9vawZ6BFmER7wy9I5NfzGAFb4DU7z8UQgYpP
rqza9N5wT565BlYf7+U338NYHg6fGyQ/2Al06Wv1WM4GC2O5kbKRVL82u4C1RYhl
d4TcDLdmY0O5TQ4j/a0JiE2jhFa7TghT0YwYGmwu451+IFGLT1kf1vGulkOiB2c8
IaPZCr5QCIgZ5wLXm9vYzsMn8sw36uiiZATdZ7LmiuGbx1IIjijh67PuT9xtuqw8
Ra/ejENNNiNtL2YnH3VU2t+CEkYZl6y03ws6a/LtXKIEMRsjEycHr8+nCC8z029o
et5pd2bviTQ5bV5d57MW0b4bKGcqJkwVhcIdlzPlDOG0B7171gqEnyaol9ek1F64
FzPEvzVCFjFHGCp+4wJvBztb5S6zxTUWXKOsT730rxJNUUvb9Sze1BVIzHpPcNYA
xVeGCqcdwqjtJ49yOAHJE5V7YIx3qiDIfUyFobrsjPqqytD6hi3WmL6L73Fg8D9e
mi84qnitEGj7zx/SinhX+YbBQ24fKWGgr1J074JwHtxUM8pRHTfSnLhBgPYbNWTl
gdYYzrGFPp1ggvwucQIRm+8b5x+UwIoZJ/DKEgQaINqQGepaKXWH+me1sYCWCDP8
z8r+bY8Unjspms1iTTt3O5yyz1wDNCel7fYUsWZA9QAOGRlDlXeiMh1zgVoqAsb2
dBBbXtubUitlOWEQJA87syt6u9NDN/SRoSpTl4/CSklJwSjvDyzjTXHno/UubT7y
1z021673kVglAPfiM3Kyf0jWg9LlPukW7m1pL5Da4vdg5wue2QK22SSD9kLhAHso
ltdi8ALP8QuhkO3yKe1JzgOvrasVj1LhQVkhIw6tt1Uj7Tjijcoi7Y95LeJLi8vD
CC0uJ384qrYtAqdtu627Vr1yTTT/00eyfcBFv2HZawWjaUXthz0Y5ncvKvPIyp5t
9KjpnZESYNXKu9J/BoQ2WS+S/mi8j9h0Ut8Otrf8eY5U2ZUBlab55vtRc4zLAaNm
3XS/2ZJgKMw2g5MLvW64NjqvCGV4tZZu19LI2cXj0fSk+em6dfPiTc9p5TlLLwct
1Nrp283CKafxrn8gIskwXxLVg+ciGXNdD5sBISgOnGkVk/TaxMeOfPTENRjNcaG2
vn6uskytrJQxeLtvjgUeuEI7zJQyhU++PCs91hZHqZZV64kEy74LGkQDbSlfiM3A
q1On/MmUR8qyyaazLCT2B+cttEUv7PpVoGu9J0FKeThFo5EAbYH+F/7LBGmnu3wy
wb/a1x3i2Lk0CCsy3S0eMgC188Bo1nH4S5hNJ7iKOST4E93SvviGdNOQlGw6dOo9
NE0NGRt7I95kL2kcvNtzvNAHPKwBxsaF1gwgVIjDBm0vM2pJuzsq/2YlcquV55H+
aYbbYS4zz3f92lYN9e7d7oamWpzoVC4Xv4sQhbIuZCzlefJToKxEsnZbfCrwI0nJ
s0ujyLCr2AaR7FVL79Bi7DuMNRkcCJFyGfdcTK52XzcxCLaTEcGM9x1H6Tj38/67
7Dh+ZY9Rsisr4B6HE6xWVlnHdS8u8PWGIgE45XWizPdTRDfHOOE+psYrZfRz8urc
okqGulMXWxB/Xl9ma8KCmAfZ+wxrsixNK4bF1xkYhqACqf9XWpRVvHG3e0QxSVB4
cPCSo7ZXn2zYce8dIU3Oo7gOFKbwiPH90NgrI0YX8unPtoYAEXjsj0LdnyUGbshW
jmKRhO6+fciaHxdNGkHRElRvRIdnKPklAWCtkGyY3tXB6eqGALFOI+KDBdp186Cj
HyOXIwUZ/IZMpG1sMo5k9dsjzZ0c5uzlNuhnwlHkeowEv7KGonajUxlR8E0kAlPQ
+dyfib0eWV40gW1R02xmXplaiI1D88IE4HsjHjMpmqar6DR9zJ+VXxdbIEfoxNpE
phtzGDo2uVoymcNidtdWL+HGpIpbo27GsrvDachhstWrLhtxhKyGQB/oojOXPM5P
5PYQcwaUgV3+QXfosUvn6KNR4X0x3ovGMTAzOrbeodxzR/MLIHnQn6dlI8I6cp6I
xNWTqM42OXTew9pxZzO5gMOxADC5vgcKXcSOIe7wNMxRDh9f10iaZDicxuH4JIIC
XVutjl3JyCx/nx0Ajgm2zzifDakRBKpFugH9nUK508qfBNkAjLy1BSAYRosd2y7a
l0EBLRlbHHJqy1rB5b8GmBfiFxvqMG5S4vXBeOs6SRhbmbXzTNl/jorAJPZ+wl9i
VOqjEqYGQdXBFd6Uo8Korshs0zCKdB+jKzo2vu20yRXjK3SMRsYQ5QC0x61IMa7l
V1ugN9HR2jiezZsktImrh+/tMvmZRoOSxQrJNLH8ACzoA0Fg2kya0Jg9olqrdU9j
XrbZke/cXxObOXuZjwTeZ+0Y644OqwPkUd9eHT7XQcH+yPmFXFQxjonUJZJRJVKu
N00G6b0Ep9qG9CeSQ4vBB9HlwobUbGpYyJAYrkGAglcaT+JR+HBLbO857JjzK8Ld
/vYxaRRQOcKkYQz6Td91zrP1nfV2xkWNw3qfJBNTJ8YHO7tAxuUDFp5iMn//6R+2
WfMtpcHCuipyhGjmv5BpJ03EnHcyWIZzIC6qmwA8H+aHsCpO5A3nHXtUclP96j8T
j2EhZYlRWE5pRg93TXn6c7c+vWXhftEO2mcoxpK2gR7XEhhBeiR305LdtWk6rY8s
yC+ff6czSOeEUcgLWseOMGVgy44z0gcedS0zFWTM56d8939Zu+OCmnre4+D4smRn
JZ8FkeJkPubNrbUJhLtth768BoUuvGjNG7AYgPq0tv616ABEO0Wfn6nJRh9NwgTd
hzpr434CyWfP7ZdW0/6wfTDWX5pa78YT5D+ZNxX7Z4KxjHV6hCeoVRhJKDNtiASW
lCGrFR1ORceZ09CESV+ybp6fmmaA8alyPxKiIXm7Ze92DBVJ3o8bFr5rmYXkjqKA
RbwalMUKnge50gN1/0KVZVUWhd2ENPXIWeHNPtWLHDezfzXUNDxn8vJIJBa0W7G7
jgrjX0IoxcvLyXd2j1dG348ZxqBDOrEejQnnOTJom3rrPTCiPYP5sPnxN+w+aE/t
MfPN8KXuF4Lz2fai2zphHpcimtDPha6N+YP6fsQZIN0B4JgyKwvJ0+g1Qzvt0ccU
6tpPACdljjONeAg8m6839pKkMIMNpnSgbk+th4pzPi3duaIVEUoDQILzFqwT75Gv
RUBHUxQb5UGwd6d61jMpCbg8H4UaIe5a3V8RzucarCTlOMBdKOIcBfYRp/wm3nnm
Ey0uHP+LWK2cH7bzYYi2yGdzQLD9oGou8BnYXcuJ15UEeh9MiOK28LwYHKyoW76u
dhpig+kHzerX2LHdM+y4j9223kgBTygDAOQXAuezzc5cWW3IOPvT8OEUI/K8ImPU
kqGEkmSQccuxUaYvgp30Vq6YEdJr+hcJzwXuwAI+RnePh6faLaVWahU/aL7GZ3z8
rlqYl5Vl7lLGrknTb+F4lvpfV1ruCXpd8ogqN2eGmQWDNRJM7xrwvtl40iL/9rJi
ZJscCDhPw+eo6WbBuS2yH/pRkL3nhx3vyBnf8IxaeyeJIy5K/RxG1IFROAfd55GM
TUSneueJV1qWNPR+pSPNAyryup82mNmKzRsBQzvd54ogIbtnhe0ne8F6lvAble+L
Os4MySFc7bV5p91dsfwoU8eRa3oSv6P2iohIoYEp+b/hb9UMAUdpOGeZKIaJezzW
W4bZscGHhHMARzEUNMGT1NOYSXzy1ZyZQ2DLNnYcvVi/zmHwK0Q+BslyBjtpNNZs
kouqZ+wE8lRRvF+p+WxvmJ3FKK/kYiuU4tjwimq4ZHpPyjeWhn1fGics9UgNTLuZ
Mw5Q85xjgP+Yu3/HpeL41mCnfAlqz1o1N7SqhWHb0vOVQuMDfqqnkL7JivenCT6b
990f+Ar5OlDRPgAXrzbZeeZFpdnpUYJ+0nXfzlino+RNTemrDYEHZt1ndE/GOaOq
TnTq6sMwzeExQKskYOZFeMpg4315VHUukln4QEeCD7sGfUho900sIpY448b5XT3v
gLMhIdKXWma9SjHyRwo12BgQJt54OKaRoI5g/FeOdECnoysSluhfvm4KBd7CRycz
L1ehyT5QomgONmt53WETP2JkpXpzyZqxHt+8s83zZWuGWkmLzXdNKKPou+2jhAjS
+gO0QGh/eEQSdzMLD+fgI1Xnb4EjiD45mT0IAFoC6776w/6qP830KG+H7A3oVQ/u
t4RnxEABD2m4IhRtfkw5LlT+KOvrFIQHzE9g+jvietior/dk/q9jIvhn+Xzv2W4l
SzEkEfvdQSZezSP+7DwtQzZnDpGlU8OjJ4ftNb2fiZXhAHJtfXu4ccY8x+4xvgUL
cnszkG9MBhbr2+tjVLtZDP8P4hDQsqwkAkCTNyIDX7Ahemgl9L5tmxNEmkcOlQYt
moCxmPotj9jFh9ffDSNlj9+nREvw2MkCcrF/2TeZ7oAUB/XfAlTxiCjR4ppELzks
ytNta8RFDtWMWi+EevgfMhpBdQNiprxvrikBEON6CU7CSBguzJAOUypBSq10xC4j
uuxeSESS+hsYEevtB4V0xwrUFAWzkmeFezuHcODRWZK0wqV4/FHmUPYvQdEWEFHd
Cz4f1MCQyFFcB60oGETVHZ1z6XbaUlQvPqNQebj1nblV6dcKiUA5nLorvljf7Zu3
27M6+EnmjqC0z1RZ5Ec2Ha7+aIr0Iokm57f6/4qd32XTpK0JoaaF+MhRoPRNMQQk
5dCNWTc0gesDOSH1uzzoYb3grYhxzsU949a30ZhAPb643uIwTok0mKYl5Wvgh5GW
dqLsqiYmmf19qd7JZdtmb7uuZK3YMAjI6E/idrlZUA12xatbhJUShpXPcI2PKrx+
XUD69DgO1q4j5FCbiIyNyfjkL89Hpxu2VY76Dz0cEqAoCUOpBDM9aCQshhPiqg6e
2CUbv7hpHU28GKJ3fyB978rhRWMwdIy2INEZecK391UvEW+daqq0ciLxBbzrb+1+
MqEQElB/kmny7WTHCVxOkNbPAOpzZTIQRbpH3lOY4d238IgUxjbuM9vcdilWqXKo
pgjrp/LfN/SxnFVXoeoxi48U8gE/AU0EMCwOptH42L87UtR3XrklXHMAHfW/GKwu
e+oA5Km7wTNCSgLMhFZp8t2BPfszc84YDqex099/ju4eWQDb5b7GxEfU9vg7oJSm
BTsY7oqGSKitMBsFqDbFvyd0625UWeFj3276QAKS0Fg+QYn0U8PpNzp1MBEmDGji
7qHsJfF2BjydZ4qKKPj+Tmxb5tqhIs+qQLkuvpx07HxTjaX+4z/6C6wk7i9zUot8
h+wYlX/5QXDmt9uZaIv9teKeqeO0j0GBnOPsWe8FSQ3fdkPsOje2z1SkoKR3nTN0
T0cR5F+bxfDgBQ2kZ/VPkbxMTkg+vRbN/GR15Kbb5gzSt7yhx39iBktbaQ1opc9j
rwHhGp9qWQO330nitdOvOu4sKQK5mhgDR7lvh8908Njp4VYQbnrZw0rUdND05BBg
kdzf4E6orlno7M1Cjo4Ya2JcskHsgYm3uQCk/N+S946HRsNrUiEXUEh1mzs7gNTE
YXRuxLRCOb+Qyl38bdhceKQ2IzPLvDoK947436xvx6pTLh+PA7yEOiGYKJGLR0Jm
lDc5PwVvUiyKj2sVlClMJYCCQNRa4puHORZDY7LKPGkZeDX4rQBcCgmiYHNsfChx
bJ1/cH2bFcJOBW3EIv04D4u1e0Fsn7aLtqIiw8ZW4w8uU8z+xCgi5hUcxhtkbyBW
tTT5nd5+MPUNdD0oBdygPs7Oz2KuIE8KZe8JJqhKXP0+oEL1vOy5Q8MpWMx32Sh8
880WQtw/uJn1qAMyoT37qsByczn7As4+KwtUxpvFzNOeXk/yK0IB2cXHPCgJsBdC
kcNpibbPzYb2LjdpbxdONS6WGvAg4CXur+fmQ6UXjufwxdJuHhfBPX26rnqykD3G
Gflip+xMW4xLkbfC0LqQrysnV6Mp3jTfT5b43L5RR3BWGAgsh1BwkD98CN4cJfoI
0Wfu5xL4exR+Ft4H6U7INWrtfFxqRsBDxyiFlxRGXuabdMohbhqBaWUcm8fH49Hi
1G+M0S91KbSI3bj/DbNF40BrqwdwvyP1QoEdYR/yX53AcNBIfavoGh5nGF86zaal
GiLjYVqNhvcFfNB59ZRPC9hZTf6yCvNX3gpu4Ly+Bw2dXeOTGmUaJB/IaRizmrVM
htbUK9NJmg3wPBSKavsgRu2H+gvOr6VWcyYPfYfrG9dlCrVExziR8bHB8KT6mm1h
iKnFj79Tz2ifom/v3RRsu3vSG5peqCxhpt375YLHbCK6xFmLSXzL4t3diUb0eS7l
a9ysJlwbQcUbgXgmLORfjvskqgpS+Ll8tOLkLtEH1iietbCcsKzKglynDIkmqw6/
+ZCYjkidrikBLTIn1nCSAe9T/qCs1fJg+qKkMmbEYcGJsUBRA3QnZj50bSku3OIB
MNxUrTyk0J9wAw9QZVFOhvYOwrbbaF636ltnx1EMBrD4Bp0UPNEtFo2mUaKZBNiw
WyYE+SRQFS8GQS4bAy+5c3Y7Jpq/PuiIQxRsP3MO7XwzP9xlJLlQtAOAcOwqWm0o
8jFL1haJBIxFiKE/jl53KEDVp1tReNgtzxl0b4q3uvRrlg4Md1proBYw97/08YrK
Tvf5deeNdhXpo9yR1aRF5jsi3YNBIZlKnmOOvRw0fDLt37LJ1ieHQmpPUKIQmeiu
tg0hI20bA63I6mK0KiT/7HB8DsWEsVYphJTs10D7hiC9PVyXmmmIJTJsbYhzVdK1
6jZa7j8p1Q2wQIWFILOnH1C+yHxLPs+O/bvPwU1TOx6MsKs8MmA87myulSGI7pNx
/I+0SKCAl7jxE64IQ7O4R+BIVh34xOpXRVIPia10QW0CpMoZIpMK9ioVfgVribpn
w1THDVzGByKtdz0PKz8pDPkIvvPvzqhvGDhfvWxXRkLcFYAew5ATHBKw9Dfldr28
ZKptmMBfBT7K3Lz6v5Sl9s0Kw1p2bDXDyD7j1D2OJZ3XyOvDFC6IvCGlHw5lbuvv
AIX49mkivpMqjDJNAF7oLFlkNeCznxKjhtDSErZLmo/zTcYHwpl2Loxoq19dJky+
hj6s0viMc5gmt8fWnRdqUKrir/PM0Pbeo6yVpYqLO9MeXArZe7hSNRCLfqP8dd2Y
DhcHF7KvQ+c1LP40lG0L3ZgDe0yp7mqYOnO+m8JlEMnq8or13Z6S4gFsDLntY6LB
stN1M5L3kHXsEoA2JGp3X10xHXkK223f3jNHYEuujJYePIygfpVGApTVRXabTuES
fRg6Tg+7CN0WbxhBsLTMB/lNz7gXxR6s03a4O06YH5cwFpx1OYa/IROwDcho2/FX
9jEWb7JNnv7UyqtDTmQcKkpt2qsd00kVaIjSVFAkivQ1E5bJwIR1kt7lIr6jPzOH
7CAITYjEFlHDRJv4iYSEEzkWO8W3ilj9oLtRR6RxkYZywRFUUscBhqvd3/OXCdxs
XDe15ckJ/+hrxHkt0qBBk3UM42uphBGUS8PQtjJIv1tfrgtu8K4rydtYd97d8hph
1d1UGRm/t7MRQOiFQSDghFzZeQ09UthGssQxZb/IMzUBWd3l1q89VM0/AyxoQUIW
ZoV+KptfGBCPFh9t6pJLJgvAWM0njJGHe6lXuIqtXdOg/AFrRwod7xcr0KzxBmcV
HySJbaz87jLDeAb7sGL+9BWlWN+fXIj52rVjBFZcKhqd16eOSWszDvUXeZMMFHtu
UZibPt0S/jAqPN6eqLPTvFulQXpbqQxAC2RG9EgQj01ugw/XpWFJER/7fHg095Ef
QohHeJgAQcIEmkLfCPpiPRlfzgIoLikmA3FgcVX+dTmdFc5F8Y/L1omKbkiPXmSw
di7bZa7qJiJ8zfTDv+jilfGPI9/h9KmEzfjcz+7sGxmZj6zRR+zIJEF7iB/01ssa
ZdDxy3rBZZ+yGmhtJWI6YryZGnlaYfv8XKBUMgPZryUHZQ4oQ5bXwsqr6ZP3rj4u
3H3KNWkxqVumFIBbRFoL2Umcg2CCAt4ZkyGwlnpxN1h29iUuPAdonPz+fldie/Yc
r68uK/dpde1Qe783DHt8CQIaHXwi7S8cwZN9Spcv0pUMtthsqX+hIM2aRpyNWl8f
f7wINNqWZ//vYD99zig9a+b6LiqW2CoCaEBX1n7vppM++jkE2GOn25Xk211xEDYt
NF3fa4B4BdWdwXmEtaeZlJ4v13r2VtOPTTRsGDJx+rn1Sf9PIIw6hmWf5ljrK+cG
1KOCPNC6BJPWc3dE8/ayeVEEd2XDBZS7RZNnB+pdacMLA6QzyiiWPbgSoSJDImaR
SlJEMLfCAzitMpdoUSFQ9NJY/E2PeG4Di4iLYXZ+v3qkIrBfzGbUXahhtdzpJC2f
cW1SFZK7Fd5C11bXFF/XDEHsR9UAHsaIoW40Vvm4YH9/mLgsrYkGYcEOfHf5ITGk
vmjY+elpMjMofzeScAfhamJRAb3fZB+XZ4wox+CD+UDKhib0ZzKGmPkz6j+cazgN
TAAseXkwEGhE7TN4K2GsmbTYQC5mVmbo5gMFXKe98R3z13qUND6AqgEgBxFBgzUo
dHtnZVLUi8AI58zZiI5MZr56sEJiy/eDczhJuTXUsBEcA2xHGWWLmKVwPPspZagp
cKUT6tjRLLVnX9eS6miW7R9IfaDf4R6C++LolgLNXqFWCKj274SN7u3Br4u83fyq
P4LlXbxwvoEps+Z9MsTGUSsXZJXw3cqvAFXzfN4oDZSISXfeRhQpO6zpoWLHamc8
5ha4P6mucFq1Qelbs0iy/MkrZlPH/I22Pc4NrsLCKNk0ZqGh8plWPCaFjzFEEiPt
SjnZbd/x/9yWWcqt/2vOMs6s76hyhLrkje+fdOcxS5rzwgKRHJvvmh2VQP9q3hD/
1XjJacaQUTexWr6231QcdWBQJ8rCN1hWZC5rCNy3bAydnJ8oLEBtuWe0le6pvi1t
H02kLfMuI7s8nOH6sF4AL7YNv4Ij2tAI0IqwdJUuwjBz8whfXlHwS7QiL/VnCs7U
ePuugHCCbWEaOVY9oBeBF8S1Y3KlNeOXCvrI01yy/MPqfbs3M2gi31QYJrZsIcuA
p0i+rAVDaDkI+sCM1jyoBHR8CcurpoYe82uD7L8pQeZXJZxB1LdJw1iLN4qmzleq
0WlMMf9JKi381abQQwHFuRyKw120spUksvg2fkEdqLWXOikpXGrLVIQpOHcBI0mG
3THNR1vsdtCSj4oF+axdFyYlFHBMthd1vLpTNaQ7yBSRPHjI7Eln9U2J84RDQgKv
yhfXedlu2TwcoBC87WjYHcyTLWs8Wr0S0En/y5fPLIjYDAhVQPkLSTC9pmvqZpw7
m2bsT69TSAiLtOdupUg5MZK6YeQajyHh3AJH60CVd1V1Bj2K5kidnO/+tZ+2NOam
s3cUBoz1OI3h/KVKhyfvfNkIw70/+va9D7P4JXd1EQdpKZ6b4aJFkCDQ8zhPpDpN
oRNijpvyKdENsxlovQKzpgDdVrxiFeCyUW1wgtRpudvAqSWS509L/aGHvdd3lLBc
jYoIneq4y3EXhZLsS/+KcpZEdrTAov+Flu+2rIhs+l2xOrjtEYHYFvjNQAfrvMSa
fep8xrZszoCOQNmPQvwGaKcxHjIw6Z4z/MlFhqS5YG9xue46I4uZJShiW1EDievl
vxc0NMzQV7rtuR/FI6+86dVt2Tua7styWHNLYIVIzCCZ4T3NHJXRQthU2HL64dC+
cUv5MmTDohvVs2CaP0l5NJMuvCkEoIMNGLfrZBff1yOuf7eA1tPLQZbOTHkCS6EJ
hqcl/dTyvfKeMPySESInO5uxojz5Q060uctfVfmYPEHX79s4lGYAzMT5Xj4W8nvU
zCkh/xGUUHHLyUyk8jW0AVkROEdXQNhfArLkkuK0fUaPg30aRw2tQJ/XbEPKJ32l
0Vwe3Cp/ybIwliFfIVILs+/6Oru752AXlFZBnwTX/8r6BZZAyk9T9dibk8WJO2iD
NGFsYGKhL5i/Cup39RjloQnPUMeGHDJniHP7K8VEi4pU0LcItedeKOsUtjeuqd2u
IvWNvUDQYZ0fCfezegK3+eysfCLitL4FM8fZFoyxqCfUZKDJxSvJXB/+uspcoqBi
dXCEzzOSBq9jzcUiHO7atqty/gvU4n3o1NS7d0+WAYNoehP8QcIdHU03OYwkVgGi
1EvdZaM5OX1Gt0GPAaItLvn0RTsV0UtD3yQptu//vT+RTUdR/ss3AqJIr3Uwyf1d
CP3c2wEWQWAF0bRY34bXZkpemLEEQL+Q/n+w6oZ4F1Ba67nSpqVq1y5vxIV97au5
GxpQRQ3m1+OLCZhnfQgQtVCV05rp6v81fuF99INMTO/t001tkNHdAf8kuzAJOXwO
24DGDBhaqvUAWti3VEhkqutLWraiOcWtGx54Hotmj70q9UQ2w5BenJLO2ZhVF1iJ
PtI9LfSpQcCNF1/Ap3z9tsvmh/iNpPKR5JT3V7iFtfQ78N0qaJH6lUOon1VqIwyt
20vvp3JhLDcQKJfu9iLfNBFpxy7msxRhXDmjtrpO2m6igYaXapyv92oAyIEYxT6B
GTKXzatI03nH/nSsH0pLuBNXZ8OZJJGDRk3uL9nvDWFdOmq7GeVK3l1pculL7ZAw
M33sMO+ynHnb7vtAIP/QtaDOiHEUmSRFXxoDL/aKwf9z1DRV5irUYCJDWEggvTV1
t7DZEVDWafNFMaKrqLYaMqNeVcX9iziX64N4dYI3oTWyTsA8tx/9ZVRIB60FAHIx
zCxF2Jzzky1LptSpobHuthJAaCItp/Uav/ZOjQHGVhwVmni4RdKq0iWyuVlzi5Qu
ZPyaQ+/TJQp/TnYgFRtf0y6mvYyJbyhuy1rowCxB9rj7OFKJwyn534MjVZBzSCjU
4o0LXUkCtXn0pW90ZX2po1iiy2VWoE60BTV697re24zo5Th9AWVBtw5muT6dNtwS
VJFg+ORcJXGj7vycwxCcg6Q0cevRzEc4M9rcHec9vdkfplMIugVEGjQAaVZ18mdo
xZ5d9YUbmEsB0FH/Th+CBK6SDnfbCRgBUnUhFH+NS2qNkVFuKgzhJIzVM8q9A9jI
zgY8iPxXpFMpEHzCfWjxXTj5JNf4MAQOYSH95HJuwgczxWpc3uY2HLMODWHbC9qt
BA7TbpsI4HJBlh0d6XUEmXyJNTWGjLmukxQetxyuXjPgdOJrYOUVoOSjarVn3eRd
pOeDX/a8ZFCTM0V4pID7cOiy3E6Ji/N83jY8IspLkrx3xm7fIKS9VjSVa0PggUwH
d3/o3wGHPYkmf4HPJEAVL/j1UwsfvGidb15Kry4CI3ljKIhu1R41jQnTVt6EMwNl
UgM3r2LnUCQ9XQpejl9H8egpGNPxhiwLIEJam5Sr7iJcxiWSNeWdyV7nzsAHxPdy
zR8Fj6AjS10vtbY+WsSjTBeyN2orC8KFzheoNXd/iyhgSdOkCXq7XPW5wMeuROs8
lQgC5AsTgWH9ECSVsg5693/7Th1TygREVZ3ZAN7AN42lUKc600KIasKhARpsQZRh
UtFESJsht9BvDxhInUuJdvIWz2lORprGB25TvgLyEouezH9zYiDFPkRIz3HthMWB
ijSvaLgx76jDVRaqei9c4CUeuwlOkx1vUvcCth0v2rOEua937XUCw9nRtmatnGnf
5kX2hxcq2ZTXyrJSt5FQt5nk3Bu6VTfRrtpT/32oZUZCT5AEQly7XkHgzFh4DbO0
V7R/9iidZVs+K3juyyFoDoMF3LpawRsaLfWZiDCrP0Td5FjNJKptC2Os1ITAPrkb
fzntOeAk2a9yhW2ns6hSba57aNTXO+H9O5hFVnusJl4IphTzgkXXmgp1VWUqUc/O
D7n86F7I0MT+E8t1d++eQwNXl8J31XIFKpb0zRZN2e9sWR+o1sDAbrHwVnbuc81P
M9fE37zEm24/Cm19oXMXhmWMDNXn3nyLVh2iJrwwtx1SyUtsvW3obf07S9YHi2b5
FHJbsNA9tzyrR6+IIb9h2c7OmRGqGyxUQoVBA0U/483VcfYqDkkLR8WX8RybDsdd
q/PjjgJn5+EyFfBZK8R2PHsQuXDRFRhXeZ9O5ihnfM3OQ/MI6ujtHJEmKwRuXV6L
0AhJ+FI/3NreXanYgpio76gD9nbjPEroyEma47rp0G8TlWhy7r5lbuyARAM3RQsX
CDZPyLd35FcfwKuBrpYKF6Cm9lNGd8qiaFYpQ/irpcyVSy+takmGhs8ER7OavIEx
UiZp94zDOdrsv2d0VfIIDy9DVl1MIWP8E8SdJlMyNXian4pSAlkS4D/dgUrCz5ZY
l2rZK1Rx33rAAmC+u0yh2LzM2PbQvyBAru1PEMMmJt2FQ/HBJroiURJ44ZFLT5hI
m3UdfHTiEMnVhevGJhQhNGiD5kB4bmBXenGGZ6fycH+eR8vVWLLoOgn3sDXl8U5A
8In3+E8BcgnqiuEce0rENml9MHRcSAMdsA/XSZMvuIhyv8BsRl2SqeUjci9zYE/s
fEzSMr2G2jkxC+1SOVudOud1UvSv0oq4S43xCdx32zcG9Cm2arKimM5IthCcIIwR
uL7QY/7SD1kCDqHybILc5KyYK9e2KKglpd3Q5N5TMs9+hHiFw7vLgUMirB5xts9x
Ff+mKj8QmRiD45oTdukA/8lLDQvOBeGQb6dzLVAE6wRzmrhpX4i6gXM3cEBOjFdP
97mEH5lpq1kwmAa8p01e+T5KdAWWXSA7xZ2LE9Z0Uowupt5qCqwWaIrUR3ivhKzf
rDy2F0iINKt9/FL5LuqcxQClYXJQ9Qp5kdW+uYwshdsYYRzefOoUXNar/05SHHGe
OrxaRNLgWzZWOLTxVSBIZh0QlqU3Bt2ykCMslnmOQqeroy+jsZPiELbLAIwvt0pg
p1HFDuDGfJPUK4FG+X4e55ICy2iZTe3o99B9f02aPf0UjP9Utx02G7FWNXS6Vuc9
dfhIoV2DW22U1itt9zHe5/AE/yFhbTfmjmzvZKlH/lUZeHmwQpYuzPvSUrqgP8xr
fCL87WkI2npH31VQSF4Y6ulapPaXpReDjzN11YRw8j8dnEXH99iTTZ9EGDRefAGw
iCgtyBkVpOesG3htd4pY3Z9S93Cj5TrJ51tKU7OGFH8z6VHCpYqYfJZWHxbkkszA
DorvBvb3oNvDwb0uM2kiYfPMSjwBsp/kNM7kbki2dRaID5dP2zjJfHHd+WAtR3+h
6gDexMC2dzly+fgVHazSnqog9NVHhXlDNY5vBLu/2oFsAYakbsyhiYcSZnMAeUKm
niX9X9c6cxcSheqt6oaHsshSWq31KZmxwSGwEO+mqpp4WH0ho5I2rFtLXr45RmB2
NsaodxKoKFblBc7p+wY1eaby/LpeaSb6jPDgEZTs0lZ4UBrJgrb6MLA32V99h0kH
19MjX8F0ynB0trGNo05z6wxrVa8xE4ghxcxj6lNda+htaBPOnhBU2ytx06bvDW63
SUHcNfZSYFgM6EEhCYtxt48qm33A0REhLCzOMd8pCswLfduBbaUALEeJ6BtJBFTG
WGyYuXuIXBl9YKNfxRuAhq7r+gt/BZbFPz2IebqUzdRzOaaaQV7ZKt4F0GHJvEcY
dAbIboGh6hFEYJFOhpb+LELuoel/fE5pHq/GmtD/cnvQMNgr5azox/rmDATnAWnk
A0CXbcVK8IMpfTzCBL2b19VokdtbCPwUhYTDonro2nsCTTUSU1RPBW0YYceOt97b
OngXu6phAcRdDvJGIw/O1nsiFPDol3WIGve7IXncBRxgAzfYMoSfa+CDB8GOCDR8
tyE5P1eGscHd8VulVghY8e6DBWuXhNasf+zgn0ANkiwh1i07kzyZRtBJyXlmNnEy
TVQldZEEZWHBMDT/fCZ+gai8Fvlq39em596PSGD7wMyAxwL42XSfYmo+kft+W59g
T5fLG/pSsDnG62zjQyIJ4gbPcTXdMzBmHbB6zhayTAmRJk27SwwcJNPJpDtONbEI
6hoTUzVhhchZdMkq3MfVT2lxrZAHuixeqX+tRjt2K0mODGcnFDqRVTaC9/UzozBs
pONoh19ClVRIcduOhzWLI55b9gTNYlJA0rUfyYbQ4GTGsvHi5pGlFX+syCXdKdMW
3Dyh8vYGj0oCLvmWQkUriIulc8MnafyNySmaKjpeEl2E+/D/E1/qLtMoYsB7FVAL
/3gLMtcai8FB41RUh9AdkoOgugbOieNTuQQ0Wy+3tGkHTIyeSwuHmvB6wbLWu6Jg
enemmYg20rWQdrPwmXpZ61iw2NKcJRt60DF/PDF7Ilg941txrDJiU9TV6Br1koxr
Iy/B/kEl9NX410KhmmaARArgYb1x0vd5qFOyPvJRYP5COf4dY3O4Fsb0GK896Urw
YU/b2CdLFrzvnHHVJH/vWsHTsqnsy/RWC6l6slBpx9rj2Q8Nu/lBZbgO0u3yVbkY
xKaheYoZNNq8fQf+5xu4QgnKixil50cs7IKEu2r2/UaMin4H79/AwG37dxEIJga4
Kz+XnBuqE5jkkKWsUdQPNMnpuAkYpjKOdPoZhl4Wo817D2DfSdNwX59kvQ7Ck+7v
AeQaW9CT4Bn3LYv7rHeGonhzY4fV9QzBkm3m+c7s/WF8hLDM90y/vOnmxB1KHHlA
f8v6J4O/O8uQ6a2gwlpx2duj6XxAC6T0SUy7zncfjOo9evony9h74jdNb64R3VUx
BrG+MEu9QnEzEIu/daefap+PTY/F3ww3CGCiuzCDGnvU2i9Msg/dKK5Qtx3Dzg9r
MxOwihxAIsWoz+LH/4DC2jec5h+ZLE+hxs1iGo29kIn6xnmOsTa5/OVXMbrv7vNM
QDGg1eeMA+/C/ygq1OxoXENDn8bweNVxbIXUkprB+06PcG2XcxsvlDF+wqLwn7Ej
gdVgTHZNLXKaLpD3/OVB35/bjnZXfyFaeVrkYM8B58haJGVfqM2UddCr+s31/VTF
2SJRxolL9HlHXTTQeNWgiJ04Zg29bDniZklrh0QS26+yQV8/eYtmMlg7QMh/Fo/9
S7W0bveyfoyA24F+CsYRPl8bhAm0DRrx7KH3DGJl5PQGORVtTWEEsouRU5vCiZoy
RFhMZhmR7NjN2GO9gx+WrAI+3LSrSplJfGi9V/3YuX/tKQcpGWNaj8Ir2e4Y08Pk
GciWZt1O3XpaYZ7uhdMWCDa1Rz1wcDJQlh8WHG2eGOhHTfKdxqX5M3jMrzFyKq5F
G2bXwvzAULwUNpS3nQprA/8tQuXX+vplZx9jj4/Nss850V+9kJkbY+MafoePr/aD
ZLG5Xhn9Ry8/I3tot+3st/mO8nXosbk9J1L7mbwxzMt1ixKeoe/VajC/3/Z+jhhG
gMR0OsxGH+fP4Dugy6qfg8Vx9eU++tn8EEGTX1yqPM+KVoMsiX35HMU46mlf/5V+
VO1BQUZVw+HQBbNVPewPiJw+aj14daMCtuG97SnLqXz59WxKHv8LwGgbcUQ6pOTr
F8Rn4ZwOCvTjwOBWLb8D41271mg/4Ag+O7YbeXbAXdWPuVOwY8JYnAK8iwRiPBea
ZUv97WzRdt8EDoN/xbL1AVNtFkLRljtTk6xP3RcI3tDkMG2GgBmQUW8by3ZYZ8eD
BA11phZovuY/xffrLAnQcegSFT1+uZhnyEHa0TfDUwoqsNpiAnmh7fxvOVK8qOgf
8v3nwgfme7SLavzTSS1CCAkh2YNpWug92TwKVsmI76VvgSAdhuOTTdqKcrzi7aRl
nuH7ypcR4nAphHAbGW9z5DwnfvmkIXDowett/FWjLd9p+noQz1ewrG91nM/i2eJH
q3GlKN3KUA+YCxyCyrZu4WxXW2sIa74pOniz8WPj+2j7kgo9+I3z5uMHHDx6QjN+
E/OLTycgZHYXiiYASakxUuPx/2wWyN2wciMyltA3rIUBvp0QhADod+C/0Yk0IDQz
WCsdzvINGmCn0ejMLVJwdwH/FXoKYdnPi+uUjr91j+/CK4mUXLUq2VSHXeGgcJ/K
hGuNOSZ6RvMcj37WO2DI5oH74+/6B2n7VFvI0QTK31xUowkmYVvESV9ZP6fzEfQQ
DmgJdRMJL4Mp3+kBUp5IzAjvi6DAIL2d4biCqcxDFFAkcJJfuH8OUL9i4hNtYxBl
RqMu8RvCsa2nmfL7YHDm81mXwIR1x1GIpyYzkccS+JF0iGEXc2eZNV7XFwXqVoWx
i9XzGbWdMSBfyxxstzzW6kWnoUYaxcDz+VtWDk9yIISpW+5lHcIfQH/XtIUejtW8
WoZ9wIYf1hTdA5Uo+WO2KOTutEL4nTFGIEwS9YlOl3/iGDlPLL3c8rX2sup8/7Sm
e/8iyFA0dVz0e34p5EmExYMu3MCSMNSu7+erBqeMb4Tcc2h9YkG4O8gG09KhH7xF
oE/EbLec6Ig5OWTQRTYqRpoIYHOd75fUSOkzX7bnUR+V0C1c8bTanoLpXdSy270j
Dg3JTkG/cNQXI+vGym02wDPqT5xrRANcBU1i3fRZEQAFdbt6kyC/4201+SjjbO4T
atjFdvCOk7ov5TLmoVKYb3Dr3J4CY4V1pjyzAmBhUonw3q3+ooX340aYNHFqHttW
Zta1MNYEZSq2UKGO8ocDBfU5kUkB2lpfEEAp1Qey+p4cbwka4yz/+adSJ1pms6OH
H+x/4+G+Idb69hMmr3L9DIFhu3jfDIbecsxfOQv54XCvgkybrsYdxEP5fbTVjliF
rTvrOdEKNFGgzYyiioUpzJdtUEQKFYc5F79TwzKC4jWVvmCo+ykw/Bg2Ec8TD0hJ
CZ/m0ta96mpJIWFbcxYjQJJS5cn5oyLk4TOtjaab2mDsAZXbQM4rewuqpvwoWJcN
cLNJfwyL190r21M9vLDHW1scHMzceS7LiRyMYrPQirUawLY3z6KmGqoEmh1gm4cz
bChSe3VEQ2QNkd2+7tVPyA2tUGR3PHUj87xNLuwr2FHDQn1whRZ41PINj6vLi95g
fRm7vXGilNvA47LpkhCsa0se+Qe7ho653tfYyp3DAG1pbfKLD51FgtsegEourBFK
KWBrh1f0dPmn0/kM2aFBMeS51zvqJhUugXgR/u9hszOcfuZy5RGdaN2PMDqiZle+
sOjCXOYzwFECxe1frCOWSxH8uI1Kw9RQC6Fka5EURLZ3wf/DC473toBo0ekNeKZa
9RRj/5KDGoWzl7DwperuQOI/F2L6+CzipNWu6LwWMs/nffJSoslBC/K7dnEmGqnv
3dLUJxmAWMbwxn5NHTmKXwltxCGEBgC7hdQL5iIBTcVXYNR6ZFUPqbAQfuTlEyZP
Zxb4KdiB3fsR/5P7Hg0WkAdtAQB5/T/23FbperKTDWzNvOgkNxX4L5nDIPgWnf+F
k4A547lf3HGBsnKRIewlZSxxLH8xW/5BqtaunDygPyJMnhfMio77/C+R2HqKUqQb
j08GkwJDhBexrobMzphkQ7NJj6v+G9oc9MrQ6xdUY45U/YkSQ0sZoib+naXH8nAz
GR5FRR4Gpgzt3VAwrqLtSSitCsXQdMlxqceZBwB1/RI0yg3Zb7UP6tqiiz39THJ2
RBWed3UGbt5MVs4icJUwQHmbLpUnG/krOtFRm1WA2cpVoXcbkVihWeoC6/+P9fKl
khYmjoWtnsQJbfLg4ddqQQDzaerGu+t5Fvbtg/GPRyFRkT5DNcJr66xmGPxaL8c1
0rq20ZpVpXzuB1oPearb0w5S75SiW8LfcPg/GI0RZ/wcQVNfRUkAjn0r8WNf5/ft
QXNZBOcyU21x0xMqqFrCOASg8SYSUCbdPlFaFD4o/psLL+g8YHkHLYnlPNZx0try
PWC0IFT2oE5TcTLHgVpcZZoqpvNKPjct+meulZJOsoYv6cvo2xT1NrSH9CUhFBMS
sr60BlbcuTLNLnCc+9Qgq1hqfLkiaRNiM7QDpgogniAelm1Vu3efMv0sfND+kgLz
AuyAGd8e6WAFqblOXI/QXuElSYmOYzATwYWMBOrxmORUOFeMXzUFRgTupth5e5Jr
Wt4raanF6pGUx6KFtFV6wBtRGzFQRYXufK0QKQaWG3vSRNyDHpw0MB0m7ZERI51C
ifeHuRjuEDK3XQ5FE/7Mly8ykpRQ7TAzOZF7r+i2QRh8rDcNlU01mVVJEdO0N8Wm
LgYDBie4eUyLi6juv6kIA+aEH3vE/yKevekSl/JolA1w36dXlp7NEs5Qtyrd9TKv
276ETK1feTUJVA6+W24UeftEOxlTHItLFcHCOAuvMIKsVNBMSnAQ3uVJxd6884Aa
Lpk6zpW0J709B1/MvFrBhyWRAt+pfHbbW59RGMQspdMZQwkC0GP3XgSsgMLLaW9v
ouCQBLo7mD0CY2L6t2YdFZqgwMFX/4cpM/A/6UjqwW1cZpEui5axgGnkqfBztQ0q
v9U+Pc+CubKgps6LJdBnitAQFSJ7HDCTMrXqn41jsOs0fclwNpwDOcfTKTu94CDf
AW6R8djebBtlEZQHmhiTihLgvIq1mXLxEUh5dl4tDfN7T6Y+fhxQ+QFe2AHawoKl
kPr8oNY+y417r2dL7nFsxSQ7/WWlawglFN8KogxYIqu4QDpMiRRuHEB4F+k0b7WP
eg55+rNspw+4gIR4oUaICrSTTt7hAQSmZFLTSakXRS58UeOU0Slpkj4W53iM+2aA
gyBkYER/omBgxUCEW1GW4yvQGxVIhmXCPzM7XiGhBdn+Jfk8/q8+fWU29SJskohb
x9+CLP6hzcUPvvq3Zu3by1Tqjxu7hdOiAmaVgtH59PdybJu+uPrSJltjwY/wh2QQ
vlV1heNA7PsWel2u31vrbyj3tJfTgj9/hiMiH4kMwAWoi/755BSGMT3TCmYMybis
ANTCn1yap10IhE5F9q75tsOlQE8acPZAEWztMPYytBTbbkGm3fZLje28fwdnUM57
Z0t2fRp2sRHxV6LBbL9+WpNLkEUuXnNpCjSwiSOQCLiugHdVg+RU4I0OSXgG7/xn
++WY0ojS/3PBGZO0Hu3xjJPguQdpENfQKWWbE7gv0+9DtZbHBjKZ2YflMIhZ+qnv
CB7Pw24kzGUSjz2DVtRQgTq/pulkuGhHJYBGHzEK58/2p7SNCb13xLcCFqrZVSwN
A8ik+nR9RGkRpAkpVDXESc+A1nSY3Rp1z5t2BKvIT1oYDg7YflKBmMN4KTqhetzl
skNkK/DD3dOlR6kftPBJ5Mxhy8+vhqLZhrsJkgcXnSEwHbsDABgrGwXs5VmeRzqK
wC8khiRqhtSMB4zL1mjyFpEkIXGl10kOpwOiUMQc0St+vC2XpwxVWtGnTbKasbkE
iBLPd17I4BxsHK9IzZLCOttAn3K9tbicne81IOQJqCgw78F7G6zOYbWpNo6rzzFw
qSeZ6WwHfODRCPvY9tHDbpbV3+G7csz3x2QJI4YbYRp6t4Fse+xVbHKF8J+P1Qtt
Nldqw9nIMeXs7PePhDSyIqry7dUKaJJCLUYSiQSPheXaZHZ88PZSMxbqCoLl3J7G
ewBbcOda1qI6Q9kxU1s2R2/qGM/8eJY6WERxUzEDu94RfinoVNqynuULw3KHJSPi
lsPiPvCWln+MyZBDq2YtZS0hqXkpvC9EPXZWhB/ONb3DI/+SFEhZ7WIuPXFWltys
O/Jr5MDQwpF6VrEMXLgHtDJHkB9wciBR5LwKpt+eWVAoEmwvpuQLwYKvTGj3TK8A
oa4LFroEkHIui+L/SgeKj6uu7cj0Z0jEavL9LhVI8RnfucVyW35dW2oGI6agSeAP
miTtE9JYEmrGBpQ7l7bKSpo1eK1mZtZDgejkNSqUaQszH/W41tayzKw7siyQdMrr
YGnzIGUMVmArOgoNFr36jfmUhdT46rlcGwsqM2z721Vmf2p+Vnnx4NN+4kvXx72s
UBV2Gh2GJRhSgF+2xavUW13yP2rzWAFZUkyE9XnLoTX6Q+PldiZNpUzsnyPD4emb
7yHd02cBKvbh3NKNcFFQzYAXImIuav7VWusfHwgqRu674+HH74ZM61vEwXy9XKhA
PpJj9ec/CJSkYGVtpugKnUZL1Qvtjst96qp9bt4R7YfI8ixlmIeIX3+iXztbFSkb
7VfVT1wm5CZ6vtF9O3PZhHPI6BRUD7eQQmykOyAdr+idHGLu5950W9jzVJWd+kSp
QX49ymVVMQ4RwXnw7pdcdw5cL2DVkn5Aixik7hsO2kJayouZUvBjQvSU4yNVeLMJ
Nbie59pUpUFGp3dRGKbJ2J2+lUhwTIsSJhayLjAf5mwcFcNo9lU9yGxAjqpvn4/f
lqRkPqJvVpc6XifWgVgbMDuZFfJgsUBH+v3CeNtZYpe/Q9zFT5JBi3Poz/M7fHxy
qIikxGejPQhEM8fiEE1NsWCHJILdV+RFlFL0Q8PyXrV02gUCLt+wEgzvYnxtdCJ4
rezpgBOqgHwt5ZZtHQ8Rz1KfdXecOTeK1VhwHf3TgKxZTq9Myi83bbOqalPh72d6
O6llqR8uxUOyCahQ7awyJJZl1/HSJ6lrCiOTqqy5f9LvmCzDo6kPDkhIx0pwzG/t
B79XkHJ4Yuqq9axGjQRMrGY1HuSIHHMDkhCBVHZI6iG5Nyd2A64z7VllhIzK7zCM
pMGFSXocGmu1tzskf0ctim1cSZtma77bVD7307cWmbP9Yl95RNqFa0i4d8jNxkCG
JeM6L4/C7VXUnopvHofplT/AnuTp4eXnrPPBWKKqhJnsC57H6E5ap6EUidpClHHk
F279Luem+bHUzeS/U46MFBmW9BQ/hJHn4q2Z1sxpyYd2EQ4bUWN+sXZmi0iUsfr7
DSF8RZfBQynseaqys6ZuOWQEve/o7YKw78hi4jaL3D2asucxNo8BUvP1SabBznqr
wBjUfHtq78Rh7Q1xf5JhGYF3Lhg3b8GsWqAd5A6bDFRo7n4LbYMJraDm3GWHVuJN
KHM4HmV1VKvvgbCH/aIU/FwoU/ADfynvRXjUPmoyG3OEPQOEPxWDxMgEPF3d3AcQ
Rl2YTlORPTW5LzZiL262uTgZNzBAm3jpr07UbiTCnz6H6aalE6BfEclQNeauabjE
9z8RQcUAuwwREAwInZQxwg+Kh57pHB5h6Sa6zgFUgaqlGTi8a9+VdqeZKKUMdCmE
rgB4vj2Ewl3R3UINN6tBb6UEjwqDO54pYKo7jAk02Le2MJRnJXRbVJzZsi7zxovi
fjlqQFb5QNTmWeA7FoVfdR4H46eFovKM+n0C63I7pGPxUJd9i9zV8zdEK5TunAXl
WZJTtyeJQg4u5nAxnHmyA0xTn5FlWVQtLNRYCFSZDBdYWJgrqr7uKaurGoodt+rI
2JSAaoQ5N9MKpzCDnPd2KQBE+D7IaxfG1gwoV3pulTgmr9u/4dGP/OdAd5xlNCM1
tXOF/KqO8Bk7uFVHG5/BuxCn/l07q1fi72K+3VuyLk7f/leZe1WAMtHhnYeSeeta
c7PGrSmxJmIV8EW+X07ARDaY0xO3haDtDW1rLh/OMKiuVE+PuTPfSR4DHQ3DR7DU
H7hg55yBPwT64f+s6igLIk/UxerGOPTEVJzQmwU2hNc2hth1HPNqy2Br3KklON8C
TCQfgwohk1dBSGFUsdPZKc8w2aXXyAHg0k4e6O52eyYtwJYF3Nui21zGqrjo/ccP
oVsi+Uqo/oOuhnZsQ0+CnNs/gGKjhI0T0a+YUd8YU6l8n5AA3cajup/XffUgfTZN
ugbnaRZHQG6KZgd40Hy7c5nLABQfSX2pdLy9NQWx/7Qyf4cf6BoW3sIpUT0lhInk
aSit1g59nw7vx9gt49PMJCm9+fiCTKKVz1UBq4Sz++1jt84DtaCEjZQkXOdSayP4
XPr0eROtbsYnoTUvB/wUuxSmKiXJ0WeA5Nd1hHWwAP1il7CfqPGaACFcbnOfSjdq
NypTAsHAuZkN5B/2Cz+VQmomE9H8wRWkksV1RyxNmdUueVkMO8PsfQmbMZR/akMA
89yCjzRd43xyXW5sZ3QLsRXiKk0KCSpCXMXhw+Os+g9JC06H0shqxPVVptYATahx
thb2wgAzuH4tkuAeHj9ZYOj/uLXzQxohzFBTKaIaMUzsgzw+kjSTi5iSr5JPyno8
OoVKgEeCBmdQy3sE/PjnrcSaGCY1XFkZUgA0Kj1/Xb1FnaSPdv8nQLD/x512E3bF
UA0pCBglB1aDffPiEHR3wLFZXehQNQMS5vnMkUMTU7x8G/NZCmLDZHPxz6eq+qB7
jHSxExCHmKlMDDk/FFUX5mgAM730e5HmFHDLd+3QiK3GdXnfraOa/BWknZqERXcz
qbGKxKhAgMGZBzGpfqblNqsR9hIqopy8cA2adKQMBiXdFrvgAVOoRNXaKTlgWXOE
QZyY19qcaRmZVeNwb7lO+/FAajRd6iv8kqAc/2ssUoPfJ7oddyhMJ2oBDSQ4CFs7
c2fREBMGca1AkLmsLdfUNTFuGKz5bNMKK3KQ320uffbxH0uW7xxFVBbpIpSFxBnU
6cYHFpDV8NfIhJXCfQ4n5ahSYdvoLd+TPqoqaeWSoktGLUE4pakHsPJaZD+mdfig
xw8mY96sAiMPnUADM+qX19+vGqY5hM3wnwYtRBcm49fRS6X+LnjIQZxNHfCB5fOv
TO6YkvZytoaCYD0iAB7rUwmixaLVceIgarWGTo7JeVNwTLZi3oiQe8WiWd5uVWjT
ldU6PkvwIFzKLuNF5EeupF/qtSHxlvzyHm4QfX0qZhIF59W/jjSE+J25VxwhzInJ
82+es3IHletOV/vo9q7OQR7sL8zNlg0zIC5ywDC3CxIJuBbD5L7y8NyPGa7FeNY3
EqMsDOydRbp0qO/6iRS4HUuX7JpoaidrUS+JOuwT1bK3/WzV/LmHmk+5Qgi6YzIo
5yC7pNSPvjzQorIafmoqF07zBdVpEugO9Cy4AIrHS4Fnj+/PP6q7XnOm1+pHr5vR
S/w78/WTpeg26Cm2wPmgkb6X8sNc/5VFbqEoAknYzYkqNiIxxnV/MihNS6lBHx3W
e3wrTNHCyvL1bKE8hPR1k8Dvw7cwIG7d29y4ZtEZUZJ2yM8dgrekusNtRixT10UR
xZaJsEEVYGDwGkkZPyZaqyuo3AqnvtTBXs+XbSLpYK/eGTCX4HZEYySOxf7GOSqu
Yby18Bww0aWSTJUUzftIFoDfczfXPfnx17M/lZMMqwy2LqvGCZ9/SFKd8kkYfM7B
bAFlwZGPA3yD9sFGq+v3ttbkIy8izwhSrOhVcUYl7/qdN6a332nhyO9oaANtFBP9
X5lg2V6doijky4HZQ2ajLYCpF6/QT5Dx1sNp9Q33T/LRvLOE3nskqXVtLjUqtSmF
vfFJpJFJPRQS0FkSygBvWdds0h0oayOSXvEcUx4i5RPgid2GDTddwv0EBeGMJzzX
hNOjTTdgQP2S5zVd/hZReWBMgR+kGS9lbetvTwZNTtMzKJwnYsmS+1tolXMuvpXd
Tof+PMzKVstHq6GAK8RKiiMfunwp0gew7NifSeGnUc/zbqfRAxFJPQViSAtLT1AO
rvQ3oYOXcFWUz1QgyekBw9wW5hvckqQLzHAite3zjOqe7zSf4S6/2AhkRSFpV2Sg
mzHfLIpsI/i1bSDY5P29JTYJDKp4SbmkTlQu3uIpjvW7CiAtme1dO0AwPn/HDRZY
D1Rg3t9KlNvffLCsgrwizp/26kU0QNKsAKsVagx/UDNoVeJofH9RgbbJRl998lRO
zzsXcDh7kT+RVx/MF4q0uH8U3Ms61UEtPPhLUnq8pZfX4IXPP8AoEmxWBCNeVqhX
NoNdwDdINDxlSK1m1jIs1SBzbUt3b+VRLb7ok8BF+xcy8/X7+4UBY/Eenp/ZTzwc
GcqpRmvcBumpJ4bfyytKl8p3OrL8gyc6Zn/r53jSGcbrQuJKb7iqTnmCU/Ws4Llh
yHLBljjILw2fao9JUYaRqI8VTVVW+Cd+5I/mZOjFtrh/x/ofr8HNvgnWGsCt24C7
FTTSMJAoQQv71C7hDS9tNtfkTz5LVzb7Xkzqm1iZUJD1ps5dEPoXftKB6YC9Pm4R
nNOD3HxhDbt0L5T1BtW/mEOEHtmVYIC3MEIZEdbMFwRJzGW9G/2AqnSMHikxPDA1
KMXVW1uUxfXkC/9Y9HtzRg6tQ5Et3ZrF5/fOOf/Vyfl5+ACu1qnTmc3SjgW02DLR
75k2DV0oi4mHrWSChCH25o6ihBS8398QM406lHQL1RtBPXEDmJIq1VE+qQiEacDp
1oGeCD+1j8zMjr/huvTka1ttdahiqAaJyjWTW32DAZwSRnvrV6kvKO5ukDn0oR/e
y+JjRetGdF1V7CJiIi2HaXCskzUViL4pD4FHEVCeuWyp+GT6788XVHpU97lUGoNE
3SR76KNT40M3bhCNu5EhGI+4efg5kIO/9T/ai7KPX2qfx4XzUioFlPhyw38vpDd3
Cuy73lryns92c0OcOxp+oZr5OwhWKp/Tf1fe1GCIUyCEU/EMe+3UoAsajQxNOq1P
sv4mF+enN10UGm1Twrpm3L9ehelnvgGMi/SHfO+4Uq2KuKGWLsxGdwnRa0mocBFo
GwZH9msAIUxg0ZChloeqlHrxcktRm3rERXCKuUd5oKbsH1cGG7djZrP8mqPHuFcP
bCM4g8SQVV1CfMzxsZWC6YN+pxAFBDAXTOwGCb6NuEbY7blYCETCftd+Wm83Tki0
SmWemno6/ztF5M+RpC3vOCLUsszJtwz++R0EPqnh0oDXLvGUucn25J2/sEpIW3W9
bMxXq52vd0Ee2Ovax1EMboQ7lENM0eub2N6eZ9dYABFXrzSAc+r9MkeOox3QpTOx
kcevLQD193PMB/Nm7diO7VkGrJc0Xw5LNaA1k5C/ebtWGMFhxcrfL3EPBDILP+BT
3vXe94sMJ2lhzYLuLcTvO32mcOwEoJcg/egMoSdbV0oCYngFuzVSTJ9DdrsOVbd0
tMr7tMeAfbsLYQWn1Pt8uScQRfHYOFgQPrLdQs5EbALOV0tPoLRLtih1ZSCen7pX
iYnVmDd2UtbwjqDRFgnIc5orY8Xw1akUrZEzX7QqzfZHp8G3Zjkierxm/wtXqZgD
X3qcuQMTJAXlC6h3PWedpfgzhvZa6zSBIVJVzBixKx7ttRZyhA+WmWSLdombl3gE
vKbOTFI2KYtcxhB9c9S9uk00tWwrQJbtEP2l3R4+1BfVVhlLXFH/tpa/27Vq6jhL
kXcjxapEWKf+iJqJxtGDwPd5q4Jzmcqwsded7QKmPF6p+p0rxlZQLSojiAXXN9F4
mMS04Ueqf1bITQ3xBRfIA1LNWxgKyvTf15jSbrZLE8wi0ximINH8JGu2Ki7ZB90e
M4Ho3TE8cGUvVnKGW323XeyTvMbBNgUWiMC1KrEPz6KHfHLE9DIwx4Xf1ZMeF2K6
g63hlAeQvDhrIWNLWWLgYMUXT999OOX/D9KXEGXMQFktyczjjbiTl+ktmddO1hLQ
MbVVnzTavyNdeocl29Zrn43mp2GhG8dHPWjrMNH+bi6aYqkd+981AwRq+wW7i2jD
XpzLSc1gChbNSBBfdQMY2PEBul/XmESlU6cxQyQtdos+Kt4qz+zjZ/Y4lNIrxUHO
SsXQ4nzkecKPDrTmeQ6XGqLvaDUcVJN3TQ84jMOJoNTbT6WnzoaYgBdQMn7dhEtC
ddsd2uSAwUjPYTlRC3bssYcwtPsiE/zGKzWZIdcaAYuY+DuP0SqJAgp6I9c+Ef8U
N+xRUCxgcfOQd3nQsk5m/wXbAUS4oYoMxAlmTrcwA2NER2Wgy/bbK9yCScW1Z+Zt
5jeVs5tzmpZhAZ3YjAuem0HkGnKlT1zeF8MZaa4GDCe55JRuIe7hVG0u4uTA0K8Z
fXpUMscWa0usdbxFLGeaH7X6jrIjCQP798L4bC+6yznuytBxIxsMOUTtzDZLdS9C
t+/kbpi/yBOBXDsjbqyExnOcUo8JC0WX52Bmemd+YIz8eyEnc0CcQfXeo23bEZZQ
MbXgEcFC2dVz/j20L30kJs3AMBF7acaSO80fW3QplHPiUI9pzJKN1Q9X2Df0NVso
y6HhFVSHUP41cro6SGDi1a511fc2wOYcYLmRVbh36lghAH702uKAMeQmLkY3rwBh
9ioVLGeadis2R5MDILtjVEU7Sow0LOinlJKggv8UQje3kUDRcvoj5Wz6RhPH+M8k
pbNyS6ALVBY4z8GrbEtNTIWGNyDb+gVJ3ikqA/0oLKwVDnS0tHZcMdqRAp7dX38I
Jf+zxQOUap/8OmDll71PW1Jhn1JwKuS4RDw74HKw+YDlmp6NI/Ju2e0YMrsaoQOH
MJcSUz6RWqIr175Ly7mRTolWXFo3RrGVyYmAFowhsNBPITqGYHioA9BVWJ4A5Qos
VCyY7+gQEP42WtNzLagcaJg/ap8bsFcwZuRXt302dY9wudd+gj8g8ZfkNBMu0xCD
nKJlK3hjnV+vRkVsYImqcXfx3VbmdQ0pT+0pYaRCEyYTLo8ZpWZmyZcpx3LvKbeR
dKPgy3NVSnhim2JuTWFCAxlcQVdGF+9iOUTmyNQqkUiBWT+uu5QFwvqlntSPTSda
PNK+bPTv0jReAARVuQEZpIjGWz4v+tgKafpwpSZSZFiGy6d5I+qaEoPV9I1Sfe9I
Sw2h3CQemPQ5tPX8uXDCpGyhA5dVR1ARBemVP8LOREL8tKaErJaNlA6mEJsH/wl1
psBthBLQVLAjjday6qEX1QYpbTOWjUL4gWHvs5l6v3yBAYxBWhoNanjH2BqwYi5G
YZgPBu35ZybXZ30Wp4sdaSqZYP6NRURAAQm4w6624DMW4KRLrH4DG3I8itGUjz+g
9I64M4VTMNCDA3bgjDCaJcf3SndGW0H0aGtihSnzTjzAhicXNw3PZbB0HW9acKl5
z3OyDZ2KlbXWPIsOVVM9FvgTy1Mas9H1xsmetAP7kHohhlEWhpnoQM0Vte7//zHk
SPnk9s+I0El1ZbwuPt1EnceMXZ8JXB4eySzvY7dqwSUVTeoB1LNaCZyksSfsfvtS
hWGrTibqGt++nscoVsXA8usLPGPw6ayCdAzVSD9IVBDhxg7eilbu592Ea0ShzLf0
rqUWT98Opq/11fyOvOKu75mBz8URxM3p+w529zcg7xdfJXLeEEcCH+FrwSi9YyO0
sJ2z7p1EUTILEfLxsbNM9SAaIVAUns1F+xrZUFfGZaMNEtuTS9mqU4kmVSzYiK9w
WhLDZ/1S0Ol3sXrr2j0TkgzI3s7SRwVhrdX/0eI0pGFufutYUesZCMfly9WC8IGY
8J8Gzml8R5n9D5vmdZFL2p4ZxP37FAI4mxiMZGgvhclY30T6lpYrkMTgFVg/Qq68
iILxRRD5LE+F5RnD+ZfbIvIVe2RYqqqg0QfKKOPobBO7Td47qqqVeF9QZz7oF9lw
Rj83MMe1tyn7us+KhyeKS5+GnRc8cXcdmo7V95YUz/eKFq+rVJmfZ3byvuJFinQX
K03Cl2H4iI1eWH07KBch1/PZbJ+IApudjwTySKxTCek7r9Bq13kDuJ1bjsVVGEm7
fuCu1IWvj9yT2iasusc0XjxM0nNfjaU8A8ixF6/2kQZoZS9mExtJg/XYegDCpvza
AATNqAn7qe2HR/uuySzviPgY60iEHyLID2B6qQAOvCQKoGH8gB6fTuZRAXrkkMLt
8yw2EZzTsR/sPXQza9rynGF/LgvIH8zwVwpEFlePRkU8QSzMMgbT1dKXl7BH/8r5
swEDezpUAtQ2D4qdgrjj2+96UxNf2QO98S090sNAEFKinHod+d5IalMrxOwg9LXA
L0LIXCaZfU3ft0m5k+PiUzDf3b8ouYsc1bJu+YxNBykA0DvMyz+1le+emdK5ED3O
ieiPhuXztXajdtd+0sF5BnTQh2QwZUGH7KKHu0jevHcWyi6ddTbybkbdB4mJq+Aw
MUVm2FCOuzkB1Y/DlWx8fsTKPzQvaLOXaEquwt0vrg8esJeR/UlZ1dpWnkKfOSCF
bvvMaZgQE1qeWA53+PneffwO+k1ReAVN8WM8pK2w4m3GcABABYQK2pgxx8SndHRC
T7/1fum36gYi6f7IzOaC7nCxBHtwFhlC5noqItxoHKvQbh1KFFcAaeD6pem6tpmL
V/pY6thNsgr5oCTa4nv2NzaqJQGSGOWkCFDiustLZoMa0XCasobhiGF+kKQv01AE
Iic1a47RcO7cP7JqPeMZGsU1xVnGycRdwqTsh+bSAdScSpvkD5vBmWkoozvyXNyf
ELtWQLHOzKuXl2lXN3y2qYbyxXTqgf+6P5QaCyjgwMsn/uTOzMcc+lCpzPmLl+wh
9NdgeuVlme+x6UQlN354YTbUUhyOkak5aDRp/S+52U2XTKX7OdDQjY3ZaNKVlk0h
lKlfMJOvPVfkeJXMw9hMKjIP9zrHUl15IA7qmH0UN/WKN0r/w8iwnMLkVvpn5EwI
87PfKgofykcO6j6cmg0Ya56CWAUgIcSZ4Fslo2iHeTZqophsUkNEYErFYy30HNEj
SpxIF+bhKOJB/zkUzEmtF2WbjgTc/Ca3OmbM2joIYMdQkWA6ad9M/N6f7XW02qc5
tWbadqV8TJk64xRfcndpwIqruT4IGUsLJmJFZOgx6KDIKVTZkavYz+hh54R4VZ2f
L/st8D9xPdju/3cKyW3UWsqPZnM/pjwBTPh5EwI0m5zH/yuLHngJgz/Zr17ie+IN
bG5uRGd79ZE3EGCiV0K7ZJT+tMV6V0w/n2OP0ePBO3wXGj8kgo6oVgwFGQYxAYqV
qfviYt+wVgo1/U7WKWeN7qZ7eXReQo9P3c67BwWaJD94sirZ4LCWSWgxbxuxX+Yx
2kl8BmOVfY+tcRq94WQrmx/QECtvxv+s8z7xMwdWYbZDwvFwzr5lBYJNv8NAcKCH
4b7MYkexitp5nM73I+TMuCXT4+F1BgZWTJac86wHLzdZRLFa1KX9UeJkY032M+Ra
xMX5+T0Uo4t0UTvJzrbuBFn3iYwg/SqjQEmUJIbqtS6dP5WgEN7AI78vtaSQcjc6
/0sJZsFa6cA9aYmcusCk5px+cCxAwpi7q6OUi/kLwueCLlJHmZeXNqQAEZZ6mHq8
XHv2qPnxZfD4d9H4z4TR3hYWz6dMmF12lHIhwclsEszI0kLxssCK1De5OYgnSI7d
SvRCLa0Gin0a7l7VDYPoIItP4jlGSA8EK9nLn5I8QQyF9GQyAaxQF6brqJAkuUoW
tfe9VHOZK3EvMQTCqycwhYkm4WF2X+v4atZKBfHJU6CVgN4OtdXdpjVclLSdsRc3
SfePNQWDJ/SPYpc8GbudF+ZsJwZbUpIvbQ0gfjmvAo8flAqnJzbOm0ogkSZ+3L47
yQOvOC99eVi/4JcUk09NIadxrlMlMmo4MXTozXQ1m8XcCgvpsrXEkqDEbH06fxIo
F9CDYz2d8imv7EkqhEDPq667aTyw5H7m+x19gxKhEVYyxxH9Zw7Hn1PAYhHn8/6E
OazwjLAk/B5xCBTh7jiZWBhIMxpgg3mKZMbgIMBbzd5D1u7o4EtEP1/5lA390omF
WOrv2UoJSE8jwEqzza2Wa6LvZs9+J3IfR1HnVLD8lFdYY459mXAJOTnWO7EWQ5R3
vC6r+4CGWAHSUQSPY0rCtOc29jNP1h44OFU3Vjj8iISUCOEqih6yLYmrMFSUKSFO
1OrPDQABmgmcYkPNHiambCNMcUmhkY4V5jQnk2Tb+4WLBKogncRCmELJY48YH4wE
obbaLFfmcQ/V5ESoIo5zSPO2hmpT5yA9Lzurf+zZFkD9LUwpHfLjkyNSkXFVhyQz
Mw+opjp8AKHi3TRmuSRbLf1kG49Owda42djrXeQ4TU74SSOYtocBc8UcUUCJA116
+c6rnllAaxYSbqStreAcBjI7dz2jIuOojMCoL09i0+RCVaQVBp4Dje2IUl9mJmKv
DJmVXP7mrPnuON7MghkzX4RR+FTVXHpqiJZ0CI7aYwPfmOKiE5doyJyhJPNNCHt9
8nrka6wCaaPHhy3TMpQbmWXZKMDdKaQKw9Y2t22EI36Lv0ew2na+N1P8cg9E28+R
fMhcv7tF/Flr0GM5Z6t1gHAnL7tUEoBx5ztdA76qKf63aIet0te+Fgbj7OZmC8OC
Jpw2Y9sWlf5kgO5baw+tVyMr32WU9YEyW7Un+hxJx3JZbZUSCXp+NQsNI0GnSeHq
463hBaibag0bn0EFkqlHHihKN+I2zpO2v5+I3ERXuffqUSOz71LdUt6gUbnncxci
DX3j5Ky0b5YTsAZ1vAl/onkiMDOnc+0br3bzp6XMtisQrZdBaQ+h+TU6xgAUp6au
RlPjr1dzRXic0QEhNCROfqX6ifzPE3Z6U9yaN2x4ZiL9QMHv/KxUJh2boVHKxATB
CnoBWYG/7tUb9kKSX8+bXc8HwOad+PQZTl7UZI2+BgqL/b4coHst6YxVN+LrP0je
3tWSCHJzePT95IVhnHOX6UJfRnmruvHfeCydI1rwsXwylqpXXZMrdL1uuMJUZw3y
z1ESEatojZAVDhmf2X3jxONO6lPaJSsmY7TsoWdqgutjqm/7cy59kJ/hTMvTk/bW
JiOzdqLy2hF2tBgZMPtbbc3t8OVk6kEhScIwnradWQG3v62+8/s1t9m0NlpUFh7n
LDP1Mwf49XbK160lrunZ0LVwxUkfDHurFXnVby9KAABeXYgcpqsvOc4xQ5sovoRQ
0PtxPXwBZ0PSH9cPCB2Ae1/U6EWCrsNok6vu3v1vPZDGObftMsoyqbE59XN5/dsE
g6pmVoZcNcDNBkmcQ5yaxmYV8pt3tL/pyRnpbepKv5mhkQHDKYq4rehzQvRo+ZNa
7/RfKDtkruhLN0OT2LSe74+RFw/3ayvn0vgW3gPIfy323kx7JkVkLtF50boxMOr9
QBnyVWyaPSdKS+bqIGZSmpuQCNvZ3+wUzvCvkGQX+3lyI53yWi73Q/gvX8OCr/YL
uqnEWqTneYCVOHND9KcJyALtJI2sp1AQzgnd6lHPBSA2kgeSegEDvs15zVYPEweV
Y6QIkEUiuGS/YTaRXWOjwO+jH+EdOCoV+CzlV0hp8vTDvukQUW2x5PWDeSCttkhR
AUjZYIajUriX0yEeTX81jGm5s2A9x+uZsXGgfyU2GyAHm4R4MocZoz/JjcQwwLme
6KWwzsEMkFyL8p67YE2mZc7D07OQyAE9mNrh7aNrgFlsBpyqo+5WTIbfwulRMscr
ooWKlFJOOcyxNO1VtAiQZyvu8Yq+4UUbDDYm6L4h/pCohpkDz2l7PHs37NdJ7wCj
lCkMbDbbD9H3bFcoFaYC8w9+wZW+bkpTLexcTwFC1QGnFSt+5ofINRLDWqiJ7ks6
kMAWZF5wN8fUyRksnJEqzxMfUrNCQH5lmCkFH4XZ3a70e151HcokgF1IwCn4W1XN
9zz5Fiz+HjuKWL+z5D+Af/ULv++aU0pn8jPjcSwnHBGbZHT6OamEA3kaEzAisTLc
ESrNe7zGsWA2/nODeT1sLkOSADk4VMBZ5S/BU60ASJacNAVtlofs8HcQ2kAhk48z
DakgLbGbaCOY663yQL/OYcex8KHqBoC0HmYDl5ERQN24SnvnU8zMdNYNJ0bEQZw6
l19s7G7+F9JEyy7eB5spK7U/wlUZmzg/HUKjaNTEzGrr2D84yoZ6zdOUhj2etpMl
2SQvgl4m5tXp7p+sCKFuNnLoonXnUsK3F5MmdKuF68GwRQK6fo8f0z4gnjkk6ybO
WKBad71qOQthOS5blIkKYPkHPPs288maVoJh1LYb8HZNiRb3HR1pQyYG5qqHpUMw
GU9mc6Fcd7dyTkQWPrUX3XlE2F1RSAhWjJm85YnSicMIfwctLBzmFHBpVBlf9I6j
FdoOCgS44hSAMeVhRLLtwqDCaLp76e7ZIMAjNoYkceDmgQTvTD4pWWk2ntYoeFwu
c5S+ngf9+j4LAtKcq5Qtfw+sGcL9sOW2H81qRCmdhDmwEB8hcO5n7ma0kmLoHvZ5
MqttXMUzRkfUJpi3Eex1RvtKfS1DzItItsbtmwJ719XY9fs34fyiuHJhSjGPEuDC
m6PhEZY6v8EzDE6JnKETWa3loCYixQIv9yPNcBFJEbOpj74j2h9gKI6R/kYDgcRD
aGCH31lLn4gck5txkUz+uh6wBnim9MiGmyQstzvtCU0GX7xh+Lsbw+7VXS4hKk3/
W3Kn6nXFHQ+QfM9erQZohU4znnypZpt/cu8P44P1AIBjQ46qFq21FQOeJ7koYNQR
l52nh+rpltdNgxmpTR9FBs5dbBReZaPrEu07L77xbdkYnkUnMiVp6NJSp4fQjmV9
gOSMFdN2flVfZE7hTk4nnYU2YtEROO8xO6BSGfxjIwNScOsnLMG4Ugy4Zyt5d25b
cgFcmPKbpBlbjKrSNRrSDPqE3BRTXLbfx2fHzBL8seR8XxFY3F5ID82E1nj5BVI2
Ro+nffZdRg3mzOV+NrgPQw10fL0caU/SrrCw06IAh+MVV7tsMW/uOen4gdtQDjD9
1akVCtztUV52kdcMLpwzToxR25m712R19++HSKWaCsX+MvUi1NIflhKznxr1gS5K
blTTorcYnIbmjAWe5p9IePecABimkm7aeY2JGE3/PLakWXDBUh4JfKytg2AJQki4
4sANeB7QDNbM1/BJ52cMLKPsW5kTVMPMVYqIMeRh78cguqPoR5zyxa2Zirf5APbQ
rxKeoqtPFQZt2tUeOrE+RMij2lABRvOr2STy3074dDlx0aU97lJdQ5Tk4G/dLzVG
c0XpIxPEyNTKJoSc4gujTsy0/Jk3KSM1uT6AmMkdOEmdA6avB76CcR0tqZ9iRoTz
IylX5Mntw7Y1FU/XPigK7M+SdVlwyCeQOZYA8iUcBmFFulJrZsWQoX0BWBekwgOH
L9WaaBGEZn4eze4BnML4EZIIUt+3Z5WfWeKLfF4URzIEsCL51ptKIvyEfFGm74nK
AbzEeaHQfKg5t9/m0u46B48pQ2vBhqLsc1E6TtqIKue4+FDID2Soz2EH2QaY7dD0
5doaMykUvwzK4ZSCp9BCnZBWURLVvMKkvu5a1pzWFg9GqyYsLdkM3gwuM1M83AMN
Pln1c06DlpJCc+5JQ8D4ZOtUreB0zgVTdMmHpXR3mxUpC304GSnTnqo/iA5FIr+L
DW8d1qiCk9AnuhFTi1nCE9mpWxL81iRswseWkX1uJDkgAlrSZqAgyoulpBBynlns
r6nTqEbh9FvVyOXn0Sl3rzW/fr5oanQxinh7Z8X3BGGk9p0PazvNxaoalJcyH0Vc
GBiB5aqjjmpVPJQ6qvKZO8tonB4mQcRSn/Z95N1sVBHgDhNThzShDCP9X6SvMRe0
By32JdfK+/jRM7ObQl9zo55eQtf5SXABBTj6BYOg5u2zI7lBOTgYACEIWk4eCmzP
/RceDVP6mJIOwyHmMOugC51El7EEfeQLUdzOEDmS8lECMpPO27QUnqL3opDtAst8
x8+NN/ESW/HmH7i/W6m1emzvsFnS1Bj6JVBt/CpWbM6TBrWLuNUam7NvtXJHn0+y
7ZvGfGY2icnaNBvqU7uN1tokIxa3ZTLB/I/lwYnvB5oJ5VEkjzeRYBoE+2XUVfXQ
XK18BPuK41ssUQzqlYobPC3LfKhV/DygQSvdctAR1cgUkW4hHL5J9T6jtQrBcAip
b/R+QeNYy8P12riLm2BquGW0C/MmfR6DlPPLGvZDfeSNu5I2S05RmbsKCBU7QTaH
ctWfmjWw7jjTcSF5WrcMvDe8yeTPLoAn6wTpBjYc7ZyZmh9exLwGd0gCh1BNvQgR
WSNZKyFD2zi+qQ8E7Cn6qajbnbgWcCjGyHI8vtT41RZUZ/uCIlY1rYdTmP7jQHQy
ftXkAqg+IxQmi9GihqUpPwmOtGxUnMvgL+pb6BOv4MTGXKxD2gRsL+mieBjczraE
B6HIBIkOTd9Tu/IADcnabBKf6YQChWgUocCj2plAHegw+OOG0fSeT/YxEZ64GStf
y/9n9/gPYabSY+NPyRQrIci76f00rMr+Vx/NKc+jvyoF0TtNDDg5g3vOTJWemWMO
6LyTxB09AsFg77tA82mAv+3ImsLS/0Qxp3F9ubZa+aHtgS/ZYroWWmrl6HpcmTjX
a1CeudDXOk+QPCMoW5nS9XjkMZsUv5vnhNjT2aeKOD6Cpyta5XiBAmnA6L6dzBbL
+t5ydm5tT2/ApquT34bBXP+v0t9brsMUvoH469AKXB9WM90TP5KqwkdYTBziyACE
2WuPK8+nouyLqD5WSWSIGUcQmrBq3FAT83jZ5BCX8uhezQYPKkHAKF4ZJ6AXDUs2
gBzcdfOE5TsrensZ80xl4IbDf1mZ3j/fI4tLZSMb/xOntB+MzAdvZQt7G5Mo73tD
0cjYVdoePmN/x4saoEtepRvtnqzqpd+cuPuR4LMpsgpAQVL6r7NGIa2wI/EnZYnU
eTe0twC6VwhDk1YfXe1+n4RNfO6/P1M7uw6mpuO6J6aH8bqUAQQPMw1/Imwynimt
KocWuxJaYq/bMkuzYGG6PlcSHVGpWTZaaNOlOupM7ETXxsRuvJ909o4nOzsRE2F2
hORmCOm650obVgcxtYVJlu6rWxdzFhdJZMnTp82brHmEIqlpnRLgjVQko1MB98Do
WhhOd40scaXtrmsIrzUfHp9mYYX8IJpQ9RagRy7FmTyjPhvVYdKlcwVjWXwMb/yN
8pwR+snaaeLDDYFOuiWD8+MPRGddMvO7yKJsSRlhTVcpB+TIzc7X4zB/RphW3KSy
BCCJ4G4TMz2Ogn6eUVcrmbM0d/UNPsu1szw8ze5pOdQxuGOfJlcxkbM4z5R6DyO7
OGTnf1dxxuMMJ17tQev//XjrxJ6AbwrCsLdSCwJO/R1BF0IB/WdZy11C3iAzH70M
V/JVpoYVOvFsKm3kODAmcG/jt1wDk5QEbfG0ks8lBoa4VMwhkuTGMKoFLu4eOQ1P
L8WD1vh/kU+UMM/K71GYiiYAIoPlFtA13AzVsdg9UkWeLswjDP9+saUinG+zY1e2
FxZvpbJMQ1e+PeflYI5xNB+GZQCd6W2Yk74ac+oBZMVHXPyi/k805KxwxcuJ4TJS
cF16ceZlxqO+Rj1PTn/nQXxwQBCZDEDRLaGxrpp2JoidD7ZRh2b2i4kAGmABi1L1
8Z1YwKInT7uqMABW29bfPwgl6N6Str2mt1WewNZFS8zLz/uVvyd2cR/tFYTMrnMq
IJvdN9bNiLBwQgxwgKtxkp7SM1S2MI+wGOymJlzPEa7sOodLhXaVPHKzdBCnpKWE
5Z9uQXvkfXwiMVGGsCcioo5/1ix6j89+upXxE0Ym/w2ZUfbu1IUTRmAQVa25m4xa
PYC/HKg4HHBKQrWofvKPUoW+SjBHkA2POW85vJtkcimsCuStp1q6ES7de7aRqD5Q
96/sM1f0LfC67ucIM7a6tcQekxw0a0ppECsVXz0/L/+n7aDazfY01EKLO3BsHyQg
cEVi6COG0WFZlS00695CCTRusf0Mxw71syw9xvOOp5uA74+04+c2UtgQvOI5BALg
OPR6FZozHWbQVJV+R7I7DijOXd79nfMSpFSK2CtCLExQlaygHbUXClZvaBkmfmFt
LcBNYYlW88/BxTwkbBskmS1fIzyqTZiypjoolmErjKAkt0sAzpT2yyCfBd88uqfc
HVZMcki6Ma47bdMtuLhVDJYGm2X7o2VJ2d4pWAcln0+yBdo7aUwvNJ8Jv4CQmXtT
csEoRiBAsRpjM5l3EKzUKIP5l75UPZT/8E0URGEZQGeBxBFGpx57eEUyLjdCLzFV
Vv2d3xrSP4KHxbHKP34S4szEF1eQp8gKxR3pklHTGeNZp7VvTFTQR8Jo1gR9ppSk
Dg3w63u56DefLWkOMJmxty/WIDY5Jm/pDCXnQhdoFYAmGxoBbS6nRakz3NO1E8Si
XCLU26GEYFX7gsjYE6SKS4eQpjyrsiU3jiACMpLqm4NzAgRzJBR26Dlfl7EieLwg
OVewbqYc0cJBdNSd4kcmkNFPsU/vMsZOzoj0SCfaOXQhuBno5/xPjDR1qo1KfDrd
ZlP564ZsYU8fljfcqt9hgmDxI0kvGQcc2vWdkC4pzkA9zMGqQpMB6KoKtVd/t48y
QnXUTWBvTOwqJJQFcUGA4eHme92KpVcDMak5G0UK2AURABqg/5tn/rYCnEgbLL3S
dwxc6VPBKcjdbh3LRcJ8xK8v11s3ghamwpEeUqSWWhti4rpb0swB7fsoTYF4Zf0F
ORMvBym9qYT2Cs+/sLrvpQcFroBZKcv5kK9VaDm4A5pvBK7qd1kNB21z9aez0L++
pgGEyXVhZRsUJD0BFh8KUObZDCNLN1qNHS1BRN4eUHRUC3B3tgxDYEAQ4EVpo5yH
HdsxLFxHEUGcbDWotOBtwlAIp/hWkIWWZHa9KXUVCOkpbHLhR+JoxlqEDzonkxIW
rkEo11JdK6naPYBjemsbIDAkKKlqJXHei1yJ/vIPe+XY2VY2F1krmD/1HulZLOF9
5TwCfLVhxDKwWEXC/kUVaB5aE1IAZR5lapwAJsiEX76bEV4ZVxduI+D4FghM0nT6
yroDQhHCnC3H+nDxcTxO3aTN/5wLMubecExTUVz3paU3a7qNE9PRwbvG/vWDqBfX
Ai2luhl6X/KbldWVkiGAyrZqSj0SBCaePMvx2j7bLx09AIDsg01uT6mGZT9V+oTi
zJ9VRlUQRXBcc20LR4vVUAg7hmtL8FzyN0BOBvfLXmEMwYccKTndAZvakVup1Q1e
ZhmDYkmbwUsllkh2LVWXe7Z1NtYVxdhEiFUvL/4PdyT4+NfbVzLUp7wQ/3P5t8tY
BzgC0kwPPXmjI6x6EFdHwy67rp3ohvQnyAw/dfaOKR8yNKNBwKrP7cr0ENtSv0j9
piclDHU0qMZ0nWBju1zeE2gd4iVSiH124N9zkkRSLO5Pz+FjicuPLDT8VzSp9UKt
VIKN3+iRFLCQZInJ08bJ601YnKjL6RV27b6Xv8jLEHk/5lagqUptWYmErmTGthO4
BvPvx0mWkD445Vva2GGVpxAuFLaRo/ORSfxIp0xijVf7Sl8S6BZ5/Fomaic6W1ch
8+5oDBiLOXqJ/Q+dF9h266xyFt7WQja6hrey59cJdkZ55/qsltiep3vgrkm5F+KI
qbX00tftmjcJb6HsXn2yL/HlW/nPHDU4OA1jvs99o5aUnJGRIEXRIBgF/zDRmwq+
cCsfJ3TONlVf8TGqPJWQJ+5YTEL5uHWWQpGdc7bVfW1FeZvQ0egqeQbDuOx+2rZk
PVb6c5WG4VQQxdPBqJMxyye4QRPcdn5chTZ0xpNIqVaH2GQ+QkDZ2WSfrjZlsx6R
DU4xa5YHvU7kadMSYExOIY6oHXbkzehry7fCLrPApKBwTsEBb4mGvYglg0VizmXw
BTqKbFqIilNefeQf6ud5482dzvas+CXlqNxi6ELnRh62swEAHsxzo9o2eMG2XStt
hYM2bDXu8HaIuUscL4+4W2Vz/qVk60rHseBj5a+MwHCbIZUCZjTybBkPlIzLbCNf
6CRlk1KOlei2zwkzZa6wcjpCjmWPiX2RgsK2qkiqM/h1AhfVN0CtaM3tzM0Gs/5c
OV1gAhsCtD92BynHx2symV8sXTTjXZO6j5AfmvAXLIrNk0TFe+kp0EqIOWE4VXCU
cfnvqjhKlJJDsmJyNNzzbSRyzYuZ33uSO61ZG3y0G+jXNxNrKP63+KXL7T1C8pHE
2y+GoYMXCVBGWpAtirgGnh6jkJ4iLXqpxwoZOxQbyuGyGQvHLOKXohAcEUxqpCdM
+cLXo88+2XeOsv2NwGwq/UWTl/lQyRd+RaoGlYiKCEXmDFmT1m33ISOZ5z8J2J9b
taDtcwzFvKMsfVGC37n45EnLg0WJFPkr0+6fbFvLd/dFc5HfvVs0lUquGLKXMDKT
7CuKlyy2vWQt//XhFMDRbbU5wUDrB/Z3x2NV9KW3X1/ZaUF5O9e+FZ2ijqmygN3T
6crr8gVMoyPeR8jM4R+2WxE0+8v+eFt2GjBsIU3gwsqHvuENlvD4OCn3BI5HjZAP
inbKMP5FburmdbAj2phYGgN98BatpqSFRdePR/wFF1s4vxifJDjkIUd+XxG8zOCb
sReE/pcAVFWAeZMafi6JllRGpXbnnH+953uC6y/GwIeVKuB8PvSe4tsC2qHmfMx0
doj8hDDNELokQnjxWgON1sQOSQ8NulIdBgy7Yrq7RFAqDtJABUgdTE4kvTikX6hf
6jP++VQO4VqqS1fokpRGee4YS5Vc5Tm5nDK4LJebPX89lN+/fMvh/MBbo46hzs4T
gJCq1Rbig0QP4/3ZERLs/WKklfi3tJsVVtgfPUi20Z8t3o5MKNmN6bbEhwajPnm0
l44/X5aaebwXY+YdhCNT7Om/t/eglnAL82AsH6F+YrPAvMDNbVrpzxnpwpIs4tFP
7NVK0ioWw8c4Jct3qL+2U8n3OguerXoIptUJekFPRT8jeTOKPL7udIJQc3t1nk/h
qiwNHRGjVW70WlLn+IVpUgLGKz2Q+oPNNYHxzkUQftw7OjCQ1mcYmCLo8dyhoVts
scQbEZpecjRFPX3tWAOEa5mGG6MvNrEN5QDLEyWJ6kqH9RGtQGacnEviZpMYRZaq
TTYjvkrA0W39ytkaSmY5iUOc0CV+yUvUb4MZC1D6hMOB35oKHNTHig2MzDNlgJ3B
CfxSw5O9YlIiVfxO57hHVoFIzxfeHGrZEugDoTThyWIbYHSMdhoEWE9w6jcQTly4
DFix+pAgcQMoAUO3Mhs95kWTPfZX3HQYiCJFD/qFacRX0h7PTg8jRX8D6aqUlHhu
K940QztB01ScY8t6eBAyzaUh45A9DEov88UfCckPx/f7hFWIwYvRa8xTpuzVOmOK
rkp6ho5lrk7Ez/6Sl8gTwbieGhHSqcN3xvKlBosk8OwtiVeyjL3YAb/XbIR1lJ3P
9zsS8I5PfD68r0nyBESa5rkQf6dGp6A89fH0kTrL1fT0zGhrE1PMvVCAUY193hoB
l3f0XTQ2kM7H/fv23yi3WAqK7d9mZQoHRxiQfh1YTknwzy4M+UOJZPvO4fGrHZrp
1yofxgByRCeXzK1oarOr+39zZ4KK0vV06bYv23CPqXitwusS9ezoauH4asqP6yzX
Cw/tpshK4ElOtAaPmXPk/fBdD0dewre52jp12TiVaAhx6uulTMKm1r7bO0KIWHjD
uhjzwh6zh+bqCF7ri+3xV61iph3v4fwCBD6aARRaQFcfU35vLyLO1W/QA4ZTaoQm
4dB+A3Rk0uZ66xWxoy4aVRhZgiyL+iMbZJUJstyZSPytlz5yjwSlvdsaH9oesmpY
NR0N6dgDgUuoUt2ZnhpIuAlW1X0nmMd5XcEO1g0ZxHAs8Q9AeDvzPKnz20rsIj7w
UrR5oh7pQprpDNhQMlbfRAk3unzJZGRBEdkLP3y4JTNi81f6En4/1Qw8TTlFinvM
Dh1RpblgI3v/XPSZ0ifWGzTGIJcGzGgOaWktd6a0KDZ9FLv4Dh3zdfYpqKMfjoYu
HW6rlm7wbvdwZZ3K5TM/rLq+4hg/FtYp5gQBbZh3R/WvAQerU5iGFIrD94vwxKFf
AtXh1xRRiuZJrJmrB32QuO5f6wmxuL9p8oXpgKx2RYUXS+Xi3lnGw+tm+puPrDUB
46HfDbfZdZmychoC5MElIQ8+AR/BVI7lI7Ao9lVIlclanZPJ7LSDTPNHbIZWgiR6
vgjbGrWDne5TJRrsK6bPuARXU//+25PGkDI/qnCPV7JxVWBFiCtNhDOhfjEs8ntN
+b/rF6TVp4kcYDbZebY7nLz4XE4TwzngrRucSFxdPcHh6+Rw9IucJtRyB1hR8rVS
OiergrRkgEA2W2ImAoTF6DEAWXv2MXZVakp2h2aTfCMO9BJZrPiBzLPCAzDjICs0
N1oLxDHDz1MEnIUn9YPai1pcqlZUdAAFa78sOJ6JUY6dczF7Mp9jux2FUivq/k5O
y77I5JayTha0k1w4Nysa0uwA2w8eBGoOv+BJ1JDOZyHulwVBbZo+Bq+jNmyBE2f5
o7xBtNRwnc4KGVmbWma3fsREOZIb3NOo5Nalh82neDLkki6JAurZkGQWxVHv1NHM
3lTOBS7HX723FqmRWrOzmEhEcLWqftcwqp2x1f+1nqqFwNGzSVI+O0WSHPrdhO01
5lA5jHFJSUgjebBXcZUNi/JVzt4++56GOqOrFPbOPJ1zVv8g7BwlwiQtLdyhlL3n
DlL4bmpMEwwScHqsxOk/0XG/VqVeQSydqxiUArA5tLBcXkixICrUrfpO/hgJafNb
tz/cdKIehMD4i4PpSK3xYPIBvg01Ur3oA4XGMaJaGp+8dC48ZAsfZrsFS+iwsqJ8
7i43/gEeXEaARxfWovopXtFRnJHeoSBY/aavot7jBEpCPb6zync7bMGvDTRkH02i
XK3PJkuMfM0Swb15vc6AuuzrRrVj2TfOIJg2XJcasOSoxLEFUkOzAg+0plzTTgpx
I7ZtuhhMzn55gIPRYu99jW7zj75WXWJNxnLdelK+rSKdY2Ai5rJzegohEdz2LuS3
q4QIOtF3qPg1uygqItUSBFygUtwXB3ssiWgw1ne0FHsKzmeq5JQR/4mu/frMnUm9
qBQrxuKQ8V1KIWfeaBgIv/2ogKkaeM0BgPUF5HzTqMcJMxPRB83mH4LqAvljRjQE
cb/Qmr3KpUxL3sNZU23b3BMZK4fH9kLeGiflYYqr3n4IlH9jFVh6CoLnAB7pZCek
Jbog0YKpky2YEP/Ev5VlE7I95BhcHLp2V/yZEWOruaBt+fL3ejdKgiWF8qQb4mAg
VIK6fETgvftT2eOd6XQ0imF1RqfSSDT/XL1zSFsuDWK3TkXXT0t9LIPjYAktZr3r
MRUo2fS37Op6YFrovYn7mhGHoHBDMBkxEYxkWId+wt6yBz7OC4bkyFbGn38mu2PX
a9dyEhhXvD0lxKwGP6D7O88omofq3YlhqvZhXJZqOTu1XY9L7CzOCNGUo4UXSaeX
v8L4h5/NJKVDtXEv0tgc1EE8leZl9tIXX6qqZc5zTOGhnsFNJwANcPSj1hEksFy5
68mAVh+BqINZZTrOOUoT5Ep0hdDj7SR3iMv4oO+TGnuhyw2M6aReYueoyDhskE7i
mD7QnjtwqKJ96ITyWBiNFymjuiqX+WHJLjbM1EGpeEFDqww9QoiU+ujoGdYX8Ki1
TExklxi7zeXW14SIrGzS/pGDLCXh3sOrNdmgg3Zj99LEBgQLRwEB7/oJ5bsdtI5W
pGjmJIZY/HKyLERlgUOBqgsppuTA7c5Vsg3Jwt4qVr+vYG6md89CqS9/8XaOhQ20
VfYWnn75lHJ8qloROG7Po12JL8wdlUpAoz4sIZApWVCaGiQexsmzO5y+eqOGNxBD
DfekInys6Clg6gImk/UsWXCZdNFNba7jPCJksgdlQMk+fWemedmH3M0ijgyqO2oB
rPK7K+a5XZuDXwqdRG7FaPY6GfOJCZm1uxAnSVcQEWQT2GVjn9mu7qBRa/epsoMr
ITZuocbMn1PyfphAF3RTNhcx5i4UI5y4ht4/CG79grDEwYdM7dXeNJ3QNmhb8z7y
h0DkB0Vs5fApFSqgBgQ/s3u80wJaRCUp6kCSUg8HbvMY1V6WbA3UtpdBpcV1VKfo
P0nlRBSkSSYSQe7qdMhvcm6oRMO+v00rZLfrZSGAava+1FONEnZFiu4S3U5qGvR7
XL+Pps2W9EobLTgcaEbto60pa4Jz7/zumy+DIeeISMSP8GJpvbH2Uh1RGlNUcQZ1
bfPcZLkg8LV3n28N0czRuw/0Iu06+gQxli+NGe9hPJfngfIpvK5YBTnHbfPcRcNc
oZRMBfjkxjlKhPzfWKyMmhmmKOpRaeYomNN8m+GWLi9kObN8zLrcFjKsPZZXWSc+
gO3jb8y1UrBpJ69VCEBA9081Tt0WMQuN7tbS6sawXk7//Tvz2IUm/GEkfstpH+c1
sNxGyucGRoj4Yy2N5T5epF+72RGiUog4AaYq2SqD5F0WIgTso2qdFI9tFVDb7592
PD9Ev+PoQA8ZB7bOs80aFPHeumVxDSmw3Z+J3cQ2c4XvnSndssGSqc/o+y+DCYBK
d7QpHjeTjkaiNWSRtozW9Oqpq0/looUAWuZe9OGL8x8uOE+NTKXIN7L6DG7SgUhm
ujRe2lALAN+VXuE49UiG3DlnVAro/KCL77k5t7tUu4TdwCY0I7VjQnjbor/tqaGE
n7CQOxTnu6UgdZWW444xrYO6QtmsBblXNyhGi29Z1Dn/cvF9C9JWbDcfyMpThK0z
GHjFChfpPnqP50bZd130ZszeNZeqftTioOZhYcAXGDRWSrS35DpyTC75n+P2avWr
Kvd4leXkFCmTTao0AY6AzEXAcHMK3q8MRuj2+fw1JM3xz+wgGSrt9MDgiOsF+sE3
H2/ir0pE2jeaXjb0PguEZnwAGC3PETYxxcoY23ImJvEstWkgjmZDibviCqB9xLvl
gFRToODYTnL+wyZU3MJACm+4OdJgt3bf60YRJ7OXzYlEhn42YwN3VzSrq5QnWwMv
ZIPPjglllyFdKH9M9NZSMC2uOJH9mAJRwYU6m9pgyDPrTTMhwt66cXBfe8SiGsqg
VM0PUxDC+HSQSuK21Gu5Z/pMUcn07qJK5yf9SXPnNoOAj6hEWRN/wmHjChapUODK
xOTYgekD3RJnBI999zbg1Lk1RoHoGZApwSSq4DzueY0j9FHzZxGlFAGDvhbA/88N
8EcZRNHM88zeUXJq/J9puuszA0n/ON1UCHF2BKNkAVQQGSW1YyTRX+5+GC4u6C8q
dxkMDY17rban/umNiWvi4n+DEjXGgphkaLsfcamA1riBHkKu4iH7qZvbqgYEzsgT
ZakJBGDQmITiChYl36YB2wyTYJ9DYe/zb0oh0Gaww98wS9tVfPSI649Suv57JXwd
PEq9Dcge2VyIMHf4hSnY9TdUexnyD/lZNbZiuQ2gW9ioBnN43pvj6J7v+Wv3Ic4r
7mxcB1jcfSK49Mw2xSR2qfN1ZxkNMznV4CuaEPli9k59fJan/ob8Ky1LV/oAk1LL
udtulm4gd+W1cRJQ7USG8/k0sd/WaJOirIQzQTp9JIiapmfNfX8m/yOheNvT0dO8
C0huLjEZ5RO9628G52EYmjerOB1QIclvOYPfem3gWol5h5hOfy0lsXOM7gP6EetX
Eq677VekRKI8BhIXGp7iMt1lw0r04VB8egEr7sbPiW/9GCHMKkVT8qR+WpBJYA/l
wLErv4e2rCscZp4brReN8Iy6XR1JAIliCCKfnZhKndlGG0AD64hr+v81SW0yPwKM
T9dSmaLFEyw13jfrNUWA9ZHhsca+7U9e3cWmaF2EWyxd6b51j8UhgWfQpvcztoy4
DnuoRH+t6Ok7Wu16J1ax07rZaDXy8FQateid6ueKKHlkXY8+A5p12dW2Z3Je6plX
FGq7qTKTw4eqElptRdRWM4cztC0wmtlqHpwddw1/gZpwvAXAeRXKBX6hRAR5Cap7
g7jRc6ILWWWmcRTNSxm8O/KuzK128xoj6Yi9e6bh3asYhqoD/OqF7XZmV06+WEQF
qfQtXXhy72ntX9vEwJ6LV17+k6vT4UDG+0Oj981UethOk+sRtr0CIymOuddUDkuN
V+vu6gbA+hlj7L113UaJOAHWcN/DmNi5djhk9BsHQYIeCDGaSNc8P9ZOIkjhYT0J
6x9geyXiOayfO5wlbwwu/NMik19hZSiGeJVAijsI18el8xUkxDnOuKDfn4o11Ttq
j62nwqhuY3A3Cs37yT8nNd5aoesz3b1RB/oGvlmArBOntANVjyT7yK2PXlltu3HU
4JRbMsEQ9g21Dp3qtezM/abOLDl+9gVZTKYtrcbsKlg+LB73UkWd6ORserijSVgc
g9ffYee+Y5UICMzyqv6XdkLJgK/Gcobi84l3VhTfLgSVbQlUp0SFeo2FnvCum7s6
L4RQolhAvFnZ3ZcnVTqmlXYWUXvnY1BS0R8heWQjohrCAbLzdEjXBMTQv59X8ZGm
X4DKtkTqa/FuYk+GqVozXIXr6y3Wcq1fhqAsSkhvtxLlhySYRaN7sv5XBXEyG6nC
swH7QAolIHJyxB5pb16A2pH7UDSlWNoE+rSPnw0X4KXzWYN+GgnxOqDSi8SpTe9l
EINsUfZbU2v+8KjxF3Dr6ksvNqNXOcj4765d77HQOXWEaVVTa2klsZq20uoJWlhm
XlzewRXmAYw09bcA9Nn+XUqhzrwP5kVrBkSDOT5wYLDTQ7OoJ7zqQWgJLgZ2YEa4
cTSm8hmSIUmWG0xY2KYKY8euvfvd/C/EbODvk6gzx7Gw3Pd+Mrt+y14Ym/XWlD63
DCCMEq0VvcFbhsKRTYXfUHh7M+VS3MjVWGvBD9nlJIdzjLRkztFYlSt6N8965rTR
oZAlj4U6mYnKRDWkz0teqnHeMGx4dXWtkYt2+X8bslTuHa7bKEwWiG0tqEczM9ZL
u2XXgX+DdDKAGV9whg9Rh7Rpun8VvNRbNwxiaXfcx8VXUrtehwyEdRQoD7kgFdea
w4zIiptmBFkjDo0p8PbtBAzdy0ZRmucuBtgwpIFxauBVBJfbWqEEmZI3/uRN9CNq
29oKzJ4MUkjmPPeYazDuInQYHyzz2bc5Y1ONjtpDKVhGfW/Id2thQE3kJRl/la68
azAJDxTethA5sxZw2mXlqEFzamH30DK435B4VZtBEA6jw5dQrcouqK25SaU6k75q
rnG/6x4y9xmVoECFMJ8qon7D7BUXyw1WEVaI1T3sg7m7ky/Z5zdKOfzWUW4/96/G
p4nfTc//AD6YZqLSv/4kSQCoavaDJLF+xbYLs7L3kII5O/uhbFy/F9C7an4jnZ8P
ys5cMkwMzW7c13tYFL7bPJNFeFM47ZIBmrO4kqMZ2DuUqr39HesaB9PrpOgpd+pC
x+t0kmj4Bd5whZ6VkAy/jfx2xv1EHUmeE0HDt8UkSKg2HTSuhvnmnW8pWKky1u+6
Jq9dL4MJl3rhUswKGBrrdNgZ6mYPCSjcripgsSxR3lcbkrCzGOwMmfYKQ/T9wiVs
kFwY0nnp3slPUc05uMIOoxGobSBy3DzdTMGL5lMrFG30HmtXCAT8X/b/8vzMxmtC
/jaZxel7yXEdHx7nuysOEuq7pbYhGCqs/Ij5TTfz1ozbPNwI+b3eLNZhCrAf8HIp
2yn1qRPPyRhzCWr+MePiYGxNTor5dGGX6qMLMoucOIQ2ZOuLmlKrX9JY7fquP/Lk
D/kYW12obVOZ6qZ3aK+zhwqhINva/Gz+Oelcdic0GBkAo2PkCzZciN6Ru942weIU
HJXngM/Z/97Dh014P4ZnkLbnQMcgTY4CdRj5jmqCVdLoOE1GGbf4ZV01OKxRwASt
aMPte717/HtzxsZekvZGaE5u4qxwGA6ETC8IXSb1usWVwkf8mZZyvLk/QiuHkkmr
daUkoy3dSSikmCavcUsmQSNhwwhnByVsyq8hvNBkQK6H6tyvhGFq9P2xHvQO+6We
VlBbVzqN7Gpto51xxh7g33SJLvs1fiZEj5gam2FwrQYYUUrRU2jSJgiUwcmQdsTu
96vo1Wln9pg58qxCEdsUUuVO6dUHsAJsE1ixEi69WTjUSUIGiBaxz6igcaQlH7ZU
fGleG/Y7DEyAJMIrZTXeBjOKshYscrqg9mpmWHjTPNCScsZNAmFAX/ajgv9QLAEj
quGU0iumJpuNGxWcTA3ObEB3dQ8pSsz1E+wfaP3RS77cZ+ymqMsDlGZIAdcJjDEK
JvBTlff0G1BkZp0eZfzYicCapHhs3j58Ktdh15l+b8yoYojyiin3rUzWqZHXeOlr
nQMdTS3WUxJHYmfLwq10kuBzEI92zkmi1OOnMO7fwvmQLaM68Q24I72kkWoECTi5
TF6MHOYha/yNSckTg79/2JNREvzUTthpVCW2T407Td1kBhqfmSTH86RM+3VBR+/8
fwXjOplPvcVxMFw9GBFLwuyz7Ff6zWQR7fbn/Tq8Bxgz6vKz5MG5OKsQkNt1JPJK
h9gPMHxfsrtg0IRIECIP7zSseYhwzKe2umnT0vu7P9kSCaqd3DGq1+dzltxMMyyx
nT4RFU6ZyzCNBTyfma3QqAmWGfso0Mp/O0xPOTMpkz1K+QBG6dgkKtWq6kHDjTj8
5eJkBRfUt79tpTpdirTMDFOzaKa4sasv5zrEc0VqSqKZdOsfe8QbjtDM4UWOtK/D
wsJJQ7f8L3PMx842M1fEey7HERByQCWldCkU3XA1wtgYoFScSzMo3wPIesqnum2T
u3kTgBBWiDVJB1XV6EK3LIISFNjzcfHtr52U41r/Rn54wS5ZuLuPi16m4RaYwrCU
/uRnzrEKzjDl+dYN7MoqqTsOESwqwSARaEvjgmyJH9//2p9kJWG7hB9/yqNdbPkr
6QPJfv05xQZevE0BiN2mrAVEiSFxvcPoGEFRFTu+v6wZwrYsQ0lbo2nb4yRNh1+C
eBcvvGRZyENnK6D0Ez5CV1wbWJ3fX85s14fz821WmpSJIEw1mBJqWgeszLPetvAk
Rw6EbdmO1ugDBMts6cLAzPcbW3ag7ue1xqjQzrnmx44liB36bdVn2IV9BztSiftZ
+QFyG3B49+B73eH9abW82pZAagXNy++D/3r/ojqmNePAUCd1wksMADsSlR1fhopL
0VnlEA9ccqwN/80APYPcq6Rgh8OnB9rwjznRjWSQHUJbSethm9CEBq+2SCkI31hF
JwrdG7K8qslS6adbCTHAcswQrMxAbhUSzn7Fy7ZQWXMpR8MAZOHGFLucgPL8B3Zn
P0HJLhjlKRRQWlnylRq85pMBId2zl1SOvRh5QHMmRMO9dducryIZMkG++3yiidz3
EUlZYtvl295VML6NybvG8tAvO76UQ/Y23qIRccQ23CM/T+us5Nh3VC1gSeTgnz2v
SAk1TkFqjs28LEKLE6nqbE3lp107foaR2D9IT1C0hfbfE4OXoHfM8rde2p+1yCEf
sdzV+IbRYgIFFycW4ANzjCBo1lK8f5iwn6qDZHoCB9OLF0bql1N0UmGjFp5G/xOf
qlJInzB2HoeUoIZE2lhSzTCFSVtMudf0ApggpWVmqkhJkF4Ytgc6LyXrFZiW9LpY
bZm1Xhajxox1Bu2vgvEh7SP74YsiJPxVCKau9lkNx0o9N5oyciF0hihYApHsTDVJ
bBTez2TcOMDUMF00Zo9R2BXRHG5McFAWwc9F3xvt3HRp1bEsDZdpbZQr8kvy7Eps
5X/IWdiYnZeMyGI19DAXgK4q9j5aOQSLQGuW5znDGv4yqdOR5ArZsOYfr3W+qfbV
0kft10DxoBDlPcs4j43WGLYpQHzD3YVRpcCaNrsTFrL6I7zCxSDHPfRkfjP6/ppE
+kERa22QBNVdUu/Iw84HSaYZcY9jnJGyyEFklOh+p+2rkiqJx9OOIaq9/SesirIj
t2rgfb/f6vDRupuv4BQ4hYxkGSYUv3VFAKEVL7qBlSyN/cM7HAYDiIqmCLOAta0z
ANLGpWnayczhFCDgXHwJzwHgq0rR/FCekfO0j08nXBD+bR9Z5VVe9HBF8/c/OM3p
8WGdwt71UoZk7tyrd8oaXAzJ+Kw1lmFbpRcMlT0P7pF7A9AhYqaNMTnRHHAJfnCW
3qZLXaGTdXOdPb+zDcgyYpaSj1eWWCEa9akNxwxpmEwesfAc2X2gXdgOIyjUkbD9
db0BIqTGjh7D+gtuUXHzET/sivAF7ZfMBWqnq9P0OSjHEChcX+6Q+O2Xn2DfH/lh
249QktaobyNIOfbhh+qMgFbb1dcIsSIoHV09/gMP7CfHxY7n6EHdO7TxPaN+qEv8
x8Sx37QVe7v8jLXVnoAvyFq/n7nccFKNQYIXQeanqpWnPAkv3Q4KQNbNgXr8dlFD
So/U55FFroJzfaCkGA/eE4AI56oCfaMSIW3yKxJaD5lPxkhsDlEYJGOw2SZIWVgu
abke9KsRP2AEETSjmwohs7GsEzgKRPW6UEBcoFxO+3kboO1YT7TdqwQJhT/IOiWq
iWo8HiqcG6YBa66l1QDNGiUMTtDBnsVjmn9X8J4Tk9UxJtHaH/IcAj3CH67k6v03
oeCgDIn7TLq4uxlRax8n4btDt4cu8wkpo4ppIlZVs+RmSG3W/xcR++h/NKKQosOP
LPDRh7NUTLWW68S3sw1RjMDnjMSIeVj92e0ZwNEBHn13UOAl2doc9M+RBrkMWXH7
B1KeqyOyHReRI/uPbeS+4HkPua8RWgirNZxUAvJT7D83JwbqKPNNO7LSkaCThWsz
djiKZzK2MfiktwdYeKt0HKoHQK3tnKjcL8XGVB33KjqYR760si+C4gk+jmR6qTHy
voXAzwWfqy//pPYbZ0R6xoZVnJmYzru0mGi3n3HDlDlWROgW0U/IJ1L6RWsS+eHW
YD6aidp6DqU72UPow8MiWJ4pe3ZLbMVK5tDY9oddqG7T4JYbGiJBcLudqVUdPpYv
hmG5htUvImkp4J9GuQzYp7c3WJ06rVjj5x6xOEOXaW5mC5TXlzk+NFiiW3h4Qh3O
8/ZOxlN5kd5Zx1wUCWvcSzwV4LZLf6mOvpl6waqD5m070VzNrlApk+yzJsPpXS2D
/PfwmWptxiHfPKoFe8Rvi/S0J+tgyZT8+hmdBRvamOOANTDNPYwAv6jRcpKI0eJL
0rH/T6k3t/tcyYQaoqpscvsayV1zPAGrsKJg2bWxWl+ubYBqBqpWfHmHO0p1cmxv
/jh6tCLW00DFhDdRd2B6cf327qa8tEtwjr8F3oY3QQWd8Bj+LxcoGBr1dkK4njxM
/wlYSjnV5COrjX2prbGttzEE6FF2UmjtPnZpjySGm0ptvQWKVWvKALjf1qUxto3z
kx4ZGIhedwHTM7E58/eJv4bXuU/nSIxrJ+2joRcEgWUQp9LT/Ag+NI2T5EIMwt0u
pISd16ClGzCgy8oBTkTwNV6gYk7cnHm96sbX/AZtULJzGFHFJtpktuti/E/rCHEt
Oa0VGmscfe+x3olE3XJtKqMMlYdbltZg36imnUJnJ7EkfXPpGGE22oWtQYz6hTJM
m57HEW6kN5aISVsT75I0I1PusbPRrRFD5CtgIphS901SLcjCVnILh4Zn9BFhbIHR
Dnnn/VCrAX7axU/sFawp1n4N6wuCamjukVhnzMwaRg7+ZDiu3kct0j/Wt6QwFEwr
z2OJ26rtf2e3U8cJ6IlCV1nHPhCzh/DtkVaNyL6f45aux5ueWH3PMp++KYy2TnVq
sXvaRQ51ZTmEZM9YrXHEKiYnCBbJcq4oHz/0IWwSvSOsBRReZZ3OrHzoWFDA9iNG
umO1pIIGLtZ7N9YUNGDR2ct8biJkEW+on5/4dtCebzvH426ggauonsv0iu0i41s4
xyOaDnnBTvS1ca7l1dZLlVmRxjx65cbHRPVNcPvqLHmyCU88voXUhOB+WuBFlcq/
29H1R2ra+yQSse1Z5wRsZ5+7ZFngFK9og23EcwFiLWx8ps7j5chlz2iwvR3x1BIR
+196WzJgCsN0CtvlNNxfkHCDSoQxHf70kF/19LDJ3PesV5Mefeh0/q7w88F8L7Mo
mstKoDNKfAQZsqpOmfRTHVyPuUA3Q+3gbkw5f1PghWX8/OSsGRz9hQfJ6e1MTJ7q
KpS99boWeolvdtzNQ8pPyYORbKeSIIodwAygs4OukNMDV8vMfLEMwDmjsqmudGAY
UN8GHuODIOP0RF+Q9GPyHoqtL7+4fVvAeDd7up34Yfi+taPn0x9ddaY3IZ361vLL
Q6uKfb1p9lWm75y3LlBWdoRJXp3rbSGEOBjs2ngSbWcOfYBf9hApyN1ZrlP8yj+1
WO2qh6U2urEDyydrdZHih2H8Q9WaTQ23KvqsUr1wosay8e9Fu3Sf2tJKQjeURT2M
gNdnKJr1p7VImndHIY4TkWmRvjc9MP3cx8CNBTmCyyP4KoJn3JrECIjh5XczUwY7
D1ipNbOy3Ff86udKhaaXGOOsmQogKoXXtoG0F35HtiXVBUtJgkiE0A4/mSxWc3TV
jmhQuNPEYOvuumIhYmzsI34W45msA2n6vX0VM1ktebmh5+AOF0bXBhax4UYGQgiW
O+WroKJJ+n3niNHH/apx6yxRZjpI4neIv9PVIwlUNdHLHxlzCbCG1z05fnR5U8X6
rYP/O9G4ll6ahnCc4eqo0Qb7JxB+jR6KCEgaTq8yYboyeEj/tD51bxCfGupXDH9b
UMsS6Z1A9kjyGIFygqkLzQB6jzQPaUyOGwBIU9L0G8j15uDETkp3En7xh68ytGcz
NNlkLDmpsM9HX/Rv/nuQtD/+nbXlbSpsKe5U7y7uy63HGq6KNWU2PePlqfrPMdOo
aJZCiX52OM+zOgmBIKDxONWfiS2IhDKNR5dkYpKlhbA5lWE5ZaCNqd4nfZiyy7Jz
anAAGvLAPBVyxppGVEt4aJCuXNyQ+B1Qt2jUIeTISop/lYDVZDymg3aoRFens8Rk
kxlF0M8LMQ5JlkLVSsNhp0wqT88RA+PpQ9ZHjg6816sqdRP+64yBmEP94hfPKgp6
ftw3DiGT6aCd4l9R17Xx3zcvdW29caU1HVAV0pMkdQqETIHujEuXFjCe8fZY1GHt
EXNEUJeUVGIVC+PVQBdAmipcSsCNtQfAvzTCyl74UeMC2J5V9HcQsXpe/UI0aXYk
ekGGcxLPYhZTZaL87anuX4HIXDWEz1ylC4nyAGmyJF2CqSNW4LRiLwaRzsu9tg0v
dxLtvdO2Zl9zzUujcTXcod4fuPEepCKome4LP0174WN3bIXRsQx7r84WygJbDKG6
qZ9Q4/zSAnBwgCJ3KYzCl3x3cKygQn0GB1YBBbascDt6bu43RNrVAHpohAwJ1kfM
cocQRw3obfAko5SFf8FuN9Z+/Z6GZj6h5SfB8VLHyOZK6Rybe5ANoriwXKxAtmp6
FBnM9UEXILbY2otcJ5BO/SWZxmXi4w//pHLBWtF88m5Hljo2jtvym0lFp4gnEyKf
LFWfNdfgPSoKXJHFcUZCtLORFoUFbWrse9o+Af01kXnJmfpkhT2nAkmz8ZpiWkv+
oOgUZaxf0R6IFkyn75tLp1X2ATRnRXKZkZwsfEU4fxxXDiLxlEUAdHep0kmWS0+d
GDatn8rWVE2OiteV7tKkK0hHdO2JKpG3dn0W/ey5t7dc/lWj6I+tEgQcoS03FPqC
HY3I6GNNfiKLyMFauuY1p9r3UKcP6niiXt4ZUD10xkhB2j0j8unsGfAxc+1N2lj0
ra4LTZRsKWg+wGtMjKbeaAitbsZq2yJmLMFciQEuzzFo3lXb8SqnWuhbOOJx3zbn
OKQDwXu0baN7kc++Iifs420ro2UBm8vZ6/KIF48zQFxznp49o1z14SWgmpfvKazt
pCIMY7o4pKQrLz/JcrSkitaSRyFE7ji5nOnXBAbdwL0gL2EXENdCxXYlakD5pFCk
cZLf1pRmb3EUnpqg4tSJ0rfFxIGc0cdTOJ9FxDdMEoPrRdASRuiMzbM3WXegXtnm
MG9Nl22KQOZ6Vg8tUpiVAyCe41xp8RO0GCu6MmTH4vzJgwRp35c6hj8YCRIVQYPR
NTVDdIPzQpMKvUiuKjlYpRRpuy9Z5GB24RWR/0cMhdqHpazlVrt6a+Dn96ZW/B5K
qS4mRn7roZgX8TLYZ6ckqHyvMC41+Kv1yMz6eEB9upaPg4Vf/qqIH9NauTSTjvM5
EHAOsIUtg9dJqSUFFwZYTePo9eBeM2DRE5BrIa0k3+XHAfaOmrXBpsfp1qZ6J5u9
nlnuumBDjJqvehTPxz01pU1o9WYHCUiymMiKEiBTKqWZgKMZ888B9j0V4l6iLxCq
QMPGzyIcW/y/UDNznzoGaH7Y+ROFwPeA1jb1FmlKRc0cwc9xwIZMtF/8nH1ym03+
Ul4SZsHuTFqGHPqoY2BNQ9Vs58StQQTY2R9ApwNEXsrkUIrkcf2kGs+GJcvoyZW+
lXwxXZZDiKsstG2Z0ywHO/rQMeaAVZDmfRd5yzCOSjF8tOPP7nxigEOuIv0BJGe1
3eTNsfM6gUZrfNaSsMppOOiC3IeYjSNM/hJ78m0w6W0ig9YWDGb8jZpEDUqwntPR
GX+TGf8iexZTO8D80opm5c2P/JFd5Q8vrpwoP7n0OIRqv6n+iGKONW3xq4+pwifk
Ltrwsk0/pW0v2KHAeWOtoJrHewRxTLkSUb7pmJ6mUGRFJ/Jpsv1LO61OSzovp/sX
82bTAcTaSanNYylA5s81RUKUn3cBREhBJBq6VWs5nrhMLQpQ8XlgpQ9h8WCQPxyD
cciJp6Lx9GdP03VMiPd+b4bAZzQ9FRLUbFPztITY8Q26LrEEy3T3nkZYg2eNsGIA
PrGWMAqJMPIxn+06IeIUL2+nj1qNGZWKDUvIknn8RVvb/Evme4jmcouUjNa45leP
MYK076krHTgXxUDYMjav/9I7Hau+XC8vgopAPrPUdXcHnBaZYYI/lPGM420Nh38j
yI+LM6DM4+TNQRvYelRiBALen3uaxhJQaCKjmOzmu66KqIJd0dExP9eiUNVnSLWp
S7gdw3hb9LUDQKj/AbuPeFPyhf6O+cxrKgmp1WY2hsiHoz0Xd8J4k3UNS+uu8/qR
UTmm3H8/MY5PJEliiXn+deMbY6vghxtssHZSK+nJDe5kSWsJ+i7YkS2aGZaHEjA/
5+S1ROV3QEN0PPI3GmF65CMH12p7SbkpngyPQQl8K4Adw4RmKx/NPB2LQuoqLpV8
EfBzRgCDCqOmyDpKGkep5IOPlUb5KdZd4sMonysmtlhlEGah5T9yyX06xThur509
loiG6G9esDGEUccCfnxsLRghoA87uTciVuZZFwbAejXbRW8QL0W/jrrsIWm9zTSE
rTQmFKBgnlMBtilxchKm3DfcFqYGlpQeNxUMg9ZOa5kHy2t3iUiChM41Q+3U549S
mmjcbb3PyCGd2SZIiliCw8fuNrQWqqdU5i9h7wZ+JahnUkz72aehVwICFgaJPBCo
exnEGy/o8lno0LThGsYNMU3g2FrYjRCIjawD4ExoQ50I0DnhtmiLsmj2yiM1DYgv
alIxJcwQZk72VnUHbrRpnu0v9OGbI7BsCccMLKcnusYie9ZJyxCjWaCaIcaWpkep
15NSCJmKEePAU6ndQkEzTCe0ubJQ3WO/aY7KBD0a3rPjz/CZizWv2R8s+wROTM38
fvG52K+Tjjp70WxWJoLURTmuskTXLNqlnvtwE4YrARg/A9OsqjyBugMBPHFoSeGY
9lVmxtBezDHABHfc/62cMSjvTEprocAPLoqfKaJjjffhqszQh7kZV/gr1o9T32lw
4n8tMJXXGJ9VRWKiCf4jFvfqefQg4ilJkJZwylZplxlZ+HUWeCWaDlXxYXaJkYsw
fmNf2EKV6Y/u4v23UCrYkkTcSU0lsDrQwwiiNYr+No/E6EAeCoCzMYUywO7e42+t
FSTEl428KOv3lLVITDungP89mEPnADZPaQC+kiZVW1muFLM9WhYZzt5V8jYMGCzM
jvFi9DsCQEN2VEB5dIyK0qfRXmMpwXMOS2SNw5eBgbOmi4mnq21/R9yENtl6S/T3
Q55G0ii47K0mrwEMaQ7H0pXaoa4WaV/mhvNMTgwG1v9sg2CXWid7VX++c2AX4ckK
EMAawWYp2CK7TDEYeae9wKqXCyvrXXzw5/imTALF+yNPoLdXP/72DOJBCTkdPLV3
cWY6lJiiUyH6zphobUsyOCTr6lkp0gDNEEJnkR9QPFykNU4Xz2uvX1U95FzKplWk
yFzrfleNiBOEhkMzwL9skuiD+51vCIUfJg/82F4lhZZm2H/Q0whzp+4NcyIEgbs2
36jNH1Ed3xwrnzh1n5piY8EC/DqitjnLtat1CGX92Ff7VH9gBL4Z7ranN3DkaEMu
ChNkhoK8/ishcYeLbVZbWMLWxqGG9zvaiHbiD32gvE+4+0LyTb49zwA7p0ojjwDF
wv5ILQDpOyflj/PAxWIaC4D3PWQVm3FgME4OPUbH0m4iGtu3IrnXZd2O/49of1Gm
q4THn3kMfOKSWVJ2FgMXqCY7qMwsETK4BohhuwEU0DZ/AED6waUkXdhyqVO1r+pG
+oRseKl5pFDUDJ6yP+lBmc2Mf/3bYpNITKWUSuK3EBqjTV+6BucP5TPxcB8n1jOo
x+jyk1X0hbbbhEEEpHOC1//ak3jV7HUz0SN7JCEgnkuK4DjFtGzo342RnCdSjaVx
/K0gTgLhSvX178cm0ZIzTquIBnbOwUDvcGAtF8dYe2kGlr5sCeziJDsee/XGexZO
hFpo9FAIYNNpB36cS/fiR9KIOCPriRBUOof7mkxZKs4YiKeNai5iCfZDbzT9Kfq3
enl7yOgJ80a2owmOTxVGO/0ZTQdWCvY+UB+CZTn4sBVLRpbDXveEVeTD7sJN2qnw
J12i6jYTKyQI3F5Z6WiDGL+MDbK/kGO9XqgyYY/KQuShocvqkNWreQO/lUYxq7ed
jDXV/Kl1rqguRZHZ74/whTIx/JQT3bHeo5qok1ixop9ZBBb5ylHUfvtR3uNoUeb+
cGIDMAweLpBrO8d2J4wTAKxWoynzG8/oFV6NgpdPFxp3w7ULltjYF90E4xUQmEyQ
UsbacjPKd2YkddivI0x3HyFPHshJVGla+aaa6AK6KqfdHecEWEmy1B8tAhmRODTA
2Xkx2ocnhl9LlxkevHey6I6ZBpjteHTu21qdUkIT1ry098bQH1Sb0Pj1r+B76B5A
3D/syYByoguWnpfJAnzILCtfo8hRgD+zX2pM4r+fYXAvuB9g8u8Mg0ANY9XnNqlV
BjnbkivJY9NP5HzMq+HO1YGNpVsmbXwzFdfDp5wEha0ndIitaUSuXXVU70YBCAAi
OQfy1j9smpCOkCLDUQli9r3i3RCvaoObHMX1t06TvnhrbBy1Sr4gul67gaQpywE3
649+h+baheKM/HC9u67RB6YI0Hswp63elbegonyyUCYjGpML9MDlkTi/woja0udK
dwgUEYfqN+QW+tSILcXD+5V9pa5qgcNdig96S2ZbKXK0p/WpQOhHufjZJ3gi22m6
Klyxnca4+xXhPLJxeTS8IGLBavLCmNcqEy+yRwvtVs7oak/0h3LUfIyaJKRQAqrE
t/vUJVCVqIdp4LsLwhHULPK08xTN89Mb4Czab6/y4mGxKXxPGLE/E9cVuUv6p/xE
lVPqgswHyn46l71dZ3TcGmHOsn2hahizeHlocYiqwdLeFwP5dXUB/jGOI+wCUCQd
vIhjaz9LqOSwkI2hWfg0RALPYpH/QZcLOczcbBs8uIo6ZFs88Jign2WUaXMzSD/1
IWHBwW7fM/GtTNal6Y3U/EbHyTVS0jyMIrHyGv7RdgE8NU5oUL1xaTxD0xLlDHaj
ddNo4pGe1TA2PkQwo0ZkYBSxpLt+ABLJSpfbHw5qunkiV56tYTqkH8iIAmYZszl+
v72kXLbs+wGVMmMdKEUsa/jvH6Wu4cVenm6nrdmEdMmzYMBGVfYCVPBYOUToybYe
es+1bSl7YFmFuw5/oK2u292ACl0f6jx2v8MIWwnRzD3CwP7pIRtTKcQHGFNUwxEl
3zgPv6jxMeCX1CdCbfDFcjLeEBBzWYWbjcNwPb88ZnsFyx84I2DUZxDn88ke7/t1
sEM7ClrslLrG9arLUSG1+JVq9tckbtFhe/iRAOz//sDip8Xpsi6jDyg0VC5DyPM0
rf+6qSIn6DjulgunnziHaPCsmZUq2StaJEsD1uTkFW6mb2rMoO5OhHx5YIaoa+Ll
6auxawJn57UIYIf32hKeOxiFz9LXQc3I/SQT7tXr0K4UJGaQB8WZinQADqYMhFU3
OKOnd1pC/QIMIzOH4Jq9J4cMlQt44gmD5VFs6F+Z7wlVZJZ9t+MhW6/GcbRC/XVd
6MZzfeHW1DE4JYq0y63FFGwoNU+ZIXlyXvu3lifv4r5bnCbj2jMM1GX38c1UkCr4
IGOs9fhS2jKnDqOoAr7IhAdOvsL+jkrCn7BqDHHcg97NeCPekpGY/srjV/y58K/q
9d5MZfsmGdXtu7k3REWRy0oJyuGCzK/BQO0uYrU60L/6+l04Bbnh7cUCVgFP+lQe
QdGAcwCBHFXIvS04iLP/Ogs9henAMQ0t1nGdXuk7G8/2C4/ljqqiFvGvBfjGyH8e
oAEAAI0ICDn4bmR1qTgWI9iJ8Hz0XTqWZR8Ca5Xp4tBhaTCLKT9qfj3KHj7e7jSN
IjlyD3Djt9jAyDuucxCSPqRThiRbROVVCT0DCeXgAAUHq3n8bGzQZeDk29RMraeR
p/6kZVE77Hk0Cq65m78epJf378inGsSZVLPByczqvHq5RScJNmzF+E0lC+PirhNV
B0UQEoNxdV0yfnGvRLocLxwdDxZJH5u5Dt6xzfLZl/6BUrwQtGxH5dG9lsDXsz2E
34c8cNQuc7YPHbA89e3hLa4RrEBM7NqXl59awGs48/MeUsjHcpvkJPJuQvgDZxOL
x5qeOsHrLwrkT+xld6uH66tqIFApqvurZb6AdlHNxE04Bd9zS3Scc8WNOEwl6Rgy
odAG5O7kfFViHNGhsxL8yx1mm6n2rGVmzgMRUTGpGO55WSa2woW8MjPbGScUqY3M
6dxXuSY75BuLupKfeDbiFPXscC6iC1eYdZ4bnJwQ840jY5EZC9Try2szmINVE4Jr
FMbJq2k5fdsRbbcVlWvS44tWFQ32wThDHzPdAcHayQn3l427MoXtiN997gZ/sG/g
eJKmK9fgq8VDVX8k1HumyX9vgrhG2bn2vRAopZvhOychQ6Ud+MrLjreDAyMyK99z
lLTswGabRVYZ0pgcLD1ahARknsyMv67JSDXpuTf8DaDztsUQIE5bCqAhnmq2GEzt
mB34VDN9eNp7fHDZCGfEUd76OaJey2jaLoVZ2D9A48GuJvj7+TBTQlFaA2BFS1Wk
SFONOoQoozL3PqX30hbJX0dcv0IpInFmViqB9pYxBT5swh4mpK2qWCyGopMfo0cA
rJN/7KMe/JlKXcmft7lguQUu5ZOJ0Pfesgtr5xWsTNHusjb0D1GPSqPaIzEOAibB
LGe22Pzdk8Kj1ghUboWtkqRFYzT7FI6vurgZfKofNvOlO9CkoxltRB/nLo+WaZPD
vXqdCNdOPSHBsnjb+BDYL7GQE6v/Ohtiu/BXBT2WyzREjvFu0OwqHVNjJiI7RW2+
4Pw1nAauZlAO05xJTOFMWIvlho4bGi9fhxboOWekXycYeoWau0CGT8jBwHPtGLXy
aXc+DOu9DUdq/MuNBNd6jmehn8Q6nG/MNPtc8vQ9Hn2JXSs7RGqDjBihtoRvvAoT
rEboiFm1Ld7oJtVBKpwaxtSzggBfUpcp6CgdcGwC19JxHSbsnjcTsgiCkHSg5Z+n
tDJ8TDGKj+Dfz2JGF8vyHI7m9vLjPL/280liRrWqY2L+wXtM7FK7D1ub2lrjfK/V
oP7mE9SEEIKnNqHqjKGVCkB/9061X7fWkJ3SdjGLyxY0QJ/Wy+hzCiwzBAuUf308
MtOSke8NQTW+bzVqhv3xt02TLcdp7XwnWm8z3GltzVrTgy2T39saXKfvLqY4INGw
jpbccbAiMvEv1xur0P7KS6IbdKF+1DtNVstOV6ZugCBk6NCeIdHqAiYOeFLsQayB
2TAtsBHrMAVObFrzDZk+XfVQctmbS28EyoUvJOO9YwWJYMbKkvhTjXVKgtf3pVv0
+n+90/ajer40GvHndtbMqM1fC12FJk+KoILYIndBKQNF1r2nQ3mh4lgFJ74MYGj3
egU9BURMNX4m8tADKcbfA99padvw4xov2qWuCdw3tNOD+Yv0LNWBKHgt8yTsG5D7
sJYhPoZZnWSYIK6LiDNnXSie23rFjAL35aJ5pQVyeCiXGOJNdjdMzAdif0u22mM1
xT3gnvJ/H5ugNqzCtDpMMdpt0Kg+1D2M/5uwvIBegiOEZV83V8pjBNES7zD11eBv
kDjkby0Uhh5fJVotOP7E39xmmxUG+Avp37SEKXxbqk1YVM1AGfCe42z4H3fPWggV
2OC1VTzAAAmg2Pr43cE5+jMM0pCQ2qn5ErgeVJRkfBg38BUrQNolS5aR2Z0/dVCD
k1MX0nwvdp1lGb2f8L9lr76n7GiSB+5Qp2mOfadLGYb/xjuxBaRSvqKJtrukGDPn
785frOJcIRZBekgfLFIS+PhZ0LW4HgvGNlnE/SEAytee+pwTomsG7KW3gUcg0buO
JMCeFkkR4fhPMQh5h1w/Mk9F8S5GewmgWcQ1v+wwlobZcx8tp6OXSeY6i1GnR54v
a0dhVmZHiTR1HXLLED6gTvcGHpxFsN1NP6KP2JgYgWIzDtcaMLqchVmCmq0bXzM2
z1zC35hbILqS9LAVp+3ICIrkJuH5J3SEkKTm0D/xxu2eJC/ftFmzcHSrWhGBmtoq
qgctVlvLnRuISyUfwo/TR2nHvE/imiOKJTuhubEsEfyey0OfyAfzGeKvzowrkd0I
8CFi9g3J5OWwRUKFCXfdVIRKMNENgIL509O3yPAX7SVozw43UyM7sm8cLFBBSSAV
adJTLhFL2kn/P94GNHu7xCTEk0h4rGp4r9sLtlYaDYW0mblD9HFNIoZ8dHROTqDZ
WjvMkzHjjmAJZooi7gCAuwGFDr2GgDlcsAlG0XhHz6+rd76o1cmqqSDHrXkojrX9
3dEKvD1Pp9AwRQ8sPydldavATMwINYszE6ZvcVMXBKFef+EetAYauSR/6zB0lZgD
rURoZ7QR1JRsLmIj5MrYIfpUBZUqlJmEo2hs/rgYc8EDd07DHQCp39SuylRb+VzT
XYkuVmdwXfOBLgxMDZHeu71IiRvQd3ADj/4D3uWqwg2OL5nrTBNQxT0rooY4vElp
i/zD85ofk58Jhg6RHPwaa6UZBcrmG+zHaqdkmWnVaUvhsriqLgmC0uv1xkbVbHca
D4+RIkAHNLIKdV1XyFhmvBqiNFInQ3a9NY2/SgSwyGHi8FtIu79pKW88/PMQAK3x
YgDWbRhN9E2IvBLneMZpciCwbaGwxkQTRJ+0RYCWhgMwkWbbJAAb8LSx+MvWk7Oz
i/KMmZjLlhZfFJheXeNtZaR+A/2V56U1uFbJR3OKaYvvxZW89oyZxzQQN37OULfM
UE9I5HG3dfmwpp26nKNgVy0dftXj36I616zbMGQyW1z+8BJVb6grWoyRTHNntwpR
srbdjV6nRnbOI2k9mnQlFwzl5Iu2oGjTCZEdyiBYjv9hB0rzw/MFm3DiHqjtH0GM
KdYFAG6+0L+BM4Ak1jdcuF7/8jeJ7mPKPCDbqw9DDvjG4yxXxBZLirqEc1V368yb
Yxk0rCAQblm9j8s022Yfj9OhW0I4XdbYghHPV5nKwj9s+h15hIukxiPWi7TL17Hl
Q96M7RVTrn4os58gjY6+7OfNzJxZTN/ARgBtWZA4VZdk6VhdgmgmqP3EoLN+lHA4
Lst2On/mhLgns7KVPWQWogmtlGg3aH48qkjvn8txZwZzMxeJ7Ibm/3DeczgF+7JP
Atan7YDh7QjX0vmqRvfoZInuNz26XBxfQ0/HaJ01iN7tGKdUjtU6r2h1LYXNJ3xE
e9IGU7ZSZUyKlbAG0aNDgmfL1jTYAkdgdtlBN9C90H1xEPdMSzTdnq+tfFd4mu82
YYLkeY016cMNoNiLxLOanWPrBd3JST4fCovZakwY5naYVclv9CekukwDzQnh64SZ
0mfKIgScYd2XO5F3FtbYSmkwK39+DZNcdCP2xGdWKxdt+NY7lNRMxyeY8cZTq8I6
92OqPbVsfAnXJ42xmOdOA61C/hUmNc4qmCiymiKmNVwNwHDEGJBe7qz/CWTW3O/y
8pLCdWoNPT13jRNC5WXvDvtJF1F9AbTXjENxP67w5h+T3aKNOCQH9LcwAexYkXBx
MRD+M70BNdvMgXLNaTdav2Cy1ESJWCRhmxkEe/k+XQuoG3eTavuSVcqil39sHYj0
OzJq2laPRLI010QB28uAEVfPGa24QqLQxUCPwNBK4+n72M6d8qH6p9QhvbgZ5iK6
VfzUzVhlRijVp2+m+GF2RXYtOk0Hh8wt8+fInMGDkw8BmEbAk6LSyg38LNEQuRyL
vbxdsoABwBexux3hREgF5eHp1IW/J2F3sGd4tWyd444RiepdQPkBxssL27sf/Vdn
tV1ujH4xltDXEJNZWD49CVq4xk2gDNOJnyb2ZKOnlsTR6rXuhY0iuRIfm2b9GmNw
aSFdT6g33eRKr87cbDVkF/PPWdEZX9jKRMYoPixHwKGfW7VlDAF8Itm1U0lXufqL
nsuUdJOtPvFjnzYJzxK1rCC6vaTYO0wKkx7s1uQ/5kqjYIZulPd0EP73ow+5LeaZ
YwuoFq0MyDmrQ8RYJiya2ivaR994C/STKf5jgUwXNIdYxi/tupG5Htt2XftjThC4
XqbwgUzxrwo4cy53kgm2edsCI/biANUQWpuNh7Mf/lif9X4rCG4AdQOrd8U1BDYE
8fCbaCxm3Z96lS5xjuMb1I7iChw/WEwc/ULb/4bdwhVScRuaLqehc4WaqEuQEhwX
cBO1szuHPourLVZyXvdUv4WDSOwfP5XONPev1no4wS46WtwTECS2oDB3/qO/rO2b
pMUcuUsr8YkfWBgCxh6HH9NxALrV9s29uRAC3ybnjV7bZ+4ZMBPW7h8MIImAW9kY
kjY7h1XeNosOu6HMYTdJ9G07rRI1s0Uj+r31PJwHU2JXG1XKke1JgvmNJmvKF1/l
I3qksx0vWz5K89nQRX+OlTUUdG0LdmUtJnV1XsE7itSYuWzZRnUQOPJ0VdaZIk4x
yKebGMLx4Bm+iSs9XM1H0bw0vx1CRrovk/iYBaDknlZWjPWcsl6xg2ycwD7q/APT
PXi8xArSYxx6+KWHNeBC+ojpFgQKBrYPnr18H7i/kpESZ4Z3PxKocqi7x+BMviFl
qXN6CQBozDT9RXCbEidX44WxC74ss5VQUqbdWuWMlwU1hLdJpTZqHGZlXMOxP/ll
Vqi6RjVAl2SLxwaBU7xmqg3nxvzATNfda0gITq76gtV0c/aZ3VGEaPFTkxeOlAex
zDytVONIf9zozgKqEtQFy367Q2HvEAq57e4oVG763saxIA3tSB44O+xkDPEELLHv
k9il9RTIRhlTxP1bD4I2W5aPBJxlzpf4sWyst4EjhvyRuxdl+KatgS8yvBbb0Ims
3O7G0dV6pSegbW4dTTbXNLA+LyOOKCkRj1pCJ+emsfSpP0B8Bd6H9zzuah5nl/S5
dvRKMClOigHt9ahW4NIbt9iC5E8OJEdfKDLUtlrd8U7fHOEcBHAbM0vh8Y955qh7
ecILEwLBH7BerVoHn6VPRztV9jDQzR1nzjHrmSIZVcQ36iAkVyz/ddT4uuqNdWtu
LoOEiM9WZKOVUKCUvtObV/rbmwfrfTVYE/jfY+LF7kGJFzAOKb06xaRgIkvLmTb9
Xdk0hn9pLDjnGhTjmuTMb9ZyK2ndrebwS8LtC+bfyLXpmBbaXUCrzTfbz2/iKSzi
iGGPNGtRgWOp1UDKXvRT6RGBswCNA0l3T2+iBjmsSz2OzcN3zlGBx3rSSrzcGTL8
zszuAORGe6ZxKgNrbBqYhoBtBQE+Qzigkg+SQDIWEDfxJyri2ZbOy6wRLmZzYpm6
rb3PmyWtSe5fAXRSGxasJiyYtVz/mQ2aTKUG1UjEOO3DldztlEHsoVNMbmwMogNA
35HJu0I5YTfgb2mcpm5amv8uY+Jk6sdbsRgNneCHmL8s0CoLYMLrBMXia4LmKG7n
dL8GnBsR+Cqn+kYzvSKKfSZfPqsMgKwDxL7jCV6s1XO2qi/EdXyuZih7o4UuzdIJ
l8cw1a8BrGBlo9wHOisp0b7WJSr6/2fTRiAQKJdgTaY8KeJ7044I1JWEVzuf5J+Z
RbvhlnOX1qv1634OCue3t7rjdhG/bOAXk5j1WfZSu21Ou7YVAXL1JsURF6lEzru0
qES5PRy32qpTYueFEWK4ebGCUDLR98A4IZU+fXCH/G5SiN//UhA/Qz65QBBvpde+
qcyCmKhZPve2OQPFtErwLib8ezz4Cu8j5WYRNoTsWZ8CKeQ2RUGbLS1oX5dUKPgw
Wruz6Nx5LqK9bCtAWdbQNuSL/u8v8d1xmsV6LEe3OFtfCUxOUBJvf+lrdm0bkuub
8fEJhQzPJtSMEmMLvNGTJpGnIBheG1vBqCvhI39EXDgaYaYoAGDB6+rN3Y840cr/
2roZ06ltn54hE1KreoXAEVN6ljEUx7FTJHupffL/eN6Tden9i0urhuhdISIJMZXV
QhhsOxCD7N8NjTqX0sHGRyaw1EOGVksygqcBNn+DWtNVyWz9ba3cBVIMyxa1QsZa
RwrTKz3Vhz7dZxvsaOFw1NB4inrqdC++HMk1SExavrs6sVoWN/Bz8TJ1RplnvT0U
9PU3OCoFqUSmDZo7JSs5uIU4KyhDFs8Z3cfS0njXBqKZCIro9OBwwiNfwXlJKJRe
eK87hbWTzc69x4UGehFbwdtXlBPsqDvoK7LG+8qJDJzJHh2SbYS+aUWvqPLGOU0E
Ze3NrqbjA7l1HprAAkMDvad8oI9eQrMo8yukPaDPNmcCNBVlKNer0K0eqGNPpMqK
TwDn+tuBLAON2/vgSr5+ghtFQHGnDzszWnvw34nRkRikRNMetDkSwJiENl8RyZLJ
KTtobr2jR0hL/dV4GdZvgiA1hBBTsEVnhAeIe4Ly+LRBxjjPlSBpQJKL8BxdVRum
eji9LEj9f7348oNdB80Tip8ipikhDMH+HSga42MDCMH6TAJ+GWI0AIobs2fvpvEH
AeE6dj3nrRB6RGx6WaO9tSbqXBuIUNwrZMr+EmD3e4YNDAxg5NEgXvnkxWi+pkyO
Wo+1p3Ju6vNKTR3N4AUcGFjIXnpAZRK6YP7jlEGMKT/KGquvwceGX5CnPADk4Wjx
fJGFqSK+wByB7qnkN5OmQPrZTgLDUjqirlhtPOY/maHWrvgg0KRZOrSrH61SuHVS
ifb3CEwI/RsTegwhc/74ScirEBzgcxFaJxR/8Yyy0VGQTRsHm6kzTIA/sS0Fi00w
DZJn/0dPECu6p9q47MmfrfQW4vr9eUlHiTYLjTUmuDI40X9fu8CaLIAhuluRQaEs
CXzViIYKcTEi47YXtOoUo/HlS0szGwjL1UTRmpzfI9+xA3bGzKHXaWfjLH4TJR2z
TbE+90P2eDSvSs9x3z1Y1xtVk6DplgILWVQygyBxmOIXrAYDK0CuUjSoctRAS8ry
PEolzUq7gsb4bK83ATLGbXdFkW81wCjmge9ZPujx3podpRkUC9FN6PjPY/MHkkbW
JqHlJCrAAqJDbgYBhnNxutV02xMcNwI6DwuoTv/0QDJ1kaSHw8LvnepkFUncMP+Z
SYuFVTZ+vUr9Xx9YJ9VrmSPrWcPFJRh1OPPCyL7yomdvQCXukaAPYcJ+Lvmf12RG
qES8wQLaEa5kT7Y0BEdsBb826IYoCN1vHCOxzlNm8lhSPoNXwrB2qrm+7/vVoXeB
9c/lu77hqledu8vUqV3KuXI8Xb0PFFZEWGLoSjt4w4XEUrA3iTQHGXU1dpgR/Ij7
fibebvVNZjm+WICAAJ9EzUMW+hoA64WZa5t6Fj2Y5PZ4d5QM0bWGGuULQf86XQhn
0tJA8sEdEEmkBNHByVqSZu4gy9f831MqPIUxa8qZcvu1DzI4aL7rYDN90T6E4o/C
lTF9JP4yFnR06uVnRRs0DCIBCxS5SbKK/x9yyceWHWI60aDDV8j0gnV1Km3P6HnV
P64IDDR2Z6nKGxw9rwmBhg2tBcdqmZVQuquyonAXOy5gv+//DTjp3zqF0+PoCzLR
d+Ut6kQE2Iv1Lg8BHlcPT1sNvf9Sw0u0t5ZetnRx6UbLfc4ZgIq0amHF7WQ25Kio
feYU6F/SVUvVKcJo/Ns6/Xg0NLHWjSPTRjmxjndybCVA2PQ8uuNwi3loSMdniRjK
7up6a4sSmo3IAzf4GTOfoFP8Ie0mYEkV9iwJVLW8eXC4kNSypX3adUK2ulN1jWVC
lwXYkoVUSuVEZOAuU4D7KbBLf7uxAjyLEJEB06lGK9Is3KNID3yuLHmRMv1gNAmW
MDteFA0YLYN0v51yKBEQjv6yw+nKn9P60Qrqsqyy6L/T/zClxElDCFFOCgq6NuEn
Bx8brfS2tJFkU31xtfLF60giyqj5BF1SPvrtbnEUN4FQ9J+wW7+kWNzERsBFpcHt
EeytzE72c3ogg8ohFOe1ckqSjvINIRrbp2lsRc0BR5nbszQiQbzr0E6C0Ad65kzb
5Swa37CHrkhFP8lNXsyohtukTQeH+PWcGz1tQvozrkl3gFQ+JJX/Ry1Pq1EzN6BK
+uvYrkbFXhqSFaWbkMFstIAlr0z9ndh9XIU9vTURc1Qq4Zn4LgA0JVXUSyX+A7B6
Tig/TKUy0lXaacyjyn2uoQuA0OgAVsOw5PxUZ+Oa7srnT248ntg+uBhSFlvGy+Ed
ylLjXFaPa8ES4g9IKev/giPl+/RxNzBE5Vwvo7cJrunttvL1XlTTuPBn2ENPEZ92
t8qypiOcaB9SljBQ0djcnjVw+bgIrU1DW9iDT+cI/GL2eeYxPnjOMa9vaGovrxYT
wKxLTYu+oARLuwYNHSFxECzikIWCBJ6NH1kYGb2CE1IIZ2woQ8QPT9NNxfPsZfbp
J+JoJzex5GBG6Q0iOYms7BYmb+qRJAVMlkcFmAf3DYucoWKcVA8GZae1ks0aSqdE
WQKXmVh2W3Au9X/K/OeME4+SyC0bCUzWHo9iWJRw7UXK+zVCbHBTsi+/vqtR9t2+
t6Jh3yovi9W0YdPambWpnz+wYiA+XxMrzL27O1INXU9cSa9U6YPeczOiN7f5CLwR
hmdbS26O2aeVGr1R62Up+WijwzYeHVIu6GYc9gZ9fq7noR6bvfc/gflsdofR/4w5
ka9/icHZ4+zOTz5/6nyFacWYB81+oJLpsX1dw79P6lUqx7G1ObXfugVY/BzybJFA
e+g7CxLT4JoMF23cpC/ztKHuuPY9dCudGCpxZNx3QANsswacojGtit2aGWk9QXPf
T/YIueBpwXWqUogQo4RkqGyqz90UgAsGYb+PEnAoytH2jZPFWBbkLpj7LkPjMhaz
QUH/3OiKaNbRbUJ2MSzNwPCYWsoCS2xUJjx++uts4lcm8GcQxBVyoItsepVP0YnF
Gfl4u0LTtvUGoCq/iqpE+h+uEP5fl3PP7c6ZklBZ16flRzvZX0AedswG5QwF2T36
yoUYdlXSM15se6H0MGvu1sXkaVMnN/nOoA3eN7teVY6bQT36dAvh2FKcOQAmQlH/
70wpq+fpxyIydh3iSlBafBkUuEWp+ICKJxYysO66pmRBB2kI7j21rE00h/0mB/qW
cPJCb0ASzAZwwc2tvjlOn34RPhA+8p2RbWDE9S7jco/7CecaeF9JUwTeZk9c1Tsh
L8V8VKOXpCKrwZn1A8JyOYN1wXE7QM33WOlRIUhg8zA1FoX0+v/WUgczZyJoKUjk
DB3Lm49OS5Cg5i3LDUL6tuDuVbDoIOwPSY2QN9eYbdkO7Qmcdjaevuj8A7SHP62W
RtPgJmke0qlzMvJ98WLRCHRb8vPMXVJqx1dK0IBWKYR4smzADwE6HbsHQBao1+6z
9Bpf4a6UlzmVnm51QmbeQhlPm9BxUFjj0wdYPlmfEbm+lFESqxafbZuZwxyA9K83
hMOUVAacIzQwFHJ10ZZ1NCGsURmygwZSRNvZy/jMPc54FHsL2J5dfM1ef3+HKWPS
Xw287xI/aHJNchxtIGe06V08QbRjynHw9taOvMryIvZWrp8FwXxyZ1yNugSKm6TC
seO9P8B6LS7QFJgHJYSr0oIzVDfD62cgi/RrQqjJRHioF0/L/Fwstaw8hXJEkoIQ
DOLJ6hha73qP7dWzE5hggkj76uU0p8dV/dMfufY24oAG3jbSnbdjWAMYPveCKTvJ
+zn4WN/Byn+ixFw+GaDmiOpdxwLkncCwFg/SUpfrH/tH/hFeaWlhqyt9iDp9TPY9
0Z9rZAXQpE/zJWKgvjBV3M8VQMn9VumsIgH+yVK/cSGTaNbT9AlNDwiugBlXkZpN
xopO+/9Q8EpQ9/Oo3YhVOZbollwnAjmVAmz5RaeXmQ5G2pEq7kelriBBmz8jgMER
GD9LaNQfZ98ea+58wL947KfF9pdAAGMlWkfzCIGdLvmuaIHF0Z1flwEI3RSO1efs
x7Fh1vNINk4S4TfiavzfhL+SlUSbncPkSey5fb1jcx4mGAEm4DzI8WgYypUMIvDR
npwIGqgcR9CqYG9leVycPAq2IArupONscxCGKFixQ1Aee6IPVCUsZethvv1ircwu
0uCKsX/CaWjCaRcNhe3E60ewe6tI0+tfoTzu6D1iJeTqDaNAsMqJ1tmCW+UNln0S
1oP8/JxyItti3VQoh1h5FG/nrtCj7ecH8wioSVLvixmGQQbJvQnW+er/Fcnam5Kt
TVtNgLzOtwremAXedM5osGohL/wBoW5xAcN3oUMhD7iGVavql6TknhrwxWHoK8+K
NczqRDQW9DtTMF3Y+TtTOWT4VUyhfzkPyp/34znJllGHB1ajlLpR5bwXtwTruGWO
uf6FB56wpNxolNiQm2A3p+2gcVXbxYbTsuhT8cijwrUNF6C7SCp0En4M2Mpp51c2
CE3WFmmvDaDveW8irjqWf6ajgzcugP0D6+qTbbCNmPDnG2jnFwTi+mzgCCRUy9GI
NmCw2zbOwkO73P1Juh6JD9IK1vBeU6CCl/aMFBAHvw5pBUxH3kf0lyeNGKHW4we8
WwCNGGyBFev3sGYn+zZrpQ3IfB+R7i5zCm1Pkvwn87OyUJMdJKZ9K7hF8dw1Lra+
379St7gdVnMxp0p9a0+d201pq5vET7OfnyhpK5YjDKe3DVuehrphFydYdxlnoewa
Pz/exfYQtzi/xj1KZz6zjpIum35xH+Zc6GuTpELvOcwRlLhXRhfKKCeCyFUvCucG
a9tikgH8MDHSPL9+WVQv0s81BZKha74NnzoofZ5Wn3KvynccXBWHsrouykv84im4
EI8qZZ7nrqnKRBuk1sR09UEBxfZADevBl8/dz8XmKHI6/r0BH6L8O2/GKO0ahELS
eg5EUAN8orlAXEhmo1LJOTn0AfloGygYVUAjgZ3dJ65IE/7IFps8ndaB6U/ads4Y
OaIkRl0XLTIXe5g4ZCJ2eovdNN13AXajY21gBSp/BGNVtV8lkx65jMav7oyLEIFF
3Vazeq4q4ZVlPX/A7GJe9lVBLl/EBVCoYByOo9DrdyZJU31kTLGZ/trzPyrJs13w
K7PbSuwSm+8Y4ODL6iPzqSXk3gXpQDCEfF5KDny4vtkpPAx/WsU23BH316f4HLCE
ct2icnwkLQTXNoBaxSdifKB9blHOW5+ACCFaW8H3prOWgs5lqLnvDoTi3fNeEHB5
p9gu2Pg9ShL6jP6YTF2nYaH3Ey0MIgN3l2C1RiQ+jZpU/4Sw0xuU4uDLQVlezonZ
F2BBHT+tNeSdGGNOvMruYkbjMTLX6+ONXb30kGa8ojBLdvH5oKBfXIs0hBEOym53
DDQ1x7gFv2OADGDXqEA2iUjSfFpnRxBmodk00g3pz1BSFa8iJVEtaNOVjivct7Pl
aboZtDEiUqXEdFDN53iwEpP8O7jObEry7SYBPdmGMGoKCf19L/5HhRzTuASGCeLn
V+qN4X96fQDCe3ijGtGJVNLMFz5Ge77QYxcSrlQlqRvCh7t4SwP8tesKoek+qMig
Hq9CgK7UguvbZgOiReUVLC26fh//tBqGXGAbmtHox4YF8L5utEvhOtV79Qxy0F0f
eX9bncWyRJiMS+0PAnRHI2E/eJu74yWqxicr9ztNib9wC4bS+wSQtj6ZsGCQ9edP
hhKZi1cuVbXlUsaio1sB7a2C2ZJfGfT4K3glE2OCmu59iRVorBRDYEODxxo5PiTF
v1qbGg7Sge7SBLBPDOxHjimdjsSzogavpkPMPXPWga71fjsVotSoD+5Xz2hwT0qh
eCXshUStmBTLuWe+SQ6VtuPfxBisIb0oRIe9w1RR2/8+7JCnyIM92V386tHH53Cf
7wbAeEOHn9N7spf4yeW3XdBiNxCB7YkurkuY6i7Sx48ZV9BfMG7KPRytG+cekQc4
yqBOttH6imzkpREffs0uQsthOX239Nc0kfThPWwaRoM9T/xE85cS25nR7Lpsd5NS
J+AbProCvOFo6ClpRzYf/NJkA1hcB+f1/yynVHXoFQKsLSeatYbZoRcLhqUIrAph
81uA5LRkRP5ZQrIcwLpebdL7OGuTPyXJ1jAuGyRR2IRzFJ9ASY+tRuwbT5o8fZsX
iaE5GKvC+PpmRnP+CcdA6f8B5ZBKnivetDYLgwVeAAtkRCVbVKV6EFnE4tAtQH2f
7YxL001DjQbKni5j/b60KvbqWVBENqg0TmzolFHHRKYQl1cc48cPvChU1Jpz9gD3
12CYyNEbTfCOqYAgtD3hPSpOs5YVvmK140bRtxy3Q8NPiIoW7Q6jT7YiZA60v36j
s6Z7ejGE6DKDJfJyEgjXBtAQjTyLv7cBPAE+IKXg7KgA9yVYEq+LXR3aOHx3TlbA
GZWkLPXLHsnsdCw++f0+merCJjmebC1aXreSaqAbb/flYe8QFpg8uvSnrbIVWds1
j6MOcnQzV0UR4WswtG2pGDoPcjcfYtH/C7rbsdpCIoaxijp4rxqTgMoXkOgaHwZg
4ij+8lVwnwWO7s0x/60EcfeI+cuD+QN/4z32f4HoWPApdYCeVQP/g4QdrFmPvKCY
ghoY2YQ1xauQkK7TlBrWBvFMXR6KU+LzmJ3xf1MrPon5A0K8LReOdyNJvFwSfTEZ
BSeEldLkEX/Qdt0FJwZr/f6Q8EyrEZtBKerleWwZA6FvdQyqs77+OA35spvXhlws
j7DGmytxrQEnLehmZ+GcjVvgHSKaNKJx75DUsWNfRfUZhvyF0Hh6MZcg85phaX6T
epsNLfoV1HPO27LCmz2IxPBm9dYkNxV55XDEhGiQZ9YxY4ZvzmLjMQ+VppLLc4/O
PsQ26QexhUZ566QWS2WgtGunhhi0Ujn2qoPKcYSMD28J3YtD52V4aJRDh9ifxHLe
Jico36WILHJfGEOG0tQ9uVZzPif9DOXXlQOhmnHqaC6VgdsjY3q2c89p/O9YbIG9
uCSk1rThm6w9ZnfRvRpV5OOT/PFr2stZ/iJN2O3ppfk+EhHIoGnt29lMxYx1/CGf
nA32dOuIGyKMrfXLbI0pm5SVubut549AG7ch0b0OV9X7fsuP0svbkxkqisMpk/3s
DOvfEDSsT4gv7peosB3H5XQL2udSS43vU/zBAHsewKxUu3NrugDwb4fyCTLGJecd
i2wiob0PY74+MwpcKAfZWerJQdImDx0cmWvIKGR7h+H9Mb3CqorwMCk250v1j6G9
l2cYaNcPAbfY82OosIV1wbExHrX8xemVIPcs1X0n1eMgaHeR8ICaDBV/ISOyyl/E
FCHO/9ooY6dTUcoDIdJeC2nb/8hrZMgRFjaOLXfNDyJ2qbxzjThXNMhZ7fQYoPUj
u8SVagdEILbDH/M3j8oCKW12bpl8WKPzlrHynW/Dh4WizmdMVzVEdM9ehV/o+/Vk
9DS+ndecm8lxkZRD87+EtK2h8gNTC4W6PUuQxsEoJ9cz4y819f7Zf63Ach0DOWmK
wVH/c95MWrkVx8d8h7fwssOtpbUdrQY8S6INsCfwjkjzZ40RaopsATS38BUy+DWn
3vHkA0OKDdAJj3YjdPWd9zZKTyUbn+hHcs2SpayY/2GuqlOLH2GfBQDT2uOwud35
ZevnwdNpMcnhkrOdkQpW9BvUSdaoeM1BTg8VTKO1Z5ohs3E0HNUlYC/THB5dXmF9
QFsFHAaEX8iXITbMB6LYiPYZW8JpWsvETnlTv/FeM4hgZ9dwZcNWSDItcnAUTf9n
rYXNIt0PUKE0ZH43iPZDDZf76GxIf0TWcLu/uIMeISg2YJE0ffUteycTGD7PWQnl
SGV3Pbf0Wg7gTAw0y2KaZgVahBXPMwclpy07hTrFcfn8Y9vrHVzuak7+o4eBWFyo
pnTGh9QWxRa9AktBc1K9cGzwi93WiCNANfjo8TSzRiiygpswwup6HFfDcAVY1v51
f5MJBJuYPaY5mIx3cbRgsHJdtzSIre2Hbt65zMqo1Qea0xVoxjWFNbqh1DMNtuJd
ljwqz4fwM4vUEXd/ZRmd5GUCnyUQwy1ccYVjmZ1bcC8J/8JJ9CsTMVbRHoVQtqsO
hjXDUVwltsFiy3kZUxFI6g3YwXBmdHtJEoBmrHCQjsVSCEpDL230AmBhe4dzTNXP
501lw/eRqroFYeFruRJ5U7wm/b8SzFJYbwjBBL1tHOveIYSkhptZwfL9ixZ0TzaC
LKZHH7+jhZyckKnVDN8HBilALBX0M8eHV21C/S8YCTXz4lTHI0r04XMW1B4AA/8Q
ca3tEoWbKscweo8dMME1w98/5qwb74l6K9E4GC/lLhzNMDxdK3aVJNr0+c2bpAK7
gVRjLfFWTemaWulfbAXyeplxJMqjpAzXgpZjzNZvSha9RZHbB3BN/gOIce490dVh
FAJlN0uzgVvkxPLhIOj7JFoP2uX9xYYqiOumOIcUl6CtXCr8TFPBGCP7aIacjF4f
vNXtqsBBCPjgvmwFvJjUYUDaronnmnDE6RwXb99q/HESo/M951TY3UM5xNizqKgh
hl9DklfDsYtZXlMVP4ev4eM713OJNt7A08TFvYshh18eGZgGjHnBgd4e5X50HGrL
NPWzuy/SeBX2NYBDb9p3ZCK9SlI3jC887QQcf10xEHcF4yK82os9FMxeWLaBRXsk
Yq0wxdMjwFfwzE5C62SxGzSwzg/CHnruxH3T7aF5H65ppDS/hkxweIgzHwnDlaG5
CTNtiRowhO2mFU3PkRmTqGjbsOQMcms0BTkn5dgJPLUU2HTB+BHFs3M9WxhBh9kw
OhmIdNbdttJk/j8P2n1f/yEGFDbxPXUQVxo4S1GbhYnXjGHZrIMdJTqmhIYBNKXR
DUGyBzypnpnN3u+b/UzvyTg4JOvXUhcB9DdgEG0Z6mCp0eHi4tw+UZTnaVPCVz3X
1FxeAgV0emvyuAzeND1E7snayfp6IVvLnsPNGL7Bx6Nx4l/stf7kW/qEYuN5feem
0un/6ihzIih9z5OFP6mapE9sd7QU1+nBXuLeQyrBnEiSszv18gXpLdLHFGrPLiCn
8Uclsw0SqjbnuWVx0LmEYLiFDF8C3n1O0r7GNvvSFwy/cP9aHGhJV7/Unr8lm8km
vuY/MfptV/i6maVqFRvO6UquNmQJcXEEm4K1NNwaPbFpcScTz3JT2jPps+FQ3DwF
FFOUT3DKsQl/E5mwDMMUOJaDk5yUw/piJRC4Z0h4MmfruEKTwJizymzXp7jODTxZ
GYXWlSfWnV/js9KzbI4N7/WILs6mi3DVLEf1pLjcTdRE2pEmiHd1bT0yxrv+36K6
wdlMgGpdFWzET3A/5LhXeYvUSK4FxAua/6rSllJZAP4zka2DEiRWL3RX60sH+ZrU
THEY5VHCUneFNRAac63vNGDd+l7g5Gl8gRsrfn2y3zPFKNZObgFatISJ8EVfPTRW
kOK/KRgYohESl6auMRLA/ln9SVjDt8/YvxLMoct2N6qCe3hEKvvi55ZVg1EOmycu
tPHWwJlqiNIfwVVPV8UgRzuavrf1xP+DAIvc2Mb0F6Bz+nDk/p1d9N5FgnpvZv2L
Qcs6/lEGbak14oGEFXPvwKlG2BEWqUzpyZae+0mNPmznzEmJomJ02Ojo5GU0oOe7
wuKqX3/qpcer022cKqkcXzbxIdABb8pEFuz4lIbshAKP0hecNQSz1RKddZmzahvr
sW7379Ap6EzgDxQ7FdipsiKtEjpLcok8EQNxgeOStXEscr/NKvu5fD1ejM/rTv9n
Znf2e1UlqALLVhUdEwzKN3c7jSj+Ci84uEgzqJrskcIZIr+6nWBOuxIyFk13qXWH
yNarVIMireMAxXlpveMG+sRjUObD3Jdsc7oa/aVmbGmaTO7Ihm7rf/MAlRk+m17t
S6xqedoC29NdbCBmUP/jL63wT4xz+Dk3UOpMfgkqVjdbiH5TSzFe8lDR8S5LEC89
W143bp4QesxYbWq6eT+EqVR40CoJpf7zjc+5FGRv2q9TKswgjWgT3gc9cf+3b8vd
kTYvzyc/++zmSyR/DIKEma8N6dJZvXpsm7um22n6IGhRNIBx236Lc6Z7vMrdXq3l
/NV9s01w3GmtcD7d4rMLhXpF30NZnoo+8qz4rfX1gqiRxBLk2gWJXWYqDOvC6Qft
ALMkh0gyOuHzu44/Z6cgkPCGd3YMjspEmSsNuWDJijhJKDpHKnCHFUPFNo0q7md4
Nslc3YV48FYgYd6WFUoUm0gzAKWXG9WrLl30YPPVQpswXoBLwxcQRbPctjv5qqqJ
PmlRsQoV1DQuP3TGwpTLSzl4Jy/AsxJugA17pHYEmyP/xr8YwMcI6jU+i4UT4oQD
EIB2W6UR+SQstLXjFDmdAZxk4HKYCTw9AzJIqefI+MUi+8mCAFNS/JlX5JSX2gM+
KpueT5Xhcp4Cx/s2PiBmghDf3oBxcl2Zbjs94fYGOz6HIju/+/5ycyEP3Ejml3bW
SCcJmmWTb9Ju1w3R3VZGvbcKCWF1WAZPLgZvAnHOT7GEMfKa9LHSljZGbgT3ila7
ZTAQWVDT//UCrjIPdrUCsr4BnT5GePG+yhQlwlXKqUgMFLeKFArgC6TmYtDRGdmR
2PtMcjNgHPJgTOvNOTf0DXLuT77HviPKjynBW/2jrWL3W2TW8qjKtlV9AR0mma9+
03OWhQ/AfbhZ/hzPHfSRockGiZhgOywqQHZUHriV3iBQUk72LSjORmohGJk4coyH
J9bzKGd1fmiZ5DDE60pXY3tXNcj2jtfC0/7TeVbgdbSAsPHGQNobZf/OuSYl6KeJ
afc/T1XVLGbgfDMaQOeL18x8/bmzTiL5u83S9KAYW9tMxCAQVsPWL2LVl22YwPld
VH8SmZ2GePXJ3CqHa4t0C/qAJWqDY3YVakEGBpMrZgNHeGEIyXco7eL4b2sBP4l9
Y2hqREzj2LbK+KnpPlvvNu6pZMgtao+ayOSgLGW8wFG/UnojYoFPEkcrkuJkc9Ar
lwlV6tmp+JjsEimfTZCiyqn6jpoTw8eFP2aJfzsiXlg5Ya1kdkhfuqD+mkRj6JLO
esVedAUN47JOcDp5wEucfIFnAz8AP2d3dcupZ0OtWHaE5JX9wWqeprMNGgr/uFab
2THW1pyRVo91DwPFA5OONkZ+D8uc6v4z11Nd+TgAp846d0Tj5VsU6YClPWakHfZ6
b6GmfzRJ/uF+ANo4lcvHBXG9dOcrjEUZnYBCl7gJrbJIMfOV4P3GRrdgcU3NlSZQ
1W0e5uj3r1K+5/VYHq3mTqo2npP3yAksnwNwPSxEs7CCQuXmjgyWngrUw4JMQU2S
EpSii4E/CJgienWw7gHJrr1LvpXCf70+JuYMXLPZo6TBad16W7iQX9zHb3V5wGCM
PJew+m6tvr82PpvkBr8auHEk01YEHeGrW9a9jn1qyp5MZfvgm3Mc0mOChWVDwavD
/f9PtDSDCfpW5uHgCTY8LPkPLmjwP7huJe67mZH3/uu7rA0Kwi2CP0uB8jiRPZma
HeJ8MhpBStFNwL/lj4rPBvR4nHgdlkFosayv5BKcpliPgDYytSbsQ0VaLgR4PbgR
jhjGiltouBrzcnslCfoAgvW2iYFfMsgyJxGpecrKguj7lKzDjAugcTktZ7tluxdF
ITzAPUh22Dc0Zx9lD4Xl07x8b4W1tVZz/qyqMCYh6+Q94hCK6a868bVWlmrh1gf6
3xAAi7z0hBfRAnBvZsCJTaFZF6ejicXd3qEyWKvC33XWMcX7837qAYXiR+l92iMn
w/1GnRJNnOipfEFoiSaHDjQKZjCWTDMdgmXiYIIbUWl7jaR0webgqg+QgGH5rNN+
n5AIz3R93jC/iQM3l6e0psnvjhhjmcGTeRM7bm4m0WSRwM+V8u0yoiLeZjdEUhq8
j80VEbFwT/xCWemKDfgVjU9OtHWS4xfcqCim7WIGOummTb5hELUUnSD+8ud1adm3
jbxQUiSjYmZA0mvfIKoUYn5cbrefnBGEr8X4zKONCefEPI5J8/LAgDGeyjiKOJKF
z7PtfUNERzEgEFIUsuTOyX3BG0E8tR0nHdYer1WSJgzowD7EBvITHQaJphF7vRyc
halY6HolaTnLA6rdcxXQvqnREcTjinPrFlwKnh9vCAtqvk+TYrE5jvuqAa7DZWSv
eo8/I9tHrZYZpMDQTzydarFkUmHeBig3kxczOpQDRKOkiyroo0omVF7ERKoI0vE1
bNTCr0oRfupS5u/gBL2EHv8FM5NVZzHeuni82/0pQOGSx4si8lsihdqzlF4ACEvB
2ri1iOV2ImoWjpXlVU2KgM4Any/FeLccxFXmpdyZO4pB/gnoiIp/xTTidIfNJmh7
OO3xkX1vuXXVYOHFqC+tsy1eiPL4Pb2dRqgsXRreXW3ffCSQEsFqBWtHcSfDN45j
FPPjK8efhNaKVx9Ko3u3oy1N8QdkbHG9bMYsB1zAgjh+V2SwrDJMYhQhc+PYIXqS
vjojrGYHrFbSF1pAjR6XrX2of2STuiMwL4xSPtm6M/876OzPdnWENe9gjvSPqDk4
dw6L1Q2QKbNXESrd1fakwBniQF/VLyx03l0dDqekvU++Gst/m2xlf0XyCPtheaun
xnGDvcwlFEcs+BQK9+lx6+eB6EQUJdyWXeyqomuXy66pQymeSkXVU33vr6kL7360
xomgYHQet0NV2mM4vRui/uHF2lDuZBojxpW/u+LAoNMFP4hsoe7yrj6MdUi31SAO
vSWny+Kkhkl3T4iI8Zb4bz+Ka2ZWM/Ajd99t2qY1wIgqL47noWJYKrja3nCvcNZk
6DqJ3/uY0i3mKmlEBpMzLqH0Gqzt2tjHtwYg8516p6ZWuFoyRhUmHGgXI60Pwkd4
pT0gzr0zLFR1YeimDCJzv1yLbi2GCpPA2Ve1lRaaxGTMQSea2GPtk3A1yvpAsTAl
U3uQwq2hOztKDcEVPyXGGoJpItbkIXD+OPVgoIo/1jPxInhhzWiiSz7hhoNnV8Jw
UtgtX7ZRkLKt5kxdshtvu+V+QE4DIP4/IykXD11CJ2BkExgm4sYmI1nV+PSaxdIG
YsRNxiu93QYpJ4bkPby37gQ8p3/sp1QM0sUlgmzpmV5d0EstEG5pUnd5Ihwzk2p5
D74RAhiFp9YreUEbaBJUr2lIuVrjj7i9A+CrstfiLFvGwQXY/sYZyy/GGKXraK04
KqiRVPTFEvl4KsekP1/bjyrZqmckAoj1FcGLotkLUHaOguI6UumXElGdcJnL1YUw
uysNr3Em34l/vGdiC24OHYTF5oKe1RzQmm6EhccQNjdBb5tuWajd1oq6WjZqNct4
0tfOQ2lyNM8irVPVXIXyT5rq43fmlEKjcTV1kdx/EJAzTTzKZMJsnt8bTF0AiSH0
xTKGDB8JiNtuCaDdVgzofmjLy1ed2Kus/KV7p2fhyj0Kf7qRuhEU9p84U3L7ly89
+D7s5T/ZaoSRWtodLNJDV+cmtnxseBYDI4UVNBBMNpzt429gx4336D/aAFxDWZcx
So0bXHxLRyax12wvo8ar5LOaBTYbGMPVXnBvvLOxG+uJqJ8O7pIP6cBh0Nxmdv0d
sBv+cPb4PC1do9VkjXd0Y7/hEegsSi6gEfQ42zwDNrlLi1yyqXVUzQ3AXI416Zrd
OkiRvbEfFbkY8tANRYdYpQiLLlj9nktICb/ddaFCRUDYWmCCEIRfBBpJ+21Ufq+m
fjaYRHoCb4kFD9+o220ABFyNbaLwBBv3pJsIhEe89+rtn2ubYuw+QnKd6ori/zsY
HKLv0FFQd+Y2wTB8aqCrOnM4YO6AYALAQQ+ayTA0xSAo7iOvXcIbEN1dONvD+o4q
C0Z+5/T3/FZOWhpKGNeNE+YFR3xS70bEGKnPWW/dDD65VpwJuPQnOYX3j91oAaXw
CqkniefJbWoc/MqjXKo6kI/74Rw7fcY2ulgODdBRdE9blk5uKGyRuUPa3Tgo2IGo
2dJz0dTLO7hwsqU5Su5wFJFGsRwbUw1d+c6jZigwo/qm+lIFm8V5wPwM5JZ2+f7n
99OIZEJuel2B5CXOvl3rtZ+SiCBg9WzRP/phXBm42+PzpTxp+2g/psY975R1dhFv
OvRsUsCEFwkVnFUFhH6y9fFqc2ULICxBOUPHKkPMMMCZRc6mx8WcKUIEQW5Wp3Jz
gXGgu3zha732CjkrDwkW0b90x4gvQy4+NqeZ74ovbHGRJkVfCdie9ZkoFyH6REVs
6MGzTPthgT3uT5g05oXGM/h46AQ+3GAjNOfO7WaLLrZt9ws0GXoTyWN59mBFcdZR
uNZfEJZ0zUhNiBK3IoT0hm39HS0YbIVLO6qc/yR/9ZOdk5UspwFj4+smnRXBenQV
zQXITXLG5isSWoyr9fd/nhy9Y2j1vD1CTkd4E5wB9VYkyCYPpFAH2hGgOubhsbd0
RCPRgQdvCFcTsII4ehuR2QM/DaQ1GANPCtvLy++8j/71+VQ0+upd8tPyWwguEUR1
SweF0TEayKMsP6ATEF3i0FkGQAsCjUL7flOAlyIDTsH1RNwUV/AmQLB8VbEyb8wG
NTcvVJwWKPNFZIebjdELb6bdYcBp4c600rld00i4ySyWLlf/yPswzUKnCD78+gdq
kjuhYMwA6xYvD/NyU6jtut66oAmnkgb+4JITAB9TcqhqREexKo1HKjX79P/Va7+d
U+eej0Gd8ZaGEYDeKyO9hjuJBrNXH/A9DElr+7yadjGfNDS3GHAvj+ctRkc9PkDQ
/u1Mf3b8bhN3NHkaDJwF5VJJzZt+IPBS6ewzQEm7M/ShEYs44AZdKMKkH/XnD2hT
kmSoIPHji7o0f3HsFrXJV/TvESixwKzAo6yz/+P+j5PufEyEJb/R0ABwYHspCnhl
Q5bsUiYAhNmsEkVFNE1X6RStKZkMuUyvjno51pDTA9f8YF0JZgM+5+K0zOY4OvOL
05svLNTVUei79T6AkDO74CyFt1BgIkY926ks6gl+YLy9RNI9sqo+aKcclMIbauyo
hkzLBuYckH2khtJj3252pE8Nj6scUEiL7W7Iy9xBpibZ8iuOHykaCKM/w1LDmbRh
4HHfjtmfmMpvwlXDF6UOAugzLr0svHz4B4QO+tCT0x2GzMrda7GH2P363nUYuhdC
tLaMBM8mJrxeBMdW44Y1dsjcQzzK5f3WFcIcgCT+tzXmAEb4hyU960GU+FVii6y8
aaqVqNii1yhiC9MISZ5Oi8l4szBK/C9sSWmR8Nx/bA/i9zlOIAIVZpLC5uNLmUCo
kzpK7qiUKQIRP4auJ+8DRl8dZRk9HYbJUjj2SYBHHOswByvmXZtMx6t6aWt9UVmP
FCt/BWWgi/pfsU9DZbxf/61GrnsskVbDkl0z+vcdqUI4n/J8jHQEXCftyz6DXOD/
GlqaFwcSmx7xupsrkx1M//Acdf8PCU/GPW7TqZ4GGwF4NlIGA2Myt8Qvwv0k98a6
u5Suxhi3ivSmINHYor7snqVohk20oE2XoRXZqAMGkrdErtCSniDI+JFSsA3qWa1N
C1gT2QXKNMwONjKSKK8cO1O/Kpq62sUZfFzPLFohgTvAM2Q74sa3osYjnIgDe1Mh
In1IegMo49m55vrNfJCkH4BZhQTJlh0iKxsCoxotu4hXBEiS3fg2QdTuAKAmXJpp
R5pQefU24ilh+hj93CX5pONFDB+HRrpCvgQ9upAVNaceKTyTEEF598ztLucXr48K
R0eHctLyrhLZFTPLc66GoZ5V1EAZz5dE8/vxIGA5U8kC06Yy8V4B7CmsOhJsbaHD
yXgLWfB8FKfd4V8iWvpXbeVRJNFW/I1Jg5mHtQDo4w38462qZ3QXjZK3Bh1oJ0j6
SrJT+IfiJxVn/DnJIcd9y2HjAj3kIKTpOK91XegjFJF9cMuT0XRmrP+VC6QqT/If
X0sYNmfq0Sd9HpdKQc2SYyiK/G4IOmHzyAGR6c1qPL+ejF4ifdcDI+KA8nXilrC0
68ePsFX6sS6IcgwCy7bT+M8+ACcPMOsf/xFFWau5d0tMR2xIht6faX81PzNAmlIW
2Tfm0FTNNM/WCXnI4WQOBahys4BwveWqFp7F9X/XeLlypMFiYOzqNVVddpuzabx9
Ys4T0meftT89QHQcJtSD83MQVGGnnR7HmYgmiCexciQgocgYdkhNsVPV9mEGIOZI
knrM5QLGotphsF0rhX0yN/qf26rVTfPQfMUeETqt+quo/ee6FZ8YGC3Cdp/QeSV0
fIhut9Lx/lKEpAv89KiqOMEWHtuERxEcI/oyoaL4G6Y5VUswomDE1fQsm4kuUBZ3
fNu4/f2TKf/iF88WJQaBvp9Sp5Sg+hoyWgpmbuFaP/crcF/GIjPWY2DjKo0oH483
KfUDfi6HUCRkUmmbgKGRVxMJeU6VtpmKM8DdXfK8HYap/yaIOS4wAFJnrrkGsJjl
TZsLk1A2xxRA21HmmcOGDfFaBXUnPl5+u4vEtaBLMJwx1nSBCO5EzLmcqsSXdvb1
EDEn4nA2++FBMdiUpwn7y0OeWzp/Y1lJuFGGSdXpZTxlEGu/EiRPxZtoNhqtxNfD
FWdMXQLdywcKsigMkVvXLlWlPSivKSyOV728Eqoa67DTV0lffm6NwX589oN6b0FQ
ZcyJwnECktPyKB5p/qKPxnzN6N99Lf5aS9ndHiwesPPcmzF+/hxKpRHm+EzqpNC8
/EzzgCqkrpEJwBqnVnBtUvbMQdyDHZaUMVDBPOGEw5SHcREVb9EBbQ1+sVndsIPk
71XvFCtTadCJ/KemEy56bgLo7DYlZZxKm1gnlY5j1l8HQQz9oH8sL0ZrW1kWXMCT
kHFTU+1j11FQ2BrgA6izg9tTgN4Dr52+LsdI6SWvw2t7XL8F8koyLaYG4v5Svv4c
dpi+YtVH+06Xo/0T+kHUGVJ21wQ9APsgB8J9+OFsPSxXI2EMvLCqLB0KgaTK4QfE
jgUXiCsDZD9O1dilAx2loeeGQBShk/7099Ul41N62TBJnNlayGjLkj9UDRlEN7G0
vYJfBs2S+czM/6MF/VRJ+sG1V/Qila3hpJeJpI2ncw9ww7dzxLk8jE0zYDH688fd
rAowYb1PDvcbsV6jZlBuFxWkKGsyI31TM9TpKgmEVsN5zJlz0zb44Hg/Z0ElV8GH
IUvMildIsGgPUkxQnUpoSd0LbZ36CqfiIQ6BB/d3S2akfisJJ0cAVJslkj3hfOe7
wi+asuN5PdJ8EhLIuUFMPxKRFEEuh0N0f9bBUzuNTSaPWQB1TGTqlbJwDdnszWa5
GS3RJeVGOJ/iFO1J/DBgLc8PczhG/7UuYFEXe2XD/P8xTlNfDox5qfsS9/730Bb0
MQyDyBbSdQpydyCs7u61K5+jy3po5h9GHpk/DDka82xUMynBDvW+PGgwNgbhYgbV
dEYwkM8QVd7KwWR65aMBmRsZqVtvGZPYA5YdJ23jikkLmxLDxBxrWLlc10KMgd0A
WCoH1ScRKcpPMblXRvegQMCJzuDtVNcgi1W+iAIu4whEfeWCrDCesLeqChQ8bGa9
Fp3b6180KIbpfg3QBfTQjZMum2SPgdAr2T1pxIbE4Wp8oSoWA2GK2yJ2XlPyza0+
WUyoP6SLvwxq5a3hGEuWTAjNdDxjkk6mQoGGWNAizP6cUcQq9HhrXdjsiLAm2YP2
nmrhmfHhvKPMTN4hvM2IqrQyArUpL2Pb+SOzUl4kKxhJ0m9X1W5YSDq0Co74yrDw
hnc6pqMzn7AcMIlJdRhpgSJyH59Et/M8pEwviF7fkAC7XgMldmqBX/l153vG9mvj
YlX05fVFeKQB1duq7xYFj42dspVE6o3W/G4RAlQv1FXZXnvmIoMnNbQFYFD0j6rL
qZCAjwLRKLBl0HzvniKXeQDHN0eDS6XVvu8dyDNNEUS6sXm4jB3vbdLZb3vTNlUm
cU89cvS4wSk3vLteOk8t1jxIK2xWVlT1vR3n1gqx1tNc1OLmGUWhpGS06ZoXO+IO
I9R5r0/wdpC1XzEBXcrUe0gbM1Y4kx0KQ5i5nEPhGzYYj2+1M3eodG8LYwaoTN5j
lqpOphBSlesnMz1rN04LE4L3xJLdIyhwNYKVf/ucuQXOJ0A4Ams7XXnqAMLSrm7W
0ebAYkS6723dX9XI8Oo7F0Dy+jnh9b4I2khNmzBnJNtDLFXvrIji3WSHayr06tzC
+pVXJ47yIJbGdP6KGsVZgxPrmocpOjFvVfSbuU8y4vFo9qaMx0Agc3B415Z2vsiS
ZbwYf+WNz13KluGd5gcU4Cjr8WIaiAsCbbtCvWhRedioC97SqLP/opTlbrRBSfjh
etDa8TVtpWhCRFMRr7hY7DFHP7YUrZ0W6LA34qyk1hx9Nn8z8MpX9bGrx7xmJz9e
+YjiyA6GSS+9J0imCpgeG6l1ECW97jpwBr/eQcv0kr3AKa+K12naY/aKFuOXHVDh
rMnBInqQ5UH1nEmqztJ4Sbhg7+c5a2UP4naa1oe2uD2H7gP9fWyqHKVY3D4mYt7k
ag3a948ls1SwTHgCngL6jDHdu1YJbQNRIFpYnJqrCwYy5QdmocRfSL9iNnXMoaKR
2IVtbYHaPK7U8DW7fIGrDjzrkwGvAmlS78vFqYYJK8FIp9haJ+5qlCZB6ab5amNo
mUo0V2UCFIwXc+Tpr1WKySTIF6Hkd15LBH1kv4SVnOQObpvSRV2du8umcrQlNdCf
T8Oy7RZTfBZGLT8T4HobnYMhyblTv5avwZhTh3r3YtsRajXofxmC9wn2mS+HtCRd
App0rN6M0Askx4noKzlTJNcK3WbiSAIDeK0vDf+3pDCdMgawDjbZql5T7Hf6raui
C3UPU6YKLCAuu38FZ3fY402loTgrJPeTA4LZavyamL8KqO4ixWV7+dNqfPha8YUQ
kND4QqhMAnnfqGlPEqdm8kun3EqZFKZqOLRo95Zrn/TfPMMOP+S8n5KP9uCQjOqI
bkKEZNsJKZe9ZNLED9nkOf62U1+hG2ZpHP3WO7uyqCu8z5sID9YeKctPGl6B5NcL
twJfxmC+A+sjeB8285fE/8tldbxLyeQc0xIptam5+KDp8SZn4m6jEnGgV3o/1dsZ
g+W7eWWKSEg9Avmyijj6YQ6nZ0Ynex0IpVd7pMAvHvELhI9IpUb1JqFs6S0u+WTM
OgbZKAE6ZFbC6FGsTHexuqM+CP8T4n/QNiXJEVXTwq+y9hlVR2CQBGomwpTXRva5
Jogtnj4Yf4trqi33Z4OaEcyW7+zNJTn/JsZcIbarEQcMf/XiEiryZIA6xx1yId3P
dPueJlyhsQJR0eO8B4xMSbxcwh0oK4yHemBYJZUnq0Ri1YUpu2EgmGeSl3u2/qTA
qp4GDxgUy1kW1s54RNFhJUGL0Y9egQUH4zx88EbYfRX0BRwJTRVVRypKU5AUv+AK
fpinYKrhYFtKl/dm2ydn8qe8IEZCuOb4WKXq4lX2Gc+bA0ALBM6i9jq1qOPowzuY
v0c9lTv9fDWXymhfzLH2q34hNGc6i09gwVN9kFr6b/wY9R4xW8i9liLEAPA3hYQ1
w77jXknDIHEbgc1jpQjVk+t3ThRXcVmBdVplHISeRO9nQZFA+eGDxg0RDr+c8BgU
sgJUI25PWdBBwgTHPvavwop95a7qxd0EzPr/FUHqZnjDO7tnOsBNCT2R04yXoFyM
M76njLJeRzq0anuzj6VRqqmd+FWbKjAO/7udmOf00oOM2phU+qT9ywvfsCKCnHaN
5IJCjOmjWJHR3OOQEoJYRVZHjqiU/ow8euhh4s/5jU4jg+FVf+Kw0Q7P16Gu4npd
M5SuzNE/GQoE5PDL/HJQDvXyJIXza14ps+sQ/PupjuzkzeXPEIotj1NoezzjGBKr
yCNNf/phyGZ6TCe6gVwg3fZXcMWKIaguU0Ccuh4QjiBnqvPrK0d+X58jibgceTUJ
cF/WbuLBmUpQPTN19zWY+upgpXbQUc3A1zzrezgf1j4Mxhb8y65oYZ1QCNtox2bf
11sPzqo1oGRJQVVsFDlfuXS7iqd+sNeaWnPcjHsWP1HVIll8y+oF8zM+U0ZSg/jz
KBbw3rcijSGjjSSF2u8a8BsYlo8sgwtNPBIGrdrVAUVcVvK5yVJm40HLiw+hUEFl
wqEyXINNN8GxCiR+ldReJot1GfbEBRI8kvjPQcHjqBNa+fwMhLg6eRvzH09kdEtn
D3Q4vlhCTcY2JsCUsDSewMJ5wWHoKmV1U1OMPyGM4gOLofY7xiBWOOhPSeP7INSj
BFadhSiSbXAt3jgGh4pLnvCqWyBTb6opWJdMiBHkC234MWB1HZO0K4gyJtL7PyW0
gAwjoBwDjw4Cdh3jaXtJeBPIxvnWb6nucJKdDb861qI3BJl188XZ3NmqL37f0Qn5
uWAV2qyMLzcGXdniUehOuGgEHHzXeJE1Q3P7w0gb/QAxrLUKWNa+7G/a0I0+vpWZ
XPcqyfLqL7xek1y+vr9aPDxx6NRhGPI6UNM7O1/FvfXHDT6u6/o7VdCpgtkj3BXu
W/c+HW/6H4X9suAntFj3dO/MiVaXdt2g6OlVuFoMF0w+B+oMOVYkxj9phUGbMD/X
EJXkEO1+S1BYRCxOGgoTYMtt8LP1pLqseFyHquT7WKmwvzno7g+2uWhmSQJ0fD2B
1ePfJjLuzPlFCdhkI6gHa8BF59EEX6/8jaaNURQJJGvmhZ24kO6yCuYAlhU9Mk6n
l66JAkchW99ARbKEAoPRTWnroc73EpgPUFdyyHTlN1vCnqfmO8xyM81Pp48LhmRl
mrFU49os490X4vxmHXYoI0R6KvTD/MwMmOwA8iZo4PwzooRj0YH/VMCVWNJOZZZp
LWeejBBMQP/UV4zTe9HgjWrPW+kWsSMql84g7TwFEj1WnNCnECZY/979Dyz552YW
M/bgO34GFb8e+v3nny8QMvs88YgHru2gS/ZP8JbFL+lwSjWZxH9X/x9aVt7spG91
sRWD5jZFlzDYQiaxhK3tgJkTG15JKGQEBqPTdWQCCLHSJ2XMm7ME8zQkpEg8W950
e/vjzyzh7YptHnflvpZCCqe9IlNKO0Cjk292mLUDDv18NUsI9Auu9yOkU33d3Wxa
c5GivPBQp7RzcnCMcFJ4EwlLqciTRg6wRDm0HnEg7vpstrbr2kcLSFCjbzmmLVHs
Fb1jSMyHRZDccZo3K60NLU5kVU1+RbgPRg9c/qRSSlz285AnTxsE/UYUUBFMQoa9
cpiI+9ie2mhX0RVcv8drZ41LFNByv/9MDZa0qi6vew8q8IDMVY/MB42R28kt+Mrp
VDMh0nGE9couXC3tFJBWCKNKqXvdK7xt44GnWbCiG3i1fQj/FLVjOqjlTneZoiM5
GJwXaNWT0Xr+5N3Q0+xAPKPyeLQY4tGK4PaYEt4nOPkyrPdNoXhKDFua9cSSX4CM
5yOuWe4/BqWdy39IkiMh58SVWzZYmHWL49JDjWlKipJj8ojwqD2WS4enJjRGd0eW
9zb7hPSgJaeY0VqGeE3jda/IImiSQ/wUKdsAEBiR8QagLiRVyTlxbhAO375Ir52F
PtKmRMNih1Fpu5LbeSUmGzrJg2HF2aR8oKn42YZ6S+Aeqy49XQFAjVhJ9KszJdZQ
TCFdZwkR9TTR9IygXRay/j+4M6e0USsiz4OSVamRMmIuvhvmtDREZro7kUQ3WMSK
WZ5pqxwhtBy+O0JTLin1AVWPGaH4zrAkGr7rjRlh/ZWJ0V2QWHXz47VSm7WsIHje
nlHix9Cq0TYrKiSxbyVjTHwST5vqE99Fy+tcnsSuZ7vb1ZZHXjoiE2skHCjMinx3
ycYWEBGdcO7QU8PrmcRr72zYPbY8yftY4MabI5mPLoBfxSY1nRtJqUtsPHM0jeX9
Fx4u7cAJbDlgZnvtG586L3eKPc8HTKIUlUDxXpb82WrHnAe3Ls2gKrW7xyHpKzWJ
lhcub4B7ORcc4ysfQT7Yo6GjV/x7Lm4ZIw0wofgn8IYlxrrZiAJ3WiAaSpMgM4yP
oD0QEvPrDX/vJqRDlzBuOUu1CbGuphddEo3dOgmwOErR3M24b7uItJ6KTI5v7jCs
L2a9kzWcD54x+vnS+w8/67jZ/0nkbhdpqYxzthmX3K764SkxoclH9vlHtPdXEMfc
Z7Ra4j682WyLGaK75RYSJ4mgk/2b4ige7LrOnHWGmTQDc8XfTJLjv6sRAAvHOpDV
BMIYpm0Nxt/ovk65zC+et8jrKm2PfZbh25+EzWcJNIHhsexbn35/wr66T8NULB3r
IHQUL/k36tfpbcu2d2wFiQ2i7RR9vRybgpJCei1uUsGqKmrOnEwqhnrrnL4jPYr4
yT3qUnp5ysXgZVDe02fz2PW2/0tEKUH3AlEYY1MjNOWdkPhq7H1kbMYrtI8jwfqi
VNF0Rxi+7j6J0yClymxsEtfs81HJ1k7IvyTAkFMW1enfmL+lyVHRMYpu/f003A/t
RHDXNCj+qj1z5j+9+K14LDMfrDKyzAtVbdgDcsXR+72eAnCz2E9dHpdLezM4OWPd
2jvBfYlYt/i5qbBHBwEGZN0yp6Ep4YgPunO3LLOgeIEeo5ZZHXt+7J3Lo6flsEXT
lcEjFc7FVVHr9ClnRKYFZktGvEV79fZI/p8bycgBckNNZcl9Gp9acJW9n3aJJvZF
s9EQ1E82KEzitekiMP7iCzBMThnURCXlsOPsnyGjQVDB1gl1hgOtwHynN+KBXdS6
Dn1pPIx7RkO+e0o4w+vgINqYevnFJivsGoH+uUsLpb3hDkD1rebZ588FOTU40ucF
1Jwutu56knFz/Us3vsoT1n/VjHZgJvDAWvp0W+JecRaWz3hqQ/OQ53Rk5KnmYpOv
qqypYTHe7NFxvHGCh+lmMJaCGe/5ECtXGzm58iXhOVlC86NFE2cocu78f1X5jl7A
dKPQbz4EO1xAPj9WqO6SV3iShQHDz5tfEM7klHMKYN9A4qXjLKyxc44p2cZ9E62I
jVdrCaEeCNK5PZIddkFdf6SOA0twN803g4bjF2jhP0e62FEFVJ8/ZYWHbF0IkQrS
VOlweuuYiCN3h3FCbKlTrCow1wDc+kXQraElKK2ibI5xkukIyzxIN4vzjBZhnT+9
8JBMJk99HpnvfFWzzgQUe+m0vOaSVF/ByAByIgmSZbEMs4LBpH6GjMTrxd6ArELx
UrZJUbHd70MhHMOfWa5wH5xqrd9Cxtz9N04MdflOgA+B2OuQckWL/m2o3V2N3qM3
ZlaMM/HQar319oMZzfAKcd2n9SwX+tmJkVAYNdWrG174C7M/brX1NetjuIVI/T4h
OuUqpQPt9v9oS6dYVaNcoYUhCbND7dD9EJyNtA2KYE9zYeLuEKryYZQAq+QeoBVX
QG14WuTasxtUPR2ebd8SUmDHgzGXsqVhIFMIE61i964HzeC7LJhLQ0sdCIb0h1js
xm9qrN+DTnwQxhjfqlol9iZSP+5M+AccWQOX0H31u7/QpT69Op7CpsQxeYbGbsI0
lpIvVcQWYoyiIkoPcDrqQUHbJmpk7sEtzQBdQCGNW73RnhSP6Z0zz2RHVDDFPd4k
zsAXKLk1p7oI+c7umQ7rEpgHy1DHSGCO/sbKiIC5lRH+meQbeFoTjC3IphXYuCHX
2n7U/F4R1DEEAZyN24BpdCXBO/I2r//mhJJyY1/M/PjYwJfFQlo3nk769fakZSaE
OZKbR3nRpuQzEDZ1LjJXzgASy3zrrtC4rAsRJKnReNqjzrjtzwM7gFzlfHpFp36S
Of2lz0e5U56aP7+tHx21qfKjffAC4hiiVGgsaXQxPYTx/Ijbdz6ZGDme7fiQiLZA
iEDPdbmd4nw0qdogRUuZhe63isH4GIb4DCzkYgnHEIgejnCeD9g7Gm8YWKWxEH9L
a9AhGuEVeYoyen+58Eh3g5knwQ80g85+5kFXj+ByFy9u3KXbpVawKu8/JI+ezf2P
iYzG17fvsrcG9m+31F5a1oMbOHcJlKwL0FvO+MS5l1WP6iFl58y4nWUG4bPFpcZG
WK3oQXMFdzenLFRLhFSSo50DkJ1TCQUrGCuAJTsBYvVsfyrbwhqC/QcGyZsYcW2k
8X7jjMyaLOXVdeh7OqfNQ72VtHMD3l/u+jqLFnp4tjw5w/QiwqglR3d+O5JxH346
dCWrwkQ8CcDp1NFyYxtBQSRzScKCprEqDyDfqKMD5B/pE8OF9enYFrB4sOhcv3Je
UK2fWStfpQPWVfHyAXiieE7zyuW95Gaw1jPd2bOhVEgtiUFtmnEv7+rKd9ELneHn
JrKvUv4SMp/q4EBnckWJep8UP+HEdQuakEL4wSMO7Mo+sBlOqOAwPee57Vvfj5Mj
NEOHIeYJVJ8fd9SC0hZ8ahE+PC6K2sBcT33eZne7GKv4WGSAWmt5qZvm8VDd1EKL
ZAg5GbErZ2UlMw+0gdz9dmXCYxb9defaqZVNtKjoix446UcYJGTl3ssNvtEtaafI
T97yVUabAj6Ns8aTQcj4zhTyhYGEH5BDddXWRr+l/5wsIkyJslLb0BRo4eCbzWYX
Vrga53WiF0KZ+vHTCw3vfdGotkA3W9VNiOUkiDUgLxbOmIOc1/Q9LCNQyfVBfymm
mT0Ktfjp1bRRTdNnGC84C5Z2hfoECoo/3ohNYf8UYNqZTkeXxwqhn5mYmbVYiMOl
WFit9K6DY9KQdVNUBuqaPByhazed4oJuqwmKkZNtbTYht/dbmjLKF6dB6lqSpcOe
JH8CptBYt+HXcO5VWFhnH8Y2P++0jMYIG3DpcihRh4NkWgoeE08t++V+jgAgmJR5
n7Ly1vi8a8C2jk4qH7h61wGIS7kgZ3tQeOYtsUEbgbA2mx/JWDWd3ZoT/yO1NDUp
T110SkOasAJlpcsf3quEErWBq3e7EY408UqMlRXzYowJn7VzYNNhID7tki30BM1H
K7Ypq65QgrpN1CYbWHl7AsKEBOiI9YyFiJyWaCuKdg1hjui3q+fSV+uBK3FR/H/G
VAnCVA1VGJF+nrB/gvki6bUHUnDCZGMoz+copY5u/IfFJ9otnlml4jeXoCYIbp3v
aQ8/mSj9z5QkraMC0ygDskc2o3JSdLa6r8EYovhs0u05KPVlb4axWb6JeXzlJjE1
Ry/I1duUNuYTm5IhiGjGjBRl3oex+DzOXeTSs05Wdj0+lAAaIlG17022KGdw427i
k5W/A4ALc23PblMdwCjROv60briazjVjC9B+8yBb2M/NWKgK0k6u4HJDEik6AwXB
jHL6FRuy2WZD9CStmUD3X63dCHEpFCtf0+zBcJN5egtkmdG08/oHtp6Gm/3AdiLR
5x0EyLLf+cc5KCiK6WKsNUsnmSzkJMT3HcapL+2VbQ/xS/B87ABqtqNQOm1XpNDZ
TSeeDpJB6Rjn5WJJR99zVEwNKyjhfzYICaXJsRFZt9dK/w90AB/resCWn8/sTdW6
oOWiB2+M1Iz2pnl3Lre7e+DRe1XTn6Ysydb9thaCi0UQn7z1QskEcxJ2TfYr6dus
fUXq2CW8AzTYcqheMDjy9zTg+KFjlOabarzfnFFqcHoL75kYG14AhH7CJI9rCbOC
+vO/6cFPYAc+CRMjtoNp28UAd06Pr/ouFvZ5iX7dFzLBLpPk4ZjhZqYetHqijdOX
K42ucIOvhnb6YPgnynNOymCKAYlPe2GKBWoKwYS7jPvgpd0ICzHBWyqKgVLqL4Cj
sk7hdIESH9TVkTtevnvBFhuZBEMAk791yT3ilrlV0osQL18Gq7gZ+qgJvpqHBgFK
K53QimlGP2ASQXeP7G2UTCnxc6Q1z6YrLgOm+qvEfWCcWxY1uQfA3G+XrsifaLoB
28WryujSShNHw4Wfiv2Iuf9waWn3c7WBJ3/0mVgjetLGAuoaXuG9s1fkG1rNgsii
N65fFe2wPv4rJvlqk5seuopEBsrIMmSDzOzRhqSl2UKpr6X0L+lePSEalLePa8ab
kYeiPgn+M4nT1t/ORle8SS1V7BKIxqTs8EKVdRfRT65lzd3fpmjCsFXPbGA22j5F
6qn+lYeNugDglcf+mOV/AhXbjkJJ0RmBZAU/5/qsdoDfSak8uRqm+JDVCgUupE/B
GSdEXLloWBoPka7sdWt+mgFIcmkSYFJjQfLEviFKfDR84NacQd9I0ljzIVE6almt
AuuZHVSkB1ktfw2ItmgVKlQT7AMZ1nTp9MOJYIjRJv25BMGlqshi+O+pypdlgYKb
NDYh4VHxMKuEoF14C5wlpfgDQD/gqI5/ZMuHtlwglvPmape9hQYky0ygiYkitu5G
aaxqQSPzzSH1j+1OlwtoFsSi3pFYYLL2m5imx12S6VPaLTLoBQuyT2aRWvnjvL6e
zodPDh7soJbpGeHQXbllZ2KqPohM2X+xSm7R2ZDvJPSte7K5l0vG/uwl66PC6FXQ
2vD91/7J4leNyy3ttZaHBFN06SsNFYW10d94ZW8HM/Yehw93FMetRCPVI3trhfEm
CDLOuttc+XNuyTyDWjbPI2Ud9snRZmgGZjr29neEq0tpD1z45XBQSa0eS1GfFGHa
xtZn32DfNpQyyBpqkYnGrS4N7t4lAynVPTZ1ZvUllI8OwgZ5Rrrk00RSHaYAgbWR
Citq8gNXMrRiJUhnLbWI7WZeFI0wI7YHVvu8cD4rrryv4FrQNnWw/17od01z7Q5p
PPNvQWNIPFthD6Z0riJImPOvouXRl2AqZoXW3cVdQYHGJxbcpHKfm2j13a9sHxpF
XStw1o80BkMxykzn4fbIEKAPx8xHVrxss+/LNItfb6Nu4VMID4Dyb5YD/G5rLaaN
q6Q/5yFrKO3OJ4WKN2EuXP4SRxUYENf0juqomUoFGkBp1EZRdUfOVUmFr8iihIfW
PTVxZ5DmAU5xqJjL+kRP0K54ajeOx1ejO4si1xZE47X0ojqtVYfXkJ2VkEmfyaRI
PqLYUiAIlvtG55OtjdiUado4xEI+XUIzb0BH7p6WT0AmaRjXuZ9Sts0ifhuVvAJB
P8/quIS+AeCUtgf8LDSJxjSaAcap3I5CrCZM76u3MvCRU3MNNsD2dytI6j7/IPav
TOxu54tEykV7jlXSETzWgUXm+zzIvXiEOX4vd76A5OcrrC0RPCPjPxf505W2QXKg
dLGBqhPR3X0Fl+wdg1y0WuYnJAao04wxUyWlLw0NLKX3XAI3VOVZX0MfXLs+CM2r
dpBCCypIAW/EaLTQAuqp94lP+CtJ1CKVVx1nImhv1yRQXV62klK/7HA7grpozQ1W
y7WB4yZJkpRXnwd/OEwS3LEu6xwqCkctnLYWbo0CD+CmwaFBZL0FcwCU8D9zZl+Q
DdeQ9P8VzIBnmve+lYTj+noGc9yTY87ODGrDNuW7DxH25ffYY8LO/St7NhTE6CoO
DbVcq54EW3WJ73zTFaNdSOMvq31bqj3WRuuGu3Et8drC1bfDjY1VOgzRXOlPVBHU
GiCR4ANSu2l8x1m6QAJaIMKpN5kztLhT5M7z4wvoGUueUke8c1OKlsxwJEI+MbMw
57oCKMdsxRQUe2iteDD9wo6ECWhQmhZ/hcJqIgD2/lm0qGEIaxWjjYWwOu+rF6nn
wr07GBIKawTa/1MhwPvSgByuhD7qcWawsf5A74xPX/cM0FQ2eOKemjnP4vRIxloJ
9T/GCpmho3vqzDODeCEXYIX+37OLSl6xSmN5o4wqaB1tzi+RQEpnB8vG8/zpDy7q
2zgm5OMI9IG9r0vb4skrG4JGGozLV//2TRrEqTQ7CYhlJUpFMktNUeL36+BfI86q
Ivh3ZFpyfDTME/8s89mg5ZElgwlLauOuNFCqlSXUNOD6nMI6hlN08PJcell6q0dP
XkBPXr8Ih/RoXxB2tbogmE3aQmsIdUy2x8ml14kBkx6VraZhviuwUgCmvmz0n3PB
pxP0C6QQBFnFRdOTGFLCqLq+6as7tfCcnOCUazDCA2DtJxwQOnnC5OGIpcRvVhc7
VYJ6roIagryiPHD+Cgz3bJeCSle/OhP2FFcTuX+RpSVcI7lwPtjOrSwQeUOq2wd5
tW+MhgsTfmUtKAWveSIxnkVYl0COOJJ/4KariyMYPL+pVqL5fA6j7gLnrB5SbXcv
Mq1Fe8kgdhLl8g3ZL043fbFb3qygwSr2vawkN5mcEa4vkZzPa6rYlPdc5rc2Y/Zc
W8JBsl8Zq+AbP6yNg2EBuJ9SN87ATSMa5P/1OYa4de7TrlwXoqxZZHXqu5jawRAV
SCqN4c7AHMzkTk5xuFwmy4S7ygVKxO4mZF2dhnLCcze0Vj2vzwEfsFe0f2ubLEig
h93LiYmrFNFm93gnSMZzOyBjwj+HpA9drRjb24CoRURHj1nhGO8CWuACMo9bQJjI
jtCVk3/SRE4yjtCVEPIUNJB7IVnWZOUZI07k18oNRqBFEHO3ai0+jaGCNaS3hGbP
GVDQn8DL+W7Fuk/aUFwW5c+zZkmU98L1c8ruq9h0xNVnlxS98l3WfamqlXQUE8o0
JJ8cJdrZvogugl3PURL/IuK/i+7+vGOCZXVk/wVsEsBHO8X7MYNhtG8Y2CHBKtiX
Ypj9mHNqxqDCm1Cp5qwHtGRu2YPjqKoOQYL2CNXdgTVfLpdoGqkjGcPUD2fVNMjw
NeUvSIOS/pug9LoKrLZd1aqD1eUKR0EnwyZGIoabFyTX11751g0t0LyF4Itd2Zu4
jNICnX2Pjtd5DctLu9Eot7nZPPBX8hzmNyN1rppo938CIyIuJ5ePGuhLuetgQApO
BGivk1bq+gPfpVO6vue0UsOVbuu2YRbqQ8ge1NGoioiqVrbcqNcBGM3JEhdijd2v
uoM9eAPiUjYjzcLo0VFpLV4orwGzFyVRr0S8Y0QODll5edGPNyxyMYbPnEZcjblM
0CdAqj6W6jduDXbfAbG34iYxcngIvLgC5X39UV+puQR6qBHVm/a3zjy45MAvq9sd
XnIYj3VkcvLNAdojm19mJi9HcoRB1N6cBmH0i8D3kxQN21Y6byCj7zWmynkfQp87
GWqEyALxz4uPTZLWN0XVwXUnZPCrehY9PpilCvBvtMO018cbuSgWILEzeSumDbnw
8zvOGFENSG0UA/Ea3lHobzh7iG2THE+5NrgVVUgUKIQB0i0yODAKN5cOKBXncpqk
TYzMRMDANwXxzm6pzNyTSJIeSbEE09PBuuCLMK5P5x6X/ejK82/RR9LQf+WtoJtW
RbxkOQ56M1qJiGST6FAQ8v8YU2PVcozNhsBNJ3TLvOlw5XhNsuBDxwn0xfnAJXGQ
2jYuQslnYwOVRsyYVp0Q8bfl/qhvTPi/JT+TC89yRnHsipfT9pIkAvuEloQc3Gt2
EZ6CjXqkyzu65BGmB8GYHMOYdQM9pDYyrqwjgX5dKFZDyMCYKw5OnVqzBosuOaj7
LCLs5qv3v11VD1FbzswQBj+INXLvSKdWenf2ZoPccdV1116fqGFH8IFbRXs3++wg
R21hwfjJIMt4gHP6htvTxLGkkIZ3Xm94Xwd5yLOWmJMZUMQXD+2Ws2l8SJ/diH96
G+YTuI32D5EGS5cUh/m5sBymH/XRtRdj/botraDiOfeViAm2CPP7/BZ9dCFHysHf
Z7XMH3V4mL/0PD3hMPFpTrw5OdMMIohfZbYbJ8kCzhkhkGGymmP1MflJvsa1xeIt
hOXMvohBwCEM7TeGRivGGTiatEuMc4rGAabbl3BxMQCgLQ++MGErHsO68gLchNtE
eMkt4mpnjnP0o7VWpin2CKcT5XTB2BqTEJsuHmdgLgxauhqkv2bsDIxCDk4oELRV
JWk1KbXgfmOLOtw/HPIm8SAotTs/qzPn57fnuPcn/T4EUSnY0OKSTdiiHu4/5Fle
py64H0n8lnYoKg5J880pHSov3/2cZAUjcD4QSt4PQf70g8x6cK3u1SOBbNUzz20H
e50OzTigMB8Y144r1qbC9ASrpJ6WNLoASiJSdlQIAE5q66bhOTof8qJ2XUWWAecP
SZWZmGm1mzfq6kyXDJ3mlXUgxvitClIlW4ZWSQsIQ0r5Jno+tovYJNRBXbiZZqxX
YyJ5v9SgsTWhR8rWlA4doQ+SaGkRi2WuvUSUszEZtJvk7EYo0LeXCOIUAXCrodHv
/hzKAnUAJxTUrtiJybcOOB5lcvYDmSBvekcDrXnnOLbA3I2HSNkltI8l/6UxgLgM
m2oXpdJHucEPWtUhB0RsSW3oxxNusRBpXc5sm9TCEwJl2udBnykfHxzmc4Kbfy2Z
ZgRmsHKDTRRzBn7N3cjuuDesXHkS6W6lOMOXCuIKA2MbYAIkrFVfRJPJFdnyhFeE
bUVDcNLYQf2Swcwny5SImQ9bfl+FxAPpAkHs14sTV18Xe70xmUeBt4jkKKxMRwDa
z3K4sG3krFiJAxliIL6PMvulwqkEfifx1tLo4Jvp5H5yWCWN+hReetdq1Y6tm6uU
ZZUQ26kKTRWnZyZFaGo6B4zm+kWpEP0/30iyF6JycnFwM1ItYbQS1zv2qTi1jx3H
3PJKjY5cMlHzBLmmGiiaV1Cjc8OPSBHyz5uqembwJXZSJZxc1u7jjt+KsesnFXVg
gOIFtDHshTZjr99l+cROyXjw+EWvmELMSM3nbLNW8lrrsI/kjw/Lj2ZtfVQBe4cs
zmx3bzEv2znnS7rNreYbqPQEPykxY3ylfvvzLVjLHOPH5jORQ4i8nlGcTI0VQf+S
j38uU7zJdw7osUQqyX0fzpIEenqIb8AcG/PjxNIDSpt1+HJZlKmOnp83ihXfjihG
1rSvaUDIgGxYnjsTEakMB3aZKOskCvC9hurRT/UOGpVckL1AsV96oFbeSTeJS5e6
9wv3WHgEoW/WpKzpMRYofhH4MAZNP/9R07U9ytXDfSltJeYElIHMWYSdoHj3YZLW
osRUuz4yVKcq5WBSywuuKRgr9ize6pdWvjXY69vTu0SMjbQIOBoPJMhH/7CS7Uor
T8vz/No6BWO7emA3ClW7fJhpYhPd6aTI2uI6EqcpoSt0ARLb8WQiWq6ojtOHaO5r
ZfON8DzoGQAb4n0jI0XJEvzKWHYMyOAaGon1l05jukH3dwqrdHlcAYFKiHRyu+Wu
2jnmzRXAPMAmWl/KN2kVJtzUyCvOQA7rf4htE2B8KGZh4rjsj/le80woTIpucTB/
r0novT0BTqWX+A9MmpRX995VvEytZhwnu6cmFuDgDszlNNMTWyTietBEfMuFyLZy
FSBqezxUfZUAlu791K+Z3UOhwir1BTSq79sxz8Eo5beZsj2dqyrLEKU8TFAA2po/
W2+Rqt04fhPQ5jDY1Zet+Ti/TYS6ezfaDX0mGLWhDrdabJJSekh0Dw7YUvhdhFcM
IiaCfo4dxyIyQQRJNtD1BLo7H6iwghGInZGUmxr0bvXaFMC4vQjviJHwpxVlgdTo
cW5tvnVYRKxIf05ls3epnkHzy7RnM5fC/w8U7QYRT6zpwbM6tSnWc86QWkSvJmdw
89ExDE0sM9gmhrl40vRFUI/iaeUR6pQ5FLx9OAmk+Wh6igWGpWymEXIAKukkoXP1
aHZ6CT8tBqlHrn3W8DDwkOQa9TEEhqTDvf3EgcKIPCPtBP4jQ3322dBYU+KOqGqZ
cs5xmc3x1/nmsPpOAZgjT3fJYXspZtoY2akOq9rO6uy+uM8JohdshYYF2NdyfLav
UcSCB2SwwuV8xd7CfWI8OSeoRvdQjgayK47oC0s81sgvOo4L7TmE/q8LyBe0lIQm
s+VM80e/rEPu712IjCZcHHux/6JswIwL9VwoTL6xnihRo6t1VwHgzMIRL1dmR1MB
rI97xxpX2ef/xQzmpakDKZZ4fVOarvDjj2J8/h1JQueO/cLIH3d2kkkooNodt7Cr
9l7kVQQ/Ruiv7winUmTTXlxCqvp7EDTcAHXolwHQ6f2zJO3MyMiXG2fbUCAF64jT
wECcMEkXVLVPgsZiHB4cPQNx77ZILJBG3yCVimVEgdUmabMn1gUB3hqPgsMYb113
AztjnYCPKUr0e8Rj+K833aWpsOczv24BJKJRodoSCo8T00e2XaiOmxkkOMHqCpbu
ytfvTPUmkfIX4UwcVOEO7O5LJZMja/DqQwYBElldoK/rIHzz4M8/F178V8bUVu1X
Mm5FGyrFy6W/pWNGhI5nIrzTgtYqdgDkPJNrwoxRYElYuRd0dixYfUDghOB2Uguq
Y9giz0/1ioVwbk1qAs/HGNPqgc7td04jHw9SlZ5w0Ayni9yWqwCa0zDA7C3EwlY9
7uBbA37CodiaQReRFXiIPOLbPvFt++L42GWrZHelUbArFEs0YMz7aaWWmDN3PLEB
rgFFvxvMQTAY2Z4QfXcznDusgOKL+AR3tevTmtJ6Aq0ZiiLRa/JffgdJoQ2BDdTV
tZpMvwW5WY2hSpntFirMPvhj567NLG4c4o9kKRehhjJcxVd9K7UZtpVbhgEN6wvt
vbXv41s3riRVkk2xqTnDo3ckHdSeUGi5saVcTw1n6ysRV/Z3LMu4VEiiYuf8S2hd
1GworbxZjUdbNpNsxp7HPIotj4zVi3Q5ohU92ob9V2wC6f+9VtFO4z+H1iQ7u8PK
TdflV9an62Q2iT4pF+oJoEOJy7dwYGmY9b+YO0BesPhispGLoiCBa1UAJ4hUR9XW
c780ff6krJqSSWiit5OUAPKxL5LZS9bPFJQ3PuoIfM1ZA9r6HBmQzQrxXi2UAPnz
Cpr2wdqdTxKu0DdpJj/vKSBWOCRH8snXblrnyVN4XTXJO1O5xcZHJsjBy4jefAjC
bMnO+L+2oLlA/Oz+1BLw+kHIqn7DUR1au0fKnoGaehibUuqyg6hI+QXh0cE64RMd
zkdRrgd+Fkk+7aECSWRQY+dpDC1eZDBYNtov9/4hUf7Y70zIdNRvpEY02frMdwF6
qqjs2OoyNvx6GoQGLQOGej2GBIc2yJGAGJ/woSL3EABg8NIGzUO+bBuPf+w5gnmb
lWcCCO0L//EJVF4M0EBzlZmnvAj4e+pCsdxcufIWb8+hdKt8qNq4D9JDShaujNrr
UMlS77JauSBRxSzJXbVLqj7dXJ8406Knk2IXEo6WTYWXqTkElfe01Mcb68aYGcre
ZlXGAcejp65jlPdLSt8ldxqXg8AdyoDuO8KZRD1bYNyZYI8+r2PmNplWwXfzZFGa
Yhle9F0wwm5L82ljX8W01sTCAXaEt/fD3/FQuSl0TPH4wdg1KdLDddZ1LTCE3JeB
5dgv1mQyLmOoxpfB5p8h5z5qePqPID8XSEynzWrYEoZQGf29tt4iokMIbL6KlzlY
DlPGPn0wM4yaouCG2/gfDUah7C+6QLmONOoCbfcXQJ9JJXIMhPOvynZEjyAuJyV2
tOA0WKaBJ6RUUN7QZFkY1yO30CGqGAszu3ktvEhTQ1KBxX4fywtoaAgIeE+VmMUf
uHbyjuQjejYjT0y9QNX4u5HjfaEIuPbJl76DEinYJniXUj5fcjLmhTrz5CmBoMwS
D/ORLSVn6mUAb/5s0s2I2Uab4rdzwOONBOGLzKED0AXbUcjzkX15LtWGv600w3J/
PiagflKQtce/EttQZ3Qd9KowE6ppCeZOxw7K/10+vc6KxR7woh4GE56txX8sipmF
NyerII7BIOYxmLkJlqVyepKMzyTuErJ4ZtFpFMPiLsZBB385QA1Z7XzxKShTnx/U
U5VRTaGWx8v0GLkLQgAKJVfTRNqPgXhSWOI66m6PcAuM81oaWcCjvXqSesYCwfsm
6zr8rpOJJg6hZ7dxA8j6m4u43JR0cBst5mHzeankWR5l7PBvlDVZkraurWFwdZLz
8IfyW5tgh/xjwDa51nwFFng2rJRDL/zHLZNW2BLJBJxvrxllCWZUTw8eZrX0/06u
vW3BvJlStuzU9e3SR9f/Fa3pbunntmAaZR3AZy6OuH4wOIrJuATp1kvtXXjVbnBv
BxAsH5jyozMDlB0qCXU3S5qElw/tdg2JmHYeVTLKkNyejxDXXg80fqeOzGwpGJXy
Z/VrFIw1eSDLhzzxRxOUQ0LWm8w6HCY9YxBG0gOWqrrucisxtNSfD270neosOESg
9b33CWU/4OGn7lfra8sJ/Grdf1l41qOmYtW54gPLB+R8RW/4Rf42q33z1ZnXGf/k
iev4Eo0mDsCxyFPt7UdnSgn/wCU/BI9tHmm7ADx7kTmLoyHi1nYUJMztco4cjRb7
WaHRpVBB94tqgsndJpetnF7Iuc5hePwdgG4iwHiltBQpIHP0w/n69TfhcbfyKQpI
gJ0zsnzFvAPh1ZOtjOzCzqt+0gUcw3iuivTzxKQTReczKHzYrnGPhdiAwkM8DTii
DGsUmGaX59HOR6JKkUWJBe6bw/s/pwFsO7awawVCPdTUiMatMubzhEtzBixbWK8K
2zF1n8A3YgNhXyNrs7ISc6Oo6mWfodqB126OYENcodzVNb8/aZx4u+99Dudegm5O
IiJ323QizYGqRF+Pwt2C2yINC+8bqhsfwLE/cAP7K0OTPX+GJwRe7w+U2o4uejRh
e+hDAlAwPqcugG4A0w3DRaGVuL9sVANk71bcVFncT/SnWGjGpN1xTCRXx6Mn2PXR
FeNbnProlIPoFealCTuL6gGapGmRk5lSunWlLwf+cAjFlEAD+NF1VhGWbEha8cnZ
V1DZO+azJt96JAdZa8BaU7uKo/W4p0IyLD4dHbS4NFPka5ZPr0xQpgAbL+7QMbSf
gO94JkdnE+EiprNb/YN9bQ9fl2WYXJiZ+h6F2+ekqvbCripv55Wj7eKFP9oT1dQO
U9FA3RwDWm2MIArKmLqAPLYYHP1qczbZrXfjscot9CkQV+pOVdq2MBLvOM6/oiG7
f+UAVBJwkLMSXbc3adJ/eEAbVsSiiRZmCPhph3+k6/ev2HL0/3kcXIY9BIEvzreI
Xo8pHCOj1LVUQ9U3hUM9/uhn27y+zo/hmB6C+V1luNZIwVa73oO6E3SYooIx3j+A
xPwq6PZZPjdkbcanpNWUWmgazDPDomQ9i/j7ZnnIELdbN2RdvcNhHuz/10nDtf9D
ZPVABY/GeGt8ziYYUfjN/zdcn8osPrDySe5yZxL05du+xDpgfbw0fEhS49fQm+SQ
hnKJQ8e4SK5Ipw57HqbUTR3jJHPV4xNDtWXnJ24HmxIxMxcI55fp0ZA7bjNq07ph
YKzQtA3VhTEnWUjM0jFkkJgVxmecMRF3nglM4KuaTOEH3HVFFri/TSyxfpHZwH97
lpDxzBIODejUvmw6nccXWPplYzC+3PeqPQZRfGpPgLHDp0VlsOPMabrTesFDZHGG
fYpGfSbUkSYuCZBnAkJxvMZkn1Aern6CD2MPeAz3xF3jKcZGn7QM9vUKsegI18/F
F9NhkweleXxaL2x7qY28KpckLA5EkvSQi3K9KDjInMC57D5Fz4Rw7tLDoOeaAVpp
uutQrgGieWOgoJXGgrLfY/PYE3goVOVHsRgobEN+aAik3Nxr57uwqQg5VW5nsmJV
JIUrh/EGsMUvE3c9vgmlPU9LuNM3jyBJ3ILxjdAl+e437wwImdP1kyah2nAE8pyJ
++LvDBlvPoH+0EGSsnJVDWpEqtMwrOiwIsVwjzsJMezuJEEOazulD9JorupjjW6S
tu01M3SqdFWTjf+XhBB9SaJCJIENVxATyM6fVCwMX9jtprIsqpY6xSqI6OoCppfu
f2rbQmEM5OgHor6T3pDjJzGRSikL8sMq7mUsDcapTRxQDD4mGkZ55sf0zq0So+RP
j3b4bKs2PUKnGuwOgWwxbEAw76zYG0kWsb4DvNoYz1HblUSQM4VvYz5N+hEZbWcX
3otRCeMgnlZPADAH72YitUwMqnwFE6x7ZIJCS7Bd7+UwGgAyLYpbNfrUPLxT26cR
3TeDkip57GunmzFNYnMKz4SV1Tm/vsm/wrsmKEzcFbjTb/AMWupYmDz3yt9q9PV4
b2P65Q46FiHhbqgq+phQl89GSlaNFU7gYn4r16zOrp8HmydEZihaBP3nrbmxaKP+
Vg3AJl0+z902d0eXrvJL0t8yt3D5//9RaxiWIyaNBBuCrt58hUCdyHrCbLBR1yAY
bJaM6nw/XFoiHzo1/rWz22WPYGwFn8Aphe5k7RzgQOhK/IAtx1nRQ8e9FoSHwRmX
Xu7YddLngBA2T7vq7+Y5f38ZIHj7awaDE1UBpo1Gr4xiUjBAsdU1lcwyMNwfPVdd
7Z4rE2OLvvZ8Mqh+OtTpk16hySYKxd0z8eueBXxJ74b0X/BZFX4q/WhBlLrMz6Tt
Je0B6fVElPWAXGAsGndY0Lk3yC0wvULYJbYbNyTtadlwiczDHVDfzwXAklSlAvYf
KB7NX2Z3gfKBRW8n1AepELgBIkWRB54bs+NCX7cA++d5Om/JJMYSAdW9b2tI1DvH
Lh7cldBY1p1S3r6U9cHcqMW1xsSOOuIpi2GHjngW5Et9s29lUbR5b2mHS2iqvjTy
wzoXmOBjpwqoYvynbhO9SXRXAEDnRU3zrMPhbYrtR30R7/7CqEuuGfJmysNAMB+V
4fzQ/h30HWrGF2LFjyAJrdBBQWxJ7pqmYPVdmN+33B3gv7xHQQKdnZpdU87fttuS
H+NazBIX43SfUY+LvmwWxIseQdFmFYZL9Ee0zsjZJ9i2t/aAGbijGdld58UlU41m
sz0rP9VEq4ozZhRU5fkztYdQqEwVZY6mcQDBGhr3cnJw0FPsqEGPf9LiASpvfBaQ
NKxoJUACfOuu8to74PdOifjcQq9IU/nuuAKqRci5TRVJr0Ea8M66yylcowazO3dv
Ssyfrlv7BE6Vnyv50WpKecvEFz4d122brTyOdRv8a7r4faUY9ykqsqgck1gTLxsG
KChPzsZWdoL46VCxKKHrsoL8qDfLHV3Ran6sX5thbPGNxcEC317zKb5ho+4tXp3d
qWDOoNAorSUhiTs3MMwcWlk0OJJf6YPz7L/vvxnpUCa1E/aatyzB8Ktbu708qITW
bYb0enimu8J7A9zL3m5whpCLkJxrSUTcflb5LBnROludEePwRQCs3T/pu1ZKrFJQ
vniZRyKCJaV7eOEq2Z9P0rD9qwX4OSbqlDdAqNYX5ita4nYvKggM3xXaa3cjXmfu
zMF0HR4HgDtcNky5wbDRCtspW+nSchY65xmzKPijrZN7xBbD61IxsiyXsoGmb1MX
4yu3gy/M5lszOkTyoDAk69h9GC1HrosdPLnG9cwqTD1PI/PaPdPO8PSPO9IiXrF1
O3ONR68UTV3QmrNj4rwvSlZ+4AiUDJEMDVutHteI0hW+ZA9qXd6KPJq1OEgucTl6
eUmHnhkO0Skujo5cOvMn4kKPB2YCBOCzrelNrThLsAPmhajWbjB2h0hjqhwJqGXJ
QmV8iTs0FvC2HDC1PK/6jvacNfFcEouv2k7gwJhMhyKABX8nb7vU02bGiNVkLZFH
VrP3dR6k/TDYl7Nv1fUsvxDsq+TGS4+PtMqxJHLRHypvV0zqvmdlmF8hRvxa12qw
Zn+Iu3JDEKsUxzUsGg1ZE+DQIU29gHrCX+p/gL2PUJmL5+4fk9gYFcPRDmXb/rG4
bTCsm9b7JEaXVBV5mivnFrPj7fFaK7YaTav7epOo3WxOaWjxKdoDUyUPbpAsQha4
tUFass8R4dSdRIVvLOb5v9WrNTBNaT7jF5L1GtXe5ITZpp3x/4/KgE19ymBkz/gp
5mMQ8hM4R34He6STt/wMF6JKriApZIJ0AqEugcE8xhR4Hc23EiMg52fY2BR8h/Xr
GHvCB3ztOYgufTfgiqicj+EClv/rL/X2xRXjhrvzR2Qac7Gh6RgVrGiUXN9kwbuX
yunbG5ilSUxjZLVqP82aDMHL6YdZMi/24oHxGfX7EOIP11D9oVXrzrKEqKtbcU9x
iRaInBTMxSnR8jcTyjj8StYtOOSNQ5K/8lqLpvI3sr1WfG7c+yGm1TAYAe2WenmM
1PIT5gOqmD1MwVwd3/+5uW22K14HIdLlppX7JwdT5GZyctzzOc31UMFRKen6ZXRc
URNK95Ly7AW8ihxj0QGxPBOs4dAxLbrLMpXmbw/mnPWXyNChd65IDIz7aFqDm1Ie
sYBT4wT6r0fw3G+GWo85JScUyvGGvDkdQXxeCo5pi41zlX0x07c4Dr+iKcQHQbFO
jJGvtb4TUzq9EEwXA6kQ8yc7qMmeGAEgTfMfnTQQ9OV/kJWkUlVXGBIwL+TeZvO0
gL55rYJC3sD6pQSeaGrrCGsxgTNwWXjoJs4TIh3Ofphn1M8yJXVhTZghxeajbAQ9
7R3EqfnixhNpjwTh9bk1t+3To9RFVc8Y2XKH2nYlu02+WXjbAhSJJOmZJON28SWe
xMHgSgP5ukXo42x4C9MQt+yKbxZPk2U/APeWEw2zQ5frAF26mnFX2sSS+Cinqr2s
CY5xiELwvCOj0LiYSb5SNNQJl9x2TR50uyaKfW/kx0jc2ua8VB8jbLerRa+vgykT
sXei8oI86w5hOV/QXl91KKPyY0XJte7AmxJ8yFlyTm1PQ3SXhgRk+BLqkpsqa/Ny
Fgq1mNpv111bdmWTbMf6bufj1uTTps+n5m93V/PYHu7LQCCwiWUzrOEur7MAqCdN
9VSt2TyyV4bI33ZtdEgaaSMi/Ifsg5hX27sNy9rbjMxZCpbQMTg7ejfuSY3ZM0Nz
lr81V6a4zLjykXtU4apQOALlUURU1dwVmywSgQzsUSneLga1ju2XEsj44HjpB3iZ
oQLt4QO9hDqyoYpLsznSv4QD9x07ieN4xnACThc9k5cQ1SRhG0P0vEfldTMp2DDp
NgLz8IDZ9JHyrVCrWF/Naqp1VCyupbABwMtwj5Im8YUicNW9+SyXuJ2hi8ymguly
D7yrzQriwtI5rW9RHNcTEp3hkz8onlBeDtRbhlbWIsfQ7b2hmarPnKyhIA/WEPE5
b0+hXu0rcahuQnixlNoNYveL1R5n3+QVw2X45s7t+Sc9EzjFj4r3Z9iRBN2+Bp5h
9X9QW5hoYnPcW/2gEWkX0Xv2l6tnogAzb4EmlFL+G82Oah6QxilnJWIxNAXy3j+n
mctaR/6cMwoacCSKPFl+cqjP7EJk+/0jGXLfxbemoBLmllJ042Dxhth28EDh+yAd
gTaS8lyvjHvPNu4pD9zubOEuIKAjxJgOXTpdK9YtNA1YT9D0wn5oIf4J438R30Sr
zymh4CueuavKxzUxZbcGKmkOls6rhXlsWCkv91weRplhGQ95Wt8/faT1QTNAIY/c
OA4BY1wsPPFZT5qG6VcErLFu5rTlfkD58C2gwvGZCTP6GBULMtYIBQeF1unPjYzC
qqAszsOQDgDTe6IaI+lo2AysCHbbI2ja1phnr7u0QljU5OxUXSBQzw0ZXx2qzd9c
DEVxHrTQTDUmm11trupWWDRAPHAlHptkQ5ndhLXfdW0Knvx/PfbX1yzZ77RCv5/J
df+zP2/i8lsSvUGuw8OHUiA748TOeZiGmT2sfzECrnP2JnFvthO8fotcUa3Yf9WM
o3Cw7JOcpGGYfg7ISiTDsUqLv2WTkJFapIPxFBFxLOIfKTuLdVFUR7geYRJTXa+P
P5ntY/F4y35aGErILMaDLHEE2pyJbMU++ixWZr3rntsAiwcLRT8ZvUBt6rpC8BkW
7HnFWwxB+HDivmU/bcpOcfMVWDUpnolA4pV0ALQ7ix/UnVDClJcL6j0MV+roEnih
07K2EmAb4YQXexrbQKW9aiSRndJ0Ipjl5+/ZN1JWTIPkrRPnyEvy5DyqwuMvtkKc
kjpyCmG6NPTdTA0f4AjxmXtIWKCBFD4uLao2X/PbRLqntzT0LoZq+XPV0/Q2ceB0
yEv+HNwFzWozqtKS6NqWVKfzylCdipQWz6SNdYV4luxRTT52YW9jbPcGxiIMkfC8
mDOLnEo87YnVyJBW9W01qscfbeD0MmtJP/YfrC4tfcn8M0s3mzP41uweUY+4bQKp
1V0EXXEoNHJZpmmdnmu7lvpWLNUTI8fDK0VoJ6CCuJ4buIhZetHZtYOlGbUdHvPA
QbS0AA+l72PG3ql2Hcyl6zWAgtR7hxTEzN9DRPctBR0Sic4MIBZidMC7X1hVvimk
iWz2nUXTW44WiAOHkhSeJxsLgzYFkDhu6gs4Z8FFfsXq8w08FC40hh/YvPbJz+h1
ZKQLNCF39i5GrTC0OsyuJ0eBRxjRs1zIjz+SvRpSeLok5Ij1FTlUQljwdh/JEOap
jPrf9bLbXZDXcdllxze3CvsyZ78a3MIYe+ziLXoJ14pnwaPCYg9zj66atP4p7p6D
fY6Fcs7GPnDAIInvByjvRqNLLno3CKOX+qg4Y5LJ3rBenXzNlwa4Yk2BTvqHOcHd
aVU/5dPyYa6sdcijJDmoU4tNppgRniEMJCkSmauO7cHDsJXaKgnzVR9YEV7BwbZO
vtsxRzCvcsRIFbQPJNKUu38/pIvp9GWZK2jHTM1qLPpSKQ3O5P6HQtw6PZlxP/x5
/HGBdS5/ElVBqYTAcil55WIXVLM5ILMgw6ir6oxD6YjYPcKs/DkvQd5FGtnFve11
s4iO2GtM9fbDJk2bYBL2b+Q9dIpYniVQLqttJlsLZf9KOq1Wps4pZ3hcGrg9h8Ik
eV2vrxGJNRi02hgXLYrTHbQAwObJWql9BUowVE8j/sYNZ5bibTNtrrRFTAsvFFAL
FCWAvalHIfnZPDABgGZAejG6QNDR9R8dytOCt90MjBqMLgx6COJDxlDHQk9WSz/b
EYGDB2zDPphfebRH/8tqi+8fP5RS9Ei/rHFskOeDdOsa9rnhcpxdnHxoFAB3AO8G
/XoqWS0ptYx8mF2C2GcDKx1uR+fqK68y4DTFIlwQUkDAGcf3PZZqZbdnRwsKIqqK
c603pMfawVoUvwR7eNDYHB90ZtylH+Jk8k1Sjy/MvMF63ZUlU99N8G5eJ6mS79Cc
8RA8uf4rZSpcJI086Q4h7nhEJKCYefmj6LopGIcVHp8WFvlKl2SXNkBLcq65mzfn
0D2f3JhQFo3fyyuI3+/OYRpHnaewREm5WVXbM0Is0YczIEINj60fn2rZi65TchYw
Vgh8SmXzjS/5bbQV7TfbDIK7DooRGtyzMMuYZDKeGtd1NnUvqa/6464VvVrdKqVv
Y9cfX9jqeK6dTVQVANZfi+j8WpTiz7Xp9CvSCims1fo5FAbSmG0nk+X7DGnDMAk4
Wnyn5+00KOXUlmLt38DefrfXzj94Ovxt/lF9BaohlSKSKXSKK4UpZgTx0vCxJpHU
ME28FGnMec04oURIstbkqBom3L1i0NLVCR3q1otKm7JBK0pG+3wsGU9aA2ceEHjb
gtySjJEZxr7i9/6zq68XweFVVipLQnAFNp3p43fzWewdquGYmd4Kvuc8deecFUP3
7vyVULvg4Im4Xxvieu+imDYUH292vghewmLDGNlhYBJV4eLg0ciESQG+4akxgtes
/k5y44OX2DIKHbXKV7neyOKZEH3zppAKxkxmBvA/Emwni945Tp6Dqh337dl+OvB+
cXxIQiB8QQmqcPCTbByTj+nkWgvSDEiBy07EvZvZeNALVyoHoAskEe888eWUJcgP
csaej31N5eoPmhCw8tDNiBePVKddOOQESeBA+LuPC31woP0PkCLBkx5XRNq1bC/h
zRDLzNeAaBJtXJ72FdMa55uT4R4rEe+AH3bdTxPiI0l6Dd9g2noGXZM5wZyQf+2h
FbDg9f/vsv9VaLJPt+jWCizORF70AOWu3GbTe090zi7ljkjhvG9hzcltRKlzh4GB
I0qOQ6NOvlap4eyAT32FSloRlusOv037zHdIi8wzE1A6zF56KpGq1+UIRX2U+4H1
qpD/MOcyfSXNgCnN5kDEOuBQQWpgNfdyIW/zrjpbpxA52pYXGpwOOOwYEy6d4E2o
KhvzMAXDtR+yGMqb3XWVjBSCxR5RTb/LbsbHvzDKgs8MKI9Lt3sb8KsC6NmyLuuq
cpBn7XtOOm6U57c6Nu6SoTNuelUabghiHdYxmCYQ0SPz/9Xnct9R+C0D8wGzl+TX
sw+cZ8fvvQoMbZDCSOsEaw3MyI3fDJKF/Zm/aXWw13ccYnJwExZPs4Ueeo/gwQyu
J+XxLSJoMCAWS/299BLH0JlFqvMqVi+zVJLVNh0iwUzo7LQOjyJg+TX7CnkWT/5a
7P+MiVokDGl2nusM/UmvR7HPpD8p29wEqX/dTbfiNsIypEi1kv4RLqu2rjgWoVr9
EBOZaCTvXwPMCmw0Ty/6q0BGQNVpkp+wuUlT9b/hydiYzqMPcQL73M+8Nau8yqwl
wgAd4kOsskEgPUjstykBNjwlZ9bKBjJNEofPzgBCELHxvUcb/JwAwDYIEsfxpKYd
bAYYPpJ8hSpO5UgCVEeekLHKdwW9k5A9wBYSXBzyyagY8Iy7yTix6o1HaHfXDuWi
zx+wTNR137A5ulxun+XfV/4FKjwKAMw5WaZnOiGjkTMdYYLzxttM8twPuKOyWEiz
TNdXlKzGAAmq0agFangXzMtT3zsxHzdUE+GwJfzcvwGodsCsqmLUQyCY+JmFZAW8
Uxs9HeJ+ctN6DeQ5QfQS8cIrHOs/LKUEGN4hV07TOI6VMWZcourMCzuXhLDsThqK
oeIDdwMxG3joP8lkpykyntTCHf8rMAtPcP/IqKStSXeNLLUMAaXunhgEtiRXpMuM
vva7zIAmT/CKZU/tlc4TY6+gy0duassXldp61wKqO30e948Gqcm0o4MzUhmiSmGe
Sn3VOmJ3E+lTOvwuvVXnERghOCtwEKSGdAdYgdufvh+frZtuLa2vKX87XFzG6Oa5
L1bd33sGfiFRmGOl7L/gid3SAKjTWDqsOclqP5Xytx3x/AFienbFrPHb7ndoy8DW
UlqmEsY82OYBGW7fT0HO6IkLEuUaDiDqbJ/DFAKgsw1wf7NwSnI/0mOxpau2NEOm
2jVW6wOtgDh/lBmnhmTl3O+C6fTCC0SWef5ulc34a9EKUHQ6InP60Ie/Mye0WXMO
JB3Pb6wcE3/L9qaKPUqvYp7gdNLU2sCPeTBPDwXFE7MFJvj+KVHX+rqd11wVIkbw
KbtzYcQ0oG++jB79SlWWrIy9BlXg4xGeZvtLX6La/DOblgw9JIMc83/Bh065va3U
4tnfyGjGGRhtMd9Cs1TJRCpsCNoWyKhbpJ1CScV/K5FP/d7ndzct4xHzxfL8803b
bm13Fk+mq+l0teWN64s3+UmWRxu+5qFCh0uXXB/AhWaY2tfg6fmvAYjKsS1O6Wg+
x6s3iprb1UPLlIdNwLi8FTM+M4oe5OAGKLOhKndoRZWAtEuLauB/meYR2gpGRuUi
yuUZgjB4k/ApvaEv1aX9S0jXCa9XV0/mkNFb8EYtFJ34FQvvuLA0zIRyNykFCjqH
mhS5k/6x+mXEMsluo6m4wZC4CshlwYdhPS7w5+pGscWGyIvguu3LYEWVgRUEa1xD
Sx0M6ZKl86O66rCHFjc9ISsl73fEyXAeppmJ9QTlvaRQPO4bbPjC3XrKW4VhX7at
OUeebS7FQk2KttiLCohnvrATcnnI7w5yFMu+6W6cc/h2zA3IP/rzYBgXKFyQUIYd
uhhevjEFjaV1HZVIDWHUdkcTZ0JW1Ri7GC+ka2YXmpxLEy8D+VBfVtzL2R/9uJt8
gqsAMHo8zE2kJZB0k04xTveQh0Krc4DZ0OYPWc1zDhfgKHd3p6wciUQpNK8MeZ4V
b2T3t0RdBcPflx1NmwkeN3900sLpkR/IfRys8+u54HndBMLWnD4H38wZ5PP+IHxq
0FameikOM93+lmk4A0ASbl/uoU6c+rv4WdojhRI1q52E4O281pS1AEczXB49zVHV
VTDK0jSIt0G5dbI1+JplXY0jPwSOk9dchZXjQxjRzYLGJha41T6ZHobsCoy9ND8a
48AHKuuEE93e36aNt9rIq4AxsXaWEzdo/TbT0f2tjR3jGDQrpZihB5tq4kxLAJEI
ClNE7nOC8rift+0hDNTTXJdK+UdOcW+/kPpAZPslmRZM3Re2XrCfCaoZpSvzj2q9
j+KQa8Rs1V1cuMcxxSjG8Hs+f/GYCT9nJHb05mgaqH06UpBRz46vAN+3alCe9DX1
sNUeDjdLy/iquGZhL3sYHj37aphkjUgMgfiiziYW4HfUPxJ+je7hG+MdSChekD1W
277OyC2Uaty1kS+iT8lGcGAhTXVDjduuvJNqVmiO3phWj07lvz6IeoevTNpnh318
hnwf6r8fEaJcV/BhxvSKNrWwlfw4ynX2CVWmuy0iwlspnNuuBp2yDPgEUVrQxaam
LpwWSjWxo9gW0ZQ7eNtDgAMMe4RCii5VKEA5uhSrVZJTq1ioZnzbvWbDLoaWXjMk
mEqiXZGv78VsdZSasARap2pPg7UoAuLSij8aw5/gdXFw9sNyAk8Eqa0WNLh0rM5g
9teXx0R3A7Bk6trNzFXT00tQccnvnDlL6jeR3LSgP8Wo3VSvvlws5ONyBlyWFI1o
xorJ6ThnVPLg0tRIMOMLCDSX9HaHQNBJgNqKIoxQADkynp1dve6+edMYjMZWTK9L
z8g3VVlmbB3lchexhFOqqEwtnnpdrXrFJbM6ZFCRc19oZE+pSdSBUTINok6CD4pV
bD/6Ua62Mjt5zUNNd27NTRUXxdX2k1Pgemo+wPBuW5fzZXmCIKUIuhSiB3IHmikl
WpztggdqmVXVMaT7pVLPIUqCQr7+ec0DqpdGJIBejfeh/AUFyNfZLRCfvdW/h1BB
O+Or+SpXcgCtnuZzyqxiBo2BGF7qnK3pzKm8/qPvkr6sa6jHt4I4iSR9bJJQR0XU
ebu9oS8HUZA9qimr1bkvxDmzoMTm5goMITnt/iCHfcNhhBh7xomJKxg7lhfU7sAO
mQ4sFLrgugnWaH+kALr91ICwbWY40iLh2rfzPPsQu/yTSk/VFEppkyvZ9oRj/kvN
ty51TSxuB3jibBx4MjxDeTvFk8r0TiTRLY5qix7Z38r9meb9t7+mBIPanAKHGRhH
Mur8DgwUcTttjC01Wo8lYW0wlnzcJe12O1Md4x1H2QEwB0gLTWxjveAOZjeT5LZC
H9KjO+spaF3K2N0TUw0D9Pqt0kEDBhenOeIjwEvzmI+bbBhQWiC1SLPX+xl2TyhX
1RxA1Y1bCuWgAxp88WSnZIUO6zeeMUkHIKUz2CE2HaK74XDzONK1373YYcbLPQxE
FANodUzV1pyaOU95vGhcloII6av1x/pKM9jXLWcsmNtskQ2cSSi8M4z4+V7L83K7
BptGtLQUvGxtRfdcLy6SldjHQD4yJqkKnR1eggjLqXoR7Y3Q7fn6jtwtBAn1XV9w
UvvkP7HdMN/FkRyapRxH+/kwgqq21108HttLYEs40j4TH3VRCIjmqbEsF903QSk2
2qm/vX8T85ibA/D2n0PCMCsoxXhPccRNiNduLE2Ji0kjkEoro74NDSIzIWQ/QJg+
gWjvHvlDLn6MPl4UH8CHclpOOQErPPVVxvGlUh6MN7sQQ3gnq7svX1UJZ1vbmkj/
/egSAj05Vjb4SM8qYBsHXJ7YlitDt5c7mQ//HTzjwRj+ctC/iOGHqhf3yPs3z9NL
hLRbkKpdUruuyDsHyKVS/VWlJNmv01bHQpJxAPnQ90LWHTGyQ2yrUzv2LBat3Kqo
cC5rWEzUHwAxmg2awHAJQ5ENNdq1gJMtSrd+fONdgU0kBnCow/y5DLLs2cWNr3mn
I8JpjTxSFi4CEMW/JKb+c7fPUHcm5VCzE9lCXqdOG6485XINU3FLd/v7phsFiuuN
ImaHGBE/RcywcqcrzC+PXeQjgyOgoSSsrZt6mvNX5D5HB5KdQ5hsOgHKWrv61jdb
ErHwVySJcVSEZOQea/Vorc5BggPk8TtzPWFbpOH/RznNBUP1aqOfqtt0uC762QFc
7waixWB+Z64CtkI7Tqc7y2a1Zy83haCo5M29uwdmYVDPAcaj0XpovNy4l1b02c1v
ROJY2Rg/9ukRZtEgc0SDykEX8os3SSZl1/IBZEUFfW/1O+PFt9aXcux5HN5r2Vbl
hNTsTz4RChhsCE82QDH/szxtCVHR354TN0khpD/6amuVEt8bsXqHCo+N+gC9KioK
cqVKXNRMmwKPTUrUzZ6pbU2f9BJnp0faob0GWT9WLHoa1w3gzFPbVrgFVPCbTCGD
G78hYkk9enH2/T1aG/KF/bASIGltOtjVPbYpPYhanvo+Demlil+WKaeIdsHyRdXj
dw35yYVNnYy+lVEtoKD26FwNTInyaoOA9FBJy+1SFcehERCrct9lfcILBKe9gzX7
JfbZvra/5y98tIjk+Tx9p97Yf3jIGEL1bDBiXZwXU0oD238vEPYHCxNmshGIWMtf
aENQ1WS8LtyM3L0pYy/hcdW5Wf8WLLeOFwIqDVET0DK8Z9ctqj+w28lwh6LX/PbM
8TaBISuYfe8Fqf6Buv9z0oOx0MywWlYnyU60rFLZZL9Gv58fFtgrYolQ7gvVt9Jw
PRD2G03u79+OOuvG2uXLOSEACNQzKuCurq4I+0Z2yqJWcSiLk7pOFti54NZ+p0s+
DoXvXrMWnREU8KoISZxKgblToe83wF7HSScWDRcgdD6GeaglrLD+ypUQ4iuSstoX
53UBHx+418VNqgTxl35Yx+efLzAajYU9I9dznUdlMR9N6Tr7qjPUJvjI5/MsROhq
QnUFQ3MLVSZEbjuM0WUxflodg7Z4m2nnwQreHQL1h7veBN7Lvr6HiGQooyxLJUHc
2wxhMJFTSbMalt8ukob2mhofxh9Vsa/lzXTCtydGHkES8D5qZqJ6FRSsDisO7135
lDs8NAYyzLPVsenwRO4YXtivUiyvFMKd9HU/ofx1OiUza4txBFnu+CIYoblkRUJt
M+q/jyVJIuwjcGXpH8PYCtwRuoJSICzJd5G+JdYjQ+/v2K3FfMOr+MYRXqiQhLef
Cd9X20mxpeZ+6VFFsoiWKr/Pc/hffh+pk/rGf/1Tni4LJZC00cxKswKwoWkNnPLd
2jarEGPlHbak3ewZIUgdchTaYDTZZN4TGuktL/WCTIzGY9Jor3r9Uts9YhPvP9Or
RiaTcx2DghuiWRVkJ2CeVwLTSUbEiKhjK6T/QFVZ9MJCqSzg4YGpY1WCP3XG/7DE
9cWFutTTmzlcJ7ZAZmnzrLLjHKlAThOOv5A4y8X438wry7eR1tByZDkY2kdD63DI
E8DdIPmZMy7Awj0QM4Ujuv6Ubgagl1fbeLv7FRPkeD9kVXufyJqbc2pQZ1VZZ8Xa
BN39ui+3ak96rc7J/s7T1lO1RUMQiBd5foOeTh8A9oZdniOZazj1Z1p4pcfrWEqS
kZeVW6qadx22UlHAnCXfttUnupfOubf+1Jgip+r8tc2w1dIpXJXdKAbnU9716gGc
pnnjsziAfuTvLOPxxtsuG6oyU5VJKFnHOYVoWVn2rwUkwzlf0XRJb8GOWWdTzG4R
3eV8NcSZRXjDo+GHuyfnToCQXuy13EeHUnUk3GhfItIsd2VH5l6jLzwzhi2xrWAx
pFjEyWLQzTfmVUUy9VjXk5gqe0Jodvc6UnY6kX6DkZl5JQgIOzmOcakhT9COKGlk
z5MOXIyjB86Cwu7BVKFqJJwa2gktz5OEd9FQDKe3UUSpirLMbzS9wb6jeXDSysOF
5PdS62+2DGlnhvlnBiS/bqAYUwNTyvwymultyiZyxyTQdm0kIdfcWDUPytdMdHmP
2wruoqBnqgxwDmpbtFlA9AQC+PMO2UT/pkMHX7ZWIGd4WLfvBaLqKwmuwT1PJ93A
rz0Y/nbiaGDuGzshORPjATZMXKwT0T+HN6vd2ClDhejBt0U7SjgaZnsnYHJGeKa2
auaY7VmQpw+kHjLFPdoUMwI4M6aY835A6I+mdmCcozxku3f80fa7njxaYGbCKFwh
mR8st0TtgRRl/TgNi1lxKAOrCMa8/tAFhjzSz4fqc3ri7fssVJutn3GSV/9GMtkH
QvLgbud/Zu+ZAPhmlHz3EkMN+qPTxqqpIcRIHj0r1mveExq8oEgq8qyi6b5DZDWf
miU8gBiuaKplD2nzRvqbY/fG1njiKP64hoVEDMhXjolXrxQxOPS0jq3lFWEvSZOy
NEY9DNJpZh6zIawzpYMwUC5TmNkuBfXjIL2pjyDV7nLz6/24FAOByNiZ8w/HS1i0
uGYiJ5SSWZIs72TdcyJg4ONvxjTYryNKyD0aQGfrdEpcRLFDw9RJQUq5P3WScV/z
lVfGDHNdiIdQRuh6yRdfU/GUQvbl1hbJ+IiDmVr6gSeJUKHTz04To/XQKrYVzPKO
xBQQgs4BGAK0ZV40sijAHfQSUMPuI5GRqjf8sia+VP2YtOwvzZH/HTBGS0BI6SBy
PAsie3ZAxHWrDm4/oy0OcjoVwiXFXLzkZDUE4pU6UBlUYjz2UYQVnkBnNhKu/J/X
F9QJI5gELKxHwuNoLpVblXft4uwED/sv2gFxYsSthlhMHnECpC1kdJEs8wC/Bdmb
udibH25iMG2nT7J5v22WAlYOmbZV0RhPk+RNzDH6Z8K7xIOTGmHj7VcrlkBhlrDk
eHXgnAmaarGqtklqJVPAV68XaCUKL6gK+sycmRLGOfzRjxOe6/6KpZmdzprZ1qEI
Q1aWuoooC1eOgfuxMMaIYJtvmMRkDfDnncWFtt/+pS8+POiHkNXYEvZ8wKLTaFHE
5EiD/cpgYn80hriGxFLZWXJ90z5GdWdpoTAB2IKcdd7eL71qT6YXwJry5PnrL8La
wxSn87E9MTwRX/m8+6JUI5MFLtmNTQFuKzsDeRDa+tWcHBYuwDM7D3/b6NU93r1Q
1bYHBLFKAUiMf44gMrRmwEd7v7t5u2Typa3oIH5UoPdbyqfykh82Strbk4GF7agL
54QrRXgfRpvmQaTHBHL3UMV+ZEItN13g/4nT+zVg1r/ewpqiWfdXua+ykALUES2B
33eEf5UZTixiVYJe8sjBb/GrXcOtZIkH/fYLJNGBogj/OBYBRSS4EnqMjAvip2UX
hwHixtxWdQR94ZsEcgceLdy6+9HvJPfUfLfi2sQhtzXImaTXu4ba2cm97c0/WOHl
uHHggIfafqMXA5YURoNBV6+jckE54ifXrgZYbrvgFDSB950TWH0vPQE7D9NXr767
S5uP6evTJcPDD5b8E1m4zjvC+dVJsFeZGFkELRau7YpM7BTuJDXmpzsUktfjuPO9
NKQWf///ft+CTFMGc+uXU7J/Pn27euk0QC18ILlR1MznB3ZS5PqqhyQkdJSCmUq5
QEY02Z6mYrBIDNCod75NkJRSuXHBSXZmoE59ly0/inwu7ygstNpFvrwX/R0KuSfA
PenjOSeyuwLKuFje8XrHsrjbiwyk+XOZUgKF1TCaQCNMq5oaNO4fRdUS3g74+3qt
G6kmiqz6nZjnWK9H94FIu9AR66eDwW4Xq4rOsn+Tu3sgTJICaI/QhSx9Bz1HAROV
+dUt9bAeDZo1RT99UwvgQJq2thXno31qwqF5emAmmtcvAieamJ6+4HRAlOhNTkMp
NSJYykhSzfwafbBtxChJa9W62ZQ+vjjKHA9tNuWK+IK2qwwUKOTtVKviOdZyVHwL
q5Q3+Tz08Vxs+XM1xMOhOzDx8LhOLJ5yJ8fv/Oci1rxU6EKH25l4xYiUXfnYmlAw
uO1PxsBo4ltTMZbZO+L1BB9QGn5DsMWmhlk17kuBNymWJ7rbIBhvDiLkTDaYak16
CfbD0nYyyErhzvL1llvj95mF5VLWfxKS0T22txE7p2X4alpGKUxxlS9QtQ9IbmRj
7LyW0HXdiNkMh3xbkok8wC3zUlm1Gl4DRKkusMScNkPA+KlpuWmn14xD4BVUsH0f
R0ztim3uoYpKhRWdrlGIKw1S6OvBVPFNpsEc9BT/f9lfC2Vfu2vqRsy+fFUs7v0J
BghsO8kN7xD/4yvwLeuYRJ3o0BcP15xQ8ui6qnK8WvqezCuTfHSsakHB6th6PVGK
WSaksl5T+jqyFiVEkaWMHzYGzdewsLsaSHGvp+hOL9f8BCZZb/d0UkYx7rWrQADF
Nog9uynP/Kzl6vwVjzqk+yMEZ9h6DUaHpbIC2gwI3cQePB5/8TefDe1Ow17F7efm
t24p4YZzQKq0FYjtHWSamGCNCrZiSRQHrjv+fkM4Cz3YwDXBG/mFZ2NJPscHLPXK
jflqpBXSBSvvekYtZu2d6lfURGTZuWQc5gfF76OY10lS5ONpo7UogXoEX2Xlh2Ww
VkydnViHi9hEFk11RUoDK7iOYVNqDd/NIjdEYcz5lPk8G0V5SvfnD169pEN5PteQ
6bDL1jj3GUxX6evBggmgZHoD2NfqXkqksVCab9P2K7202rlJMA5JoaVrt7ASzDzQ
f4RODqqK3LSBwQQyYBNKcMAPz0sd4Ge84e/khEjWp2jUvwePbMhLvYJE1Xcj6E/d
OOA46b2x2NOI5edbAM3u4BvfTRTDOdwcMZBxZeY0c8bC3gudjWoaMH26Ac+21yRC
Trk2/mvwWWtdpg5wmCtSrrwMaHMkRdRFnO+Xfx8I3Jt6UKfFtW0s5iBieSenYWWk
ly5JWrfGyz2UDQO5HlVakgpTpud+/+W3RM7r6mZ3GdAST+ftZEz6NKlHORFhLn0L
FowM/wEYFS10BGO9rIhaQpCBJN1j0l5ioT4d0xjR+aSUGEJkAnp1zTYyglhgVKUG
a00fd5OK6yJqriUkjgr0vIFVJwUeeAmQovz27y6p2tjC7656j8HbxPU7iNa/g3Wg
tZSPGGlJjGuNAh4fCYDrjEMeafvdfmU2MNllswppkhexabNP+2A5FWXsXPy27vPY
wyBt2XRMpT7ZcKBJzSM4LH+87TeZ5EnOD7zk9HOcO8xwWvZFPiqzOwozehzJGM81
OKxnR6qXVkfKtfuNaP8/zAH04ZgkHI2JJ4Tcr4C8UWM0DctQnK9Bacg0otBgs6s8
0A2MrvLjf1kphmTtg2A31EGiFko0ha7IhrqTHWcjWIGLVshjlg2DqK3Pl09WgO6F
iRUvMi4hTngdseqdkN21xuffg6HtuXcbDkAXSFMqAnCcdEEnL3XeHuUA8NhfqzPo
gAC3Q/PzIRY00RkhTobsvhM0Q+cndLLIrKLL6w9tJ/XOnoED9eBgUQSf1oIorh+H
+Y3XjzVSSdNZqLFfmT+kuS9FdG8gucVJzhg6F5mY67vCsn2s74bvdXFC3pzizP/H
AbdPHs3VQDVBYRe1eyuIQ6qZjAqnw3Nt83gwy29wXyb3Y513W40Y0/KjXsfV7t7Q
Um9YxeSWlBM5zqhE0cOwCON7xbT9AWAs/1rCFgXyNQf/A9XclLzhzqbKjuycanEO
9nxQGPrpVTSSi6SFJvrAHCauLM/Upf7Z2R79aAXAO3F40J58EDbMy/sYvg+Bf5r4
zRZOtsW+aTVCPsjvXVJ9hnS7+Gfbt5E/hyDx2hYcuVen4WDrbfOE2+cU9IZoALvF
j47TFJu4Bvcn6IpQMWRu6hV1OiA+QbIW9fd/kR6Qvp2tiEz6U/KOymPnzWX2tebp
K+H75uT9Y1yUt2rJAJlhEV6xtSUcIgMQEZHSiEge5K5HuvenFg870I3Q5KYd94YV
xqxz2+g7p+VyR+oFwPgV3Y2NnUGHlDjzimeEwtZ24XaVKSySw4D38DIGr79b2+gl
uVKxwbAq5s5NbGKYdEbBD7uDZTAuDMRFbEKm6FJAHZCAsczeAPAUy2oGTU4ai9Kp
7fLnMdINR+hH+fDBxKYf3YOQEfz1ufap8vydC2xKUVmVMa6r1mzlZNH81BApGrWZ
xuU728VE+ELkqBnbx/Qs/9vSoRPtXLccXQWkEURhIpHvOdG5fWOENQ5gmmzkbv46
tdbS833cXlGBg2ZALs/yXrv2qBSRDrIHkTJQ41LH2qTFtpiSSMKkM8nMSAfjpWDN
D88MYkQn65etZrdIDyRg6vAp2ISfjsYCaainmHzAPrQqcJrW/NjfeHD1c+zxkgyu
bqXML7ZqtI0dpvXto4DjSK+KXpIqSyiLUV3Lgqoa/nw+Nhpd1T3JwSXTOlhQs9Hw
nzxSfThayLI0a40UdjxC/s8CvvpmeQFI5hZQ8j2JjPUoAf4rea6uNIkKY/wQk49+
GAa53gjEERKrILGRjxVGAsjvad7iJ0QuI4lGSrhTpyahTLjSDywkHmHxqTKNprmT
D6owWzrx7mvqUM+ljhNqIWb55Ksgt1WooY5yRy3efX2utm4TlShe/GvScjwQCPK6
1YaI6AITK6nod03rfME3MK+aiivKDbIAh9yCpu5ZDyEUdaHsnMAEG1uwGhOLa8Z5
5uIMs96LS7vfrFb/wsAo/Y+rZrfJ/6Nr4b8Et9w2h7RXGQ/BvrK+HZdfxvryW/79
TC64y8I6gy7Lq7hdrNJQN57nwwWxaqcNj9JHmHPHfNFA4PFqNCt0BZP07YMa42zd
qzZVOWJCYT8nwnNtR7QfR2/fiO6/ALbjNlwTS+YVSdV8JOQ1wHbZ/ZsldlC64JKt
WOiPZQr4JlBWY/yGutkDgmqb1i+dCvrmILeWCJgZ6CD5LbUPCgkH5CDY/2e74yZN
OEbIlEqi66EOpk+t1D85rrh2C/skzS4gOdIl5GGzHbsInkYtN2dDHs/uekL9jecl
OMm0rzNN8fzhqmbLaSsUq3Abz4KgK63xZG2BgCza4DI35hjz3KhxmZhx4gETf57c
tsS0/mYuEppccDRjF6Bxy4Ze2jynfYybeEtq/iwmDiDY9shuSE4ata9UXfA/FhXx
IBXukPFNgihkg8YTKOQXuOcmrvhbE/KulyHfbBvN7wVqSAajeYJEvR4+FWooRw43
/OMUm5PCe47Pk1+iGmCA7gFERRrJkpU1H4vPRofzg7Ejtvt2O9iOLSaGZXNWAeDJ
QfyufyUhbCi+7VkXd1RKm9ok1Wm1VetvDUXByU546w0nbYxvFyTgaqsdqI5E5uj6
hnC5/qoW7XvugMxCpcESA75/CrzXqXEB/AhF8TLKWtnaf6t692Rf7QAUrmSCKVn1
6PM6Us+ODNH0aQjfQaERziBvGtY0Hh1tvyuLbUZOZWrio6hHfe5LVSPml2hrRhXf
AIvBz67EJ/Fb8VeBRRk3d7XD0CxlPRm5j3WBJ2rpGfd7AjFjc+3otaXOg5nbGk0q
blKjJ7YVrnb2WcIf1KTRy3uUssbfL8UBmMp+8oaMW9Hu54vCpjCs2zccs4Lp92Od
mgb2QbgMEkrYd3MErDoNC20wv6WBmF3Xb6A4mMb6FJkEixu6IZKS6uywR8jDReyi
4WQJ+awx/V0QuhKPx4SG6LGxXzFyMtWPEI+9h0gWiJEyUQJ7oXM3R89Hhr92Z3Zg
1NXJ4x4AXt7d3wQqtyHpN5I8aqM30BG3Bl/JTSA/r4/edZfb7RG63K2lrExTJIjJ
vD4LYDSaMPrCO/5G2G43hxY6YHfDE4HE2G5h9TAunAlbp+ShCQUyN3E6MU4mbsBM
ikAvS5oT3GjpZf7Za5RK19XVmGUJEPlEpAc/RTKvbx4hXDUd+gjtBvCnJ8eVKc8W
U6c4vwoIYaEvTnFEU46LrYDAC0KWz/5dcRJdaXIWbCeq/VUBODA/uwv0o7wXWDFw
DkqE2mykk3Xz7Nxw+oxQX/6LYekHDcRqNKxnFnGIP0AWOC2Ih/VBFTfBWgIqN6ot
y2/1IuSdoS9ULy0vNiZ86kOx0j+6DKAG4tUZ9RQ/p1gd4EbKCDhLiUtzP8t9fNBj
+qJXr2Y/1IRIzVUuc2TawBjFNJt3V1Qbor9mEZnr0csBAJyLFd35DnGSGRqKWhe2
CO7Iu5nYjKK1WwNe7AqVNFEssKIiOUs64Mk+qABOeczMWwH1ZAPT8EKmh3bYBZHY
PJnYMVm1kxr6r0HZ9T99nrNVuOYJYNiCh75Pgaf4v5WwTfDJckbfv1AY/F59dvsv
lhyi2U0n33wKXzjzcxFsS2f4lmvCrd1I6ABxNtb5YC8cDZn3PkAtA+4+63qAUXf8
D2gtSsfBDQSTrvnngUcKhNNAxbt9MuKjFCnWNZ1aFRxQMpSddWP2Y4YdAE2pm0r5
uo8NnI76lypJIK8OKj3rBz8gXFm9iQWLGEl973YWns9Y5NKCStHqjx4ObhvSQTs7
B6PgMT85uZVyiQcNXqkRMDkXySkJMxn+IkJBKeGwVp3+yBXuCtz0Eg5eAl6y64CJ
LqXgKXk/EJVv1zBHipb/3bpniEacug3t2LDRNRYm7hh+MtX8+0YsUzNiRTWMXnrD
pywk1Lj18BgnGS+/odljN53OUzmS2SGOwC6IldZDKb/GIihULinZHuWy35dy7jZt
FYreRyAvcikzKk8fEJSJv32kqo3dQBuUtzPXEr13axJ+PkZFktaC6ugGmNXzwWke
/XskD9ovaz/1Rpn/4CRLL1TdqMagpeluZkPYfmTftNoJnsVLX+QkbYEzj0HHCgDy
3AShMcEijLTsdDw3EPWYfjXHlSFHhshSEz2jQGMcep5xkFvOk+jTUM/J+NLfrjgu
L/qvNu9Ja4KJW3BH1wWt1+JDLPIrnAvxQK/GUoovGqZhnBnBDcPupKUq+fICBC5Z
8qmFceobIBR+CQvr0AiLJHLidqVQgJSU7xT7eAu3hejxY4goiAxXzlrZXwVGD9oY
7s8u/is/8/4pBYWoMJxzARUuf2QTJDVOZ52GpKQ6euhfofr8AhHGMbtm/GAC452F
nf1oBDfWS9YgG7VyNy+b22+y+HLeiYzJDiXp80BRxzsOskMH0F64LAF4cW6WnO8v
z/Nzi4ysQPp3wz0LQYSUFLo0MoItb1CvcaiGBvlcH9pezUobmK1nIz1p2Vfnywjn
sXI4AOeIPFpbwi+//guPEmz96q3gCobEAN3WHjuGGTtw68KENoLp3VKBK537xWD7
n/frO4u5enLV9XjELKw394xhq02cjgRbU1GYh4HFKQuSMRELzS51ZxMHhOgNu7Y4
WNcltKAJ/4nMKt1eAe2cNBF9wZAwVeeaon+Bl8g+Avb1ZyVWSB78sqPfR63buswB
guRrpFWA2Vpub6+Er8fb7kdFBUcl3WNfyKYdaE0w7luRlGWhHatuLRVKIz/DQ5pU
LyaIMf/CfmzCLLItcdC5JzohYr9srJthuNz4wKQkKoi1LU3SZArXXxs1FlmA0CVM
wgwHhtE7wMSj/QLRFh1jO925xH7N3v4WHSoMq0Lv7xMVxOouZRWjYYJXQDZb46sY
fi+WFcNQ+P92WjUBdIQs0ACgedM9/UUESKsJMJUwpTc5hJApD/bAFCdsQNYmuOGP
XxmboFPRUYZxwfZ14NgxmvNVzfMcvQMHrmpdQ37vl0QOpf4mSwNLFAILC4oEMlvL
caLW9oUZvfztdmST7bcUSOEhIYqG+oK1YhjqpS9EJ29RI6cntoAIKSx2M5mvaS1d
OvHB4shocrg7oIsC8i+HrwYqpy1a9sZeuYhJZ1Tm9jOI9RKaaYn7+jP/bPXmyafy
2L/XCMQ/zQ61Z87C9zZa7KA8YRxondEsu0ihv0nDVo5Twex7IK3cmZn2kGNzeFRE
GsIkpt6P38L9QUMUjvIe6xpzix0cWuYgrMlu/aFbX2JleXNsGxqnIL3yqEvn54q1
/1qigfPCsK12+F0E1drwPsfbjxcWVtIAOIM7RxDOKwL5fvcKJvk3wtEnJ4NpYoza
ZhLYQ+Fn8QS7Hf6+02KMbpjS953JCn2YMwagyraLMfAXzd6hHyPD7iBymzKQKzFR
WV1H0eX7hQk6PApPAwcrWeogNw1WMozPQvB2RQ6OFV6H1SEcrHbJj8Qa9yaVS5s4
Nae5vSo1See2OmIuzkv5GpJa0vCGbrYOZwLokjIFYOM7zDWnEuOUvRUtpzg3mZWl
NeAaFt8AxVSAxbPdusYvqn5uqDMJb5BQT9Xb5rqsEZToH+NvOqCtE4eR0nqhbJYB
BQHj7Oc9R2gB5OHcBz1SViSutLTaYydceOz/DAXrFyxbfOyjL9l9ESzpNhYFvRyz
u2CF859Cc4fbTGcGoVZ/oQHq8KtlYADovA/5aPycDY5H9vON9fDFEVrHSYHPhF9u
tCrD4kWQXWKrjGpTIU0pPXgBrBP9ZF78vp3m3QdSZyA0BspvoTAIZoa073D+c6yq
iPr1eKXbrGJuazF4qVd5W3qY7isqTDPhog9kolVIwLFcDMijqdJusKA1POOXj+rh
mMWc95+03yl/yVKNhQfnRAawQxrTVtjC2lIsGi6SXoA9ZLUkvn8KunFnaJ3E11ua
uZoqmqv/BYLXSbPODs2KPVYVzZHJdm7jaWpAKBgcN+TVZR8REE7rcMHVDfev7qH8
QjppTb5K6Q8VTwxXWhzO+NNpm7pwvKYkXlpNDK/9qiyjlwdLrCWlw4u8rklI+gKl
3JLteirOwfniuLA7B/PLu+zqoqCJlvnMH9P7nAEx+oxNxtVzYt6vkfb8Fxc1f3yq
BPXbM1/FuZPXV+n3YgxLDwMt2gxH4HWnHI/cZHhvhpGL4hay2LmLu7P8WkVXdHUN
bynAn+u6Bhj3uVI2AaYA7nH6A6sxHVm0ZOD3O6SvvfdPLY0IcsrJyLkac71liEWb
kK+0DLNJtgFLVLS9vI0vI1hjHu2X03AIp7mbPLuVf96D+pkyzZ8PedJ6PtQla0Kk
zR9lvXpJPJvBcpLpgJbBsKZX0oiCh79Bk2JdvmgSjKCOU+VzaA+CM6HRWmDT3l8a
KOWjtAJpAuQvtMVS54qkSXs9rKqxduxHfx1paYII/yphLl6JDHuVj4gLNJUYKPyx
Fev5/5qBmp9SZe0xnPXvUxSiYtw9sE1+kT8153Tr0yhh6etUBiZf6QVmVeDveGMG
u2qrVlQO4BYYSSrrgJ9aIzSP3B+21ha0e4tcJqAWRbr3vMCiEgNJ1628rQ0+gMSB
JwW+LpDRb1H367OTcruIWuteiglkmSttrYgojHGEJTjuE8K2lfIzuOSAGGsFBIAq
0M2IW+Oap2mUl6FheoQNd36kgOq8JA5tn47RHcKY429rqCs6x+NQ5+z5yd6hO6Is
s/Ksn7KPJULjIzEKXrRgNxxg25KBzV6PmvtZNT05yiUpMhi0JQ6+2z4L8of69wSU
+MwMqigNV7wKjJ8xLw1/cppTakQxmhpvMCqwhxwQLELl704vb88a8ZvK0OTIG1sQ
yuuZq+lsyT5/M5B9uBM4utyRLVpkTJkIZu0RTcPsou7u3reKqRsIw1m0nLo/TlnQ
nMPpBSk68qZpYLT+FVo4jYIkbPtkRvaVSRJEsu8x0eEizk7oKWLDPDpgzC84kNJ9
d/J/MOJcBsMJxDL7ZaVrEh1B78TIVlCEGmyjHY8NqmOIlYaKGW7/7j4pZhtzn88x
4dvbIUjf0ggAQkL5x5cPvv/gtCSloBnjs3o2P4ayjJMYpxDsD/YbbHJFTlaFwKNk
oEVwHcAB0ytw2zIHlu/a7rJed6d3bvGXivHPYCA1GamKtHZWv+JmqrkEOkA+zeFr
/aZ++w3I7A/IKqCGfz8FppfLjZQs/t+vzCeduV4YLfC2sRibWtuVzGZSKANqA6MK
zdohS/9ljx78cHIoHgpnZfg+1N3admWPt5mpBHl/a9+xErQ95RQVp/binAtRv0YY
RFNwZsktot6/sGiKt8ucsB70znepdhZ4PCWutPA6ye7E9GezfNUTs5ZiCAr9ARUu
cllfMGHrq6hjA43zMhNaTwyjXpWyIyA9L2U/9zuiW2O5Qz9Tv8bw2juvsuJAhDNa
Puhz+ay6RET9nZBz8TZDhQ+Hf95i+TG+T//IrtGiHGG01cNiXPSyHBzVScWF/053
h4ezi+WQ9BWPwIcyLHtjZb2I0bAxx5C7HXsJYeilMlVZegkoeAMExBexd+RtP7Ct
xGsjn+r6Wtvj4Q2xbcZlPLGJMnzf8ZL98dyzYWLcou9IxJnZFKh0SbvqwBZ1feeH
mHTIKs9Ij8t5RDXUuJTfva0LFLiglhUXjlOcHEubHPrfN3HPr58OXtRG5SHlteBr
wuW3z1nMfQez7+OVC91xVWmhG97m/Bmz4x3AMRq/i/Q1ySovHZTn7UkVi+EJg+DM
/BL1AySrVTKnRekzOLreOe2eMUFClgyy7LV1b+iUE2hnED4bC8jZlnSUpcZs7sXe
hYv2dABAUnf3S0nGE3aCBqFsOtMrHIcmQF6UHllJ131ytgN0QwIV9PnzP3Jgup6O
tjTRFiCND01uN2L7mrcGDPUEsFA2sUJ+QR0yS1o9eqf87VKXSnPryWLnWlhQ1zXX
S9PMZqyL0Bn6KzOuNxVH9DbKVZgdX8qWxKxhzzQdamEd7IVruNQRH/0krZbQ/9E1
aGc6NEu9e8z6Rh2nuiQmWQh9c8ff4R5/GCBw4+nRCuSNttAKB6Y/LkUhwUdacRot
YnWdff1UmT41sghk2b0PPyOYA8lEtck7BsvIS2I2oCVuRGFMdrUawkXuab6kEzjI
HM03UVAddc2fKJuvgNtwGDZxIdFoeVFe30vZfemjygvo8EUyk5P7toOkAx8vftX3
fyWfnDRq2uTZwiS2VCG5UBIeVTxe5Fajco46CJa0orQmSZJeVpTS0DB9vCjkSwQx
YGIwY43EfTRBqvkAv2Hw1U2JKYy1hrt4FYUZNvjehIsCdei3j4RmRZ9N5q5JGPy+
IXyRfBPui1nuYicAd68vxWIuS7Njff/vl9hbTfpKUPQ4kq4HSgN7Sqlua3NIFTqh
PCA+ow9UorZ2IUJeln8Fr2FhH8PqvkAkIIbNAxIFoA1HvcJGsBNM++BgfFjEhKjB
YjBF+D9F6puMp9AkPuKvUQfEX1H4RvGqetzHEjjNNxZDNuQAro7CwPxVE4LP0qwX
L8An9fZJyC99JIPsC/2EAXWZO18Le5DGGNCgid3kd1UTHJaaVL1hj0HPxWjWYXYg
5HfSUc/u4w+dHp4iVvI5R5aV6VtQc+4NjDkQVWWUuNwJIfJ6D6XKufNA/hBLP2Ql
ACLMl+Y7Il+iHRFNB7iiT+/PB7ZoMoT4VZ7s7qJ0Hp7AL9iKXRCJT7mdHfcS1eE2
m8LMzLvc+DmqzwHMmjr3kLctfs01h5yed3XOgPxtUhVmQ92zHGWURpTiAa3jABoy
8hZhDmwGM4QnGSInrmzCeZPs5iMgE0adzQzsT9fmxUuKrO5/LA12AtCJQnVCVCe7
u1qwPa3Fm6LIZWY+kDZE/KdV71kpZpvVNerpLR+WnJJtlB3tOoDk1EwMqazdrEqi
Tyl9Gy+gBT6Tc98LK8FYt3SdLZodsn1ntKbKQFQ9ZIiRrjLuglC1MmvUyhuzwj/t
OQq7DDhIISPgDm7bgN4pL7l4/QCJpa6UZDSMaRb/2zhoHmrDb6uf5eyV2946KtMa
xv46HdUD6M7SCvxH3s7knFw1OUFDMpTLecR72Lgc1C7mACtZOjGO8TPGjgmIXdbn
9oHfNlE+sSLrAm2fcEtRQKIlmgeWeEMAbwrLuO16EtuKYS5yUFagcYZbbOPiOzmE
+GCc/H8KZsyzy3405GYpv52pxb0YPPjMtVlIIGe7N+i64FEsERrVtFaTkYHhmxSC
Wv3GP8z8eA22keZraXzpRQ2Xa27bDex9pwhrhB+YSUCeUrixmlhdbVfFAivgwZD6
hIcmT2eYSAGtu/c0IPJpdPEs6GLRlmFAYgU6R9L73vZsUG6QVzX4ZaULN1TUjlKN
q/U8Z1oSlyVyYKdW9HD3kMpvKSC1HsZ4pu0XfQKux7X6MCjyfPTfgOKCcTHEHUnr
1qf4UMnWMddVX6JtJT//y586nq+j42avK+mn2sXsqBZfB+f9GYi6s6TRHqBb55BO
hsbc7akxOtvVBRtz9vT/XVP7Si81JG4vzaz9Dk3WPtmPnat5hK4t8f4i536QH+vH
nfQO7pyHa9kxZ3WBgxdk/QagzakkmA3I2PAwJiNrOIsU9Y0aRA4BG/NAlu6SaChQ
b3YTKxO19MODHMuuoTgVGNOijuP2RD/rqAydgMrcfUetHM9K1xOj6kQ31uPsF2Jp
xHk/CeW991LSX6FL/MihHU6cVuiEYQtaL++um3HPt1gP5WwikZtJvfxS3Rh86dn4
d2ayRjTOdqvKVHamR3f9hmFdDEPcOH4/kxV/lSkhC/ry7tLszTbrJ3KwuIpmIoxd
fwo3j0vsyQ4Fu+5F7qYPCrBBY6ToYaf3AihNirJwIexTtceWZjbi4HvDIJ0ixKXg
+UlTrwpDasOORHJ88N1hg3iH0H82QyEfzw4aBh8iACUKqZGUfv/pzLQ61ITHN5ci
DGYXU2Od2Ypfd6OtNaagMRKamoUVIa/YbOay8l28NMpIayl47cug4/Ni56jFgfbY
n1kRWH+Cl0z8e4dlTLWrLcC1RbafounfNhTtO2XASB5jMJH8q0tfpwdOEigQepCU
8ndnMntHUC5faEsDDudadA6bTIeVvcbfbwvH5zuOfWDuAc6mNoZ6kP4iTOn5ueb+
ddYzwmJh27B1H/IL9g0dnIE7zz+pO12/OWS/11U340031ymH1jmCDq7C9s9GcqYz
E7i/t3aVRTmSQ3HeGqvwmHOn+1r8Z3hn49QyGWaJ+FfVEMlzMdT3wemxciYvRyKO
sv9a+J+FggUsO+angNXbxzqyuliKZ1gjabWmAr31Tt2pHdCKHlv9LBkl1Iw7aC8O
jWOEjmLOzgjB/XCgp/j3kMDEj/nyzLbEAyuB8EgLJpcACZsP8ZBlq/rbDiyvkqUg
kQvjOQQyqqnvHbl5cXws2hJQKiBVrLcdOR62q/Am0JyCSQLJ/ZdHAJi0becKpIXX
Bo5zdTZxp+W6SZySkdz5eM7aQ7AJmAjVHGhJyXP++tmKmOGwPseLU7MBSkYI+UcQ
+22wbGEdT/H3dlXad3hcGivxt15NRJocFtNZxsq9Ie2semJoIlj3Q8VCe33vVQmL
XF+09VW5MwM1gVLGfNFNEAnAmSZaURjAyg/X5weNngqaAXDmDRK9d6YcfNXNmsAW
cVDuufZT916xORRAMwi49S2xP1pDQ4qK7u0LAtqnocIgFEllIEQCJZ1AjMsaEdMf
eRsnMt88ltN2BXPly/XT6iKqz14CnFhvq4i0xqsNsG+jnKn3eZC+yaJiX/wJE1Tp
c1WwvltC1QUsrsqrNsYZqRm3aLVzY9XpuQcq+78Xv6k0tdp+7y1vWZe+4fIeReI4
Jemia7dL03ZvR2C3yBcQ74chufs8iChhA5n6cHS8o70IB2SV4D0dM4BtXES5Yf9x
fP2SYN3zjRqtFVh3VPSoPEHnMcCNdBzGbfPaKygs8Gr/gfDRNsGg9D1bxJJOe/kW
1xx7+FMPLxx0+asc2WvCf+o4UCe9IuciPMf9Hd3S6J5J6gIVMecNIUb2mN/I6kHS
38DqUCP8+CxP80IvYt4cEh2EccEhUScS6Ta7a58ttcrduiDPpXiYVwsLrS3w/f4K
l+T2vHrdJSrqiju7jl9APFIb09ZmN8RQTn86YZFQNkbCIkoQqqu6OMWaTWC9NN4X
k0y3vmm9eAGZdV6NLiTrb0EoFETNPG/0FHCwRRLnj72K5EriK0mYh88FRxnaV4YE
HWh9UyZPhh80gnenX/VanYD/dM+mUBAMSr83VJeO54JAAQnawIVQ+wKdUuGZYJYX
T32U20IAniZItPDLLNCRgTPyTOdN8NjT6XVqGnT6hEPG48NuNrnUImXLNayEo9+g
IihOD9tWmjiYqZtenTUJfyrPVL0nT5EVJzPlzHRI9tshSmxNU+/pFaMRs8Avz69j
ApU0mZeZlZdOkg2woMdRB306TkIPadSvVLHwc/rO5IWXAMNKKdsTkQMWDLKTIub9
JO4icTgHdBuYRhRh0k2ywCMqr6OxJnTzCrECOTbOrGL2WN9Jld1LQA6osYObmmmZ
5nl6UYWN3xbvfwDdc5SWYWJDWIITiNu3wW7ts3B5fCNLoGH5ufFJ+H3QQeIGvBLk
pub4CjHkvsG+lx/w4KnohMyZXRv3xchU29VzxfiyaiQYl+rsRby/jBXIbwhP0SYr
EenNxyFMHU52bg67T9AiZTaL+vdSqMvR233qbTW3kVTM1q3PQBzjZIqF0fHsWjEu
+NH2wBXu/bp7pI5qkt+S37MBk4T86yBUIbG2yYtVPuABABFNB2t7BpbbiRTCacoC
9soD9dCJHOdW1cXmPcOAr459t+FhcYTT0hPg9TjD1Jf6dAe09SWAuZk/ugMQJqJA
zcl92k6uu5nQeCvmXjNt0jyi/bP7Djv7n669LGtlvBfZSBgldpoMa9reGljX/605
z9pzIu4mESuyaaVdvpOuodO576Ctwy2niG8jfrpPIttFGB7xtHfChggwi4Oi/fgG
ggR+y9xjNBSNM00hLS++/Ldx3XbDg02eNfJgqExbfuN7X8kesLi05K53oDpguqP8
SG7R/8HhyLUkXeZcpHCD4g2YB61gxorl3XD3i03ASvnl+c8XAV85BDr+l2fJ2bTw
DEa8mP3c/rgONY+5B2VNlosqGH2g4c4XCSgotPZh/BiGX8lvTsa3rog7hNaNpd91
/OwEoRRDGDO3OhF2vOCF7i5+U/31GEftcgeA3CZvXtxmixNTfMlrtK6au9gLBNov
Nx7Ld0M9a6Ap6ChAEQLLmGAPBHJOLmxCrAt+eh5O8hbBqblCahTvMUQ7SgsLREjp
RWHg8lwKStGqyH782Erdu5m1T7jPCDUFAE5t4eipQx87GnR7DNEystDvQya1VzE5
1qEIQU4VStketJ6e8mE1ZxLPWTizcoqalzd7+d/u6Bihf0oG5NpHXV4ZzbnH9w8r
iHxMWQoIsNsN6zzStBe+gJ9gchNHY+cE7DgLJlw/WBwkCAnqeMUYr55cp9BJb0fI
aS+6yhY0oGMHj7FaCZUE2eyhVrtJcoXQwqP1PHBbZ6wBTmkLJMODOL0pz3zOsmS1
UajUUSLO8yKoTfcdvYWSznxamGrEX9bw2TtmWZtwfg9l3P5PMqkSWW1voDuK8s2H
Hm1474mMQpG7z0F6MLwr4Op+eA4y15sSk6dYWhJ8hTwcVDYONnN/Oh9lptIKTgrr
nehVjOJ739OHSIc/QgYBYfteP+f7LUoyfn5dRbfzRTGfdv5Ds2Uu4D8zCcjV3WX2
HtyoyfScvkuCNVUYHHcuOeurK03kPzk2cdWqziCqEM4t3LloD82kI+zpsGjkHd+s
NKeAhLsLVDWOKSDRUjXsxQ0ZwQdcMghrE7eVYItmjmbyGt6hQjgzogZh3G+12CmI
Ds72FY8UhK8UxDV4Wj1BZN/01l+4Typh/AcAnIsL9kL68vPFNzExUEJLGwQ9AHC6
h8/iesPEeHV/brlu3BXBSCb6sAkcNLmQwzp6z8Y+irXmA8DjWVUg0CrwHQTtwfQE
P51j5tAAAAjF59b0Y1sJP2YnOfvuxrYsWt3cRdRJbrOspiFzdhXQIgHynDEZhQum
FTc6qjUyPofbmwPvcQbu4o2vjBg1esVa1OjAu7+8tTv9+O/FBwUh3Tu+i+avAujG
cX8IELO6sCpU4CrwxBvljAPVPlj1h+eIwM5MzNu5TvIhXe8i9QDOwOVWIRT/dzWp
e9in1Ro2Z65k6anwUYPFOIM2pQAOz9k2isGLyeqDzdglptiY7R/UqVJzPlOQQouC
AQvKFlY8Ydv03zNbR4NsSbnXvYrJGw1RsSo8/YP5yDE+qleFBD7sfjbwilzee8hO
71pNNzevpF4p2uP2drgsYP9ZRLPdPGhrNfmUv0cED+sbx7EmTQZnYsPTX5FNOB3k
eFx2TPRVMXH4FGsQHT3nrLZZxVQqaa214HFIC+SWpqmi/UY2DxQcTXGio1xkepEj
nf7GeCdisNWsjHbrnjLEBwP1vTn0cWP8560r2Ne3RlqsfIZ2cYhQ4V99PBuUB8B0
Em7c07TMqxrc2abINeO+SSEzVgtKdDMsJoznYbgEm/2Mc3ATV8ZaYVwibNxQyo7o
geHQQA/nnJFogN4rQUusKZx26yTtxUVo/qheLZU0Nj2oBb66Uuw5Hc2hV7o+1i4d
Tuuc13SLzcNxa3ru1aUOE5zjtvtBBmc4pfdkoXMAEVhQYg9/4TVvZ9zOWb2hx3el
cLTIqudOwKWymdn/s22BJkk+mZpAcP92UvZfUHhxLRPc0pCQ/vZNzIQMxNjMSz/U
/nj/fbs+hACCcqA3cY/cTskobuRoFMweNFcFCzSO2tNELYm01pWurg5Bbr1jzcjG
IzQSO5W6Z9Y4FZDknktf5Gxm1oMLBpWhxxJlZezBO7SdKRjQW6qfGIqznXR1bcKv
NNd2haZODiwqZsT+oJ4H1c21zI70x4fb+svlSIYYju+teC2JTLIBvgMNZWgA4x9/
i0uZOJ/dY+c9KZvVQof/ZS4zqWP694ABMvsrrv+lMQweUmc/6g9aUo2ULQc1H4/L
+bFcgmBHMr62QOjqYk4k1V2X4XPSeOl3vR6TXMabzeo3YL3vhYjSXuTUm7Wd1H6I
xFofKMP+twyr7USEbIoS+VGZqHfbRhX2QwpHgmYqVmthfAVk28KtUD2bD24xKp8X
jGAerwNGiF6InyRn73UCp7+U4LwHU47Hc4u32m+p0BI9OZZ0wX9HVyI5vqTF3Hoc
9/rBVaIFH9RuX1NVSlTsQ7w7nDFIn5ZsIH2D3yUO1SLWFBsG5TzZlhJ5PVWbCx2F
H10eyiKV6Rzu+UKjTkxaz0SoiPyFulq9dTOPrSOgQZoUhy0eE80VYKSxcmV8b7Gi
CrTzM/m5Bxfn3HapwrjByGW6gU7GulbLKnQSNuZT6U72+0astzza/CJKXqiTqO2p
TQ/jtZ1Dgzm5tUUUtbiDg6eS3SIqezSAAtdQyCCm4+NAbm9tHQp3u/zd/ssfqOjP
8aRiuMyBOyzLWdJcfCS8aBVTo1Z4FvKdW3b9jJav9LiLo/5rPJTfv7esDbZHmgGY
c1OmI8OTfc3HbayqmVqxkTWS17e6hsebhyv9KiWYHMzY/XfWSKtUAkPHLFuUWgUm
KGtVDWvinqOODCXtTqyRI9UWEgGVW44Am3a8tk3DQpOpWKqNTEvKggozt9xhYQDP
+A8dzHzdIfmaE8cOMkRPHtg7CO2/GntiI7LHLLfkBRMYd4klA7ea5WaYou5DKJTZ
y6FSwXTnw9fjkoDct6chzGsdzoPYpCnpTgfNpDlE92WvEKMOCa2knp4UwCnAsn2s
wCDNBDeVNlFx+4fRCDNPYV+FY2PIJc6cGxpdWEx7fI6YmgvAvIgslJLT/M+O2klx
w5+HGqDryguneYdssQy8UBKhd3tWEhQNS3SwLMGQyEg5A6Ru8OAxxFi5abA5h6cm
un86PQUVmKQ4a4hNWbVP1doDdmwbj8LieVhctSq6OgtF/kLZcfCiXmG5lUtyxIj9
Kn4kVDMLfgW5hBGtBV9dNz2dID4EJ0kjRqYB28BjyVjdUDFSv6rAx8YvZ7QIrXwz
3c9Osc6MxcnFdzgrql3nvnw7Jrl9hKyO3Xq7oU17465PXyy7iRnOipVXOSRcUcWW
6qJXn1A/ChLpcRv2l61CQql8ePXr+ARGscg6CmylD/2YpDnkYWhqG/6nxms5/IRM
DIt7ufFrDmV+st/sP/SVfK/JLUF0B3Xhf8oZRRBZycldcIHMWDbyORrmBYT2taPh
FsaTND9u1Bwn6o7ZueF33YPMHG3cPaxSOF6Qfubi0GSW9kU9pST6vkS1jiaB9tQy
Rude8ey/eIqe5lIdyV+N6VIRT9/CV3matVzMXLPENwatqUbVZAQJKV7GZzoJ1REg
2/eT2r6jjnlquVvFFIQZdWfnJdlZCoZ2yEGILboz9ycv9PHUm4KvfPd2iUY5i+B0
Xm+8jxPKRNRGK4znIvO4CEicW+e7bLt5UDQ9c+4V+wYgN7/6czQu1ygROmsudfwA
L5eLWIdLEB/3xzIB8D0fiQkG/wUBSDcWo3c3NosSrkAYguVqmnzMnmiYUJIsVnvg
sqhSsUf6f0zgq+9U0nDtcolOv374fqrRzTw3NICzY8dKVPz1OtZYtZAyKw1NwmWU
qTQklLewhuEbn9F5v7ZiYs6Ekn1lulAmDSQAAzQ02sBKH+YFiCGmwU71o+/+35hI
qbmsCEzCB6IaqCMEqm00VFjiDNLKmMWqI9eOm7wIDKUXwwV7PBOVTmGBz90Kh+fl
k05h3xA+ETTUAnGnkXAZRrg7lzKMdO4dvXsG3IWLbpm3mmjgzj6sCKneGqNsH49m
UD0554BKXNNzkkQ451T020blrgwqNNCzpBN12dLd99jnpa2XRZ83hq8NURgFnNeJ
7bigJPdsMCjlmYFSNZyAu5aJ7zg/PjjqqjXOyh0GSjpcd/NQmxZttnyMZsrKqNER
qeeJMQXy/OiVhxRdcHEMuWdD4EP63O23DINUYjqSMu3Ap/dqr+jTdRqD3kOuoNCN
Cc7AzAoIoF+g6bE6VHthMsPZEwt+DhVwUMzdVimKGjISI/++FBK7T46JWpJ4Os0e
6ds0VXpSXEiP7sx8D6TgGIVl1Gx4kc0iIKJnKtHwcYwwUjdUu7LXMwOwpfXXqVAK
Lr6iGGiUryKCZcyzPUB6mQ1F6e1htd5jIV4Y0/Dquv1A/qzYFi6jVUtAqLLBEI+d
j3hk8a/Z7iqAq4kmzhFyKrJZ6uU2zw4AyeuOooO4byqckJB2O3pIQ4sehPl1ei7Y
kS+Pqgbp+jefc+e3pTa7GHhM5TFDTtsWVGly21hfYy3qVp8UmDosP07/m75h3Ka8
s+LX1B06D3wry7yxcQhrB+g05ll4TLX8oq8cFajn4xPK3TBG35lP+B0w8sXdYA4w
+VXAZlTykKme+tVTPQKIHlKCREGPs291IE93CXPCqjUR9SPkN9LzIInLJI/RbJhw
f8Olgdc7itboRT/2mSSt1XqEnszdPZ2uV8BQM/KtQbJKeUu3vXtok3dZeege1851
0xwLzSw3dJvyu2glDYyRRYLH8WTnFaqPaoaBeaRcPnI+72JqwDk0nB3GPj/qBef9
B46GWUMaeg3luVc+jhJNqr6lpmIonFCSPX3UnNspPzv3Efq6CrmnYPobpZKtmYSo
k3odrGAiuwz0jtgyDYvPnf4y2aIYnoINVnscEPPf+6JrUFVNbfjHhLjhd4CvqYT3
d81phDEamSH7IjDbfp6w8n0+dL19yJI+j1+/DfNdJQsp/m7ri+aT2MUSjEHowReo
ln3h8Oz6xJyQpPIlPl0a8f87ePd4ghbuCJ+pAcEsOVcdZnfAODk96WTMi5bdGd5X
a33uh7/qUPuIU2MO1eqpXyzQWHDCY1pjKWHlsMJC5+CKnfNW1DC4/s5UKZrlD+2t
cGrKeNXu9uT5+yt078Omr/asHNatsLYgcapMPO9AoYDQ2ufhdGNSDqFJKfrKr4tS
Nz4zibcNsCB2RXhImC0l6BED74C8g7ZMKwX3Lmg2Q2xEAoAeRp1z7yOiobP2rTR+
Cgx/B/53eNI3KHDdunzSfjJCfUz68rm2VD/CbgMOzx8TClzSW82gGLEkvFYCV98m
eAaW7S/BotuRbCTTPw2FpzDrwJkD3RzZEnzRD7Mgpqmi4CQhFBarwspUjT8Se17k
4NqRVweS3PnghCL//L837/GrfYS8oQCX+8JKgjanE9ACGfQzNNNcTbnXg4JnPTLf
eQwUCarLBfGCr+86IvQm4fZOyS4puSE9RBqbMkER4OsIit14jKavsc3zKJO+xPSo
PJgO9I9c13sYsXiCfSGwFeg46PU6aNswXUp5wrU3mviTdMzffWLz4F3BMD7jKHPe
BKlvNZ8IpIM9ZTXk3PvjIV8REmK4AyrTiUGCACOhSR46WMiX725ootRf8c0h2fHS
4mMOWZhbg5/HUaIGnZTLv5l6DHYPNeWuXMCd4zPeGX0yrbDtoDY/SvTTeH0F8dnW
RXr72mkLg695RYZjXPWj7tsXWcYoKrhXIWsdVCJpIKWjgM7N4/hX6yIPONcQpRq4
lKBTiOro/31CEPf+DG7G76L0bmxzogi6i2+WTDWfpQHuDKf/r9L/e0sfi2lWE2wo
B6x4ZWoLgq74LJOLK20W78pSOekZF6EXQtqpSIbcY3nuSGhYmyF7Nxunx9xk/jmh
cCYRHOL8QoVf4OVeXZD+qNlApVqKM8fZHBQUyd9ZnxR26skJtM26v10vdE818/IY
WFnYKELhpZCO7EpmOvCLRewh0rAfjuJSLiGH0HG0TlgtKq2LU3enZEtXfoxSUQ8Q
zqIya1O9Cv5bk/tG+DBCD7rLi5noNnPdhxaJ4pTyIWpvBEeSIhDnlKPCfdKBxSVA
XppRB0kll3X45etnfXsSW/iS6qJdSd9ORGKdMK4i1fhZY/1z/bLJddDrAirZN/Sm
Ap7x6dscCMw+76Mv+5oT2kXxu6geKoCiIxk8W0gBowiOn5vBzIbAU+Ing2hZim8U
NDBoDChB6c2intxoc/K0AU1WHA1eGTQGQY6STQ+OBP8avXUZjFpH+9VnzKpk34XI
h23nrLwyQdaoJT7ADvGNBCl1mDj6yaR16cjPfBGlsYKRHDSA2HETPvyXrH8R4WS3
sEZKgo9DuG7czWtrqhVuu/4lXYB6OluEZi34U4qNB+wYQ178Bw1WtMNx9geXOeC0
u/ok2op0aMjl4n4oum3u9O/+2msLbMLA5wG7sE+KbXntB//3yBT8TDQoEZ5cHpBn
VTumb0J8D0fy1uqVkIqQ1P0N6Hk1+LC+wSQyQx78IGzKIx6YixHEMmKJyU7WZz2m
tZE7NxDNDRoCCHRwmXqeDQcJcVA/wu2pnSZ3m2AhMLnwGuFTYpuumZKXlUdAsBJn
oBuSTDXUImFyZ4MepJ4DQcNp6QBILP+0soi2HF8BX+MSRl+vsFHoWyQCpMRvGH6q
CItMQYLOl9FPpSu2IrJw9wJxS61IEA6+4XIrShvglFhOI2Ux8dQ5iU9OPlVJwII4
o9sqgKJo9TlOhp+p8V9I2JmVOj7YDsCJucMVwbANfkRUADw96vU2zGkGGiCO6bph
N23K+qNFlgZdoF8DKHIdcQy+eBRMplyvSBCx7mpsfq5swBEXqw1DKr6OJuO4NXIi
96VH1GEFeu8RJqklBjadYT0P1qQLe1zMyR1dQwa4Cdf1bAiClgVOxrpoaLj1Aycn
C5bvXTsKmbJ0+mCxJMd7zB5bHOwLu8v62GziQw2liNHW7DwDWkJv7oWTzO9wFl62
YldRvZz0GIytK5bDb032fYwOgz0QcLtiwDLNFA1QchpWp+QcRjZb6tekIDVSeHcK
l66888PY/wedaiq7aehP6idoN/A9M6otkjog9bt0cPy/L8esyS8FCtzQ0uobE6C4
Q6sDCJSy001yjlOlmJSbjgdaXf3XO1U7JcdCCzxbP8niuTtd810dH0e4BXAJhh1+
jbO/uH/APS+aBefR0rqREmxZ1quST/wH+VWi0WWSVNgnx1mUWfohh7xOcDo6vKrI
pPaJKxvQ+9imX6XaSfSjKSBe3dx9JLtwK6k/bUkj3TNuw0W2oX1B+kcfY++VWwLO
vB3p77qiZ3+ZE87dvEzXi060tJ+QBcttyNFSeU96DF0i3jP8RhdNZI/zNHr16B4V
ZdFXUvV8Kd+izXp5KPyzT+5udP027V6B9nQ7C5NIgj5hz5X+fj/V4WxJkc0p52X0
0xTpQhbTGg5Z+WAcTikTqurLO/GhkLIEB8DvgeAGHkGlG1M6rYRr//WKEXXTG73s
GwdDsJ0C22jCuM+q+6UMP8OphYAFhi8jeFBH/+ZxJGCIerALd9d326lw9P7re7IA
t5DLPY/SFMYjIb/RTKVVOebjtBpfcej1BZGRATszACdL5+Wpv5Yj40Zy/fjUg7ew
KYLziIqDD3fnLpD6gIJv0ftKgKxUld8jf2OLPlK41cnbAYFcZWHgs1SllRBoFsUp
BjppdcehuWyn5SIOcAMgJMZXk15nC7FYWesBZk5+R8grHeiybIkbw+XNVQOvqdTt
p9sJBe2c3jOKUe/VVqVFEkB4MCdid6C9hHj3XlzwQofURBAoLqXzyI7imrydC0ok
JZur6g76JezdHMa1zCIu7ISwD7tw52iYlBrYJC+OFElFkC/6weCjZB435DiHDTx4
PTFG8zaLw5hPjeBBb/0L+hZtwHooNuUzmH0JGRzrSH5DRzONUoG5FlD4CO4tQt6T
hOfT6y/VbL1CGWqgl5TWU87ASbvB21iFf4JrCsnlau208J1u4uxyHMm8pzrQLkQE
JGn7uW4VZu8hkWeV1CYWWbzO5n4ewi3rUgZEbj+pO3xa+pSZrakLPGGSWTc5h87B
cWYMe9G3GYQOUKYCTTKuzHU2OeB5rIdAUNiwjNybakftWPp7zzootx+CMJlNwzo5
36m5qy4P8SAS28xGUIH7dM7AC1Gg0/ym+x7iTVkB/3L8JHUAGkK5SPawumhfs6wE
awXK2l4KTfJ1KXuEdthpypUpe5DnvLjfmxilAhTjh8KCI9+3FwMXaKA35EfFEp51
jmn5HXy8TYIKH+FFfjNzuyvLSXHzYiGUWMCFGJ55aMjMqU4egVasYqIukNgPyUle
juuY/fhXpt6bA1WDhnpD7FW4EI/Dfpj6tlgh5aUklt7AC1guneS8eCMZjMx/JkcB
qw4NpilT+uwDiYqCYA4GmTrGnnsN7sX1PshTFLrA5z1hR9jG3aMakrhKwFg5cQUF
bJ9yEqEzOo4DqLgE3lhCU9jPo//Qd/RTTJnWqCpoEXzTTTUBHP7Loi3epjJIbF3s
vVj46tTrHhJKSEhbBaojf4QY+jDFBKrLHbDs2rPQLmsS/iLIeUR7oZ4tCv0Ft+69
BL0bQcGSceqWzolUkcF+RayftCjov9Miqax4+fw2yqjtC0jeHo/k3xR1pzRsMM1K
bAs95HKNHTYDkEJ/a6dcLYgsk7iS/KMnq7ncrJ3ojD6Zuf0yFELq7UM/2/sqtKGk
0nDVmf7BjuqXZYecprB4AphciC6T3Gv+EFikWJUJItWbEKS5RyKu5Q3l1up0k2t7
WauEypHeSFwJcXNnEu2ouSyRVcqo+3tMg07lkPal9VPPXKGVvRA622MTIkDIE/Fo
TNM1Zq6QKaesjAPIXem+4LynavrdwCUUQM27PFEzNupPjn1kA4nkP+bv53p9fQd/
p4iE4qiR79YSZWscAeCwGmtlEi+5loU2W0uaDsSaI37RaKr85JpY6veCHWMO7vPc
74HbDu7TctObEJms8Ptda85FebXaO9RNpxA5yY6IjsB+GrZiDgvpzwkm37urLHCk
OaPDxj+oGsEZVNFexq92/SfoZFkplh/88NXh03fCe1N8m3oFlezPytb+HQhHIRht
KPMzC3fuSP+LuTVDkE947QoD3VBq4HgWThMYv+LY5BkCl8Jt+g5Q/lgK81yECOTA
sXgCCZZ84pax0YUo42TsSIXbRx4bKCDhFlcQsjOe2Ihdy6G1Fs4VF3n2NzyJ2+1k
X1t+0fAG6XhbXqYKMTS/NISDhZqhOqugH4MwgCx/PULyJJaXzROgICbXwzktZ/e+
B6155Vf8PfxoVPysEeDpT1tud3kaGz1X/8N88yoPLLyASr7gYYbBiWjILSVHRK0z
qda7671nCvl42/6u/1ZJnSBB0qPeRnhLqk/nz9ZLbUk71s2e+t085eDYz5gOMUEg
9f/3eyeMexF6uI3uEPb0Wuo0gxIlcFrF7EttWu752mO8koVryTmvlPvtrJJluPCE
twXTdj+ySEA0N1j6KISpztHWPyo7GGTvhqFTy9zj7MsL96XKYyhmBreUfc9wNaIz
xofYM/xcrhAII/Fhi8j9AcgGOFmDuOsmDyt8E1RtuRC+7BFAT1Gk+W1wy8BcAq/E
B0FTb5n3gHuHhcA6+f8p+rG53/9hb9gfeppnq1dULId6/639zaTjeh60LcB4VbBN
PdsSwq45zo8bMV0/xeTeANwMxAkhacOo9+plPS4evMmZuQVAsWHu1HTMrOZdHelY
5jX8gdJL+4skuDNEWgy6L2jRZzv0CmpCNTHsotcBEUl+2PzMODKxwFvOa4OtQyh+
xy6DRNyuRVISvaKXtUsgqb3YhDzPbjelOdpIphmRCx0mBTxZwWGcuBTqlpLwp+2n
nfm4R5vZTMEwOggnPWPKbnXJH7stCxOyHR3AS6v1ztsTJc+/xd85vn9ss5Jbdwe+
7jig08RDjeQfco564YcR46UmBayfDD7B/ipQFSnL7wgSQig698vmBf41oN/gaRrn
PNo4AWVzRHL6g+wvwJepCMHHJn+l6DRY8CpCInrzyFIDSW61Ilv5bWKGQiz1gju9
K1s+Gku3YpQxew7J6qAPwX3wgy9VBbNgck30tUjq6PpdAF7vmO7awadFPDfTAlIF
swNh4nODQbxeprCe33MDUcNdJRTTsMtvzfivihQuEMa1NV14FcGLJ+BwLMIjUzGy
ck8ms+BjaAtlLTVAjOvcn2OegBF9Qeq3hS3zQHIcONT4je7g0vmFNI4g5BOCt2cR
4o/4MZVUldNW2ZdObtaaPxRC/C5h6V1k8F5JQU0HXrsN8PUTDK08mgE+YaGe2DYW
rHoETWPdUA0IC0yMsVTHtf+GDmCBn3jpwAMfDjKjevBPpc4AHabCs5+KeIKqt+El
vBSmR8tgpBzbZkm04HGzDvU+Sl+i/RKRrW10Q4MWNm5zMZgyTOloT+dPeWQU57b0
b9IH09D2jF5wdRN+cYuaNaeyuFLdTUsnxLOvV/CQObeOwKc+7GVlHz9pHMBH6jaD
d/FJ9weaxJp3li9Ibw1wrfQCX/LlmqyRaOj9Iv+nOBLZER4S6rWqIehEqZVAsgOA
hYV+3/NxZHUXg0Ur+Z9scvmJKKaG2usqJdvJdFh2XEST+gyLXPmPVX9UWfLBaxyw
tlUYlz25Bsn8PYAstLilIpE9jTfNDJh12ffd3dRXmcLssv47i+E2BIfw68J1geSF
7+3RALR24qEiHetB94SsbHSRGriOdJP9tFneq43AmhQIIaZjDvQOXaXEkkoYG1Ly
Cog1oSf89dj6qKugmalv90oXMdvzLT78KFlVgVBwY69BowfOHcmDYXeBniOrnztn
styTMPzsi81qMWqAKNpjMw4t4AMskZJj/JESlJiyHDKZY5ksB9T6T5PI/L4EHxUH
QM+1WIK1z0kStJ3Sg092H8FdCOLaKsohXO/hcoPLkDyghKy0jBNwsbHLcW+lzRr4
ogp/I+B9oR/+oEv3bG8VOG8tqwde0Q81NnyV9po34+fSeZX1re7pvUF7bbXzRovU
x/ZcKna4/m+zePMQAVk7qw7oXHua3YSX/O5/V2mMhPBIPnbz98OCJAOvFP+XJdLV
/HGlTCuJmDiPJOxnod2w4Z/74pMtrvVHj3YKZHQnohu5thtHKvppyRBGBXd2BaqC
cWyYUFuW9qorfPD5oJRVfrLXZmc9XQ+rWRk8PX26W3rS2oecz8eDii0zJ3IBJIMt
QXxunEgwAlTO40gHe/F8vT+/8snmReXuRu8IaTIgztEg5sZuN8PJXp2KEQa53+L1
kAWAXt7xDo52SQ9JnZWMqDpx8H9On9Nb/dki1eDjmBnWLfeTvhwgT47qzJxGrKxJ
tDRxcmYlzz7C//bCj4Q/MmmFzvzYfZXhioybPOfLCmOms4jz/BRt6HVx15qZxy8C
NUjMlxzEKCAmT3V2KCyMqmqu0SFTX5paHhPBQEawJpqiWCtbMnw6FNs0Sr7HQeME
mbfw70Q5uNzDjWF+e/Orw3R/latP3Z/8lQ64VQkSdxkGaa1EkcSWL6PIJJgU7W/l
SA3mbbLkbHayBqw9CcUQocXMz/L6dO5rrG/J7lW/1LYGpQR0oKnH6dT9BqUEmfTc
GWhS8sKYVJbgWBSqejSuMP8eJR9zZjmoEw5YDZH/IaF3JvjBkPC1/+4io2nkkNw8
aqu3FpvPuEa+jITkxx8RyYU1WhyUxho+fNUiHfr3srvtdx3eZfSfmSekUqUM851O
QfUfq5Ppv9gMEK1CM5vzSQl60g2yMfyljKD8BGU+ZRb2tQQIQ8wfHsUY9JnENg5G
3IzPOsRV9MbMHekOgtO5eLfuNtWPUi+H/+Gfv8BTCwvXD21EM/sEUFuGHhff1H2d
66lx71uuZ1/Lqi3RfKvhYPihRf1PG1BIDRTVNH0ZIWrbdlTFwPFjl9ZwH5/9ypyW
yHpmkOqKUWLm8ivbEV6QhxNtEwYdWPyF/JfzQN/5UnrcGOBHyR21WUkdlUjv7J2t
DJhsVST4Kl9OcMBKWJIcbbfjgFKLxOrQUP02Fd77/6m93zy1kRCc5NApVmwpmGGA
Kcrz80HrdngvU+ZtCbR+mUWoWP7g6z35CDDC5333pBvmCm69aoQNBCLZ2PbIhFsQ
d6Y2aUBOv6CpucyaLPqOllYDop43eZHGfaWiYox4oEQjpCLH1xxFzuz6RadrATE3
syaq+w+3ffEE8ZJ6RL2VbAa+ifOm2WwJ+Kb7AHGaW7vB8GIYn9FomwVZt76uUgdR
EjRouJNjzVTwcfFF17972Hz9fqvkacu6+UOAHD7A8utdJNvppAJjD4kdwMPKpaqS
klk6g1qj51ChFOiG4cvadCGeVVY2FrVzsvbbO0UkBqGlYs1KPfYYqPBxWaAk5Qgr
fUweELShuXM9JaojTXxQZBYQAYTkPO/1XpjjG759eHl/GAfR5Sq9DRclT97GWJJg
RAbiIJdeq4OJoeCFgnFRbC7OaMAHZK+F8R+0HOeEa90yTHv8cBKjN4E+qjBsrF0j
009Ykss2Kqu6itwEMqYrC4JLcYQ70Q1k3zDnmEvtqI4q2MTXw4mH0uraSRfoWYBd
IavP/BZzWNX5WNlKWnsZNqcnqdS/sxSTheXX2s6j5w2RrtsQ9h61CQ7Y35VTSy0C
uSS6k5OSvAdkE5lk33gCKBoTu5LlRCjYmVaCnEx/ytxPP3lAsVo5ji+Thkd32U0b
9m17nu+BfIPWW7zF1vNVL82220mRud5KqKBIYeWTYECB4zA4IMEGyAQlcfN016jQ
IfUfzYSDlYYyqygkNZQLr66Ixh1TcDJgNWABDr1lXm7mhwuxfMKywGoWudqojDpV
EgYbKSKfGWCSxe4ghEWENPQ+sE7l7+yaiDEZHCX5n5rMLTk1hnXvvn97sa1h54fu
Soy3Rh4Fq9J0aXE1XXruBWRmujSVjoUFJN+TQffDPPzSecvq420uLpCUF/PnaW/u
/45QPZugk/DHKw/tTmuvA5HKh7Pu+e0dW/oleSUu6Yrrd7tQ8NOH66GcJCxxAe3c
kRCdJl4HmUNJn7sgNLEu/1SuS/nSB1/unWfOk3GHK3lxFQbNOjTJnhMJp6O3qG6w
piLPCS0vkJArbDkRWPI1FmqjMvHqW6497msfzovaye6z6lYBL8UFW31V9qANRmcB
+8z1yPsgLFqiEzWH9p01RLo0y+BCcWOy+08up2D6Q+PEXOOo0n2cavZq3Y3qwqDu
/eeRWvYxpztByDoLphQmrTzceLzdtPSO5DI7/YOUKtB1tDW6YvPZ0PWOIoUzhZgt
wVq+G4wRyCtBZYw74qa57Kheu9uq5hpsOp3IB9nlPrSXQbCoIIi/6ijJV/uYZNtg
mfKnWa6N6bK/tWdt9ke2vYK4g8IFIde+Dg/2hmXKMM/AxAPhz6fY2H8lbrig4tXU
nQLcoYfBPTgsgroOA1acs5Tuv2PrYozIKy7Zha1ZR5oYeDUDa3a8/mjjFWSX82El
Recpgu8CvEzN9cZS7kWZpPBFB4ApUPUigOjrx0G/DoaEaVKyeJA54/zwlaYDg8uo
gDdgLYPhZPTNiYTotvaLXJplTqvDbgb/dxmLto+ti0Pr8UmhQIGRL/wgFw+urCof
aCj4r+kzJuN0X+MCVsDknRxAVS6fBRLC4gZWvBwFrhNRGUP319kzigoBJDIbrHpI
grvSlRhFXgYIF9RlxVqFCTl4SNPC+c0pwbe4aZ05aBzDHWBht2bqsQ/efUjfPAwa
GrHsZlr9MjMg+/nAPgeiA5uLN1HW84jMb6nsvqYXyULPRIMzDoHEGtcGa9rozmK2
Jj7yjvCucIcTuloH26wqvrfRzfkKPEZfmrUWSoQ5cOqTKOsiYDF3k9Byt7pkGbQX
Rhipkjdt0gylo0zmRCim0NoQckPBUvBmJeeT6+6iJabG7IZcj9Q+YkRhfu2QzPIW
RB4nKK4+tYSydijWDewc9jR4HZ8YTa2aJirYu9FaOaBYQT8Vkw8dvopPVc+ZrjzI
U8s3QhuB+hSVObKsr5jwEMCqEc5zuA0vENF8dMcCX7KVTN8c4TVgRfm0D+lD+0IX
PtNNVJPpVKVe/s+HMlLG9s6MP47/6hAlDFtiZnl4/68hRy9eEPs0/KxzYWlHNbw1
+SQPsr+/uI74uZYROOWD7n4tmo4j9ii/xP7NLGJCnPBoO2Pz+GqH4pxG45F8Vav2
IE+f0SMdbSRnYErlCwADgK0ulMQBrH5oX0zVJxVO5Gnp3rYKoe0FLHKRGQ/Fsti9
pvIhrf6Mu/0JFSVbrtAPyaDycBu+5nPdDSd70ugZ8bfL++MucRWoJwk5Kbibzk1f
LzcE4sjMtFEWX65cHKiPSqtig7gxMztlRUHFVIPNjO74TTlTEGjxnZLCF98h23gp
kfGXfHLJcMZ2ASEbQGDUnEbEd2Lwfx4b4m+FldccRRJgCHtOv7ZnZwTkEwEFMN0V
TuEUOMcHnNACxsjMXCq6QBq3NrQbdQ2qGb9e742oDB8BgqKiJWZKPV5GZgbkXW5p
FOjCccceA0zBtIRZ9S4dRRrIqchzSWf4FCRLcRV4tIUp9Fe0ChFa/0UAtK3j53CH
cqTX2xmurzuaM5dOskkVNxjMiSkBhDN7ZTG4n8FsIF4x9ds7NpWJxVt+WiEeSUgy
2PS3bIseZBLxSpxO9e35RP1okaCfDZi9Fv0QCnM7lZ41RwwqsktMcYTN2adLQX2O
gV+fHDh9T/ORQ8+5tyclL82t8eOyXRaQJV0Hyck2wzwJZmuVx2UIwWD05qnZ7Wsa
PUU6Ja6JtY/XkWSv0S+8tot+tfyhI1YgNRRgwIDqpYT7Hgg4od1ZgGKcW7CDJ0TQ
apsBqqbKIfyycfAOMS8IgTqfrK9lA9nTwUIJ95UVTKZlfDdKbCI8bivVxKSp4pH/
/Ijao3u1IcLL4/DU9CFggKyvpjC0GGbB9y4UmJgX9q7tz9PVRxcJty+esx7W1F8d
/cOG1XEaK0tCYEZTrCql6CRfL7J4L1SMYWP233UfW6Ikrej4WgLMhlaV7pA3HYmb
ybF/YvL5nnEyY2A862syz/p33h0vDEaqSZnZaXTvyoAAICREZFV+GFeyv8aoy75M
/U3QldATi5gmIeCKi1qT4ESsSx7kPJTp0Ufzob5v5XuPL/CiGObyC9gLgWpeZtHG
N02G8QWT2llh6l0KtQ8+7RzPD6i0WGKv5v1lCvwqM7rc8EIL962ocCEFThRqbCF3
8PjjH0rd0r7xEh7ymGsfUR3tvX3dRuT6km8DVBqfElzGK+IU3fDTeUdweUgEF+RB
ADFIMwpl6c8gCE06vPh9jBeEHIFi79Y8Ssh4vE3RwvNJXca3Ze3dT31NGdhrc58k
sbLvtKnYOz1L1WZUWRWgmGMHt5SVRiBGj8BWqk81YsLOrtYYEdZs6J1/tpb5Q1uJ
IrGOnLce0o/SdH7sgntIvySLhGXmuJn4j48GnEHJTDCsvSrhpvX2V6Y12HcjdCar
FoN0M4AnnaLu6u0E7ziCRCKtNsxr7BOpoNPN6KjCNpgvAushhNzqcH490GjxZF0H
mtqBzPmftZJ3dv7JX2c0H/6DGPaBrT1VNRtzQMcAFCdrxuNxmiPZvo6vpCN9mwRa
1dH+FQzlp8iFPfWoZ1CJoZ1k+yyAMDgWrUcKWbfDaZu1dbu1czRBZkFo8WE8BJNk
dF8NUwN/JEKeAvRvvqCZh+OOIED1nypdRlREGpkAKaejp1vVOH1R3KFNkauYAm1U
4GCuudU4pwLeUy4OCeiKaRBTHq8IFbQSxBC0LwIYuO12dZfqfLeYwnR/SDpwiG3u
bGfRj6jTlloxFrPnXE58hOcXVfJZis820/j95bXfUfimyqYeXLchq487jYF9pB/+
sqKM8Fz68/n5S9ye4H9CMwqfl+DPEHI1jZUpX71vJug4BlB59mhugjfYTaAW1RPv
0eWVgHYmb78YFXIgl9Wl0IEXUmB5m2WWXLpGsThiiInvALIAtaSGInBWnov1UNzy
p9gCMr55rxJEMJoA3j669+2Er0lG8h7AoJ2Vh6XuFJJlGcaVlmSuR6zUWjqCTSN7
1OgyE2zj9LRbs53+jokyV69+iw8zShyPezrDs/2w3gbwL7HVPPi5AxdRawVMBwYQ
Lh9l/UQW07f7MEkTT+UflCu3+umj788zwDiRc5zf1FftG2bmwNdoFNfgbhwhKZIc
ywozitjEu+Lz3dlbRCNCe75/eVOBvlLdTT5Ka/e1kOr2Y/X+zdhNRgug67763maT
5FBgDD5qGQCHI9JyFZpXnC/U/Bk1u0F0c46z41U+2Vlu6aZtN7Nor1Y3KVyuTCJJ
4a1koimnmYwQEvUD9CnjGW74L/NSDpMyywl+zwJigsixtDIWyGrAPaDPe26DpaH9
06kUJMIqsf81AkXF4YhzGzd9TZ3WSqHCXJlp0Ww/NXzSbtKznW74KX6bJP484Wh3
ONpgmzW5nb/e8RpOOaFXOsxn790DaZUjyUMAwstjeERIQNRAxQ66csUEQ9Q4LYOF
ReuFenKswqLTS8DkB605NNxpzZrQQoQFirEKe9VgpJ4OLxtspgEoftFBjwpl0/S7
NjyOz7CP6sEfKxcN2vUXLYM4NdmfhtoEgswTqtU+EAuVp9EA4y7EWkeUBwk5qVUe
+DFO+dPop6g+cb8tIcvKLcb3DBbDXdK7i3sjL6N8+PDq7LKWrVxR7/Lf6mRx/GUd
eQCTqpmiNnby+MoShvowuCNWV+caOvkBgRihxpgJ/4BjOnfpCkr3aZWM5nlSvjs4
3XU6Wm2I8aeLDE1ySgXrT9f7Zrzm9uIZeDQZSR+UNjgRhVnPtrbyyqnzh95ITctL
xg0jS/epY+Wf9bwg+7DSJcE1btMsThYbOWMmV/V75iRhfLbaBo3ACumyBPATduLn
fwx6hjtFQwuEaiwFnVGFaMvxoZic6wx6jOUF9zEZ5+90hFt5uGBZPXI6jh5hhlSP
gHjIkHi0YcEIjKqoTe+akEVHYzYQ+Twj5mXtjCX3FWaaaLVVcv8DI8QKb1Up0/ON
Tudkm646XMXa0urshOBNAUVw/t6dSZd7XsjWz/Hr/rdMCEAfLHlhk04jcU3+/x07
Ww2RNwG1HliA0nMGoNvnPkyUnDxbAaQ/M+sl2hGk8URwLHi4f4pCWaA3dVqUGlPv
lc7gJ7jOjp6j45/IR5HuGJfbEDkSuZ9AapnAWAEQXNdCqiGu61w38lsNU+BYombW
b/yrrEpU2xuMkwUQXTMVvsqTa8JKvawtyXe5uyeAHWQpAh6gqwBuiVbYLEe+UFdT
tGf422pC/VvqKzov1E/ZO9QCvIc31KjO6vP9xhZeZebimnLDte4odtLPtOIb1jv+
yDbqbH9Xkb+7z6cmqGZtnI0SdSXUoXBUakocZ4ygca+ITBKzMt5wiEQIW9hBZw/2
G5mcqL3fP6c3g5ewqV19yS4kuvo1VRykneMHL7j6ztuNxg4EsAy/2rdP1ey0ua52
XhdgjcJmiwKjYbJSJK6SHUTXssWQuy69PKAPOE7oTJAlWqNrvQKk6N+ZqBfGk/Lb
g4sq4loa59+KYq68TNiq6PNlMOMYspUk732s3k9Tc5yP9wUeUnw2E/+vn5Vlm7w9
KmKzgsbliVlkuYRwvXOmqfo6HdYcDDnuL6nVWliDQSo3Uj4OrU4lRicMIyuiUbL9
Lq/FtNM2DiKyziGMCVBiUbZUQF/5ESMkJ6g0GwwyTmFAIpUGsf/n92XqpgUsh3LK
NIvMg0szR1yXXkbrh9APZjM2c226+4Bi5Wv/mhdSa/s4rVE6Eo0xGcbeeyOOj39c
2JVDCoOLLcomBvRcqldxrXq9jBMGtQYpvbjuX5vHjQteTRpf2Wx6sNJOXe5Th/5e
0bA4PGPxbAINEC27Rns2DAEU8ozyw7NA/aqEMgfPomyWSmXFiGQN1k5XjfVdX8Tn
BpCGe5CvgniF/DKJ9xFfhtdm+8tKL99Fm1hyM39HSIPGAGowjfsP+To/jyf/CirZ
VKkG9UhfuKABxazFV/i2jxL1uyjYZPwNN7cF44b4BCl+2ozJ2qcn3fK0+GtK+vbB
rYNeKWCPnJYJQz8LVmpdNetkzkIwIq1A8bEkmx7Z2nzufGv5Fh3jm0SB+a8Oz7mO
+wtPFHf5aggALxkL18RykTqJjpd8zokLjB0tznsXn/CRToNHOMimTobc+MRQzM3S
jw7WprId9WFFvC+N/LOioFOOWiCoMVhkm8TUyptwiaErQSkNoAmKlPywTMsTWf7r
q3bMFQdrURYo9qqxIwlXO8RC9T5bvJez7O6SqEjmi8xMaNyaQkZh3TDDwx3RS2KJ
JHh/oLnwCzx7lTlqV/va0TE9rCdnIQwqhzOdFshzy13uVRDg8zk+QSvPX/FADnJl
lScRGK6unLcai/pPhlRlzo52KUa7db9TZdnk1FCGEm7e3buwYbvCMHdbauTK0DoK
DS7fppgzEkNzCgWwnZs+spxWtgZbD9EQaaegUCqu4tSptn7hbD00RtNlBGQaxTUV
8oektapwHLhyUiTTsjRFN1qgz5LBya7MfhxbpRQcKhwnLCgjnMItPYTgu+AWO67O
M51B1YEtur3Ycq2kRjGkP14ZmcgIWruvIW5fvIYhSUJ68plZQAhPBCage5zWqDr1
5wb3TDHFYQJk+w8zb9xfuJA7acFBhn5u5pu+VA+CXKmdUSncJ11tQwp9IkFZwpCQ
2gPPuglq7PXJz6jYhphglREh/YkyFKKIbG807mBwt/h4mimzEMFo4ryqPSJ8Tpsj
Lck/iCvbZprDjVsTFOc/gPKo6vdD3taHJan2mofKpetAq7Fgy3iL/PbWQ4f4kNbv
PM691nJJv1mJY3b5CKJh0ClMXf/zMs9VVJs+1Yo9ipsI13w8Ro9dHi92sXNKuLN0
XJI9C6ShBp1VNgfRkcLrzspVO9dIiL4Lf0sjSArP4qozUZRlQlCHSbq/UG0VptJM
BLgYss+b6d+sq3p57TcuckXrKAiaTCi+dEvInTPgCxUINtIlRJtUd790m5R1p6Dc
HghCILLU2dgMV/xbYlixLYg+UiQt1MErvXqcN9clCuNcjflOvaSLsH5PSeQyxw1Y
XfL/FiWW6HJa4SuCV3tgyVN5dHIyLZEdgSNNv+73DGbe0YRkYMy/1cjWibqkE03N
bF4wPrijhp7gSF31iKKznC+OPXi8qMcY+kTxNocPHYAtQDWbKgMYkGSXfhD8Mb+l
5lx7/4h6Fc2kbojb3g2CNT5tjMJrLxxGR2ihhHz5Cwao9xR/bSok1iNzLY0moBc9
RKN1JNA3vRYJxxgdEwPyuRCrZBHJznIhY+Eacf3SESigKi8HQFbu/vaHbQNz2jDx
qdpLDb2K+27OwBiA9h1GAnrQJB1nt9OxcPSz6+RvntixZtQE2WD01EPyfojgstIs
5xlr3ih+q0xKuX/S5W/d6QyR9uL0gBxXFwZA2Wm5L9bRuxwJmK4inb4YEpsXNmz1
w2Ejvy4w5kGD8N+A1HrFwUJWVPcWrdEGugwXc9zLxP186Nil0hgVPOoxgxdvoQnt
Cp9xinYONqCXemYQtdquk3GVeqPYo/LUmUGlhUbPJ7orEA9a3e4jkaG0sc+t+3e2
vlo1ImvqJCpDrEc6E6ntiE+MWzic6lI2h5CIl+owYOdIEPSTWsrO/CdXFcW89IPZ
odxj9yCaiJRhxhthAW1axwpSi6qm6bqu+B8P9DXJ9yime+qoWtjerUofScNz8F1Y
MfBufZSoR7QnUdLKvqDpgvkqzX9ydCY3QeNYh7frTNPTtRuBBhLo2s9xtIeJksMF
IMTwZmmHMEfw4WZ0Qsu7D8wq9m3zR3ISZcxoOpr/J6qC+bJhZehqu479HLXCdajl
WVTby2QuA0fb46znLnTMgzk6TzdTHZFwAB8pJ/ukRErZcMA57Xb7P7CrRqQ+qYwD
ZZUmSvsOnQUK0FOLFbY+tfJm6RQYV3NcE0K87XrkQSXjcPcOkP050P5pDT+sZNMO
ls70QP/1g0o2Cf5jp3whZKrsfJryH1g6SYtHlMVjszv+DCuU0a8ZdLNjUuiOfCc6
2zTzI0+3R1MZ1tM+UxOk4bVJMpZLrNiSFMKmbkvdKuZeLzqMBMhM2/i9geifPmhm
jBxOKaBKcvttoUTU2vMzG8V7vpHe8cL+i+4OY8RQvfOZzOa4333F2rDCx//KUI3/
SuOiQsxy2KD0ZoZKhoYtkgZLPQBbI7mOMgAd0lpM59hTmNJ4Yt6V7KoiTA/P0BZL
ruh178raaC3zgOTQw2cw3KX8eRWzbh8luHf4t6tWq+iW2t+so/KPRrH2kvFZEvmP
SqBrJE+/TER3cEGe7B7n0M58xaGlSp8SBnlmg7hO2hn3ClsuqAhvefvgwF20UYN6
ZlNOMUIt6CHUYFqxOgqneoQdcf9AANBRglQ4W1k3coyFUO+XzoGxz0ljqQSh2jqL
34cgDb6U765EZb0tOurk5tJxLXsJcRiNHQDiYRBm++jd+KidGSnSLh3ZHiMzeRvH
WMsb286NWPn6pl40om/VPzB0aa61FJP7eX4G53Cu1+1KKsHaDQfgXMlESdUN8v7Y
q7EFEoawT3tdKgUDx/LNS3m2R9ouuPf4xnu4ZAquWPGRYdqKMqoSpNM/WFUeA9V+
6FKREsHg0bshW2uL0evrTKQkmqi3DS1t2RUsjcSMcisRj6MsPEAo8c01r/SKdR2n
zQOcS6kcCHGkv2yHvq+ydIrK5Jdo5zx6YgmPeO5/6DsYTRvmR0wBj8WWwXLuiqoP
bFEZ3sCo8Y63E0mq07PnK8KcPIaMxtezK7Y60tu+Jcz49hOq6SXgEOg14naJZqpX
RFbVJPiNgTnD/ITQC+uBu1/LPerRB5IU16dWFeRgWTPZumJPC0zHGtxVaW0eBhkg
KBLE2LyE9/nwEgk3k14/6AZTwkFfbvNz4yazaOtsILy/zvfLnysbrR81zepn0i7m
SCSW+hE4vVg0SkZar5JG9GzCkiQBnbyca52liX2XTwKoXJbdJ1hqHLjA9/c443o7
EYbBx+x/wDM6NIsAJ6R6Qcwic5pNWkmOoJ7H2KykEubiMVgV8e+dFbnwY3eeKOHL
/LLzc+NJM4mL5bLS7YESq06onSiNTkxPOizu1VgjMI8Emgc8yijcou0a61PwoNlB
49IsTnZrmZj+Yp9fJbU84HMZDjznumBChB8dXTJxB/SXdvi4InLTO6k5iurnG+md
fwAXP+12j0+9y6nO/ThChowYgUe9Yg3F+q0/Y0GYHxmCZ9r+Opgk0C1vhBXkv4zz
lON/GfdXl8+A5sC4nZQjCLPIQ3z67IaTehhFSFgppz/1Mo5+0s6vBLRfBu88a0Uq
hVplt3om7c1NX3eGDJtNtoAk8gjivzowAxPEoEe9TuawzeEgBf9HCQfUXian937N
06Zc8PWYU6WkZ3k0eeQzprss8vxD3Jg9OVLFWztut6xqRFI3QMoxkXGHou48/25O
IW6kEnNydgX189VxjFViyp+nWUNm3gN1v+vr5VcWCsOZkaQl4Fe6+vDL1jM6USxC
ximmhMAVOd98fdjiDHnLvNJagvtcJITXntNI6Kg/tvd7wK1yDvCvEDEtz9p1+V/7
W27Xw3cM7wtyAMWd2h9HWHvcHF/tgUIYU0SyfGxSEqoJcfYy3f9I3VUKqeNLgfYs
O/XpMl865Kf7a4J+Zpn2tPdFJbkzOXQwCe0/m4/xEZZ9M6KS4qHCQPJKJuq6bgWc
To+8DI9rFfEF4a3OJtwZwTsQw5UlzuePx3aDtzDoT4WbKQDIWadzJ50hJ5+IOH/c
RmC0Cqj6H20kD5D/XVbBRwxAHUCI9ItAJUe+e2ORJ6lpGfkc/iRncqAcpXCxUGAm
IYRS6yU7WMaaF4AXpDxbt0h0d42ghnpMr4NoX8PwywrEKYCvNDlZgoY9sBmUUatu
JyJDUf+r1XST8CUQ08lMZRIVB6jWIVcla4HKlgZwpjot39uIHbsulx6K06XFbm7K
wdbufjv93HvtuyN66/PhHBm0RiXXQsmjqks1zYEl52H6IdafQIe3aNpimtq2y5SG
IfwIOUFdhBRoZxrWeBuIQCj0PlM+Y6wvWxOqqffQBMWZEEUcw5oq+GklTKYXEf0V
bnTU2tVa46jMfLOSJqDn3xikxB2UCY5rtuW3b+tKNL5SvtGxDzNvcZHO7DpZQmA7
U9P+1HUHeto6vGI2LqiY25XHdGy8Me3estalPr2K2VyMCPQzg1ENvMLZhBZJ9OGE
ockFCI6zyUjcjdS7XztfqCwfYWlhDEUehAbgN7+IVbw/NV37ZcPFY2uKPK/tLvDa
6thwHAIh2awlstuFbIBM0gWemhfjJ1FnQ/A53WL7r8qVmlfi4RWf/tbXYIqcwN7I
BJGHostQCOPvD+Lrs2mM/K1CMXSKIGP/48zFViScnPs3uqy5O+NofmQiBETW5ZnS
FTDyxpclXbWkc9TOpfvgmhvoxTzou89s+PVkQ01FmSOJNWO5Q2lHQW549+NbL++R
WKnjjRb5aSq6DDV+xCdvVS+Gze1DlfAN+x5vRnFyKxs/fXXF7eoNkm7U97ZBor8I
nWbqnPbQAEA4tEpyp6GaL0rY6GjX9/WsJZV0E38rTPf768WIO+09eSdJRn/EC+gX
mTEdRdig2cq87T4Y0CU0x9ReGvRdtd/u7sLox9sdpPPD5Q4A6WSruDGnm93e98xG
uq0NOROR91aprysxbuRJUrcKa5RyuU7bjgdQJzCA95Vz9yOG8gX5O09NKTjhAPV2
ZeabYBJa3a2NSjTAJwyox8BLYPXLh2XV0PolJEBQMvnRNShxhWa9sEC3wDotoQcw
WuM95rpbsA+idDl1pwKlg/sf3453mFtXSQNNcSjE0c+nVI9hANUgci20X1O6bszp
G0neIFvLBzcfDnFChoi7s3OSnrwZRDRyUH45cjSax57cM9PqQLMXOaIRplBss4hT
scU13/S7fFA/wrW84Tyx9gpHvWXoDaZFUF3DDaNTcoyxNIV3M8BLXobKgReZuk7G
Hugfwc7i+VVaC/NHycMt5OVtGX5kkga9nI+izVaSJaIdfMEi96Qd39Yb78u98yIr
BlK+O2AZ+zKJsAtfud3TV3YCqMuYEQBbniQhcoRqlPRMqvkR1dvnnd10LegFBEsQ
2M6xQ05W5NOIaFV9l3ueKtoDWWSvuVwGvi3xCwgPaQ6r0SUx1BDEObfvgKG8+IF7
XuaFbnalVUjM7eQmfKMEMeCHm/LbSdfVpP2szxNkobSdRwRU3GglkcS1mxxMR+UA
vwrpMz6VBqhb4rV53R78JG4DrGweye+A7ZGraIg/S4+piiVta2hQw/KFn7VrxLFs
Ez4nV9uoApEpmNV7MpEDkwvSo88c/3SX7bOc1zp2tEV1nijhY1wy3Hof1+KO7t7K
bpflJyhzcAtOodiaP+zCDOpMuhXfGg84dXnR5xaivxCVpiOi8HEimXVYItx7bvzc
HGNkIADuAvje9OaYpNyQI3V8qaDLrLKj/2uZz/YPzOVvVfL7po+DP1m3DjUglUR6
M33e3PQ557Ioh2/eB7nsm7x3WNKuVtRSTFjPFNKKP3Z9Ek2yAH4qJk/PrAUJ6ZDl
6ecZgQrj313ou1pjh/+W+H3cOsagtx5Ln0d536fmjtnINAcZTVcSHAgeH6RfCT8e
u/H48Nm71d3IR/rQDx9oHhc7PQpKqbzTfM/nWYWgnltTK/usz9k3EE9YPZNMdmT7
n+6fkRctT/Xhbdaz4y67yJU9S7Teqkn5N7RIjShnFrEdwBT4atGoHzE2vQmagAwy
iJ9emeCb4o0pULiUygcBEBDU7wnkCMeR5IKwpu5QKYyffAyZu9FRi7CQDj/jRi+H
dkWwe/b+RhyDMNZ2ExFbm+TNq8gnHvt+pnhq9iagxo5GfSSWU9YXGOwMolP8VjZh
4U4aY6dhPPXxVPZDNTGD5P13pQ5Wkx2Klq8DSpfAuRh2YDJZKoZe6QzPyz74l2kH
3qAvo+NW0l2dMjSzO7nqyPzHLZFCwKEfi5UPdbwqJML3OU8ku6AwGY2iwh+/2LzD
yYhBBmdbpzQ4w0w/spZleIN3M2eMeTjzTwCfW8PiMVd9Mudt0Gabdz55MPPAZTln
upsJdr5Um+o3zmFbQWwpWEikDg+DTG/Ste/Rn3opi/BOVv3PMgL/DnKJwLBJ3Sja
7xz8d1Qyy1CFEF7z08uaFSteL2YCDQBr8K/hcZVphwViMXaZBa/wh2Fr8G9thJnT
eVdJG3RY+km71rNdzt+seF5fiNwy20GyonTTty+/Gyfy6ZyeH+zVswEbUdxuHSA0
T4w9T820jxSLtMorpsA2pVYUvCMj3zEIwuq4RBuQ83aZL4Iho9JdA1w9n7WiiZUx
S9Ziafw9JT2xYDlH2RKGbGzndeGJCCfCUfH6uz9FwKNtMBziFaJpKelwqeNV1b1M
ce6F5RcbpFyQ0oNLMZklQrbCakLUDmry7daeYpGukaJjwwqLuoUMHEKSb+WnqwiJ
nBMJyOg/PSc9QcloEhemEeiGpRlObWN/3J7eTm+cAjdveLDrlTNj371UHpTuCYMO
FbbVqX/mGPeDVQ6B+5UkVcywXIy1d7UFVJ1J4pqeafv9Eqk5hyTQSJQ0mZeoAtE8
eXy+KaetNJzRlZuwM4FUei6l2Cy3aJZ6UWe4kzq2TeGguFLUpNjXud7EuknKU8hH
BoCX6p4aZOQtkcZWP4CNie+S0leFg8ZuJ1xoT2EKWH2rd2z7Nfen4Za83HTmHxrt
etHdt7ag8j8vJJ4kimszkafhejsvc+rCjUCCCGZDKwuYHtvp4Q0Hu2jgzopXu5Mv
dPXFd11l134BqDQzAjR30gnZxqu1p8rpumr9t8l1iw00xfKerdwWiQniGk4Cz5f3
q/kLD9kNhOex/3ISd+ZG3/xTXLnbWzZpRZWJzjL0tONFXlYs6ZfpplV6Dcd1bcRL
1rv3kCyzSV89t0Tje4XutBHosBe6A3V4BxMFfR0/j42Thg71N23A2TmOLFZ1pBy8
BKvhPyp+CCoGHC8JMdzlsFs8vrO7qfGHnUOd/+Qxx0rZQZiEtZNbMBpCPkLp4W6N
bi494/HeUxH8ZajjD8YrAGsPLWfk2wL+EouY+3Dz1sIQ9xJYIiLJ0r9uy2euCcIj
yfFvKatcAY3r1yg2sRAloQSkBHnZ24BYbofNixAkXVvPZVVN6mrAZsviCQnIZzcW
tdUu7z9bTW6w3BgE5FhOyp/pXLFQjeqxgdKiNUbq/LCCRTs7Yn6TZR0QrR0X4Pk8
F9KCZXzQD6LtNPe4J8zjNmk6J+IwOk+XjeE86p81IkafIaur2aiT9ALiibqo3SEA
vcVWKliO1BZFTgOfxUIrQHD/kzatrEUWAsEOopH1LKrvQkgAQEst00w8hqJhX5cm
91+EcHowdBKNsKvLr80LwuSTTz0yzXf2cBLd6XG/V02V659KJ3qWH/EAobfOnaZD
NXPuqk24Y542ECCDIXH956QFLkcaPJJDRYLKAWCKSu1p1wqqwxBffRy7ou709yu+
+sY+s3TC8vY4HWcAcKM0S/9qD9xivY9jTahxE15WBOn5NySbrZezJ2GMdXKoFEQw
31BmWBbtDVJiN2wJbP8pptOptshetV7iyx3JcVK2QPyAVXRipxgdEnGXFKQtzLAE
+NVGak6yqHvQhtdvvP0tYe9KZOMTO2/AMpppvyUJ7ThhJ6McDkuwdtset1eFDp5Z
9QUKyoxvYQfgkLcvrNI7tZCsQ7jj+7qbpb15z2iM4pGzUX/IPW0gul9bpr6HWxcg
D0NmyWDOydrV4TM6BUWbnzJzCx/DhxZ2RSLMLiiMfrkPT2jr/S07tkFiR+sVxWUX
l6i85wMdd0oagz7cmeK7RY8DLC0e4t2NNjov/rzs6mMvh/W1x1vcEMFccVg80kav
ApPFJht1b/MgLTr57iisVHh7c8nc37pmOnH1AtFmJuC+DAikZh3ayHb53gnwuXT3
uFw7o17RY0+xA7tGj2q37OHzONlHzkPstYLQViebCXDuc3P6I/FFPSHeTzt64+Sg
e3J0dLM5TzCwE00LnwRGMLESTh5WnWd2AAMOXSzwokV0VYUrfGNRgP3QtkySPS9G
sQFckyNETZ02uUoiBsfDrfmIu6qCwT4UsuSKSYWv1EjfU0FgKjtgyqSmrzK0RE2R
uElj80N9oL4izAPL91tdPpIv1Y89v9QbCBjpdFiB4+DnxI/FG70z892GpmKebF3F
uZnCDEjG6W12xZxHWB9X9bA9UjD44FpW5/BVWRPilM4y8uWvUBEAa+I8ycerEcpU
/V2PN4adG+Lz8g3HFKfEkyhLfalUOiaJCg63xZUi0tDDlDWQKYLzFCBru9ZupcDn
mkwZa6nNkjdcKdavlZx9CJFlfGfaLOrlgInSTdZAKhJuYZoQs64S/fh/HKUB5fdI
JABzhneYfvATBRSUcHO3OlzbRAeWjcbppBVg0iWYdZ6HPJfMlT6OGjjj1NRkrLj+
TRw9nLFAeM7jc1IWc4PNF3IKHRASM4cDVxWqZJZoWDsJZ0zdEG/L3TEjUpN0M168
+nzMurKgzB4is/9d322L4PHR4T4djpz+0bRRMc4OiB5zBFtRZG7Jtm6NxOvceuhw
eYluZERTK0F0o1fbiO0n/QIHnWSNZoJn52DVvldI18c1RzAlDlK4Ps7DwUlMDl3D
dOkHOiHI3I259OLNTWZU2kfsQfItUC6NDMlLEQ0FZhiWQ1j9n7bVj/zztMEVdLSV
D+6uo3VtnhpGkOn/az9uOlPwgcksimr3lTwthCR1Dzf8J4TwSRj/SACwyjayoa3d
WqJqHrleU6p3Bfm1mC44HrPON32SnQfE4qQFpfjyohZiCUasJ4jsAHEoi3ihJpt4
8NDbeSKGR7bDqojT7Ldlx9xNeaNzSxm6rMV/sRCeJ1zdyuEyuPsIQq6wJY0iOx1Y
aAz0JihK8IZnkIQh31dzF0Wp+6qqf2pcvzqTdvwcKcaeaHnxHSvmtSiHYB8xmUR0
o4K2UKPJOXt/gbpUmfqtyBzV+h3CNXg2dee9moZ8r54urTPLIz9RBGk5/sBCRcR7
RrF8ZZtb1OnDhZc6GBZfxoBeCbND72g9lCgUR0Uf/pTMjTVYAYkdqoFTwo+tO32Y
2tfQais40qMobPklKfjeVEAUOpZUZACY85FBg6OK/bnPaOJo5YQaeC/i6xL1RA5c
dRKB2ellXWMlO02uUbocUtPulXj+wIj6Dtzd15bcuNPMckPJcK8wHv2XDx/fwiRZ
jA3C24hWp2l3RPzHqRgsadx+3BmZ6CNlwGXNHcMqRJWM5mPoLkkZbBo6zscapLv9
J0KAWs+hh9PcF0PbNYwuSI1QOHYmRxXyAcMqkN+bBXbPsdvPpq2TURJ3CVu1zrxs
Q1OwoJn4O9JFTWtQ1EnK0LwzVdOkcxjwnjXyPKdH0cyDq0h7yi6M/MB2qW07yf37
xHXytGUPEmRjdwTlJTQNMCGpsWseovIVWc8jypvw2daEU/z/GFKifyoGaIcecU5Z
McvvW9qco/D7HP63MlYlLNSfpOE2fQcxHAr/0Jk+1YhXLpU+4ebYjN3HNkxTPonY
gjpkJALXcH0nAZTZq3StSqM8/Mqv5lsu2Sny8sFkpoZOu+VNuQN9L7iZRfitktdH
a2dCgSeeM1svYBUgFBSoLFQOqzrNmMFy7CDsnMtBwT62CpeTJRcYT7yX6v/CgNrv
kdm0vpx/tAiJi0tjDVzfdBzuQ6XA9ZZ1pnkoTAhctFJ0cMu9jlHKAYlZDVzg3u/c
PUjV2K4d71jrvs7PWt4IaD9806JMupVwNUV0IKYYj0VYZfSF9VnlK5Xpob9sCnZI
U+Ihb2DK1UZGXx32bozv3n0b8rfDK2j6EgwuR08jBCWpClqFBFmxuQFc01cwVmQV
yI97kPIo7QEBJUdIRHPLSm2oszlsrziKVMHp1xtB7Qu/U8VlOUqzGJYuLDd6WcN2
nesdO9HCwm4AebM8NOmd5ihHthV65tJxqU8NOhbA4QYBZMOU40NGlF2hwdMInWL+
oSANFmmvcvEAhI5Ab+YKFOZ3ID6fVs1jWDnHvZyW/whvZAMsc1OhU/XUwKvkI6cq
aQHNC05O+n/PVs6rCLyyIv1tc9rheioyeyvJHzJsNNj6cbnOBd6ryTLrLHAXrwJ1
qTTJ+8BRIXVkDvdD0x2RqAiuItMVPprtJl+7a2c5ZZtTWrIkStzwjhtN6VVBmp9T
wvLoWn8ZTNqlVWJ3zzrD/nyN6MoI3bX/0iUyJNF/t52/airZRzVEoSwzzQFofSYY
BQVOw5HEJqLYBFYSjLTyLhy2cY3T9Jx9Icqh5xYIwsSzUldtsTN6K/76iNK3RAFp
2QErha6+y/fm/GO9zU9naORdAQr0547EomXM4E2ESQ2ErgvxH6/61vVrGdKRhxSl
XEIhpcMvWLHitOYev/3lFYNH2IcIfBXTOvnZq7aZYuHFwIKschFE9Wq/L65Ammpr
cnqhf8LnTLM7YqlhHcv3AgNadz+EPEcaSlldTmfTBlJ0aF2RC8IGzdDsC5O/Evat
LtxdClrzldSY31uYlgZvdf1XwxoZQL+HtYmPk+QfMysniUN4dX/i63RHKsB+Di8V
2KpjmoBTZ8B8oZYV9yCsfgPNQajSmonwpMW3wz41EH8lhcU5p+SWXyMvL8AHqGKG
bnL9S+EjdTSP7jGv1LXQE5CFFUpkCXreOdL4N+vwd7dDG5OgRs6VLtx209zZ2Rsl
PNorxoiP/YNPEh4/hWa7bcelVIyRMw+Pzm0r9v2QAGxz31/+ZFk9BMRtHjuCsaII
JHMQ+EbxbZopuEK3RLCYHEdbnBu5Qei7qJbZUsB06lM/K+m+vh1DCsSwa/r4w+WA
BGFlUGvtdjK1/JgoPAXT0FYtiSBBUyFMsqz9OSee0KU69HO6YkJ0tpr+89u2hoqF
rsT6/pRFpJCI6zm3X/b8rZMkhvVfuaSiAsvZyJdlq82UQhomdpmS13aLzlSmH43T
f2WII2mPRi0XmIkOHorAi8PUxVX1bgL5NU9h2OPFn26ssoDUzwc7qU2ch4hTDZJA
9TS6bBGmq5Q5R2XhK5PPEvFWw1BRSpYk+mZCNID1O6+7h2OZ8rH0LtFfUmjppiSq
cfkl6+d2C81t60mQezxQmBKlwb5S1ygUGsfLrEOLNCgbeCZl/19M2qsL0zPSKPWb
kmxjlePlBnvqavynvOhv//Fsl8XNyRJbAbKnqLDY/CKqgbMm0O6aZ9Z8mFLflrbe
LaiCka7656d8PkEzXWXKz78DExTKXwuUnYc5h6hZ/6cnbfqLfb4lgkBGD+ItrDNi
JxnlJX5RHMrV5ngXkO8fg3IvzyaUVdnYjrYxYrJrArgJn9cqTt8Ke9iUrxyGNccw
fuBiZPFygPvviRS4odsWPjGktegLfh6IjpVw0tDJ5khaBtkXlE6Jsu70uySNMUA+
Tz37wKRxa9kZSmsdDho+JLHAAR4AppkdDxXYclV+yWXRNKpACVJ3QGN2XgJHAbd1
6mfADfRfbsYpaKwiSSYIFiQOphLg+lm/tDwxgoOJkpS+WZxlG+HCGHK/cGbWiTLB
+FnHc+LjY9ZUmeuXQzWZrd/tAYSFglIE7MA9VdcA5X/v855BjPQvgWI8SucjFNlH
a2aPaJ+sk88gg9j6iutkOGsmuv7+yyIGQpjkDkfRXqYfRIg0ooSz3PvwTbOzzUGE
ZwpsR9aanHnUAunitv03OPKzxApJiSKVNAYDGqO37mi+ZndPVkfmjISYbFASej5C
Kuug0yGgaZ4eMGQO3V0M/mvU/jAIguOWq67fFvX+JZ4W36pdtUuRRWQQy6lfercE
IsLR+HTtCUqc6QC3Akk/zsNpbObP675RCUkGKj+UTX1Rvmhwsfre+yKyyXgOPhnL
kUL8wI4aAz5tGAZwf41QS6QEYhMLiJLzW18q5sDaAHCIrM6K0rc20Nxjq8C5x9yp
GobtYJfUTHsanSPaSDkUuJdRukZKU2F1YXasWJxsFWP7Hmyl4SROhq9C/xUcOh4f
0gTdZ6p02z4KHhQ3375GREtYo3nqMOUy9Fx6E9MmfD29dsDOOyRsujihUHZ70L0F
M0V5gIgC2Rx/XdvIDDd49RNSdu/4pZFVf0BRCLg7hRpnrbt8MCqjqbw8ZMvhdXPi
xPHwhP91mg00NH/DqnJni76RHhhvFSTaCXHXr3idTtu9RvUM3t4GAqavGKvCckBL
KfP/OUGVp4Of4S/G6z2zyP/ALVEYj7nXvT+KChSEWnVozLOAIAIZmrb9Fg1ktDoU
v4bsFn7QvUxBSWo6OeZMUw1+NPg8ZXUKkTuFPrxOEjSIS+t5nDv/5WP0H26HXVHv
xsnvvGp3eq0BDXyxEYyqxhGiGz4WI8QUseuJvM+0YLD0jC3QG5vFPdjGQb0K9cyO
fELqxTTXw8H7GTmI0QhVOaInvrVXd7F9Bvk3GxawpQkT19DS5weXMMC4x/H7xOjp
NaRLBPabjiTJe8kX/pQFK9toC1j5X4q9glfh6E7+GL3WBkmqouWLOkFeGswUMbIO
5jcsTXlpYXxnhoUJORL2QrJ0yzsVudT2K8izFoSsvvxK7Dzm35VNsqlE6jbpx0ag
+RpPf45NWsTDzN9tflIuTe7cEEV7ps7sQU+iXS7VimZU+IiyLnBdXnkH7ZX76xkK
QAUdfBuoPSGOrfuM7pb6wTHAfbLbTwQukUQjaCHkaFXaXh9hPASKNcXoAI8/FC2X
ChLTeuq8Q/OnOsHHGGHJiE3fLyOnEklZ10JMVQ2trv8f3UBFnWHnXqB8yaVo6mGe
E4vk0qkMXhR73PGbTeWg77t1ZKIg8m/KfkPyiJ1Ja1LGz2e+d01TdhlAJ0yJGlKa
iYU2QNirjh5FCxT8Ajy9z4s5buEkxMy1tri7zhD5fxXR6ZmPUmCPlRSs3BA+goLx
rZ9fu8VXJD9ZnH3v5QZ9kckabS9sSwijTtKYWOwYKJVxJO80Qxfq45Rctto9XHV0
afGGX+yeRCQUq10Z8eVpM82xNL8//h2sAujzfCCs9TZqrjSblPCMq4uJO38nt+Z8
pWos5+XEEhPcKQ1BdNZbfTDJYXh9P7oiQCtsAYEcixQ42UUk2rRmXjg+Du5wX+KB
fj3tx10FbQHS7WQjQk9wOyxQ0AeerjDz+0TCElV2yT5AeqMMMHidxxQihU6uPCsz
WkuGI6RDUNU4cMYpRXfoDdLDB5xrRFk+5jEi8XrmcDRGFMufPPyA2GrW5TSBWDmp
hp8tvZ0Vnhyig/c6jqBSXCDqAx8z2mCY29EI+2aTYqm77T/QIAF/eoDNPocKV52q
+97+LZVvbMr8QYeCyaAF/R6RqWIq3o2AknZatK5WD+rCV2kekWqJq+x/K2K9WzTY
xMNWEylUODcf8rgbPlzUk2k3lxqUHHX7oXfyS7fi5RhKpAYXq1JuzUGndoBgunA3
3rtZQfWdLsYyQXXgLvlAOod2fo3dDQ6PC2wSL/46V57e5eiIpx3bBvtSqt8ERACt
Tx+iYm/BRjKc73b6OEGj/cQKbzdA9VJMHRDma6aYzUtAm848vVE1g7/Dav/LurYR
8E97fkI6brToi7rkDQv6tf3Yv7vsboHXa4qgMFeMz8RAtqbVkMdyaNssFxMpyhj0
Usk323eZZslLb5Kdv6AXuUSEjo/ovyo3MQkbcWAAVsVfAAwuVj8q3Y+5FRKtLZKD
enY1DOwf3nc7yOKnaqDnF9p0qlD8uciAQ4E2zcTs0UtZo//lsOA9Z5/IaJ82sUrS
YdHijvgHOSgcKFyPt4W7Io4eyKtz2B5VeXoNQ4fe5lEJtzdHMZw9ov+z80xwWZWK
0EiLzrYq1qg6jvmajIUIGJfjglawJINmriVMSXTkdFxslpM3RgMEHwvabgYubUYb
+o2mX9o/e7q7tClpdDUrrNC0C8XF02lkNJz/yPHF7qhoLrb/uiq4Qq3SVSjmnYB+
Q3N/iVJjDphJJhOml78E5GghYMWbCP+uIUCfDZ6b6TpEtZUV4n6jYHcKhp1HzjWU
wIUyj0kuhZVF9ub1ajUoHML0J3s1OXPwBG9stfKilMH8mO8FrjGtvdaUslOo8sXF
U9v+kRLERZ22Y6BHlB8X/HYVdgqYTON3HBc6fGA3kfFL4p8/y57+egaNw0BFlSHZ
R6akEYgN6mY55PkkcryFAAajeqwM+aQcTX16Ugb9BpoSLhGex0bwY1CAKOGYqwqB
8JHzC0PwZgQKwbtSHs7OTNebthLv4cwk5T57yaaQ61sxDXab50zyQJvb/PNcKWgL
08AVMDqhTLzziqL/CLbIQLXw3hjbgjLIALg6taS2UON4jr7ehfPKlb9cjkLfI4Vl
cIeAWx405ubZjD/alNe5t5g1FG3vVpv24nxwyOluRCwBriJq3dISNqSvjMo38L/B
48KGDugvN+pqSqwIABiH8shF3hM4LpTbCanowWVNrydc/S0taoz2haekpE6FlV6S
eiW0KqSI9xOqsllreqwwu6MdPefC8AW7zHw7PG1AG0hkPZGWmsZSlkiUntm1KJib
qfDTPPjlNTew89dxKu0vuOMPeSLc7Lu2Z+v/dJiwvBBrAgB6JobicO6/XeIH5cfl
QwQcYqx/f/2W5XzoeJL8f4wOfSIRyx5dKibOFc2i0D3qjv+Fl+3y0Smo+zUiw3dX
ZOdThTjbqpKIyHYCepdSpbBKougV6nJP+m13oFJY/YvWN+60Q5v9649rKq/PSpQl
j3/yyN4BtInMHBhUiECVNAgqmFcimC2Mmj6pNMhD6BjC65NuO6701WMI3vDMpuQn
0OKor1wFzIQP8aSeb1keAsWHz/XOITOhiAwWi7y4M0nlfuglNT0AMxug/lKyh/xq
YU6Ko48BAsgSnIZPqYFczLARmKXx4rkBpdpzvgxQ6+J5vNnAS1dO0fifp4+SaHw+
8xGsqPkMObUh/GvNlGAz8BQBS+aL9jjL9BZGL+r0CvGDqLi5PujT5gg72gifeVXg
WWjw02OknhGH5/RTKhoM/ALRRpKEmfzw6Yxldg9QdYekqTnr1CsYK97cIwGhW+v9
l5OgfPRoaMwwr2wuPZnnWKsX/ZwAqH06ev7BAxkQC4fYpi0t485lDrYo81hHswfp
esU+ZidiUjPE9+YR4UgDZZHSyh2ip2DqUHLOvcHwQKbjArSHUE13r0dl8XQyaofZ
xpqwSnYZJImVbh1n/vE3qGgN70LoFyS35OSRdFKSqCasx2jWBgiEzYhnc/n/YkU9
vkZDFr5l8z3e2rV5ZlVDplK5CNy4k/07pu6cgZUolNCAp4uSDHSttDqzuldohvc4
g059nN64w7O2jx5jJSw3idht2/PrA5o9A3AJJXmc4yj+EcGtzVROPvKQuR7TxyjC
FZKrWEtehMB8GO/Ot1Y+MygUpvuXF3zKQOtTGm/rREyfqs7dDF20StNdMKBY/gjf
8gH0EA0BB9meZFz8ZTPCb4hLEUXpsA2uBuXH4f448STQahi3SXOOowCAx+lnUxwt
r6O8Foel7s3B6/+MTEL3L+3dAqRhqTmN+gqFEBsbBWSS9oWW5CbGNK2p5SJWjCgY
cMIyf6cxr66l4X4NDoB7vFb/LW1NdWr/uO4HFWFM2//bT2v3dleJuMsbzFIAiW3N
uKg5OYNzw9ssROT8QchRjIQqAboqSWspV9CXup9fbPoKL1XUQnFSdZrVAXiARi3h
B8qMfLJj/5P7l8L1+zYja/82Gxtg+mQZ336xt5d8Q1604gI2nPemuJEcGdpI8fgK
3j6vEfU48jkCPESbXMuM/Ceuu983z4xVFKjET0ON/AvOdhUL7XxUapGHZRCBKrQM
GSacbXINTDJnDxQoVegql+rO+uXODkHTh+N8NdMALLM8ZvBv7psgKSv+mwVvo5OY
t4GDlA20435SQpinNhdQydPjsL3FpKMvYrCf6B0LdpDOVrCrTgF8yl60hHIkN6xQ
8oE96E0Sew07pJmcHExr8IiA5g7mYkND4nMjzCzuFHJFZSRqV84HqSylQC8YxHo7
vHb9NvTN+WRlyH5/O8OhvLznySmjxWptx6ZRYXcbXmV1B+i5xpp++wv5maET+Iyk
0+OoOK9kPRBbxD6qpXPbpONmxseaXzf7mVdr5yuYuzprzsT9PUyz9fFyZ87N7+Y9
f9Ng+1QfMVXp6hY7Gs/mne9Aw9hT7+sYyb4nmPc2Gm/NydGAQy7z1SvlwL4H1/Eg
/mpbmMEDwWXX8mipi+jbtZX9oGb7hUmCrjPgsK/otnD/egZokVVwr1tOXjbuJJzK
2adzX2JXRAo/ltwY+Lm0yYlu5yFlb2dIkq+rVZ68f956e6XvbrBf6P/xjigwo5yA
jpVjGjgBW0keb82Qb5QTj7M7C9TL6JLPwKR5HOzjwLl/sYqUZP4LFs8HYLVY9zsn
E+3plmKrpRv8BTlLsCBxjoJlagWl0LBLTIDrCy+yMDM7WkqM2772rgfvjUf9ejy+
W44u86XO+zGEHzuimA1bZhwLMXSk07j+zhB85iKlenR25iT8mkqGeE/HRSTQQ/gw
yOypUS1h7WikKmDzi2wf926gCm9nLT2w/o6UYBFtSRcH7+j1i3mI53QF//Q6FHfI
GvS8NVsxy7WE+pnozSnqhc9YCAqAEjxORzGMx7+ryqfRqpAjOPCTKtJsyeM0XPGc
UbgFYo1dsPAGHVt+kVi3ZbZJFIV3opObh5fhtXxGaRCCBrdZKfPmHsl7rcNmZB3z
3Gm+mzmmkTv+8GQAvb8xj5G/caMAFF2Jz1mnkaGcifV47kqwJq4LzHYZOybR0VKs
YAYZM6NvxiKOchmoZjnQVHMpcRjj0Ts2b+tHx/V0QY9Vm6E6hPV4ELposZTRkm63
bzwWMkVu3PLqqObk6GUnTcmoopgmUo4ULFH3IhkdGrB0H8KJGlFtW4CwamKtbRzN
LGjQ4xOldGwv8qWjcRsxVzOKqx16f25MXeg2++TWKKl+Dcjk0PXkHzfNe4NxAwU0
PnKC4rLLqbdI598wDsX9z+a7VXRGA/bcYbzmZnvm6LdLo2aN+Z6ASDsmVpsN7sSI
TRTnzkZEwtEC6KCz0ej7oxHqRe8Z+pYnR7OJlPbdANiUc1mPvrdjmMUrgIfTlrpT
6yVV5VQefHg6oI2kc5wL4nBaEFZflGKCkJN9ZQPVrAd1782B9AGxF2X26E3X91Yv
KkqKWibYVjcFw6I+CqleEON1lWP63SJ3b7vok5vzi5RcVT7txYUS6h6K5tHcam6K
5nSrxWdWoKe4OB6xFoBW3cCKVUaDC5wB5i59+iYwAyPYDO4XA5/6B6MnywsV8GCX
qdWfALQsG2remtiahwu8xlFM/OZNuMomVyNflhb39vDAOr0h0nqIALweKPJlyUvh
Kx4WGdKvYkBXfPZ0fixmIblmoo9aeK0oVatqsCWYcevaYTbhuXLKkl8e6QJGH85i
iAPKHPjTXoXQtMIj12nzTcWWsjdiO5kbFo+gnSAGZzaMfUUkVs0I+hkCDkgmyyYo
ulxbVdDFMND4NtGukch7FFi8hC4mECW/sI32n7ab6QFH4MUz6U/XBUKJ/HZ8UnbL
oMgO2zxDagk+IN/VEi+Z+Gc87ooancilioDQUIbFLq8lFjYwCgBRL+3nKKJCaqj6
faY2c9xsKIcrFCHe2KLVi9T2oi0hvxyPiE4ZiERzQ70gZFdrzgoVo/T2wT0LeOwj
uMmBltIDaU6MGGhcWtqbCHErzxEVPwGjqZg43aeeehJuOtdNRrDPkvVLoO/07Oc3
o3j8G+4hJ4HprYguYMFAIPtv8cdFcQ+5ARcUWmxsw3F9vA5paT7IvyRO2Fw+mzJe
HU2uW4EMr0u4ouwTpHTQsLYRnYHiw4M3Qoj9mpZn/rH1F/rWLlkZklsWSvx1q3wO
kmsC8s6OehybSTQW+BQxZhB9tBeexxwVeb3hDnI+fPWL/sNdIqaST5g5ZXob65ai
fQ03+0byIpkltU1EeKBe1oqkw7aWWnEix5r+8SQ9l94aB+bgSz8mfIKaaqYfPBE4
yhUkdPSxd5cwhmAv7rSlkplPw8mcKuB2FL7Z9HySrQIbQVe5FzKsfqKNqMKLQZ/I
EVPdUVhwNlbRrgslHgMDQaCh0V7Iuj5qyc4gTyajCaxx6gEJUkP59Y+hBe+7c7Lq
fE38qD5lGGYg2oRLIl68b1VYnhQsSh3hmVNhNBcOU2PWQzbAYoNi7eDjAzdCRFZX
oQz4B4rfUkttnkvdTp/Q71X3fhkYpaUjuLJ1p3UbvI6DsOh77PeJnfAZdFzPKEja
oPex8qQwVU03VlkPcbO3fsQYC11lyALoWlLtkU+Yl9znDtRFsvJkQ8UBoMANI/n/
znjTxqI3NNl7/Uu+I1Skttfm8yQQzXLZF8Y5hae+e51GzbtlpyB4KivrloaCrGL9
8aVWlDmiqsnW7evegOWYyW7W2SZk3VWzPeVjJK9oDLGDZX51/rZCPQMT/lxMR/3J
o0hx6pZmDuFIx0gc5uk5Cp7/BsW60v0XcNtdai9fgvhzhn3oCpLJrIRR57Rmqtcs
GFGhm9DUQwohGSogeRK92tB7rPOTPQ3nBXgbpJBBKMsFlQr2lT4ihX2PsKmFs38W
yUrU1jnsl1rohlUL71Yb16RqlNNTD0kDWpCtXwlqIU5V9eJwfm9AuZ7gr+53rjOl
LN+9CvylJ34RBTNHq9Pm+H6NqNeM6FvPrhQP4EX3nrJ7Asmk4Vpna0Z0qvrt256U
+pQDNyHjdOC1W50JI+0hfge7S32SgN0rPXHNlaIiZfVmYM7LtmSvA74+m9QSplrB
IoALiRt2U4/WzUTvaq8GKWv1IEsqAS+yOfDi+LY1jfaEQehNYznvMdi6kzzpuGnW
7ScWtofcOkKN9iJ35CvDXz+k3pTfVOVoOth8fYTEELTKyrxOaLrefTPr8uHHmexS
3yj2pNh9xvOYArne8AbrvRjAC9kU9nC8NuvhkqVAHAr5k3B11XQ8UhjYA5zi3nSa
+AFvAfXEdqOntfx1/1+LvYFwAU+UI5fs/r8oORT87RLqPacfBbLZR9s7rhM5+Mjw
yLyiub4EgVLYwm2/ltcGSD5g1Ku0WdPfhqYqPWPffUpITI5QwzEUfdeb1vjdKtsO
k7XcuFdTBmA22gCxtaKY2sXmdfIpMvqEIjwjVFDS36u3ynPb0Rsz8iy5U1RCmxSz
8Tl78NRRh4tosYNRCixH8cVLqBxUM52Xh/RAUfTcjqLjj5wnp9xD4khBaJa1DGjL
4oGRaQOYzLFbKltsBgOqRBEnD5UyJOqQt0tgAW8ptE7j9jlTTXAKiwIiTqMt6ZUp
VHFx/2EgVR3G2Hvi4hLFxyOxUlpa4aDczvY3tz+xWfsbSarFAbpkPrfmyiESd3HS
FyE3elwPgxkn0MzpB1yiem2Cy4Prku9LTb8SD+u9TiBzMwEcNAkQtuUHaYbTIxu3
++KUOhKziUnbJP48LrXEGOIjfEhBtSbvonMsWOXkt3rLAsbdPV3/smZ5Wl4XW6kZ
r37YJqw7Rycjm+JmYNu+1ytFLJGXUir4ewJNZ3zPpgNLkeinp82zUs5Hnh6HBrQ7
TrfaRWl1185RhkT6fQ182+MT65w3OGP962yL6nrk6rdoBa5X3H/lQrxj3VE3lKYP
v1gYgnerbSIpNYQwbvlyskQ/zEpHSLPI5Dzp3d+c7ESrbcdzjH3OVn5+yFeLUPTI
rumBZXQiLpvtk2Ex+2k4yOLR9dcml8+3Yig641nsV/FNPS9BY5ysONu9rezrUqB/
kBKuY8xU7Pc/F8zy0mIohGW33TzpK5Yz+AoFLYWEzNF8AGE29fzbSKKk/ty79+DQ
wx0V6OwuY8079o9EkPgKGfqUhX7Rggno4IPHvu5Ka+efQTx8NtXUW2M51rj2mupK
kflp6xzNiXle20XmiQVq9TQJtOYjDIsfHkutCp/Msu7iNh2ihYgH3/dQOvWJs+sh
z76wcjLGX6/oaCDqzlq2FoZAUfRZNud/QKww5gMu5cm5P7ZLoyvPYS7mnMRJ0iF7
f1m0iOMTe4Afkjo5liugqW7dx3q55ama8k+VJl6mLm0+iDkLNl+wI/pu4CHieYox
4w1Z9cw5oQ8aOjVmn9ErMBV+p2JGVkYJR/T9dCAEfHspQ1oWBDTzTF9fHiTQNQ4V
xnX/onCkuCFF4hC7uGRuQg76RTu1N6yN0gKtovGG2nAQ9lSfqi3eSmCrF+kneuRJ
57JP3MkI9GrGxutgunaUHonkxgwO2ccetLzuEB7knFp9zIEabD59APD1zHDErUrM
sq1am6ekTq6ueH80fGcj/4Ls487lTNwPz/i5nEpRbA8heRKUGnWJe7OxLY6DTevM
bFcuXZF3yMW1mz4L5zUsD/dzk5ClGtE3Gw9/hGsHLUv5ohw8URCOLbLbauBcngsU
CzJZHUrNgqAHnqaUoSojnkyrtkFznWHk31ejeOILl9BSuEDvzfcBettmq2D7848S
0dyJFoRlPvj7AA/m6hWdu6n+4TRgyc81jCA2W3pgF2ah3yuoreUZ6K0yNvRLs6/T
ix7JKdkTkeOq35o6y5Ri8p2t9M9O0t5bk2xlQtRVHLDrtUyqdfQhMPllj6Y0Kt9+
nwfS02pYPOkiM/nxDLcycDeIoyOZjAW4hYofNNrPI2vdc8sYyYSohP2TYKZKuXiA
FGiU5S2v0wdXLnYRGdPy5xm3F4VkBBA3rqRyobbIotBr1d3Qyh1QFmUEdJVSdu9F
xUg08Mga5lbeCia+0dPzQc2S4qRUk9wHqG2JhTJWcuRJxa63UJaMcJeV6Y6PDxRJ
PbMchQhS6wQNXxoQ2TBnvTAURE7mkAjQOuAUqKrqp9roP/EY6XPocvItwS5cLyVW
lHLA04FUwTlntczXJBC0h6p77zG534uSDKIvG81heKgQfjXcvLWhG7RkA2krcx4A
K1V5Lp3gj1Q/oF0qj9ar4IayMCfw0aeCtMAJApxoWa4SALPivpwDP4vGlQQjUsBI
+GzoCCZVSwaxzJyFYq1QoICvmn6w/2uGhzxysnQT+Q0XW16qcvVT0EUk9Sfv6Ich
iARZz2tL3GB09ggaVdrT76tv2TsiII0cwHOMRjq52aTqVwd8SEkZRWq8q0rpw5jV
vXVFH3f20CakBXl+BZwecMeTodQXIovHFNwFtgJeLIn88basBA1+ptIneiXc9tuv
ewrDTAy45VTKFJv6mHBHM8nt1L0nXLkKBd+0S7DRa8+aFjKn7+UYjwl7ofQUvKwN
qXTw0r5EOInVJMl9USHWBng0XxCqvd9YOp5zYlU+/X/OV3a9jAj3ZAm0jHnfp0WY
mtETUO5SM/D+gNyYf96nSbgEMlitzBWUXiiYpkZrlmJpVj9ndOCpXm+xxQ+4wKus
+hKDAFlAJW2r9CrHzGcqqlXm0/38UAE0N9/NMXdZcmruUP/Qeptupq4XyJt6XtuJ
tfan77HHolBRDa5sgEFwEtSak2EcMmE5HoK4Y88s08C2CyoZadIgXzUmJ4mkG98y
TpJRtWXR8HgVozVKmkGC7wzRSCaw7XKxssL9/v2KOsDzNcdR4lWZvORduQYdw88S
zoLjiQWb3iVb8txOzboC29Tj1FGehHOAEsAk2lblkfv2mPncpkBIYveb455KeTuG
Ng+1PsdonJIcbsnVZrBJ4CFaD6oGYMtNfaJQpTruA9DUpbMi9eB31NYyPScsOi69
QSMvkX9N4nsHVYy2s7mNO8AvUBtzJAzRBJWyY8NIv2xqxL6QN82JlABkiBaZb+3G
ixOrA4wok5cSnKeX1TmktIAAUh7yOcynh1N+l8khVOjfQg/zXm0VMDh3w6qAAARw
Gqg8CrpTGBkBnFmiKf037QCbcFM6OlGf2QMd9RKzcwV5hplfHtn52w5HvxSiPSoT
Temt6cMieE4XV7ueMb7rAzW6tLf6oGTuvV44Ebamk5SFB9w7FOOHIjM9nxzrKQQh
hr47x5UoizyIrnTu6bH1NDILXRycguTqLCNR9EhdfSZDCspPXr9ooELq2o6wYtSo
ia5SUhHWgWjd/rnh5osIjWssbCxAKyKM4hiB8M08/RZVqLObi00ucW/SjpIDiwct
mTM0dAhBOKG+Lvnk0OVLeLg4F80cjL3c5nwYSEyBWTJVRYyeVdQ/3CnNjLoY4Nxk
DJUSOd+GIU/5WbZF7YIMM8ESaiUZLu0S+x49HRRO1As3LTsR3Yg/2bhC/L2EUz/V
+drjyCndQCUSLx3UUnOLivL+mK2N73R+8Nf+Sf9T5qfKRsEfWBnVSAvujlxTEBc0
2A12h7S30Go9q1yOQ5yasbrnt7U73zaKMj+jTzA6XMcwPa4vGbiRCDY9jAlcgIhX
udbTq4B21Z9xNGBJO/dB22Ym8o/5C0K2/cdQQGSdyzoQnb3D0sZxmB9aGLMOrfWS
pPxD0S6nHm3Lp3cedH6M54UsElcgFOJsId9B5xVi2srh26NI41egehaGQp6Drgyl
saIlOTJqiOhobAlhUxCGvUm+596G3limPdbuTbYkbMho8B0IPXguKqWhwxJQe2mg
r4eiaUT/bz9/QqA84DnPwLhfdueyDXRosKlAoYxVacOypyZyMKMltm3WeS7YVjT5
AqqruSpK0NgSVCD9EG/c1S3xE3/deVzg/0QvT4+14At3l4zEYEq7M0OoDaHf2v+T
xM8Ew8AunACfPfYSi9d0NSQarTga/uWsdxjiNRwVsX1w7XTH/iqUsozorE11HoYZ
TuPOjcemIgtoAzFXBAWW4qs0Up+X3jQRHl2/PrtIZTK3Uug8hrJOCw0IRdua/W9H
x4FK3uXcB+SvN4T5UNJgOyFrs20Vqmaip4YKhD2cxC7GYuglau1oRbUVjBVCcb1C
fARNllHIraun8NbZIJITp+rgGfJ7/H92Ya16guL2pQyShbzE/L0VPbcYIP5EOl9w
4tLgnC/HaybK3cUwQ7jUrx8gw8cg8V2vFf/IH+Dh5BduUpvJBF7vATSOKSRM8Er1
cByRhqKNm4DXjfdSC6/9yO1GkEMcYspJkwFPvn7iAYwwGRK4o6Sw+0aEzEgx4AYs
jVuuDwwUea7tpvUVVOc5PM4IIi1sxatA6+vRusVsWJbdR7PPIhjlcN61WT8JKzvL
BvQ+BXMyekSsNhNg9NDi68W/UQ524aNCB5gbbQNWmOcm4obEMIui7TwsLjlaRnV7
G0hqeJPdRD1UUjzJalHaLY1gBkfK7J0aZMkw11lLv5CGdZQbWvGguvP7P7Vq/oXi
LeCsywNtGQEcY1/+M1CaGNZJE050o04txy0AtXn0YMXB40ZhcDOqcrwMnGhesg10
0E4n/Og1OJRNU/dNGJ+uCbN6hbRgsWz6ip6HdJ0ipV6ZkDWBFbTqQM45pNIADTwq
lQd2vFZ6pyF4SSNp7EU7Fp1Hn7PLwAnUv3mSpsnz1rehP6GVbdcH+l3Q00XlssU1
pMAGHQTYCflSTIvpoO+DGVzBj+VCYn9FKSpcQNw5RKRk3RhlLO/fszW3NqAHj/YC
2N3nEvnclVbjxax72nKPsY5j3MKDUccJp4p3E6qNiwZNP7Rg7BPNh6dqrEWdGwEd
6p1uOyAHw4s0vhw3z46ssEEdsZydRwRuoMh0X/W6Ljnxa9iv9TR8jHSJM4lC2JPB
WtNhcaExDFEPGy+XePAFVR4Jv/sI1xdDn/YanwXwEP+bP8rQFRRfmMc2LHqxKxI8
Z4EOXg2I0KvkAC+1wEaRKVONzAN9KCDesKBKbMeV5CpDye9Tyky4UECwmN/vPDTT
x+uGwjQ4qSI12u7TvBC6zwrtNckRR0+GP6ym2PZdhLgoUhpeRyzPHPs5KfD+sFKo
ppn7xYhTbexOOvMY2W7HQd2Al2TBVWQlGKA1YaJF8Mnzl/6c7NZLuadcQV/kqDzF
P2tGUmQnWWLgePvEZSMcgrRsweFXz+GUqD89c9LuJSo3H1YpO46y8xjKtt62rzli
9rG+uvF/Zr7g8vViBgNaaAU3kr/wdzh3XVmeKg3kEA+kxiW8TVZxyNdLhEJP76g2
i3h83ICungd5TmS9YLLwK/8gGyxpkw78TAnXonyjkIeMoi+cqW6QDkLm3OnI/Ndz
FsKX9XEr4SDKb9ijanUpX/1KvqQYEK6Ou4Tbu83zkuSsFl8hU6Rr+YV4ktP0PAUR
Qw2ZGC5r05VJPN03OISYRPzN4piS5WXkRQI370fIdXAwDVkQeDDKbP6XNNIeTh4X
N4gUNU/aEu8BQ4vAK5x7S4xhE86p6xDhvuAm94E0JkDLCBozzCrlQC1ia4MmFNRf
dZrXnUI7vybW6eLj7Atm2xcSjobaRY4wyGHtycj+ntuUJICi6yWaYpP57yaeb03r
W61Zp6jaqvSNc8YPyRUzdiC2kLrIeSf/z/fUhiD3YfGsCnoldF2Npc0uIyBQMT2g
67bH+yxh4KZmSA2bdjg/romm8TMY4NS7uBEeUir3MQWeyc80AZjfs0lcy2d2hNLL
zGs1DAjiWqq9LUzvtkOCi905NAEr+bXuanAfTy6ReBJXTHtOUTh12OEkPycXgrJa
4INpTA7l4n9RY6rCLQ3HQUbOqIdSAvhf9FppcYl749LG9LxZQX3ziK/zK0nDutHu
1GeHHvx+9b4YHm3qrojl7prgg8nqVoV/HKZjZVWN4sTj8v/cfR+HE3EBoC/VJwRb
ZTEu9Uih8a6o2eeRavLSwEUp0/JKHdfc8lA2zyQSv3CqhpJTLjNr+3VIQadeJx9G
5yR+G/cWVTDTfe3nt3xnWVjd4M4sH0X+GMnzhgwYQnwo4pwiwnYN+SOggK8qbjQn
SHGLGACN0WDk4Cb3yIVLrhqUDAuwbopFb0i5hTNC+s3J5y0mTXIJ+PU7yEP0Dwr0
+ky4/JI8at+kdMhcf0+9NRJV/oMg1UIzFCtJ6+4OZN0+DMG3dDnBiUfETfxyt0oX
BsVDjgdXT5z/GnZlKCK0VbMOo3MTidTVvgQmiqHsMz0ejxFG1JV9Fibrr6AcrV5/
/Ia1CtgMduKQE9NVhi0cjSGUNg9m8WXLYDNmmFjt3vqycHzK6GYB76VEHcr8719o
M+w0vXFf7HmmHBkohbifXS31IF7M1RlTWjhs1wGoRmxw0VeczMxkpCmfqPAki5ou
xZYMro87Q4Nx54Gd+ueuhqAOiumHXrEmoEHqekkOvE4Xaw2Q489E15Y5IZMQP83C
e4XMIdirRaJ8VksswqDktvIU230QRNHhux6X9j9dHY8a1PggNRQ2a1fuNZu+ToN/
8FEjNUaOGBgFgdDANBLr7UUcTnJ/AcI6k9Wyrm219aUrbaeZzRJ8mdDfY1X9NOa7
YBDQQ5Ou52blR7vyYgUoAEVhIzBWIdzJH7oCpNIkKanWxD1CzdS7WsChjTOAaGZH
j/ehFl36hc/+0MO2xBn49VdDwS5vL0V9JGCceOprpfuZbD6k+6PmI92d36CsE7W5
2Sr7HzWKcY/x/OAOXy1kS/cZNMqWiawvTdNZyMw2GfBRqyTE1LqTV9joVp9V7gI9
Jnc9DqhLMMcNKD+FA0MT86zAYfeMOlyzI5m64bmkpgsiyA56kPZk3gOFye+N/UXa
a603VkGihTVOHNP/2ImJ2YvOBbyhg4HdLtz2yYwookR47wYh4tlUO9YVhNqOa70S
B9ztSYzre8h5kvvAl2zEocyeFhxfBcPDcX+3zU4zAGMkBpFLFixPy0GodPWB+zPr
rn8CMzGwB0TnzdbhrZiNGhIFZt6b60lhF7EiQzjInl1Q3iprWNAJF41GCZx98uZe
S6V+6OtQGiz70gdVGSHxP24c7+bM6iPHvDSsAlriKum1VDED5olzrDPfe988ajba
fop5TFMovlaTmqwj393RlFZiSSqOtlyhJBFB6G0F3tySatk9176w2Kwa2pyTZPn4
53LCwDacYZBkUEOvG27oM183cuGQP0LX+mfw55r17OStycyU+RYAUneiOqM2HyqL
vk/Dy21kHSPeLmv3DGUTc/hVUs+Wvzm3kT3vhvZC0cfsRe0ARdt382lZTLap/LVn
SoDAIJRbJhrQad4jmj+tbvm9gyLLlDNfhSOngxoYnKqRNYvo4rgB5UZ+hVY9sMXP
SHiHKlxW3Zcf4Dpvk+JyNHZtUAES58sMaVw1COp+xmAQlAy/QgND6fz3ZvqgSRCm
Nn0TOOlzAxGAB+V0q9lgZKeOCodSFgSwuNNTM7JT4db6ABcjHixHM2hYWgkHI3dt
oQjFT7jjxz5Nr7RcKpF/b/U+uOh4n1o9TyyOPpBI10y97ovf+fjMX2VUm5xGD4bY
dSIVOuCKf1FZg7rIfyX0/hu2t+sMGRYQYOuKJdLKUGsSUn8l8qIs3SEgqpXWETBI
h6VGaWPK/tiUrHN2gjbj8TxdEaMGlGVLmEbubld1VknXbdl1t9SO9JgYQdKPoj/3
Es7Ml2QYslQHVUPinnbMqHh1mbf9L2kq9KaPfptYQD2C1vG3FI2L3Soez6pHwowi
Ovznpqg7S7+b5r2XpbiCGxFzLqStSFLDc43poyHxVt5wh8AqpPTUVHkBvn8LnoFv
ka4vHJ2bCWyySCIB6X17XP4Mx8N5q9gqLpZxYO+VueBXroF9roubwX3EjIWMzePx
zJTDOHsGKJxhswfuIQ1Jm663DChH3+hszL/5bg4Kw7WrGu3ZucC/IWVePQNrNarB
75M3eb0eSPrsqX1VQ2B8Ss2asdkWgUtwvDnEcoifyApDiz30zeGOHUHaNE5blMvr
4vfdPBrDfTr4/9x5G7VD4y/hoSTaK+q0nUSfqFFk9IfyLS7553WZv9QwFkA/MN0b
OeZny6C1drGr6UXilAQbzbMLAEmisOx3HcJRrmR7A1IsE7ZEZXIb8EGFLEZWluq9
NpMpMWLYk3xlx0e3uYXpDKqHe3qSoQHo/Q8QsejPLSSbBNcMAMkRREjXSrYUBj4L
/8/IbGboJz36Qu/H58TIL4e35ejNWXj+eOH7yEHgd5395cB/aj5RUwqnVYWBwf5E
wFxTrp/3Mem5sTpk/cfZLfakAaaHfFEMT7gEMml+AbfAwCwIilKE14u5FFUQdc4J
K8zm3y28ftUEc0tv12cf2A4C5bsj5Vl78Krpk+4fFrpNyryI7V3W54UnEU1463xJ
BryzOtuMt/zz2xhmfTmThANWiIq4RXjU9rTjm4aDZj6w8s9j6Ec/BeKQFJPV3Ngz
1NyhbnbGzorYk4NlygMsiTJ9mDCaMMTJuQjLTTyxqc/Uvl1+033gI+ecw0wDlAnH
DlhpBtuSA7OvtxC1U8ql081TMuBxkmarUdQ2PAT5prp8XHfllzTGDPcicFfjvxh5
aDZcd1UUq0JC+lXPI1buxXoy4rUN+N9iniktMyAIITenWWaj1FAYStgrIrKmIMLm
XaAVT08+ajKSdy9P3C+sG6Hy+GBkmno68f9ALcg/keYa8wJ5RxckIVoyOa6for7K
emZespiCji1k9Vh1H1DMWJhcj2E/fmDc1lzQzbC48SWMJSzFvUds9uuBsb3+wgD+
YGueBJPJ2IvZO8ak+gceOe0RBoEsHPnGewwZTpYSiMy/w7GD9zHlGiOQimgut0NF
S3eWlIv4Nn4M6SrLyhq3NwX3HrHLAvAq2VXJugoCokXkUCvnAOxstX8F6j5UZqv7
ULLBv1nAA1Ro4rBiumLnE91rDHCDLbDvTopw0y70+wb7jCfQzFqgjqfGG+v2Sh/l
UJa4vWKdWjJpaCjMO4DGnrqRHoDfgBl5ouBH0xOAMvwIcdWThN8eQnNqkOqJ9Cq9
WfevPqPSP+OOISN8D+qn+w0Oh1YvE5okym5UntnZokrJ6p6s5d8M7lUc3G9NbG7p
JCi63bbjyYrcJG51fISY8TNW1iZsGteCzjFaOR0wEdhAx508ox6SAEPuB5YPMGDE
6dy5p4y1B0eTTfnbo/WW8bBu/5QecusIJ9GqhTdSuGDc8Q0+0x0mMl9aRwBVHM/S
AvKSHZYS8RsnGnviLb1n1Nh0KoYSSE333x4icBDk4ZrkayfUX9R5OZ90lniqfdAe
z8IOtAOr/KdBkzePgJ+F2DjVez+A+U74wf1mWMWdy2SjJsM2hmJ7mNJSNywDlVUF
YNX6X77IRoEYcPzlNnliFWEo4k2Sc86JbiAvVfQqd3l71rsRoCG8qAp0Oa7waPNS
vVQEUXe4ssC/FdPrsMZceYkVG8jb2V5n5+4PE09MpfeBniUumRMGvSXz7yEavcsB
y9kPCJ3BIXiFLwktvf/GgEA8/tEpOAxnIQNa0Jo8Ru92ryKk4xbpaSMBEHLCM9zY
irSLxWrnl/Rl7RSV81Tsb6IpFN8YDGpnQFtOhbpd+LmslF8DKuyhZvHH7OVMvFeq
biroOQX5tSForqyKjZZi4S2mAoHXuZoeMPj+iSJ03Mnc2M3hvYguqP7u1O0pcHVP
x/W/W9cAW68OKws259ADEmH2zwBCaXtLjau5mnZT3cyagRot1gKlrvpwaGc7MN73
vQr3bhiuaOC+eXxmRgQb5Dd0f554I2oyCYS/UTfkYOYBrFy8aaNLYvKVtqBQwD/G
j7utKjWQnqWuz7u1qSdnhliSo+Q1tno/7lXV1duac6SduIqCUOx1rqM0ZZSBFyyt
LAds2KFH64c5vCFQu7axxb50o5OcNlpj3TZbD/B1JSZE26sUxNO2UWC9WV0KQ2A5
Ege5C45hrmRlnOZwwQrMtaAB5/DRNiWVM1lntYjwLDkbUyQG5OjTeRm3AhrNDPfT
q8h8nB7GT5IzV+Rhl2Pcbf5cpiUys9lA6fAMvbN8lTdazCaPwYl10LKVfDdxZEb3
E02ZS+Ez0w8o7DtyHVI5xwn7u8bv96GmlxBmZxq3Z3PcZ8txvmw6TfHHwcWn9bWJ
bimLZITyDDkw/NhgQ/ZN2FPHyt94OEbgEwzTXNYqwLjPtt9nU8JDi4H4IuJYZQyJ
S79XUlFYDxh2I1EQV3axjsbiaL375AkpPgL87i9B9MocY71Bm9zUe9aB63xWhHb/
91Dkm2i+eiFb40PXcvTYggRUBUyC0rGLb5NTSpvZzFcx2pOFEW9RP1DBQXJ9PiLS
C5Qxhg0AsL1Xp3XAL+ahjQqFvD7fe+p7RK/YZQLS4wJFnUDF9KBBFLu865vWgSrx
jjpkFYJ9+5p05WscN8p3loyc+NyzTB4fMOxBUo6hxP7naavzGj4W/wop+y4feMkY
zoEHvR4MByMGwSpgIY0BjUsA3TqUI2AOnPhUel6PxN7LUODab3gBYxkL8N9NL1//
7ktI3gHydbgDvnLrvGsl7YCllS0I6pdG+hFn/Db6v2XYNv+ChENvMrBwiVZHEDCJ
HtdiPb1q6h/pZXlSORVue3AEyfcVMiPDRQol8o0WOfCx1cgDtzRfGf/Sm4UBgrlQ
t/EeZ4rIhHUpRvk1GQ3Po9Dcwmpi+WPcMlQeGcJPJNhCvf6/Btpi18rJ4aHpJGPv
H/aegaMNu0350dlaf2M0qxUrMrW54fXAxHVFgCUW5MkV+3OENgRbzHZLeRFK3Zs1
ibHuDPNAz9pPSkgnIcfzhjM0oHw9CyvQloMa3iwcdP8jfyUG/awEntFC85O7cRj+
zFoHGfSHIh1LSTpyAuY7KhZWRCn9Izp8MLLWdMvYScc64KbqbPOiYLrJ5rXOmNuD
GGkHU6wk4qZfZnS+SC6RE/F4NHbgRW6OBXYi0DUuwrHnHA98K7uxZU2AMzQweXfj
W7/gC36qy+wBA5ygXDSzVHJp/bugsTYmnY2qbH3IjIyltPziWI989fJorXwR1400
J10tOVir0ADDDwCB9J1NSf4q7pDuuCOYpWRLTI8eCl9aD9GtacooqcA5RkOVnc/N
BP79JeFtbOoNJ2DEyvmHZ/zd9pLDu0bIgIAMQmV6BOubgWSiix/EGNA/4hzkvyzO
K6HvP7dxG2yxwLMstfj/rMztR67e3qGQTg6bhd0qSMgdfsMa1zaTXi7oMAeZByUX
n3MaMO5tMlgVIyyJdkqbvYkipSMD4AkBUhrjnjKtJ00BLt7R4Cbwev+b8hpyig7J
ljMr8bvVGyVSbbn+BjZoBD1N1TwHwruHnMJwCmKozA6QlylOgq7ky5No7Qg9ZxTZ
ECfmd4mAbljte9rTZkBmG80TsvLXULqeulLoMkOSHjEGIFPHJrOtuS+8OfsZKbPo
f50m3ueqq4TH83cknxLcKdhdK/A3RcrXGoFLsvJpviFJmXlfDwhCD0ztwfr/aga7
iuZ91mFqmBsPjU2hIEIikzdD6/RO2VaXh1dKIX+yfphnXiPRyuAFRcghiHLeNBoT
ea+t99BhLi2EYnFLwhUbBaAUAolO+lzIJkhkMejO6dxXxkBDM3cecoYipv/KtGNj
sZ0bwVnHmmDvt5lBZw38ccjNtx55VikShWoTwJhrzf5Q9++AoC54Z4WsW0xLyvkE
G9hoMe0iesrzDaAAZlyqVlLNFGA0OqbaaBJ/UxqsO2Wqp8TCUi0U6GRICIuHL3KL
t2RJouDCutdn37R61EWkfPAF8dnn9m3XSZH0zjF0wZrfuzW3pCHASjgjtkxkibuo
nY+r0GaGvICrzMLTrnkpU9/4RlWeRStkVZiiSK9kjuFjKHjQcs6y7Q7b+K5L9Bbz
pLlHFRtXV+ATPCbYpsVIFOvxzu+Y2HxSJD4WiO4tenUITfkQSzsubvkfgP2C7dAI
ZnPFsU84yWp++ztkdy8x08Zc+uEvmAMaYod4Z8VOLNGKaqO2uoJ9+WYExYci2or5
9RHJJ2Yyz6hopGdQuvO1KHswhhJo5+uJN91lqv7P/dC28ibJ/KvzduFwvUx8IbSL
Ir3+6eZQNKNMhH2bFPPcN830iKJTLTKdK5MvAizY21dPAENf5r3YHQ8D0R7wRS3B
5vzGTo0QSjzEZmnmIyIZHpL0678yD8kFPstyLc1Vbvus8xFtlj/xr1jT90vyx3Vp
czKE2+Ac7qK37JvwTBiWBj0Ki6eJo2ErRdj22XuTs0PjgwlgWo/RppZzy7iyr2cX
0ykcBIqFsgWOfVvuLdNxQSOVK4aUwK6TklEZODhWnn8nHPRF8VrNzHv6t3O11t5r
OFeREKW56dCnOMeCf7qZmO0YzhUagj1LfJYfQHROListXwE9Nw4eSKrPW1wXZ7oS
bTqReuxNbXu7dqeN5FwoJiqODftGiz+63L2MwlAdVx0oBckImPg8ZyCMcyH5OUqU
PimbAVFywDr6WfYjB7d+muU07mXtKYmqJtsRhr1/2Lp33tAMnVfSEfy7AiJGTotE
193Y50yPRJDnNwQNu/5+htSl4Kif2rAUV2JES6FAOnzp4UlTPT13EwhuuUjCnLxL
xTWRtQO1IUCuhIrTByshSqzuOF1Nhj+MbPIw5lIgJGdOwSoihRj/H4fWSGa84bvr
VMHm1twIVegf0BQNXhtLvIctDJH53jChkXLuHe+J6E9KFNJn9SeAATPenTNnBW/8
945kDEaIVImVappOYXSIqst0rFKxR9cn86OJsHCoWeusaTrEfR+bQ/fdeH8T0d/E
s80ksx2fQS59qNAAVUl4XXmFnnpC/dco8yopBkO6XluVOmEfjVQtpIIh03xw2bRL
or34GlUTZVZ6MewdPM368zLDyAGwAH1oSGFOiyrREa9rAip74CQiwUovZdn4ACyK
XioQWrVcOgJfGlRXwoU8diJiYV44pfqI2q0cO2IDX/9cCGwyNEoZ4M9rQbKp99Kg
dq1ccsA9K8vJED6dRZi7os0Qz82lwGpJfmXfnC4hPfa4+0U1DZ2gJ/PuDW0jjsmC
OFRyPhz3F+FlcvDXCSsjOIYLG9TkIW8q6WXUnEndOaiSWXZWCg2FI3c2a3Vx30yz
CjBa2aAw5coA5ZQglAq3DiKlp6VMGl2yYhu/hmGKpUvESPpqdPf4jSo0AAoP8ZzJ
3H574tqlI7t7jigqNlRanYrpsJ10aEsbZVuyhKuwZQyw9kb5FOZZtDJQdIA4vX1s
Ed4RknBVW62TDaRnsYbQZ2OsAMiNq+gpssSvsTIcOYzPA7W/B110p0SSQ0Reiu50
FCl6V/Tj0YD9CEcixR0LOs+9yPtk5wQfdWDUeKfDPLMnGZJ6IfwFpzpykLB9dz9t
KlEj2G007ZoDFqrjrCQGAH0QpxLmeSvWD5G0UWGKAIKAjlVQeqZAPkW3Er9p2D8u
5X8fqOkH3jfoyDOWSCim1xu0h0geZEAW7tbgra8oXGt8iImYQfRG2kDZMYfkdHsS
TRE4cfRh5KAog36pLBap2iGjBjCUU+vg7wixqHzK0+t6c3wN7RGs4srOdSbvmTLC
sC4Z8OQX18f6pDtNoaLTWj6DylKGyxHXiPqH2t6cqCiQJB+S9qMhPLSq2tUAcZgg
kL0KmScRhXnRaYBy4Zg61cd5j+JB19RtEixvLm0LHb3CZ73T6Z0kcSGQK/f8KxO1
1uSqoOELzFBIfHHs6OhLquz5mwDOq9EPc+6z+dsyd5+YqKbtKBINTzZfgkrC3EKF
zwOLQAf2CIvkHGErdPU/tsr3CbP5OWZ7cnrGn+u2noPs3f2a7hwfKEt4LVKF2mP0
vbYQ84lmYhova8mnVL5HAv1NhNR9n/71zmRMoEIshp2eyPUHwJmiNF83hL9LSqez
wulPBtuysQ4tEMdoewDrbT02TRHKczstAafJvr+1Z+PkVj+3aCgZ9WC/WKx2bSb4
OKzPACCAOLqEIgFJFx41ANFysC/BWZUfwM3HbpKuI+ZbT0ZlTLO3At2uWOKBvm27
W5l0ZwrqAeHjWXVhOPdExE/vQ1pXDKUmDLVqCeY8Po5nF8UFoCSctXnVBSoHu6ia
MmFrnYEGb4SWZd6IOU4zzePmkvv9Y1REytIvpSEuWLr1ZkJAo3ZLRrUTItpzAmlX
rR8hfZrYwsJrJWtEiNSv1/ykLwrzs5YwdtPOmdPJKufYfKxWNW916uhWtZTQediz
Qc1T5yiQFTlXWVWo4VAhdxtGsIcdfxXjLoKwY/JGGrZMEaYzNUqtlZK+6jVfU8CD
iUS18i9oMBxIkCTSumCmoMwc7Ubif69psEef5+wpawjTqh+mQmMzGsTb6GLAEdKA
CFuVzMs6aIyu6oJGzJXY5QVsRqAVAguSLgTuO8Q+Xv0yhDI3CLQR7DdaLrLjkEAE
wcC1iukwtpAfPfOS6XaLvAnRffSSDEzzjFy9MEgq/OMiBJRjM3BG1ES0vOsQ7ooN
A/gH8ZH/XSczDG1pIOwtchWASUy8UajiZxoNWFbNvNrsqc+gei9cwxQGdXqZnIwJ
si2vbNyiK4aVFYLW934fenMf60pTilFIv8a8opL2xeHji0osFxNxfU5X0Z09yM6v
KqMh2ICnvOnPeDo0Z+ABIJDmUdj+hsKpmXRPOeyo0Gjk+wyCdj7ORrpUppYPI4xe
W04W7Y9JZbhoD4jHJNxw6cYVAOvM4sarbwSYnfGVcqmi1/G45obBYnTaXJpUue1k
E8qFhWXZtQhUmijKw5ViX/AJ52NnfqJxn3DWaHg+XKURKSobiy8ohsoG/opO1+eU
GwVubfohnIeH7bKolj8N4xb1c3/ogMWryf8RV+PymAzITe3o2qfCuEXqjLQ087z5
o/OCJ9iXRz+7JBB3bJxy1GSXeFvx4ZHzImSE0R0Yu3SQcViI1Z1yOTltnOcvWamU
SzNaA7y9KM2urRpYLbsYAM5GXWFxL+XIf8otAFTnl5mCzthjApRkHvSeFvVLE5h6
K2aW6/jSeDiwyj5UI7PhICWnKoaNGfXC2mg79fBVVrLMmztzT2td8gpb7LfWrL52
LApkFmqTZEJVQnKyF/tC2X7e4ebDBxyQR+ad5AgMFuiFg0VvKH0RkhjN2DWxGEUC
gcy/oi9ykHV7VdMXhAIQNWdUDPBJgyuJWtcYdAP8MJCFNVb8LS6IfSdT/s9C7NXo
S3h2U3GDbGn7pJikGBsPvpOiCodiFT/ZE/RB+yjMRHs1paSd6n5uE8DCPVy0B031
XMnCIFbKPNjnFIn7x1LHcvrwjkYnKd7iWvE8cDc5z8e7MvhzWnifNtf2lOssZCDA
Ho7yIlmQ7mGVFaWHSKPpKGQysCtQzI6OKyUHZSu3MhIlddbon5xcPZBOeZhijdrb
WKwsq3ieocbu4QeAsHmcy05h/H9TGqbiKnmPNrwDtqRZqIpOKnDXWUDrp0h4Yk/B
pEsPAsM3kTlaxjD2FXfqLzr4p0EfJRwThL3wIC/uZS1vsuv5enff8YpYFlqPLzam
nxLmZW6HeCHxIO/TDpzOl/p/O26E778tpnx+rKF7YVQCdEnf/U1RotMrsD4mgXe5
513xVgfxV7nQXWiguREjnWOXAYrYxIvmHn9P8662+YUmLeYqgZijWmxvBsAnY8zp
PUKbFG6UeoJ9cv4/ySOrI1YYo6GUdSlMbtFy9Iv1jiEzqN1ldudvivLvQ4lJWkk5
IezLgF+rRvpwpljS1y4MKhhsskE/yX7Bz/n7hqEhu5797khNGcEmfsJhCaHbpol+
q87wo4WascPk8eAO8P7Q09fYOEQ3Kokj9gIusLPZV+iVrq/ngZJGN/Nws8y0qOpC
K5r/BicM11XK4Ayf9TUFvsWByI0/3AdZ0Plhsts46oWiPmTxpDxyNHmplm0Bmhxv
LwQANIyG8KqXey5qxIpfTEzOAT0S3OWBcn4w2NEa9l5TN7+VdJ3Td3+INo3O12oY
+7ZCD5ondjGN7NHPQckV7Tm6u5+FtG8fGmiEupUqfsRWcrLlsUn9a4kL4wdy2b9N
DI1/zD1MwZQYnJ5EIgGsfZOdKRGvs/eLXjHZBRkaiaMxAEfoAQuLHzJ/BTlWVgDd
CqracPzZDzSZWt/qzRaf4q4AD/R6z5y/3DRCM3Mtq6EqiRzKod7G0drUGYVChid5
TTOqX6nVxJ7+pUth61PJ+656nb6D17vOPUVnyHv279/yqvToDDVqLKmzjAmOAJ/6
SCI/+xQCYipDHdSzLVEIxwMvFx3E2N1IQncf4zQZOzYCgwqW3SutYI1eUU9+5X/B
7BroD+dx6CCC6LCe3/TIv9EbFFxTKI/1gwEOEeTbaF1e66tO3+fFUrmOrbQRiccI
q2kOi8XHvKTH2mDQkgXeCDlLw+ugu2TpfBSmO72aD4yODNRAGIkHIZHxs2TnmLAH
ZYLQ2AGeNFM70IJj3TZcWahzRFYMLdjqVQFoJsJO1v8lwxqrVIZEjCGpgvbcZYtk
ETpo81uG3C/1YTv6S+caBuM/EUCSGXMwiQxT7r9Av7Nome40R/7+YthkA9R9hW0A
m+0rtm6KovNNdOENR4h+NkybU3vPFTnsGmjT5Q/QEaYAzO0NipDd9HkNVmPT4ZRo
eoEDwHBoxq1rPhfkAcY/B237vRaQ7VNmIk8WfwSiL9UFcd6rz5LfciuBuUSLwBot
tSpHGOlgUUkRy0mauwrcAHxRl2IOmOSZGWDNEVqOe2m99T12zHRNcz2EipWid9C2
D+OgPw2+tXUbm+0+BvVan1eXkj/84wVPDFY7C0/8WnaecB/RDXnPrtOcvmBRFWjX
oPgqNOvSbPiUgiTTgHtYDz+xl1/i/xq2yiXURY+55h3itSPZxQSCm1vzkCjOnuHu
OUQcc6Bg5LkOWQygBQXHsGwdpKLW7TrY5QaL4UJPriv60Suz/XXaH8iB0ZmhqEGp
6hAdKuTtYZQX+1MBjvgguS4IW/Zv+Vm/Rh7JTqI8BdtX7tM/RrvghDsxzAal09dB
lw3bSaozNa/NCfauqvE9A9XZU0CCFbv4BN7HDOcUo9xkOTe0DZScpu9uwTh8OqCF
GKkoYcQ3JZbJHTsG+Q+NR5zLjfWA3COmX+1T5c5M6khMK6gx8MG7ABSGLiA+KvL2
pcf+7sYLZvX3nWTCWwfQ7ad1sdDVKPfSnNXIH01ju5X8Mt5pmIvv2xFY5rFh1jd5
k64T845rWOAO7CQjVLo6acp9yPOSt8WbgPsmOQ7TgUXFZsfFC1tBK5l7c9ZM5Xdj
2wYUEBZhREzuM8fR5O0TOtKT4FIVSEJ2n2xGdWYjfnf/+Jn9BiGH2YV6h/z0OhvL
1XK9yffHxry6nK3JMgSVWEYT8Tev3lqOfE3H6YOvgWsb2cpFqQm6Hs7h3U6Um/kv
0z7UU1A3iblc+BK7M9UoDatXaYSViEGDcYigxq3S2iwtH/IfjEXvAkJQKlNjhjOI
s4q4tkGPGij1eZQYRLurXQWZnfCP+dMRx+YthhCrnKIzwzRTISG0PYg4sF3r+bSH
HcaxH8Xuc41nrSrl9pmlvqvX9k2Xma/0I/EVs1uaS0R+ic/k+0iC2DKsHes4MXkt
7X5bnNP77YpKZz8jMReKFvzYNYEfOhctEXbF6LSlD9j8WUwWisbVfdalhsuHROGC
SwzmypPwENwzoSzF29ymknxGHlWPbBrgYxzdrvbnckMR98tgVEGt2b4HsAlqYiRR
FagII0tyxMShhSqr0X7N1neAD9SHJphoSMhL+ddHGUx3NnoTjBbdjlllI3BH672b
1XNHcWJQMNVfhePo9GQvAe0xN23iCbkaeZPlVVwTthyx3/xcqDBh2nRLsBNcMam/
2AxDZIMeSnTP6oIiRQ7XoTvPYD1SNuBymG9XWMXubRcjx6UpA1s8EfOJ2XEPZqha
rgTEPj9rOEjsMRzyNU7OPZrbwp1Bl6obZqL2mqtsOpRPLq7y7Sl4Pxoky7p1UsOz
GoT+GcEk8FN2+HrBaetpqk57zL4uiqFTcnsLEo0m6K4rymsBXD1gic2vSuaeE1Lp
EYDef6e5PxKnGFiTR+emezcZWPIhB+YSX8wCpDR6SwSx+5SlICKVtUltaUkwi4nt
pyFuKv6bsXGQjn+MXYxdcYDPp6iiurDMmsKYIQDRBXY1gk41l2iVvlZuMT1qeR2a
BITA0JWVGewK2Ki99QQnk+TH8iGggc/6N2kWcN2J5fftBY4NlO9o2IWt22NJACdA
OoRYyjCQe8inrLv+iOHjveYYA0/TVhDFcMaH/K51P3lU3SdXEGIYNr5Ewm9fbz4O
IFZAZZIaffWP8IsagONzbSEZPC7r0dmtLngLz46OaZqC2B4AAoJG/v+UnSLfiq5H
UbgKWlVEpRQHdS7SkzNCBp5/KhCUekQH2T4PowPExRAlQ9PwzFreA+U2uBxEfxkg
TeYHwmnmUGDBnQ7OsELEka9iaf4K1D3c9JFB4/tT4Mxb2RhbK7Ho5+9Hc8Wa7Mfe
Ych5krsi9mQRvYKDItGLdcVNui+5uWG/9aN1LA93fewW7qYPZlq5z/H4mlimAvMI
RTt3uavwsqSiD2s/j3jm9NSxezEStptdplvZUz4Y/CslRjWu1YIJzO0YuLXyLBTJ
OZNHGNPJqjjhHAVoPyxDZwWBnpMk/cfJmXNjLNaeb26qmA11DFtocIVgja7+hA7b
ljdTOKfNJgjGJOPXTiBZhACQBZRVDbK9YJeVafrXrgd5MXzLuPkVYYkvyTuiqhQ/
AyjOyrhkdxNK3L8sCj9AI8WG2Sdfkf75sF4dYJagSNk6T3o6wACtXVmF2Ckv6XF1
1STyLBmQNeIketHZrC8zqcW4Y+6U/byTluorFxdntjx/zcnw93DqoOvwCy8PuxsO
j+IiIkGUzQSyasaB/eGAbMacyveFYp5Bm8uOnO1AO/JeBnNpb0wpzWpXOpEuI2re
gm+I56kP7s1c7co+wJzMivR3kJKc8Vw+a5vPZL+HHRqMU45p8m8sYJLwJ07oiNBQ
UzBr7Rqp7w5TQKPiHoJXpHrp0kZYBSYmErsxGsfeyRhb8O8eOe01cn/w27Bxumyx
dIZyG2LQPc12bU9bktOlTfEeuxmpQhG1AhEprsfWxGNOBQSOCcR+seBdgTww8Hyq
iXJ8nIdiv1p2eY4rQHVbzi1oOOlCpewiiWV8/Y/7raIdQgnuW6gSQADSzOkv/W+K
i8jLQC8WXZq6nV6MlZdgn0R2lvtsrH4ESsPBdyUlQgLMnIcMF+Or+GF843cPVnC9
v6E+bVYqD1ZtrvWW/bV7mjjHw6stySFboFBRqnTdDfdGMIcrmfmd23PkChxiNq20
TPr2wY/bQ/qJQ4ZPyKp7lwYdaGzU7HkG76klwoFOx394yIOIA7/6avBHV54czAT2
x159mVpR71HEoC6a1UYsSZiybhqORGmkVykkSdTLs5YIpMWP7m4mXKC0mVVbI5iA
r9BNuiKGtqfvfWRPbdZn+N5NT2je6IMC2pdN5Y1l79tyVQxwFx2dK0+C/M1U24dI
T2JKfApkGYTYdMFTj2Kmt0UmEbytGBCXz1GPbVBxeXEliPSLxXDFOx69QattCIOf
ddC2oXvUNDayh/v6P9td2DUBHcazD2yaxBrWDa+0+9UWCAIqYzVycMjE55squpDO
/ywd9qisoeGYHlWYWcGjGolvIq2A4VX5KqEiMV6NXjv1SlppMNZAmTggsLvmsFXL
srqxxqQ7Uer3spENklxwAt48bf1dlIYD5BKo40cOhzO6y3HNHlCWGmCNLj2sWuq4
J2QFfty96pRvlPeDMaasfpNZUJWG08tXxFuzfEKwwFqlHYa3Q8WZyLVEM13Zp2xV
7bFzK2Nuk2M4Ec539deyoOwJvVaaRPAF5Js7FYna9LuEO+D2E83Bph0uEnZ61L1H
yiX8GLFTGiMdFEaCIzutZsfoZyqlqlycxt1HhnazoK9e2jY1Pli1p2AznXL2Ydx2
e/XYHs+et8s4/MkKcKTjWzB5Zp0yHWFZXDMNq6kKeIWuJK4MsGt69pGgze5H356q
RAWL2PxhANv7n7EaljwqqMAL9XFFCuXJZPCAWWyoYwSfXEZzyxyL006qfqQ+VHqu
3CUUAVXfWPy2FCjG0iKkn8iTGF9aZ2urtn89vwl3zLTn1vsLdKSHbEzfmAgVW7f+
XPjiWUenKHSk/UczGc0mp1FYjIqUxLPEOp+kIe9w+MW6kP7vSdeR2XybhYpcc54I
Rv6Ficd0KoZBJ3I+lBPHK4V92ey5qBhIp0iJqRC5dQUSl+9EcuOOtXh4ldsgZQtP
xIY9jH0VHWMYdHlH7ZmW0uWDNzOOVDXlfXr2QI6kg1xE94Ep1+n9NzHhIxEdQwRf
rb1Quib/CEtNFUlJFIPWkInfO3T/wYAqL8eVCknhiy8Mae3GU5lkIaoorPULiQ5Z
jIJxI44cCD5GZI3TPrIcMamqjaZliAv6Pe6/MG6gEEEjYLPkfXPsELkmswByExI2
ZeRflLFXaE/MDe2NRSx7qOaPQNV5k+v1ZX5J+vuse1Y9UAia1dyklumqqDCIjcxu
yGToONZzp7/37IjSsJe5A2OlRRdYx5d/ouFVnl/DDQk3rn0/PbN9uKaLOF2DP3tv
i2YxbSxgxKdLubpA+yqYckwz4iRa9c36Qkxp5mILfJR7lEHh5XAeqXwHJq+JMNHt
GmrtDjFYKBaGMYj+qp3/RYe+4slIjVEqsncOiUhocELdMAHvkJTXT16bzmrTZ+B2
pf226yEazcn5VhKVDt8gqvvnD5BEjVi+5a7NsTikYezSJ/m43+22LA6HKVqBTfCX
kESjTdYem5nA0y2DMssHyvpAeLVGK+J4t3rbp8memu45EXuMkp4WgIO/dJTfCs8P
TG8k0jSXDa/x8EwWB+V3G7pRJRIahlbnUw5aiFrEiweaoJkDEYbuDbDKNJ00hGuK
49/20S4g0CZwLKAPPbG/jxT629eWT2RbBdk0vwxNsj48zBUkE8ngd/1xE1e9yvQ2
cVof7Rj5AMVSCmK8ns83movi2p7v3v9dT5G96AmtOUp4MloRPz+/3Miklfszwmcp
HDWv8hA76S5nefuHJuBe9mmHW+sRXkWxD99skKHGAFasHF0b3YtwhBWpjSsfhkcH
LrnI7xOHaQCm8Npj9aTVGL/Y7sdz7rsWrYdMepdMREZoFSvCShm7kkR7pXhFvqii
6zZt0csGVcVdqp+36fveHF3qDizoiJRH636Q7AHD/LHEkl0RgVuyomu5b863dCMF
qAufOML58Y07WAdfg1jppXgfFei7MqeDukTZ6oYvBmYbQoG2o345sUFgMFclL9Ik
2LZIbQpNYyhKlqJPhze2IT/MP5KnQU7h0xvhqxMsZNT15PEYuI2cBC5hAvoqTyF0
/uhdpWXNxfBoTtZwR5fdSH5W858v5vfrkZp7XBh1+pdzIBBDy8kw1tsCi6Uew5Lm
wP69veo/yznIB6yrUvUIxTLluSN7v5h3oKvp0294vxrk48WyxsGmLgS1ofQ4uUQT
RjiUVZfrFY4owpm+OVJkZN7OIVxltxEpvGnaAGFuLMK4t9XXAY4fhY91cMHEv784
T9GwXsDkzmEE/Zqp4BJWEjrBY1JlEpQZoYZTJ98ODVkHfVJmfFMN6q9on1LQ+ShT
PeHE6RaWa7qv98ScQ0cgQXfiVNQ5+tTtgUcCM+08K4mD7jY3/84gz4VKsi8i3RFk
iu9St0g8p81GjHBOyJOJy5fC/FgS9RGx6RtfJ2UvmOMDIuAe5aPVcDHRq8j+0wbI
bFTU9R+X9R4wdrUEYg7klSdrlMujOmukGgeFDE1uUAHV/2mqtsIG9Y6YUHzRq691
e6koAkDrhnWZXCZN/XlU/uEKU3FAPD+XQQs/jQHG6DQgLzU0+ZYxgAiH2PgMt1Yz
fqrTtKntWmUd5FvtAs1LH/154ccSkua8EnAXIUF2eqs7k3Ml0W5kBF3AVzVvo+kc
Kzei7N4sSERVqSpcMDgO2D//49HAZRQlQ3v+PawY05OdHkPz6nbfk6PZAYU2fLHG
YODHsJys72sbg0HPHjVra/5LYErqE5N6x1O2b+xBeuNsnhhMmx0WCkFqb7M03HoB
hbL3nWOSwOEZAeFKx7Cpe3aTIE4tp/zP6DEOcEXhUky3O1wMvRp2GQAhy8MQUEtx
s+m7LLxBxICXAV4Md7RJodmqsv1CyxEI0VxeqJV7YtfcK/Yu25YLQjm5z4TK9kDb
YPK9jbXiZiRvZZ3b5ffVIQSn/IifceZQ+ZbI2fqQpRcMzWX5yeVtKsYFiua1MM/h
b9AuXEaFYcfGyAMWpz8bI0b2zL43m6Zd7dRMk/Mr04IAFQlauz9SJnk+Wmbyf9Ua
S8+Z5xXfx9S1a6aciogNJqgPohYxGOflb9Hkt7Dz3570iJYVmhH9OYRZZsI4GuWj
XmToE+cCNWIx4otCMrqh/jt9hFAigOeCncWDOmaaYBQq6pLLM67TTWB1mBseF3wr
WAoDYJ/77g2RQvLMKdrhCzB3twzdCruRCegmRdl2bn34PvT/A3phn9AmqBxYT0G+
mmwwkxj6nlovpPmAuy04WFNuSjw27QPjtNzgEmjp/gkHwbrVWS/LiY/m9WtjRle2
JF1OLEKun8ajbIZx51hooolhfEbs2Ip2rSi6YBbLZssnF8nXbDAwZm9m/ef/7W/U
aaEUCkUoBHkY9+7F82ezZF+BQWB7x5YRM/8tgJMyIQhPX++sa4Y4hTf7ixWQxudW
hCYqJA5BC14JLbLSjuu1RS8/2wCVVTJPYyvudOZRQcJ1xB1gb6oVc6VfzzfgZC1U
Nhpl7JR1biNcDDYyz6yvBhvPCSrgqXGeIuX1h7AhWPMTYxac51ZmZ1fLwKnEVKFm
XhwLkE3mWi0Mh56RUOCtRVsltkodK/NMGQKNx9pqoVwmt9F3Jptsiva7h9RncuCu
inYojAwgmcY8ExNYfq7ClOROFC/Qqj2pXfJeWfNu4Z3UQULwCz3lt1UFz9F/8dPD
Fg72SITOMXdaIHku82P6gdInIc1nrXgd1WLpty5ta1cY7jQHDL8wMu44vPu81s1W
5DVxTw1Vg6njp03dUw+B1E09LLLsNZ6mQNdFFZmf2siWoQidCZ41cOHqRBsPEOgr
qJk5AHjyK37gZXfqiGNoYD0Wday27iKvuql3xT29FodY0U2rHzFuGsrMx1SuEfQZ
gZ8G9qWA3u9le1g9xzZKSjxaouv0YolNc1E1aZVD8NltrAcdHezfD80b6fFteRkY
nt11woSdvF7v3X2tMZCJnc/B6TUiIZYcscJvipFjATyxh7fVWyo2juqXJ6TAZLKb
MA4IB8BwSuqfB4uePzM2BuEe4mz2BCDQHz8zI/K57JGWXRzo0A4Q2yxNHyX5xUi1
G0+kQCzTfQf5LWF0te4jRoQNok3dM1dfLQ0yzX8pQUyVlOMf65fGVMhvz+PhMIO1
i8mGEOnS8vPgJC2iJ00t78Yi0ymClEdb4ZsdqdTZXaQU/8dBnEOaIxpskgimNvnp
mrfNWZoT8E7BLmAk0bqLaMLFFMHssAkQqz8EFRIv74s+WXBNb40wlvZv0RdzgAQh
ef5XYWC8pKT2Yx1Qn02FFdOxlAb2lmfzuVT0ealZZtl2Xz9E0KvLqs3T9yImJalA
PKXOtUwSkxJ2G5GA0aAOTgEfqBx54xonOHoh1ZDl2ACQq75Ex9rbMYuyV1Vr6sGb
CLiKrdHPNjK/NHdt43eWKxu590dnY3PDUF7YJg995WTBcjuastyr7dia6NAgllqZ
2HYIH+ADj7thpfdL1xz+PmcBmX/VCnH6vtJDdj4Ytimk1hPtSiZHQAmhzK8NP400
dE1n5064BIeWBpe0bVWxrgOM2oljPqcdfk048A4EAzj2tvPu1NplNzT6Ytd1+11/
MTgzjty0/87JN/bdEY9J9EV3SKngc9neoopcV7lXjHTLb3UEUYE9U4ost2aOfqzJ
OVO/l7kwMSxmn2YNoLykiybv/R6twsbwkgepzd+GscvuBmrXErcSaiJxyrLoEFos
ZWMjLasT3jOlkHE5rCj0DjsDAy5uTNEp6Iiu6TGr3R9eBzBGqTNUfSHokQMntPpr
XnSeWSODnr2SpPttNVY9rWvXE8vAXBtRIGZ7S+W/RAVK1MbYsFjgt0cRsgUbccMT
m4N2nIGTlyGodKzZqzp60XlgZirAm8uM/CGcjXlc1ZDchXG1TLSDHnm/SApfBHQh
BascdlBO24kwu18HN8C99eolNgr+UcNk/ztV5thsmexMYO2+lkm9xBCo1xaXqDoh
EDJnNv/m2ZipRsn3oKn+8XCd+blcKiBOL1CsxJv47mo3cmACT49OhxuF9voQlkQ/
jEZzCuUPuAj5uN+etUO9jjpy88rFbW9VJys9cBMrp0ET3eRTYKmILzdEJ8FCSUtA
salauydkrjm09jSBySsBRs3SSFRe1AEl971dhgKwMHZm73Y++WBIGo8zDWPGCugS
w/OEtItX+ItedoBv1rqBdOX/s8gdIsWxGHGPkJJc2SLaZoZaC0EjbRJDoQc0K+/L
OofdaVKShfQQZBinquKTrk+gE4IoILurDMNr/An1ORuMSvixQRUQ0S2WR2Fx0Kv/
BpwHjnGDQkkEkG4QOghSB8fv/VP0DY185xnLki0G691V0enDclcXcZTeSFVjhyYx
slRj35bcpZYDKKN7RIkLQQp52lfx8rN+RjGxwoAMzSvOnJof4AjiPNlnU4I/tFkA
FOrlKiJSFrDiSC/o+9AOisxSG7iwi+ofUHUkbZ3drwESAo1WCH46fxuDIElJaHIw
LQPXwn/HoCaFz8kIwGCdX1RX34O6zayj+VZtuRUG6/a4OeDFBTvYNq4ZgmnTnzBa
J5cyEYAfekfrVZzDRvBl4lFO+NjNHHcuXGys+tV3Joot9fcG4Y1DID+XJu9Wpdyj
gkm/RxQNQx6OY8NkaY4Q4cs8CFX+STuU/RD9v9GYlKAr+JhJ3iuMtrLd5ehbUN+u
o6aGwn+cCTBoCn4ZVfsXngJGbZt14TQSfRQjvhsV4RpzhL1KC8n3P7HW1G07zRIS
/Xdnux8OQkqPn79FrrtwBIX+IIfl9s4Dmlx1iVcy+qrrHHVjsFsK3hujAcX436aO
j5nYZPZ4mg66/33pZ89VQeR367L8e8M8ynTKjVEIEBBPU20yrS/T2PYYFjPopwQy
fIbHSLIvykygf0IG0JSxHn7Ey7J4dNlMq9qoHYnCQvc1UMQQMALGnRsvm/gZ1dH4
31QZ5rC213bf3lsdzKvXup0/WUjj7Nq3EiSdc8mGTv8Nyo8ecIY5UvtTbSPbhCfv
0Q5ZxvMZei5lTJmW5RsBO+E1L3ATHHAyI8o0Bo2KVPI5FgWV2q3LOIfmqxg4XaDS
a4iFB3muwfifx/qy0JuqaXrEKWt/YuKEfhhhJayefSUpIqZclOuUKyO1LCpf8sdO
HYZZ0P2amak6u3joM5HqXuYAQCIfqRREMV76Wvqr3ZYINvX/sjs6SJMD60MRRnKA
7pfNB+AiLeFH7Fz4z0RRQq9hsv2yQ4AIqJqPAetE6omPj51MccxQofzfWWdBxd6z
TJocbU4q/qi2tBpTBfo+OoQFDnUMAc/ARLPYMGjwTjc2xdSHmoCz/DGJvnvk1WGj
38QrSAwLZupiFmzRzHdmRt4VDG9ChtlorQu+npygg6mvkepk+NZrvnWqUNUYNMHR
ktoZ7Vm7gumyJYqo3y5tFWTPgFrRRIMFckY8iok9EE82urudPH62MCA7E150pFDN
VONlDGH/S2v8puHLHU+1oF/GTJ+phCqu/YHkR1QibUc1/wENuixVNEIEFojQnRPr
eI4jMAVVml2BDY3UG0FVkwrVqfDhhEiI6Ss2gVmjEcw/S8AojMyreeT9NCePRK5M
E1/U9oImY80ZIZV4sCagVBlaxu0KCGXNj8fpvJSznLmcT/pFymqRfiUQHGQa32NZ
UDZzTHaCHrUbjCFOdVHpn24JX36rBma1sjwY3bRcTSykXh9LrlfLPkOmK8gFzz/V
cbjFvjzmKgV4NI31QEmu+hmiam/wZRCDZxtfwk0q4YitpSxKkvUcSNajdNshLCTK
nd8UHzQ5R36JiiDH3oEVMu1I20eggopYd0W1nDOJoK+9LK1z7DzS54vuFrZOiBa/
f60vDyuSx/7uhV+rnS3tWW0rOM/Lyuj8DojvOTrau8J6POQxDo1aHTdD0+xiAtSS
C+pLru23xsP8qQcEfGMNi3/TB5E4TZqEH76WTNNfkezaNZQsGxXuo32tgK6fE9G6
k0HDF/MFrNmni3pSSw3r7MVP3u0mWlRT3eoe7y5X8SHydSY4t3UZ8w+ABrNkRO2m
nubZpUy0+RXudjDZvFygo+W1gSYHVP6CD9eMUn7rTVCn6+A8PEd3tCY//oSsoBlj
gso5sjglmOD7WGMR8gzs8mo5lXPzryeZQy/iwR8CM7M51HaqqL0vUWj4FM2cutZ9
qMfutmiQYmclA6l3ZYq6QS17lPRzev98e4gvHvTLbUZ/YaSMd+/j3B6i5F8KTput
aRQ/JYz03PCDbR6zhGG3ia3ZXZ6A1UwRGp+QVhq9DDZbn2SUE1cA6QZgL2nOJKkQ
UrSa+szNTBNbR6T7vwwG7yMySXoPv6a+WCGeMGOTI5CGe0fQvUfeRhggErdXYauv
xT5Lhasq8wNpjD4pve8YrdJaAkN9qrbSpuXhc6ujpGgG1Nk5tG7bGzZ6j059f7WG
z1w6nrBkzefTzzmkHajkqIXthQbSm98JZLvhpQG3YFSNSVySUu53WQMmCNMWEoPe
YPtkmT51ArRpe4Qnr/f4UdXPvrlmkYypO2Ugh86BAg7Th5SadP1LyW08H5PB6M0L
0yB5kyQY3Wc6SHlVLtJOW9ez6jB4leUOBtJxrwrTGZ0sZrUV8iqVBxYm06Ta3wzk
OgQLyEm5Vihvv0Syy1IrqEj0kl33YLGJMg4KUMAyufd36kFVcXlKRJy7uggdytUZ
qwv7WeWZT7E6mRM/LneslK5LCJINC1SQ79qiGvvz2Gzq+iTyanuHobnT+hNpZzYq
0Ke26xPI4a/L/Gk1ZloemCg3BQoC06Qp2IjpCMRcpD3rig6fSzUSxrP22mLOkykK
Hqdx16EaWy3y4zIiwFk5F94GvvYUbmQhIH9CKhhexV1Hb3c+tau/3ZI5v37A5rJJ
SlpRnv04ljmckLXmd4i3UiQUmT6R+FK+yKiCjcQzUCAV2ZDmGSwAFLduBuYXSu1N
dm2btjYbDQwQ142orfU/mCFlMaZoCb/0doYUgp8qt9v79HIMUkYo2Ls0wP+Am7As
SbEsZ/U01Jv/AhT0bLc0xZ9dbjCMINVKRmpa9cR/rE/jkZkyZbVEroqphPvPGv16
CZ8X6rXVX3ksQW+pYnGAYI8+VtFAF+XHeePvZMTalewa9QMAGwjVRnkw/az08Ety
mpa+GZ2Kh7jYm3O3i2TRZ1OiF7IRlqQi1MUFmlSRJHbBQiB1/5HVglTPVt+6hVBa
QjogKN1W/sxaz7IcbCY2RpBMYiqBx/cCkDaECqq1Cuq2ARKb2PyfdFjvkyLRzRw8
OAlADcyWvXYW3ByxcGIr1zA4GiZCl9ztNwRG8Da0O94nVz46WCHZF60tmyW6skRa
Jp9WrmExJYWxs8MQa+rZ1KAYHPkqx8+N1y0yRQ3q2LbNrYQCAB+eHw+njIEIbRW+
I+yRLjzlxS5rQw/f0QTPLFFGJ5fmawx5S9MkwCjNgrk+hv/CAtzbdZ+7WSMrgR+a
V9zFKogPQQzS7ZrRrgOPOmBGHkH5KubsB6bnLTKIswlacqSshrs7IskWmhOAkzND
K/5YvA7xtyExGYVfuY+zk4aCuctk0mbO8STuDWplipSmyElBreQQ0+0HELMaQaIx
4ByGeHYYtpQlZDtibY+jLiDT7iKdEFvFihtU3bDfT2/QQ1+lh0VFYkPlCwUFx57m
I01Px0vV4gKQ3x1ebvQ8zSb/OOi8Jh7Ufp+dv/3xb0KKoi+o2T7McHLkPbM1EDgy
Y8FFuGqMM+F0LdiCiQK6UO6y9bPLN8NgrvxOGrW5WOylH4q4l/BYbBPmm1kGppHo
O6LJskXOoKOVwKRIgplO8iv77WnL3JELdGQ+dzs1LvtAiNEIde4FBVKYWzakG7dC
dz6jpZPKb1eSbUMngOXtZKWh2/D1+OSxR30Iy2FshLMh+IlvaS14sGzazLFLxQHr
4/X/gbN3VGXRUOV0yxawAbXgB6byLIinG21yWI8mSnmaH/Hmu9a6IB+qMWHNsTuA
DRU854lCDSJEk+xEke9eFxBsAaGKqMJhAYJ4cvofkLAdKQVko6TXEgbeecCS50S2
ov89hB/HLCqRUnjKooT1gCOzSZq9MPVs5DTe0imxKTUFuCZkGQd/zupDSkoA4lHT
Hyu3gn5ahG+ye2iZmVWJ9x4UJCTR2PLCAqqZzj4Ka67WnyB1MjwBavtEuHFgnaIr
tad/onqsDumlaK3KP9Yhpm3X7bxh2uFFXMSWfsPazHcOaF6UG2D1A5gutniMAaAw
NybjPRrRMPKiR+xC5JgTk7PHBnYyvuR4TN8y9GhhKt3rj0NRAFthpeyNt6gAkzjF
tCGNPMQZptEj+mnoa0o0OhXT0Ob2kC3KmmxW2UNdjR/kzMFQ323+wTDXwkQVhfG6
elZ8Yl6qju2DbBTbuGPFmi2t/wylHcW7cN2SQN+eFF42Fpf8D7VEQ2tG2cfeZQPZ
qUdwvqPj0zhjmEE3xrPQ8F18Qk6oqNEtCSZdI/jZO0CBJe5AD7uUZvqA3YMyebdi
5/U67K5Pd72ArzeXwvQBSWYoY2wJSJOGP0nKcMb3DVW0ISgmEdq8AeD67cH1XCkR
ISsq/V7qizAslwdjvrbIR5Yp5my98SNYVjD2JX56Nmp8tSXu7J2fd2bmeU4ZOga5
I69QS1VUcuALusJFzF/zmMVLIyzOksmvB3KgQazblMf9ZfN2yJXvKiKjzq+rqpHt
BpvaX8Rie4zWUu1Aw4q7IvlN2Avx7nI/HFEfrp4dF7wFCsjyVn+Q+j95jCIh26z2
GnFIG7KQxHWhv15tmQioGyAgD0PZMDpw8XUf5yNpvkml+gzSOwr50I35M2pOgjvO
lz4pRZ9BSAR3fVUPnze0zneDAD2PVHoog54zGYcXwzmgoJEEHIDLOHLFEmUH2lpU
h9zBRftF8gCFtX9sNVj0Qr9pnMMNYhhe1FflLc8/HixYiq88iaBxyBnmuPN9wOaH
4bY0pZXvkacB4F35y+NGvAIA+GU5RPshgECQdpwEZu5EsIObvyNJKQp7Kr7uWN0c
pCTMCalXK0gSnq6hZRvkzBOv1qOnEInzcGxqsSjT4Kv62Tx3Dz+zdpvl05F7GZEt
R3Kyra7J9layG1wN31P2xy8Y1sjMFzeVeiJmjKI8nqEAzPfz9evvCm3QV43bAzF8
ZflyVCrlHCq3TozYtUWnYGDDT8lJhTNvOkDerFdRWzg3XE+0qqmY9UkvYMu/Zwpm
VfqRGSNxodG41bb+L3prtHqZzD2M98ZT17lIarp/Q1ZAOwST1icthkGUEThUJ3uC
t7T9TSAlyrhGBja0BXIWLG99W+82kvBZvtvruw35z6nr2eGnFsCrFZjGpsX94Gi1
B7G2LkSXNrOMoHrVF1uChItilmeN6MyHHO2iPF4tsewnmKoesIh1vW917qo48MsI
2q3tQZEcB2uNk1nC1JV9U+NzrPVN5tjKuTY5/MScIK8jqQWurr55cuYrAj5aUBwK
cvdM89RvK6vBjWbKyDtFPbptTIa6zfthuX6HC5idyPbEejqPd6FjVyFhqkD2YDhN
+rMJfvMMgUCLsjaWtW3ve19zACCeov3b0ygotGa0fpvBXhTR40cbX/0yXj596uw/
Q+3lpprcnKdsPu9bvWYAnbkyYkUX1IPGY0SWK17RvXWvnJkWu76ozJkNOlZo2E/n
zGzxPP/EHffO3e8qG4h8oFY9NY+XCc2LylbTLbwpqxUeuICqdmSLqdB+/8LcWBS9
9dQz58G5dIogvwCa0yavjQcPBZzGoBiBvDSzRxgmGS5wNDtXTiULrb2AGVJVRquM
PYEqiQPrYzUKjMh8umyq4vKqz4I6vl4yXV705lNaxx81gNjhjkXXlue18K7IxcBs
a9amdsnGdwf9mmwYIchHNbG0SMFZxg82UhEyGAKZ9iZwZVDp+RLsOtzOmOnGza21
uS+ynsBF3kJYM6bMR0D3LGnkbAzWBnE/QXLAJpg7mIVV1YNzdaUA+Br/1EL34Jdk
KtdUgQRTo+5CSNKWuaIeQwjUMieXNytzcvDoezGiKkNKdqMB9TjIawtM5EX+PykD
icaoQ9ehqs58lEDrii+09EncN0xCCD8yUxsY/C5bLXUAtuAy/b3QtJO+eXCaJmvO
jp7HqT2OpZWi9hEnGcX8JGrs83t1pGVDxH9HKzAhPg9L0L5govarGmnVUASyT+aM
fTaZeW2UVfcWT2ZvjnMRdZ8Bg3zyJcLs0dHeDNDACvagcHTZYZcqiUP+Pd6CFWjS
uNbunxBHWDXH5b2ir7M3vSoRNVl4/tQjytx0JcPcQBg+JdH6/S1rInIgmjk+tW7y
YJhFJIICvXlW38apjnim1uVe/pbfV2Ky31gflkGABwpYPqNpN3vywOTlU+qJsoIZ
WUiCuqY5m9M3KJQ/WGSO//rRt4+mBpK6WTeU2Hq+kzEW9vu+YH7YHAdcDG//IkU1
6mVYA+NKgS/k1N7AAdStqeEMalgaqd4OzRjhB7iO4hDgXE1obuVH037H2jXfPg3h
JKvghuoLgrSpDZOQJqcqiD7o2JPbPo64/ad4hXTw2/LvrExtnTyqiNmShkAZWGLM
kPUudGL8DFaD/tWjjw2Wi5tOgt/ypFq0hrVaklJby3quFTpwxmhhQ7hVuI22nTfZ
WRyU4flmCCO0/4u+vjWcylH02EzCuhmmge1d5LKyM/AVaxzadnA5hLQHfoHsnL2i
ScywG+cbYDEnlCl7++I/gWF/wO9V6O8lWTcxcV/M5DjJU82xZbeVrpEBBVQjh2Wv
ie2KAmnshmjnAWqFOVJ9e2v02d6+Q7rQCxz//Ur+yFtwBnd3p8Vp30GbkQU/8xoq
U744pRyFF5VIf5zy1iNjNzP1EdtqxjeNiMdWNv43zuNQMBYk9v1d+4An7bebBBnJ
stn9MirqdDfR24umBxaoKnFDb9uGxCIhKeLzSqJoaGJRRzj51Tk61m44+t89ilti
Iy6xJJ1Oygyp1zGnJcY+/CSSTpTkiB3RCsu1ODk5etdp8MaYKJ7RwuojE9UyweN8
aCIfwmxwXCbmDrPRMDZA/hwXgmPuJnUDp/W2I6czqeBaAcOhjr5I4A9f+bcyq+Jz
ctWOcJ7e7r+iKDdnpoT6boai6Gh4xNZ8lMTD374kQ5IpOqwgXB1qN9o/0Qr9ymAx
9lAc0l4V7MrtVIRkQJu0i9x+lBP2N75/om8Ov1QMX/qEHtFSuf3hg/mM7v+E8z1C
0k2RoAx1e/vhAw8yil7g5jEbTLeRzdjl3faJxPrMKWxVkEYSLZEYxAmSxRTgpVq4
dPc/3rXFJLhAIKIoCE7TtCAww/qMPu8oXyoxQju7mHA7dgSJ8u7e7XiFhaZX5w/y
xETh1hEspAtF225cQ0mR29Q+anfnZB51RRlCVEvVzN4tRqXAYOa7tBS6QjJ/BsZ2
z9zW6/UKZezdBIJekvlu0aaHPzmSvh9BtE3TeqeGkoOn0lU0IbU3HWSBlLwjuwzi
knd7rzUI/VZ7iJC8ONF7jeFDkJaXtan049VU2bwUVe8gx67xFWs/7sdC5jj94uVI
DAWcE1gRJUtmike0Lzr5BQjfcL8OHki2NwGr9Lz4WFuJGcIqeg+5OWVFrZygwqH0
oLNqrRpMk2qAtUxLAXSdnnl9yA4l7d5hAz74w0QhN6kubTRMPWRaEDPQe0/7tP+D
MV79WYwH94hTuVmAa+kCh26I4Jgy9q+2qlngsb3EmsOeYkGGwguSeyJgFmMELB1x
+Lous/V0Web056LWYtsZLXybqt1NqqZBhXfbXjrjy0E8B6auxmeeYECL7YnDknz8
nddy53VXbXybQynZ5L5G23ItP690F3UZuAN96XXmF8QWpKDkbefRHJChGJhr0Vid
yK2NLCRoeSVzBinE3ciiE3hoMUQ3jn3BrTChAssXVC9k1WJzwt/OBquGcBFbdX7m
Q2jXIIu4znDYS6zjHQ4DQ6aGk/wJGO26guFL5Z/nI3knMw3G91bAb56LbGgN6Yaj
9tbdhZDeAwgmYoTLRnQPy2DAkBboRQHR05pSgS3ANqdC0Sc7gX0lnvKxpjGcf3AN
978T32L/UMt47FJVvQMaUqST9q7Hc2Kj7hRI+0/S1Fg6Am3OCeaG1DVIFKvs+vsh
F+fmpLCpl1R/Js65IlzPcI3LQuaaE520QXSRJfFFd7dj1zmqJmkJqsFxIZA+VbUE
6enYVXikFvy6kXEp68F+Hu+W1lLRYxjRPu659zyPSMTG3SYOz9+hYePWTYy29L9X
GuoMl1W9CG7/0VUzyqnW228qoK92hJ5Od2UQvaGhiYd4hYq0w0POVXfvxOluNZMH
A+m986Jt7r7q8CGSjy9ynO9xDb1/IseY06wspo7k2jqOKrGCHPbmsNxZ0E8vnRBB
QFpesFRvAzr9mGVLR/vkwChcRDx7MgVKvuyQqdL/Fi0nxQbppLHH2slI6Ma9TooB
yQOYHGqkLv2EihTrKCvCMpylEr6+OJ3F1DcFdKmgdFyytSKX4G9gJboTFE1lUfht
KI3KxGhThDRXTvMlKf+McePbGV8hCMJwj2PYL+Ui8Fz6MmPLhCSbW/BHnGBh/vUp
UchYZuxTmMicsEfzV+2LQ++IXgx3oFDXJH65P6IN5sxscUvyprXVrgyqlaF8JNs5
4WVS2ji1WIWB5apGZfACgqYCGpUXnGfhyvxPC3vQ1W9SFeAYZciJbyUeXZr7/2hJ
aJiZApmogb7b7dH5hp9LEHi9ib43ItjNMdDfik+IcTpzOgFONNtEOmZWvyS1zCWF
s0BGnoCm3LTXyl8z9JyN4o7sFrRDjCZqwoIpDhjm0aN70sy2eEWaIutsdil4PEoj
uGDi311qBlJ9CB/TWKpIbXNjW7MT0/LT9AKVkejffz/aPuDMdV8lw7od2QkTWSsU
NNc/K2gSi8u84CxXMu9PM/DFH9RzCWG6qk0cMoJNc7vPOsTYBDHa33LI13aFq52g
S8JorRQ7r7gjriaFGW6gs9G4iBEusrIo4N0KTr2UbWsMbB8Q1TszJGLQA7Md/EMh
zQSKTK7OyAdn259b0cBALATBM+CurBXVwCiSlPVYy/VDmDHbAiVcSZ556Q+cAtXx
Bz2QC+yeIV4C/71jflqC5yEECoye+4RthyT5OKOIJntFO9snqp7bcf4LwpFYUExI
RGCwT7yCyU9Wp4fn0Tzo1IJTuBTqEj2XSHju3R774aGhy/QTdA68XFU5rwfAgK67
dXWscfg9Bq9vQaTWtNy7yj9kPEXQTtgEe4K1Hmvbc66aVEFGjeqEUuv+OLzzpf/O
sGwBb5mvIcW5/FTJwherwhC1Vq5C59dbJM4qMgj+nFZzn4RESpDrunCsaJI09yh1
iO9Laqzg8xEhyap/n9/boMbnC6fT+TKlySPr6BCYnx2ii85GxsIJjMQdI6/5zNYp
uYrZPkRubFSkk2HmJN7b4O6sR/M/OJgdCrTWz78PS8qNr+vBpVie9Wft49TkgNzz
+GQUy5gRBsTOHa7XBnsuCBoBJUYenPsPMFQ56eTrWzqoMqgXW448ns3PjAZyTXh5
tRLtPX7elOHm2RzfbLttLY8AJGPic24Lzc+68EAriC/D5u1zEU797Qc5ubXopCBk
CaKXtG5ZngmOARMcBJ87Hw08IaayLw1dSSTEcnzjyQ/8rNdKL9F3w+32848Ky0sK
MOz6bm0H8uk74nrCC5SxswXly3mERTVJqm1xeZVvrWeax6ZkOhoOWCEf96UBt7bB
T5r0YAklG18ow9E9MOWOMvcu9gqstZBbUtVqozc86KlB4PQt6mdQsPTZN5prJSju
y7zfFua8QnOKhSC3dixVPBzC4SJkt8ffyAL35pnO+PYxRNOQbI4c/0xt+bgBICvz
3FT66IGMXLjrvZBJocttRpcc4Qs5YJRaR3XymZ8JCwiOf7a4G479m88F1YILCRmr
egd9Jm0+NWuUooY7QfRwlrceep0CeaQ4IfiK2RDyRpfKXzejU8e5rQjVuU9GsVNx
m3ko4RB/uhEUq0XwCWZY3p8MM0dZ8TLkVACv1zO+tC0b64L85es/Bek5PoLWSpMk
rXsrSO3iKrPYemrU7bJ+Uogo4cUqZHBCGkKlBOuhZM6GNmIi45By9ZUQSZHS+Esh
jhWHmCspfaDO4umUQ9ne9430DN85H7+lO5pLflopVjn2Ro61rh6U5kn4+agFphD3
GfaA9w+iqgwe5IhmvO+HVkCiOK8Hcv+jD97taeRFr+ShoG0wcSVETd2bkK904DmN
9aXQCDiD2usveGHvcituQKsml8MZmKY/5Pjbg0gpFKT4ZXJc/7AnstpvwWQLdVwJ
Md/mKuv3PpkLMImN2pTibH1dV7hfFSq4080xn95kzyYs/nQmWVjZ+HJMZ1qSwsZ9
/xHT5OGvvVYzx56kp+f9ZUbvC8HUInmvdQEoRlGtwhzLCcW/vzkFtSjuIk3g66H1
jgA9mQxipIJ/XfZ0bQLzTCPvAekireyAiiQHnCMJg2c3PEPPy4TRgxWvGFuHYjVe
4wuk+UJz19oiSwf7AM6uOhea7M7B5BjH5dgQ1A8Co5taLzCi5mw04duazdSE8Pk3
vz5x4lh5wnKBYpFLUHSkSgVTR5R0hvEr9teclRQslU4FtCPJnMVO3dTtYb47InxW
90QzbmvnWQQ4JrrbhgcfZih+Hlnax+lu2xtekfel+pmwk3lzR0l8V4Bnnk9xDjoY
Y7kDKFWrS/Cxh2IFXAYLgfRF7/fRHTqVysYIsGM7KqIY7r3obDIhattwP/asMRF2
t7dl4F0AdqfGVDj750na2dfuXJaI0LEZK0dY7YrWE3l7+BVizqmOLEd2brKdFjxl
OQ7Es0Zq2ObU175Jd8QSqM+TwpnLzMRZHu0BWfhq0362RCnxF9UFAJXB+rL4VVzU
2x4GyAoqxRT8dPZOa9kMz4uXZcLyeKaDjLPqn7Px5vozXlOXVYl/JES0D8jCRPDA
WGsyResSU06z10UtnZwpDsc8KhxtNVRGsMroE9yPuDCbMR3XaaGF6qygreEELEkd
B1r4tv2wdiQiF00an7C3Y76TCBPpsj2kcwjh+mje6Ce5TP0aexUpcQhLDX5Cs/9G
7yrn3cOmbDxDvPNmVxnzmmUX99XUD4aOy8yXXLtv6jT5OjB1tkPRfiud8ApDuGq/
t7TNAICHr9yXfxAB21+oh+gVkvI9Mj1rWx/Wn/WJoE1PzS7XfjXulmQ9q4iOy1Ho
DxYIlg4ZTMACUnVF8SkvqMfaaIxs72qlNpd0aR1BHmJYjwaio0xQuTbbro9OVGB5
Jm6fugj3JaVPPmqEuEk2J5BnXdzhAyrcMUxOlsSEucooM62c0a9g70toJWDC8Bma
pQsfrTY0rC5Z8NIRabiYLQgU3FDXmoNob9HPRDSLRUJntw4dRQ29UN/cOCtA/Xwp
Awr6s2ZCp4CdQCTcErcY7v9fZCEGNrXIMhc/f2B6XT/ytDQjZ1us6YRxHRcOlIgn
D6Fxdfn0xQfdRbroYiG9ZWM5mFyzi+KT7R1P4pr59Oe/EYBqZoT5FL/5K/L0/BKf
Wyn0xbSsYT26mEeZZnafjtC0NS4X+lCirNfj55bmF/Klx1Ui5N2QGjqjH9zemwcH
tyrbFI+e4+tkJQ42g/2GdPImFGRCs6f9ZkB3jMUUCkoV5jTuDAX8BNJByP3VFnvA
e4DIWqOpU7RLBl0hA6NPAc0RidzwnnPGdL9Ojm5bpr8KMW1aNL/hdfNJnhWdgxQL
CwseuyuRTsqkqdoHD+6j5MvlvCJ3+k3xc6pU/J1sJNhqdTUcshJC8UzjVmQN79E8
tAyCZFFU90+T3QQ25ojlkZo+5RJBHZN2ZK68FkNIh8YVayzhDOVlJOjM1slOfdOA
QIBVzb5dc7TXAg67mCGB7ZvhuVE1EwzST8+NS0GMqiWmSPDGlxqYLa9gBfGL14dt
1vm6BQsGQ4Rah0h/B51ss6OwqSFeB7qwGuksi0RVZhgcIhne2xCFBltqsDq3Trgr
WUcy6zjwYccbJYfQ1385202DOsVqBz4MLZM65kLPjHx2lRKx76M82gPhaHqs7teU
70W5kQE7pt92/TO/rxXYuM4BLov29/o/2E7X3f8eYcSUN/c+LYwNj1yGj8CEkTBk
n5R7HPdcbocUf1gJf+FAzrwOkmAjDkzrTt+3xCdtp3pQRVUhBfpxtD3SohKlBACk
D0yc0Hs5I1yl1WQ40eimXTTSmR/Y9XKhanI8RN8vYyH7V4pTIeT0V2yazYDTzuEi
qxWuW7m2CqizHH0QksQc0mVvZy/WtR5isPdAiIjhkDGSP7e2NM1jA1sCYcSKWS4A
PqDiFbzjV/Vdm9NcdX9nrCBpXfhlLqyUzpYalSua4qfj0BU84SrotvNb8A3nZPNb
jzcbaloWkMMzWubNZl/2CY3KC2m0hPijyzk4zRFwY1RxTJCU4PxOPzlpYTsnKhhQ
3o/ktMr2+2lG1TJUFuJEEGIJD3JexNCqLPkLgRO0AY8eUl/ryDWayArQ1JDHAkyP
qQ/SAseDROp1SgHNhCMgwxcsNTxW2hoJMpD1iiak+th/Yx0mcXBij6luZWzf/Q+/
N5t2h2kl1YMi8O0GqKEaV6eR99JdxBdbGNkqQkhdJX6cz7Umzs5PQxyREX1u7Y+V
Pq7kPc9G2aHYaR0a/NhoPzzewXoxizbc7fOLiEBfAw0cASqDtCD4vksWnPvRtytk
Sx7m1aCkfcsddS7rg+5tg7HSXY+qXgiGydEJ1qEO73lveOQl3tuCEFvobAFEZJOw
yDdh/wKuq0mRohgWhpeOwOLYtxtJPD0H+6pEl7dIu3LQzm185YcZWaidQs16nxAo
qlrvSIcWMN/9d0dz26ioYu0nfkb3tP1y+Yp5ALuC3RCG5793VBip27+hRPUIppg0
q3yJ4fgoYFr2+9BqHyC72mQDOb+CooPehTtqtIT4TFwsECYi2JWcPI4qqnAkEHOr
/GdjdLjIZtBjBKWM+LBRDohWJKxjzNbwiwyHyxsXSRcXYuNTz2LzAW0/Vk2mIxL1
Msbbg3Z8a0zgcQriyR5c2U8o5uRkxpsMDM6uiijvZ95wKSOX6EIjR86pUbFhiPn/
cqOMSpu7urq+zivp8RC6fpdFQPhYA1q6OffeFlQ5Aa4BGTJkqI7OzdgqNYYt69Mt
l/Xe9LsuNZ5vR8rce61IjDBw5fxcKBWjiiiLzEvjMFzrFLXFu0h584xqK1r/dKGl
e/CTr17wXsCEeuKgKz9oMk2tc2Lht+Gv843VrKAWuuIQXL77NoyCb9twUOjpyX24
79E3CAY6n0SmabJqFzoQwm69MPE+IVZvCfRJGpaaQxYZKvmUrLbYmLc7+1dKAFQ4
vxQoQzQlGaG29IWtScvtLjXFg8CdWXVaqPrwOCwqK636QfE3rVn61NgbLtGvaU2A
76pe4w11A4Ic68Whw7CZaQGbldLeSQQ9mjBS5f4Qbga0Rff/SCTrD2KpUID3bmiz
W+VPua6ZSS+58bepAQto6KxrpTD3/UMBIF/3uGmZ9zF8VBKvenGqYUehnEqeqXQm
pFyVH7UcC+Ju4OdVTjBQ5wGHYKLC+KDJGS/m6CqWeleB5wJZJN4AXubuco6WP0Hm
CfGu6TGC86tF3MkbSopSwbVihmWArYDGAzOqSNyU5XYZodUSvC98quWpfEhJAtmm
93wauUXzCpwOawKrC0w6Y6oFEBnwn+kjfbpSTTY/xJI0hgBaTBg1RJCKpCDrifZ8
uiXmdh3QFrJBkVkFDVPa+IENfEXEsGbPDAaq+hN6KqwSIeAOY/KS9jHRvkwaJCB2
u+YYXGeDwo8NUzjLYjP+/MWV0Tk7ML2Af2YanAjHFQTFS3QvaFb1xrx7Ic9Zj8B2
n940GJP8Wj7sA3IwKAbwJhg3Z5Jppl0dxT5DcmVs/KpyHtvTlan49xAnQBR/Jqtr
4AC3XsbQrVeWNZI5xL0PLLwMSbkFDOm4WPyZigWKvVoGOWMvavsumJLY24T1M4Ei
+5gcLf+49iLKqVTBRHxYwKpsBT63pUhfgPnzzlrDatrIUBiPUvlYmos1H5tw98Wa
u18xfhdLOlZiemDyaWVckX81NznG1c2zptOHSo954vs48sak+K/7/vSV7hiTQ8yv
i7j6A7UWn/teKvWRwU6kqeWsZxYyDMRRhxi2F2R9bNvk+g20BgM/uvJ3oWrirV+Z
9dBZJrj7c3qXW0fVrM0t3dIDzQvEExKQDgRqTC9C6dm6Szxgd9QmaIvnZ0ZcLrTI
XzWYJCzOuXATJZE9fXg9DWjWDm5KyPCCXfUrJSoA8kHRC07U724WUO8nJffl9e+G
6Y0llED0CoAAB+zqc5EJsT8WRkuDrA1U/NxMcfzCY/J7F27kmQHK7LVCYkTgCAHp
ahQU1hUhOshN6BeX6+Cm7r3U3NfdpMytDbXAqLWuwXx28tjDlfaIH2xbD4hbUrHU
CBq+MA1lwHOPw2MMZIjTSVEQEfMKWFau2hYcRL9X04J3h7zRUWnyi5a9vFTZzQpj
8igny0+C8el5q1ujMRRKn7eNaS1vUANxXCltA2CgBXAIqOp+HJBb4e0XE9FJer+k
L4MuMNsK07iFtW91uU+9fGQzeBJoFFHhfH29aLTHkxKDaE+1Sz7wTBt74NNbEOGg
VsiSIjI+0ulExtxb6Cp7emkppSWNF3FpwLZ3yY52yN+x0SVjcY7N+xAh6j3RypVv
przZz2rV8wTxdmPIN7NgIFKXr1X9s+GAWMtXn6rfVkxahgQKfcsVU9G1jASxrSN+
xC6hNa2JwEnzF/rXBF63P6He7Tt0uRZvDOa7TxyvjB6/kJxgSEVWW+rvlKx5T4lN
r7JGT2BS21UWJeTuiHd8NKwHmOutUljiIPb462MSd2/LbmP29wViCHdhCDkidGgt
Ouee+kJu1ma4md2nHpvxBDYXJcIH/pCNOl3Xt3A8czGYhHfJIoNUqMFmV4fIsWrn
wbghiVzoIzOClpZK2DkoqTB5/ITJgCTc2FhE/sJE9Jlbu8/j0ZnOzREoyVpdapan
1ZlNjk2dhJ7VYAO/LpaXUrwIaX+RxOPhiKzKlI0YDrbc2xbuTrnywStyAQnTM0gG
r9WuIyyfVbTyCn5rkWeig9cl1KR7IpGozrybj+JAdxN77siULScOepvJl/O9CNGO
udXgMKhOYN9kADnohi9o+p+x1Ojotq+PaqFTRiGdtq52I+81U87hQyXv4aQJBhzV
6qgsnqiBXaOevkfdyhED4JE8FQDa0lauCe0r/A+oKbRG9MHapIsZyNqt/cycJ0tu
9vV5wS6ikwOJmuiW3L2WF54xPywkRSrGoalvRjZ7p6tuRCFq1pUlaof/8/WtIjVR
wBM8y8tkOsm/vqcRNhhBn4QOKjEXHxEjOP6OA2JBFaPCowhqA9QbVSd69ykPW5WQ
4IXwxWeLtjhvYcA0E7YmXzTh8H24FVWCQLU5Vf7sX2GbbtMQ+YKuip3BPmbWQUQ/
wy0nd6GIFAektKgLW9D7n40jq+pwsy53WXI1rgvCGZaODNPVA1xYHGwSaQYDiijO
GjQBEg3ELY9j9HwSuTWcFBzfmzyMyS3TQ8Z5+3r021/tflv+u5tXdoGJdMd93iTV
x1QTXzYqJvbonSHqrJkMHBH6AtNLlAY8FabSwYk9yXWQPIssZSMd65vqT6lrz7HQ
wbdivahy+yecvkRKgN941xnUJ7kUDGdBdDzjggmm44gmd8kT5AYh3KGaAj6hCDwq
d6J0YRee8gZjB0d+gec4qxY+NZiIvlr8lgmSPG/FlaV839LdfTBC4/i7EQ3MFmQ6
4c9zzZnW53MLfLooNU3ff+iZiCHjyJlNr6EVChJKOPmELzaorp+5BS2vEt4bDgHj
Y1Zmae9JePN4b3iktsEoLq1bt8w+1Y7rJnIsYnjGy33P2CmhiFsSrOjoRIyBcHKW
k+OEcyaOgTy1dR6QmkNzjIDsuve1IVvgBHCcpobKNZZs0HfXG4WgAUK8rWQd9mP2
FBhnr67G99bG//FC6kpMZam8uTc9ixWlSccqAJwpbddA6eZRxI+QXngOuLPdnb+p
dxeWGpRliA6aVrneSC2gLh73FnMWxPJRWQTxvQx4DGkVKe3auOo11nrMuj1una/v
LhtXBrIYBYalEHPZZl0nefaLK4sQfkVRWinNE42wtji5Hqm/kEuzdnbMsv82pR7v
+j1KQ43yGHvLOVOgHYW7l6quNlWufgt+CO6AFyjiiaMv3SMqGfclR5Cgfki8Mctr
MLFQZzyoknZ6PTyWfN/On6ETrbLQLtLNbc2QeBpp1dBZihjy3TXtcC1BkVDl9mbh
4YZ0j6Cg+eQukwOb+IX+vp+MpsLQwO9UurGtScItACzhzSfexRVVczbF2Orzqppk
hVHiF4twifQX7hBDtiDIZJpkf/TOtOAZm6UCnb3DFahRo8jKze14u0etuyS0K7Wh
VwQo45e4qD573Z8/xT7co1AaIsntnSDk1RmHDLxzgSjW3zvAK92pfiaQ6dJ6Rhiv
Ys/6fcX3INTRE8hSZTDW0+aDJ0vTDamrKWSuik92fdp6s0I/1voKzNdsJ7/5J3zg
I3vzTKRQT4Aj/8NEu84yendSeyD7kq9cu9CrERIenv6d1l69UDy3ZINWQBDPfVfj
j1neddq3Uyz9HT7gxlJNJIC5i4P1HBTELZF3T+GyOoP4kQhBatkyHpCW5xwxuWbQ
YOx+UYx5uE/zYu7TSo7m8zuC+ohv+ylUMZduLI23Et5mpqdRLQh+Z05OLzbTw7fQ
9FPECxg9mf2H2OMolJbpeCIBXJv+5w0SM9X+09s9DIHtnxoL/rOCEBUWnjPgU1Co
XkC8wSzLE9JwvzI28KZe2YR4r3yn57dOsYQeWddtp2RuZRhLnz4w5rCKNN2Oegow
Njao11cgkHp2CngumPqQ/Lapu4BfzDj47tpscB8SbVNgitaJqy0CpJHb5NfeJLQ/
tN44NBMwWCnBUdmpbKYulA+dsUBBst8zuISvaml7+uEUiEjLTjO0jrfBZ5CgOYYl
9lW0jGWagcQWfIKs0agO/W9MwtXTWADh9zkKBQikAr9L5zeiTna/mYZ4jBn+vO24
9N+eTFpXO8QwrOrTMt2x9aBMWRrcT94b8KBcgMZVNpptSDcZWCG/5XuDuwhJ0TJV
GT8Y/TVfrhZQDQLhTHr9W51V5sMSJBXKXJov+x9wIGGKE3vFH94mncsDpiYvxB9+
nQBHdnzH0sFwFK6p5q4kIvyGnzC4sYX2pFPloaPuTBHzibaoTFvoq5ti38cQhdhm
uBzb38i/RZVqUhzeCGfIIoMeYcdHKMSG67ae07Fiv1LG6DPqtT2bZgmf59ddVpEe
kdh5g235cMjcFy+tPwXKZe/JKfJveeC1a783xDstNAXXXcb+bDPtOwRPcAxJtRTN
1bYHBYaHo1YheC0gN0LFJCgy7k5psOeRNomN3MP5hhxhdXH135wuRNUIH9mxvj7C
tCYCRSNnqwToxu0ESIl0t/idoeICFgIbER1/dH+Zsfn2idnbA1ewy9513QCeWotO
rn0tnvFIlMzdew8EAYwa5P7OEE5RhknVp3qj1LL6d1PmoWKx3pIeB/h5F8A8u2Gn
7NIjuvZEFMptW7ufVJ47SPcBjNfzmmyiNDNDqgnTpNgx8ukn68Odng3ZT1pD7lMu
uu4sxRQOUPB+4ftp5XWHWzZh788k/Gqv0WOzlD/1JSw8+CurhBuP0IEvajS/4kWt
516P0K0xTDttWPrfxYzjVjL7jjkc8XUc872keZJOBt6u013/wvb7eVYShimPdypY
dxLQj7Q13lqSQK0BEqPAsoKjpB37hm0IwjiwDDbVZghjxCgy3EhJYX5mD5JcuL+m
Al/sNmUqMxkB+eYDY7OqeyOIa0v6tS4vTsgyryOxNDjPArqLN6E7XzftrixACsc4
0WdVqik97Y5UqzKmK+k7gAZiMyxht3IOF6GnaiIJQ9if0MlQuPpOXp32IUw+da5M
Mgd2tnOk175X+95mO2FwSNFk1cIIB/2XvtnkcV1+LzuNXMIlj0GbPP03z7M5EI0R
f7FETopd93jmlMJefTRo269+7Rj3Dx4MCMXoVjpAT7FjDN0wtLpgQbKIsN21k4AG
u3tkslYZlb4lhZmlXa90fYmqmLdDQUISOXTmVZMNk8Mji4dLNKUdxVQVJO8Bqhxx
2zpLt7+pYFWG8JJSjkmctOdEcw3FhLsx425Sgb1pUZIfTzOFpoVvSf8rpbXFOTj1
L3xvhNJUOkYz03oWwTuvVDiJdx8xgOmuQKpTxhlxJzCS6ab/3Y7nSbyMW6og9JY0
GPMJb0RT3zDwwpuqq88uGO0ryb9HKiGvqbkEsBfhOUq7xb5+Fd+stxwwCSqqfcTi
0C/TMAdQWTiSqa1Xei3+vAk4afPh1pYQYcKBN/8RTffLgxdDZL4Y6nlWpb0KXuJY
kiWM+sqNS0EMbKjNPI4z5vwjKJiR3gXf3O4smEHFP0WnCIWjMddSfMfcQ2Y4kN0x
7kyl7xw0BCOPf1169B8CX3RHE5+Ku6EZMOrj1P/Psuf6tokTIvdVJxMNhqqzvXaq
H6IomDdihZbKcdmdIi6/nSIlqg1Dx+AM016WJTDkSUGO+Oq8OPm77TaAZ0rKPepg
hWyW4adxDIXCQjpOYSoAKhQ49J97wyeQUGzp5I6nUFZRMaO8cGy1XULQv0yvbGmC
Lw9Y4fWqTbWONDxvg8citGZEuu98pFKllTlZdFPRGCsRAFePYFEIxZJ7C3V1J8ty
hiPqCfaj+lZvAomEI7Ea5ZtGkCt21byWA44ayBPWT+RECNOnT1ZgUeB/hw2JmySm
1epxMEXPldKiSsTo4p50VaiIV6Mhk5q+EFJFQ8TQYKQBicaFnHzFBwoYRioAq5uW
tyafv24CrAkC0/8RVkAkFA+xzKtGjJ4+Y6YU4jNVUsCd6jhqCNprJxKStzVbUoT2
jp3VG0+hTIdMLJToKkfes63oWWl3tnHrQ/ZTQy7XdKf6GBEA32A6np6pxFN1L97b
Ab7W7OmVks2aa8G8d1t6XNiEAHMD7yIvAKy34Tpke3DkMhMv0wvboSFA3op7JyvV
P7IKu7sYALRemZ+4ciQKjgLJWuvQqPSTPaHDFbCifuIue5kvRoJkWZBkDg00WY0Z
ITGfHY+YtM2oLjzzUCnZOLy39HvaQwMQaCTF3jKkiiPt1sfm+5zQdH2oWaj2ngbG
BsV7ROnRzm7FqhUiCbvph0+gYoUdVsjb5Bt66aP5MFfvisGne3tliNKO9DqmTvm3
eqDLYE61mlJ22L/+1zuOfQa43GHHj/ww1wWLnHP6hiIrM0z4gxsp91zaFFzQe1tE
sO9niaGZo+dj3nZqOKLelKxIWbUK7fhxUlfGu5xnaibTBc6IebZtiHm95MpgfaGW
8YqYAGe4k6CrppIjazRJZYqLrNAomlTd6awPb+HHmmGpYOxjrun+c6ii369jT9CX
NkpaIhDN2vT4KgGUmLpWyyjoS5tp+WIej8oaOiwOsQx9q/GxsHp8isO0zqjxG6rq
CvSe6WYYiG7/CLMmiFEL1PC88mrKqTDnyjHbsWQtP+smxOT++SQVx2IeIY75/8VJ
e6TEutYCpqSEzf2sgP856vPb4gozTCcYwefFf9pynd9up9CGIkr1WYbze88JguH2
4qUnEVJM+Gk64I09/Tk5nN0tMKXhilAE+5KcvaXqTITdtxeTXle71XtaqRZgcmgK
D4h916OjolPGrfHuDOrCCJfru3Ei2gTIst7P6IXXXS622fAzXyL/BBBWEOkcbzQ/
WjydQFna5ef9J9fCNHxgIZGdTZCnHUNNK1MVkIhRFVGBORWPiwIWNG5TqxFIAfnO
L8To3ABvzns3wSl7AVbNBcOXcgKhT2JTZKclV/yS8BfSHejv/7d4vd0Vn1qyz7t0
O2i/QkXkIrAYHyxCNc874HveGke9yJq+xZobrSNI+mJo4CXEjNF3ZezNX0qHOzRf
79KQe4I7Yi6E3ut+5CgZAGBWBQi9qd3y3wAFqV6X79BCLgLheYUipOlmNhmswhzM
06ozVz75XTXmxR+HzHmxo0K2Y9IFkckm6J1HdA0VMUfHi2Bi4inPqpwmOS9kH+U7
JkN2W0Dd+9yRfi+YZUFMN6GNkgSZbc+nFxODK1IlNRIPfS3+mRAOTn/eDWiHN/bo
0Y0398Vg47ttxAIJS0q76DTxEb5X7YRcK+8O7PYMNXZPVK0kN35fGDEf+EOzl1SH
QuKA1kiYOysu5W3n45iMquAzN9yyn0K4B+c06Ij//Cpym6XEPRYrE2CBXQ62FtCx
CZJwpkCZiZPMjDZGxOYmOAVXmxzRoYVgfOhdoOhvm1x8AwwfIrvHA/U/X5iGfaLH
6fq0Y3Lmz7KKPv5ym637/1Tf2PtXCYSEb3O+pwaRIddKdh/9kD33yufBR2lJOPRc
lSLcsId4qfKfn+z0C8tEss82qpREfmDH8h9tQtSR+S75yDNvjD1b5+2i9I159g2Z
xj6LSGGxIydDgjMT0zX4VgKue7zsxfuQvSAN2ASegCWAnES1LanuVEUMS+MaC+Gp
j48p1fSN+/01kjUy/++/qOvxXdwcjpp/BJ1rc3zKUKB00pJbPAArLEuJ74QZrywM
tf9OltF4mDi7F2JWhCFkScq+wBEmtO0u9OenkkOXOPCbo2zvo7Sd50uFqDIuYV0p
pS4PelKPUNEVMqWQ0mY9Xnc2GeVzRV8FFcUS9BoTKVPJy+iM2F3DKpbnFOlh1mZK
0eLjARhH4HA6DZpxj9pgUlGMi4g1lMT6ICxMq1n1rjK6MD3Huf18D1EgpsImHEHp
8CUum9hd3lW0syPX6W6PgUic4OvDGeF+LjWUqi+0WCuWqv8V83Qaq3C9TDwd/Yo1
AbGBX3jwUloC1jANN9czF9tG/Bepf/q//vtYvCv2/J4rwBFMC9AYLcTCSr3hekI1
hPR6pjQF+83D87f1hOouNygolHsySMHakUZ4K4t62dqKN4sFL4D5uoLYCieOgWeu
txUYfQQ3UuYCywHnon3447MtisqJSyWGu6k/P+gnvB3e3Ok253KhSoX5i06ABmFA
lqOKjGmtKf0ZbeZs8odemrZxeIvgzQJWUyzlugA7eIXsr/6vj4q0InhvauftPpVd
wiawLsBY4uGGVemv9n3H73neUAsz3A8N8iZux9kEj3NCz1N9iaVvXskSukNYODgL
DBUwRGZR7HYYAYs/e2KqEQUKYjxZB+F1q6i2AJb/S+ve7IwXT/yfw/PxFx4h3PYP
lQCUX5WkfB8+SVKtUQ6pnLx93eKMdbWv8UEP+F2JVTOBauIMDrQZvvqqexsXdRiy
I/DOKwVqRdSWkjSJwseWD7iC2lEAMJ5dUjQxcffkyYN4+TDJiww8WA2rCKw7f+Xu
SYwCw4JsuncnXKEUs99coxo8lOtQOmAd9vHs6B9YWKp44GD4SBDMMD4M01HM6wSP
4hx/Vp/QLWZkjsIUpktuzGAYRP/aoEg4A19XuFDRXpLuhIDKxDJdX6Np1mq0DX73
S9fZEEe0mUSXopz4iCZZdihGnDiK7ajzF+NgrAiXYDflxWWfCfAMjwkjn6+fcVFs
YG4ky4Hv+GPLDP8BPl5zrD4PeS/mszbZeen6f2o267iTdPkE7uqnx834q6BgWcOk
hqmfO9e5YfnhG3ipg1p4mf0PTRR38ZiUYAZLTIcAiritFwjay5mnUWC6Cp+Rhlsr
0gVdTAgEG4fvl1wRJpnSNMFB6kUCGUp4wXyJfRvB6Wzx4GhAJl4+6gseURPGVsfd
kWjnjknFlvj7lHM974Rg9Y+hbXqyGxB5EgqdTwA1hnHVHjJWhsOHK2nOxXSq/GMr
ilwgUnnhOzaX0x1kukwnv9HzAGHvRTnPo6Z1zYqv+InlnjfuV0S6dP6y/X4TRv9p
oqdR+fl66qNMr6EZS+4IGCTh3+JblkhqSulXcP9LXm+Ks95OGqGqJ5K0Pr9Gzd7D
7aqIEjuJOs4nK1znMz/ua1pTzB0WwFBytsfs5hE+Mkm36qfi6FGKn7TblzKlzDc0
pLbObbhhaeyLzLdAjV7tDs5Npjz4iBthm8ZU1de/uirYj2jlR5R+UP/C/eorL6fO
qYlxRDyT2g7a0xcs9D8gbwr7ViRdTgTRTW/q0QGTFAMq9IbMpNdV2Mh0jaIJ64BT
R18V1B/mrk2BMuLOIBER3H/MhSTXAY+jkV34GeVEvzpXfepJgjiYFqvPPinCt/wv
P6iZubCQtbiT079GdLkc0FnjKpuFeARnae2fXuLAA5b9guZwLiA3DUZtjlcYuPnC
LeZyrF4PhbjgbXSQr2TMYiWSLlV/Yq5eyr1IdbpeF/e/6+OD7okVOWnd8ppWbGiH
a+txgAcsX+gAv1k4g97UsDrvpDot72cKOBqzMbT0XJx+Io2NlA7dv7xCD+OEjVhp
y+XogRhBxfdpwASxFLamTARadK5SHvY7+ZcLCPtc2Hjuob9rP7pDs3WulNM7z3vY
oKKLGZKKshE2CNnR6fUfzKMseSsgAJguZ74KuGIgCrmE6IdWwjkgrlwT9hOnrLJk
ILJA+pE0S3iYuhsy0EDggUjGS6nVS0FWqze7HOCmAzyp/qKBrjXXFP6FvMmnbFLC
Z3uuU3sNNbRBw9HHwpXzFZugfDyaQlMA4+7ww0u/5HwXp0WrR3pA9b4P8whxH07q
x9IpVHhyOCpTleD+sM3gn2XXzS/CZU6V7Cf5Yvl/Kg9FRtPZT1Z0rsNxe8dQhfIl
YRdFKkIttfxEUVg54psyuNI96odHSw9BQE3dN9yiOu649hNXVzsSBRN4rtabpAa8
MgB9CzN1PJBPmEhw7p63WhW6QV33lcwd0ChzdpXwlEyjRjBuolxHef2lvEuOhpFo
suafgDBuDSrWmS0Olv82Suw6i78YxCuiQ0eUaIzuXrPK7klrH4zC0fAGjM/ItLMs
EhQOW5VWOmrr3FBITdSh01PyHyIDd5FE+f3nuMJccPU1hQnUBZRfhQ7Ag4J77GUF
E2N5iCMmjM8cd47ouK2Y8qqkFc3B6BLFWVLLOBZeuVw5HvDWhnffNcGdiAHfbE7a
+wpFlM7geGWylfTLGJfwin4ACoz7Qt1i6V64ffWFTT8pGGt+AylIvUoAN6Dnojr2
41mZm9ge4LU13cwMvcxitkJk6t6wMQ81Y6cyldy/hn0/07HHsHatXPx6mAFh+DG/
3EWT4/FhcBAzdA5qm8IhDTiFiUtgvtAF/yV4MWiJui+d5WtDWaGvVJQMoWd9NmeA
IA+SKjdZgKPE+PivaenQXRhNAfQ0HQK/5DjPx0fSci2X/g/dYYVc/oqkJNQ7e5f1
5Dr8bdxeSqUSfs+cnE6vdJnKcc/e+NFx/pCGnqxkMUCxXOsdyL+0u1DoygzfKf0D
50uUXJib7UFSLijH1PN7dsZ3lqFg7lIcFsoy5rUHllmZMB6wBA2bbn7ExEtB3Gza
3crHX4Eg5PXI0f0u6ZP6eyVs752HG8j+Hqp3bqgSBB+wBvCwfJ7AkQGFJQjQ6xHG
XCD8h9bD0jX0yDzYT/YvPysP25PG0ljSY3h6jJioCEAgQ1jdw3dMRpON7xx+GHHF
2pjzsN6yt7aFBUmaXFpmNqBuqHg4LXqvBjmEd3B4w1rl403BxXDea92q03LjV/tD
/NxG8+zhQ87TYcwu4eIlKFbBriG/vshrOtSMxWkInlPt/yNug8E34B6VTfbF/8Jb
JMQH1afv+4+kQBv1Dq+WFZu8pQn2n+kCr3eWYArxLM6qhYMDeZV9ciWzMbO15Lym
05g+WN8B/ANpuuSg44RTeaKyJOZG8eh8bQAeVGW6ENGF2z1gBWk1XhN5P3K60MH9
rDJyQll3cffqR7iGon7w+LyYGArYpxkHpDZmWA0aJ4vEohdTmvjc11vDUVJJAKsM
BTpsz/YSClB11eNuUACfsfJ/zLSl8bimZjZ9vNn1voydlQb0YNurz8XQtLpvEFw0
vFCpj32BO5Y4G7PG/BMX6GUq35TtpD5iDVSY5kHBIZtGvK8dsRYh6FsxfvGT0BuN
cCqZSc643lAwv9w2nE8CC0hHdptj/Tn/Jta7YxdXmtRiBAKfVm7J8x4D7uj9KDOz
LeuDntqepzHN6S4HxhCrGJKPsKljKCNRzKryAcg3bsJ35OWPMEFjy+GHQUHS7HIT
huZ/naZXXI8fwmxdSBN2yJSlczY00FZV0Aak6Q60HewOuX2i1wHxSgZewo+C0Xgy
3s9e+hhjBYxwVAJonH4RZ2HCsDOEB4YzIyacWj5xqRVmV9bV8r7FlFWLLwdi03ao
m9MoyzvBVrtyN/6JQYzf2Ex7B1IfhLuKoluci79Xc0bSliMqZZYqFmnqHuVx0WCz
3ZIpaCmRz0ifJHxx9T0Oq7SI5fVKNz6ZGXq+fOZlmG/RIbgigKHkK3Bv5trQw5+d
p0Wp0B7fQtPxVtL4dTLfxZz0UGvGEY7SwI61cjseONW2Nz1jVeU860ghJ7U8XNlX
fmhY2WkJ9aLHGxiltU+iovJXq7tWg30NqsH7sygOj9KIu9fGZCozGzBmq8b1Ca/3
JBhLSf7dWr5w4mtAhIkgt4seSY4EBznj/OZrDhppnh5EaEZYHKriGqnnpM683msA
KoyYLCNqzlLBgjcGophh+qEvsDy91f80qs5tHEgOZo59iuVl/5yMYVs3AxVomzEs
/glFViNXJZoiKgHJDdh2K05vz7yCOzewZ5kZoMM4/Pm3IjgO7b1Y5g31+mLM4VtD
GUQjxpEhVRO/vZVhvw4vpTnpgocVkSCLg2pJivbcRiH8S95Bhpe6PxZQbHNbQ8t6
tz/e6muCBq/bhGHUFgm6+h16jLPFZ6pZbn0mZz46j7y3hcF3/3gJXSQI8im0K7FQ
npItISh8gg4lZPjlAuOALPChYEgPZnz6exCRMa6VqlYBau2PPO+L5vHsJAQZqkGd
neZ4tJe64zkb6C3ZcrpIEpidsEJuc348rHBaAE7Vhohfn9BV6+tpWC4btmxxb6x6
vrLt4w7clqCAAcaNCBfde4Qlh6o2QH+YbtilPGR7HlXN/jl+otg6WzOA2fJMkHFv
dpcyNVf+MEAnVByP/p4zUjqgNf3o0mCKS6eX10Mp3JMOYtFOuFC8mXoftt1iekZN
bVW1TBf3j7M62z5MMOtbC8k4pRFR7TMGIy+VpdjQrZDAzYxG1DHzYq24Az1EIdTm
qS1Tbwmnuegt5fR2Rz6PEs2lemIeonUcjKAGSEvL+QN4eb2VHtRoEszGUl7Z+dEJ
xeyM/FGeH4Pf1Fe4LdlOD2MsbUK08MzLL3qoTysrXKbiX8ZDzUEGo98pGD0zrYF5
h8nemxdbUIT20SiqUVtg4512p5Vhwsx9bYYlIS0upRRsjngq/x1D9FlW2t2Zn1LQ
I0duYDb7C+u7W1OL7XO5YNpUihD+BEeIaLPwIWENQEhjUBtVaFl8jLuV+0wC8hdf
qD0wE412xhxF52o9izofqosXrBi5cnGqW4P4BtUOv9Z4GUmoYFAk6jpu9Gw2bsES
RY3vT6gj6UaieJRSE/8+a3QpCER8sbnRIhN7M0sYtDMBkL3FrslFBf6cm3YXK5aC
msLvU892BRJM6LFpyDfgl8rE2uScJUqr5pXr+WSyAx4YKr5n4NjD8N5he4CcULtd
2AWkswZPJkTCFcp3xUf8E3SnA7JNGiOgf+HxvoNAFcCqG4iK+u+FyMq20K+24b7B
9KHYCTQPBLdAHkqnNCfOHIT0xDpu0e+RfJfblwhB9f/PljgG7chyo/efZEYX3pfl
zZprFyr5Tl4PysXARbzxJTVIpeemW2w8ZabvKdIqSrbFiinBeHsO72XdRAWTxDbK
KX893CTE7zKyLMO0jiA0j2s5Fihs3FFmIZg8Yswk4vt0Z9etCPAiuGmyhgHMTq97
O1VPj2Vzxk1mQ/2id7/PesLLrat5Bum79PG2H/oaMWKd5ZAusKPY4TTwT6gzVTIs
RlrguPK7uBe5FMDn4VpKnXlXgzwkPJ8VBE8OkBZ9ZB65inD9jqq51kIXrF4UT/mC
D680jTUWhnotxIygpO0w9QWsh16Fk0PjqgQ+lO83opbpMqybosACH+5peudSRveA
QxImOiYeefpJZ16LXuxLr41GmFKS16dwgbhQ3QIcGyDwtpHGPCCZtvjFpHemAKiV
CYNg6GAZEbjLBYFYBgBq6Droa8KU0jfzNXahirZHqxZc+wFX9NPYQf44uIuGTvQ8
8SryPAEpwRlLBC6k/IF4SfAy+aodA+uldpCZkhE4ZuW2ip4vELPEuYQl1TF18t78
bLQWdCkyX37b+FEo2ERDmkTK16ZgPMB9q82Ot+u1pQXtNmiHgw2DYe3mmcfaDXay
BfDPJdgeDjytYiJvTPitK8MTnehMVCLHYLesAfSF7IAVOsEoR5wvOakP1BgvPOw3
akhGpgDeNZ1ed7kNFNsps9FNl/SJArh/i0GurmLsE6XEYYi6mVdbldcl1XpOzvF2
bnTbZ6v6legjb+VMR/8tnXkUMU+7y6c1kLUzXFhDrcr4vo5zWT7pFTptStyWvKAR
THezBBg+C7yZYgU5FInOwKsynebk4Xk8ySLu3+7uvVKfk/MYTxmr17+5M9UKpMYe
EUOhYs3v88hixaW8nZcDMyNMEEl8p3kUUCNyAtiM6fwqyv4doKLEem001Q/tMM3x
KY+CS2uDggvULraBlw2EFyBEsW4DkAJpW8m/DHzbTCXUih8Gi/QO6uBvMQsVjnGW
uh95IWmNu+eq/x+FHH22+RwEf8OvNp38WU0jNUVhj1bPBBTDfpWF/Cj662tRgAU+
o3S6vh0QjDL0fdqjnY7IiW0uc2BhmRKcc0PUkPve3OP8mSe2cUOk1cHBmSWNi0XL
WOk1wCp7MJk9FR50vQ9AlGY7sZBE1TeeMMiDyUjvaMAMAgeawfplDxhSEiHD5YsO
kGjb5sJG2ftJeNE+O32/Bhg5XHQsj0VlpwRbu1xY05tcmICFI+3ow1uG2mEPciif
cA6Bi6HScrvT3u46eslcr7AogeDLB815ueYjCtJZ5z6BZaoSuWdxVuQLnRuZ8cQH
PnGrtnL66Aq81ECibwXpOyebuWjQ02wICFpDA6rs4Lo1icwq5vRU2vB14YLY2yup
5g9/8GwzcKUSnAnqijAB19BOY5wpckdlWjVm21z0WNwn5pE9i3JtZWcofogc0bDx
5M/fon6pDClYISE9kc9aRF/Daa+T5LNqxi/6QryMT7pap0dYfBZWD30IMxmKx5cX
8GZoBFJkSUDOzjywmPW3oYtkJv0V6H+1EJYwLcOv9SyzBarYJIlUbn7bRfH2oTXd
O9Sw4mp9n+MmK9V+PU48H69ryYfQaMHmuhR9sohVaK0Gcw1+Uv7r60phVTrJAsp1
xTqT1p6ufj2UkTrRd4upe/U1qh20T43u1ygG8l23YijNKDnaUEjfrdDPzLeJtAMZ
umEF78ovqIYMhFhr3FXZp7ozzWaIlbLoZwVwCc5xGNoS7ThTgqJIBs9wngQq3uBG
uQZXKB8Xz95oDJ83DLXaSFHEau7QbFAuH28nfzC/KcYsnswOuAMZxzZ5cvsyHLub
sfaCNsSFCHf4sdwcZ1mbMfDVswEPxMCMTefaBM5NYO1nI4Ux2ozbA8v7ve8XgGax
EsMM3LosKUClLpTKnHuZ56r+S8XKzVd6ljKwYyNROap+wXpTo5iL/UciqNMYK+X9
tchPrfrK5FvaUt4pc3R1fcZsHDFR7Gh/SbYp5qTxO7uusNBwRTvl+4HooBSn9V4y
BoleOiv/q0UNDizaBaPIqehTwS3sEVKEJ1kQx4A2jBI+lv4C5sIS+tNHSU+enXqW
MxISx4qENkhE9Aqg3UhrrizcGj89NBQP+yG18uwkBzHV0w+NI7ciEY/4d9hQebhE
BHQaKCrmzVxYNuqKh5HGOm+HzigPWyixmwtxz7QtSjTnNwu6oxNCeRjNoAGgV6cw
1h0shf+E4M8ssDZ+ur7CRDM3f4zoc+XcvG8FgrbqkZK9M2Gje+ny0d8agLQ6NrWT
lSGz+WJo91/OWF5GiExzAPpNQzuBUAo/8tyFMcUTTgcdPA5VHKTF5rfi8Ru+IE3G
+Z9t+fg/mp1QZ1d9rz4l1yTHr1lIn2QEW3vO3LZRD21WZcsKY2r8zwxZ7y4T4inR
pOu6SPNMpUa4lq4qM3fwLdwG+FXAZ65C5keW8MDlBQMM1g693iS+bgi9q4UEwYW+
ZCutH7aWyBFIp28mSioASbyallvQuooVijk/3zTpLFtg1leL3Eem9YCh3EugVL02
aPlqVYzpULzY6VmX2e1qT0Qj3PmqH4So281GxIIBOsoCjHXsw+x0DGtchPSfIGLo
nysnpCD3jiuZPD0TjT05AYAZW8mqGAsHghGV1DDXepJyAsV7tEh9BCMsDjjkXKZH
O9XO6AVINNUYhmXqhwUVK1nb5+VS48X74LBC8BSlPc2ID4UbYSoFEAn/fu/Kc3Ra
9JYdXyOQDIW6see4CsrS9fkxuK/q/kt+fndskw2BMlxrnHstVwmoIiqKixROACU1
dBw/ZyfBxXvbgqS9d1QkevT2DNXkPGCO6DGJeVrjtdDJd4ERbuiUJEgFjR0uDlNR
UplR4l3Wgsyed/q3YBqNaCE43SPIrBpBK/PR1v2MEDvsY8g5Lskml3/6RMj9HcXc
BEcAHE9KcDvcwc5nA1B0SC9VPDymuR5kLtHL8b9uDmQYY0C9pNwf+kMJNHvmDcFk
iIS/cJxODs04Brul2tr/rfyTSrLbqMqXoYS4SqizyJ/ehm82eYjyVx+Dk04vyh9a
ILvv1NXSZ4np8zpDSbn7RZzhBj3jriE2f4D9IRQvTz+oKugrrP0DqpqkfLsbOZub
RP5BWEf1lLNFiEe2VWUsqTvHrsS0sIGMLNpG/4P2ixVIpGAzRHma1ll77GYltTyv
wHZdDeyGS/1AzpjIf5PWD77e/gaVXgpnNrsJBTV7DSeTZlNTuLx+SLu+bH/4JiTc
+Db5qITKPsk8L5nb9OnP+P4tPn3zfMXoj0eBJjCOqWIno6jjl5xm1Y+YJCc0b2tA
FTCZ+lefSpodZ2F4UEhfOduUCD9ZTioKqbhKBZ1cGNWCbchb65yMr9C4vqRpcY3e
2gXvj15FQosTydATA/iaVSkuiAVPilzn2tkDe5EwMYbadYhqfSN+nmlb/rYzBfak
h00COJfAb5n9SdEfAzRAHHUN3f/jZ8VMxa20V3TLuqzD817Jzu7+dR/INBFdgC8o
3bSxWYTbbilpzUaLM7qhb6w19PygeNqt0lLOFOoKAeiuYrN5VGk9lpWgVp69BYVf
85qbeLBEdli+5q1dHlBwrQIbN942BbIwzfqpAVC61GiOlEanYKKnyVrVUuBdKrdH
1sMfQALNtDW8IX1bti13dkiD+YnTiAZVdfaz6zxIMOhIeLFtMI/GZg1rZzmaB3MY
+u5NR6cZlOIQ4IBA09V7z7ZlAxy3ay7Eqx+UmWdQ3HP/iRSHtwsWYOiOMBlKprRZ
1EJqAwVCYdunYt0SLIJsu8EnlJiVKehTR/b7DD0OodbXex0vZOLkzqrz9vZS+Xnr
O4tC1Xk655GN7AbGm66SVWPcre/v78iIyveBOBNX+27TaYwWDeFINODma2gVyu9f
jhvB1nFvCMOoPaEBW8HNI+zIZ7JbauItD7/ZVmE3VFqVCwLT3K1B7HdFe7dweDRg
2EOomVufIrAr1kTj/KmC33IH5rJvvmWw7IaSJYsv4Xl0naT4CJaEuNk1ukFiSP3H
M5WxDF+CUOrmaeTn6klTE4bk73LrPbENJDBdtJzmM9iBvEhuUMyPY0oSUq8/wnWd
hrV6ta280/aC0bHkTYh3UT56bwJnD9WG27XuPzHulQGjKUw3jGBN8D+XyWQQhcdN
61P4kUmKm8OBK/jpjXXIOIkOKB1BWy/euR5lsykT4rV8t09d9y7HT/5i7uxv/spF
rOPfwdcAg9PL9xqly3jhPlRivAFl+zrrRa97hBklNTFREEZJSlmTzDDkEJRM8US/
J8CZgm2saHW3WjQlfUknPTlRwf6Mvs9yvHWJqOJBpqqXGZfh+jE3480b8saI8jbT
RfFdSxq77qFwTeiFF4U5C7T3i+BJ+sr497gHRp1TBeHDmZ5ezN+aYWIxB0cWEXGt
rCquxn1fWSGL+DKgfniqQ7+vxFG7/i8mXrZrUhAGAIbYT7lIqkAeeso+Ppvwb5Qz
sAFWI2oJ8JyKfuwHJJalOJgjeld7ju9BuexHNPjJXRBvavvsx16TfQHrEv+qnUj+
Q6gSYBbseVIlMRXr5zog9HTNZK+5FsbLwy794FT23NOB8TKSW18ywhsR/oBzhaEy
ZurWfgmkjgRtriIat93Xew7xP0bIzluu3u5v4P+4a0EZ7LeO9gmHzlubu1neL3W2
49DpligRpdEUmpTlybIwU2o5t4tfximD0TRudEa/+usM/3qM2lyIOiYFQUbRDDLi
WUp/bXyxoGf+yEESGmxFqAeax4OO2QTxBLWe077+69mzgLQtY8uD2EfQci7ytI66
5naga90Mmtnw4124+gJiJaxnVL3asX8LbPqXTLbDIrGKN5F4HA3fBmWGpQEN5AtV
VdlpaEU7s1WHADrdGp4I5E6RQACqgYWP/FEvDs+k1lBet1FhMX9MSJWBzqK6u+SJ
V2Vsu+dZBv7kWDQeeFtKsqYGOcK2TEJ01W1gasOoSJTgaJf6BWd31Tx6EJj//J8v
wfxtIaUMZwMvrvobwa/hcMVu1seQT5FoLm5Ga2TSTv9qiIdO12aG2b5jpytaPSbd
ENCYWBmQqZYPPcZGmzhnMRES5i0teokzwyJb2MVN3j/AT+D9uia2dSF5Ju68X/XA
XTNiFDcUoWvqXbEIdx0t+N88KxsmkvN+d3gVOJ5GQKFG9wPXs/B3/WXQKElzudlj
upLj3oj6qJOT6lggYByOr+W4VbpcxgdJKsxfeHq/hqZ7ovGUbBLrV7yPYARlFmQe
jclWemzx3h+F6p2VvtOTLA10dPPZOlbQsvBgrelpXQISpAeX9DFFEjOenPK2SPLL
osW+NfC5G8L6Ap4dUN25WwShquBTeTd9k7XqUXTkr5SuY7Dd7RZjgRmBZ3Q1S6Za
udcHwDtd4BW+y7A1UDxzkhMI8HXqywcR2MDdGI5W2Pf2DMfdiA/9PXmTDKOnGYj1
57gR6bNvQryruHtEmMq7RKlfPXzdlsBLFdGPElbXNwOoNuTUsUk3tAaYVbrXlQnw
EByquCp2z7Uk/Nolu2RFG6+kUOXPGGm7lw/1Yjl3EzAsBN3WeIAD195JXVEeB4Dv
ofRmV7xQJLq5XS0F6Dzh+STGYaVh4YFHhwrIGrzUGI989EU63oq4OA8EC3Wg11XN
s/kmxmKo/iY+vgxj99S+tI/BPiDkeK0lR3x+n8CrxCT8vjVM8bEhUQScM2a4+Blp
oGScshtRvuk4UAwJg17NSZev2atX/I/gMoWxY9tTMMKjX6OWyPYPIvSnvUhKo/um
S3WoZ8R+zAVIg1CZOzQvGsbgC/R18+m+7Cr8QZZpwuTonEZCNplURJ8D28yY9uvK
BJQOdYcuapiAPv6TM6a+w7fNOSnfE4V7eGcsOjpkuajRb1BQ8yRSJxqeJSzGCcrU
xsD38Nu6QZPbyvn32wY+1KG2tK46xfV5x1NRT0sdUs8nLoBr2ueKsuF06POoiWhT
rGkuXBEc60zJGn6DRLMHezCBOb03HCEOmn4jQhWgHSaqVst+iUFAckNF0MV8KQDm
5iwCoUI9SslKDyZZ6kWozbo5SFo01vuLsPvA/HediF9z8bsfDuedB+g6kd6zRlLN
UReGv6BnWESt4bVjw6/r3tx+uRo9+ui7YpPwHek+U6FRd8LwmNbhCCQH8H98M4vh
6LGsfKvs4ulPQ36NScqRUGBcUQBqx239i6SX8KWprBEX5pt6buvUOP0k8vxxHyN8
D4mWlSj2SFAD1bC0ICXe8S7JHkzJ+EBtqeAGWeVXauYqWimgINdSlTQXPDflsB9i
ugUkadHOJV0EX0mFSkZhb8rneD4yBkqXFLY4w+A+nsns0ESj3mVhoMYkw0sYlf5x
5Sxgb72hePq06lNl5F3/81bJlUBtmNIwIrh/Djyw32FI1Gb3a6saDW8TWEbDRnV0
rX4TXrKQrRHm8f0KzF/HbqP0SH+Mej6FeoojEN14wYmAAuizeRqITC51FzPeRk+N
SNQzyIuRZ/3jdVR60vUbOr4NI5fPO2eju15R2KZx7Hb2Hf6mvf+zCcL//Mo/exgH
u2y6w7Draj9xcAy0mfw9gBJRz+uGY/n/ZSSbPqdeKv4uT+i8ac5M/mp4lDUpHJwi
TooRpfsbM9O/a6Sx59Rvwez+3bdpXitWxMHhZnNmGOMZLUVvBQZawO/aEe1FXi+s
Bh19cVOuiVhpGRwaSDBniq3OP31rEm3DID9KSCkxglv2LklrT0EHYdB9X18p+5px
OIe2nn9Yt8y4yxxuM3G3hjWh2YduL6/tGIHXi/gFKh7PUuvhJPZZXo8sbtyQZql1
K1XEp5ejpObN1vkZiyIBL5U9Mpj8PSobem//cZG6NlhC8tBk5fd6UmUFGpXlS/9w
1jHWBqTWLkNL8Ege1Y90/oyp2YQSXqf7nXos5uOB7LMt2Q+WvWRwTyaDxjibHth6
MWubaJGybqZiDIBsZV5p3KmkJOBoJMUXg+M1ltDtGYEmMFC23DlUvycUfydM5KXi
S9EHEn50ZLu8JTt/ouYxPHn8WKts/9Is94BjAtkqZZGazieT3KGGZ8e+R9QBBn1V
vL+8EDohTAq7P0Omq3VXnJe7xtlsEl5xjByo1t2N0jnqJ8gbQH0TrtxfGkpA8+F/
Ksz+JqnEFxZILsfmIPKCdJQQFswCuz3Bx8NYJFt9klDOTCtEffjwbOlmhIvESB+j
qlwMGQvuVtUgyfWrMe5+tYTWXoRL1SnY4w9E0c9xDM/pGj2TxtZzXUw4IkWvu9g5
c+PG7rvzhMv4800A4PclbNOoqE+291W5p8dnHzlN1XoHrmv0a1fFGqojAAFPlgT0
XrqHQIyZ8TL+9pITR5DFBp2x0k/VHgrtsXzKjA+W+C6cBTEg2rKSyp9VhdGvZWMy
oNIB8q+QnpeNGZW7i3J/sNdvKav8dljZhEdsYmECsM+JRvG0Gf0wfSLKyknER9IG
6JiO7/+20PEUkZ4lFtUXwKyh0JIBZDnk8TWZqOXCG2c95zbx0kZgEAyrmddCjNh7
A/j6q7BSxqKz9uAPvBLNlKgJE8K9IH7kbJb7Fkp45XJmMyRltWAWoXrAAERsXvhJ
v/ipp9FGEcYbLzrtoCFbMD0fOxJW+bAc7cYZAwGjhBf4BHPP5SD51LI0h0j+UuW2
ZPSkg296k3tjOYvmKLdAV2ISOVVRzKh6NUefhDMPeyUUYlj75CGd3aOkJwCNhuGV
ZPBhzwFxwZ4xyfIXP9DYhZyQnVDRkGAfSzypdxrLMzaRM1gwWTiG6Ll41vIrZX8x
dGHTxVNUXaJ9wTSxTCCGt9K9pQ/8P1JVKZal8yPGXRZgR7DqkEsWc5GkPJRwVxm+
oduO9TL46xWi7sEDv4LCs/0UKFl0wqsNRwibAERz80KNK+mwumle0WCn4ELHStUD
1qR5ywn0BbE73VzI7rzLUtTKgPKbqWuu8tcTmjgatj6KmGToOcqShAm/4cvbR8aJ
MzAtxvFvB0kJD1gj/GpBWU24MWfJOlfJYK6jQyjel1QK8USjKvYCQ9lPjLtyKJ4V
NGZOqAgrS//iw9oTgcNDHvGeIb3KgyPu08TdYxCtWApKKQfS/1UYb98dD1f9ywjz
T4S48PFZRsaQe5IQbU9Qn7E1E5EmL0llR8L0DsTviGJy30NbUQ7l2AaYZpLxjSYf
OpcAnQtu7jz3ytbG63kV6oy4hqCU7fXNSuI0IsAlcru7hnaQwg8YvKZtbEKS/dIF
OKp0sOigS+QMGIcF45lqacK663gKVUVscXZDASpOiEj+p18J8GKxo82lH8+o75qy
gwgqGC3BUolMJBEfZKSNg3tNbsY+aiJQ/eQ6HaxA1t6OZyzhDjUzkDcgL90Im/GW
0tR+RMWXLRm3cCO/C3+NERboFJgk3yQV6LRONiOu1hNDW4M3KIKJ2TxArBC9bJrk
oC07nZKAPBk9itNW+2v4WbqCzsgYpkddn9w3A/LkygPCzixueWY2V5i6EMaR2ZeV
fiHlRBFKL/AD0MkZAvEPVnUF/2ElPQUKCspMnkyp4dclSUGLI35Hc/BxFR98GfCZ
0I0HcIrYXoSbFwioSnvF0Kt4WkvFURzols6C6NGNYl3Z43AbaOn2pfcUktZhIrVO
+Bj0s6d5mSDsCRnbJpNUbjM4De2cEwIKPe+DRPeak3do5Wx8pvS7AF2DHuqt9HM4
87yft2Lt9Imt8bUaZYWtMIHZAU1XzkDb22eLdHa6kkigOT+6MTrQLCxl6iRaHRdJ
QyZizfJSNaaeEUlaVnhYFlQXfnGOVvmedRPPifpxcCL303JK2SW5LkVe9o7cQ40O
xDZHnrFbGjGExtcjRufHC4hOQ9Dstr7ho0b9Qpwzn7ew0pTM7liH524l1h63/aiN
lcqIGqQ1hcL9bwt4CR3WY6qeKYOW5Ru+sk0fms1sQLw7ErjCTYBURkcaKBZshEcJ
DVJ0cliYf07lh/YQoIqlpz1hADvaDzrDqCzxVGkkk8icnB3jeaXWrRgXUMun3X13
9C57SYrjci9eJC8wXEWkl1830Ez+f8JDemtHjicNBCKdj3ldniTlGjdecRyNtL/V
qav0FQQOR7gBsvijZvvJ0vT9xDJV42wXrv4JLaeou7WRdtsNSF1XXnu0H7BLKT4S
rWFnebPtWo3KzroM7cVyoo9QNVDaCkmAXmyVY2qVDfW660F+BPCVIKHVBtv14PCf
uQUBAPy+xmc0iJ7toaCkVXGXlWj39OwwIhTW94GGNjiPM6W+QAtlXVuRSFdkvbP8
5MgwtjxBOxUy0ZARVra4kIUOVekF3tQrsB51Mv6DCGYaEADnSdEF/z6tHevap2I6
shmQPTCjcX0LCXVDysmXCV/69MqmwBrmXxprDU1g97DdSwHgZxayDQu1LBA1TGoJ
34drxlBI3rTyh8BdFenT62ZlCeV0NuUi2UyS9G8yFKVFKhwPb1ll/pa1WnLOVdz1
OnBA7kFJh8X1/BvBS58IoIaCdPebC2Fy24GFJo0+pD8Va1LSCCO6rehH9urNpi99
QqaIqrI7WkPQMyi6ImezV7sqn5nJMC0xajmxpmEAb2dH5YeJXPcXG3eusVGlrGfK
Aj4QN1b1TcPPIY9wWFmcTlxdJ+/lqrv7vi5ONAPGnvbZQnD1v6JLiLcwWMzs+4zq
tirCOTxhV/D522bTuKEU9eOlDWt8G4DQzZp11wsecTaT2jIIg56KKR8zluRDTz0W
+EeIveAA06d+y2Bgwv8PUp+VSIVY+qZZNS7o0wPDLmsX3K3N55Mqs7L5V3XkMcdl
eIZE/148SkdZp6ZSPydx3lU5oGomO6LhQnzfYUYtc6mrQTJF2Bbgyzc4do1LusCV
Hzlv0fp0sZKXWQXd8ZnYH/7uFgm7CQL3xTmQx8e90KQz08CEwJnGSqlt2+CqqZJy
lJPWi7RM+ET/4otwO83MjdpEVczorLwETvEekA8+Y3VghFwlbyOcRooQPH7GSMMe
Jsc5oqKFIVUsHFs4m0pQG/S5SbmAu+kV7tfqv+8lsAk5oxxy6Ev59XREEdKQPWwI
0fmGpIKJj1eRnVh8JMIHd3JLtrh60JlGkKxi+LdLJ6O8EOWFQuXYRwM7kqpoAWBP
VWahYQwSEmRe56KBjZHcce/ks6ywIfEq5qnsHNciRmqGdCCPKxnp4N6lb/I/pqOY
lVzcuR075o827xF4LHmFNZpp9neEGd8PPRxURm/IjvY84kMzKcP1EePAncsbOZxT
TTqCPArTtndne/m3l14ePWeFDE9f2kiM3fcB5dRLlG12nrPrJLkA7Ppoc8dsPm8C
RegQhRgjhuK6ShH3nXRfYOE1mxsB5Y8BG06ea8X/0J+/z+Dsx4EIahIYhHdeWGDz
w8F7U3rgS8MNaHQUtaDsX1GYEeSpQbHbS8QGCce3if2B/vU22YMhGL0JeRpFx68q
G0/X66KF/HbcFMmnrCHo76CVCawkG3C1aa2eawpPdxfQ6IaM0XEJF+XKo3KOw8+7
pHkzXgiDfhUka5nV5xBz47WYDn6QU11xWUFn1qBl2Ox7xnXxtONdoZamb0ImMqX4
ST1fCp2zQ4PJHmmhRk+5WrAvLbooPIGr4oRSB6zjPHK4wJI0+DGgQFRoYKpuNKTO
N2Q4X9nBe/D17u24qlmitYmxt/ag6QwSL91q9S2DkDqTOnDBQpciGDKuJKGvKdGH
t3vPKQgGq8xIyeHdiwlgF5B9oAtVNVuNd0s6PBi3AE2RXa068BBOCYn0A/F/JIx3
IkHF1UDnKhMFa52RwRY8kIg9lBRIIa9eT7W739VNgayhf8vtDCSCFeQJ9p3wa7TO
+9jpKolQ5EaJWqQLWsF1hO0W7qV4MLpLXzr/eYbU+szrK0AgOxPzNNQ+gGpX2CY9
1al/+Ut9fS8RQCnktgoLcAxRx8PmVElFSE6uG5P/DQiUobsyToOmuOhVsuEHRah+
JANSvuQ/IZJeLZScWStYT+krFP2iA5F5y8P5o06yHtmA15fNRmAAxUu1K6Thr3SU
UBI2zAdmmqbvZKFML5o0M4i2jM4CjinRcnjqFERRPYpQn9FjqvHZ90gMdMtyUInE
AJlhhEUQchihPncvoObp/djZmovQER8GhpzZUq4jGOCrMK48v/I6hM9YdvfedPBy
spZ0CpDOubdtzuOilg9V38oPt3hDi4MNKLgNxyy70QKQrTRPnYAwXJU/AS/8lIAc
LtW+iJLsnwpg1uGmfghILFqjzmORtIxkEzO71ni13UL7MGZJO+zkToU6xSF9hraa
V8QWISA/kyLCnbYw0jTCWDYZmMXHtflhbmFeVLjWC+zXrVquOiKgUyEKkSfHfufL
88ic0anfs9lJ8fgBLu5IFvWohOxDyNUGE7tgrCkT2atIY6sKnG1c0JZqQPNTcIUA
0QJG9cxq0W26zcZw41jf/X/eCwsVjExr/t7J9xvo3pX44EToln8s9FHqoE+jMff8
pIYg1odvKc4k8SU2ctuyEyD1aK548vwmAa0jVY9StEDMQeGHi8kbeaaNTN38sXcH
MjfqGiPS4+cn0gOwe4k72CDTb2vu2vwp9W1SnU1azSaW70UeoyjC1ccD2R/btQRj
GvAlsmpNncNlOom3POTk6pqquF6JAg9sXM+FH09jt4MLL6ckrn0zqlJ9Veyhh9j9
y4bgREbNI+qNWyqAbMmIoh5D6Advmh1J8EFqNe8LvWNn++TsHXB/HhJQ4t0Rl8E8
CbaDBihQQgFGuC88gRCP5ccSU7s+UKkczHfW4i056RDP7qCRlsqINVtaKIz+iI5r
INbrLPTtZ37tMWP19xvgA8TVufPrBovykhwLFV61h1C6vSQxwjDFphEnHfDnkOVj
VDAw5+zs06I39StH9g+7OwE/N6W+lAF84oaVXCFx4gGDg3NYGt/Vl6rKEZ0RwKTy
KwattFetgs5Dd8TKaqu0L2MzI8jQUypXu6GrX6ZYYFEvHkuyeSGFGP/Io3m8+ssL
/8nJc2Wi4ns5y3ZugSzO3knv3Bwpbq/6KTiaLyu7m3xstpvKWgMgF4kueVX+UpD+
TherpYNxmlswMrfkXUs7gPy0JSnnK+2QxxHhBEiQBvg8VUTZ7enYqq9A0uFsaSeq
0BABP8hc5rgJTcYsZZIOfkPVypiOGxsbo9zN2H/+ei26xeVexxEA0pu9imzLIa/H
RGBZEckRuGSPdNbuyzRb8rNzTEHrLJgIcnA9NIGhbKjIQIEGgBnOj2VKFBgiEdZu
p4O8vZLYxj9COUhG0OQRSqwWPIx3czDXnngUobyj81t2lOrrsewkhCtIoxDPcISw
QJLgldHgnoKC8mFsFg58vWznDCkx2WNT1BmNHVLADwStuR9MwOfavt04kvvFCh2n
DQqgwd+lOG/z4gsGrJUdMqNesDwE8483qdhmchtTVFYFUYEKDYNUyTwxuJCn0Bvp
AAAjBnmnwuIqhRg/CNFbxg6ZpfL217u0FwYwKFcSAsT27+tUwZOs2h7Fz4iRCmE1
oJ9Vdtzzt0tzdctMkBxHbl2z9HPmzQvjwqsUIilhFIikyl0CluwpKb93i92WekF1
vJD3kVi59Z8u9z9AY8/uA/Y2FFZPh2eZlDcpS7OjPl/OD8udQt3TI76ORTKxZ3+6
cD7Mc9mc0L2XTxcNFa7dwAWQJxhdU+KnVwM3cJSK/pnT0n9IssxO46c2Q39222yW
vG7OeG/jekW9mePm5aOjrUYg5FMMt5I3iBalPIS6O0pXk/dooDmJ9MXL4j4YqjSW
SMuMu9Vi/bfDVK4G7HIYrm8VW5FSVUaT2jfPQ6zgYiTfLBBeStF6UcsJ/Tv5eCh0
AB6M3Y+VYSVQShhoLVs7wjHSEtsrGcJajDR0D5p1yAL9TFgKkkw4/7+hHHLoIATA
H8C1/vsWCBr2mXmDEwxm4AckJnvURb1wmflVbAEL7KletMQnlD+mgmG5oiX4+c4Q
dckQ4ll4JSp5WKmBEuxEB3htHkjzXWBlCmLaiPbRIKUELylHN1QBZ6rbIb0fnenv
dGmZF+1JdyxPjssz3YSxStjNm0Z35tl5lz6gsU7Lr9C6/MUxiZe6psxJIcws1YsU
5gAmc/YbMT8Dz5ehlXkM0PiuwLYkPJGYdcErcatJ1YwC8869Sr+bN9L3P2bcc7iZ
gQ+ox1yznauW1orWOxqDfD4JDOxOecn8330N46huAJkdcqp/n9MfBClITzPmc64I
XVK5oK91lzi3It0wf3PDws9M5RxUWtOwRjOoz6r+BIhPY4WCjducDpVtaFhDLWvE
iFStRKK3xu1/N5Ph7p7tTNbAQTQJWf3FKYc7cAm8JXpZtyzVE7PJWDuSCoqMb6Bz
ybCGdlR3ri78tL6HckVAjs0XVHQn5sqmW2gN9HrLlmH4O8GNxmYkEmFSnDewyFAB
mQOzi/DgQa+wV2vQrsgmGcK8RT1Z1t/VRvBJGxy4a4J53iblRqLTOISAL+WhOtqx
Qw+V1Lrb8+sPfvVdDme00oZgyjLQPN89p7AYWkW9hi79i7FAZVkb80acVlBr+QAR
2kHPn0o3ZKEsI8KLT+4cSdAo1+3yBn+GQKKIyNfHq/cNwoR6Ox5efoCHIsjNGqlb
lKi2jDzaWeSxU5kZo2ZfK4hLtsMNipYe+zBzJwLK3bLcb3WHKEmkMabd3ry/SAn/
+h51FRX3UPqX018zqxYjGbrJLsNAmWc8Rzl9dTJYtvZlgVJzcOX7XY05QMoL2pFI
zRN83g3ALHlN+RJxLsS76vEUKcgOfqQnW0+8HkbWSXMQzqVAjKKWGDEfi7N2iG0k
Ct2bAkInWsI+abM7//Y6V6x3TSqEw/zvXo8y6YgVLVQ5sQBr/7xHXtkwEJXQrLq+
JRlES7u0JTOcebdMTEiMLTp8xqTVYcoBxNEwxl3n+3XGWyoDIu7+7xyiDesyDaX3
38mOSAVND9r1aOhl2NkV0MCwT2eIaQmJYx4ZO0wTskdcUzPp8I8zSXYm7cs9Bkue
5b/3fa53+W2CXD4zA/EeSTxrZTzuzjEyag9dzhG/xmoUUUcHKsp58oeDZMS846ja
OZi1z4tXn2YewRi9ep4RAZUjaniY+hYIPDLW6shrR59BNVRtzmafXBSKhpi/9+9O
67SxTM9o9ME7bi1QAjhF1zmFULMWWAR/VMTnmvEFuReAyaOFPgpX+nI1h/o0VeZ+
v26PMP3TSAKvvv8TiY7+2ZCF+dlbRG3MVRXy9Nh20N+Wqpqh0OCh0goPBXwhadSy
lQfXjjM2sHkUFcvw0l8rnyhE6ClSJH66NyQvR0tupkmZq2maPuoYPu8Cpmf1dofm
ldkrK4SYwdt0O2+hdvn/TknRazfnmKN545xkp2yLb4sOYa/lm3ox/zz7EdjQu3et
G2KoeSBMWD/wtfeK7zThgEx02ctG/DTybKPgZVStnbuqNrNZdy1q968uTCi2+/4K
BX5eamVsViq1R4Mhg2OOR2253XzcpafCgakDQFUCodiDQPaL76WBXBOuQs9tfPR1
61ZDy/10nWxgd1TmYlMF1zOzoCeaKVADa0Q2XiETYZQT/rh/SRhJLfFhWbAI86x1
qYeVGTHkQ06kiKBDquV4Ik9xth5wmHQyL51yk1nXw07LWDc5S3vzkT1zWPgn9CKt
ZyUHITYFxN6bKll6VeSPb01/D9x+jWU++PbER3G+3wsclNFuebRQavslqucOTQcn
KmeLG2BVqwKiXmHkqvOaqf03MHC+YS0703ft0JffEHUyAQkteS9cLrYj5ZmogSnK
F5vv4cq7wCUqi2+qenU1tdokXpTeLnOwH2Ko2+jIMpdAu6FEBVUS2VUJg2+fmALB
c0/Xov/lHM0mCyukyCPVCU7lHzounHMdOHOcGvbOSzYOO3oHB5KbjPxouw0Iq7+B
OEuhgdMrKtkcY6jmia+L/MMqw6NJ43x6mObECJbm6VBN4oWWJ99pgXN23nB74fbV
g/imyMRPg37rqbPTBsPE29T2QSBbjLK+XoSzYZ9aXIwLVW1I2gknjnLvI6zOyyFz
Ancy42tDRHit9WXkBDUdsx8SEjNWB6/R8KWT/JiHbn0gnYMHVHnGmN5rMHA5+TPo
tTaG2SsPpTkqjNUuQZvpMPQ2dsLWkxCV2RJLn3yYdosyNhAMxfgtWY9P59BT/Kbc
Wx85Q0H9dKVx+WFWcsv4L7Kn+HuZ925E6N0IKl+WKl6Wy23/E8FSyp6ivi0j+YkL
YEJTww44AzTLQi9TbiYgTNllxN5cSCijfQnlJfFs2Aysz3s9yFd0GmsLd2GoFiW5
GmAM+r6596fnaN+xcWPuUrZuxrTNzYLJubw7f/tGFeV9xy4j4mm/RoBqKMr84wkM
aVlUtB8+KmjSvpWIBCbTv9agOBZRxKetyyZ72KCvu+q7/CWE83PhxofJgxWo+UER
wnXrq7Wid6XMRxK8xi4kThF8SYvykEuFKGSnjijspHmjIQ7PYtnUP//42TY7VGqp
gXAmLmQMgeWKJDXvWefu7pKhqtQUG5UtMtqXgHrTi+30VW/srCR9zUVLa2Xaerfr
n2AGNlIc59dpfcKZZAN97LwWK1NS3atSWD4CzaycmEhMgmcjWnM/WWTHyIxjeczd
GcmnHKAPwe8zkptvvQuxXmLdk/fM2iQ2Ytgr3/MqjufZeQzYqmDGfziJlyu7P2jB
IUTDMkzl10cFFajvMnMdRtNn68DhmwQ78TIJDVAoQBVmXHCnc+BsPsx3+UVkNCmI
lk2z5oc9h+kHoxAsjI3OEznomqhSg8/3qWnl8zVjMjE9wP6SdDZ62sWh2ISeXJdY
oM1gb1nodL2S3yXBH9tWxOv0ajk8Qe2tTBQpviFcAuvCrjAg1e6u9CUoqdoH4gmA
jzp93STsACLmXOPYbJWPp/koEh6bezc7Dk/Y6V2nuq1vBqiuCiW//GmdcAPtdHW0
Ea2KB2Tba70GpmySOxQErdBZId4B4kY7evyZtWBD1Ke5rZXbnleAhzKdaNedKdMo
GLiSa4l2n1SsQakdqpzxPEV/92BDQj+SGBAi+put5vBcqp0f+Qy61AT7+ZHnaQdt
uMa0yqkD54DVrreEUjrrh0pig9aq6trQ6i/H3nEP2/wHSyW+oHztNte49+UhvhGl
Tsd3kZh/Is9qY1Zsw9N1CYG3W8qT+//v4q7lTYeqhbNcXp+OB3ZQ1oDNMkW4cOSC
OZ8l3OYIvRgCxmhvrk/nLrF3SLTJScKB6OtVnuYS5rCUw2So1XLNO/Ag9yDutHHG
fY6q6X0DsG+LPoCWb3sMPbJPHXZjGgH9oK/f4DTh0IfVtvGqRYElVfoWfA98lM37
dYQPndqf+I+/U+yNBMi3UkjpEL27nttCIN0E8Incpd73dwV8BnnT7dJNva276Pmv
P78ZawZdwDX9HfOdrCeWiWrgrZpLiUP/3Tzl6GxNFAf24//luveZn1O8cinNNAh/
5n0JDpC9Ai6B2BIA6BEcbZNu/ihlzw7hIXaXmBrcTWkNegRfUAU8xSBZTzpPIS4X
S37N1a/H7XFf9KB7h3Z7E0pol2UAB1wRw65oFGuU4akTFUhwQspIKj5gyKHfeX8i
T5XmSSpTY9JQVY1w+wuNWCUzq3a9dk60sqZ+iQznRDPMZ3KkXzNtZtu3qQUhwjrZ
dAGfqT8uky4o82egzpz4lvtV0BweMTFlGb5duM2c9BNzjzK6LDcohOxs1v/hAn16
VHMQEOW+/DywEinzYH6asrL1bmpiNKHr8d5EGnAGen2yMlsFnLc/E+ItHC7q9wed
h5A9fXFRn3hczBng69TYJ5zMXS3nuoePsQwzYg3HC5dYRhQEwBhp/HG69dreaC4a
D9rG11Rj0oU+njm2y6MgUZtLDXcP8hQlkAJxpN2+UaIIH4aZ4vcDqBa8E5R2YYh3
mfzSkFG7xr+rw8pwf+NCso2LY4myaSoWvVqBGX0l/GX7d8d4sWjK70Og9HsfBMC6
PVDc5b69uPbsaN1vftfaq7HclNFWXW/c4rQ2YkA6qW64MuVrZ9/NzRgZ1jouqI1X
TsyQPS6B5P5Ube7CduAZLnZh+Sa9BwFzj7Nb+DH2xJC6Y4eMybXep3ZFEh8eMGal
riHEb9MKsZEpjtwK8PpFJDoCZW5AsYzBB6mZI7qgTC35KBYXYwYGYnw9SpKosvCF
TH1gyLthQbPVWM06/NzbicOdN2jORlw2/sZaBGBZXMZkNZwwApONorb/0B4mSn27
oHKM2WhQYaWq3otJ6JMFeChHsawd88IhhSAvoj+J371q54sQUzznF92LS3AVFTZL
JuHxMFuFiIcPHdKx5A4LAdAUAPYPQNcs5EtZ1eiH3jameNIMkab6pWFM9J28Z87r
SQTTLKlBkaN/bft+e7da43eAH6Qrq+yQj5H7he5jWzEcW1W3YQIyD6YuV0wkv63k
2tvko4nwc+ECidvakBIuvefhHPYCR/iq9ie+JpaVNWxDpoA8zV13NHze1pISw9yd
qiAalqNHFc261la95qKJ2jxaKWsvHqha3IaJd9VMswqNMFdGuhooknOvWfUGipMo
ALV6/Regt4I1b45U6mMo6a3VdFybOgpNYk6n9LOWqxLP2flWzouM/LUJ9acIxmfF
JKDCI+58jxJz7uU/wIbO9wsGskq3zypQTOXehx/4vYRbNGIqG7N/e5JmBgz7jatM
2+w71vBDWvRskE2axYzDYaFuHJLFodBrXgNC/8dkYix50nNwKyWLc7idtmh1v25S
7rrzgP7Zzs4lo//lIy0FfIaKdldW2aK9/7wfPHjG9gWyo3FrdGZIE3Je56G6sCI5
6zXjY+BD9OwGvkpBe4ees3kCeSDPB0KpIn/2jLNgep79MXbrHuu7G8nXW0VRi8bf
3439oS2CJhNeNcwYtF0IGVKoW4+7Z4i0QeT/t1+GxFzuqx0qQeJI7g0Cam8/XsJW
tnl2FIdJ8u5950XjljaX8xz1DG8e2ovq7EKNDSyLq714B5qDv6AVASzjeHT0/3rE
yYp7C+d/3lxoZzvxlkWK6poLCSg5QZ/eIC9sptVIcAoQ0xUMCcuQDchmINMVRs6v
24TLR3lS08/QvB0/ebLPakU7QDdTObPzywnryghZ8E6ON9/Jm18mOUc8M1ORJF1f
icNYyOX0PMSrB+IyCtP9nGI1hgLqYWWvzEcoTe4nu6PFjZTV0gY9Bf2FCk6AtIj0
9bOCze3w1bRIehh7/YQINhBc1BUqeJzR5doXVUJqxpsy3AfyXlvM9Mlhk8DsMj35
3I+EExjtNa+1rSor6/ktRnheMNRejbKMBh36eGhNc7845OzL2Qc4eC9CACa20XUm
PgXdI0uPdLgHhK5dLAGvm0lt4dgVeUxb2YDWzqLAn59/G/dV576HwEtCD2aHmUym
C/nllcfQSBGIK0Kq4SPOTo3WkBFTOIkYoyKLorSI1oqZVFirpkL6pN1qLFaOX3c/
glpvw8PWl3pISmikpLMoUro2zrtNnVCeJN/RfR2rqvEJzIic7PPV8ZUApQZAFvze
Z3v71wVWQnvH9FpU+0+kWBZIf4xcZHrCAlfeRJUvR2KWKb0bH7Qx7/hlxyldwZnQ
ewWMSvBiKmhQLOT52KO5wgJvyBTLrw5bldBBMuF3BiEU8T6Wx68mzjnwBfmKV6Yk
8NEBMlwI5YyDIGnSRRVKeRnRRMhOs8C0ocXl/M7B5stIs+/E3kxIjStzHvR2rpMg
JrXnIrmXvD7WUhEX2aFJpQvTwlpG6UfkM+qGChGrDSECMVc2SoZGuKTBjlEsIapj
6SCIj9jfrrek19psEP+QC238zgj0cN8n1CFxEta25IUcOofCHu9wHZtBIQf55HkF
Cc+WJdhuztVNWgX14u03ZZwyGWmH83XKlWx0PwIV7E0iNdQ38pmvU2T0MXbjXFb2
vbR6LwwMd1yq52kI3YTn+5qbz26S+30DpwwNeX0zW7SbHS9Yz6nlvvdXcMcpcsV0
afiD6OXWnre/YluFcPHhH86x2bva7ZHrmTHOYSUG7dFv7PFMm/FdjpZ64xU8flff
GdUaP+F6HcXkIej9x++Qp+p2X6106LaONHokkLJRNuIdeqmKuZbn/39NjhUr+Qp4
bf+wFx5P9trAzBQKvXDfHDU/5WwPmcASUYhJcQr1mDUedRXrKnC6vL2vppmjDIY+
IWUrBQKRGqttyhxGtNKOusPAudqTIUMM+uN8xbH2Eocl5gTjwS32wo+dsvWpJy6Q
BLXHJ9Y2tDmBH5z+Q/anoQzIvsIniH849ADPCsHCMO7IxFEfb/9rrvWqRnPVPfjw
VPQ3phDy+zQEdFlgSzRXeGuB48PLaJWVydQz8LJ4LqgDH1T+bQZ9kQqrkZywSwq8
YHiUi5gVJ/T5jf49uP9VNavbnimPw+cz7w0zCsXKWK6ZjN9YN20Zr1sf1e7uAwXF
pH2E3oW8RUGULfXQS9usPlKgW/WUydAfYKh5UiC/pXOrlIYgLO47ftTJjYD7YlAP
KrutKYG9LlXP9o4lSS0H2+IRlB4LjzVjxHcZ7BEMk6WU6vu2ot2uex4JBTALyjxY
E6ZM4ZyemRW6GsRV77xobOOl1zRfgX6Uv7wn6gMOo4XpuRQEMpeSIUihXcZG/iIg
PYuXrn2rmBtreLOmLV7WSb+AT+SVKJVPoPn9/zKeR3+YUkhPZMblccjCtLtdW6Nz
N8E7/Ypel1UWwYXqHsThouCM2FRbTf10YlNuBD2Y8cwj0QGYdH7t1CHxZ23y8uve
+M2Fw4u28wSeuO4YGQNKnE1PNYNUM0FElnYwD9f+CJEufTCuF1Gm2q+PWNkmlGwR
UVcpfqdFrf1yPosdgRkgqyj2T/FSk0/iz7rkxPKOeRi7tBRr/Byb4VsHd3FOVkL6
FqvJ9yQFXeOshUPdfAU/DHLRIJ+WF3rYDupISxkvp9ThGRyXRgM9gEEwbGhWyro/
ICblUwgkah3JKaMnq/BECYD/tVBivZuYGlueHkA1MUjwBhvDcigSRDyH0k1LMXX1
7pPIKYRRqCivnMz8eH9KsSlYt7TdvhEJWLWfzzApb4YeeydHubRLgR6qJNJUObIt
I4Zc72ReuHcRH6OK0nt7KtOK8X1b9pcFlC/qvKUzgWUOZdSiHweh+Uz1ixQAnFsT
3jzg0XNbPMF9gwRGRi3I0OfWkrLApF/gWICdfNWxiX+hE9AlaoylhlbSFZR/NXuL
vs0dtQep1yoqymZA8M56jJAoCzEStbAV2b4E04TeuMbW1oa8qs5c0UgXV8SJW++G
enspzw2ZU+zxzH1wZ5/hCyX7Blr66l+NbZQxTzQC5scPk/Eqz9MGiOYeCJE+ntvP
NCINKnnz3//kZ7NfWz8I1oklYLGJeHjPCaaP77zzsMdnvvLgdZqOgRv/RPxuVBCA
d708lbN/bf2mcG9bds35R9quP0kIq2QJJ/hZtoA7c9hGu0z190zC83waTP3qAgzm
UwdG16nPQCFcJbQXWJvz2d4Tkdlkz+o/AV+lQEv0+PHiGmeVUPa1qO9e1pQjdyHW
Bd9KRkERUE7DQuamVW52Ee2qZeBOr7Y08VdmykDYxPAbVLv7+LqzgfU7SP0HeV5J
K8BwbXdH9+RER2l19LKkpt9QX341vCGZPVoBThcPqn4b+f48w4n13Mvqd2kE10Q9
7Yotpww6gJ/WMqO7zUqS3rGYCVJ8cbjhGIh8o/gpDfkMz7FX4VcGl5mK1rMtKN3C
2D9JukDmKAsjcGkfSVtNek3RP7gEwJLjS5ib0uGklIjpSoH4dJ+Lkg7X03bI/9Qy
allJ8wcob4armqh1E6HWHK3e/0t1DQUTN8EWZVOZ1caHXOBeXNL3LHoAd22VY4u/
4QO3DdSMOm9SBWhX4L+AgHIEG5t9qCuqy5qDOBv+I/1s1kirvtUM1WP0OOVuYXYl
Axv2ifMKgppyCKp9uMRc34mJHVoWokoGbIrGnhw3eSCaPS5YKmBcYu+NlGqnTg7c
f6LrrYAavhF4C37cd6GQKkUru7KK7l85zE9hxGhVg5muvfFCdTnoPf5MHzJvonb+
Lo/05jlqENZpOb3TxC27eNro5YiB3qJG290L5aSFpbSObYVrLw2IeLIy9FMcerk+
qNh+r+6A0fCqzO3iOW+lcFp2XVu9adp3tjRj3RC9Q6vqkwAJ2OhVtbRdbzRtvzjO
wZwgGBnyaeftkUVetBchP5ZYhWFnvUI/GU3EGv6GT3/bGsEtY0vfTLwB2QS75+rP
1xct8TZ/I4mekhU8UhKe+3moNQRiRtbwEHE7gNtnu0DKrqIDMfT8s4x1ot4T7k4M
jZcloLKFcfPjzkQUm3BedXgXNOKHHYtVHznOiPrP7KBKkQf/VVxrtDShPobSwJZS
hCgJOHB9oxxqeIrZAOq7WgR5O9NqLkzVqeUOR5lUOesiLmkgoUNmVZYDjsZhbkG8
igv/Bz+cWC4H1VSIBw9e4o8p4mmYoPsYtoB+Whnwy/XKrq4vV42n92ebFc8xqxyg
y5pSi2jb0s7hHpjwIeGePHSfrEEBJQXKJr/qfulAo4g+kdSUzYUTGZapV0wYxz8B
WvMEjdrkh9ISzkxn533lPnNg/+YK1NjBqGZmKfQblYjYb25M5QJVWo91z84gsL4Y
NT7/786oGIFZjbWYKYaLu58Id6Ioho+4PwYBbcurlDCsBYp4TjlrCY2woFPR9AUe
mATQfuvumJjzeM5vXlpGVvTXM+5SsQeB4EWJQj6ju0bDPUYRtD95WfXv9NT74Bw4
2+p4xeR6P0/hBwEl9hy07j1y7LOHt9RxHGmTkIvt1aqCMjjNB4LYv6IyBWQZ1F4D
wBYQBRLp64nZ5I82nh9gbrky08PZiZut4X08URUVjv4Ne34sf9uIoo9zkV157a8p
A+PrZaAI4mQCghE0PYJhzxgkSO+imtZ5qXDLiCHnleIhaCkcW7xmqcnN3SSRqnxw
/B4bjxIp/UEpBb4D+3O4pGHyHqG3+E+EmfYuzkX/KaGseLUlxNEM1upibqCsZrVz
bEk6PjhtwghxgHRHfboUJN3JKmAoCG1OZ1vikR2tEyv+ZJID4+Kj99cA2HxnF+R8
3FE9N7aRP5RsZrFUoQVzgrO1zST+F7GjMSlW++QGnA+sPdFbnS6IbBzOI0iNZdC8
HQV4A09fRCCc4Z3iwTlVLX27sUNSzllcfx5WY9Ob5sBoCtzK9DWSz382OPuwFZ1s
nnypKOFMgq+LFLxfvKqOuaTtO58GgCYm6XEArQAABFRkYY23rPslbLU4fpMzvxSO
KJ/3EbRbvX9StWFaul3XpBh6NoEqq2XC7efW6mHRYvrvka7YsYw4WTu1ASdFITMw
Z0Xgz1K36yJkqaJSCByCNMxp9qLMzSsbB2BpicnPg+2P1Lj3ReAi0G028fVQ7dgI
vxN4Tsip3U3nsjgiFdXv0X9Zzm3OEL921NOBZHYLiLEdHIDdZCi/99NPOh5XG3B7
L0MbNIvivfiWGoOa/BJVsf2IwHNpYEZ0HK2ePQQmxx21Vtk/JkSRdEqHop50mFz9
5WpTTPXVTUqbt6BJcFUc713ec+4vMeUqodSRe8b9zkEqZj6OxRRaaQdkEkFVrG/J
Wi4XyzaZXVp5PJhO77YLhYaAnMzTwthdo+ijQxmnhIJ32wQAGoWn+c+riTEqQot5
7SCeD+ftAHJGjmz5F9OzH8gvVTTP4anPc1P4E5AFp/JR+RD0VXLQ8cBHMgqxR2vA
P/Pd2sxMAyLh9YNpWBq/8UCbKBaD57WXm706gRW+ZMdCyD7iWHUyJLOroelQ1am6
pP2NTaYOZfY2/1PGsyuAs4vsj4aeSaF0MA9rgBGiE5+szbczVG1IyK8spXZNP6Z5
AQFnXMZ9dR/Mvt1NVhOvAR1O6vcbZoS9BiaWCqrPOJRRqrp8+N7PGMjH0xHqGc3a
85x6wytdYoWro6thTVUjmkyz6U5XIOWyPEWfAJ8ZadGiw3S1bd8qKebCqTEWhc8x
CFA23+0KEdSZmsdH1plL3b3x4suSTHpTIEn1A9FE1MksGgar6ptlk68oq9WPczvb
4esLga5lA6w27vbXafpUS7Ol5siTPhsuDI8azBwy3tg8j5py45z8mxkfVCf6nfHF
cDRxXOiGhyAERKl0hkgFiXS+cF8yLA+USfZKpuFebHsC7FhNutLPHpDIFstQDV/V
rkWmW4uhSDmaq4Jjw6QXiXsOWQT6tU3PPWwOYaBGAz6RK8/skGvMSTmIHxySd7C4
lqYXrRRpB6GIKkae8OsRYWcW/gTcWzVPnRT8Hr36O2Z79xwn6OJIG7WHS3ZVLDI6
oJW+tuSrqXIT/vAbJWLkWN4X4WXClgTkuggRtujS69qXStLznZTq72VXZr905Xwk
xvmHQuso42j2Nz8GuPD+Gzn+5zBryuRoFTw2tz/ub3MlCQ9fAlzPJwQsJF9qjhEa
Fd9A9tU3tdOUw6nKmOnpACBGMBkNp2Wm5tGYWeQ4mn9Fh/0H/UrdI604sFxLPRu0
w8yCCevHc1YiCLaYf3MM2IMITKGfVj58Mkqdv3RhEUk9bnvklo7cKEA0FnXcJabN
z4U/ZPyU5Y7WKUQkXQLaMaR3PmsdlpCxAjaQMobOE1aTvCi8pONq7u726ZElQaVq
De7h2JwVgyqDW+boC7H4rBs7SQQLk6dRALW93uzKapvG4rW1cYm7a+BSCnb5MmMh
U8Twj2u3AC3FKCtfbekzPtfoFsIgBEHPkogKiE+mL+itxkhH44IDQDj15GzFAjHO
LvrtIqOTeUB5aU586ZWJJKzuFnIclv4mXUPxceCqqJYXGYFg6q9RHJPM3bsqXWZy
bWv1veL/w2l7hzpBL35Jm4dABx8mkgu0HXulnNIIlIel2ja1kbu7qLx6Be9OMeVv
FpstVJPsARgjC2eptPbjslxtdmmc7cog55laA7eSIklXZaIqpaDDRn7a4QB8JNsJ
o1GqZmZnRfx52uvZMvnEkr1aNXU8QaYH2Qx1U550RFBolVzn38H1bVyHqkoSRBZ2
Cp8MV7J7UavtuS/3DhWjCw5qC76Ek5Rfa8tVQolr30tPiXDBYXHP45P4r4GY+dpm
W+Xigt1cValvSjuA+8oOkmsGeGJaEZ2XgiSfgJA4Qg6Z6yDWBFSo1H2pj6utfMV0
KW6Cp1jLYhLkY+cxoSGGLh6Br/0OSmOHBm7gD2pnt00r+jbfI6nN4idw12BYezN0
mFSjwkjiUz7H7hk8/1BmJAtb0INV3m3x3+MLOC4+NlaHsF4AvO4/6djkmitzgVMf
bYFViB4qbhS3631fT3EWzomWyFQSKS1FD+Uj8LH8k1J4k2v+w0LvDbW8o1Hk8iaD
v74bB7goCWcISDLB+poCTh6cH8t6JmthQDpRocYgxAtFehiEUaUNuq9CakLS157q
R3FR199+7S0JkFmZpwrVF2Pont1oSC8Ow2Fbbhz8B2SGEvaVA9cYQ+r+zLWSxx1n
Xaojv9VtBmG3WX5fX4vjvr88t5o7t6k1XQH+r1CTLy7aFVRL1KJx9UDaSxxiZgwC
Z51vSB7N9bv+jGToKORVbeydsGBxPAMYEBsI7gk3zz8ttNT8Bngh1c417nrkV0FG
z2lU/OCvhgA/fU0skGf5lJ2vpkuS1gyTBfNJza/5ZV4jdhL4gc47wawXNN6iuNPg
3uYnQL/aB9s+NzSlbc8LqxzNP40EhHI304j7fl6V2CMVbngdz+73eJM2664NUjz9
iDxi3QQESev/6qHBw/+BCRIsgzVT9IkGIbbyKvQxBd8GvsvqRwJfU9ByaprY67e6
/dO8fVvzXVdY9fyRA4osJ/tBHOCJ6zoaqjfuzRHuWKDqAsNkTwu3j/cXDiXziG2S
aqo612J1V5E+yOMyM5hzwR+7u5DQbdbnvwlljpvLnKCQDtU09Mtj7aWu0oFtGJlI
UUDA0mHG/zgLHFzT+uqp8hsr7l1ZPDsEFtc+m/HVFD+tel4x9dZ2kOMb4ovHzMzk
tXcB9RYPy+QWTByrmmjTTgKTkSHGQH3bvLx+E3q1YbEGzBCojXuFD9/EfyfyEpc0
4E9fw0yV/aPAAe9QwRm1tFyW+O40OjOGEQF5bU1rb57yzquJAZgGaDkFd+rC9O6Z
+qwsMIi5PO9r6NKIhnpqBMrEgzM5uXgHJ6G/kOkkf4iXuEM6evt3Mzf/7M/wpoBy
ZDyVXPc+Y1le48MNoMhURzzydMCaJFpcyPOozGJzG2dkEWrnfZrHLVOd24OL0OkR
sG3IwDkvoB/P++aakKQWLV2djkqHd8cMKzsdAtAjctIW1sFEpKEw+sNHlbkV8BOX
svvKeplIg3INORbMFkozredYASihODutokYRLKk1L7HjePtjS4IC/iHSBIy8/fEf
FDDTVK1anASIsBrbUk2YVd6DrLnGPAOYMqql3y1Se87g4YwrbJ/a3+zrseobjWtj
h5di2C24W8BI7jz3iQTiJHbSmUtIgWY4ug0H2kH1BQR3xcHaDA34hEIvDBcXG2g9
MPsPfFzEe/EUA8FFa3fL+qMNAZZbIKmmWlSIkuWzGBKo8wFxg6kDiWyPFpqn2E96
sYvaAIW0aIrUb7EDsN3/QQDoWydJYyDthS8aTnTA372a+cyAm7sm4EStG+M5jAWW
1YCjlhAdwIDSkjo0UINNQakyyCIrTpW/uxbVvM/8FaQTOrYy+K6w/wrXJ/nn/P2Z
gvh1cL9UFuwBDQgvTfxIljXfzm/M/+9OVFtmF2+yEj8KdsIHaCN7hl8cHMYQ+Tdq
Oprb/wIc29Y3df69SeqqbqHjMcl+h2ZSz+N4wV64i/YWT1c1KOcnqbg9muxuV1Q+
ZnKGTJsEfmO0GSy2EXnHqLjSsrp55/m+U5sgB+z6FZ4+W7v/rETahoQVzkPpfYMm
R2etFiHCWPxyDh8SfOcKKMfO2SDPomvdHlnuMgt7AYYI7KcRzjBEol51IZB/KiEG
aaMaasyTpZhPu6mgKlEdRzT6iYaahYzfx+MAAMyf4qhgmRK+WnlIzoiqpDDlhzMZ
/a99O9rxMCGWe7rQlBXEYalz1kIfRS9vgrkGxcHviTvBIVqiVnrgI1DGGSe3aQC6
D86VI6VZbNsNN21ojvbDu7tXOW/XaIrwXAhhD5216ZOl5fcaqyK59nsecamR1s2r
ZWYAh1oNbVbgfNlRi2L3XfXAChsloAcTdXam0FYQloxNuMLAZl/sn2HCr98peRMs
BqcOD2ciniYHuOJxQgIZEsi2XISCSvOEMqbcGPK9V0IqAHPpBJ2eEetPXuefkJQo
3TLTZIUXmCaVLjprWiWYJTdnOL9W2vpwtNtJKon4Dmy+W0+7iFhDBcvIMhOqbmJx
43tKg/iQxfWYiIKmmPNGAKfNce3X6qy1FWZXjfKo14fVTI38UeWDSg8LoTi18UCd
9M40M7kWn/hCyYiLRNcUlbS4mDNUtGZNMiplDwADJ7dn5L5ImD/EZ/9EBCmAGLkg
xrk7ty2N032ap/cyN/He8MXm+EbW2zEbLHZ3SIWygtmENB61b8qJ4YKttRohiE+a
Ybv92PcmRiDlPq2VkwdCEK+NV7Zk25RawmTFmcJ9M2oXpKLdh+Tq2Qm1uMMRcURV
fZZF5XQBq8BjGCgjGF81w4STsXzicbVR1u8yqlcRjxd984yf0UlT2NsHlb1gndpO
wAcSo/JhE2kqe9jCVTtyn+W71FV/CgjQIg6eR2yKZJPSvIrbMfPDtSKRYyQOk3z8
D3nObckp+84eDqRdrKhsNzFi4E0KL8Bw12XW7zz34oQEbB07jLs3Z5rJTrkxnaWM
50oYgbcuvRXM7wMi8hqpYRX8BDN7S0573OTfL/oAakRMdUX9YYwF2MmUnkFE6Pt6
p/kA/8KSEjcqB3DXvPf/1mW+8yXh5Xzdskskk+eEhHLeEt/byxkAajwgE+fI4+cG
W1Ra7ypeUXk2svNEfx/9i2MMGFc8pNREf74JdyMr/hy42YS8K7RwEYMWCOOrdap5
5gWnPSNhbNfbyla5jyqvqWm3N0PwGAN5/bQn1ny7wXb8th/Up88kuUo9HqtiGYUN
xocdFeGJC+5El7X3RAmz1Yr7C1Sw99rUVNI494Nvl+L43phvl7UvCUFfOb64KWdn
7/RZfbZwEkM6LxfkGBCaMcHyxom5IGiV2ofo5o8xOWBBVqQYD2UahQFDJezSltLS
TarHzr5Cu2hz0YWRZAq8SG1p+TbGQa9YL3C9nGsXunpD1X33BCDX7catYYcs042M
NbH62DPlwIpIdFaYHU5bGqo1GQZICqyVQnGNRcqwJuphgAgwzyWdQ/F0TLIJ92O+
Ub81py+2RCNng6U1ZsmYOEf666oHuzlw3kRfjd6hU7jZjUQuPlhTVnSuCrwxVJzP
t6HvLasMXcJH/7kFK9JVXLrJyI+A0EI1qGGGEeESozmLIFcJFJ4NImcJE4AepdWB
U+5YB2dJCb7nTdB/q3/zZSBWpQc5/ECCA1Ldufybn1QZpnYorBDN9bs5fOGZ/tRC
Jia8mvH5WwQNZ6polbBDecvdLTAtwfIgdQbzGunVe5EoKlgvNSEcvV39flHqjU6d
opCe0kKuK4/T+IffyZvENAPoZ/WR427dYTlUhvNugNmySXRhiC6q7FQ1QpRkNUlA
63Z8qsC3M7ecgIl/P5l5DF49SLbXrWnc2schyWX/rTWuC14aNJuQZz9037iqbJqw
JxIW9VTO05dMJf4+Ha6YPnrnfm2RT65NM1Ggm91kKcdmgNW6t2+OroMlZwb6u+g1
U+YZErikQaZjRYpo1/eonCmFiL+j0FnUtgRvhI4IrTCuRlY4EhfmpgnfFUYAGnMB
2hOkKSojXIOArFyGih/azWcog7/uduTo5RFcmWcO+W5hH1INkslRjv5wfuVxyhFS
3K4M/kQ98P7aoJTGEs5lJGTsxUg9V6odXPTkvpKctoQPfB7zO7blZr5AOci3hrdv
+w7j0DqKBqqW0YZnTrOa1RLSsemnuEQ/57nVphXfq47iq3Yvo+ZArGVYECvbF5Ga
LsoQTrOE5EaG8bLAdpIDhuGx1qZrhKU5eK8AFo5Dw8RovgpBj4VmBeoZH8tM37+b
g4P9ycFvdYbgj6i9jo1iMCaaAT1s0uZd64eq+lrWLH2I8EMWn9I7ZPwPQRh5gxS5
qKGahzdHDCbmqt8yXMXez+sp+PkI/3+fhSS4tFM64CBnO6ADTLh6BMtnm50HM+VL
cNmrpj9KCd1XyT4Sge4kEJcmSZKjrhPA4iKeyZYiz0mFpSt89PSrOVoTwhCjovTR
78R7CLjmIBotT8Bk14dfBJMuP8l43r8tl/yZWACJu8t+Xdhvp4i6aIvgs0KDkrRE
NxjGHpUMtSwbksCVwwQVawmP/VHyPUDLVYU6OlhGhHHaJi+ruPxIQHbk+s+QnA5s
uCcpmFsgddLMT8YW4dFpwKFCqi99mnJ7wUxhDNOse1rba9LyLc3YUkcPZ4jc9NTh
QQJ4Qw+GalXV/sbfrDLitV/dXPd5ZB73a/2K2HeAVPqX9dwWlGQydmXn8xoKV/g+
zBYYp/xyXKbMeyfL2ckBVadnRJ1IZTCvOyf/IjAueLJzU/VuMabPNEwGapGmPC8I
NTJ7vkTVqOmgT/SU15FY/sIWXgBMxHdR284mCupstvRGVhy58o1XXqGOie1iqZkd
WlgA9OiqiLPG9gJZCX/ReF9uXwTx9jZSpfVU2v8Jh1hdg/tPTiXUuWoeiuEPPgL0
IIrMCwPxMWmbHyYk/IYYlPXw6Ryy9WgduPjDTjyiDRkEPrr6eIy1K31VqymfU6lR
z0QgTOx6DpO0EX2Vou1LN7Cv7dXu/SbdjidAa7CH8+56sDjBHqjIOo6HItCGHr5j
+IU4+F+kvLT+Ny1TQmvPRigo20mcD5ZHrDe/W1yWqF2OJ2dv/9ueofwbyo52vxmV
gejN4N9iKeiqnnkSoz9VzJ6Jwa+Be9+pzYXvyKmlIfWHoUHRli1/Icl8/efWn2G5
kOUgMHnSktwG5VqWP7/sF5EZGahED4nZJKedcMY8qWWq+/H6/26oJ5vujUaOQSl8
Epb0tQtEmLttyWkbpQ4O0x/oBG9jptR8Dr7wdXuzh6s3MXsoHdZ9J5wnxexpVlic
133u58oYwxpCSzn5a6MZjCUHoAWofwEvq17hXPlH43KnATJhjTuMWrVGTDQwjNMv
rHc+F4mwC0ewI+4uXtt6mtW+AfVb1MYVHnXu58nvmYQkYJ53Zk9mY/jhMjC1oqRJ
MCP3GUDN2pPXSrvJyefTl5++EBnY6BcKR88gJEGcGhK2Y5p0oMRz8VU3PlDK8Yhm
lEfj5dnfKLFyVB4dRR1NI+X2YQQCM/4ReI9I6tvgtHx0KgvTXfWn9Ad8esPrdzh8
Y5rtiRR59h6+iVnL6WrZv74izk51bqOcDH3hGm1XB5hMNo2So/4gXwqLI0HHIEe+
mtfX2/mY19NGVQOyKEdNMQuEjk3f6jm7znt8DiS3WgKQQH9DLyBjw5Jr0IWIJqzF
lYgZhM/EC0UgHlXUGm49YtRK+FwA8YHglq6avfsWnn4eWK28PxS/v9lYENxxkdGv
g6BNxfvuRLIWC5LOt8hHCyvQPfrNatPO7NwD8qlMtihta1256qoZt7B23nKh3F+K
p9ViwMkyj4C5I9g4seLGwtWPMRGglHa7FBNNEObrxxM95DM6s9G5r4fcQB6U3tmn
CI2A3PB5GzPUb5nRKFm4mjHM4T7TS9MChpFbm6P+wxUs3jnJCbHOkdyEJRvVGcox
Ks2c6yR3nJEm+tMCZM1ybajKhugOVY9bToUVaeD+lqxLv7MGkt7sKUggt0WQHoU+
+AZTl9rOaQx/xHO85RIJpM9SaQUiQdWJ10KOX13O7l7I6DWCQ6SFbkkiX2RkxECx
WaIurnS+PieJ8szeq3Nc5VFi0Ssr0aTvm8GBxHGp4G4h1GOmSGSQinrbfDjT6EeL
Gobjq9JwWA9Ub31iyBe+yH731Kt+qTrzl4IsK8Vwpt2ozcFDEJ6Y8noN67WtDuEC
moGJ1WypOnSufBEKlxRJWH732udZMSGGiVErFrUp1JKuL0IkwIzi7EXQBngbuJun
Vmq/OJcDBgeJjduUarrIZqeTHoTmDQpzvuicSlPUUApKS5ZrfLR45uXm+bFH92gM
t7C8IUUFj+62KwoiNaX5ab8p1YaTn5V+Nhyv0lXwsovMRtKy6WHR9JvuW3qIFol5
pBJZ/gMVr3PtTF/ua9/q6qc3EWJMMe+GCHWcwh2JjXp0FS2o8NPy4UEsD5Lvo5Uj
aR5xymMGeluctSt1Anj+Gdv6Z41HOq9SNZaooAhg7fjw2MhLgzwLcLQEMkLY6M8/
fYqrXlDw4zPvbzguTTy+MmQmYx8lf2VH+nr97oYwMsZaGMynb8KwmRHLFLB/O7GR
7LrDRugLJaqaFRR9HzFOGd1WvMH2XXUX4Ge9k6Rbcrj2hmHjw35XKWDp0BU5xPw+
PZC8Vh9CneSinstbyNjV+Q2UV60fOLEKUdydVCjE6l9C4+t4x1i0sjII0APGoHoZ
FM3TIaU7oMMebm/F4yJUuaY5pwXVtEQdXSZOarBfT1Mvvfc+Z0GqT7agdeACt1Av
PYPEOGGgRzDoZzmGEOvQ0vML+X99Ndup7Kx/b+VDzTEYs0eiIb/bzUTdLQh10ZzH
02S285TUgMVDtgSKrdSd5H/rI1/Dz5Dtuwa5citZljuoyhNPSG9RARcAGsObW9P6
eWqwH65dEYye2//ZjURCvhis771Dzem1ozYAVqI3WQbXiDzvb8j+8nvXGfpKP50Q
v73ysXlZMkiI9vWOqFOHK7f0Oj8mRxIrWe3XueWKiUe4yh54SDfIPbEb0UrjV2sM
a4mfmzkuo6NhZaj7UvEEo5WsUAxH+siYWLZTbDL+Gg+nZwQiqJaZmVNRkORNaLUS
+qg0TOJvJbewVuootlcF2KMp6Nah28CsXLTcoslz+qFuSp6SOhGhBp4ZrMfxmvyK
Mw0JZp4ejV6B8WiC4mv4IlrtB4LKr6AR40nykEx4qZDmZkLkaeKTnq/gmPQkS277
j9aLuBVDB5jxo/9azkz9vlfnPBhB8lqsyWAus4A3lMGqc4fNUG77er0GVdtDrdjO
xjXv81rTkhWrrCxQDNXs0Z2uwmFvc7PatPgaDGVlw0qmRT7yMhG2PHvJcGIQ5XWO
ff2bOwCoFBfwORj3mEwLnSAdWYdQm4eVrNey15aAomfdReHZhOtFc1zM3VGC67RA
ZNn9Q0ZRV2yEF7KRYdTuymYdhXrb2EMLVBDOA/IKmHBtrvKoHzvUZ09te96hkNHh
mNbRKRepv3Tvz1bjWbUehja+7zw48PcVXh3jzilw3IqMVozqdtz+goSxQYYwsbCe
+XKrfh6UDBqkALcGQmidndjpMpigB+X0E4bUidAHpVyF4SxIGaAleUJnyVnjjxO5
oI0wvNbuPt/NPvbMZTqhP+WDP/ym7ubG+crkh5LqzNvjNRFmaDaod9lA10tYnLuA
AZ6TdOFtkWZHwifP9VMV3+6QuGDf+u7B32dvX1q3pfpjhYGnqa7ldvibdSIG8Dc4
cwTJWasCZLweLjgoMMMGjGQoWN9Pz5bkvUk97YG1wRCpFu+zibLZS0BdKANzmgjE
2OETob7sDfCjZQ2+C1eZvSNzdwo5rOyzbcjTML33ERR6qUt5cNs4OjZ8LuBitJ7B
6XJsUL9c0Dbs0jvqAvsAa28tc/EO5OXrUc6eMDZ/ctqaedGUUAlUTyO9TVG2LCs1
FIHVcV9SHlKKJNOsEOnRuBpShYXfhFzygE/CmeLo6542cLWW8GBt2GnMJ3aP0T84
lm4reHM7NS83KSpdxI56Cn1ZHDjiWywALl8J4EAHJ2zNYnKK1w/ZL14vCgTWtG/y
ZNrGg3fMuGcHzV197EvSwb5xXgo8PixST18dowUfZWlIMTdKkjF0wk2RUGMUStZF
eEKlPiUl+BbTWD+RBGluEp7xzZ7Im8gYSo2+00qiot0g2gZr0m0teuB3EuP+Pkfp
yrfZxDkWns2h+J1iBc36VfL3nEmbPgNbKop3eco6CjFvnUo61uMaKyQ01HIvN6NM
yRtBrMhl39pz+SeZS8Ucklrw+cPI+XjG814tdeGEZ6jKbXiFTM9xPr5QhqrWwv17
qoe+KCSfmbA7xB6MUp+UDQoJRnLYe83gLORT6LOEotQ9ZvIsf6hKnLB948BkUNkS
lBUCwEZzqe1zDnwqQ6K0FdqB0FKd96ns4pwQOnZVefuNuV0eLJgRNQ/aJFV+gtZL
SqicBP/0mVpRSRAai/xAD5fO9Qdwj7Tpk6FgI+1zFj02Hwj7AiKcegZ1ddHNKgb7
Guzu6gtILW5FU/9CttS1JYrcUhFY0gC5iMvq4zegzmrV8zIDlHaWyoV3JDd+OEVY
KFwjt0P4tb8aWzmnpAjpAEZHDJ7XXovxZsThOASdyA4D1G+U28OAGH2RDQak7v2d
joCXZkacTptT78RI+VrYC0CFkoc0EUJ6/Oa1HOxnYdqyEcV3p4NIxGmx6RF9AQ2S
bOq6ss23Jfjg9cmx7rM2e6U4YzIBNJuw8JPwevMQIQ01rl06sWuP9Xes9+jNC5Ri
0gMNHgfqTxGcli7P/QQDAtrD0paG6ZuNzi+0ESHbK7kSQvOrsD3A0Ai6W4MZIQce
6QBUnKSjDvKHDiV6jcDPGUAyVsbvMR9uCTYYex2X4a3qVg9bER1FsSJdWL08qpel
yIsWY0T2jmhkFQoooSTzjknqRGbYiNOa+X4LAiEn7BcRPek7tGP2DAhQdAoEy6Lt
Bo3BspRzIOHJ31MD0xUsgRvECFJSmhLbIKetNH3kzcmiAbNy382quLtMYgk5Z719
+pp75jE4Hs4eI0gkVf9wPcR6oZs5IVmv5MTjRo61Ochz+bjETkpq5Zp1oBiylwTW
rs7+X+W6SLlGcn2+/3ZJ8q4H2jo0wxRICwqbuadQ/Z8kCmtYJJOMWm71GEgMiaiI
1CvvLPB2QljUk/q70nOi1CrYRJy/p7ZB5FOpacpSOEzmZR/EM5RrLfZwYjwf7Cfj
vLCq7TL/Et1XuKCts+wRDRSGvjZ4qNgzELrT3ruwITdUs3VbX0BgYE2Kwl4TXlEB
WkEJJpdOF+QxX2br4CDMwPkCVj+PAnstQIDvYQsb5k4Sj+S3/fPJRPdDO3zwAk5J
/4ItCDriiD/EuPNjXa8W2bKq6Yjfb60IOwss1b+TbiJo+zdKuC5LjZRpnFAvhZLS
l92S8NHSKk/vMwdDZiDcVvxZ8Zs9fk1Z4hz9y2FZrb9a6kD/GKjiMiWRUa0EnRU8
PpPzws26g4jUN9pByW5+UMm/R4DAA36F2A9rpooz8VOrp7kV8YV9AQsq1QFgfEZa
/2cXdSCEkPBDvDs8IB6ONmJ7x2HDrKgZIAAwdcmkBaPq3es/gTThqNAzObMfUobQ
ayTS56g/2/47wdKpheJYLsABU1VxMP54rRZOXSuMd+83xOa2P7gCoxvGRjzXFIqh
QNav6S5Ws+SWY/UObRaAcl3oPfyfxCzEAmOF3PmGRB1XLmfOS/r/92vRjaqaxWIC
CXm/yKrMqOFyDYvh2xeauSPLERsNfEpUxfVETGEJaOCxoAwcpFFXfyY42cTJHf3f
f5AIHRMvPt8JymmGCA6RKx/jzSoK0JM/D0PNAf5c+Jy2NhC3L7eL2rUmO9hrW28o
xP/xVHfemjDDuWbsTs5okjNbUNlUtp5qzXttYYzkLietVHAjLPiYOp33aMyG3+Gn
N3ZSuMI5pSCAv7zCrO3/7XttnSGk7QjrGKdI6Gsb6J05LF20G48wkDGogq4dvDDs
s0UlkkZsHI9bgK+6VoyYyn/Vhy7l5TKXXpBeuu8r0Y/RWvEPLpHINyiXKRFcN+Km
XrckiAhbtOgRFI3gnw1zUroqx5D4rECqqNe/wPuil2UdgbjN2spU9ArFg+DUCgXg
aOlu6J8gTrtX0GsIaKHLWnyR4Uza5AJtamH09wSCgxSh5DbjB/RsY2Z/hEvjk0A/
7sKeJBd1BWfVr0EkqIXd1Ed2WvpK7DlBmM4fkqimzvX5BlB3gbXx0EGWUwoo8zv3
XHvqmUVHYwyO1gsVQE4o4RMTqrBgr6ZLQ7LbuWxPzui72aexJEmHaxHEciySL7MF
kiwiVOGa5R2Ks8qzZmDgUO9ZgRQVIyYVgy1BCCCPcdGJYDjcqFpENDMgflrIIPx7
bXabskQEsCWII+ffpGd0a7xsgKta+rKpisqkBGhE+I6tGq+ZTA5WkLAvQi6tdVny
HbMlW08v9aQqZOkxiPkFLB2Hx5z5PfvzJkP3fTM+YpvhHkQ0tUAh+CBDj5lj8sIQ
iZzzOWa2v+GVKSWGdKy/+rL6f5A+iMi/0jc2WhNTocv0sODFNxhsR2VQBsrCG3JB
E8LNOFCVPSeRTbS8Yu7r4lsEsj0fxnwZqHZu+mbdyji0+BX2kRmK075EY4bWZIw5
5dzFKHWGY52+7wypZYr/D/40PUvZzpABo6faJhGBJ76C3maVK93nfLAWtmi2kHGA
gj7T1c99oSVrovj/rWUFTm9DDmLB0RgMWPvSuQb2HbcrV3Rk5De0CWVGp9eEzpRO
Fh4kGKYjj9aEeH441ZuAbZU0jKZCiiG11xdhvRHBvRPPSgAgHgY3MlngPYrZsOFj
6YxqpEOuYCht6FgmZAFykWPIMn0eKPVajhJB71BmIzRUVrI9mrxXQvR8FFhO5c3V
8bI3hDoffXz8FVcDzM2zByq6oZGmKf2PojtOlzEwWKsXMfDANRBIjPivmeh34QkZ
arTgFZQO4lYUgBSo+gOHdquYnbfD/Q0UuhtHlcuSlbKNdfFfDW9Njh7v2KAY6Ug5
HLwbaQuSbNUk7sxfFpvk1/3bHZ35OG2SapcEpmBdapSNzHi4cIinfO61EhcMmDMW
zubi+bGARc5f7S7DG9qNYBwy1mgMc0JZsIPmbsS6UwAUMsfTD8yCYeb5TYIJGthy
zaAgejsr59YLI7E2WjXwV/b3mUY62Q8LiB3rT8hQkLMg0JBGA9slA24ZKEaUOqqa
uUkp/BeJLHFIiSADtHHMwKmRVJrvGh1+60oOoWicuQCop1ToXwE0YPDJ8GsPPGYX
ePo1/hU6NYE7ECH+DyWaNeY3NjOpKvs5ORHSX5g0L+cYwsqc8LjRaNCnIkm5134i
+xPlU5hYqIg0ZIvo7rwPbJF44QyuG8Wd/hWWsQH7muhMX2VYsN5GxCLx9gUOPULa
tI7TUcSiNxM3GnUELBzjM/K8nHXO0YeCi4NHTtEA8/ydeuUW6ZBvPDRyOON7h4jV
K0ywFTSRvmFTwC6NKAd4LgeDJd7YyLf5vnmJiUOy0yBpK1Rm/gBLoxlstpIiOJpr
o1MxmMdvnOe9mcoyqfvIANWl7iQk1YhOfFw4Vj/RO/5mpnrVOQEpJ6KQnW2hJzGe
njX+JVZzv6qPGSRfJ8gklGZBv+NNXqCvp8mWZj/XXXlSfFHc9sEcuW7Lzv6qjoWy
Y2R4cfE/gSkDpzjXO4UlB3DmgMVzqzW99v6FsWnthjO2oO7up3hunxWc2Dll9xvC
JJC4waxFLhKbu63zzcRXPLOLt/dk3VNzyKvET0dabgOYmzq7PyYD2NNLHChAoXrL
lvl+BKmZeJ2ZeXFGdPcBdxHeudFrRznFjZi5A4wcAUJycPEgnz8GinuXIU/CRxzR
m6jE0Mx0LF4umKndPNLVTfXYvRQTm8Xce3kIWq4lrL1ymX7T2wdxssxCh75vYRJ7
ukF7eRwspCK0kpuQ1M5o1ii6WoKVrpv7pod/cP2R65U5DvpDuk9tqRQpwrQodZBb
RpsNDmZzDeM++dQYjqW503Msyg8u18KpY0qS84KzM9HlXxmYfwf6yVhp8MWf1qsW
oHHZifbvRO0mRdPLd1bn0LzX0wyP7sGZT96MHl4l9Ewh9Bu6frDATcdnFEgn/cnZ
h1Cr93iz0m0A5hlRCeEe8zPJmgT+7cB6QmDJeLX5DiYnrmQuGCeaCsx1rMkRhHYG
xVteIC+iThbX45r7PaHO3srT2AvJKD+ar51RukvI8sO3Do9ivtSzmyP1naNOarPU
hsPNumVEK1u0E9iJ4EyTrPa8GYRzbvwoNB1ApReossklOGbIQgPhjMwEBULzLuzo
pvvzi5/kTfyZ2RtTNGf9c7H4QIeGPRsZR6hBUp+WPfBfv4d3bCgSZ+OK4wyP4TCJ
Jb+NP4XjdVMDlCYFdrctf8fXCiuyEN7OpElPcZRdZu2wiAigmeu6MVKHhS74vAcT
F9+t1pfs48LNY5KcCM6QTpF5r+zI2FfzYKzR09Rf0CVQZ+IxnwDUjBfj3tuYNNNC
z/LOmdRfEpaheQ51oSQ8mB2Xvc6zBYxVcTRjDqD+FQKl0QdXMEXenZt1DL2fhk9F
Oia2Wnj2XCUv1hn3ZjfWn+2bYAc7/YYAzgUxXDtdYYTfrfflTPwQtLNcoUvGCSYq
xbDQc9U2V3HJ1GpRL5cEGYdwieBYHQ9zNQcUvYZLwjRVeYP07aHiq61PFjDmdpOA
5OBcjb97bMcYCWo4rL5qY4uvf3zqft9n3CzXaqS0pgMM16tGBVIQ1WAeP/Xv+un3
tfDau2YdwjW8NrLgeRJF/SySXgatbPoNU2d+MqIftKoOWSuXqFLYVyxtpGCYa5z+
wp3c1Ml62tHLPoOp+Qwbkx6LZOQiYrWNk3XoJuvPVPmeL+p3+S6tw3PRpReuz3Hs
RU9I/YBzltfSqGtI+BmApSIfzi2uhaIQpi5gZ7H2FYXMUcfUeU8mUXtZNWLDDaVE
eSiRd47ooYKfEOthgFWeAPIopHlfqUZteEZp9L+4IFAF/Vo2fn1gQoKgsxrx5ek9
37dSUmoEdKFuKvVBleNUi0mcKdt2V2v7/ZjxI/EYv3pGdAPBZNZeMdkc8eUcmA0f
2A44sj11sOYI525UaJAp4t9AE8vsk5S3hLV/3mjjkvxSzN9qMhTxu1B4c6QUxKQs
k1VPkmZKlCBAbwCkiPZetF5bqOIfityT7FPaIEIXTTUU+a9Uof5Tdh4gK+teHFZs
5f1kR+TmdNKmZjvdMq7FVOGGqS2IzPh7z9VdxDYsnNmQgFXOBexrffzDV6oBmuKo
c1o10K8WinS6WDi4QycQuriWlGKDCY5Vw4PnZCHZnw8QmLziXL9RgXn6T4JycBaQ
6xljG5swhd/C8jD/IowZ+JOxUjwVbU3fD16VXk2CtaWi/ihhmX6R4OtrzfBo+Set
+HUAs0OVNghaq33UwGxq2eicnTTYIw/y0MECe0TPn4Kg47Y2LV9//5ZGrVpSUu81
Lt7CUOFYWRk/KpI+SS36C0oT2F3VlG2/lL7HD9ddJc4+qvKSSK21MIoteJdz4b/D
0aJbN+irUgjK+YYK8GO+Au+kQkx3MNkMM8N3sKAW+Ijp/RXQRnFsm0LsQbjUxLY6
7sTlEQzFi9KPIbRqinmaKeFDlBTnpmAMvHP4AJmYpQA5jIvpLkaHL6I5CXJZBfz/
WMu6ohm1qPLI4rQflw8eylK7CSeSVI9yM4C78/5i9Nfh2aTIqzxKFBl6F/kfLVEo
vT/zMUBZ8xrl1niPFPC/0xHs9l29rq0mkW1x31Y90bWFkgPBqYriMWySHOmlMc0A
TeQENbfAQZ/eit2HBu2zsgewjvdIhwoHhP2uxcOY2KzH+VOstuBjE81IRRuoByhh
YbQ1uJAdriU2g59HZEKTvnnPpkXuchvoamwYZBUJaYcrTRjEeHjdRbnzC/M0Qgo3
1ayzeDDQvw4glB2IZO64nLapd5l2XI6ZmBDqsZIPFBoJD6pQLliWxRREtuQLKw4c
UF5ghoKPYlhFIHXAM/o2qELz4+UNxLw+IQOR8ELA7rVjJMcPWZe0rS+raI7viJWN
Ld+A2MuDUO/FhS0PW9NNfrF5n23TGq0lUJHBXqwvIxwXabsymDr4rhX7XZDYVlrv
c32tnNwGTwiyUemVCbGOrQEmeKnL+1qxCKVtAywlnACaPFaBgog0RAs1fhCxoBgB
oXd3WgLbJPDYHiVNlq7KwjbUQv4dGEBVd3jOfxtfWZ6HD5T1awB4Sty+prF74Pjz
3537I5x7TANLcz+tfCDNy9hCFh+eP4c08RivggbQaABFebZkegtOyBpuSn2iTrVp
quohe4u7gouqgTV7ycSz8sz2I1EpdCETeEynTSmaCDgPqE4wEFof86/k74GxojRE
FruM4F5fuVCrVJftaM4VQVYB9UHODMIjKlE9pzAnOXVCoNx2U0vB2rktTgEfx+GS
keyLrGEi7s4QO0MQBSRWlyfeMoUOUa04aMiLRmFkredxGzbhJ/5WZ1buz6CnKVIi
FQpIz1s7vDLgjgRLFVdhIQWwK7wr4AhTAUT9tRSpRshRCxZm5eDQRi3sAYYUGwD5
aLaXPu5w68sCnbP98ztoi6QQH/pEaV3mh4tHIZslod0HL2Z/zePGnka1n8c2Zd7F
GD+s7vv7ZHJPlNZmaN6oLV8D/wg64KAiD1NP9pSgB0Qy9f3OKOfKVtHo/uMVZwDo
SEqE0w/KtCNYlwz7tunQNXIZSRbn4zDZ8Mp92Aek3xvjxzKJIy0RsW7EO/HcdtPM
LftrbTbRt64/8LpNxd0g8eB+rPOugnxiy7y5JAv9K8GxFk3NNmZoTxMmdXAR/jXh
SK0TkgGTNAgE5Azay5A2XLV+TJUAT7lhZmltVWN+U3ZoDO5V9tkgzmDCWC2op3Wb
xKeKoWjCpU1me8TGOWoEeLQw0fMWZFLns2xAGEPAr+hDMxWcuKvuiM7t41ACXSq5
lf9ujrt/22XSi63UI+obVHOAdiKMrQQdnw1kNvE+xbsqIp4U44F5S5NPh0EMpe/+
wO3BQ0NpK8bYLvLZTgl2ClbOuO3lyvRHOv+XbfmBB/PZTLoXc1i2kIe9iD9MLaMW
bJPRnZ8JTeWocYzk+0gw2oiuGHptR3Y8WnIX5O8oxousLAP0AaTK9fWgta5OrLv/
rQU2KSZXhfCoYLRRK7xuAXVo1DQH7gkB9GFr+BrjwQm80s/etpSx3k71M3YYt8hf
5BhhHnxfThrcZedfoELqKY2x52oTR5uiRFOH7Mc9DpGvjiFWcnOnV7Q4uK7EaOfw
zrpCUgU3Q3q0uR1zks/VZB4QsSTTI0sWqyLt1107TYdBlQ5iyt0K5pUzxd2bBK5y
Dtb0ryRHZZF4n7o5sw//Nf3rB9ZU83cC6EO/2yvJIbjLJAP8XxsdP7p7Ya5IMihR
YeXItp4/JL1e4J3XCt46khT3MRoFI5wQxJc2ZHJfVQgrDvHzdXO4aVRK3sbQuxQv
VzZMxQnhs5r2G6UJTHnT8Vt3rr7laZlerngDWAif1q2pmPIZnZayCMbaz3Dnl5Ac
kQMqCs3H5DjhHcSbKsH2WjSJPt5i3hW9GjFen20ZY4Sh8a9+fc4jTejyhhiHg+sE
GBodrUDRN/HbTOeyaF0D3ohEGvlAnQjoI7mMNNc08dG+QqIzHY4g64ZVKhppC5ue
1BXEkDhCnm3rj3zibnDo0jXhLA7SUhdD2GdW2qSPnW0f9oHb7XOAkHGPMybya+HF
cqeweJs5EvMRR2c3vKwlUimjOnb/qpa4YGm/1Rzho5gI84j8WA2ZKd/zrMmN9aGt
nY7t5u3AgF+4aB12+ZTsa7ZqwYEOTC9NCsc2BcSKF7jB8WRiK/bNCpqRJ+3ghbpi
46Oc2ZJsRvVMTcdQoT6AAWUNYdqLzaYhOrKnd/LBstuoulMWS5NkJozc+DZ2wt99
mp9b6j0cbZNwRekanClNnZg7v1hOimuSXIb7LMMo3zZEQE+zw0ffnVF0Yx1LWc+T
3QvBRQrQiKayl1j25QxF5vozXqDFHse3cyimp7fFImkZeIdlD5yQe9cWscASkaAP
wvrDKI0FfL+u0moxit21YGi2iLceyyk9VLecn2mDMUTT/bUjzgqmnTrcUoX+kynw
vUYJyl1x0KtLqwgw61tdQSc6cvLubkz5GWJgpup3F3XeFKSNmGwPK8JdjrNw64Hd
z6J+pCclxP5qdlSfR6sy8XEOrbzks83zqSEXW2ppPiye5uYB+IK/ZBz2SL23MwSM
ao5hLk4cnda7NsNlPqlB+/8AhsotbPbmk8uWIbPlK3f8NbS3FS9Vcze4MsqRLB38
FRrvOImg7Absnz88joOVls3sJlTEuFasUKY4c2PPJ7t2OPIhOt4FSyfuPjYRRmTs
KTFCAhK4NBLP9aEuytRi6BX2P02dn5bMX3/HRG/5JZBi5NHQVCT5xHxHMjc/glZh
mDb0zOmA0rxkqJHduiz6J5J2j5iX5/E5VV3++IQlm0rDtvLO68qfBSwgyKTBWshX
+BNB2UW+dJS42vnPZgCu5WFDBUz3Fb1D/2K7DkW5PJHKoVmPMEhPG4Rb4/m6PVKL
yvfFvHJ3iGP5gEUlhRIBmfLG9HfHVgs9ORwZqtvJ16wOpb+5whn3ecz53YZMKJdw
/NP1s/Zl8bZXzQDi5U5Sc9ZEJ8dpB/xNHT9rTuIWSm/MHn95nrgzoL+qwFweOVxB
PlBnvzheGUQOuxXRqlLJowCtDC8DWw1FJR5H4i2sdFseAofQhUqn49p3g1O7Uo5R
t5STvf4fPbZb7XHygDSVnr8+ltctiO03zx3PCjDhjpLx+fe67TjgifFt6Jwlh/wO
AWPm4IY31KOfMmuU4IEtRuxWFxzK0NvwpzOLXhzigsg4o5oyvDygeOjtwcOKQhYJ
uPuX0anLqu04ltxwshl3pMyCZC6fiayjppohNfzWUpG559yHVNUvQuHFlAeEfVqr
Qmm0798OWlyJudO8+qTxgGap+xOGiFBcmqAalazHbC1EXhWUF1QoEHtqTqFBbGU+
a/IdGBX2+Yl8Jx5di15s7cpb9x6hVrFtXBqZEZuxXb1RKan7tpasWaG+rvwxvLHe
vmuctAVxjJ/3qkFVe08sdBJj8wQlDMcicZGnHmI/aXyHWG12WSxrjZbY010wKaDs
IsF2hG980JXijWwFMsqa7m8ciL1kpepmt44/7XQ2tk0ghF+VjyD0ehQS/e0TJacx
4D+XMKHUJJUzbTM98LDUO7Z9YHV8i5GehuW+qA3A9NsTxOPvsZdRzNZcCVrGSA+9
Pka8yXEweFLOzGENbTw6wJzj7isKoUmQ1jVmeWm26z++q8t6HCQlXUamOozSNeoD
NpEv0cUdH76j+/QCGg6x73PT+L3DfLqxulx8rA3AYA+mzZNgCvOqI+aHDJD6OcUa
rYcWHGeFFST2nXd8xMFJA7r80xvWCsDajdg2Penf6gga4FXaIS1zRkRgoiEpVBtG
nJ9M4YzoYomlrMnRvhgWLw4M/m7QLXAdNdLEs9pmNe3FM4sm5NKjuVoPggMayR1C
pewRAEL3GRBltx9KN2XRlWj974dpYFXvEaQ7laFaaop2zHlAyIYgJmR4Jr7Y6kb8
0lWDVVMLcOQvZUpZzCcKma9xXc9kv7dcGC2d2ms3686LajJ8HRWDKdqcgfhzSaEw
c6Cq+4E2QeE+IZdYGEvEWTjtsIf1WlaorugydYMomJ4OqXIwJ/i7iwkk2OLNiK3A
zsrkMQFxstFlKV6pYd6GXzhCMKoYBR9b/WnsdYLK5aF0fO6kZVidtr1MGvWpLFG0
7cU9QaqcOM82mNqi5+WXY1WYQGxkg+mw4ffWQuagn+L1wdOheSt0fXrdc3zFWmST
sjorrkiLOY1FT4gytmqFGOMFk6EL2HgpgLdvkMSRu1IUEktot1n0yHyFr0b9IiaH
zoxclqS8eIKIvhgwe+94zU9Ar3g3dVQoOdSI66Eh2Mbipf7C6ri6EUg3SZ3+UBnr
DdQhBsv7erNKr/jFw/rkWwn5L06Y99pOp1KhlXROiGiO7k1z21TqUMZYEUmHEP5c
MIAJMr6cCbTogePxrhG3u8FVy+jUf5Wn+Cfu8n3pbHJmgFGajsQhgjBzjDpHYi4X
RMkhOS7ak7KxgeEZ3ML4jkaXfj4ssY2gJH3YWUIaGzbZs4kfm0uIM5sa9g8WZk8H
FzVbnXKN+clxgm60XHHBSDnon+z3asDvD4zs3jDa1+B05K/oNabFWNSBOBPyqIf4
k0+EDjsVMW0WlSNESsI0XvV/TwecuUodzLF4AoCCjNbncTpAcpYY6rHjP3ps5aq4
vMfWiFmXYL/pDH4HhuIyCwGcWoTtlWHtN7kLmN+CW/xAZt8/YUrNfWAwdEDCULE9
aUr904noQ+0bUH8GIv6RkAyhXE+beMwXPHbwTisqTfF8p8k8oughOOUP3+TakJ14
G1/OF4h+H6Bsfx7xQMeGeP2nMYnOxLuAloRzYt0BTcNgwE8ao/g4zdtCZ4KQogLr
Xpu+LYGIQ3vbTj0WL3dg3jFcASZenyoNFPzoz4jnLLEYHF+Da1cr44E6RaWu5vXo
4yfNmuw2lV92p98NVPo9OBNVWnl8KjU9w7Y0yTI8nQKTdyXIDbAPExWnAMYcKXsp
r8cWPP57xCeyGtsuDoez3dyCgyMBK873jbsAPtIoVIRAGSxd9SuF/9ifBDETyyjP
eRqUVQPzN5B82ufsNQyHVV66ZII+DAgWoWy/ME80Ijuj1GKomKGtl6wPFhUREZat
FN4ip6l9W3NmDxQCWFIfS2rK61hpheZudV91kRpZPgjWAfWCVpyk8N3OZQNvn2m3
Ysrc6T6PhUCVTrp8E0zE/qX3NIxHnB+pBXCARHZw2pBqprYG8FzOQ2PLn4s4dCut
gDWk34W/uE76Sz6mh7WRyyoW6nZEidVnR304rvhGXH7G8pXD1geNLTbmVeS2Rjjg
DwOQogcIrcSERGwpRAABHnbrkmbNCD5tFGELHde+3KnJWXE+8IEhFVgprk6ItO/+
4zXLxqDK70DmYVrQoEgYeRNIymgyZV6W6A+eKcl7Hb1wlw39wBjCT9Ct3cFuFnQW
BlABByivVvW5/WVslAHwgDl8jJJ2xgHA5s435hgJ/f1lYnfQdb1dqqkUo/nu1pcA
LkM70CZaIemmn6aDFPh+2ZNC46lrZYYoOSp+cf+tPkLZQzGLjuiisbv+sgUsZDr9
PC2sSRhtnDVP0D4HSepmcbPjKaGdvMu2gCi5YDEdHQfTLuCTpKfqSYtXiWhSy8Gz
bITKgZcwUwtWepnqY+KJVDXEWMk4n3EkY1kQi4G1ISpQesJlJ9nQRr0TCrDwPSZ8
zjimft8Y4TQNSr5LbodtQI58eN0yiC9SMEccZ2I2r/lZv9nydnnF1XqQW/bpfZdA
XtvovsbNRph81Q3/oJYa7e0D75v5R/6zk8dqzlKU//JRW5o9kSaMynkVZozKBA3i
cyqkQe8HTZ3f9GFEtJvYmt5LSoOrWmcfJWsR7/XoVuZExo1BjfPmsRsSO3Cmv0F6
g/vauVdyV9uT2mC8Hd3lWUKzKQJ6rr5SIp1rqs++10R2+WcRj89D5tlmL78gHpBT
B0cNfh20klON5GEshC6jYP+lGuci4++QL/+GRmgQb//D4d3mFvwMSuHKF9sCy/cY
5siOT9tNm99BeNZpiZDVT1U4cYZLq3eeg5XcWqQa1eqaeC5obPm5SPbnToazvq1S
EmWNAkWe1NBTRM+s/2zjBoH5G197u4KeLvPEhs0TUqT6zgoSwRDN+VCzPgvPriSE
YbYO9EtFaa9LZ5g8PffXOt+/V8Q2o0m+tptxFQVHAtpdINALb3II5kphQO6NYF5X
rWr6OLxk5AAVIDvidNBtGqO/3JuelKgZDMqn5oV1zkp09HtQ5gD0YOn1DGqaVN1J
vvQG5LqYS6FHK4JGRkR5Eyg6oHfNhk0Z19v5W+JtTweA0xAlTWnCUPhr+eNerqN1
ay8UZd5Y6fPrsn3Kzbqg8AFYsuH6nOtRQk5HQNILlpEcaRrsHyywkQyjiT2AfUfI
nUjuzFsTBZ7CDt7e6I52xn/gri0LOnFc32tt14SnlEGsZvIAda5kObRv41brcO39
ZOrCP1XxVPoQ8SmOj1h9gHiWaru8tN5uOU5EnQVev1mM3DvIozl83OUMSzzFuxpB
YJ3ga3fRdzRRKznt4kKhUjMcqKis9zGCrfgKa1PSNGDzVQ35eB5KNElVKfO7wJAQ
naY2OFEbBjcMa6I9K7u2UtjlILYRcZC7QVohzBTbWM3rUSitgkDeubO6/Qw1kHSJ
Dl7gKegeHcZjFSAV7svLY/brlmV/7VLHjeWWeOO4Hj8Z3pM8ZK/cK3RTZGrwFdoK
XgwrTMUTGddSWnTAjQ6Qzoyx6bnphASZU6nFJY9QKqMsZUucxSE5bvSqe/N5h/Bv
PfsK4FpxtErw6N29zSoU7yKZxwAZTcSxVmxFhtisZoz7NWBlyXBTeyiAU3s1clM+
vL++ALVG2OVmPe3QYhb5Z534qf/kIrt/L/nvGk7/44//NVTCk+yza04zyoB78LSZ
7ypFIu7O9lvLSQ+VjlFwYg0DIBiaCGMPDDo+S5OJy3OjcBYTlT4CpHNtu1mCEK0M
UzaJFUxoWy/CsMcjGuUcqb3/Hm8lWR2r/gckRhD29UTlRLGwYISYHn39JcYHroG7
56RX/zgxzbiMJwE7DNRgGT4i+NYVQgNTzGDZOhuUkZaTKFY07KIzs6X/oqcQ4Ggk
gWp6MkiY++1QfmMPqC62fE6z1tkLhHvYB/4igNiOYjokZvGyWH87QNp2EAjN5e2K
KjJpcnO7k7WkSLFE17/bJSGLuUR6ZLJjc3nnNQYjqCYf1VOt2ieSy7CEDe0Cwvxk
o/VZP1wdNv/Ifa8jIwV7q71eR3xwWsTPVwuo/qtgpJQTBnAqYABE2I+XUayvEE9T
BPtc2IZ6WvQgm50avTp3dGvkC5Z33QILg1SayhcsHVE4RowUSNlLGyRa9s9KtWvU
7lMd1dii+D7gRroYzItu5ydyPcax590vrHzdp4yvOmGCM3096HE8BPB5n5SBeqSe
Rxl5jHLNOb7Xs4r6UZrFPIEJ33mWklJ9T0qoqzCddZxxcBMPWf+wIlWM61XK+G+g
U7aO33nt5M2waSSgo++i3YBqnedOhFii3U4mH7094Tkr109dP7d4KevzwVQlwyU8
8Bqd+GE46tAkjUId/NzAHfghT9pZKu6Kut0g+SBoA3dy/CmGTWtGN/CTBbb3Fppx
lpJ8NNSZaxaAXo1L63U62rK40J7yrUP3MjU/xlg2N9q3vfTj2fHk4Ckv74xC4ut/
HG5bEevXwgLOblvIsz7F9/jkNhGu9fnVsq0UktJSmrlBcRu0pCimptuiHeGerJz2
16JpgjAT/oQobkv7T6K8WgLCgy3JPnoMf7oF8FwJ61bno5kaAoIpqCVoZZCNykyo
014mIUPnL/nygRX3CLHLmfhCt3Awka17WuCKlBJ1OxmUVvvjY7fBGAy1C0ovHnkQ
jimFtgvMfDQOIl0/Xa0t4zdaoIOVS09RWIOkGuaAWQu6rHrjKT+A0twTAJBvlFyG
ZtcXIRwZLC0YQZeNqfH1EEUo/KOs8o5gUgM8c4KtSruwFvUnSfoD+COQFsJ3t7L6
DTu52h2S1+qCUeD1OX+XXig1H3jzfeX3j+PYFXjCXjb77c4Cn1SbIJM814wTHuY7
f0nKt9SmfwmYJFPY6IQZNgyIRhQceaiw34zeJ0fIKzBce9k4rNcTYmaak5nZYtUi
uCYTeuryDFcxcegvpKQDONhySEGqHqVDbW4JztIS3nFEbk0KBcLii2ZHqpTvnb24
eOP1VfwbO1YtWgxLtLgWb/ThJl62//K14xm1tr4H9oD6BeL7pfdz4veFVkax6hey
PWQhPscE9IVbVc94gL1rq/n34cNsET7gV7ez4ctvQ1dqabYCZklu/Oa4Z+0ydK5D
OgynujmQ20wUstf/Xlnfo4HTnPdfLw31ETXkwH6NP3s1X7eLTuCg4M+Gs/vNJHRL
2pEyLOSN0FmtkkUX9wVgXp2S+uXvjscmhOHCSFKFMDKB3VY0YA8YsWtiSlcbTvoR
ARkHqpXqX31F5Aj+/OTq0Y2zjbRqEJGttr+OR5xTPPPwR2Mx4xkBoyRjwC6XfeBC
YzKCwTqymRT5G+x8v9DJwrxkm7Hi/3zpJmaOMxUm2r0BIqm6Dchz8lcKTS1Gz5DC
E1loktsqgNMqJ3Yec1KSKFEDD3eFFcVk2QRn7oJ/t1WHzUV/IFilDljLRsAFrddO
CB7tCRsG/lOr0EI88+Bg26bn6Y4JlG6h60noAiGGcIYYJSQFGHN2J0+7dWSauiDw
XYCUKmMy+v9yAljMTHNUqScXYo3fXrMdAZVS4727YRSKmMboHDwzgXkLvdaiYe4/
b934BfAYulDv1vfC4FKXqb8HpB/x7bdx5CoXMuO3lqGP2nyY/q0UZVVQRwKqVBej
2A8LKyFuyEEvBxS9hkzzzDp0B5tu6CgkD6PGd0AGcL49bpxD97Bik7z3vzZ+fvSR
0EyPOFJtHPKONFCAWQs+AxOMhk6dDQ/DhpJRZ5b8CXFrrd1so33B4sYvL88CofdV
neIDm76bpYGC9PA/mbfIWI4izJ7W3EZcpWvBzVH8B4DCY8M/8gL1q6XVrUsPVjRV
XAq8BZ24sOVN11CW2xHgG/wxyOEpM5rDWaD2EfjJ8c6ovJh4W2vuh0CyTeytlnDd
cq2NOqSa3EKK2cY2cWwT50fm2md4LRVwY8wBWzkjoe4lRF5FiAmRh7RUSfTXbfFz
pSvB8UQFMAiKZ7198uTksr8hljolKC7Vkp/vLXsoFqoU+eqQUIBN5rLPXK/4FSr9
WqOu0wsCmpXZiqtvsIjaCvGY3Cx3CGoNqkQ4JNbzjVtee6mmivObe0rOfk0nHxjW
DhwguTRwjhajYlI8CGR3rjgIIO6hoMWN/gEYSdOtx52n0ihxA3nWAGKmzFuhgiF3
6J4VlPcrevJofPBRqsLCKAJf6Oa7fCREHHHYp8pshM2UZVWrmKOAQ0o2ey1t1Opg
QAH1EaOsrsm44VEnC1aSjbrkA95Rt9rWGTxAEbLYPCefzRKLqxWKrd0br2Ic/7N2
upruYDcN2QGBeLdEftWiwXGd23ZcUSYb8BY3T5kSvQLuIkBW6Uc46Pv/PT9qbG6y
rF0lqL3sVyygy8OUL/kSpX5pmyVXifYNdDWYa/eMaVwDPxbwB99QbN3i62SqEkaB
WtWFrnksZyJMmjW/U9pK7H0QP4Z64JGHsET8l6Y9UyzffrUvCPNl67esnqVKqyzX
Ggb0di+s0lYBuUuSd6gooBEUhA0Eu+fVzSI4CRyNedXrIQMnFkZ02EvS8+y0B2N9
7J1fYYBt92ZMfmvNtY1o5zLEABgNM8Cr1F/CCXPgt+Yz7Ta6Z3Eld9KLP+Qv6JQa
4qZZYBqHTlsKYniMofqOPmSMKYnfTrogE5DqmgB0QUlv7dstLKkpRmEK5Z6SDWJk
FnSCkmNUTVZVK062jf7iDrV0wUEW9THSfTKw4Q0nMZ9RGJjFiNil1bacSo8LAHMd
HQdeW63wKpSJGzV6kPDcgx80zAkmP16uQavKUr4wtczlMVdo/ophQJ2hcNFPuvr7
LVAZosacgAfioYr4UK/PEMDAcYfClYaHT+pZVx0szSF5mvXH1MTlb7KcDpaYuAjO
0/co/j7iMLMvcQf8DI2I9U19IXDYMTgd55Z2cac67yYOLQK8drgTqnA/lHKlmEr5
R6jJ6j9sGXQvwEcJjS6xMvHAbaGfJ2WXBti8ePxQfyHuxeVDIYJteyhsarZyyXyS
y+aQA7tpaQTJa2VjIaBaIJ8fUhwru1r6KzFmmkjApaN4r96rfKChVDTkgckf1SIs
newf/GeMclxNF8s73ampzfUqc4CnZsDV9b8688W9/qgOSH3y2ZMVhmatwUUrTSu/
mY0CHxDDGJVrDySfxYOdl3Gl8pq8KTUaJUXTQV7jbSMLbNay3Qdat2zoAGbeeeCJ
2/WmB1OQPBDujuZwdjKcQ6ISYtykl+ffA5PTKyel1WI3bgp+FdiRpfYXV+cB76sD
CwiIONaKi2taeFLhRRubzxICiFTg3g24BwYwlOjvgkUpJAqvYPXngV2/TSgagWQU
ZOiV1PvOVIYmxbEhgIGd8Jm0ZllR+PfpnWirvLeyPJhEJKeylncD2cS0DX0i0+bF
gJEGDUTGKX5HksBhfro/NTP1Wm+N0WcBWs2Dj0tcgeSsY2pa0iVyqVKCrbB4QdlC
Wl16bQto2wF+kgDzvZVVrTaAR7lcNSCqj6VoBBIVszW6oIXH0hfpL6zJUUDzv39L
uh5EQvEuCqRXsbXsd17K+1cn8Zi8iMFo02pdkzEQkKzlPmDdiyIw6EFwij1x1tdq
T7AnAcW94MTN7mJjCzXKV56y2A/B4bU6QStABlxmTKMyCXS3OjyakzWUGCQRTJW5
dt8Y+e/9SAQxFYfhB7eRhpxXf0x9oVtcIzTLw3Op/7dFKR0CZhFkxzsI6UyV4alu
KO7JGd4zj7/gA5A/Klcc4mx+gDPsHxT84J6cdU111533zp/m4jBjbhLf9JY4SuQ0
hSh4K66lETyObRKzr25aftcA82mU8PvwHgoLKSGStFA97KJehP6vsCOU/xs5faIR
FEzzz9od8L8KD3hsbT5L/OJ3zzI4cXY0rDRCIOL/fOtUUUHwsydROkghBE0cNGOU
Il/FqLRy8uoG0IkWRtejBGLP+ds3YkSCrQKYerpHlxk8I5bgNjYLmDOmSKRbYgGR
kE+FmyJBKwH8jgkZUTwfsC/qB3wi7zf5+CThiQIBr6cq8j7x3JqLXc8nZ/BmDIit
NttIWHu1rfrBwkYtJKXlt0cI4O+8kE5t0TapWqZnKJ2Ea3Frg2toqyG102xm6hcy
HGglYlPsnZnpDAXflmClKYcWmuwiTP5aX9tPJrbSt2/7hHCAk/8LA6ZtD6bmhKiE
IWeTW4L2sQ45odUTEpDd8yV6XYtkLPqu4gKCJz5VOvNFZuEM23hpz9wWI0Ocd75M
r299R9T/zzNagbhc1RRZZwX1ANxrsJpt/XSDqLHxgyMqFr9mw5J0PYLgmeJ+XTxL
fTDDFniprwQQa93ND28/54XgatVeG1Ul2jq1jrERiWTfigx1lcZ+kZo6dVaDZcOi
YFUvjQXD/1aoyElCy7p0j1u70sr0hFfS2Tojp3Dq9H4f/hjl3JSLpVwVw/kIn7kC
bOlSw41KOlsxJ0QaOM4luyHl3y6wikbtKKU99jRnEtQjoQL4wTJC/lr2DcWqywcN
2anDDxHYBIo3FlI89R7iawR1IUwYxQI0xBYe0OZ0uat4yiRo0KwMtC6nADYjY9bt
s+G6ysPYhvKD/piMuQ/pAWDwYaZ1rfuYUmIfxejAgP/lSAq0Tqzcg9R8VD5VSQN+
fK/0Oxnyo4dGb2Hn6/3OQ70ghtnXZqK1dKP6l2u/UFjo+nXsZDo+VzUOmCbQ90VC
tLRsyVOhe0nb4n+B3tVduANPxOdBTfxaz+7yTsqgYaXlfjVE2+Qvnjwhll3bqaHZ
0gySSq8Fp1sFQtmEQqaJQnYx/4n5375CSL2SpbXIts4i36nnCGAC9Z0W+90mgavC
K8oy3yPV+DC51ebeYS8cUjuMqjUhOcPUEksPg8/TXs9xV6ZHOQTQ+yivnkJRy5RP
zLYrhF9V3352RKv2mSvkOynsm59KW1VVsG4pLdTbQnetADE/empU9rxtd0+6AwIE
sjrYoTFXKAp915bE98gLZGFP519jnHI0wWxZTtBFLXEcTLa0c0X8yoCp1V81jCgw
aSlUM3LVkHtg0nk9eP3cUijJ2pwHaQsUegD9vzi5PVgdl+cKL8k8TWFNtxeOfu1O
631G6XWhnZK7iTO1IlHn2C2B+k8dMkcUfDNyc607GyZ7Z7lFKBa/WSDyfFTnE7/Y
oLezlv66Swa8dH5OKGRQnNTjbHTZnhfmGioH60bNjvgPSYtbevIrzPixKmH8P6rn
UsCWLUdWmH4rb30iGKbHADZClCxJgSWk3df5FHsWHHQv6SRnu1sqveBFPBFWny+a
mgBC3HBmai9HY3c7hoTaSAQxG2e8j7GngQSkSndD6LinSa7zoqVtPqsRffVQlt7A
7rVzrU9yUdPf0W40yAx1D86uZYMJZ97XIl6vCEKqQcKoeZ8CV0LNqJQRe6/Z1uP5
kekfBNSJ0zTWdRGkZbCA7w6IpFRhx1u2zA/+hcrsk2UKMZOBsFDP2N+QvZoo4WfM
jiCsPheFNKJolh/4MzCoP8D6l2KV95AqjLpIcZza3Ar6NNDXA5072ZZEMFIChHgR
fp91aurCKiLtxvIhgGMW2jB5EOFErxvEsjuFsX78dNz8qWi8E9zC0BiiGxn/3yC3
JUe+LmoeSrn3HsdkVuj+hDyypvzVcPqlT08+kfbqlzc/85NY2qzMYD4B4UqMPLNo
m9e/4kislJMzvY/wYdtZLKPOc94rPbKfVYixlUA0kMlWlkkStZb+Hqf8/1+p/BZA
FGC+cQARVrjVG5QVtOioEYo6EZu7339EnWxgBsuI/mBjK0wp++lwU3oEtzqNkhEM
kNbXVSOTfkuqaeOK6POXzb2JUuXlUtzKvrAv1pQzEsOf1Ryiq5XnQoSg6mNxlNC5
RRZNbZkiPNk9pLa7BbAp+elkewgHp3fUJz+2+rhHyUajnoiNlO4USh8c2q45MEYW
aFavTgDJIuwwtPhHXm2Wr+44TLxewgbEzGW47Qw6YSX+6/bpkMrhvxAuPrjgI90S
RIXrzVX2Oz8VgurnFs50T43SxzTAQtW2eIQUZmDvssPyOMDxAJmTW8FNAlT7XSmv
8biW3kUCaTTmANBqR4QwxFjmmv94lQCKKjBdF3hXub1h6pGjmg9nljUlATF2TTMc
V4xcbqob89g6ENO2a8hzpnuzaN5D8xEgPBhOI8fCtGOhSu+pAxTnwcqKg6DcgtLr
2SnNDdFzx+75tPOAQLRt7mlEa7sGkOIuC+85DtXalAThPKg8/6aelTmYPkZ66SBH
HxA1/vO7AmugxHXyN1uDvCLfo+0ke17xtPAkzrRuMOL8Sa5ozWdY+0yevDj9g+qd
1Xfm1Rt6mgpK+2+9KCfZ4864VLk/Yvh8pRYCP6dezjwEiepsSs6QVR7SkgZLc6jQ
bdBzUPSx1qL62t9sPZ7N0tIJPz6uXhJhU+QHQpHU5qjcxUHRwjjG2Di77QL1eTta
8Q5vasosYx8c1FTlkTLC9NVBQ1TXNDPDiLRTcUz1jfPf8gsSnalybBPbIoSGrSNH
37FdHoOxtn/CSD2kdPMJbGykBdEcGuLRnAdcOFvKZwemTlZ1vEtmxaoFfalB32o0
4MxuT0umvwWSqd8aScKKuNRNJJX8xfvrit1F2+9pnnoyFgBw6dRALbpOKq6g4tk3
qeWga4ZNF06/9YQZSLcd2HHJKrg2VaCd5/gcEfWmHlLaBjtc/beTb2VzxV7hx03h
/JhgQH3wzKO0qyK/aqc1a3adcF9H6gT+ElcaClhMHbUHNZ9rRlhdyTSIwfadHBkv
4JW8Z24qQpsNZN59H2GpZseinZnJfuzeHtjEYp2KB7CgsWAZ9wcLoU6fBxvbdgXv
Gy5Lxiv/yilvZd93u5YWs4EgJF+YRMxjEDo+8qqqKD+QJplXws3PeU4dgeMznick
muHBoxGsBUnFtwgg72XAVKqvFzF8GW1JzatSAkCSlNCS+PdVEQAhfcKZJA1jV1cu
/b0WKUXQjs0TzUdQ+wkR7qRF4w2tj5tFzNKrXjHdVJWKrZNU0JpCXdxOG1VVAbl5
qDxNqbwiVQhUAfW/NlekyuvPvsmX8IqVtpRyrJjLZAkw9blABfm2h/fP55QyXTw7
Hi+OAt6aHIgjR8ut2o5Vt0u0PegV8SpROUltaLDoBDYuar2C+oT8FJRN1Q9ifSS0
s8vUsqqqxSqxzZAQezt1K9oO6STCbukYqiSRPYzKSCUPw1E0lFUNU4jhCftORJmf
OHApxLEiLZPkB+/qpZ9Nv5oR4Ae46eAmRWmyFH8ntZ/IfkQn2+Spbgj+UxtVviiW
wSYF6jRIyWAKoMKbqV9aK+pgkaucxP5nrDdOMqK2OQRvBVPgx8QCBw/m92HGV09p
2tz1f28rjQMZXpDin7pMZQvxZ+jG8Nwp9P7kxKrMwsX/ffai+14XN5u5+SnJHpdr
m3ccNgUbADAVf+PJr8CAF84ELzGMzCRQVae6Z4JZZQsHo2XoDF+UNILIn2Dnr04F
+AbVd4OqLewTfTV4i1ZbokpACljqOV9YcE5OHjjrfoa5vVc4+e7u+4j8DNCjo07t
WuaTcddDuWiNHQ7YpK38F2ECQDjxeoKvyxUB+xltNLkJHE70xg0qqFdu8gXZemN/
B5aRAlX8bWrs2W8ltN90JMt2wIN2E811G6jXlEq0x/x7p8KApSKKO7DNdhbVk3S7
Zk465dKcRzUOUa5MdKdifEm6iVEC6HunGLK3SlP02p9z6TPYW9VCMOlF2ogZZmyS
eE9YenHZYGo+oB4DuC6+1PlgZH3/Ygbb3sLvXOVe7aESkVc4BV+rKJGinZlOSwCf
OVa2XqyZg0umZqIWaWsId9o8fLwLxWjQDCvL7a49FABGQcjshtrCJ7Z62YZ0G+eq
KPcsnyFZEy5eQH0UD1PazNb/fJu7DG+tEn5BpYhpLFMN5MlNge/bUjWKpD52JZFW
SPFtZ8EWet4ALf64eXWix0FxxYFIasD7QLmkhe+7Q3ciqLXXKtDlcpCXClM3RrZT
Ga8Xy1s5AnhDpbVX0bJFOoF5XRkcyukt+HFZW2ydqZa0XiiyvV37VMeAKUYJAKx7
SX+SVBMYAJ36j8q5kE7KSAU1V6gMyhRatI6tLGQpJ+ze3Un3mG7dOjyYvIe1wyef
hufbXND+WwHyS7VRdkNl1BWqJwbtxWkp6T+Of7Ny861boAY3NFzTgI5HloFXtnTh
4/EARhy2HjfJfLPo/WI+lFBxMw2Oz4Qb8SbBmnHRZxfXipElJYw9nzLNdyRgVvV9
WQyZ3/4+oSSHOSvj2+wtT40t/ESCfBZkFxr92kM8jAt5oi84dOINrR2Mnq2r4FoC
taQJK8SOKk5yNTUR4jB4W9QYY+9+ukjZWH5u648b+NWMd1L+I5zA5cw+tkiXU8Qc
2GB+B6wFE2W39w1eyTiVBqlSHvrK92BqSk3uja/kwjCOxmn/rMjnuJfFn7IYQGi0
T6ItSnPATKHB9Ol0/OwAw+1dtUqnOAWwXOq0371eDcy7OKWvSP1slKyOBH4f6U1O
NXHzZFUW25oPrqrxE8H1o9OVwl3NBG7B02GjOkky4OfoLf3L3zQtcHOrzegUz391
bTeHbVRJoTWLYxhM8wE1t1aKn6MLXQSNg7SLOZ4eKkJ6jJx7J682ycWo8xtfccX+
dWDzQ/8uCWRPzwUUuRDClzkBTevC1TiWl4Knrg9MVQl3AHRqJh3d11/yrUIYjvFB
CfwFanT9thNmvVH7l4Yl6CVFr6ZCRMxx72jVdc9TOfu2HTTU/iMvFJZA91JtumGZ
LuRGYSJk8A28pswVpq4vLsgRLOMQOJLWh3JX8jETbF4N03BTviMLQrOtLn9LCZoL
XQrLEVYtErFkzpVQij9NJhIbEqKZKFDv6O61KJoHVvnNa0ILg4YRUkZXBy7wjpGg
Q9AcI7NMVli35BCh9zaHz6LRmT4meQtpxSnYbtGL723DXAXVQqJOIHM/pwz/nSca
WTeaoOPFdXLmbnZ7xbl8CVTkIFAOTE6FWb7vbghmx/Ypm8pNeVLaKRVPvlwmkOX+
sDcs5w7M0OnHrSN/9vQygM+BVIHp5gDUTvUCSGFE6KY/ChrJbSbhkRz+m9HGL2bL
YaiRqXIeJhvohHUon5vK3d8264qcTGLEQ/uTvK1ni1Y7hCkw+p0ZpqQZTxJzj4Uo
7KDOQXEDTPcQaZjOjAbOOw4HTd94vy21Jj4ts0LiJBIBepHDwB2Nxd7e8Q4xOt1S
VjktvBdhpN8VXbbi+Qgh/nLsRGcnSasli40A6fP0rGPwpnUzRkCoO76B+wrg2xDE
knix5w0wZp5OmylNyrvEdAzqPXhpJtAhhYrg958BWgF6q5JemV3kN2ZMPKyt4CS8
45nObW35RBq9S7cKPTmHGwGoYC7PbKU9Nf8+VdmWKuALCPVPBkT9u31lYmsR6/9J
W7YCEofiDNBKm1ELEfXtZ6l4Ozx1Awm0Th8TvlmEd9PLktp4f0U1DcVYxdoOOaLx
eO6RhidUUQFsVhUavbtkjOAfyXNi3BoTliKmrzWoCoXOwhRJQ00wpdPeIT+ivOkC
Xh5uKzBUDpDZKOuTPbbhluBAfJFLfCPyAkLfiATLwmiZaOngoMOx+z3Wz36l9FsJ
xpx0qLW1r/zCMpynHmYWTl7sRtP8KaTxkOuP8OZ9c2Ftc8boTOpXEUCFqZL1Txn+
3Cp61F5P9AX9iEhFj+N38eKeFMIieXg4AEvij9Yr4OETezSP1Vxvwy+f881yfagt
r9qgS+UA66ELYV/mDDy8G9/3vDhG3WKbTMwgF41QiZZGFICJttqO6awHrRs8AXXU
rY9YSrGlAG8b6yNmU1IwRIinGQqXZ9futKnlRp3zZOa34YNbBIgUbaWZA8YzGl3P
Syu8Bt4NDicH2XoXHphOjbe/iDY02KraPrRINyVbnORLRIpZDe1ZqzfZF3beW6b5
twQy/XlWO/9uFcQXXPOef9bSMjPVXl6Eiw1mTPkDHeGJhnGUj3Ruvj/ubpFMdzOO
eoe6FCSBDRSESRqicZhxn/+Hc6VVObhDTT/j9j6pHruWJN4HB5s1Y0TLKAQ2HwRV
hOxZPL1xTMjDt/lJYcrf5hrA6faOSsYUpYVeZP9ARqgaal2V+x8mhYf5BVTiURHl
G9MMzaca10YiKHk7sWpRzX21d9rZgepjYb1Dkt+S26KIUqXXVWpdRMZ1ViFVC33Z
69kxbaANKZE2yoXNdvDua6Ymy6KWpjbo5v/U8CxmcK2cs4RPjpFLIInkvc7zf3q/
CFzD4QOKOI3KBJmhgNVqhgbpyyrLXYlhKclWYW/t+vFWsIgXgywVLgF+JhXmWcVR
p6ffVsKXm4JgGhLyUGDmL0mBF+hw1e0C+/fh69XWafNgmGMTH1Eln+FZu91NVx81
gHzrHw8nVFG0vwEWle/vDfS6T0cfbf9EvBEfK+fUfm7lIXu3QflG5kYi8MFXExdq
iZlDS0QHdF/CTtg+lojOWd9txqjELPVfQlL5rIHg6X+G1x0z1VHVs9OYXHZB4het
zWm0EP7yztillJW3kJUAnZQ6VtjXZkRbF8Qn9lV5X6aGk4zGHcSOi4+VsNjhcgfL
QaesvNWA1NrQs579lUT5UY4Hxq0RPBC5lkPsKpsUoH2nkwJi31HCVHzzx5VTwr29
4+TxLfcw9JRhAvyVOpp0ISVwqB/+IuAFtHdiKNaALyV6d035iqzOnwGuUCu/ppi/
+/Uavxe4kNXoAdJ2KFgUH2xSOGO2/E9uI3bNRGrASF8M7oc6e8TrOVgBIK9IRDnG
jiW1ajOH6HIJPHcVYRR6dfsXrMF7d2zhAqXuV9s0boZ6qu5WVJ0WiCpOoQ/B/WwF
Q5VpTPIf5IobOV70Gtpc3yIK18goDWNfcJmFs8uTd0YVySGelHLxJfscEYbG3uAT
OVVLqzUI8g7bIKGhpjtM8lDAbp+byEKhCBVJqLhwIvBqVFrIBxtNBAfJt3KH4IDw
JCYwTDb9+pwB0OtE7ACPyBB+MpObuz7X0I+QJg/dKHeRf3VgoFHSlqk+xqHbdeb3
bOlf6fedPGGhsMJWr+P7LoZEzXXI6KAhdbEGNqbz12mW3cAC/TKMjJDZaE+s38VT
3GZ/CNBiDDD+3rTnFMG9is3Ptd+732zzHmSZ4roM4QWTy+TG7DLkCQj1n8n77rLh
qzP9gSRYIgRj0HyclXkKObfqOLrHQrqWRo9Gw6RcI6zrABsiHOjwRCWFt+MVW/h/
AIw/+axNpKLusiarXnKLdoa3rRB5MikTDO6UlVwkBSXAekuFpoG3EixVWL9Ht8GN
IqrmzbuV3XNq+6o6biNOpwAf9XPH4ymO/kqqb5TEdRLwbkU4pcnN4HF9BVbPkbU8
xNIyOgurgF9WyU6omck3RFD/B6LrzlpTkhUGZga/8wtCjzC+xMLYneKj/cvX/wug
3VkBzAT8NvZOWe6KwGO91iczbnKBxbgVRURf5pkT30ugJ/XbzfuxtYYiBF8p6bSw
XNAno5PfYgOrpTwR8TLux/gTNwl4LQEo6Jndic8tZsxacc/xl5pTB7UMppr690YA
EjNQq48dUwa5bBOe73gvcj10oCZfbf1MxdJQrKTICMsHpFHFOj1w1VwoYdI+mczF
XMboNL03NvzDLeayKJTEFUpSfQhyTz5htqx2a3JE+VNO/QfNErWn28QnM34PxvcZ
5FwRIvHLQ7EHod4XJzFQU8pSbN58BAEgVhB24PE8sqcQelgygWz9I6630D+iqi7I
L5Rt9d1t6XCMPWN/wTgwoQX4JNIld/aHI7L7fPCVj0wxqbn7quQGwpzCi2ubohoT
RhA7TN2/UzuN7uo4qY5Qk9PryyOX09UnVFaaBrMehaF6SNsql+p2S4ZvnGP89r37
q68EJpOqhPk17D6aDF2ifTWuzDINq68RC/BrOeC/4lQxdQHnlxO9DQ5dcLnxd7Cg
d+fZZLez/8RS4RRyrzEXgc0ImT4iGDYnMfSZhy/ypHuj7tgw+5bNyaSgRCh1o/3n
yB57Op5W/88FHOcYZPBvuOEcp36BcYHrQ4fVzWwMa6q3lsSMKfKO4qVHtC0iO0to
WSLD+mOqpoW1ReuLkSl0ZggQATuobaKK4nDi37m/sAdKe4A7ND8mXcGc6TGyq/bs
BbZu8TX1/HCojcyQ8c/QoSWxZuHI4oEz9QqRtRA0/p1r6jJpRJ88zTt3vpQLKVHK
tXBu7k9rxRi1iMGoO8pjicRNo/p+b5JckKY33jvAEmlh1f/iTm4deGIOhD06cYCJ
yXRE4x/k9L1mQOqv2gx5OnWhtew6LlwI8diJJiHebXvo1ac3wcZme+4IzCuOoDWf
w09mOO7+yQXJrBfM7kOX5Kw+lvERjyN8x5GXq3Kj7gxETcueleQl6uZOiRjCuWBN
yGJ0UzKAN6rbBRY3y9xMTD+QA22JQNrZnaQVksigPGhpcFFwHZQLsI7mWZnPCH/k
jf2roAWdXfzKj/Yu6HtcSW0GrV0r2O4x0gCcNHr1owFC4Fw2Zzu37jENG0RAyYD3
Vr7SfvMRYFyvzuUaM3u7gmJUfSG79WVHF/qE4ysMq8CLS59l11voBJC90fV4DX1l
H4lYF6VIS74jzdp0fXGoXAGvPspT5uxltLGGei46a4LUdToD2JLOnovED5FDJAGu
ee1KaWwJjJ/kLBKoSLJx3amYsb4olB/Laxlj6q7E/vVM7DOXAhjpoC76goj6kps2
cFJlkIyRm1iH1FBk6bIenvREvYCZ+Zz7ZQrorEa4rGQFYS96nxxin92DHr5WAzyI
tvrltDnMyrSDwZu9xUxoRlMDLgt2iFploz8nCco/TLpdRpgKqTvSI9I4czzkdZy6
JrRrSMqiDOA8s7eWO/T9QddZshTmEZOwYCps2DVjk6EUDjRHqFp9Mk9e/voRItFK
HfNirO3rQiSS+mab/9/KMLRjkOLzgmCPII8+6tuoqBM5wGpKpgb/XKRcVhZA22PY
rvhfr3AdN+Z1mcGlNJAOJ8SsdnX098TDTLtlM0KeDR6kCvO9ymwrwxVRoL9yncAX
id79D9XsnLAxKZt40pMJIQzVXxDN8CpruN+sTCLh9UuHJmpUGvx2gj5KaeW5yBHW
PujhDvKPX3Sk+3DU5YA26eWNQoTOtsaTYQS9/bTDLaJaODlJhck0SmS53imfipo/
9OVuN3tnlX5MVrtAj3xFK2zvUy/z4JO1LuNBK9+GqcWCWrRNhQd6WrRHPtW7zXEb
GSJptYuRkQMDF5vAByXZIuwH5fXsI9h+sz77TMKLoy4tpua44CjQ3WWF/uPUo+rJ
4Cz+Z3EvRurD/qUZoGv6RxYtJB90y98m2OmW81wZz+K4sy/nSCOgtrUIy8dZX8nm
dwNInO57vMTI5VqLVYT0Sqem4fTz7WkSqLvsy15XQz7dBGRvj21jSrKpx6usC4l7
pu84lHSRP92BiOfjlM5j/8f4E4460jlLBWW5Teo0sxN6Gnq5Ffc9wMBdWCHy3op+
dahNtKONhEv6C7cfqQOrU3sa6AtaBXgR30OBVAVZQDwNOy7QJw44/zi/1tDwl+fX
4jcxgZxuVqCq71HIF61+VFY8+khhHdVTDBq2uySMlRNJX9sOFBhYyCWHznf2zsJe
cI+Muhmq8pzn3BG74n2OyQ9VUQeWyprawEKk85aNLuNhmu0PwVSLBu/kBQyvGjZS
S+0wY2AmnHNhEfyuayCdtw2PKLnFlwkRdi8pbwxsiAKuCoAdzAyWUr5gaFecf/fJ
9aMl/5n4yvXtbU+f0jHB//DT37Ou+E6GSY2NWfE+FLE8hYyfnYOoFfJNYDrwxi8W
kKX+DO3R3mcwsRKY5ccJMeQnUzVLHTZQKZDKVgWZWSc4/k6PgrMDCRfE/SH3RCCP
D3LZYGJ/q1hAY6m3seWbN4zC7z7M7swewdDOQe1U2332y01Dkt6u8doicGs34aEs
V+9I7xd7mjBaAMtwg2cQaVTyOAodadU8EJVwZz6q/CvGeqo1gnefuBGdg6bKFkTy
Ey/RnTQuMTk3WEaX1UCsdMGBmQCh0HFUla+jwkuVOrKcFb8KZsxGz2vho5m2NA37
ctDBmY8yU211ckISMYzFP45RsqELCEU/P0L04I/c7yPyqGZkDBYQztpaZmX1MIU/
pUsht99CHZ4NvEIzoAZbkEm14VyVpJQNGoaHWfnGKVlyeOzofhVPXg8SMHBOpyx8
Uq3F8VCTEmiFVfQDvDPcVn3Bqit2Hiq9L6yOjgbEMcUHmqhlFnzljHZl1kPXov51
G8WDpr0qSliclqxzs3wmDxiUk8tL6UjfJxiKq16Oh4HxW5GOIPvKIdRMyFXBiIe3
lOFDBRwuHl4Z1Hobh+wKIXVt+SEEqVpjYlsi5K9FoeuDg+DnopYBj5MrjTuHchO6
Wf9b2EXpmaxMxc6OT2gBET1ONz0CFs4nf+PmQf9jSyOfGHcjisDWbTVbYyN8MYri
A6ldErEi4UHAqY+7VOewmMXhSINKGBTU/xFxMNP1kH/1dlBxaqsF+yuEfAH0JahC
8If1Tw/OhOZwdr/O2FSI3pN9e4lueYWf1FQmJpGX3DN+FpbM6dQ4kOT+FpGMK5t4
WOCgdslDtJqwpUr9mjSzyQcLPtuRzFFuq3Eulu7fYb0R0YAGajW67pA7LIVH7kVY
MMEx8CkZzJPeqv2Jiy9CNG4veOm6pgUi8glU8WpDv992w9EG4XPHr2w+uf90Qcji
WKZOTl7jsZqzgchk5W/WPtgQTAYavFbjf3uOce1gk3ChztnNp29C3IdYOtUSGY5G
gMw3t+9QQmfTOLsPeL+IWry1DrQQqQGcrfnpiMsywpMpbG+i2fZStC2p5GmXmUz3
s4BVNAS6tl2WXBTk71HyLM30MwHZnZ0Cp4JU9HeYEasMEUmte5+UAzS1nf7Qy04V
utbQcn50i8NiqIiPMLWWLhl0FIcGa+IquXsj09dtYbx+W/QHb69/dXfTw9itLtVD
bGPwZ8o8AMliTYG8BSJyVHWoY3p0oQJioJ1ojocrB/Back0t79tkvha8plJxFrjK
0rOjjrxAEJsa4ocMMjHZSUg+BLNr7JUDA/4m6AolPUKuCGzcwIz90kspjOGy90Cp
ZillwDP+cVbqJHEhPscnD9vGNnaO8EfzZfb1n9SG43CPootWhpZWLa8ovSKd826b
wtbjqIRUiRaU9xWSSzHC8uVD1afRJ3VDVXqqD0WH2UKBWVq7DpYVabmqzKWAmcaZ
bR1Pr8KgATmqCsvm7UFBbOSPphUdsB9apAJPCjQNDohQNogEV5VtU6O+jZ3t3uiX
5H4bfnOHT1JmN76DS8j4dIrQoiOC6Z0JFlGXXTPScjtLrxNergQh32MXyPpPOJEy
iQyYZYGN2876VVgrPYKNL63iWBAqqzl5U5A4IdIGdRa4QdZB4xjpAQv1tu0TESIk
wozfdlrgt+h7up5YAUujriOF+7cX3yu2vIRFagBfIH1c6f6BMP5o/TCFWN0W4eVC
1WpwoAc3JN+g1KVXI8J86yVp7kgXZsLCAHBko2clWaDammuMireTKyuo4uCMyyj4
te/60evvhPvqjw5AXL0sffTGQdzQX/iqwBWPSKovIleq1NuhJbxAjFS6XvIJjhlR
IB970G+KsgwzxyLqtiJy8o7gCMtwQGUZ4P5GpxhdFpqJy61kFR3gZKvlicN02cum
gtSEzN8WDtO+j2JGOpQENfINiKaGI38iFjk9VYy8eI6rltxzf675QbAYXkk+yFqO
NVae0ZC0IjS4QQAc3Vm/g9y83RE2LzTkSRJOn369BShAc7bwDaI8HpvuT6Mn8bJz
GelPMjLCmm93ny79EU8KlKv3zMHufseuTnYsn0Tu9XNexSpZCcn80kjIYQcaw2sM
VpEqX4Vm5y0OsXRrv70upFZP3S2gpr2CS+LGCIKtoZ7Ptl4dyFGYSceRbFo9CuyS
Xw5vu/QU3BpJhV6BohWZHQC6XnfgGgRtZ7o2g1q9RTbvd8r9LpK49E6MbNQM/a+i
KKxrNsw7/vgZgux4yLAOa4P9m5d5Sk07wvjSzZTNfxXrQSI6OAR63pAOFztUlgap
PfNsCAiY0q5RBDe9iBVcuWh8Bd8Ib+OoNqaM8sAiyn127fXNMM5XxTqdcB29YDJ7
amm2D3ztCVbvAJXcTBniIdZ3AjGpBCUvzhGKPUO46fmpljbkzYgmsxWqglhptxfi
R0kCIhQRFa5fk8zAI539H9L0XOLZO8raPOD/RlyNTMbksI/kaOxYNBBpEg0CKOM/
OFl9x0N2w9b9z37LQADGsx4TpA3Z1sYCmgla36x96P0HEr81YmjRFxxPvmQO0ySz
lXlKO/4+HrEwp4WRt3EwGRIv9GlgAteEEnrpNYo78ukkxhkSQRnyeY1Sk8PErAHp
7uBRGnEtb8Nr4LiRYAixol4FTezIbym8WlqtYKI1mEqbC0v+1wGZO2Vosmjg+k9Z
DRRxG21Js6O81AOn0uO54ORT72Ogbols4LkW5m+XGetP/beVPJEbJC5kN1gMhkJJ
8e5k3ITN1WndaK8vsNn/FHvV6OHLWsLVFRGKSfep8rGqkRxVzXTjxcsgvDhvivEJ
A7hMP6tcNoLo8Qo7xJ7mfQZ149/01sebuR3RkwP9UPjyiX7BwLwLKlUN347nG51T
6JX4W3WIkXdQkeQCqed4RDf/ysl5HkfKg4hqCR91R4y/YL7ipNWXTT3964jyN1Fw
EPm/Z9aKknZsqOjCGy/H6XZ44Or9OsE17aiWWdFptZiAVwENwghKPJpxHZ3sK4NS
AXeYpVoxXytFGWW/wZBSi1CH0woWqL622P+Y9ACFwVhdm+VEzW0h0k06mKaIE7gq
WSSuFjzfojrRMjCa7W1++XoL34MlWO1L+XkJsanQPilbfxxkT0QRfDQY3WxRXGkk
Vvkylixdd7ArzXIh+QhMpwMbYXr37e9HvRtAy8+7JXsOdR/30c3Ix0MEAa4kYpOy
+AsKtlg1eRYNnZbWJgmZd9kfvHO+SQfIXlnvsPKBUJI3Nnb9mLtdgZHSeYs1hXeS
gaDMhc0BMMLwZnx0AVwywupewTB9/9QIDzs3fbQnX3lsXr5Nclky9E/hHeChiS5g
9WtANVA35nUxGMYh/sF7g0sXiT6SipMXyBv2uwISBrkmC5A1v//i0CmQi2ht8ArY
aZ/XaIN1mnNGNlK5MWdCaNfIPBBHbp4eA9xGPpBqPmuZat7VLmLsysxmL2KVAhxA
sRW0ZaheJudKVn/DduSq1tg9EzyJ3/HQzuWICLoOcLx5pQSprZ+bpwpm6pM2te/S
LOLqXxK15k2rEquLj39WZis2//36o2oZ1euzeEIrHWLca+WipvujaBVN/L6FiNd2
PoFbt5dZvfmoX8TzDLQovGg4Ul3BgmTCDAh3N08QpJpKpNlwW3K/OgjoLnWSVK5+
N9PeCg7Pv6s66SpA+e2jpvIgBLh94CqMttIux4XdfPdygGiUW/jpQbnAOhdXueSc
6zsAkRXsrmvdAoHDIRa8v0xlIibRMpDbAOuTUVUHagTwSRlHg1SQZci1HmSMA92K
BzyFXKayISugMkXEYQvLo1Lz7FuBGDQNasIMcdVAsYuZ9Pn5hqzoZf+Uj3URfgHo
EyfUEqizzaGKar47mf+fKselyDJvKLHsxKHL9zd7q14CyVOL82KtHoFTrfcgj0LH
EDD93YNTgZpG6Crnzx7gI+d88K92Yg7pyFdq6jAXbM1tSpP8H2uX3+pato2J2Ofe
cPVVVv8krWGbQdwH+Wj49NiQB5NrOqCp2TAlG6ND0mnQBhnNbJl5+CcL5tS8IzL/
RTYX7IKGkzTEJL7vQ/+QN7/DOP6zqmU87k36zAsdrArEHcCDTuDzcel2T2pSKQua
XuaXC2iMSTUWpS2Fz3qw8K6qrrS2YCrM8TU4GFL/UhinNFVarJJpd3vE9ItEDly5
SrgEe/mkifNo0LdbUiQgG5L2EYfMDo4fepaJ+HnH2N0UE6wh8e2XtbaRucH2S3g+
Lb+2gh1GKt8X60pbU1yO1jq4I5XAJbG9DMHTH1CYQPUIVn7lZNWf0zpIm96DMmBE
cSrFzufvCU6Goj32IhI1iSsIUS7lIE9043e0+7+/C9UqEyhQbxEFBejlwjAJsT1h
W+XZBWQBkgVRajiNAQCGTrNx5ckV8GAn9Gmnx02Qi7OzUy9lTHwHfT7dSlDuorAs
1RX7BVt7PA9cwPT0tiK+3ih6EaerDYvqjEfRrrtBkmeCkBTSw6DmAcOBBKNvc/qE
/ZucwkGIvcyolF5kUWIE0Gv/1nrt3p7NFJjAsuurYF0xGBLI2rIo0+l+iyIXnYCb
6AznPoYro/g1NllNraluSg2YGb0pwu/ovjHB7ttnUOVUzZap/qh1EZ6sfeap3LM+
uNwTcs+jFma+qtRPXMLvqjR+6UkzxqmZtViTyK+xIw2rUHwW2K2kwUXX95UBtqKZ
evc6KejGRmp/Z3qn22jAU9DNt7dPfM4uSfJXZCfdodEkfrL1CgPndQhLt6j9X+kT
wmJkxHus5bQz+874LrFoexZNVgpW6KMgL67qbX6VEZv8c83p679zkUxviSi+i6pL
FvwGl0afPIDfAbv6qsQCwyLneBhtFzUU1WWhvkQRk5H2/I5ptjvbgctiLq1X9357
xlxLsDKqwaSoB8d5doDQme9C2x8TcErweIWaHzm5RQ/NBsVd/bLoEaC4mtF5eF0y
+aYgDtIRQXJwGecIvDs+Z2ayU3B2q1q4rCCYmtPqxNv82sBsEwsOkQ4sNULtK3IU
ImKWhAtzqt6pMBu+BWLCa5XSVfcGoYJ5nlghDBqsjdJgm9bel88zw5OOW9+PiDgc
AY9fY5uk9y2Y10xPfFzQs2Uqm+6evVHvxEFfB0LaRCxLn4hXjraVhjux0LpW4tC2
1Yxnnfv3OI5RZrnIm+1CTjYJbaW2HGZqd/HrGlX9uSqghOTZ36+MeZaYhGSqb214
3Lm8j29MoJOfifGYiSxJiRjGBEbJaqiwaFwls9V4MfEfTx1BH9OoQrZlaVJ2Z7bE
mwcw273/xyoIW81NWE6CGqCqvqVVyrwJQbJtEEdVJBnbKG2uqp0cjwSQ+8u2N5qE
aBrDpvw7KJpdAv5xelCcA/DQhFqvhpNGjyB/4r5wVm/4AJDi/pw50YXDXlCRoXw9
DUWB2mZPMzajJQHPQvqTE50CiTlHITGakVMNT/Zz6IMWf9X9fP01QRDXR2l9YnIr
AGbhUmF2Z4eSee0TTxtMB7vMhMqHT0JFwL//bfOA/6R/876AbMMjZvlp4Q3wAUaL
gFky0Ei4UA8yBEiq4QusbrNqrM0jLfcQC2enZbonwzh+T0AsN9mXoKw4FqWKUF+K
GcLRSz84vXG7GMoLa7jFZfY4NmKE0wNyOMamRYojDSxG1hAazHqvaq2PxVV0LaQI
F6RKbQTRO7xZ/FGtTk7emkFe38hURJMPqUORWDTFGi6UxhtQPvJSL8CFAyZfr+aq
z6jwFAgimFfVCXBoxzsr+BKqlkloqsza+sG4potidevcu0TmfsI3lnAqrHJhc1hU
Tpk0PrxsHIn+ZgwRKKthJE+aOVEhPkfsZ9niIxtScl4FtCilPVjUBLfk58e3Oijw
K9zrTD/34APMj64k01KuNZi+GFbvVFmEtxN6lbGc1y6LTjVYMvaviZB2ZZTmoQ9M
GLlPov7klz546MhzUfe8p/yPTcN/3xfZcJDCzlZC4iEiwm+bppSlBMhY6UKlKcaY
lam8WCIwDTFYghhljozf/i9IBCwlu+cDAojdhpviTBWIhQmH3PEcoU5ZSfr8ELZm
mGE3qsb41mEwU2856SfF6dh0W3OZXXtUNWiCH0YHsd5n3FiIyTRTGDrQSOxdbiNM
6kPOo5wMWtBVoO9bnTc9nX2QQqMKrjTStOIp7x4hauQ1tcZvIeChbHeJEd/5JaGM
CvfwYJTehbSRUvSu+sJvEJUNDAEfcbAA4nV0x1o9+efPkIjAO6nvY3TtHCjowQ71
2frMaOZMqjLIufQX3xZhkuuxiq3iZtwlevauxF/GjX4lQAdxAVzXJ2QqU3IWL+Lg
YMCV1LHvJoICNFXXqWuRk50na9B36Bkf6Pk93rNhn3gGtCNqfc4WB06YbIogULpN
On4dUmvaU038EpR4x71FQvb6zQcgzdOlP841GFuFykM7cfAqWthVIxOvrqQjBRka
fGUHTqR9BVF5oY3ennliWTE+DUgNLidWjISPgLeNmS/xRx5UWItWyrvPLQOnTb4k
gVxt4cMOmcKFBT3D4lZvgA4gDJyV4WU6J2N0hpVUKuVb7B8PWjHhrn50S9bgWFvm
WlVdwpSG8xky3UfAlNy0mEj4yOXDtq5JQp0V68AiqrX7nAE/m64cCWhxCJG9ht5G
6sWph7SoZJq08N+2wsTPoFdlSWuU0AicDIMJkGv/7txR0+TkZO8JFfm9ebLUGZXn
my0tlckX1dWZli9IjxELC8bQX0TJ8AyOAkGDCxPC7I28GF58beP6dIl9Cc4duzUi
T7YwMtOQOmorEn7khpwdsZpd+aMeeNRYDhGUnUQ4XlIwgNLT+jdFli38/8ULBxMl
wfSkaE0ns2HjKrWh6xiSEqJ12di+R+CmjXuSkNrzWh/Riz4RUeked1qMpPeiZd07
EGjnfIoYRbHX4jyZk+/iihfHMF5HVzF53BYqho2zhEE+MwpDqlsAWv12wbXaemRJ
k875M5EkQGugyV8ZgDMENi8LtaIZwSnMWEAhehVfkOMFKAMVlCBCOoBMu7vQ0Yj/
nhjFdCpvQ5fRHPz5C4L/icJBr49G8BwrPNa9SqXKhRvioYjuCvNY8veHjQLFDGS4
Rsu2B6M8hAYp4QHJ87obSKXHig6zXmBvywcBNWRckNIHz/TgS9F8JOSfQq4ZK7kE
wx+soK/8nkW071gdQxJNho0aQQu6S3BGNs2cdvFuILkuWDtf1jZStCIgx+9QmmJ4
8B7wPvd0nxLaMNLOBZu1qD23RFfqKYMnPJSQk7zGjJvsCMsxQYJtBcerpvHU1BkK
GUTJUfs+L7kMpaqhLf/7ZF4GYSjZr/YJvm2aPXQNSJP9pn/i3jtF3hGwr8b0GXrC
uZS9pqkUqaOHxTkHfbFBvIVxvCdxibppeDai+83HMxZuJGeX5+GNt13eSm2Z1WmV
TKX0w7lOOcY+Z/tRIPSnXnu8kIojSWR8ukz0VumXAig+e6508V/wI05OQNMnkPIb
EVG0VNWekBaOMvuC01WHWnnFi0BHTyQi+RCi+lEBD+brqDUwsU5Bic/6OuSq8Ngg
kFNztbPFEbMT4/DxVo5awH56N/KgTkQjauVKULuh9fsVnBW85EDZJG52q4aOU1TA
kF0AAYZEl/k4zDd/O9kCuVwb4kRAcZ8XbfWbn9NSiXo6O7TiJog0vFt27Pi73zK9
lXzPHcNIUQ2965anAtg6c9XWjEPAwLg8CKgPWBrNEDpm8whVh/pHD6uJAhuJMzn1
E0ravIdw2G6YFGyQeygwjusMPoRoiH7Xyb7rEgLip1SbIe/UswPbDY9KExnXnE2c
8um90aN0rfDB623CD2xqI7/U/NZcD67P+ZEqtMypBszk9yd/vpMWtAVEQ4TJWeV/
94sR9MVTCNMxknjHudiwkugEsy88mABgvoSEUSLcvZppr0uzf9b3N1xgKFe3NlZc
m0UR+zg8ZYXxvAomvU4KZ/wCJYhtsMwwjErAIHKDJhw6ASYDTYzw+guG6nS+vPoq
mKHEhTB6u1BACieiQsLUnPs5d0L96chGXJznAMwRoJcfP2xgqxVbVtItQvVjXiFE
In7+1fUzWToTOMV2RqnhFxznp1v3nGXFjD0xWXz6j7XF+gpPASrlSFLiJb7FR4w0
+qziYFc5YBbM+7SrJM2B6Scmzh/KNpP0DjUjV/Hbyx+APJ+xPIKvQohhjukzhn/a
H7CqhQhZY4YUXFERI9rUgHa2FzDR1ExbER60x9TmdJ9OVikrrc2umvs/+GegqYdp
cXbqaGFCMoTnAt6xFUIV9wIPMCybjY60e7fWM+6KoPnUvS9i0p7VDE9GN703r5W8
jLxnbu/CbWaUYRq75+XHdUnVpVPOEMeM0Q0jqN6hvBBdapkqufNNE5deWSyQCETL
8j1ib88BQBICGA6J+CYt87WtfBhjHL/PvSRvo8P9k/Nfim0oNscTNvT80qtsiauz
9XbZ+U3dmPdgp/2uM8jmj2R9ze1IVrcPsI3zU2fDurCkpGTD53d8aFKd8v1O3Bs8
0lSnhF373FLL1QHSiaPX1GlYU2prPo2cD2lfhVyIDpLogDzlov9HM0I/wkoYqtiP
yDqVOO9Jo1PfywAkpK9tkTkSGxpNInsOs0S10HQx81SSKx8tdIsLUpSNsLEMVNod
o5w8dVwBYspgxBpW5BBYq8xASphl+ARjALoHM1oYyjtjpYScllAbN1+k+fnP1v8Y
rR0CQd1NU3nHCNVYBNUOTo7Jxhk/dm+3fAoahZjxrfpla0CJChw6EHiEU1qbpVbh
2AiyO7B2qjRURogiuKIMguYNXTOrvy+XCTOnzxlTmzE+5c/H4eE19ScX5BzyIaOQ
SrHd44Hu7RtrRg1cWkFRJmr5qFspIsk1YBTytZfEwsPeFA3Sg3ocn9aeZnREjUzd
RLGkRKvvC8U9ZxIiVEfXpHCzmE48Ri3tIKt/P8C5XWFCXjbrSLyjATK4GvUi0iNX
NPXGJ3c5ycsgA/3jDmcyK5BvzidKDen1VIvDChQ0Wsn2xgNfsLPBgY7j92Qj55bw
L9Wpy5KcupFJyZx0smUyr5r3D42oFsa5afR/tJzP3N5jGRxwYXW3i3NfKKw34eiZ
YeoZKzqeJm/hgy9M9eETdJGKvgMffPhr+J9EqWaJ/ub9e2R6WNEkAaV6DbbSYYUi
0tWjX0mtODwPefGxyq0guOG/HX2Ka4IRzrb7eEog36P/QR1083CU4KNjaUiosTCR
Xj9y+V4KQBKV/fZyoK0rRrUPtITEUkzvvB6wDjQzzsFzPvBMJ2Jm73OcG4FQ3kvv
HUAYY5pCyngLhTTwbPlJ5mVzXaUIMZP54vQhDsdbXglxjJdFE88fK1dg7fJSLRcq
sMDZwriZvPSJ+TOHmc6Znt6e9TRG7Z9E0TkJz/MLWK3ERYd/8vwTBBDH7Kql+3kN
wpBd89Bj0kUrVQfXpM02FD7wW86VoDdgmRyugfEqIlvQq7m8fZOE+FCaEJNosJf/
uO/DExb0OiAILQmSSGOy61OfL1xih3EsEbjDWVLQlkXeHXJd/zrjjhFDgxw8iHlu
++1fL63npZBX53BCodG40SdlGwT6I1wXS3kE/+q4O04VVorF54Bvdf3erpIGGxjC
1mXhOXFN7Ewc4T9/V279idnqtUGPAQg8th0odZWWgeMp1pqC9OLzLLGpaeFl0jy0
U93/TP5P9OT1PhPmLP0FSvLS78osBMwCnh90ZoyG0qiXS8dn6xLVbu5SBENRm5fU
Ne5z6KvgTotGoYSIppsQB0Pb/upJz4i1KCA37e4z4rmB1ZmrbWpjSvuuX4yloRMa
bMQaD1DJaeVRiDq7pB2O+4YB7dnGujh5ewhPguvSPSfanNW+4NWFNxXJDPsloN4Z
U6fWT+hGqZNa3u3BDs/uO2Q1g6lVkzWVaJj1STqsDmVkla14/vAZZugByJ/omjZj
P4rI4uxA9cJsE5hT0WDtgrXJchJK0fO4WPyNuTdbTHV71rfSFxpGbU6F7+hCZC6P
xa1G6fItGBvauzzJ17ezg+Z5wI9H81cIgnu/cOfuEWWstf/221IPes1u657od23m
ZPlgSBvwEWjHQqQ3+yM18m9Hd1TGLGPZ34PzQL9tcDdbHybmEiFjZk/djc47NvIV
3XysRmF44UOfaZQ/DuYpvpqNQonVTNq77SxscWRRhYirdNpbU6GBpZo2xyMgAoiI
IFLXfatisKTs5Dt74Ta6e41yLyCjSssKYvb8iHgRPTto0z1uT5EEFdm2W1i9+BaP
sUi2XBC+Uv3nJnjbt2I7eiXEkFzAdO6EgWNLqobTXKTfHNLqg4PFOYYRsiLHMcLw
sjyW9BQFEF8TXMy3XykgjRCe7xW4OumIPfL1xWIgQkh0Hj32TC0EUoNt8+YdkHCV
JBd1mPKTnjagDMAbBy5fv2P1q5v/pPgZ/Jveyb8t2teRWnZiM/1pCLw3Ob7SqWq5
LdqeRRcoY3sV0ENofLJbIi+zyaLRHE4eUQQl2kvbsQ02NU5JaT5HYfxNpEfSYiCZ
qFUspHQ+xf5KmF2Zo16XpltJ9Y2EgmAoln6aK0MjOtmILSskXrqVeQqabuaSa2e2
QZeupkPGTDsaPRxv9XsodLQ3yT9JLAH2S866e14UFnxT7HvWzgVbIwtGrBAPuV9I
t6BLylRnm6n9UZ79AIuTQkmunrzGoWbMyKQOA9iQCrCt7niZtzIJHHbtz97/azgn
zQkYvBUNELr7uvmAIKT77p9JJwad/opPoImN1r3/SQRQYupvs5J0RI+bgjyqB5pv
A7QzCmoq9qSBnb3j5SXMHlZ1wrdPkJ7MoYuWe0iPg4hrrF1JXxYKKYk1m5M/Cuvm
b9LvSpuxfNrq9cC0VDGmMRI0bQmrWQCL9FFBOeOSFQSCEAU5xheIkb0VrRDykXHI
zVP5yusG2IBun8sE0k1i3B51yCNb97YxhOw6QNNrVNSGEIhUHoa8SyNk+C6i7iKy
1/TQAvKt3iSO1djaJP4olUDPyz3ElLpEATtUR/rgC/4+N3v19GYTe6CFOs18+kXk
WpPfhugX89l3qCWDvPghK4RbLVWLmgwkrqPiiTdvziJtibdFZCIWvyR1MsTgbke8
6TIDy+0IcUTA+2xxKuxHk7OzLBi/WZ8hm6Ht6GEjoly78t5VtmV8LQ4nI/9cwXI2
q6tiQEiLSAt6gUwWwsX742Q2Ef5Cp6sVSEZ4NQyZ5pMttqib5qpty4+2AuWONlBk
pkK1BJdz4mnQVXgNSqewvO7IDtrGIA2yA4dhhKjIfdio4w/nURJb+syume3EiCnz
PM+7Zatt71SGpOwjL5uaitlh7zB8nn/yxnBSmUKsa4PcuExnmSVfFN3nqROxG5rl
DsEYmlFxl6FYvYeeCzryrf3sR9pRbvTkt2WKF6M6cnGk9QxhLGl8BooG/X7365qg
8WW0KPy/8Bf2xMkA/c8ciqMYNQJfgh3Q++JrK2DFic6HiVPcwAdNP2j1EernH0P9
DWaH4uVcas4falGxZ1fqJrEUbxYopJ9yFc1e1oxyonW7qDOOTl6m7TvwiQ6eF4OW
KqmHVu3s3siae9T1lFJqZPW4HBy5tV4dJWBqcd4NgKOLpO9JoAFGJGOGXH8dRlbp
lghxvbeGYmfFdotVgZK7BjxWna4Y52c/WcqgMSCRpO9VevxI5cbSxbl9FV8S+x69
64shl86SFpaQIJTePud5YeXR/dOwEHk2bqf/vAwSS5M3zMttNZOxioh9wxm+3QUn
j6bArYji9o9LxJo9li5He9q07S+DgwOo+dLjRPTzI9Uy8vVBhTJqKESOMf58UBDL
6/s/OAv5O9/LqjU67uLA5MDVLw1TP0YUpHhoHeGLh6vk9GCHJGGPEKJxrhDPgBk8
gPQCNFlFzQVm5XNejeept+c1q0ShJ+GqmqU53olVDcJB1WFJIz3Ilkzu1pBhO3QZ
NZOwQN5XsXiBqWN3s38Kv6EcFzPLXuchv3XQP3/cOcQWNDIVBZAwn5UE2cJtOdm2
O71/kv3Nu8F4ZZ3DrC7hNzodBNYGdRolfQWtXQfw3Xc5IaTqF+5DUMTZM/11+EPW
usTRZascYJYo8N2jEmJAQHvZUExCjd1soi00oh0KCMzDjmjuncwiZsYOvT7npfgQ
d8QtbvKopBLEdB6tH6wW/B4X7JDPWvGcUO8XJ0Pb5OGnRwowHoUVNkw+69KXxdSW
5KLGDNxiEUvHXc20ZDC4CKe1S4hofDEMrw9RqeRVu9WwSrj/D8qceZRVePEKtY8j
RHKm4kpDDxrwwf+hN94LzgLjyLnmZW7oFTUe3jwY3uYtRTQ1Di0wdOUZnbnLc8Ux
qmfz3eKVHmqCzB0Lu3NqyJS1BBHFBjiEO61IGoTVSiTYEThMqBJxOXuoo6xvp/f9
wBZqpCYYMKdsTREuOc3uMLl6bE5lrJk/mPVJju1D+6LLu4dfmUp8NU3tPcDJOU/t
6W/Frgb5XMBFKhEO9L/C49bT8pVlcdqmprcs17jn7cEWtgZv5NH99xLbP0iz44sc
EpqKrBHgS/xYbfjA7lBxiSF8WiDAF9yLRumT5mKya0EnozHDLzg5gKOthJhJjgdD
jDHKPtrlO9WaXYImB45nCkvSv5h4JUDlXOl2FSsy6Gl8onwuvgFyuu6akyAt07Az
8/jSwp2FTbakY+xWP7lQGhyS2pwXZmtXCrQJSNcXT3DyN7O1TQ3kM2Ohob3XTvaD
+k3PtabXtUSDT5bFeP/K4trtmS+F72tlcmDWDYUAZlg1u/TP0lV8kcUItQoU9NZw
STCY+cuSU0zE57NaOrdTXVIOOEUnIVam4Yq472WDdTuwxy86tG4nBDuebPOuI/55
8dySv1UjoAoS2GI5kXmr2TOp/kjtKJWNgGEviHSqjO+2QIh7DEPhg/S9JS854aWy
1MJgipJWps+xkjU5Dj0TU5ktFF9cG7tszfWoqDvsal1np/L2tskxb1Dv7plL1qll
GBZD54ZfiXBGNRpxeWbctF3gz2WoreDMxqJl+V6PkJlwQIYglLn+zAPbJIL4C6YK
M+Yr4aPwpQ7qMJBmdwEXBSoXguqABJsmlbN7zvM/buSuyLU5Vx6q3HeE+vB8vVwL
/BZBsz4rMLqNlcqAy1LrusAa/WDzINMR71O9JSe/Ktd+CW/714c5AtwWFDdxy2Ug
J2FdqH2yahpQPlFtySMpmFV5H8tcSulQVJOVIxBPMyRTBO2iQx0tuYAjdEtoXktV
SDRhTWpvbk5iRHPLTJ7+CqvluiXKDArEhrf3829OCzQbsOKerrhBABiVe5/19Xn0
s09zt/V8ZeSVuD0w1IiLLlve4lK4lxadHAAot8KLwVmk7tLuULXvVngiDZOv5opQ
8IHrt+gP3wAk+z8MASxhbVm5GYn/duSgcg4H7jYm6COfNhqu3BphDNrSybYtQsLp
2xupu6jdmAh1p74NCP2dWXb/apqZISZwCu+RjbWVSEUvTm7s4jTixbPL0S40kt2l
tJ5wq+JT3IlXMY/lkHcJIhSy+UOO0bK1KJu5FVW4ACWsmJh798/0wRdYq5QpnaRl
OdcMvDt8UuqObTe6q8VC77/PdfW0phj2DE2COvH8rgwwcMOaDz+OQ+RrERVeXDZm
xGqUbvoN0ej1Ihone5UaKgHwHN1i4gI5jBXH0bFpwfm+arS12emurervug6m5Rcl
nX0wtZYf7UZUCujoyB+pELAyw2YsoLMvhujFuRz2J+0Nk2lQAir5Xk1FO4LaAbh/
mcmhTZGHKkGoDsBk8MLcNhD45Xq2x9/g0237xBlm6YdMSyScZe7oGkKbkQzlHKWr
Q0ggN0bb06DpC7WZKGayQy5NNaXbGsgflG1QDC1ouXiN0xj5ym60XwqD73FQ3AnT
dk7d1NJoxVDD31gdsOkSga04feL68lpqb+hBSiVRWXn7V+ddz1KON29wKn4rOTbS
6bD87cHUUQmGDAjod2BxUAR9Kvj8MojS17oNNaMjwxsmUTYzUWGGWjjBG3VFvXO6
5dEaaJUl7VlInaAL3MgiDgBNkcuifTgIOjsqDEbBtLML/oHR2qhsBuarodeYeh41
JKkadQJnouoxtUsi/z85wZ26OXIYsPqS7OKRNg2PqT/BlYubkzGBJTxW8OlnVsgq
J4SIlWaAspp8g3tU8OvcGGPKYRHlcWIl0/S8HL+GA+x0GviMSpicHHftD+uvqsQY
vP3CEl3hrI1w3YRDHJ+EE+AJNZ3Ti2wb387ZgXGufisPTGo/X5KLXOUv/Yh+TuZQ
52d8LwYdVFUa5PJfSKhaZXCZH/NX7vv3SuZYKQh6OWOIdZNl2AK5cUEgWMNvOdbP
ZPbQu/UoYcfEhsKlAeZWJFjuCnR6cTF+IadRVzC+/pTqMOg5l4s+BWlKuEwQItz8
W+qCJlRMiYZmB/IwtMqUyrHb8Rs61F2BwKXi4L+3gKW2cJ9RnoaM/DVIb3ASVUZR
9VpzKykwWrboCAerFr1tNkov+eA87mKB3RY6HWl7WthW6ah+xoPBcNlQ45vSX1W3
HOIVyu9NBe2TA4HiwKuq3k8LUXbujqFR5epx+QABCJDHG9ig7HZXoy/paAsI8jDO
jZbBOKb2c1mLWEbINBK4PrxcmjT872hg6+Cddjolhoa56jI9AOO1aUQUrPJ6eeWi
Hd0f/j8Z/hB/l47PrTew/V2piGqXVAOlJErMoHjsTmqNpsbJmmlzXRRlPRa8LxY7
jfZ03U3Vv0hVVpr2hWEjxFA6oKMSHMoBvamrHNN0Finr1bDxM9q8x17Sm12U3A/c
gk2NrfQwb8yG8qAhmFG2vzkKnvsjHzK/O92IwvosNol8H9pD6mnuJmU/YwgIcG2O
aWFUkmWoZd+6RKOfK2NmMdxhsSCOJUvH4NtK9uj6V9RqBDeUzCEimbzx/lX+HtBf
ofBTavRaTLYuQDAcx2WPr+5UVY2CGN/JunjrE9ONwEnomkqG+ZiAnWBJeHCajCS3
Dqg9OnBJaYrkAOOi3q+TGyzpw9Qda428F1yeEHNWYM5ZC7wHiVMvk6xs4XVQbKRX
Lo5L+1MnUUV/CEBQOwirgsDS34un53c2v8qQQR1sAwrZVHhv3SSdsjka0Rp4kSfW
NnpQVeTnnS03hXQxMCDfZtSShRhywKaOxJQmfkDQ6PaHbQjgrwgWgf7tbcSJi0Nf
U/G97uKd8N1wbM6qRbUenJE0VSu1pW/ZQTSD7i8GhmB2YurqeCIFEESZb+w9SL5Z
L398e7sbNLWx5CZtgS7P3oQ7dJZklzvqy1xonk/IO+XPJWo91g0Ab41wuoWw/6go
X5LPqpi2XP3Z1HhUfef5H0DNqzjnEea5EW7GxqdZfy9eednFBugim13JcFC2G48K
a0T7e1YUjUBl6y9Bi+LOLcxH8S4u1nP2mn5TjOgIisjq+96m3BALvXHH6+RsLdYJ
CK6/Oy+sOB3de7EyFdog1bKnf3NNGou1RN3/cZeAX3OC7fNThsOjChkynOJZsWs9
5wpFQu+ZF81+xa9GCW6ZfcgLz5sAf9mFNfKmkdHrKlv7GDxwkZErnSNd1DueuaSV
zQgwIMfD+ijkyoED9Li1Nl7yA/N7xVZbk7YjfliENM6xa+qwoM9ICcORvHoCbdwK
pg35s5cAAhTELkBY6PQlxxMRGPcpC6GeCbMQOOLxO+RBCWl8j32ve09YIAvXiPn+
5SRxJEWkQE8egV1f5izZZ8vVnRmQWxf8NPvkwwQw3ehJDd/YtbTqlYUGhmO0gghd
hGzaSLk88jxq/tdVWY29dfrANidjzNQhDYv0N6h+y/ZELQD9Orfauk3R3N8IZcq6
DotaGoARIqYs6X1EyW1aVwobKVQ19MgY5nOsbxrkVwY0QeWeiSVFII5M9vRxfDip
kT0XcmPItTOsDuMiZ/K/nW2bM4AKEE5uBfcTI4T4xOESWwuA145p+cdhemy21WCn
TqSoUQD+GN859ZRzus+/Glhoh67onx6k0m9W20WQ0FFs3Tcmnq7ETdiz4UdO6qhw
22r4//MNUIHeC1KTQNDgpUOVroGm+f/l9T26iXgcn3PCix1+9cp6JLZU594JcDl8
Qq0ks3VGu/OiSfSiRzN/PvZGTJOTjuSy3WoQOuWrr2qNxY8/8iTbRH4RyI3Kz2PG
SniSgPLNY0WnbnlTwSpzZqHTolP3igJ6q/eHtxON3QhN1tchodjSSjYnQu8s1z37
rF/Y95yMqwQgMr0uc/eLPMOL5PEV8hG2MW5iSpEtv967ioKYG6V6f2WxvynojSE1
kz1J2Hb2fs44hUmOCXl+NCvIMyypf8nr/aThTd0mI23Hrbr5elJB0VSJ3dR2LI7Y
nDeoYqaJmUTJXXVpLDs0e0FBjY5T0+LSBWMRrFSS6iuRCKFXvVUBuZc2/dcSQuFZ
dXSAfXNUQ4vCi9lQt2r7sqVZ1Oebt28NL3QVUQluh1S/2KhZIDoIqkxeGoHhplAX
sdKcLaK+hfovpmKRTZoo8jQ9J+EC4H6KAB5XdRBSMu/EZsMhgfy+7FQZAKZ7tkA+
6OF5qD2RUn5ov8DwWvNq43nP4Tw/c5orCtd+hH5TfA/4m+vEBKx2HHTPMAxi0SuC
NlyL5Ba1i1yuZOuyRV8eGV4bE8Vjl1OxnplLEnun7TRt54u1SR+X8ANxSylAxRAi
ZWrJNdkRrj+kMmj5wZdG5/eaJgyMcee/XgJyFfjqFGtb9T0X48eIBG+qiYviRn4I
a0pjKsfXRc4pc3VUDC+lEORf57eb9FSiRLVH8pg39roq4c9Szqf9I0UyPls4nBKB
kCffWOaTDzQYMQqLldlmQeZsfSR1fIdT7BWBPsYG+mlBJXT2c/uvb3CHOiAVe+Y6
d+b/TaOCazHda4WIBX4i/oOhmpkeMCRVMeLDHEIO7+tpv5G7F0i1v9IyVWZWkXgu
tf1HotV4/MRuaiP/6JY+OFzxAwrEoOK+M2HeML/caC/izXhue3x0w/Kq028O9lXh
aBSUOskvQRhYDSFx0zfqSqmCZiHTXDtUfyzoHEtfYvgsLRZ+Z5NKBFiY9R4b+mTX
RIVQpx1BwvCqYZ6c+trhnUJUHnjQJlcKYUon5TNHRnDaSr55+7tffTYiQS+Xurbx
t1Ng60UWoZskdJIRbCSGtHVhc3lyrGW6i/0x+Ws38CAYmyn6QLXB8Rn88kiCWVTA
krHHTJVX0WjdUxkx9KmY1ckLD7EDhqBXk6TpMWt4Yunw7dbFCNuaQxaO+P+z9S+6
KM4CIz8R6nUXWJ0PI+7lwx0DN/ZDwAIA9l+gvCUgt7rsfhbkDRiAFs3cbFu7484H
1OD1nep8nh9oPaq4O1T/i8ZMw3JQSGdvevuFrf7bLsW5vbSw0hcX0K+ERiBqawWT
zjXWK2OANEo6lFNBC6lUfI3UxzXYQoHGpaDF8h2oFhT9RToJR8tWqHtTiNuB1men
2hRfmKzgdsmKMEDSl5h3RSECaFVccvMzEbZyxxXJesZeHW7glKbjSP5eCrS12oQt
/LTsqdoy+tuEu1jrnC5TxbKdP67fV0ZfzCc5to9F2SeVlz7NIAO3B5kBnwDCGqOU
IfmoZot4FEIbO8xc8POZjN2dmbzCqOvboSl/M/y3gulkMmdVNThyoFnGKH/HdCwL
U5KntcPSt836L10oMz0KG4iFc6IcZ/IMv0hYSchOOeJBAx7ywqQ8ffpwIu7uLGBL
AM+IidEye/EC0xGOKfh8/CiNLYrmoMiXG7s2fC8Eoq1ZHpuO4y3QKVMQmhXhGL+D
sjteozBiiNToWpumy52WE6/a+Yv4gX6/pTOd0bcNYNqWNA7QHo/u/DSlqUWBacON
U/jrLDxMM0eFKxrGMY+gaKVzInsD3KMb4zm5AQO4uTcM+4tb8wZpVXyBiiYxqqWz
Cjb6aQknMAepiwOBvYsfHgp8nfw9R/boiJ67KxEoZ4LALXVKqNKectWwOOk54SeU
grYvxv2aJyGmI+52cdEjKqpR1Dw7fkWa/qVgzp8BK5DTe/SXeuxUIqKkV5azI9zp
SHt+HZjV0yKbXjS+yoYOXJ7CJs1cAndxHYAhFksev9q0UR8E4WppdfSUQuJPnCxc
PSbnpy3RGIqzBSvWcwGcnp3O7mSMbS8emm9HGWoHGc9OflRuGOS2nQ2wFV9HQz9F
uRq5Yr5frQD44Kdhh7YzpOWTvmtdg6dS1SGk97tOesoC6cMk1afkf8PZmryblM73
zrK8NputcDyLAN3f81yB3fi7Uja/t+nkpXAUZrk/hEd9F0LzSYL6KuS6541NC8n6
H/shjEBvuygw1sMYWROKFj0qNy00/NO0p3hGh4B5rbs2gjDrk312QcRy38jM6W+c
GIC/paiIeKvu6DtnIWVL5NqwokstGM+RI9eA6J5X3lMRReWs/4lHc75TAXhbVOzY
TaEeuRB3qWVttMEuWv8xPHtA1Xdwr0Dan/AJTSNNp2fjDg/klMzOqJ/8HM0EHpPy
t9QaY6C+Yvj54RHZ5QSCS9U6MkHcP6ylDIp3Lki3AOhN/BF6j9BL2LdtiY1ibPWO
OZqvMMBq+OCYeHyysVfI9eb1jj9IPFi3fLCA0iXZ3x+0EWB+CYa0wrMpXus8J3Mx
ubhzHEp6t0PAFgJxPsbT8pkRRljGb4+LOkTToNgGoMeZZhDadtu6nJnOX70UO5QK
RAD/hy/JAkRIP44tuC6MEKiInQXxAS24P8xaeQPLd2g4u2X1sKs3aMitYw6oo5eM
Zva0ZHAoUQ9cwoLY87B7xFSKamUffyayLMKhI3ym3PPcX3aAfc7J7B46+RqxnMCh
b9hM/OHreh2TfgaddwkFRaJvxn17sIzte961DC2J8xWfxBGbwZkS/PlgZ4jOXVPD
UnkgfgWqP+bhJ0/E7ZfxVy/HNZczf2fDNENaZd5dMzyYOeI/2L1g+Aw9zYtet8n/
/KB2nUGzbfrqB9JY25x0y6+jwMCuAyDio8BiVLRA/b6AjJENSyjRxfQPszpExhhe
PoKLXg/j+kXeBbs90FcjRzI5xtiQzOUZ6Wxv7SH/qDtObHc66zYCcm4zJQ5oOfjI
fRWN3LA8rs4Z9v6cZVi4Vt45se4MmKXme3FakeLS5OBbxJbH28aZOd2RMmxSiaHC
SsiLEPb1u8TeKS3+wJ5qNU1NvTOXG1blnJFNToj3RIxPVfVQotPHmC5r0mKn273U
pNeqCinCU8aNPGbp3Ij2Elh730M8MC6p+wfVyAivPNZchrxz7PbvEXdAIsFq7dfQ
G1oZij1nD1vQ30+WnVSsfzGqTIApnUAsy2evx+282lxLF64q77imjE8/vVqJUWeT
6CtIwPZ46Pn5DOCgu/vMfYsoNVPn2lFGVVo5EQWbZgMJHnCf92mJCiv/4+/UHjBm
uloYiLBpWgyeIWCCQnDMfXE7NDBOmWz8lJGVgXKdCyBr54nO5ldFY1Wcd4sO7HRp
s78ERVVt6ncKomrXqUz9IOmFalb6PpsD4sqcsbZC7OlELG/h0FfdQADWDvWaA8Zv
iJP3Zdj7LGl/dJgCpfMv27DtoYlK7Lbb0u4vuYEVtSzdHR7019FS05JZdcursQRG
FflyGs17FikUjttnNdwGChmVp9pm/glUr8j1XH9Q8u7r8FYCIpXblWQmrp132rbZ
1X0UHQCDv5FoWmfno2DAHakEoRiC5GshxV7bQ7oZIqb00HAySruH4NhVY+dSg7us
tq3mXBdiCwewL7MDcSKHsCMLLsL2KND2zxA1JsiNE8/7M3DYje0/YA7lD5VUd0ti
mKZ/nvGUFl6qdfM4QbZS29oLcPBo1+rQIUf6DmYHyCr2mJML76Lmu2Y9PuW6Ma2i
m6kX3W93VZM3QUXQixYdl0JLoQe/NG5rIBmPVgTAiFox3QvsxPqjMDHMnpEjSvRP
OzvQfGro4GpMe4xNSSOW8Ydho4nif25moBAjPxf9jQ0dHTJ+XRgY4+Z6Cpi+D2IZ
o54Xwo/yKLHfG8N7ygqPwsJM2Dc6V9JCnAicSiqVhuOhgKS80kcNNz5lZAR2pZY6
kcCdlK5X8YLKUi43qbU7WXka2APTm3H5ex9WoN5nzlyIOixtPTkduuqWUKjIMTB5
tk4kOy4+f0W2mFskyatlqPQk8sgiAYf9C4DiDSbHPdQiQL4VBJy8gqIeGXRkMlxH
8glixsqBTB0zHX07ELVMpJ7xM0iWA85ux0A5IMjQjTIQ8NP9fzMuggRGLA7kpUpY
C6F5rKCJ6aMacW96LJRT08DQfIRby5FP6aftj8o/0GbQMHJUc8pKgMfYuCEc8YXK
yhuaefKuFM5io2Ta+I5VmUUM2IIPjTvFZfuwkhHRp3Gtq06yNcSWcTRQHYlngUK2
Kpwh3fU/JDwYk7gY88SMILMWvpDsaCBUUTn0KQkfrseYU+bRC+de7LWBG3CB2FSU
rMxxHNItrYHSCgSEEDFk9APJe0jDRy+LraPyy6J6f2otbXMsOQRH4fBhvi7ImmMl
FfVN9HEUij6mvQz6bAkYdprJN94KYlfeF3c+ffEnL7y6gnyu5EH06Ks2KbDDtj5P
PxhlI1W62Bn+IEOJPeHwhm3lw5LUBx7uH6emxyMMVLxhLFv8JbHm3pXJwpt7obnO
oYnkxF2RcOdGIwwB73iS6bMMEu3pk21WLgFkAZykcMcM3tfHMJI8i+r1FR96rYvA
uXq9lkpCLF9VuUJdJNVhsCzzGetlxoFM2hgeye5dUrs57xk8sVY8N9JSlhN7BzcG
q4a6N7dJZ/5k4FCliL1yzCGuLFeTIDhKwtnD6asGAgOY5HYDvPERKMXoC3ABjL6A
CMzSzAQw463OL3ckboDR+jp69fkmD22k24+O0YVkecWmUeC0KVK6p2MBeSArb7Lw
6mFiYaILcaOxyW/zTfRQDRblCoklsEeW0lnTPKQWx8hZF0xepJNa7YbCTYIhcjYO
wTV+piSrSj72jthYYH7u87i+tacU0zfyoRqdyRenwY8gjs1CPylN2TOsu6YfCGKe
TuEOQbcso5miKi/wmElN73IA2mNKTROmapm9QHTqDseR4PcFiSy5ysV/HvGwx5Mf
RJfNaHXXvT0OCoyREUilKWGKQdJ69eZFWzgPfEM6w8KbA5ZRbYOHOrJxzoiLYRdR
nnuUvWuEuswE64E+vTjRcu/sPxL0RPK5ZURdpn2xBKMhM2Riys9pocL2R3rMpkw7
kQ2h9++D47cD0/rGhFtTDLvqA3RyJ9HkQrQbWjFX5d427ksDfDbGO40BEl5TZ2iB
3gjvEMWz+sd9dn3lskX6Im0kp/nm9STaS5AuEFvZpQnMLl2bh5/lwRnLfl8ydCXM
nvC6bpjT+/1i4gbSWvsARznWf8UpMQkpLuG/o+cMAx1CcviWiF/oEerGvYL3ncWh
FYNAILjPQLhWYKEy16NrYQULEVeSrgjvuoybxCqIqzCmK+VDHQEyCngm/hYeBZaL
iUZ2YYPHLP2HBxydjojb7m9QldkJx1BYlpWGx8O87ZjDjV1zzxyCsi3NXdpz5egN
bb4WlgpspGses8EQGAj7eRPem/oxuKh0kZGFqDIRysONGT4su7fBJe41qtEtJDfA
gsldFyfKEbynE9Z/Oj4ym1VcyKjfun+5CKMAtl09QLslVvSDlJhV5Tri6x3C+D99
z3EInrNS5oKqFS6AXsn5QI770OPSd2h2o8b65d7TWfLst5PEJEPjmLojU7tIV/zC
G/atefRtPAyu2pec3qPFAmaUBS1i2/rd+FTH3IeHbeNzLYfYGs+pKZ8Nk0LqhADn
SIWyWiEmjN2mfraqwuFpvUDtBLcjdbuNCm9nb/eFW5Smpiw7TqSsQd8DTBLULsxt
tF22rdGzlBbASHPzyuK1Eaj0thC34vg376BY59jU0nsHLCY1NGXcTT8qmo34HOM4
eViTQq9jGTu2z3CjpWpoi4NWyC8le6cIHjrePp/3Lpff+p9YQ1DFLxt37QP/8Zau
GkQGKlDzWkyFaEiqJ0dE0oTOfcKW+iyBdhrDHi5q8Z04qjfs0doW5vcnHaKrCmWh
oSWs+IAOEXwGzSrL6CFdzSXltpuaJO0eI6sQ29TOFrbSRWHoIkF/+gGT6qhHRnZj
86eS1hf9u+3/OSPIAonVoFT42ZQo1BzzYi2of0OXT6dtlXdoOcnybZkqaLbkoU3H
Ab2x59+YSYjT9a50hVvmhKqlcypwqkDb5MEUh01sSsh3g8paIAKuLfBFryivg8UP
nC0V56wnZV3yxCy3aDrrJ1FiEE6AQlJSQseSBzNpb5O2+R3JOhR47NkaSkr2+9Z6
km4Fa4NJgdm7yFJdtifRSrmz4oas1iPvuOeiZA5oSncDMzYmXMXM6c8xbUDmDSg1
Paq2I8tdYayhCipik9IK7mTcYdLydqXOTaxN11JLFiG42s4Y7e3UACMrsd64mPiS
gy7oiDdQF2SzyZtOXGXvm5Ica8ofpvTQ7ruCNk/SuOqx84ca7zIHhYbMuUr7+X4R
mPSUXrjgZIzVk89WCWZjGE+zzsDW/MJG3GeG1tx970sJ/RpCsePLtF1CJHb0sGol
1AYyXdbOIzm+oFQvw5PpbxTdwllxvcr4pZPDf7PVAs+QXLPw25R/ftGoTm7FxsTj
nzQ3fQOiANt5LAAIPU891ea0/0Yqr5XZfG6/9369TTjj0GSmJNfzfVB2vRxSWEi8
jaTZNYxpfFLRptKXYVQXv/vpQjVHGMvIVivl80CJxK7wRj8uMCl0yFyfxNj85x8T
iR5/ksKHOV3YkKDKEVAyiqMh+MobKas2vzeREr+b++O6jLQiypruaGf66pTuDXUi
b5GzVKQ5gI/xSuQXqJlPNCIqmS14X8udKx20Y6DSh5f/2DeD3Pf+n2dhMg6EipNe
qZ5/SKgLWI34HKQi2CvgvvBY5m0WCQW1CxwcELUsGsjznieNgzVnmWjfp3GVu926
naVxGs79n5BqFvX2FgBbsugSI5zMppsg4yi6AB4HiccD1di1QA+N5AgtBcf99gdh
5KelpWvbsMYCrLeiqjU52hLrjZbKM5cZXq4MxR1xyhquvEQ99HFsgx+2aaELQBSw
xsoGkX0QfFAITxJwbLmxINuq5/RzN0IsqRNbIR8R3et+RVkK3acrSMzas4UhItE/
WRFvMC8v+HYoSOk3pwJRxFcqCv0EJbrypC1bzJxwR4B0w5bmYvMGAxZQjSSfTkiC
pZjeYWpzTRZtVmbF34zoyrnnzF2/0iMBRhbNdJG8h4dlV+5XtTIZcpsDlVEAIGbH
QbZp0ZvCW0L3ajU0uRNlrNubHiYlrRWfqWozAuzZL6jdhRDcnb8E8cmQ4mwyO+Uy
w0zHMVs+Gh91W7OYk/5kbg/iEZXN6oSNn3LV6N6eic0bxQ3rBnC7CSmMVDv17VtQ
nOXszgOaaVZcNk1lBpRMwV9JB2dEFogkQB6cg6hKjw+XcQpw0Sj/zw2SKEBw6zKA
eRyNi17Tcrxtu7OVtEJJEETF6Vlw2IPZK8au6laLc5VQVNyto2pvOfNoGyJciq6r
ODI22v+lGcvTy9VXVoBbb5OZW7P/epK32xMohKExxksnnEoEFgw8grPl4BFmwuN4
u/TckSDcSqpoVT5hB7vmazonVcQx6q5uC5J1LJQk+gagsZHJdbW+Y/IWBoiFLg+Z
Uo3y/+uHaY8yYVINGjKV4nwB0WiD8/DMqbir1ZxvO7gkG1c/q1zt0QLp8rhrBbp2
u3grew8IGD1r6vsQBNnS+70XnW1mtEwksIUnTqKSxXcdgf6Mg31lk1hE+gM7tO+3
Eyl5bIRInPP/PHGPz67fWnBCUMjdRyA5sWCs6pfRO0ak11mSmw0NcOWXpOmGgUFW
7d0V1aq3qrwUQjZkm3HWr/OGOpR/MdyfUF8YZEtXFOlFNSoQUmDtHRmhSPVhl5NE
HuOso10V6Ojf7zeTLmHAAtD0sNBHpx9X0+sCR0wD3XSA3wrNO68Wb+d8r8BIjfq5
s9hu4DLgC8x2BonAfshe/6rC8wMquJFyTH2BN5fq10CYWbSwXc8V0685PUAzidp6
V1clOFey3sVPOIsQ6SdV3Yr3U0KnQLbJ5b2UI+q1hGPJ+IgeB/dacChtPZsp3dvi
+TPXurIPO4sNd3N/t8znMVKu6lzjIeUQkigyWQdMTxUrBrqSabgSRqnZ6OX9p+iO
fE4qlmWHyt/0tde3gIHg+cLuEgp6MMznF8/3LW8lo2Pd/g5o5gG1iXk9F6kntHPt
dxXB6TNbxyfxCFz8i02Y4v8h4TXRrOFx7FwVUfkDfmfaJdRuIemMh9oIU08ZSR+C
HfGIKhEQArzxQB4mwmpkTKWfxPILJOY5CtJSGoEsxxYmx4XIcpwk3hAAEWGL1WrW
k8eB3HSAZ1vwGbgV5SKBm0EjV8nJKLe2WkeShks2PK6lCb54B3TqmacZP42OVxnF
XgUNz1oaIY2DIATxw4AXOO7ch9HWNMBYLZg3usaYrNk30XeBaqRN7rpZbo8TTm1o
SSKZTLEuVmAGExKwurI6Vd1oJZafDfjIYIWZMrOiMqEuarb7554v9iOIcXYhFh4F
cBuey3bvRchWuzsAOIXrn6alkUPV5I8Sa1n8Lu9oGskzLKSs1NKttZbG3YcvyEjh
eGiKhKqkuarZVCckYUduZ6v/9NdGRqe316CDQS4lgVkN9Bi+LIYOHcxjJ45pkKV4
mYE6VgvJLSM5CqwA6kUpiZHb1qxM+1yISBW4Q7K/XJAbQuqcoaXn9n1GyF9oI4E0
PeQ7qCaQIWpFQB00IPygq5cmCfsBpNer8ve6oQPYea2VFXT0p99G7krCidgDNGi7
DrqB4xhVl0Z090+wUv8MUd5TxG9DA0RPfDADlE4wzr6vOt82c7I2/vWkGpYtlraL
ljZy0V7cLOQ6Chojj7XzSy5/VwZ650hwu0YgzxekFVjLE4f4O02WrrcwxyTy388k
oCpAwrdigOAmFcjptpUDSfKHN51hvRIkCcDO/o9/JshsnhfrtsdJDqEsppDrfvsZ
tyGnDJ1c+wEyZxHWlBWlya1T3SdUyxxsMSMIBsIKiTmOAgi3qY95r3vbddl7MQsl
fk+WBj2F5NwNNg5dSqoJ3ZuIyhtyKjz5a0ly0xT7z0CpPJON5mU10QpQc9E66O5z
0ylMHLtGbhjupt0T66l1klxVJAD7OGMJ2KF0UzXquvdBTtG1XIUFTZpJQ82i8mT0
sOOEB+NpzNRFH9sRip89imeARRW+HEPC5Ke81JeDpwXaZ+VBbG4I1gBdwi4G1chD
OqZbZA2LRC+0QRLyWvoNEq22cO3OBlFsiUZodHfaCzXdl7C6tUSqjPImW4VTX4SN
v9XEWB9k1ozlWJxrPeDpge00Zdz+yzVY9hGcqRKEM7yMR7Ng6VSJLbvEKhIbhisQ
BfmcXherGGEhH7EQowC341m6kAOoKmtWKdXXoTABr0BD1tDzpl3uriFG8WaBUqBR
oNiqnj3Ejtu/MXLKugUHdzSW2McIhN6pVrnrStj76Qk8l1+N6AP4F03QyoFloEoU
X0TieFbi6HjsBj4qVEttu8k+WJMO+Itm7Rut66RRH558av9D8X4UUr86wuRRitJ5
gJcV1fSLQ9GYGXGDFeRrVl6i7SnjdNSneoUroynNaaYahfjYyDFdEyGE/9HH1q77
ELk4eYB41xD40jpVVFDXhN90cu6mtqNy3N/0Gp7IAhZhi4QFbhmtemH3tPRbtw8K
OVXKn1jUuwRDmHmF8q4nwLMgk6+7CrMtHrt+DfqZ+p14AoqK6qrI4KObWZot4DmS
xxmocjj9QgzcBbZnMq6xrh5Q/rxBwEuY185WGpImkD8dRV9gj+jL9l1/ofLC/Bdu
YF0xfQKfBQUz8q8W60jzu9QSQzCPVNfqm040Vej5r6beLA4D/7zBhYMdrF5WiA7J
FXEwqke/UL4z075onf54yYhoSGGLZdmfB2FGT0pIrcSaOiByI6g3+++/tuyf6c+U
aHDhFuG7HyMSF8CPZa2JaP6rZR2W1owA07YfgS0epuEguTljL3mc9RQRNPveNUnx
shTT/ZsVbdZRns8d8vX+vbefOM+COmgycp4mgKiS7tuYH+dyRR/4m5A/lHunV4iW
yLGZ3EPZioO3JVMQrvRUTB71SQDNKVCIkd2gBqkE0rSUwUupLnKhUrmC+TkTQY8n
hJgssrwObkvrGIi2vyLY7YV/AZWLbc4x1CNKgQBubE6Ugt6THt2ooncgJ5eMoEz4
iuOWAVDa9igVoAHC527Cnaz7ktDTJxUFzgaFdni8s/HuFnbsVjJstE2ESuE+tHUR
m+GNOu33TVf7598J/wI9D82/oS8DcuUZSUwcjKWHKkdthfS7X6QIv3dUdUao8SsT
7x42D4oA7CKyO6CFMYPgrJVhH4Xs8a1UdKD+jjt5XSoY9x6a9QAyj5cZRaiMy/QA
KwnGjD556hbNYAvTMqWwPQO3I5E8y0zeK09sPK17E90DEr7uFU45ZCc/aaqwMSOL
U418L14nke6A7ldxbkhTr9APMrO9kxMhc6PxqhaDWDcqnZbUi2C4D+UgrnfnZeqI
Zh8SWmC1w0BAIbsD4Yv++DZoaSqLb4nE2bP0XLsqhhzMbg704zda3IO1npCCHIg0
rgeJlDP5DTvqdwiezcbTQEON0zx/fnNxoMjrzR4Pfz/TANnqXTttNbv8owhGvVO9
Dwx5c1KzFF5YsC2toC/+zZ+Ub2b/VZA4oHivG+v3w0uCESAIvnp13lTVj9I8n68w
gPI5Niz5146AxBL7QNpf25xhno/wRwb9mPLjTLosdlHoNsCIpYdAE/Wn+hdyFqZH
6RrwWYqmAVKEsBswh3aO6XLia3hcCZL2I9ZGeC4Rq5V3nBdWC17Z+HJfprLF1G3c
8/HFBeMvudt3zXunznP2MQieMA7hnjN4zjFsRUctst2Hrkbaz5RFbBbXJ45IBslu
RRpbtsuuwGshvJq3NTny7J0Guz/rc7N6niQ1fSUWHowkzWgK5ifSULAp3JwaCtNa
AshvdJGViRno19NLPjPzhNUpf3M7lD8l1xaBwTJwaFKmJ9ZDZVh+QALIk5kRsYko
hEAsuBAojyhR9GMNmLBNhnXRhT2yfB70X9Hporamh60yUHFSQd9Tc3oyWLuI7v9P
zhQI9u0YXnZN16K7sC+0UsCnqLWa7z2L4YnxJm05mMcrLpVDPERUaOu04opeYDjT
NHLmy2pbfa0zGQiTf4NcT2UPfyuBS3Fd1RMuvEbWfgmcMUH3hAAfW0UOBKeCoHvA
P5gwvDX19kBLB7ejiAwwGuOCb0+JERahQYsslp6Mr7nPUxLgxRyCxh4PD3I0+76Y
b9Vko5cVH3LSzYgS1DxuA52zDgH32eqXT67lxWgKsroIz+j595l4NLfx7PX7om+l
HLL8JxxSKdrQQWreUr67teFYUhvG0g5Cp4P9Zh0vp9notA6qI6ymnvuJmLFD3cYH
yxZbWCvTtxs+zi2IN9W+nqT1T3ct0W25BokhZcsBouyNCJ/C2chpEGgnwHnMy+MT
OycOOcn8hjQSH/R1Mr/D9rXfz083OkQfHv1rxxEigcXQ8sXbUaY8Nb5QfJ/Xu29v
M2d6vh3ey0JAUBwnc1FDNaeeuJLN756NqGqbrqDXuTRAS5ycGTqtMOBBGPae5FeR
3ZwZWZaAI9TP0Mes9b4HKe0gWS7lrfdUzNXd2gVsEx/eZGrD1EvgKW2P6CAYj47i
XxJcCh05fp3STkxVYW2OoeJmHEB9D3zdkbo/ak0IqXEdoH8Q/iW0KneBEX2DvF64
oRPZwgAov+g5THzEfr95GojXnEDnSjRIdLrzhXAPeYaU9zp3d/4aICK6QjiujhfU
0/mGZ8Bs+XN0k0LnlCczmRl+vaLvw0VwUjKUOdWlTPNNTuE46Po6OCEWvtSw7Zm4
3vtS48eB8zZF0ssPgytyhA7RCHy+tXJMv9HymSMMQ3F0w02LaHPMxsST7PvYipqe
qHOOhg1Yavkq4mCgFaP5PtoLcMiBasaaN2xUOGvgRiZF9CjwfyockIE3QPscTGHG
ZKPlAFYT7mKBKA5HWasfb7ye5H7BAbdJ94C6Vl1DRlFmOMoMv2EtR2RQL8BE3PMw
Yp9bg1+UqcaFO0qOSXEy4/lP5qUnfz7My4F86CzVI2wUtxKgBK4THEuZ2eNg1GeT
aq6fOIvSGYpuAjfIqkwcl8NIJcd5vINj2maoV37v6OgoEOOJJk6g66R+hAkvpw5b
Bn9m5j7tYxzqu1D4/X+rrqkEc6QSHLFeWPWdXaMDFg2RaKT3srw+BcTLjrcNtkpS
Qx+g+0d1l7UDKy/rq25BBE1yJZqNEjfyqBk4UBIrMnw4dFA9ZHBio5PcsylN622H
xbzPV4SXK3BkMRoFnRTZU7p6l9w/puaPeSpjJ7i7q7UTyYJPrhkdOU4dmXYrmTe2
mAktRr/wpCdIdKP685RAA2491/gVY/YIlWOWv5DWOGI7bR4GpKrwbV/MVandV1Qq
R4T9Ro+6IUywnWhdNZkYYFY2z15ttkl/9CYLMgOAIzqNAZH0P54IJIPQasS5D1eh
SmUUJhT6Z8XZaopOBfd2q7vLfQ94L1s/v5Beu0tpSgYe4W6dw4yFZfSiuVAUDm0D
4OXQM4J7hk47J8dnfiXVTfIJJT0Z7rsqX1N0EW/w1iVA21UENn1xW8+0avseklf4
Oiq9lm9lefIW/DYMDJiuQphena0Lgj5U+q2HtoEuKFkOsq+4QF5/X3CmiBPTaauF
JGA8gm4OR8KbBKWPlTvsrvn+RywSeFoPWnDizVPyOD3EPmk+nVAXde2b084E/Hni
8NWRAFU/dbCoC1zBTIPiAlQTmgwj0+0WobuSQaGFunt6u8efhWnz3Cxcg+0+Ef/Y
8TmzJJIVrpvaJMdx+Cozoh7fta/mV+obpHiQ1uHYzH8/Yt5sLK0wD4BPyBqnr/MI
MchuXoKaziWLKsYmhJSFIjrMN13RluIaeunm92k+6+JBlpAcPFAqM7g5SiqcPu8k
xIF8ECSNqVyLnJp1LikoUgFNMTHExzsZFCznph+PbbKqT7fMfmW66GO/M16QXLRP
FavgVYt/ttqTNBxOz+H8BT3sHLVunuJXTzAbLjGFRNIt+S2WtlxOuliaCag3tIZ1
JO7SbnLhh8+GUqQxoRi/krH+xrDtGLOZqVaDR1wugJixjAUQFpWZODKpRWW5dbsH
na2yKsDTINpTZSEWKzqQudePzbrrfyc2Dcfc5hNIX4rGDnlhcn59k5vLvDKZfiJ/
49rJ3vEutqGALn+lidk7RQ8pqyf8LZpG09AwQSs5/mp9O+RWJfTXlgyNWNWynuA1
kmb9QDnUYthJJt8BIF68q7pxINpShwhw6S68u2ufLUm0Btocwfi/n9/KNi3vjOhl
8TT9vjTZwItcrgzKr8csvAtNzSouik+HZQcmTznAHJ8nIvyEdEXxhQC4gkbDp4MN
9j53kyPbjq1yRPKo1xMFEX1l57k8vnNe9d3iT9m/Ya0hYll5hdgzXnFy0K9JYOfY
twsRBVhWzh5d68j0kM4AqTl7FWWzk81P2GMcXyRERlV/cBfDPZtoW1qok6jJ6qyS
gS6rLbs26X9vXZofgzMUtE7gyqFD0hBWC97wNBnLy6NDJShlhG73GBpxqZ3hduEL
6j8ARPsERhSXPvJvd0op+jSIsJO1GBFMoDKa6F/dYoEcE/xO5Eg/gnbTZ9N3nwpL
DI/rFQLGqTLGSNDQjQc5qKvGXph3o0QOjqaZmPduQefC+BiKASnj2S3tzj9GXnyA
iWOSJV1hPLbfBYX0eG3OqiJT11NVhX9iYNj6z6tSbxoTp9Mex1obh1aAy0HyRHH0
AQ/kBLwubTFXgu9zNdzb4QvPNuHOmVWIC1fltCfPjBNTlZv96HAottb7z0u2MRue
myWDGUoDyv7U3bzhF/bm7Mcqd0S+0YkGKeMM6bW6/1hYjFIeehLGLOwXQN3HvC/2
8ZO1b+k5lATodmwdV3Ycvteb+ENEe+9kab2TmWotWM7FaIfvs1G5LKe79B1C3ob0
wi+E0HL/lD8w4EyWlvAN6qdHB72+stN/oVBgKVSmh2PuPoUWyuYstjsxdyoKI2ym
Q2acxO3dTKxrUuJzyWnEWkysteTds46xj2CCuWoCPAMu7Qh0rRbxzm7TEOv5F62E
fKESAn2W8Bmc3ecBLnyJGNt5ceHCidzvfT/MyiqfAkb6ZAGx5wCtllsk6xbW8uoS
4nFO5LYJIeqk9b4H/vifLQGza3kLbp2XI3odS9ficSele7UvuNvfotbumobE0IpT
C2fv33jbOo8d8yujf2F6ECuqHB8YO/WUME2BFzvbmnAS4Xmfr1MFo2ep5sJNsW13
El4sctQhoOx9ZW6ZEEIk160kVo5QeXyWNx163LQ7SGIPT4mH2IAFtzwgJ559l5hK
hSKs/UpeobOm0dzlc6OXHHfM2TxT8Inmq0A5I9jnTA4cuj0aorPPbKU1sP92lHol
nOZh5xVGRSNeYxot3DtpkolwGLMrR0oj9hl6J454iXWspxT9yTZFIszOQXXQO8bE
1nK7xal1n+XKGzW/Wj77HH0vemvGFekZ/vaYYLFEcsFRi/7OXvHr/iziezMOzA+Y
DA86e+4A4o2PSWAUc/009bufTwqTtNYWH5URxNqz3t0ldSFOh6ZBytigNM5KAQP3
ejzOpBI6RCn3K/vhVforGoIOpaNC6asIYjV3QJ8RCy6UhoWQLQj9BGDxyquE2bfR
ZhUDDo726ggy1XFcrK93fHojd+s6EAdnXF+Owqjaq8CRPsKqvr1R9n0kmrGCXZ9n
wAH5+TaFN+dTlMLf7FEAQ50ssB96VCd2waFLh6JKwdJGnODkGb5q+85cr+e7rTCE
1kM/FS85cgWxAqfEKzwGTSH6ObvjsFMU7oh8gSbSKv8HJZHuCHEHvOvY8yn//fWk
PUeR1Km724whJ5saHeEjowibwfkvM0diICAIBmr0rW0jH413fPpWttMaZZ2UMgTL
FPKMO2DndrrZsjkk2qbP/jA8m0hh6lynn6u98UVuqOYK9CObONdsID/fC++UNQKC
lUVxuBEUwxp0ewUCX9qrERS4xq8RGJMWjCQfXzFE5kiDsTlYtUe/MlE6kR0QDtiT
u37PWqVvpzyqOUDN/A0JV7p1zmPZjIK53PgzI/KOgWtGreH8aHaF0z5VHt3Myl1E
nwqzFcPaZQw3w4DMThC+LFGT6e0RKVPXUCwMaZ8aBZYZ5WV/gNojCrx/kE4nCedB
jf8ccouJPUPEoikiy34xD8m5I3SG849TYcE+sG84qPgjGaAyAJWLTRJ1vZiPkWcD
URFrqYhV7c5vaJAFbekGrQLJP55AyVmTO1tWkh1PwAPNAkVM5ofcVSXKcuHIfIgs
iQxkfMhOk9kzXegZWtiOi+miLsnJcaLzuSTeFhvegrLVgpsJIxgCDVsebZzEIfDj
fcP6WF7DHyWkPuhE1grdm60B1RhcxxjVwp8xYgLNAqp6ITg7JP+rRTaYCPi5avT3
ICK8Y7gwwvquMrm1s/bZE3LzuCkSCPQH1DKzIbS9lnFazQeFqs/B6Ii6Ahjm1PuL
5spGmgysm9b6xBmWw19nqV54Ofm9BWIA1S4P1Izauj+PYP/Z3ow9IuFDv1Deu4rF
uwVgsxgdmMPIOXrUv5cGKm81ug6Vxe6YNYl88wQ5suSAhgXUOZRXHNxC7jEZODD0
bQqlkJMoAR39yac3Nh5Z5iAM8ziomSylQfcWrGBwf25w3gd1xBxSyp1lav4kdlwo
CQZQ6QPUYkDCPkGdwHMy0ETFJoquZY1HOa+yNUhwoe9nP5era/mWo47g7o21YktG
5jDl0ORV/1RfNZxoJcqXqQGdrOvod2zgTdHsBT8YOYAhKUka0D+Xzbl9+YDN21Mj
Wa3QHhNH4sGgotvIyLLzM3nsFXfQFaFRywiTSwbhEV9Rq8agp3tkoH/EYgpHTT1S
nsLe0y8ZNYUZh9OtDExiQegq6NIBeqD4Y46VxknHEud/TjbEDhUystidssK0whb4
Ly7nfAUreFvaRzPR7cEdO7vy+Gz1nYvtlfCwVFiWE5MB3mKZIRceu4C/tPtWbsLi
R8Q3bD5Gu6R6ifaICUtMxG940rdYlI+DDRQFycVp2N4urKYeUYrPn76GmVzK5dZN
EU2QzrvetIW97yvvUUv92akus219cxPMSFbqNngfuk3Qmb+hXkE7L5wF2Z46hE9s
+KVT5foznt+ovsT2Ljv2QAFjgVjjNHjwVm4HSD97jCsvfJ3qa3tV4UEnxBIbWUPT
QDKgoknzGrSK0lPqslFgmXQrSmlxouiMZOP5G9C051Hj27zHfnzehULs0jvzzY1Q
Em7pDHGyvpa1OvRE8bEmzh1l6D7Z5ZrG7s1MZRqjtWiZf2fLc92YESR4JUpbRV7M
GnnKwFtp7aCmWAancrY8z5WCb0rPRU35xhuaifyStt6Lfc1BCkPuBhY3iTjtskYs
jydppqnsfS6ka1X9dy3xBw/+q18oqM+lDF9NdXOcKMeQv3R/vRRXFl0Y+yCQHQgI
V7eboPJPTnA/rmiCrNkNFV23LfngWfJDPU11wlHWgEI2JryNIrGe6toG4yJwS8iz
Uj4AtYEk3pjfvjDX6Pww1okwhrkarf3pnTU5USZFiFxvjCF0uM0LcN6UsqHI5Rni
X+zyw6SJuwt9bvtSX/579OcUrmo9QQD/mbPykgVxxKlJgWWd5Lzf8LXg5jdz+VIX
wqkeUa8GIM3fsn7q1EWawOK7tkoLV4BI/FEd8vdpdGCs81L0Mn6RtmotfuMzkCcE
U2dJFsWrIeMGiwt8ioGlB0tbn9hZ7P8Y7jve9DhUAEI3Z0Dq2cG5WttC0roRSoYQ
vIfov170Majp5vwJ/Ab5BcxBqDW8IulYenCE1gYRwsva6Q29ofTRnWnnyWZlCgue
VY2f9KBaYwbJ6arvk4FVq2zX0NAdblmN8oiYAMeebyMwoWKUfzXcXrtXQ3TL7QoH
EdFsPwbACmO1Y0CwpO0YO6fv4EQwZWQKaWXVtJzc996BGCfNHXffFoTJ7djEI+qu
cfqRyZgQjWVc8WmSdG0lsseNYHYABe707+v9ixXlBlYZmuR9LoxrP7iUmGhVv+8Z
Aa3tqO/5Xm2NBfuQCulM+T84r1P5zIBD6lp9ROPRLCC2IjnhHbN0UqQWC5DZ29k5
EQCm+QZppU5TvutOGVXKXuTjISZRfGSPzyxagjROG4SCT1zyhh8mCTI3gbZUPfIj
v40uwfOaX7CIGANOIdnp8NB8X6/uy9TLJGHc3ASGWZ6D/4cnf5wRuOrwMQsTnYst
+YIz2WDaUgjFe0DmjPQNJdh8/g+lA7vnjZkhHSoGhQpyVYtgEANYXwhV1zC38oO9
g6wS4Qmfpm89j3qBDKxGAI/mOSGZ05PDu65/+UhcIrE34W89kMzPdMAkBgZ6rnP5
IkH6/64ToPg+doPtyKDoTkYjCfT/LIWdul6SZnLGSUSKtILJlZ4QxJD2JRrMlPCu
iNvlpGjGUaJcczGRxBxwvXNGxBWXjKzjgnmTGrV2NmitWaXpFzP7Y6Ity9ppdynI
k57c8hJ66CIBKzCRcgfrw/Tdh+e+Y4WymQOLpbPnp3u41U4nVTVaycQdV9d0XuOk
sQByde91546+/xEhf12yZsgEB5h8wpFBen85IMVZ0mPfrrkXiOeTTIv+36aPUnr7
3Xft+fWcU2V/jL72ecNFAGvu2eNgx8WJvmAO7/5BmabdFceoJ9D9d+FapBzM4AaV
ktSA/RCV8HNfDVT9xvprM6owiTfJYNVbjtOYNsP78BYbOTatvccN6IHIJNdLvqFx
ooPpXOsGUpD3w9dTEgJ9hBJ2xsRtcFrjuPa4uk3mMmcqcLgF3Qm5m3aNa2Ii2TvP
rqfBrNqNpj3lWu9OmWdoXfcPba1k+7r6oVmzW1vVvlOyR26l/2A84o10JO3eeFsW
ZlxJaI1iuC0H1t996e6aSzjGBRsn/LsQopdBnzRSUwnB3Etz+4avc3x91ljtVf9N
G4NlpTz1aGe5P5b+yAyDHOusoWPlFEwzTaxvRG8exndeh4jmf5ymGfVqQ5c144Gs
5VUZ8Zxcstg1kQZfiqf7XsLPAqCLR114gcfH/aAYQ7xpqvDaJ+g8s1ZqwkBU0OmN
j6lhRY9MDOSoicXfBocYvGJNOi73mmr1ZWh+L2P5F2lxCoEzzcFbbiTK+eHgd9Te
+xCOiHcPjWatWIsvqaclVn99f5nyo/QqUFYvPg4lM17iV6Tg5hwRU+0xjZJSGRjh
hCJj8oGgcKL3J9gwZDppLut84FzUXip4ZjYC9Q+hQ3t3FqNZdgp6GKlCs/DYkgIm
ey3EWMCLOhQtF6v9WczYRJKLNcyOt0XtFou3OF+f/cj+Kn9RMFprkA3ZqY98XfYN
7y8grFFlmpPjMfQ1r4bdxrsFjlbiSNxu8SQxrNiUBr7mmuTldI0vO0KFIGQ8Xg3V
jz3fCcXtXc0p6y4K0Exw8yw5Ctf43VJ8jUF98L0ZpjoqlvJEwNYjf5K56DG4zigG
FRX/eKfjYYDbDq6Y+DsS7VTuc9cBs2pZh9kNAwF9e/L/MDtKJI9EbhYdYmUYWjJc
wXYIV7mhHTiPM/kXkLuCD7kqeM0KxVntv0EeXeSoE0PVM1AsoRhLgIdWOXyBh9mN
qj1wLJYMwMtorzT5b7dN4pOZnUsXQ/Qmd0AdLNnRS+A0sVeE/eoBNkqyJ57NSjYO
3DS6kEBOM9HXi+993UAcT2vBkP2AvHf3UOxk1rIXcFiq6d7Rspnyn2U51yhGVpTu
xLeNAW7W+xIU9sc8YO0h/hdIm9SdMkfIFMmG4scJ/BBPyouN/PaJ0ZdN9g4d1/6f
4+3chv1agYXTMCiFTJ0/xEun5dm5OYbJMNbaeFdXP9EYOUlsgJsxV/dckAQMrPTy
FicvwzSzQR5zA2Jhi4oGPIfAKQXn7D7aS6nuVCvSxgjcAiRHHQztuX0mT6eASu1C
9BK3n2cbRX2/4lnicO7OH+2QQaX4Zyf9dVjkPkL3Yn4NE+GSmfcQys/EI+AwD8Cu
rEMUbDl21i8hpASnp8iY6/On04Z2e+JSL5R20DytSruO9Tt4ehaQbus/rvP2JIIA
9PItgpsYRxnks4hn9zeym/WkfgNkjgTKiHOtrS9oqaiJCKcSHXnJmis3fqYXn2kS
nFm5mJhnxn3Mfb2sQwHRNqdzl9jNLejgkwUTcNa6M+LbPHQVOPGXk+DSqXocriU5
G14xPMSg8VBBd9rSGz/7CFTd314z1VrZtm5wVptR4apLZp3U9RazudEjtzG64Vpf
wz8MjShugyhh8z3ks3O3dkt+TOLAV5UlsbI4YP38uhdFrgy2gumWg1iR9MgznAg1
1DXWC7H/Hp7kI9YE+wx89DGc1GcKiwEOYQBLeQTr9JqrBp4ROTc/81pxuUcVQOIZ
6RjfEuAlmtWrkiFsuTVVLnkvsnPcakDgh8yOCOu9p/inE61Ka6LOoMsgAmsxb1mY
rhd0k6h9umTq28LCkbmPQRot6OlPhy+j1h2iG6VhJvmLcfoKOaSZZJYf9OaTIc12
RoGyXreoQUsT9PV1hSKp33zeTjlzlmULWvY2P0NUQzW7g1CZKEY5GB72NbzyOQEi
0FOc5DTVVq2fivHR2yyVGKlzT2GFg/aJINf+GiX+vfylpRk0/yNuB68UaJwgWPP7
kOSheRKlyG8iv0alwEuDYjwmykowttUhYTs1cztZtAT4AcgWgkc07Ea5kd8qYH8c
a7WgWJ7aPknl0uknea9zXLBkyICpCbXqLMbRIirvZNVTvu0pgyKo7LBpnWuVdyNH
cagZBscfZq2Lf++VWpUT+jrxa99OxJtGwVNJMcJec0yw+kpcPQfB4mAznfRNd2G9
FYOsQJ33Lt9KCrLEQH+7+Uj+FI5hOZQfIGKwViq7VZ4ncSU2uAElEJu9nk4UrDrs
/KXZ4Rsp9UCta/w+U+EQB0HHc7ccVRImLSddkg3FWOBC+DmZne1bqK0lUN40uAwO
yuQ4xIvB6CPRgkGE8DtHHMrFc+8Ivfp1R+xDl/XxmY7v2Eqw1Mjp+7Kz1cDKqOrf
ca0WBCHRPdMDqcApW+FWUe6m/g+bXvFFtInjOljUxbCX/Jv36YRAQa6duO9JHPKg
lL+eZVk86T/ghedrD1QcybDQ8xlLiVhmrCrqj6t8hoYHErFdM0yb3W4CdOMoO/gU
Zyphs/YjWytoJ922OxvXIld/wjppjpGSgkhWVaeRXsRwEma5r1IquIjs8nfGyWh/
bK1n6fJYrpW8W5VQWkvvhA5dyM/3IkFsX4Df4sziGQEpZn1zVGy2pzLOxxDtzhwY
9sFy3KGQnG5CRYH/LCpyhh5m7lo4ELBxn5woNZieovY90+hKjQbyn+Y5iZt/1JgN
EBEVQEmz/qM3HDo1lWm9sJopA8PuNLuzVhaiRlqZVfIC8JrqcQh4HzlCU2WRUl3i
uwbbQkJduAKxyCMqyeuhno9hbkRqcsu+ZNVtkOjc9ctx5Z0sZ61rrKyIUMbSaeGw
wTi6GiebL8ns5PTxSg98oAs/ckDdKAah7adGgFayUV3ODXYf3eQxRUHG3QCIuMtJ
sCeIlj+ZOyJoTsacPnJn+pqCygdk9uGSSz5PXnVXAaRroNRie0KbO6uPkfcU8nsC
cUdIQqauJ1lkug3/M13mZcw9Oe0EOf9xNaQ8LBrtxVDTItOSlhnClBNFDAmr2Kko
pjBZ7S3PEakFFCN3o13Ewvql2YU+dtzYJYNCqSwUZZ9fPjvbrFXA/KbByNsIIjfv
nP1iKIeN7Oj3GoxngNB2AsZXgpT9HKFwjm6VY9JIAp8oX3l72f4ud++0bnZ5AkOL
VXnpVeOrSLR2BojrgHkHIn5dde+w1afARhsDU0F8CiSreU4JaN5xlRFozDJj/BX9
HKokgshWKPgZ9ywukIy9NUkEl+Ee98Nq+bdkq+GNaHlYhWNxefXCa5avqvjFnPtp
Gcc3g4wPpCRuJ5g0l18M7uwxbW3UScVpCMuYLNF4j29Iq5QTuTsLRl9zUQTpC1VN
4VvbEOxgtVQrQVu/C/uH7nz52nhYvAz0K/6zocHkh47amrp3yog6FnixhK8HF3xm
RRo2bMlRnq8wD1qjQ3rHjH4TX2ddt/QZItHfcRuYrWR4eDghZOJ0a7rbr0c7+vSy
3jruAP2BWe26zqEBT6O6QRIuPiTIYlfuScDcQ571bOy9++G407TBlEjZNgUCQRvW
+Bw53uMQAZ92Kjfq7y+Z7dpPAxvthRxinDgHyT+Te5tZbYn55NA1/3/brPiZe8M+
Gy5FnVnCsZuXmYg1mSVmtvFANkQpuDbVs25tqJolmVcPrUk20NafHN1zR4UWuDHN
RKHxttqPZLf16T9J0DdbBygs0aiyYgLa7I+PDVkufIJxGm0YnuwTJPb8O55zlVGf
40DiNUoDZ9183wTF9yU/D6lFYYbCoNycRiOeMVxZRGWMTnRYlz/BVZXdB6KbUcyi
GTsIu/gh/Qw9j9brkJJgG0etB7nKf+05hmm0xnkYfh9nKLrGYFTanuje33EyLAz0
1/NmX3lo4diGAnmYB8JuwkDP5H4FxmTCEh8b5JwsK5oXR7eiZdjjGheuqj8pioz5
RR1iF+PZoqg+rS3EAuTMCAJcp6nMwWrlNfy51UjUsy6O94RLZTJefICmRGtYvIKE
9+SJpRKPqCwpy7LHJtnCNvyfdOZCe6kWRuXJMYsD/1awln6zg5kqyZii/LhJcjME
XqbZeHp9JKWTVWBupj2CGGv/074iwc6MhrcpBCLkdnZj9SMhS3iRTOCpMfg8dzp/
YpFJRDcYSkwSe3yP5pVWIUX9CoaSykqh7G5vLYpJzeD0ZK1jqhwDk0KWjsNQm8Du
QeCdNgK+jBJvVSiChzjk8o8tLzglkHUGIRrSsABdt15KSBr4TwQ3GiEdD4xWEJkB
7PPjqiwh6I2iVl6x8YBSzmNTFupnuoTJx1oogqPrgp1FtDAowbSUbZbqZZcPecMy
FHCT0oQNvGZQUBb19L+aS+YnGgFoFjUt2G/+jq8J+zdmXMt5teofQWuM7Jzx2sYX
pxWvus17sUunecnMg/7kk5yPw5nOMYFNKlN6+lWzv64ZadYvMb87xgeoLsOvrtWw
/wk1ohWTQVXRaZGh6C1/LYD9CCK/66i5ltmTFHAsbShR3wrWEmTsaWMJV8AVYVwk
hEb55tGNMvQ5er0sDpGQG+1kB7yYfvlnk6DYN5jvUB1GIPgaxHuN5ZseYx39gVnf
RDTwD6xEK7da4eX6mILinmwJ/IjwKI2rA4s5i4yGgOGMQ23Ln0JC/xmM+Qjr3f7a
n9JoL+kGEMCsGbkJ+bylaDAzuPArXoWF8Sm4QzhkiHpdZpUVwGomC+pdoy71MA8Q
//c0m68qV27/o7pNjvE+5gAc5mAqvay91CtCm0jbp/SYhtijDY6iYsk6t6DaQoXx
+LljwH2bdAYBtojDDJIeiRqtaiG4J+iJRJ+fy2FxzlF7MrkJ1062pyo4mnsy4+gT
zDd6eJtdJhNSNKTKbHlzmq2/5o/EWvLF7FsAqUq/B7Rh9uFgBu9xqiZyVjndy/Ll
qRBJN83/xfwHZic674ZIinQ9T+onS6stL9sKx6R8VrWiCFPd5R7iTSNKH5aSl0I7
2nZcMcvwym5QTOolotO4oEomw+JaaQC7QYcKEOvA5LR2cqcH0RKmYnt51dMXzYNJ
DmwZSixpJtP9W1D84IuMFFLUYb6rLFV5hXB5LDkeHBRMUBq0CjhEDLO/HZCPsKQw
n7StuDUIu7OExE+khYbiN6jPd4+80zfuXnOYULClho9nxbjypTKDMhJwn4AcSTG0
Ozy7vx4O4g35KupV884FRTbp2+2iMc2kAQVuYrWaS2c5TdScCj+QRNKkAXmn0Z/y
5PtrUW59ZbCBf6qvWFwBJNam3oUh61CD2j9ySEkquyYKAhVE1toVe7TWo//9WF7L
XmfVSuDJaHZ8jSH27XlwIMMVXv3T+35oRwlY6YJOjNHwnZ9cGdHJFHxaubyQxEvX
/DeobwE5iDGflezk4iwdSzDKAxEaMY7iF6ulUt3G9aYl96Eenm1EYzeATqM3OOQB
TTtXrtPUeG6UNPRF21eo+0tfUrKlVqCYgzF4LjtIytjZdNr0GT9BwayGH5IKin1b
Xrr+9Vf8EgT8eCJG9IiMuT2Dik8O3Bn5bEXouE0kDflQuiL43yU6+bOMM/83pbKr
HQgdCEFsFdJRgqqDAUTcwhSREw4FlElan38kB5VWpt6l59LyWCBndQEy+DtHvV0D
XYxiKwD5WqezxYi0VR0vg94J2bf6cdS0fJMwQl+gNzA/iuBeheLFPea9vedopdC8
Gg809M6I2LRG/DcJdp7Rd+KmKHkfPf93wmLTtwxZcDpJH1fjxfcwZGVu/0pHaQXY
knZAqEfYaO9eUrYw8gbXOJm80Mtds6bwFhxztJZz1GAcwHtjET8V3o1jjUh3Nfc1
BnsdKWy5kJHmReXGe9V4J+7SCz67K+akT01W3Wkef0OAkapLajemr33UbJS1RMDI
F3Kzfi0Khj/+n7bYGZTMFF1z3ow19EBum9LjgebRkjJ9qH+tbU69UkKQITSEv5vH
fQbNnrYhb9lIOI8KYNbssx7OtyMGO3kgQ1+4BcK4AxVDXUIKWH6XWnk/U0489uV4
7UM/OxF4KijhuHbZ9O5QSlFlk0cA8IAUTgUaAYAuCPASHXu+xLY1S2Nx17Vi4Dxa
iyisbP7qFE3qtoiGPcqOoQGNmi5ojSd/WVGa9WftM6r+ggjry0Fktt+Ru4o4Yos7
0CPE6wRfXZSs/CWUyQntPHp6KCUketMIKXYLATCUre9JB1I53TM5AyDH8jIxzlN1
xLhzTPyAkuzxNx1ZMb2bistEFoi71fHXjLkB6NAO0abFSmhJTN1X+s2HxcI5MQEd
GMSTn/3K8KxstRlWBX1THZlrEgTtYUSfrHR4DrakLBhxkRufzbEe0HWzc3ajnzhm
0s1wFIX6dMn8CU5UfbL8mfmpWVwUbL4pui7+kNM8S+z66CF7KMqaB2fOXw9jyneB
x1289f3vbSsketkRtU1gJlHgq2L9bBk8WVrFs9WlUy4AtkYP87Y1vS2Y6Zbj8HLT
W9sKmj3rhxgrvyzEcqswu2fkIPSvYOcmz8TPZgLi4nEBRFa4X5cfQpd3oRm//PsP
g+jNhie74J4/+ykKzhgtgrklxZPUzx4DnPYYxYdx5iDl70aqzoz3O+lJ3g7f/LgV
iYY2Q/20ATFEic8abEyB4xSo6UATjOYEyZJKdfKG/GvPiH/7SdD7w8CJrLx+7ZpV
8hw0vyqOuLLsTmhZS5h6bOWDEyrmwggUiI9R6PsgnxZDgwqapyyAchsCME5ph4Wg
WPaqR1VpU/UTxe8Wkf1raMcEPWnBa3ht2Dh1EOh/ZRgXKPIIPLcwHOJk7PxsxM5f
+4XkW3ycEOyKC/T7PXHt6EP7k6bTrLjBhEAqKnsFycVSIadhoimqXpMwpksSpH5O
R1PmOfwxVxloAg3pv/Pl+LHwIM+Z9QQyp5Eo3uhLF7T4EVAndOk3diHN40DI190q
Lpl2ZklsstPrE4YMJSPKXM7MDd2vgozHs/b1MRpJHvZk8k4rnp4mSoCutd919yMk
cUjS8dsuS0Qoy9mg6LTJtHGTBXBQyqz9Ny6HOtYiXgK8LZa9nNVdZ0cPG5mfmLVC
Fcn2zNp7TbNIaaSwUfxexoolz+MLwlR3pWQ/tfShzZg3KD+ocwpXMfyOsP1FFfGX
x7MkoSKzsCEoHXFRZ7G0ebDew0kiOR/EBaRLx+4ViQdqIcH0DzETHfbpOD+op3lI
QGklvLiKqD6gcnHv5q/FE6y39DOCqUPegqWVg18e9BqRIG2ro1rhx+HVW1ymvnSY
CNLQLcu7RvSdjkoHCEHwJw1GpYQK0NAm+9jxQ6uJh4I+QyOV2uVLAWHOjUMoFQe6
Sz7hECaXtZlHyoE9K6QzJ/k8KWVUH4l99NHBjjBDFS/KuRdxusCrBHZ71uGsoYeq
UZZ17xMmDNbM0J+cuNhpTxIoL2jr7hb1fLCWDZ++TUTITuEw17ywzkbRuduB5W1h
MOPgMm2xQcTgFeCQGvHxjPdqzjhosdxF67mlJTwizU0g1AKLAei+UjGj2P8XayMa
/a3JmevPUnkhtFJ26j7XdmZbRiRlPO18TC3y0KwGi7syi2/mG/2kZ2X1I78YftBQ
j/BraGZSnPnvE6pNl8n4sOr1+x6p/hRf+fVhCozmdh71zte76cDfmEz4IiyJroEm
rKvZ9WdxtGmRJt0ukGs2iv8YqzEQeoLC5JhEHEq57JJZiRqPbFk6smJFBRWXPjl8
1kugP6b+9ey4ce8EZBxLanyFKzld64mR6ffY43b59glF4DZkW5kPxPAZ30JQYH9b
oRTKu6rzF7v6ikMt9kxTqWS1RoEfrQkwAhY2jvFNz/NnEccKAuD/aG5GpEmjn7yW
UohFJX8s/bVK7WWtZaGRxAJFNCztTRHrXEyIUITWSL/2wziss1kixwZvUx5ZNYmZ
jydANBG8Di7rQS8DS1ps2Cu+MInG7fFDOnJJRP6TuZmUEvfaDo1Scse62rCkwj2W
kznmR9ZphzoxO0dsnuqUqJYKecwkSS6DtpvXRUjQu0XLXTiA2S+EzHohbbX4oAUJ
SfwHOYhncRxfpxdvmaTASVLF56/bOz+uq3/mRN8CjPttL30eHv2LoGJ1ZwFM4ID7
Xjk+e5IW3oEJOqqkXfytaI3xF9pGhSzCKAE3aUjwiu16RtkHcMn/3U9jda0gesHn
GY+h5v2mIKryAlJxiccWYkOwGoUbqVgiL/VVuu2D2PKTnxTiGtH4DoS9RKCYieuM
ieTEudVzQidFLjG7d0x8YYHuICvogR8ClUVrhPlN/7yH1oNvcJMmwHJ/uCzcop/p
2vdxOpeZqR+Mj0oToVZy2edw8r5hM4s7feVcFg11Rovsb9yW6zobGKP8DygzaKue
0Mp70dpV68XnXPFnu7TEExE10P20xCf6d23aK8bJppPCJWJIYBRqlxeeMLKW5qZA
tXreyELO7qnrN8pkqUXx/tH0KugtcDZIukjW3Wwl59kQnUZHEiBrBJu47nUvydPl
27xyVk74c8DZy6GaChwyBbXgjkwcO8X3e2h3+xdWEgmvtnPOhMpdHGedaW9HJk80
YrMvVLtZ7j4bdAZYP9s6SWKkWGqjYRWgp96rOXz2zmMVGkJI0L79uwUP7KxiVjjI
ym/fOdcCzwdLyxbGv4lLuB4BUd05BNRBGWh5yR7+KAtKgjeIhfGZP26zC7tU6Ycj
nUQBU0reA8KmiOfaiSwQckOR2/mR/a4jR/mScRiPM9MoXEqQjykIW7ecxs9ys14V
putFq/DWWajXgriOOht7tIwCHY1DJ1INf06c7nhoa3xseKh5DvlVI+XYY1CMCj+l
Jj5gZX5ERPJ806Ws6wL209bjixg98fr/in5dIYeJ2LfvaPal0UCy8RrdPbcEGMZT
EAMWH0GtPsWjNqAOx2wk1+il4VKNWl2EX/S8/tJvPuf+Tswy5vp+Mx+A7Q4UZmjm
ZAEkdiwdD6eEk2r9ao++1vz1Y+t1/Nti2hEmgVEP8d2LUn10nAlfl1fLiBdPGAit
iDpw4KuJJjeDYoZnS/msxloCQrdJAKlI5Fa7mfQWyrAfm9ETHin3VK0Fnsge5XoN
qUMBNtEUVOjsXeeN4xJ55Z1aElLYDzbXiSGcVerlaF9fF7CUpU9Y3sWFA+vUo7MO
SnYoa2lu1DiL5j/Men6eLhWjMPflXRfAhUfnX//A0eyfWHeYwOTe59b/+KXuDjg7
D/Mw7K9ZWQBz89sAh6FLbQroNjL+62VRYVq3pYbxVWWnReP9P1oVCUfJt3PYqHe6
YLz611cwnQWXihIdAVOouHPerBKDF8/Yw4vAe+LVHCpacoKMIOT74kC4GuLHI4s5
rVqQ23QVXxk1a8bpHKQH7xY9x6a/RdhQAsD1HvQMJXZ1j7L55zwXVxncDDfuuAAa
OtJnjtD8OAK9nYFlGp2/iaqAMA+kPJukh0/S+DurdgI3WUIr3IjQCOT2UTAhD7Sy
GsYtJj/9N6JcyLW6SRyiDcqQ+DtSnzSmGAtKAEa1UoNlyWjd81jEOAgiF8NRuInw
adsy6djkt7i03gBgmbvyx1N8mbubdYQNyq+V5UI9wWlG2f+BnMCuFvCOHTMaeYQL
5q2WNyEKFFq81afxhT463emjhzAzmU+3Ts5V7dZ67AI1BT3CQyBFlD0ybfmHYSQY
9ffAEO1K92rBis07JBa+IB1uocoeELxOqzs7DXv5JWr7PF5ZbNVj2/qCnhzg7o8M
mNvO9K58nxOAQ7fKXsnvOkyWgYAZbKCQJ3mUXJgUArFV30HYQ+dJFWCFQcdtPwLI
eYZzs7v5ZVVK8r+YpEJqqrQ8M0n0ePLEf8FMdST8rLK0uxq0N0yNdehCkezfHwMM
wp9ERaw5dpvDLCaAvWe74NeA89+MiJcLqHW1mpd1nwFZ+hrsCogEzKXwtQR1lK7e
lBDdEXDCKDqLzayqzboKf0PjVHwjYyp2iLkLPWTQa1MmrXLuoA8MBFABaU1QQufu
nZyYVmL9x0DqFYzBG7AEArV03GAw1PZFIf94v7CGUvKkydZEitXWbGMLNex+l7rx
d195gkvpU5TsDoICtU1FyuAgbhLTV61ECcxL7GHk//+0YGG/YNmEkoSh5Zn2JIP/
oys3TCQs7bi/yxolZ+dcTIQ8njAjjI2IePYeMdzPMYbCw2RbAWp7kOf/G3H0pDGP
OFvl7gczf1uIJupJdVX3jCJo9E+EGp6H9ogvktBKpMoXsNULyjm4rVxVBP18V8cw
yvt7cVDhc00QEIB4LyoqbMx/rG++lpfMqoONinQL1CZJcw+mA2iOEOq3DoV1yZAT
3VfjF/ZiCXld9yCxWQtnmcFPmlqzowaKiY5vOdiv/0/1qcwHpK+svOjiHFNRJKV/
NV0MV24DlAHvfk675RKxyz3gq0stLzJJaVkFrF0FiZ9YGJ5H5HJnD+j5fg8+lHCb
Z/qdSfDRZZBNbU9Ypc+g0rZKo6rNm4kQHayToLRem3pnCzvtEBaVLfvaPFz5XHT3
W2S9VjJ5LPe+XCqlvIwZByBfel7uRGIYIYlju+00orOB0OplpwbMYrTbIEe6YjLv
ltlYJ+318a3x0RThl+yst40UyHixEnw0OKZ7yZIFstVCvbsduutZeMp28Ro400Gb
hbhYrJwKxg5Dooaa3leYRh94yz5XZhIWhIrcNTDPMsAur0ok7GBUjCQuvj7Ys5dy
iN11FTzMq3IuVFdwMS5K+lAEvT7/XqCjqyNawihNWP5e+AHwmE86BuTTXdgmI34l
ASDvdt+Icq2OSMrPaBQCUGiTsUeAKhHNGVHTEW9qHj9o+dndCC+kBRIC8W2j6mMY
Oqp9C6ArB5PQ1AnSJAMXQw76p6e2dNEHKjV+cleO3tEvQxWjhK2ouSd/GWlEVw9n
jXDxV2Z1iO1UNTYgLXQI1gZ7FUnvee2DCGOOORf4R0AYAQ0ksAJ/oNTJI6pO5P2l
VrqDbb/FpJXC3HF0gLkvsL6+uydZsABQ0fMv1dFUPSksy1qv0074GW2x3+tayqWG
M89PsfvNuL6/HLdov5vHuxy7+a6cqqpTI17/WiZYySUd+j7e3a02EhhhJbgigSsA
0mHGLHqq2GJQJddiXYdRk0Oj30nachqBKjczbp53hBK/PYWPfsvzGCnZIqtptQYR
WBTj6bB48SVB+5FlXK/8OpCxXoxE5WjIJl9H0BPH/AWhN0uu4ikEJvW6FDySM87P
WhWavMreoXe6ow0SillpJGmdcy4b/rdEBnxlC1oBFm7cHnFasLLphxZA9JxvPAHb
PB6jOdc5HBR/trHxVrxTJ1CKLOMIzhds267oYvULi4c9d2R/2yBc+XlBeW1NaHuV
FVghcRENGjY4eCGewk9AFVuJl2xAca+nCBrL60nY9CWIj1f/4f7IxAGIpC8vk4BX
RqmSucLV3ozEuu8MUuTENuedKRpgkb4gI1FsRAF/7SGKilD6PilB15KWcOw/DrAv
hdZRr4hLPeTAzaB4OIdk9PBYhkKuB/f+GVSRplGUrtf12qu9ETAycv1ao0k6LEtB
MuV3hrj1QRxwfdmFl4Tm9RhMCsS54vynHRqOxjzA4LmbnQ5mQkUPI2ZfZTckMO6E
os/FD5OBCjnd8VBuwjjuTzooaa6SoGg62pTGM0TC1CRbUiTTkI4h4prY7fX+Ng8d
B6ylVpAieA17NbDAKDcrFDPg+ENhB142KrINTX/CZZUWOYRWuiEXLv4xZ/nBwQv2
2SaZEi/w+Mu0Lnek3yNJ+bRbP6qrXAc+OqYa5JGpQY0byFicOVWESLrFmgTkcSdB
cNfeRcUj5q/WF9/ZZr4rD0b3O8hq8aSBEuaVRS3wxwlT5YVoN295OprZZ7kslXwh
HYFAep0s0NOn0BassmazTTD5yLKE7ZuW+HAlMvVEfH1l0zl/1jipsxV0gAfxWm0i
OjFqBbhdbQIvJeanG7XSrMb3WtS10VPNxbtTzDEdrPiG7XN1r2ZHFt48Lb5Lo7BI
Oqi1NiYc5htY5spzGP9UuW+mFAIVXNi1t/spQFyddbJcIVhmwB/rppy1p3Yqt/xb
pe/9UkbJD1ewwhmudjRcN1Jyc/c+JColECsRlVyjmoaZHrLNk7LWe0CUrCtIdMBP
YO0BBAXDU6gmC/nbLCSPeQSKT25JGm3bRjfr7sg2UpFhK39E6tJtpPvUnhQOt6L7
oixVY4ZNdXL/8fi+juAx/kzOOZdSqqlQDvvj6+sD8+u1eiQc0DWFnjHH6oKKTj5x
yyEIzzGv0Z3yt7ohCwLUas2xnI8Uqun7XHOHFmE+tRzfHGFZ3+KhTHdfAOL5LF+S
JWdA/PUDW9H6zCT2wuYVq53w4fQsLZMDoXVq35pyZMkewGJPlXKX9tBfkTWsD8Wa
FTHc1dlWk/ls1f6kPyIy8/e2IMM6ZnZUPNLx8iobwtaq720PxH1PZWj5HafcJZ7p
J80XVIgLYrqlxcv4PbeBHffho5aF2SpdEUrIoC33ZLDAX+exRgi1bwa2WS8Jnwb2
730vuXSGxXoz+zuGvkE9P0pyUQaZtZU8KHLqKCmOxvvR8lTtbd4AZB80tR1em1Ek
OV74OKjM91pxJ5OtRkjZXUzqn4ipG+jt5ukbxfCch5z2Dgu2WMi17tDwnCtfawUg
eorCvQmv8gDeluBA3xBjLORT6nfWy19qZTy6y1Xa/+YyYfaXZZ8ufpuUUaddOnwu
rKfhsKI0PHZQPE+wkTj2gSzu5dTwT44CfQJ4HPiTwFHZgyUGrDRehd0PLaNX5SCS
mSgdHGpAV/nFLKBVAyWspZYNeKxnlbczsoDpn4lsOyRVKl4Icu/ZWQjbLFQy3+6S
BFri0iUi62LDEWaMto5k7LG0BFvujYGpZTwq9Fpzp5KMv++La+MchnIeuYMlJAxx
mJ+utVTb55nYogz6MtpwdGGuVuGR1+WK8r4A9DvvpyJRXMPPLtBGIIXkGtDOOL9A
4be3ISuJUIVD9Vwz7NLvIkxBZvw/ed6EpHKz+xmJk42dNj+T6BCOTaQ4ngbfnv2n
gt2AXz0hx0ovLTd7zLbUfssHw2BersSYS2EiTh/CbdsiEWaHtFlAu/sDs3vdZci3
xfB5RGar5u7dcN6dMxXJkhXl0XWvzZ5kOmhVRYQKS3puDNkhR3J/neKvOnXVDj65
6dByRfUHQOotVZyG0MLeArlr8o5XwvfT4sX5eKe0yIhzk9N77rMdENckDpiIWrLz
C7Ai/GBp/61SaetPer3Je2Rh17ijhPV2tHeGuPB2pbJCSgy0jriaVckf9uuSuRtD
dRE8e9pl+0UIS/wcDcgclDaKfxb/R4wRvh2BBHyvOwkA0HgMNpm1y7c2RjgcwNi4
i0bWfM1BX0vswMnkbQXWvO+XqtCM1DB/BynlulDvqknUf0aKsgZsmGphsajY3YbM
Snm6WVUtn1WfZY3dtDTOZ3FwClZVg5vM/NHK9U2D/DkTGD2y6W8r3zChJNB+jF8a
A+VpjAS0dE9e9M7QrFwql/ZDO3j2molpPc3N9LO0XPNmfGKQNEaNJgVHe3JVPJAN
NZVTIqlPIhXQQVQ6u754elueh6MuhGMWxRh+RO8tnTIiMSh1r8K6qSxkA93DcJ8m
IqDYlm0wCX4KMxAmA+QBLYye+SGwnnrlsnaeKIm6eEz0GIdzitdVbKPo3QUbLdXM
OdRikKABxn3YqOna6FOiT8SCWLxUnI8NqjOoRvhy5nlGncCMFKRa7QOCsKoF4qT6
WQDrBLd866auLXZuU93wEr9bqHK+SJeUFTb8oAOshvKKyWUGLS1AtViY/eLhmt+x
BXRNc6SwMDslYVWNy4tpgXoc57qjP/X2FrlcQAJEvGbcZIt64T58tOv+RUe5lAd9
i/DgWXG9kahfNdNkWwyOaF4hdLHbDkBIGwAPKTckbUlvGpfq2u4mhbPOvsDY8zYp
sKRRfBtnm6SC4FnuWhk5xnilHvTlHAYYL+93EbS5AleXrvN2hgC0QO1eK+PJsE7B
+bOwokPXmeuzO+DcacbK0c7gdzNsgq1NFwx+l6WkM0TJFclB4aMBzdIEfokJmRJO
AUTY0XG+W0teUrh3NLvVDnYQmM0y89B3qGMStuUKFunXraQB+drd9AEbisEmS7ny
HR1/u9EGJ2nZWxAQw1y2upL419QLFOXzpqmnvREHAvJC2OQ7LbEZWtqj1JVfdnFA
/bMLhtBOyyW3bUg6j4vh+5nvui6WbeH0Qqrh/CSQsOB+aGR8mG4Vdfpc3hrxVFcN
j6iECQiSU2VlYLGOcmBTjkIyGHStm375hgSFIzGIwsffYZCRKVIFHzdPr0vOc96w
8djm5JXA9V61zMNk495aj2uq9O0I5JBsl52iEATVAO8LdorB/VmassVuW4rV/eND
Igs3rmWF7KWbltfJ0cZiTLoF5nsYaSsPIbxKvAEf2h74tva8Y+A22M+5VpkVQoAN
+5FVy9WPZz7rUl2N8OJnXVYvCHngfipPKEpQZo+6kEVi5lrNogxmGqsXBC4+cLAT
8sKJ9p0qjrd5ugPA1JFCfZP2+bl3OnmsrGMFJGiofVcuU6ahPPKT4TFngxR06Pvn
eVvlVWnEDzBgfQj9t2nS921FABjVNIPgZtFKuvrJmUVbi1i/LUR38dP7v/sJd9E3
4BKXZXVnRKZIQHc0/olb3Dk9iqmiZFt3BJLlPmEUUfP74Ki11zuXB1JFPELGuYcI
wF7PINC4PMzGcn7CaBOkCVoaCI4rHwG3OAea4CD6x4ISKem+8z+wC4JPaI98UcWw
fDcRI4Hs7kCY1UvZUXXaDSEIerZdh850Jj1VfLZnaUliXc3Mca98fdhl8E2DIyTs
Fw8t2L2dtQEGqKkMHHvo4goqQBrZaxqPeMHDM1/LJUA+20SNgJkzCN+Zs9zMJxez
sRy6+Ulgdy6+2xrmWzo/Oxvzwkbn6md2Mjp3hFtVyZ+Dd9y67QdEYyz5rBpQAMRC
LlyLtXmvvxn4sl9xIHq1CacqhI9cT5kSN5ltPkJoUipw8rIrp1E5kgyRYvfkuv9I
gvgT5ZxsZaRsZ2Ju4SgI9PtYRmdY/QGE32zimM+javWS15luANJdsdrf91QquqXv
c4dR3gW+WRRnrPJiVOXR1SjLCLrRVQBv2fa5nmlX5QIoz3BmGX7MPNZoedpOzoGs
ROrtz7M1hAEhTSch4qQkzoE0eCWcCBsFUNOg3+S4A5PepFcW88MBCk8kM/JECyPc
47RHnlpt42R+NWmFphIqUtsSuhzwyl9EiPLWhbN03a0RTPbJ5TAtA8+JKNGtpfFO
3E9q90R4pskzFZTY2odY0Zz5lu8py4POo7YmvnpwqlQbru3LI9BBhnWSJyZDPLp3
H7bimYFUy7jBHbhbocq6HRoWsEc2z+DrlxOVQ72gjydUC7FAAD72HuNPQNAm6hun
nnh7BrFu0I/SCbmcoN7AYt4+3Pp5g/7HP2zLBrH4nRE+CYAdTL4CiTCWV05ctsNM
lyMfiLRaaeG1KY3XgM2FV+BGzT5ahrAlbJKB2MaMtVO4/52iWKq7b750E4VAE8Av
TzIN14XO6X97IIAKb5FHl79H8WCGyueqAbSOlxCb/CmFNunzKoXy8KHAsrG6yZDH
ZdXAXhdJMAFyDwNwHPezdebk2k30iJHsH9URgxi+CY8DxYVCjCg73LfwhNGYOI/R
IadE8WonsZPsNDC5zPCFKTEtY1E1gcEAwX6G5qcIOdKvSE0uMOYUSONcMCQetssq
q8ebSlIkuUahIOcyDih9o7XOxvSz8Wtymb++o+uLnaBPOjHLZQtVZoez7hDCJIM5
VMQVVC3ZjpUP7syzIeFZ9cdhMujX8ELHy2diYpcvlnuaJhncR8UOqWTQsOoIgL1j
TpIeHtw0aPGtxEtZ1JchVMnYenpAe7HK0pDzTIkwc292O6Xu48ahibeEaZlkRCpE
KmFKY7ehab8Pr1jYXzK4POxtwxQSa2ZSKAqpRn2IYLha3oQnci9hRpZL8Cj43Np9
fJw3HHoJJsnehmCnE4jIuOXxI2c6liIZvpwK8KeGsLwWsaZYXCoAt1avozaZahNA
CcVW1l5ujMjCbWPJ1XuGRy9lzwsA65a3S3Ts2bDCqDxCPaB6mpxs7KmE9W2iFllX
I3p5SKDrVA04Y09BLCSBMFJs49FPXCkyfROSCovQQtWGLNyRZM06LQvvr/hSqEmk
pYfcVnnOsZ8LIgLNZJnEBGd1uS2uOjVPRukXeSwB4U+5vkoMfDDo7HNHb5QgZ2lx
SulJqriuZt2280+ySsGbyOIhj3Wa35ekcqzIL7PiiwJaCEkpRlGZwaWzDp2od6HR
jd2lYKYF8uzSi1RvX6ek2T/gZupVymQrNpxKJoinHuP1gVP8wlnoVUGa901FVr1i
nbbmts1eveYWbmqceL6LUBY84UK+VOpmVcvbuZjS/Nesc+6E4CxscxyVdZjmJO8s
omOhN9996Cggd5+HaCtcQM5QUgWkUu4ZV0HYuBrDjzZYme8BX8McmXUXKEW9gfyi
IErSzeulF/6WvOeh1h2i2EamjVAiuk0RdcR9eRyBA2j9NXx3pZcBbV0rl0P2gqhE
fQZtNm5ARHh5CixBJoD1988n6hZhnTECGeuwsn1PPa1G7p1R8XllVJF35xTTqCSQ
crf0cJ/xfthpmDtwqWULxPiGexFmzw2a6pqiL5+Jdm/I02uePiNzuCPCYarUIsHf
fn7OfkAVJh/m4+ICdbtnpaD6BWRmWPjRYZJIDWFmUrmVr+hPeb9g4d5GafjyxkcK
ukppeyZgSRXy7te65hx+EToieRp6ctrhUlBssXg0VEAriG7hc2jNmJosYgNUapea
1Bw0peELgqb5fK3VLix7GzJg2cqgWXDfxHkgeCCfB+rnrWeRu6zUTI07XOcYa+Bq
ZP/4S3esFqmOJ9g5DGvBNRhRaa7BMV1NMXhARQiI/kXIq9Dex4r81Z1z4B0d5DHD
B9F+OHfE7NfmhlV3yreP7L2uVac1DOdsjtb5CePzvfda5fSPv+emKFT4POkebFFD
zDfNHCQZ28RzA3A6YUFQRTOtYoEvczc+r7QR7jOg9XK2Orj5kqFW8R1oX8akiu9a
OXHk26zdfHJgPPhkfOvDX9JMu4n+yvewydKvxAbx6rledRdhZ2o8z2xcHGwFCYBT
NYfQoVqCTQdboEKwX6UJ4uo4zHa9fYqCrI49J0UMtyJsKOfUb3MMLwoBisdETVSU
hkJQUTIfiwhwq0+GeHSqufnO1ahapP74YBH0KCUB9XV12jP9wH2KhCACHeh3oJrm
gMcfWatPGq76ez3pSKsIwqJBYsW6Qx3mKoQU7xAVrzzma45hW0KUga3w3Ps7YVFO
adGBz3Lbl5aiDTQJNCaB5+foKPEjK6JnCxpbWZtNdyzmrRRUya37W2qkVN0iH/Ri
iS8wC0Bzvst3cfuXUksptjn9QNpbdjBY9vnsh+/Q8ojteP+TTmHSPjXyt7ubP9+b
Ywon7z+7T5oUM3T9gSiZNP8Ay6bozzwc+vZmr4cftBEDa/SIPs4vHXRQyScdrzAX
hczXY+4+yDuMFjb1a+f4kJrf1khpVP1qYhcDzyzh4iU7OUOrTpOMI1IBG/fAF5Ba
rsI1/UP4popmr6Shfh/babXLG/17z5I2nnTAEB0+sA2M4EDEjGufVK+/XUoC/XDB
OQJ/reyHKuVmxsxwN7peO5dbgWLk60PKy5O1mfqfHcZSR3VvfwfYOor+xAl8ZRSk
LQmILyNcEpFSWye/EJwdT2jdgoeClbShtoYTTraDa1KrH46GUI63N/P27gv0p5GE
DY9t4w6rNerM0LNV9XfCOMWsPYPDyhO2O5Uhc6OmxoIRLVz9trJEkb7k3XBM1y3U
XKAtyiXy+sYtfa2D2SzX0FWSOovmeT1Jy30Cky4HjOGImn74usvGNU31G9uFqdJn
god3qx0iq66iKos4IV+EekZq98Xb2Iw2dLaw95y3tEKl+PMIzfh1ecX2LeNuOM7g
itGKZkYpzbnZBY/t0zYmNk4oc2MruJclczdYfd1Bs/7Y0j9IhuehKW1WQB30XEx5
XVIfPNk/5Vlx/zf9SqdMNVN+XzltUXqMl8pHjRlMCk78QT2Twyfm6xZY6aeyFLf9
mERTHnVv76TqqzOEtnaFnPJDB9wYEW3CqSN9iL26LdyBnaj51g/qx7kiNGqI5Lpe
TUa6TGzQbqCJdScqPsT8fJN10lQPUMy6jbjBcXeQeHqKAYtGw9f3bkTlVD0B6rCK
PjUUgmS86sFMhoBr5zdIQxK2n0/xskwMMIQvVoObR5W3+eyBQqgAm5btJoDwjlKF
eImKUwDBkicxOflS6kFxbX/3kVWFwblCvffB56DiwZG5Ef0hvRSURuRycO5MhM5j
K25qNICoxJ3IF3h2YoqD0/Ueg2zGCcIo7yosG6vt9JpftVWhgdClqswnywhgf0ZP
la7Pn76uib+l6IC8MDQv9DzyE0nIFCqmQFT7U+MuCT4tIf8FkktNvZOC0/j0JwFa
7dQWrZAeSCkO0wk8oJ7y9ua+bJ51MeK8Rkjr/t9nGzzSUSCYvrLv/bZIyTmmwHXE
su2OxRmWB3U/nSMkmi1VOAq2rutqoChP0vWNL5PlkejFzqtZkjM+157isFVI0gRx
jog/BX+rtlo3LgX1tAJZnI01bt+po4EPwmqWUzGoUhvIEltlx2siEmklWIc/FJiT
O1Y6BpfVwHP2v5oUCiuf3XiGTJd4r8W4LYTRmk1tSqDTa0OC3DZS9GH93vAjrcpb
W+ED3eokyr6/whMIz2cZjXtagrcliBfHkJOOeOVrV9PFAlbZ89owQR1Rt/cbTLcx
sNEkEIoWQc1S29iCqdE4h4y9gX2T4r9cG3IhWGhjiHCzjH+UdeZxXXFwlv/OajXp
Y4V0Nyu8pgyE2fbPpQTjREr5mzDyWKcQdoAG4TkFdnkgnHcwuiAP9u5OYRn28iXS
7SjMwNIvbXNcmN2c5bd3K1VVyuBYvrSvRAMluLfIKY7DvsFlA/immNA8jsf1FTfS
vuvMFtbr6Y09KxiGeNGGX0skMIgRmLcCJPREpv4PivVee3PUhEkKBj3ROkpCi597
3DdmL3nlmVXM9gJrTDd8kmiwEjXh37DP1O11qQ5DUmg4kloncGFz+N0v5GfsWUmX
j+qImFtQDoH7juE+8IfL3Z0tZFrvUHqHn+SaR/g+3DZR1cwb7k1xcRhW7KxVJiAo
dhLCsqoXa/7I9Lz+f7qsd3Gx/Sn8pYO74V0z4syQgpbhTHGinLpD8NKjShN1MIfd
xd0IeT/biJUEbHNNHG6TOe0vIM97E/twvuNxeKm91+UUPHERIZaa274O0IDTGBk9
Dbqkfy96Sgnx+veYLPaVvqBEEJOyQkH0czVuGSvLp7TD3xZxcrEhTedAUsPq4RS6
VZoED4AuLbKa3y/ffpFJ+iCoBdGHR0qZralOoJrUkNTLrnU+iUKt9AzcImVPl0t2
SB/uzoa5i1hkatFsa51lHoALC1VIrHkS6RnLnMAuCIkgnAvwpHPd24cbeiG3RApo
GMQe5unyRj2dpVOxIN4zQbMRbpbzOAcpZLPV5LPNKl7jvirwcbDIOudckKcv46od
MEuXqOckrffHaxcwv18fslN4pyyH/fLRXCw1vH9m5KjCpiL/NV3s51VvY3ffcHVM
zEdaxsJr68U0kEJj70e1vo4KVH+SaOEUHbDNjgItfY3MtRjGoB6KQ9nEv1izvWlB
VW+HlqfRBu6b5MWALgqZcl0HQfMox569vAH/Sg0QsrKYHQ7ueA4UvATnphb+RCy0
WZvF7iq5e8quUgtu6i6V/nwrT6/DfoHrkh5KBzYPEMSZiKqDuo5j+823tMYuxrlZ
cuJZCN+C0m+CGGArl9AVC1HqLt1vwED6zL5NDWpS82QatiUDLqVmSpVNAtVcDjxH
FW95k+IFYlH0t2a42KUhvTaS4fOtUymHhH+4gITRUxb0KCAZtO63LX5FoaPXZx0D
2VHrzGHKVcJlmytzBEYPVMU7Hn7jG62oK1M/Y+RbCSN5Bv+nkh7pkZG3pNfYiTu9
tVH42MlG4vMhYx/9BWVRxz3LxBlIcwx2fvVgrIBn02tkD+AeYxPIO/NDofDLoJ39
svXmMfcCSNpA2/RupEFhNGfzJy8n+3wBuCOAoi5EqPTGIHMqp0gn0en5CTkntULN
KDYko932+o1tJoMDTuPOwfZwdqs8hOA/67XYI9nbbWYgxQpE8UulF21AaptKhQhX
od38PDYsUF3MXQEI9SN6ILwkQ+pyU0d2sstuFlNADjSoICaM9CE/WhtrRxGNuqVJ
CaGUyhimTR82lC/rFUvnnnNeOIOj66DaUkkOkhsEEnZBms3n/NAAA3gIO/CgZVz7
E3lR/Um3e140ODHiwsM/vOi66DbrjsMXjHBNvipDb9lWXbi3tJybMvl69Lur784W
kUqnLxbyHqZTtQTKZS2f7FKOFoAtCLdXpYQPQOlTVZ+wArlr4tMdQR0qEbT4SA8/
5Et987q2I6X5gDI5W+1eOrquJ8BlRhO9lBXe4PiB26YOHvDHAwOyZhjmv1vcne50
0qQNFbyVR7r4/GOxboQYaHifK1jcTE3SIH+/KxZ1Qz2RDm0Y94rJyzJJ2pAeD2fZ
SZQSGyh4IRsoSFWeOk41TwcBmWItzpO3/rKq4+xfeF6BfnkRbcFkr4bKw2uye/Zj
7OdkAAHGKqK+d93HqJkTHSRV3gIeeAChHf92k98JdVonnswd1S+l+V06PkpzVB88
W7g0CmUR/UwmwooGzb/cIpnq8DHoY9fI1RdWAeFKIrG+EKLpESP0F5ZN7C7m4/E4
ePZe+VyUYrktW+qH+VJa7U5eDqvmWe1Dpjq6Ukeo/YUAx41f4HN25/u08znwNsOU
hPQtzZ1GPZzqFv/03J3XTyDBaXc4vDZedrs4oGVnxi53/ejKWj2ucVaqahDCAfv6
fztueHAX1Ur1rQW0ljaSu+Fq73ySRj3QS3TofjVSCIMyAas6Nxks96l37yLFigyD
9Es5O2bY/2HwjeY1U99xsZ/h/g+fRkJHQZ8f01w0z+nD2hw1jPFoi3r1a1vQwbiU
06vlzvZkkh4Gl6lmw1Uzk2tL4E/jVvfdbSGUAhyHMjg3m328X5bzHzsKbHIQhZdd
AuJkd/rZ306aWOOR8ARegDEmyEzx1Ql4HSdrQCJzR/a1K9aOnguTynJDpBhjpCdo
ISC+k5PQk7qdmVJy8SMHaBZBZReIKC7XWGwNELBaPekgSG+O0Sd8rpnhs0bUFEKd
1mnwo5Rs1QNm2r2abVyobfe0PUNKdNo4mzbuORDvZYqRC2IKJIJJbfLUyh6Kpfte
MYRZJcYp0NsZTrQcyQvzGEoIxOhElkv1seJG3Nx1rd95x8s0MPLznS1a7AUNmrwc
vpysY/Il01NkmJYE4sW1sgQVofP2R/8Bs0+Ymrf/J05YgnXFvVDjsa63yB4U2oTt
loXb1QHBQgf2cFxrbzOcDIKNU2p3PgG07F0YVf4qoY7rfCMFu0kjJCY2lpZG5cZG
T4dRO+UcpKHzElr7Eauzy40YJNN25odoFJqfgTpUFYXNKM2/nSx2ApdP/TROURUP
LHsEfm7QvCfUt1Z4jQq9N2/w7fqaiP1Xsbt6kEbterf/WaVMJBTUm2LHKcCPZSKB
WrxMzdtbw2q2yd/6+GvjRAFC4cxLbjcZ5VMYOKQ5g6EGoqzc+zCS8EMbWWIWwgGp
cnk19BDmU0Xq/mUhOS8Giub8DaY1ckLLRvXrSPIIgJTqgSiDtnqixPRBWNbno82H
fFeQUpHtD1msWmhGQ5kaow7NGC9OFFwS7H/k1331fHQ9ImXJiw50+4coaVTTO8AR
s3vy0GfBRyPKMsYyeP0XwIlgB9lwjhRoS0t5cQborSJrXnaPeipMegKU2lvdmx7R
/QlSlD0M9xkDJ8Gy+S3dmVR+zliCnwjHGvikc/mpVGZoNd+GPp5XMcsXZMR3j555
nR3uQwfLq9HWhBGI/2HZ5SDjjer9960YMPDttdzb4JZt3CQw3zF0T5AhUc6A2oTt
okRj+y16C7wyb9q51HE6g+IFzdgCEbaviYz0Qaf0Na47932YnrarMMlPhFuB0ZlM
/iXfkrMdU4p/Bou8qIg6YhE++K8jR6AvmddN/ghaRnJhM6QU0u/sGY6kC9USA0jq
wwFYjfEanWLVGCFxfC+peR/IgrPNz0QwBpMcpyhVNi7b4lQU8ndJLY9t2e6NvkZ2
w0DWpdUeKFtEyP+GOccwe+1NRuJFQqFOd1eYigBIsoZr42hywIhgdByEuafppMw2
tmbIbVq1HvTvCc9xNEyRoenj4/aGm0iLPGtrRO6NIX0Gx/Vvjzz3m7isNz/jtidy
Wx3UA9Oilln6nyR2D8AtTkv9+wUhY//XKw8MRTy47C21dws6NAEQlic/CRU1Pj2e
DrPt7nmBRr5amGoNVvioyvoIAU1upirYEPHQQsu4f7lHNlERoSWXZ792BgeSMkTS
Bl63edbLLgf13QW/S1yWppOauD6pWYlORvFh6e/M3p74N7npbcmK/2U4ejXjfWOi
xY57DikWpQvJ1jhQQcI+6vCu1SnmQA/DQwIxIuOE8ti3rirLSDlOGB1y/leUZzT2
LeF4PNR4mxFGiWCLdkvK7/O2GULM8s65HlyWOujwdDKXKP5Xkgrm+p1KlxA76JeV
aHMSQZg2k5FAEhF0v/mh2TnylwygkomS0tsClxeP0Q6NTM5e8cN01ympt6cnNBNY
q9hxRlbaVwmprLkPgM2Ssxgh/5fXTRcYW2SVeZwHCW0Mi5DLHhxIgq/tekWsUxou
PN7ZHjDac71b6BeZCpWnS2pBCx5AWOWyMIwgIiJEC3BnQWI8ZNkKTpUc1BXIXMIQ
tIJ6fk6Xw/s5XxGKKHzFVOSfh1D0Lrpkf8GtT9qVB3gqAZ06J46cGK+/+xYrGiI/
VAci0DicqUc8mXhlrjxX5C5L/c6Ync+zwV6+HwQOBxn9HszPiKwws2/U2yO9QQjB
gVPkP0FkSjEWF0QKPlRYKtxpvjXwwrCh7e9PWZIHm6EgRWhapc8lFqQ4V38g1ONC
7mT8oL8QmxG5VZhjb6mS2jfLD824EMLtSY+7xM/9YnfZ42bx28cxsrmREe5aOiwP
x3p4pPfHUKl8zI6slEap6ZY8yKAl66xsM7E4RVFHgjCkA5uuYp+whH9oUYFR+Y+R
TwbuTv2hxk2xT1loCWjCcIMrYjtE1yi8vh1036DieRetr5E+b4shtolUuQow04am
5qRoO0fqTNybu8/++bQdQMPSUIwiJt+dHQl2TGFMLpfDSusrGyNdVBI23Wzc2RnL
CreA2WrTjQCmE/Cg1vAw5yy4TH6s61k5qb5P2d+xvBPGDnIX+16XWl+gNZdfsliO
Q6qKbWFq5kZASEY0ZIEuKCbSttISGKnYJHXbdK/gEMxO201ME+U77/bAZdDHh3fe
Rzb+gMWMwFyssA4ByXwvhdft2xr+kvHfnr6GpURZLvOg/RWUgrRlAjuHqC83bGnM
Y5GaGHlRmZUMPZrswPFQtm+ct3u4XpfJj/6RvNlq6FdcbdTX6rjYYFu6XNWFbXgO
tsV8KDXUyvlGR2KM0/PdQ0jxtZDokHsYM4O+q/MV+wQRVlcLqVjKNOuZcQzMIO1i
N09rmBVB2r5HzpG5+PO/NWAk/RGSvCOG3BFqeqaQPEaX+mzFnCZABED1HvwkkWBL
ASkf6Vv2EmFGD5Jegpur2srX6P+cl8I0W8qUJPqpQ4xoTCpYJmwVN3+/5swzX9mt
5xkLgiqkws6y9thpKw8qGHworSQ1N0OtENPyECcLKUv/eo72VverfUCuiRVBx2G1
JMHOnYVJwFSq5FMrDCHtSD0S+NUhPkeNdmaI4AO6aHiIKJOVJpvOgAaO02xL3ISi
iA4cLXdjSTa+iWxGin2O28pxINa2DBYtfRgM7Y4XX2oMp54zvQm9k7EoojbhSpvY
RGAkWbVKI3bBkSMHfLW6l9vkCTlbxKLe0HM5PFDvfIMmLd3vEuuuvtcczDXy5CF4
6BENSbnmNxeFdX8T8c7sske8S9nHqwfZb1USGISKGP9QBaNHsFL1RDD/jKRaJMUM
PSyjTCkOibVFR7b9pqsxQJNWBYg3fgCJ7GClLPB1KrQaExESyxekUFXMpbqU+IGu
Uam/1SMrYIXBzrCLJthU8q4+3no+zccgUXuFFj9fiXfLABxUMvJs5bclTMVT6XHr
sV4sYx8DggKh1uQEGZzDzAoyGxxzIwLcejFzU0xhTO6nvWZ3ttj6fmV5rCARpXoI
qA4k39zh4qD6XgWdpqdqXvjyR7S6AE/bd1Oc4zT8XTdohtL28Ibu2fNpYBDQmvqT
iPdWBjy5KM2c9hZpNtSieU+hIs1DWIC8M4YMx1w+8dbIALrWKtk7Xx4lCWORQEXI
NxwztJkdFPm2ikk3yN+se1peGquj2bfcJ2DFXe6l26U9Rinm3mLdo5rc2PDv24zt
bm6MYL0cGPqPhWtfH4LaqPkkc+cUSy2RiOahwrAWJ67htlysNL8NziUHxUTgOpmn
RCSpkkyE9TjbMbeilb3FPlcrm/tc7cUSHX5/5vmq2Z1dxLqgn95IynRUEl69Fkj2
kBT44BhitagSvUeZEsjOtPaqI28duFNWMgEqJmBJxHU5o/efVd69GNQRGuXwZq5B
6HZ8daIqSTqEIFVR3bqkTDCp+4cYxHwDWzwYaUxYogGtElQjiYwuOeCIDvaiERL4
xhyibVDj3hPPGTiNGkL/zazra1t9srqTdXxq+t6yA3oJN1xsk1TnBtqPndLAPDgr
Qq1u5cxS3i+/KZakyLpjIkJNdprEBRX8UVZagBSMDuO792EiBOhuR62vh+BBNzUK
hlzFDckc4S/o0Z/3e24AArhKFtct/rnEgnD3ZJv6j5rxV/Yw/U4dwrAt5Cry6BQ/
0qK+VxjQm8h40mSnDsiceBQp9Yqsy/0fLck6UH8xw6ZaIvWW5K7RXJg5LDXI3x4X
uaQbbTVCUq9jpjlNYzP2BxVq3Wo/KC7cFFM7fuJIvMqr9wldGKB6cftp2RfBAnPN
8UlrBvdTBPNkDFy6EjroUnt92KLGcFyHx0UHT3zkQTZHGZ2iZwWCZZ4pJcs0tO9H
Xlk1B1cjF5nRfFXngkqSTY/MhWwLEHXnzF+XJp0bc0X2tBjVIoNvwlaa6DVwOZvF
i69ZmI4+bMaD7YxAoD5usnl3pvf85QAl6S+qMkpSFK95BKsMzXF5tNvr1E+KlNTj
71cUFdV2BGImqVZY0kz7T4aq2azAp6m2nQiTeU4FLzjXfHx8/Rg8YQy4KACZHUr9
ZHYhx1xz0gnaXEI2SRp4I4sGq+dQLwtAjSgOzFJ5knldFyc/tXjwZo2OyqXUGL+O
BGpxxtrLeeRkT9w4Ddwao3AOF+lCyUloMvSjSqF4N8vV3Os/PQboscN/WA8DyXMj
8+8jMnkdPATXF5F33aZ1ERt2hrj7b0sn1vX0YEPzwZ6cFO5/4XA3hkLv1zkpWSfF
yO5JbSe/UFwuA4jH/8sA74ojyZVvYy+ZzxSGy/T7bInoJu2qa69hnCo9hXJgeSyr
tS7f7+PMBhEs4LSORCKyWh1YgPQOqYNbXk1XLpLodd3WGWXU3O/Gd5bYDNOpkwSq
iKVc43pFjcGygTK5UZN3LL7dJj7VyEV/zTZy14CC7J//1ro3nU50Qg+2tRd7xDDt
tk66UzZtwqKFPBNjh+gERCkxrBbUt1gBn7IsRMyZEsi2yLS6jCOSS8E26oRHdJhx
ZcEedflOD9Q7BcHKqkW+MmBv9trPXQR2fCHJpz8BP/WdIH6+52fD0WQHAd1yxAg2
pfyKAkTjmSVXibLUCzJDCWjmtpA298gQd/Nm386A1TUElxWiPaJOuANj1DP1kBf/
2VWZSfI2ePPt9bTKMKgsEzOkg2ZKrFMKvfgZCKedoi9JtJar3tsooMW+BJYXhJiU
RIpuTjqhZWY3Hj430jnnIg3l/ZnOSteFHw11M2Dfsvh6sRkd1FvbsKt9j+MR84KT
hCJo5dryfubyZSwqKk4USeVkRE+Ta0MgOiZOFdcdvSln1JwkKZ9YoHG+HPrFP0/M
tAzpt7hQvMOHZNwHZB/ajRtcOivZ5ARYnN3aJNKk/BjALXDg5vqLeuwdpNCVwvDI
rHqBs8YJOWswaRhPA6catzYkbPOg1Pa/DbPEEWOv+0dTcwDFS+tnW1D7cU0xjWTa
smQr/cFplKCLc7RofZzOfhwV+l7njuy0ZzWzVAW7CiRjRPEqzXpTjoj7StCjbSDZ
hGRRfMScneJo+/Tk78xyjuu91qaNjP86weOug6AYx1TBEf/k/MNOkPrphfdFyOPw
xPlmTSyyNW4SgP3SU9+MbjRyzR2Af0LLb+mxR6+NHryHiEFvcbLwIpOVEABwWhMw
s2lYY47rqyzE3NrhbiW/DrPKi6wAIwiiJpa0pZtvVg5sya4dkFXdOz9WVLA7RcHM
IArFcUdkvnTDbmD2DVwBmFJBg3hVrlrT5TWjPTkm71r9DnjwVy3cLGAGFzd7liZX
Ro+h+roM5r8HEAKW/KDuKED/Shn7bCo1KFPArqNChO+JKO265rnmwTdRbhpXrLxB
9Gd2PUPxdTTFM8gH0O+v76t0eRLdFG9kP0mMh6dUrlzgF8vLuqDXQwr/TqJfBFAz
SUu4DFUabZUMClu3xmWToDzlRhCVPFz14DTp2rVOgXPhk5INosLbIq8fT0/fSHOU
OJGdBATLYDg7cqtkm7qbyI7PuFeh7KTRNovrojd3hyCsev0jztZbiR5Ok3VdZCKl
SB4lwonYhO+Y8HxWcUsuFnNQ86o/Ja7qk6boie+4Nu3tT2Kjn0ygQQG0y2vHsNP7
eOtM3hjvzbuCs0/MrOq1pjOU3/J5GGIyEe+uURpTXNmyE1zOMvtF35U4Q+ajGj0D
VMimMQKiUZywp+EPzLo7NSjLw89khDS8VGiQWlWvWEukNQhFxQ7C9nEwsCZ1AbGX
rpFCOwDVaCt4AQpP2PsSLLL1gCGSmBNSPoMgjQSTFC+uJNpRrnvbXBZnCZx63JSr
0W5dk6czgdl03MP3bX6gpibUWph8RxX7MzdwohDLpnpmYPdOfPLP8Z9eopkW2M/z
cFRqWJQdg/HvtZ5pNJlEN3aotFppKwd4PS6SBFPiBQ2Z0KAspocCq+48Jp8v43np
k0sbSbNZ9M8ykg4qMRg1WiijiniPACax7md1zDgIj/518MOLCW1U3/o0coDgN5wL
fllQVSzjubAvB1N89zPIo0sEUl9ssuiEREXHi6TjgiK36RzOZj1GawlCbJrbGsdd
WoWO4fHQ9Z+0L5XxGiov3FDpECHXRUKhkdIbivdW5pQdgTg8pHwNkOqlVbIJIYj1
tQaEsL3kJPOHimS+MsyJ2l6AjclJOsTtUTgwdZsTj8X/zS1MzbSFgXKIykelafW0
mI4v+tqa6aE/QAWBVUISgrcu3dalG45PY7nNWaPG2op91fP29L+k9sLfnJYEwEjK
gPUzhuRNYEhMu0gpN99N0lp1Dv1uqFjexeKVl2sNdJACeK3Y/j/ylYmQrHzz5ALu
xXtLKI4jIQPR2em2yxnG2Ffci0sHQFX6zY5ouraD1szxmfINbiL1P9o3f4RRGpke
pQnpayxWLhUcqtEqA+GBled2rj9+gkK6tmJkPHMjlFSFI5nBKuMsjCHVCxC5DolF
wt9oK4AsQJNFnFERztYWiCtEwSYHFcZ7a+GicPtvaYGbzq0NSleOSFb7Gk9yuGMe
SOQv+flYKmErcwox6rnS+9bcGmkiu+FzEb9WbRnvmSR06ZEPy68ggFh6Uwy6qzCI
9R+c9AXIkc6evSDP22iPVcO4XqcJFic1YbiCLutGh/CnQzjbtGjlpX0+GJmBSNQv
yCcVqD8Vfg73F7Ol0Gw0fr5loBSHVZjCTkBq/L7WwbCHmQ04/zOVJIiAmIprYGXI
l9C4vEO9koRBVB2MHSIAvwla+0tG1JkL+r/1MBnNXOGlag2MzZs0lpkwGLI75nPF
WtAcG4WP0rjXr3DqrhlBgLBD8e37pR+8nBatVC9tjcgjiD6k+VaH5x9gP3eR+aCX
mLp2AiHwlXBEI02CUQrWGNpEVVxsjt/S+IM88U7zuLDJHolwvhEZNsXBcU8QkrMi
0+vfGebT1nwIY2GJCVl/B24ULop1Xy1j/LwDC5en8hCXTsZXHJdUF4CFyCvCGVOI
abgR/84ctZCBIUbH5QG1+mIEsQ1/SpLOopMGqq3P8zMm0ggixBn7IVCW0DLzlPPE
P5xO5kbCh9PA8geizPyWnmCKUS0MhIRJ2L/QHU+ezksl3dEJV28ykjUZSdZH7+x5
8R/AaSgC8V6e9ml2hiEV1eatEr28b7vqnKexjyorOqOhfxq3B6bFSlHrNQSQ6/hC
zKsuSgM5fL9y32H+LBHMiIE7Jdssk8bt9bHbgESIPHG1o57R7aXEijBKpKIkqA/Y
llNg6Gqa2nM5pEJVfMBskdl1wHp02pudSLF4WGG25J7oxoB1zzJfsAlV9pYQKEyT
SYvX4JbwXSizlC6VbPc/VBHOGbGLlWwWx0j4N89VQd6cZRj8tawZKKEL67wRdm9v
TL/MuexCQKcuXI7jXdjBuDTTrE29jH1UJiCFE9n9vwuIzCLpRApjgBKYZDBGaFKW
n1f/OpR7sbBKWyi+LEjpFhOs1JIJFdeIlKA7WhqoUJVWyXlxeCpgwSWMpNM8Xj2b
4gqRplSxbZ8i+NHd6HqtkkfSx9TEh9yEyKYiDJx70QynG7nak/DbzCTXS77MKKPE
LYIpAg2ZlCx8XghmsBUwbsx1hFJQP1IeAsYfFVTQdoURNoSuqAScCletc2eKmb07
hNOzusZ7xYrEJViWjJUc4wFGOHvVuztwbI/ApwoiUzifuQCaIfmgXQmZdmJgVgEH
knb3AyqIMrUBNyPM68sZOxevy8y6m/+7kEo42gs3+5NdPSN98QCnKPqjJvuJDqTz
EOilv9TlJE1rwbL5awJblBmfMv75/IRdtMgWZdPu+zJxDG1wNa9qidzc8ohOmFtm
lr5mz7adJZsv7NDID1Nl5wgWxaN8JXDKEfGpp+DU5jmn1u7f2NulnLTYQhQkjByf
KYwKKBPcoWkf/9Q0MOUInzvOVSMqWNdSxklYkrZDQqE03qluMfFDbZTUSVGo0rig
dozsjVxYWImCiZ64o90ymuH0QhpanHEd/fcnUoLZOWViUf7/2xRKMaAiISLa4lQm
5t23sI4npDlL+kdqsXauDY9P3oTvVHy9kUAK9GjKVNXwVdDR6EHIM52Tt5x1sTVB
xfMpLX6IhYmuJHBcCzPFLdUtfZc5iF22WHGXJ/5O6kdzeQTl00M24BR8fxdLtFKr
JgsTk3j4nVjw7ty52AsM/s43hQiD11I2tr17mrCwzpcrA6gdwudAWgZARemsZTp1
tiGHamoh1ufaJQ7K6e4aic8LxpNdY2lK2aN/Vvl5i0FKFNYM0IFaSGSjua6UID8Q
OgHdcHz5jd7UuEnA0vap8KkRf0GZ5+QugpbOaxrURqAJu5g9WXLomE7EyprFaQSd
FoJx+R2PA0iSKAl58oW+4YxMvwVQBL/QB2O+ft0bo36yFYMzhP2KlcNkV7IJBR7N
puhaGHGAwZ/mFhov71TArGh/6GtRFCOc+lT0CReN4rlWmbe5/2x37vo2gdP1CYJ0
hRvoPjkpLEZAQVPn7+/xnf59KUA6LBLgYiJM4QFTMuBNYewnbKD/N9he6/fyyXZ5
dvml4GO4Dj1n6mUXtthAxoks5KeXkLL8MKp86a1KH0Uo7HGQawvlfT2ekl/Uf1Yf
kMUCb66hRelZtbB9StpbO0TDWYFJdNI1CFU/OIckWUrXk+6GpoQvykGvz14nDB9o
pE7I/CTyyh3cqGSaxR2K+AZ5/qSLeR5AwDd4FIWJtDONyJSnDP3yVHS1tSto6x2s
7FDhfCXrCfyq137q/Gtz2quhwwa/m8nfl2s+EEoyQY0ckE9vXOlWSySO6h5K/hJ4
CCnsIFhEda294dFxSiCY86dq/LLaBaYhmpt9jL7SMwPscarE2VomuEpfXQigv5gb
DM0nM8oYtq2VgpCD8LZSZTRkPlcECO4G77RYACj1wfuRwRmdY63V0aGEDmgr65Be
Thm0ladX51pSmZVDiEL7KowZCcZW2i/d4KiAVFrUAF6GEYRq8GOPWqE4dfWBMJVM
UJhRKkvvxeqG2D0JFNtZMN9ibjflj+B7o/rEgs4mdYsGP8TsYqEEkVbLK9yl07al
7ffn2CEfk9VK0kD7d/2tDJ4wEDGqpJHlDDCvqzuVYOlQAPGLrjNrpFv79p0LAzoy
x9ShTRxa6FYS5k7oRIevWg8Wzh3QNJ9MLm0WXqW4onlTO4hUk92+U/iSQ4gv+LiG
xISUwSU0w1jDtHJTZrQa9dD0yx6GxffhXOzYuC4flKYoIRMKuDRhEbYa/8Q9CWGm
eqN4tA0jTQGYwUpz+O7MMQ5NmOBF2IlEQf5gH+vc9stndB/eAj1B946IYZUAhtf1
XY3jc0DB/daErmBLbLMmN4MlBK7riS7fRqSVagYDuvGScGceTlHRiURZ2qqa+eKv
q+OamIGxuXDtTmt/IFtstpKSiS+HRtjczuHfBz6q1CU4hpzPVakyCWFmjnJfGw0y
13y6MZEw3d6OhpmRZdr09zhSfGCVlXWfz/Omv/yzBXsTmT/frIeF/m9bIBaCcp+Q
sd2C7CbiawdOww3AygZarCrCCdTuzYOtE/voZmS+3avM1lHCD8QhuFYXypVf4eCD
/ZYuHjJBse0zq9nzqf1Ye29y2+hYRHSLTj6q0sS8Fj0P2iXR6HQGlHpsa5R4tLzs
aLvZaXCqlTF3At9q8biyqgYc3yFqZXzjUV0HVC9QXeoOuE64pVSVjsQ5rraj3hNT
qZCjmrPXkgUVZOtTXIVMaIv98v/qhazIEmQNApF1SwYdgQCh4LKZ1nukpExQYPsD
SJoSToNNrxSL3pDzAAariPUjExBc6RQMhU+uvU9hHncqV+4Jd/Rp4lBe47oWl++r
1JOqYKWV8cIymtuonFr96FS/Ry46y9Va8KinvmUIYxPUMmzdFn1Vxx9/DhSzjjf2
yrosHKMnkONq9RLezJVpfRuUjxJK5iNgqHnOdI2lgMfFIoLPG9/SJn5cLtOq1vSb
XR79Ip3V8RAm2uExsJm++0iHGk5kWaZMH8L2rJelgshT+1hYnjmXwG4rUzNAcvFe
reVx6vN4+f2cLAtuznq8J2YazCl2Ajnj9Dh9Or+fAgJfhUat3LbSZilfWLXAx16X
12yMSk5dRV6idlWOijHEXReat/8CmpNdOOC2L6owGNQuDKCJCWlmRH7u9ss+NRtB
+i73eXTNIEqyZxtzJUyh4Odo7ArurPc8iTTXwvLBl1hgmJntD/phf3DRFT+7YYu1
9BFco4LXQv2J8Nib2oM3gWUfg8nDO7hjUH0zI86/3LJ5OTIl5sxbxM4wLXR55/+m
i3EItJo1TrOFKkZQnx5uktA50SiCP2C7apAl9yMtqdH5R9ytxMitxgIydd4Ku08g
NOe+P4tnxgNXnyhlXHUUy/CpqnQTRFexl4dcOmdXHU/dMyqezzaC8GLBAuFBIJS4
0BXLWOeNsYuCWO1cQlzluklZ32RILlSqKOeAFskCQuxgipwk2BuOKck5X8EL4hXB
TDlVfZyYFEnogoCXA5htKgtzNxPez8Xq6S7JifeV0pO9jCSwzLdIKkm30BY5EBQd
MrTQFyStlKOfRMKhpMqTtoweRiMKJqfj3nGDfdZaRIcWS2lr4uLkCZdGO8OD+7Jx
LGQUFZrOV5+1+VU18ZJShgLSfibv9/jQrDWoc7jFxxKO4DMG1SjM2olZ5mHT8pgR
W3cOdRMq+qI+fLokle0d+NNt3f7QYP5le2qEASndn2bmV8Cnj74Y9GGVEkCBtSqG
EDfLNk6zdMb0l/T364o4evpUiEifggdFLUz/qlixHr6ZIEaFmfsU+j0QrSuTNL9o
I05fjUiyXLyXDdSxB75L1dgDdmynoTEG2WiMqTeL5TpRMAdbg8O/0YXPvskPE5kO
rztobooM+AvChL3k95TMCGstjjkHtgxQ+0xiMfJp81ynxjtFz2qXeySwNEu+4zji
3T1fPXPNsmcx8/w2kM2iySZo6JakP+d2kH5EOdXu0HJ4GXlsotUPpUoDHEtIrQY0
vH+N670GOiqahsAZTsj3j7PSKBFlpd6p5xVjESOu14CE8j6yEo+KT3QwKenetZgk
PIwD5i8LKnBSKSdlpTKTE+qpzXh2RPtpOYLIvtK8TwBnbEspWRlgc4/fewnPhE9r
Of+jHCaZ8U/AuvNEfabpFeq9fh0DRygDMfkmUT8TxllUPpcoTZgb4g/t4IWFmqI5
L0GxxwMS2Ets0cT2DRnW2v5/oy96rRSgprPzitwAKGhveIwVfcq/W5uu3HDmx1PA
uCm0hoFPBVGRfz23ufNGe4Jhu/EBDbC3byu0kX1Tn4BLKSl+mPLPxTvLUMybWypX
KZQz+xtc/9+xXkSzNYcDJbepGDj3fGidGg+7KqP57vo4T/zTBGkbZTtvrQyNQCpu
gQ8xZ1KBzRwi7YocOl4z5JxwAX2H9Sw6EbCCtgCZlyS4b2d6L+xEOu0ms1ynAmIH
QTCSRsKONF5r3l4szuXdJgyaWJd1bNa8gwWbMe2Dex969KxCvFVOvrBq/cUTbmYb
9AJF303p/qJYu5+Z8y+cLJQo+kOd3MCizVF2E8EGNU0mGwsKdIkgpkNtfn95Amoi
BEVea8CnWqxdygDdbk89HTcFG+gTJv1HYDNkyxCPTOP56xeNvg+szOV5ILaCQmiU
q8mu/QzqGvuctbL5WZeFEkCuMqhYwIJZZlKLKU1GDc3m9wtp0Ng2trpIB2+epPhA
4RQy8mXB9/TQ4JGwtpXdCv2vqL0ZgHex7T53546NFERSo+RWT0IU4NzJ5qz6nSGp
BpBuEtt2dMZCDjBg0a/gpFHfXlGSXgr3x8Z7bZqqjz6p+RrIZuUG80lb7Dgtvjji
hSXfnK8Yh1YH41exVtzqewBS7j1jqYVHBTHH+5N1gMjiPt+Tk6ILPWQgGi1rq0qq
hDuDd+ESRKQeujabyr3GxAUDRoVmZ1fCLNIkFY5+eFvn7ttrhOTZOtY2gF0zUpfj
8tddQKDz2mU3jhy60p+jeLBIo+h/lLyjwedjbV/RDHjAF8+SpDjU3jwuo50PY4wK
tzBd0Fu/itWXaZAmk5UM1DTLMVIdJTi5jwcWxOEVCyAabI1q9Sbd9PE/xM6+DMkO
PmkcPXZHDrQoRga5/KFfZBjQ/4OaO2GooX8Zr55yCEuU/cJuLn8AanxqZHLJr82I
P1j/x4NQrGRh5ZndITUbW4UN1NV4FCLcZZeOChAN7Nt7fEEn9kgH6E7D1PUlZOP7
krHqCmlu+o/SZ+rGh7V986ncUzu4fT6T0lhsAJYGPcdA/9JKDGAwxyMKFmtG5dc4
ZTdkCzx8LEvnQY2Gj6OvsLk/09/PdTJ1lDCp6JKWG5ZKchvR5j2Rx+jwOWeUsrky
6depSH6ciywQd8JdE1t4ySwdXC4tqkVFxpZ0EsEiJVEVP0LiVdrac9/c+wBoU+Mf
/Uxg+Ev+Og95qALRF3zKJtOMqgDbE8YhjazmiUt+IFgLEHXI0ER0SkvaFXRhT/WJ
ROxiLH2GHEqwkuLGJukm+F4wpwW2Lp78EwPRiIkBLm/TVg/fW9SDNzvfwS+R2kd/
sNwlD0AbeXqqt/8YFroSZVBbY7p8Ugpiz9OuRfd3j4q9kKMlzf6vWK8IP6AeiDbX
JqAXK/suq9kLfdRuAtkYQAh7VQxDok7BR9R34A9ihJ3KK12KSDOEj6YbcBKIJBHC
xokvovvTqv2kkgNtpnvJBK4kqGugTfbEvJjUQDCLtMfgEPYZIzv1+ozNKnNp5d+C
HhKg+kypVpyjdxRa99OTJfdGNWrNgEzsWUNSaN/VpSglIsB6OWunDfdTO9WTQB29
V7VLlV+N5TU9IsBW0q6JN2aNqOs5u3ya4LS4uGsoCM1k/ux3Y7i8pqESEbsIZoDY
57puhLTlVftH+wRZC0w0Z/6BxGJwPcyJG+7/p51+i0SfDJZK7T3vWDU2vrImiZeW
cVE/8agqphpgKdT2BDxxmKtgbvFBPLo04o9A8IAz2HT1l0b3UgTlIDKyjK+4JXg1
DwExGkeF0nCaifm4ysJJBdVqx7Jtjfpe72UGDjxx8i51io/vPHrWSxbdPFdiLRVl
P3TIUlkXH5ybr4n6JPBExznPl60+Fbde+S9YLmfH2uhlVGuAa1pikbjer4b56SdG
0ZMEW1Gvz7PTfYgy58U3KFJJhh8C0Sxmum3PYOD7/rs4nJQQcM80/FvzbU+kL3j5
9R9MznOKZwSRUqB2RsPBsvrp7I6BT7nAsYPxlP0FLeykNDd0tBZl76tfqO3cYVKU
Gj3xZkDn4rP14Slh8BW4/yZxBSn3OfymVa+lx+ixvx3J+yXU1R+7XFyvkFqfW8JM
c7E26nrOsG7GTP0JyT7RHRtD5iLAdsAq+Vnbl/qMRRm2Pv2UEW7sPWDT8RLYqZyi
x2acXwXVT0RnaAJGsugNPnhnnlLNXBqLyvh9noYnmEKYsIwcIUTRdReQwbxSV37Q
EDIprH4WJOM22aZkx5lsgTM6l7D7p4wF242e+41WDaX2YbPgW5rApwFZqEifY+Ur
zcXf+arpYo86bJ0mS9W/P1WS0rDsMxxNHcO9o2u7Ni/A9mmRyzqUeFN9rS8UCrAA
Rl+MX5kotBg+oGVpwwT8j74LTl7wVRZ7ro1aQqqxaOiw244m2Xef4IUxh1ri16kf
nMG7q27TxkYuQnfBbNw6vUr8NgGXzBM1CMqIcFUZ2ZHgjasZUlxE5R2vPSkkAU3S
u6SStVkhUDqxzlDa2f5AqB3FPTVFcP3NSDfuz+s6QZjNJ6lh68VURJRcIl8uUsjM
7VBH/39sHQEJp4mYHzEompGlb6Uma7QVEPr8VfyVoRRb1FG9l68BMu9CDKuqxCIG
NiKqz7gMGua+nTRXfiJgfMjmhdmfXIE+WBVEaqVflG1/lHzWMMgcXMi05My6ZTT/
NMSJjxzbbPDll3kFRCH9Hf94ln1QJAckOZqvFl17jM6joQjvRy2N/vEgD+SnxRAz
ppA1A46AtSDlJetxLKRLGl/Dcq5omIVI97DdYlgEgdLGsMLED7RXoh141spMUIqC
3t40GuFMbAQkdrmlhSUwlwd03ljpAsugdB8Gkqxe7OQCkHIiMQlwJgZRqCNCZlfS
XEuqevMsac6WO0n7xjzi0wr543nwpu/DMkr2A++SU5Cv6IBYgGTgYSF2xThsAxws
nxor4TdVBknSO7P+RblTKGzmqUTgrTckiKu6hbgd6+ljNb60LhxVgEl3Tu29NBpw
VrobQrEGqr6dBxH+3zJoY9b7T5E7n1GD6e1u8wXJ+1YuAV9HmomDk6M/lgQz9J7+
AxfmgnHYcDY7SJ1DYE3hFFjoQXflu193u33E3c1uxf9ubXja9Ygtit+E3ITZVjpT
+IDxh6P0y4hf4XbSIXGMzrqkLFJM2FQdOrGSQMwXxdaNq4iZJUd1Wv79XJuwXbSG
YCJ8LoP77LVq0HR1yYMs08MaJA96PimrmOs0yUran/goqFuqQL046B3BpuOfnAST
Jy3CuHuLGoFz7vZtMX6DKGqdBWpV/Exq2HeLGF2jrqORPoqkYsI9tJD4H2fd5Vun
9139Qk0hXqAhonI82BfhY4TBe6ugaGTXfYty1XqG0cICYfV6aQNM/UCGM20/8/Mw
1mbqSgZbQZPyf9mllrQez88b9MIoYW05oDxNYKFEQDNFmJoUKINmNMcVdLKM140z
nMQu/9InBX4zLfu398jiQnch9ehH/+5pn+2KqpiLgWhyG+4gy1hjbvcUHdQYbdWC
jbR5yLcdVneyf13trOFOQCmBq833O2gay1QQ6FH0K0igRNid+RRyjL10mb8uYlE1
YOvJp80JJB4YR8Jl0IVGuN7FcrR86GTDKOXHTWornhWOGzV2qJvnKEqHe7sMDp97
PovNZn+xAaIVE0D2FZ5ryzt2FSQBs5Fkpf2UxytJEqd73KieomXgOZXQCdMDmBNv
ko4Wogbl+tObFsutQamNx9777x/pnbG1A7atmfbY6cuez9bqnxjQwLof0E/o5nnL
EGOAmb2fiZQOt9JH0cQoCZiKKYA6sLc7NcYKesfYCbWOHWMJt9361iGvaXxABB/y
+UMyH1oHZV+YRULk6lshoEk6jCnXH4d/VDxq6adYiRDi3JClD0fx769RQXPX4c1E
ZXrus9sXqejduvyXlxWqmbP1LrFN+U612g04Ap2y2O/GOGCf1tb1CwftKY8pJML2
QiZJA+VzG09t6s6+qdiw9//ZdYdzvU9YW4uovSBxq2XRYg5RRwWc35sOXLPhceI8
Cr895HzLpQMuPFdzszSgCwnfFclOh7zqWMVB8pJHOzW0durFHUeFmoGl3Hefv1NG
q0wjaaZAxoSBboWmGk3yirC52pt3xx6rtUUnS9xtsbWSeqq8cMe8Jn4RbU+T7pOv
DyTVE/BZOz0O5377XLk74v7jfc0sKkZkzFIYJnC/4VbyGlUHKxaBJh4AurhYK9v+
dJFzi1oxKewutUgXH2iiRv+gGzJsCHTDl9PBksCJwrwqRrIF5ZdqIJ02BvpdPySu
ZX3P8dwTbVCRAgH0FjXDMk2hOaY82ldhrnSBB4h8eqtqB1Hmi4iAmEjz0GiXKzue
u+36WizXFdmwd4ug7HXUCP+CPmG+VdEkXi3lZcFUAbsukhMA0qsZfbl21ei+zPUq
FXZ+CKClNCKJkVNEwdKrWzSay+2eMLTb4fXNcjhS1nViOzVxSsqgRd5x5JlVYMeR
2KKqymGEVbubLRYsK0T57V7pjNtbKrJuTxgYskMKDr5hvSrIEsye0DG0cfNWjS6k
3N8/CTZ+vY8kkyDIagskJzw4FSuZbwjQYX5Qhk8eChak1N4luGszJ2P/D3ilw1u3
Tkfz0RXW4ZDH2W9E0J+2n9yOUTCFCG9Q4RYeGySywPxNJ9XBm9LpiWTuNgktlJqv
HDVRauRAqjAYMD3Z2f2Sp4lLVQllXCmBI7+XF7Dv4DRje+L3o84YKIIXmmo5PtVf
FrAk48GKyARJQ11AV/F+ZhD41CfESl0M+raRNKLGPigPaSz0Jd27PF8905hpvKz7
keXm2WOmvnjasTEvOpxI4+M9C3uOW55EuFC+cqBCpt/UpTsXg/pIkyGFtBAtrJc4
B5INSs6V/bCyz3s/6RTdtiBo80etDlOQpTRAZAophYAsX53hyWZNvObP2PAo8kc5
CExCMkiWAOU+8kINwv1BMslcpMqcv48mkdrkNK9r2tThfaO9hdvoTriyq0asd8dz
VWrvBeCooTyA1Klfr0MoXczydgSf+v8r2GOR/BRWVll0JOaQD5mt2xzGK+jYlB0V
IzccH0Gx2mubV5nJDzMcfLAmv6QdZ5gpAWZc15j8aKRgyq9y366PNLr8j71SDpul
1EsmpunsU0QxImkv3lx3t+b8VG4Cpv5ACBvLt98MCvittH+RcOhlynt7NKC1U7IS
4Znk4115eAtINKvp6w8NrGaNmvw22iUMlrnnMhzfRxrLfVl7exZERH1nYKpZAJtB
/yyun6D/Rwlls6NKZOoo1lD5V6LVAC77pj/p3liyXeCmJQZpDumbzIeCmvaazTGg
b2KUlCWbGga0FfPgx3htAPXFwiAtI3lWmSbV2GJltxmJpn8rWnT6X8u3PseGIXGS
+Wgc6W6BGEHs+D4IfiGJPNA9zpofxGAe1y2nO5sCxkgl6rQiMabaM0WHIlxux6dH
3eJH0XUgaffoqIm+4xBPtG4KmUGxAEiaK4OKR2SOOzvGspZIB4o3otmRyanhgbss
QngNd8Hwt14xEkTrRuLz0J1QF4EomPRX9CtaO7xEBFDc2jgS9XdefcVmKxTGSy/Z
gRnQuRI9YIlOTzxRVkXnoCexvGm34mKYAnOmZKKMBb6vhd+a6yTYG8+DB3c/jGZ2
wbAmnBkhT+IlV+T4Nq9IzH1JSjygYcoFd4fWKajnDoJGr6VJhqINH1gwxDJTYvyf
MX7B44ZaCek83vK1cQhjWqqGFHgLA4zgjt/6DBB/Hp1tSy9mt/NDVIMAYLcWcGr8
HiM6V6hnF9dWu/ffpzAp4//aHC/eBmhEXc9EiF2iTcDCMYQ4vGlsO93YiLq1H6tq
kBx6BR9pskyHeiOygq76KUEluN5nM92kwqTcFiNEi8BHeOTdMSRfEgArXnK0/CAh
QT/BlAoCkcTJEjYms2tPj6u/ml09NFzbdU4+lacWfpQ+2gonOqPO3l5b8b40iRoe
owHLkSf+vH8yAZT5nS25jz8DaHUjNF9YUWUfLQQLWVhxVD2ieFS3tD0Kk+TR7QSx
VfCzlJiNeBmk/tGx7XCUNT6r1IuA6qZvbl4KbkFRYsorA+lzn5eU+tvXa72vT5wg
De+g+zRC7lRlKD/e6WWrVGLzFEarSP7Qo6MyOZNF0y2RIjpCwsc6jm557sQFNXWG
5SGpPilLyuM8Zp17eitFZ+S9K7ajFheoM/FudUwi9l+YOE6dBdGeiIQVeXpZZaW3
7f0xQ5iaFGWv+Ke7xHGEzR7BtUgXjPVHg7t4Mz7QaNrJ9tFuUg5WdI440gX/BAFY
/ujif7qBRqY+U/6QlZT9G3iC1Ko5ePsdC/DYZ/J7b2GHmK9qan1WZ/0SKx0c4Jyz
E4EKls8pB1drIjCLuA+wpyMZ7GZNsbpNtHY9dwFydiHvCjw4F/PYdZF64f4rauN/
O2ZlDuCEHovD0kMWTD/KzFUC06fUsCEVAtlTozAe+X9WGbGXYDYkFTLJ9WY5GhKH
6aUYrlSJLJ36Ei/Z3QNx8T3uAPeeVx6uhXbNN0nNQ5FtqmENvLc3fPMUlfMj4BUU
v+knRNL8AcUQReyKjn4RM3AdiI2ZEeTLnhbcT9I6fab2uhKtSfzZoHhmn/nxcgGr
w4S4PWug2V83w1VBMKjg9jNajs6R4TXcFjXpOvV15ADg836B4HSrsV78S14Euvk9
HDJFDqwexdyVPecQOsyCgQeY3UImB/KRqxr4TfPz209iOjvLrOUuKdfnYHTKL3Z9
DPXEHdzQUPDL3F4SjIqXgmA4su3vnVg3hSJuscl3v4lKRUXSb97Tx+P6SSqgRfLM
9KODpgCgchdkoMbFVWgakNRxZ0aRAL7Rd+ep5vTE27c0hShUapzJM6wSwOKIY/1z
KGoxWh6MgG6woDscCs22fJhT+/wIx8DEymL7cXhOEEwkyiDsOaEofIKSPbsL7qaU
ADbqMnnFHjLhbish/9Al8bxgOtVqRKTOJDHdhytxdxVCe5jmE0J1lkQcFWjVksGd
tNGxvDgNVZeWMfJ1l2eYCJxcmpCGWePIFYq60pG5xN/uFAhSHzAaxlTzlHfy2R3g
lAnNm1ZZm3eCR76KUO2Wb1TjRGuya+phpuXrfE3qTbEhJyLoBYij/WhUCFxvWA8o
LflOk4K8z6y/PERESxzXoTwfSTlR8TldBl1yJQpw120AiawtweopYQJCTipbM7CP
zefDN5ehNbp8LX0CbcmpxrfAUF9Yo2rsZFYdW7C2UOD34cWhwzCSSi3F+ChePRUC
g/ZHipURAHI7dlEsGI9rcTalrVp+WOCt7rsR001Fhk96mvM4IcGjUGrEOd3guHUo
HwjMgaidbqNInQQXJJpwAuX0Wf+Ry5igbLxJstZQtnRiVbxgliroTgQeO+UsK1Jg
++9cHEOJHwvCM0HClcwn/RkJ2j6JDVCfqb41KTV7ucCo6tQm6pVJs5tcOGhtEBtt
lWkcmWtjIVf8yBnY8mkgYkoMYT+z0UTpogVWsBNqVgU62gvmRlI3hyWKsiQpyljA
rudrrO516dWmakXB+zLH8qh+ZV0HtJ8daOcN2ue8sQ10owIEH39gKI7OBv9lktOf
7eOcbdfRGvyoX81We5lrl9NvPXOMyFpsGUUX8iGo4zyW0+0jewJj5ncjMWTuAkIb
QZBf90D3erZRR4uSm914FrvSKORGytkaQViUm/gpWAPZZmmWT4tUSHjGINtQpZmB
H3bDlH71Aqf2jcSIT3Ltlnu4sd0WW0w0SByBBoH8XKMocYk8uzSmuc2u3Xk9eirj
9H9WiPJov9peKLYedJ0vCEzXd39gFi45ETXbNMmJqnOPyBzzsv8FtWqzedp5Xboi
QsVahrG55r9XAnASFdV8jIoasIwWuov8XW94yLij3dghdtfJCfRf1S0BpwYT1QgS
sDDJOOWAm8GbpSR3wIE/gzmG8cy6GdWvMGg6Lstuu220yFccIyCX110EcbRUFvrg
QtefGqY5PU0wBVp5+pssHTlQURwsplXRPSYuDwfN0WrZEj16ocQC60UeaGeb9Gvk
/o0rtahfEgp4pTxgQ/TaxDbm+sMCVvbifVCvj5Jf5DbfW4wi8CHl85aredx5CD98
ZTv/DUPlMe1aCNU/Js1I4HqfPmN6/V5J0bWgaL0kpxI4ycc0KNx2Wo00lDzNXJd4
FZRy9WOoGDbYizeFPVctPk9RhcXiH0lCFv2tBFt4sUK4jb0NpXJq4RPXWKwiyK9Q
kFQqBnbJWjoBPRCVTqmpPRl8JyHPJ3wqJFN4Z5B0FsKiAdPCIiHvTRM3a2K0oajh
OJJxBUAxlNw/MHlaOHEVV2KxT9RYszGZKGcxPi+MHnfUC0Oi6VHiSLQdq3cMl9Dx
aMhwx9SFx/TbhiLpnOZ423jF7a0RRV8L/q+EpqXWHlSkwxc+UqV7nuynlJIMcjnA
qqW33iClm+5+pWwpOtM1hPn3Og1Eb2e+9yimS8EWHUcvFlx2CulyxpQA+adDdLVQ
jquSITG0xOW4ZAb522a6wVPiL2rSQS6wlLWKZXD39Jbt6t77EH4/NMFCwUUuyWfO
ju53CccG2IMhJkuQoEkGN2tvZNMhkCNLOBpiMCafVAVuIUo6qInty8MxQ6q+XAbx
R4vgDt14qYM1PiliwNXnSbZiuPUGVUlX9Mjz6snA7sIKfiaE6aoC8acvd5adqpki
e9px5L97tTyLWYSb/1BNiup9y8L5qbil4SS7+EmaTZuFqFpaZspO297x2Tl0Noyg
hNyu07QMwXMGxP1IOxeRDY26gldY7tXJouIIxBPZqtBiE868qBSfYi1ue3HpGOlU
T7vpUNYSIftG0sXJvfOWyb/29rp2ICvAqydqDg2Ecsp7kDOQuA9Kyj41rutfkWx+
HHuRUUWw15jpmGW2jf31OHxmDRkClUFIA1xJ6ImvZPBD/03v1vfeQnB4akpiMN7m
5RV3kPa/LfXHoRXFZRygyoZ4L1h9lb3BTZ0U44pP+mkWTvWMTWw7ym30wS0tgx/k
VS8C0gGL5PASd0/ATcZ0kGyEGxDctglNJLuAs/Z70RuZplMD5QQHEyw0fFKRwLdU
Ch5W7ebrcnDTBxh8FOf04+rJFktoCq7p27hHS1chPlII4cJ5Eh6q09/ODBD1CadT
FHKfNg70PywHJkVHQZQGhB30CbZomqVcuQD1EtILqHIsDNwVJTa/RiHkgNXUcRcx
DP7q7XYOcAG1Cg6xFAFu3BAHUGCE66id1KuwbEdC1CsB7mOUyLoMJtct0PI0o0bk
4ntSw35g4Er+9Lk78WD5KjcqNy5SsbMXv1X1LQ6RzcjDG9CARMIlIctzxvhg03Oe
jzAC0gDQpJMO79fAX/iDPidv4PbUkiPDDotsDOJ0yViWMECttYIE40TP/CsNI2pr
Oganxu0A46eiDbI3aPYo2nhKb75wyatc2xSE/F7pQ0tKzuKVAsYUCxxseUXVyFbA
x9oqXgMU1mKwwA1QX9eEjC1PHQvUMj90AOMDYOXDoeBnH7w/mkdIIOnjmbMPP79h
3ocnu8DwOaz/ZePbCsz6DL+8c4rydPCEkCCRUBxVuLqmk1Qb1/MpeACnmwAnfdHO
jmndD8B57TguAwTE4c5gfg6avpg5bpzDVjpLxDOHkginE6AjLFD4ish2TH/lXV92
zs6S2iDuSweco9PWY2CPY+juUSFuQjM1H3D50+leOMjMvvHbK2mVnuDZFCLw7Zo5
BUv77WFGuddT+YOeHXZZ9scMRtEB3kXcvBVN8KlhN5V60Vg8p3ndg2nYyxkzdPsv
tXOnBSIWFVTyGBJgdgCYXVh/Ru4v7rvuKvSBW9lClhBX+ijm0YAdxf/UbX4Na3KN
Z8IGczLcjloDcB3sibcQ0Or9QQPFKyTXL52idQVkoqnQ6wZg5Z6I6hkFt7crvVI+
ltVwcCCDuUPAolJ2EwYAA34ajZ6bllA5K66oJyXDMgoT1CGGQVBnmPV8R9H8xbeG
FdHonjrd3P2djw9qf+0GaPoq9HES2TrtPOyA+vvmpqrJlvQqFk07xAyjBKC+vZ0I
XIvW0BlvAtgX9upqQBNSI+ScjnNFM2wGTGaKqvezWe7CyfoVwsDYK2flAoc9I4hG
jBUdm+343/S6e2PSgEpsBUWC9T6ByzVxjykDJOnnn1UpvoPlSi8AMkGz58lsu2nd
v3vi6prhcF+Dte5eDs3ypj1eEZETEn7rteDjK93abxWsqTw6vlRUly02Odo84gnU
Q1Uywr+jnwJHW1uE9+2Z3VZEFRO2Sh2o46xPNcqTHw3OzrdTQFNTSoCBzlq7TAKI
dG2DapqBd89R3PrloLLfUkr0tkDdwrNP/6RTqa26mQisi6hnT5fXmlChF8VjtGM4
nnvLQJ+GWIz2CQ066UtA0WMDnByPzyKZ2jC+yn/aU4BBAddZ1bF2zXR8GxdFzfYf
Wggg7Emsq2k7959anwseSP53tDszss4D0kLNouNocaog1RbIe38a+U5G9B32iP2T
y8jen5XhEx9EbP7J0dFG10yLO4e/fKmQ8C8xuuFUXuCu7+lhrCvR5W8AdL+7/vRL
1Pwla+aQ1Z5F6vEWICnUmycj/r4plZLZmKrrldchTCHfRYKuaxuGMX0euu43N6Uw
DwPd3jKJssUfJzo/3g23yDfn4aFtFAbs6X+PFLHbxXxvL1wJOhENfDRXQFHIR67k
gJEvNf8sng2oh/DYFIrLsl8WvgozK/7Vs4xrihJGKmRWbUvtbJWANAMPr7YaxtDd
liQMjGjJl7iyN8KJjyJlDPE6m/1fb8s4Fz2IhOWzZ3Xoo7F1YjUjU1WDr1QM75OT
G2cQEjnX/PuQD1cvK72WTX6zStG6CtZ2dQELZFsTHIqzAyVDEp3HLf/KZo10IenK
SG9EeRXrbXcaX8FAoqTMYpNROh//sgTo499qviVr4iub7AayT6Q7yS7Qnr+Q6pZM
/JskTT/LsmH869LgYK0Z8382L75Ld6jlKs4FTlncuHwHUx/KAGqUIzW5Jmh7C7ZN
dkCj8kTjRh7oN0bWaEM0sU9t5jECqifMGsg3bAXtRpnUgHfyD2kKd9dKMRNsZOwo
MzgBvb/1Q08J9FVtlcPXpiKQRt0NLXhs2v1Tugf6I5SLW9v/zytJJi4q+BLS3QgT
JqHNJgOVwlOIwo6M4BysZ61dpV/7LkoC7yiAlJiJMDXp5GjfEagMreA11NKYjaTa
dS65vgukipoAUXF4zlFrwUyjpS4kElIF2avZM5n6DctsiKdArsRN9awxsxtMFpoE
SXDKPsBNTn1O/T1uid6rHwblioOq76mJYlSYiHBX4Pcopmk7uBji93W/mylu77+X
iQ77dGmKgxO8N1q0dT2LkHXnOGXcFwlhFhsJyPxv95VVwprfer68teg+3o/tz6F+
V3+UnfZ6hZk1j6+zbnFteSHuEwW+9gYI9cgXCajeFWQkCGKlxcezlXMQ6SnxtCpm
3OfxUGBhEjpMKXiWCDN4bqy4jN2Uk0W2a9pq9s2fzVaoDJTvSWJiZyIDu54SSGsk
Ou+MuVUpTe9lAKOPQ+EKcHmWtAOVUOnksvh3THwemCSf/+xeqZDBzhdqk8/UI1mu
a9R6OnRttqywb5BrUQTc6bXcu4GyoCsGGIYpHDY5NSYHSzUcxfSqt4dkVVT7zI68
m/fJ3t4QFq+wA5+LgRXcejRhWSytKi1UJhR+oCijClwsZixHtlxHJ+YJqq0UIZJx
7erEyQ5yZ0G+PUfBjZ58LQ4/E8BPiwklgmdU7HGDP9Z8RYClJQLmpzENasSoM/UR
PuARO+CvuFzkUXRjSN7MsevObP8ExmYJqEyanMiC4f2WlA1q0+UYWMzW+arQWfky
dqtO/X+Pz1oP0zIoXcZpdX9pg4Eq4d3iSiZxVqx8kbs8XEQxkbsoZIgQZ8jJ21d6
Deo5jnUt4IWili/993uaQZVhwCqIOpiFl5ke4y/Us/dXo7+ENfVGheazj20TH4ax
odiVeR7AwHUC6gEHNY4DtO1lu4VQJRj1PUHFpBNwXRUKKv3ZQRxbLwyPATKatnDE
8DjTs6edqAkYHtRWyIBjyAWB8TlkzDX0nEcx3XpaHUYtGQagE6c0OyR/nGFh5N5G
KtoUv1XGTbgnSPzbZpDuBJ0XVF6OafvlvozqnVqQamk69rAEJD0kdpjjqtAA8FQY
5Y1OwkT6eBQslw5LpGNs/UW+EaTCRkrKyV3IA+nkfIvnhuOVb091XNSNHyvJPNVW
iONT3tYau1zRiV29F2PyDqtV0g+KwU8hzpZAYzwelB2wL8jwgiChRJ04LQhMaN4V
AMjRH2bZVYPIhOlYMPFAErwpzf2NVNlAt+x63CC57F0Sfv6cZLvbXUVxyAYqbIzF
lf/VKzNiVS9l4LRrdBtKZrNQcBh6NY+gg8fc5eYueAyb7sINnZl38vG6EKXHNyiX
goqA1959jVvhPlXBwzESwpovSSfg9cI6kRs1G5klQlD0YCs/E/GTfUeRGp5UI4ZV
ypU7jfY9LTuwL0FDfqR24fLd6fyC8Bofa8mKfwzrLumsIrBzH+c6AkB3OVLc/qa5
TmwV82DBRmvgeoGdhyDGuLsauiaKqE+zx1xODbO7uAnwQ8UJ1XiTRs6bmV8Xdg1L
/fuPS3Is61eI9MX2vZkW8mraFH4fkCcI3OnZ5gYtECNDa87oQkGsvvCRC7ONMo6U
guD2mib3wiOFrstLDQVVieSvI3A9K5QwuYgvM+LAbZwCWDS4fA0d1obW8X2wKXFF
LMre5d/4EwEKn274ualHkypYP7VWIaYdFmuldr7dKl7GoITNtcETSTvG+jKLgzbt
mUPhJ8ZTd+vubn5qs10/i2vvJN9muJghDBb903hBE+zs2P7r0k4oR5JQwkxG63o8
KRQXO26AhLd9n5xe/RF4ACE1M59+jIibty8OORYYvcGm0CaF/e8ZuInml58vZ635
RQcaJKm0LE8qhXaB+hyX+yniI6CuxAPnp3bvUXKFBkgat1lwYPDc7ktXCuBNrcOP
sVv4E1t1uvUPE9ISqJP+7bN1ya0A/EQSbtDZXzWUV8JIMjwdxZWMXQBjd9TCRyp0
BOOkQCyw94tfmxhLLy7qusXrgvlaUKrw4AQ+jOHLJH7bU4EYLjQl5DiUlGLgj0Lz
mXYhWngXeo/MXPkQA5GIctORkNB+DAcdP0x8Fuln982GEJlqxmNkfTLd7eOyw3tB
lih/Fg3HssI6IMpqTcSr7MutNR3YBcmfcxkMNpadVA2ln8AGCrEnt9rYmpqf8ehu
2n/HmL2JSDBSqfFmqcj5OjFdKHKYuOn+6+0Mgd2D89M2pf9AndQZaClB/jRK7BEY
8P+JHKHIkYy9pCK1IUXG5Ubd1iGRjkXGoY8fcxOQdDshltU+VMD/KCaXYR4M3ctK
1fkuvNMr4lYy/NHMGSfi0QZ+iGM/cODqZYX7BlXoAAqTSf740eOG+ODIijMmLE0G
CD/3ya5By7Dq2aZaJbInAdKDNLHmkkvT8HwwRzAt2t9VVgIZsTf22M091gbQChJ4
wX2uPksxlQlVX5yP6KfUnfhdLP0LyiUBlIdwqrX640sMtqO24+LwRHEwZXrt3/Bq
ephFtSkEbeeDBTi54c5f7KNZR7RDnH6f4tGSAedTSwUZROCqmf4fg/PUDzIM7GH1
3679EMdKXq6wvO5bJZjqVLi9qceFeeJtU7NSvFcWURPs5IRR8fpbKVGwFLFEM49p
+/npRoqa8fKMLEd1WE81ZzWECQ1JLxbi312H0YrkSdnaAfKduk1CWsBpbayjwBD3
GoR9I0a4vPn8DKSdsg7eM7TVja38RRpxd3w3bBDNo/eFHQrJZVW02kPbHEekOywm
qzd4kuzKa40XC/cc7eur7+BU7Kk3MfyzzOKjt2QaHi9CUiQJu1w9lxqMilg5KoqP
FJmX6fsFRIzov9rAAgezsCSuE+MdXgAfpFm2lpPGMhozs3UynFL6JbxfGqDdJ/Mi
yRr/xw0Vp2XOMLzCYRckLu2IsfkbuA5Qhbh1HX/eRsRb1ynE7ibynxA3MqlFpb6W
bCdQ2AFwGV//TCPsZq1Qb0/UnFXM7QViMO72+4/fvNkUbksf4X64RUVVpyK3UXIn
AJIq6QWdsDsbmkQQ/S4RAG41/AQEcuDWxHnoPeVYpukvO2eBvxWU3WnOXkCutSfK
zMKVOF8jLdSDyahEdgrf4pZ0uBwmHu5pkUElMEBfEUqmK1NU7SgWdE5UUwmijrDe
HgVh7jd0idvRGZLCFIgDT8mkowzKLhuj2uJza8y7SslXxeh6UX585PWvzCJfGO9L
G/hFNguSUANAa0JF4IZjv2fLS+N2I4HetW3WZRL2Qu0hfw2OSz/rNAMoCUfBf0b8
26S9T4gxPUMPACDjLwoNUcd9H4+rJVNjTaJqvBuJHNZrY92sLhDrG2EdvKq3e8bz
WIYqNSwXEBtuUE6y6RPxzh5pdZH0jzp7pvBhuIrmGEZgEieQcZ5oplupXpVWVxBq
Fqtp1AjzTPOM6lEUDMjYG/qsIMIFn3BT11D1rXGd2oO++j/u1c+PKRiw9BuHK53X
M4E3srbLYLzlLzq6koAzGNrSuejbGwKBaJzVyAh9sjda4NBHDV5foeKl/VR3gYlQ
yF0Ed3KQye570V88DwmwT8eOOMWKlMVTKGHwvdn9FcdF9t4jD0Mb5BcZoIbKFjSy
m48alV9YUr1Nprc2x3/u1rSCwU4iFjFVKbKwDV8mGdl9UAALbB1gahdpfM9ZiKKf
agbEytplz7T5Tq4OFStwTshXKfHzOWQ57AetN83Z3vH4Og+MS5BVY6q0/iKEc6Eo
HQyECd1kSvKC6TGeb65881WzmRPgu5ftzfazG79WkKiwqNoGoOa0jGAJtpHONXoD
DUIpG/CsbCiUuSLFTGJcs58lryxlULM3dKDG3KR55my6AalXyupcxF92yHr9ui1m
WcI6+DJekK/V0ZJg4frUc1a53jVaEzDk8j9qfeiMAf/zYEcao1E1aBDgiMiVvVj8
A3DoZD/xjFPlQI/FhVB6qyiUE47FqNzUlzzYwPXuRDwXt4vSBjnOW8GwR4F/P9H3
6M5rkkBrhPjwFMNDyu1NZTeYlghd6cMrcl0HOowR4YHHmLpT09/DHSSUpplEHbcD
d/1WgsGclQlhqmx4kslqIBsJHJWuRrr0JW6rP+KeRmFfIIrCJds90yD+QmBKSg4s
lpjaSTKyTd+eKavSHjlv8Xn4C38AYmGBuHyEuCbeCpY+1/MW7xPWDeMQMaLTk7z0
DCgtkCUCRfwu+6vmnrtlmRE2Tuu/LUy8SDJtWV8NGrL1CmV70LNWEU8hwQHPqazv
a2pwt6oeaLzuMyAclpo9F4hoXonMeeRJ0iElxWbbB5ISoBX2iYKHZRA8gbFMeoUC
1sdocCsaDgFSvsf6vSmDBUHss4DLt+0MU5o7Li/IdTvUO+4lWf+YHaZrZV40SHTy
0CyzaREKZw5qNxrFW8z8f7OvLlnYFzH3kRzkwxDub7NtQLZJ8E8GLr+u7mETkGO3
NhhfHSFq/mI81kUw8UiF850M714ZjD3GvJNu1dg1esFsty9MIEN0gYN5zrIs6Ax2
gG0NzenwWVXArT5BOmzr6aDT+U8KZSeFkKT5LigCkd0dQHsKkB4W0+3yp0LiL4Gy
GKaKBcqRGliQkQkETdhnv9bvhHzUUg0U4qdW2qUNR+qcbLdM1oZcrPquFDY2r7d2
xJhShV1AO07/qyKFrjxgBvxNnZ67CQiZSHL24cmO0yDIws2+AxFmlG+R47NRd2Co
UrWxr5X/b3I5b9Id9sy9JG6QbSNNhf8H/iAZS8C1323Rso/mbqf6yM7lE8art/oe
5IIJ4ouh2h+KqyKVW3kK/mtRBaQbMkUsZluGvgFRbndBjK4rbJUz78Gur+9nKqTQ
CtY1l+uJ4Ppo/npzrrVQ6Gbc0rAs9A1WZlkYovViZIfLUt76oeWsSZ4arrN3jAun
CJtoWdgN9GX0uxYaonU8vJJFL3O7kx3RNnzby1PaBHYwEP/HtuJZyHGkPL8drFOW
Hkp0rge03cinyUG6h8Rz7GCghYvMONeNA9Kz3+2LQvcTWt1QM6FxKpfUJrVZK7H1
nVtxLCCrmwciNc/AJSoiAwltPiNCChA2gxfuvR7hV57pvCW+aIGjEGSa8NVYeQeB
9vSBdqjp8IvqaqRhSFQ9p/+Yjz83N4zBW1XdDpQufiEEqzU2Fq+RuqdwXiRifVNV
iBTJ7uHnkbVGCi+wjHeTiD3MQMyfnrPUgRJjquBRFryX1uIhRG6Ink7lIJtPB6Wm
1JNKkOgGxLKXtxVUkw4oGvjEoE7hw9sWp6HDAdGiXNLI/NlQF9LSnewMKwyxcnj7
6vpwN0cxAXwk6chw558di26QpNPX59dOO1csfuB3OwZZyZB0PvJb3ksqBF7MWxrg
KAr6HjR98h46Tg06FfnEkx02bdm2jlFeMrkHrTZe++Nw/tnYYPBPbsjIZHNyQ4a8
Vyidnx+88pmg6CDlFwuTgB1oKd1qAS9+Exmu6RgZ7IClBt/qGyhcB7OFtjC8Mapg
5/qgn97gJc9DioIvlnHu/ZgYG7TWrImkd3wPbD5uRmev9OQar41q3mNi2U+KQ27v
zxXcBxY4nG0+rr2jsbaSQnKFVHNItZcVJMCVuVpuCvzr3g4vOgbkI/tzx5xdMcOg
Kd6BUwCByyHyR0mjVUFshJDnq62txFFgwQMLzrDQk91kLouAH1bXLUXu5rJ4jFxY
gLl7+Ah5e1wXCuuhsZOr9kW26vD572hcjVTIla6KDmDTOwX4HgxlQS1cKWOIX4LN
Doucxft/cXdGkyRzpez5Ukjwki9v4166jGVPO3/2bXjVkwyJ8czc02HYyXje3zfR
z47TY/mWLWfAi2bi+LZ7ESk3Q4odYU8EzHAuA4cKBibjawhQCVwypZ5AWs1V22Ky
jjP6A6hOERAQ6z0Zh/q9bJaNV1yIAGaIz8rbgCKxne6CdiiT6SnmzWcf1/JWuSy0
IlgdLqHnm2F1AaPIOVkvL4aTChrMuo0ifmUKBJkbUwFJnKMv52GE/9QCXCbgTEfs
cO1boOAdcM3cvwU3UxukEO2KRSFMJgVk37Q+Ori+ueJhQ5HfFwohjljfkiB56e6V
GP3Tb8yhkTK4SWjT+ACfYFWD+CIWRiJNAPLm38uO2JXmPSyPcY1QH/WBatIe7aer
hUgryeKTsGIhXmMUeXD5NPzgoMggfBVgS3n6eyyYHF8LKRQyG6Cd3H3xmDzV3lr1
4+h1uk90QzHaJVV3eeL4RMvxvI6kuP12cU/W5qAlnpMrpKLJwmBAn5Fqyvvsfbyj
bdn0As0bTzlmf/luw+cPzpAkmnMNAq5Q29P0R4AJu2S5KYRkas9CWgDX9wn9C1tM
AJoet2iBjzaJOU+Ar76LR3m+tAMHD/TTAe3uFm8JHlbEE1H3o07suJdDt8ORaU1V
coouCbufKcGYPQoMKaNZRsgl8fVPWKmgeqmcQ92TOerCibde7lnF6aZtQYbDiH+B
UTSGlryr3PrFuqCP21QBlf8OmhCLZ7mdAMBxtCRA0XsVexL5M29XatIwksc0Cwvj
HW6WuZM/fyK5Vgb8LMy/u2H6bZ6/xQLPMHvSLp7ZZfePllKSgKNdUdwY1bNJu8qE
2wKj8QbkyMV8HWtIF3uwylN+4kR6t3v70lrisWtrCuaMnp0QmsvDTOwlXSmK/Hsc
9CyjaOpEES/EsfpJmlkNwfxxY+lP/e0LtE7taq71sS0nrV1kdEDKXPkLExIcgDzE
UCvlSwLVhdKcbrn1t78hnbMcP0F3CirIpAtpf+EJE1w1FwBTk++glYo1ObcqQ0BP
NgkBFlR7HQ0yMrWZhQIS/DQMeMtS//X8LMZIoYhbImVkC7iLaqowoJ9wP+zifToz
WEsREARByNjxh/LcGHJj43v0ajDCN6HNH66XBQjr5rGY4flbQ27h85iF7im0F7AJ
pgZOcDE189aCnybG86zh07PzbM1jNjVcOw7ZdkajogW70JCU2Z8jrBC6P4aMxDlf
ebQeCK6uxxoZzAFvXONVuGLfDqCCyyMb5XVuQtK42rEN6D1CDiWqwWFePgIwaivO
7ES1dm19AmbqpsYoRn/8FJxgzKZWIGtU2uD8hxK7sZHvpxfAgN5/5QzUXRrSw8ia
i8GuRN0+mEOZFPJr6qX+LXamXDC71Mou1eCZhZHzrPufgbwslF1Pebwy9STHCOPL
b4pDlzDbNsVSJTdvhImNfZKFBOo54Cs1fOkv5yMOfxE0WTxsuy+dcM+HCIF9kmhm
e3ni6K+r/T4ghdvxrTbUw2IeT6xcryD2Z5EGm7pmwdJwKQiaN7BxVrgv5pf97Jyi
2iMjwB0G/0dAtns5tLEkKO6mrybmN49TV3HMHX5JOjj371tRcYmwYFIplRBAoEl/
6bHnsTMYwFQx6gz4MUnpdwFFrHB/sxY+lvvvuqyDc3nGklqtCwc5e8+L/sdWXwFd
AvUro9bqqPGQsCWvjEqBoxEXRmwpnjWLJDFjbvi6AhFRvBI1/1w9kGORbdTPzvB3
dIuZozyHUQSJowKct0Kw0Ylr6W1u88ZwuZGlyIb69f+paSWxId3rfblSZsooFTNy
BdM1FG4cQecUhl30QedSKyqu6er8gFRCUvJwp3Q1ZUaeelzlPKbRhgl8GboQkz0X
1KRKZ26t/nwdTtyJ3eBm7LdDGfBVRVkWs0udwUcnCnXqwr2Ddpqofv9Rrn/OX+hv
oBt9C20B7SmDkM1wY4kcxpWSli52vdlDNB2RdWlye0GcjCwZSP3IFTVOqCY3T1rp
mBihDGrjXQJabt9BaMQr5vX8/rzjgQZcECa/0J5OO+HP1FXPuwdZyJgoYBeRW0a/
+z87Va3Z2lus5mkzpdyfq/dGa4i70WUE0RtlebqeUVSg9jxw+ovIO5kqtUtYb/P9
MIQ1NhfBS6W1tdGOhuX3TKgkTHiNK5l61cnkqg/IjQRpibG6PnyWKTSR+wUnjF9a
KCxqAa5UWBqPSPGJBldrNarsS27+NltCrSevL/LpDgErGCoxPl57+IauBuY/TETp
wMnXex+1Yz4qsqvpgDDK3gAHmE7BYdkodBvXAd5tsCA4qEIECw8vu8LxmB6s4vpG
psBaUgpbAgLzBjTL77OZ/bX7mzc2BhxBqMiXIul7bLgmVMKSSi1HKfBGepxPDeq9
KNu9nnzaQU+1ZpoTL5OV9GWWP39gaLZVF3o8Es+ljEv2b1uit11le93KtmNBAAJu
YX2EaD1rkYr7wjqZc/QsDYnZGYICsIgc9FD6ZFTwgA86zxjPdnCwrzdmDBkBgpJm
2minUg3E78GfqIZco3SxW6UBzLFEFCLlTl+XFB/JPRWKHGSz2NEHy4x/0SoS0LWJ
Sqm2dT+93GlAKAODNYs+7UfgZ1Gzi1yH37de4AfiZSLVoNfSKYoQ5NE15kVQaj6S
tWk5xYLGLdFQxV7rf9dhbOkvSmugFFqiUuXpm5zJZTG5ZyZ/wsscakWU1hJTn77T
QN1n7FoyTo/ctYoW457tLP6iqfH7GM0DKsnQvRYjsT3rZpiS7jXcMj80k4nuLwmR
+RgtZuSktztmG5FOjHg4B2ifkPtgOFfYAu7qg6uvzHe/0G10zv0d+3Pcg8einy1K
NYyTHaFbNUvLwehWB4MOHfb63TsdmekUKZAmn68+NCT3hRKD3YD2oILdD0wd+XKP
AB38uKncexr52dMJouMMMfu3FBMiCm6QV7evoXUYKy68xqgBnHGaK239N4L+v9bi
THHWUVKry20uQ0Ecm8nf6WMTe6siuEi0NoLvmU3ihfYM+utW6foj2skLOyPsFBIZ
3/HHj6MUnUektahuMxUQ6WV4TXsRTSow5XLmuPlHYP3a3PDe7Z8J7uFsG+9+N4gW
39PiZjYZ0Ik/wedw8Yv3TPj5wGq5EGcnXP2S5r78eI3wapN6mPbaNoclx43C8aDJ
tu/HrapUI3cIOk641VTLDOYLa2MDfRkeOg0PQ603w1+flYKOgAAUtQ/URif8irD/
aY2vaabXQlRRFkpRrHTuz4ZiOc2CZbZYmGmi8iINv1EQVzqqb3Ndyc0tsK7RhS+f
oYkmKnXiFmk1sBiVS7PKcpEYexnevMDYSNzp8qWtCaKcPcons59asG5fMBR4qm7E
tzqBR3RNEwKoxZIEBEvpqLzZAMjuy770p4KQiFHUL7bopfIBCDVkZ08ph+AqK4c8
vkc2vaNLve1CTxgDwneHlPBrOZ9KzVOW09Rd/9IFFfjmtZkuuL0YC6GnW7Dmoxho
b+pgfGdcF0CrH5T5xURnJHpsQlHV1zivV1vFMKl6Jfs1rpz8H8vdSe9OvNSoS1i7
rRsYcrNBP6GcKaVzqIClWG38InpMfUtGQLfo2ilVJOEv8fBx3LExaSQ34BNVa4T2
Du3cMOqWNAIujbrzCn8Bxcx5k4RwRNrdQQMF/0lN2CgXzhgF0eyITnuvn46bsJ/i
iqivsv/AqPehY7E8pVVGoX0BG3Lf2eNMSzK1/+XWsrqCf0z8bcPAJkRub1y8NiIl
bnBmOLmPwkpcIOPZPTYG3ldGWWeqoO24C0/8zcz7eg3dIrimi/zVfHuz/yAkA8Zj
BLTZ7DQLFUKVBSWiJHY4oBwWDzVBzPs7X4NYDFt10f3mYMn7e866ZOVQUhb+c7yh
7zY/FvcGf1I5xC6ZgR4hBHtGKWt1RKmcVlOi6h9CRO6tiGQy+Taoy9X9mLDpm/xk
iWijYvkywPVPAj1aC23j428gwXDRI+CInDDeP5+tmp7PnOAE+oHY6U/JDk7tS8SW
+vzQHUrrGFK/aHIhH9mnGztiOYlMyA8ayyGckR1hGho6GKbT86JuOAj1Z6E3HRdu
dbzvRhGGqcTm7WtOsZ0e9tVcTp6vHfz0wxZ87Exq7dsk+uz11r88ppfWfAlhbzpo
xFnJ5WRTM7UKhXKJYAneq5uFS7O6foPQVFtAN0wfBLs/bV80i0fAuNNlz7NQxn4a
KmIKyLoDLIdPoMQlpqq0NsPCE1WAOT3pH5tQtTd30oE16pIFk3TnnZEn5kLN+f+b
DpN+MWf7IRGKrAZJE6vfteq729KV0jtfyBrrtjwX98GZIUecwl3aLD3Otn9cYs16
0/vGhQkSX7p0W8O1NZQ4m24nkCQroWc/lG3R7gMSIsHXF01CogE+EGBYfJ7mdY2r
QVSSZ8OTLfw4x/1YLCWGtZ97Dij+JCmdjEmWS+GqXC0R9qD6s7gKHo1MUSMMIxDb
9MNIWTrnvCFzzY/SMXYGdeYwOxr2aQ6HQgNCo8TOb9V2weSXn2jq0n+lzeGzXkd7
y8q5pyo59mkCun+Vxj4Zj8segdVl8R0DCZTJ8KDbi/S+rzVhAYXro+8d74zEtDBs
jK5Ii5QuZmbKgix6ym9Xh1VvPlQWHLKFXEZ5GhDGhtfFBmXRSpekLgEp3D33i+da
A/O4GQ9mqRTVGJ8tNvzH8PoKgYlNnEkfY+a23JYEt4+8oNVd7KTaZlS/tirHKngm
iLPhlhlj+4MtZFtzrdLt9w9rrVc/w/84CYPBSWnXtJdcErDj8lIqo5de/4Fol11V
EJkf3Vl/u+bY8kVLGKhq3xKEoGePEZMUFVS+NoIWMofrTHdRy1L8DLzCEY3jHgJu
kjqxFl7WmfQaoP9HcrdUnoVVlwwMQyYyF8lBsfnXvJAHPKPe9N4x9iAsKcn2D66N
cCKA6jLN+IRHj9WerfhitrMAhWMxCSvTXWe4BASjnDX1BcChnrff19+zblbA9yIR
+QBNN8JMqepAYNdx5BxdFZTnBk+w8kSbatbSzjx3xfykfq/+7hV0/VdKH2yk093G
SrgCDLlM86Vbbq5J2lTGM8ebB9bc8yXjOcx2Wb5JjOpdFbi25V1Do9QP2oItvtML
LMxcEg1UyyFDqE1BuS+ljqmqI4XWSKB/zi9itAj2lGsh/ZYtnZ+iuyt2T83bdvlM
4yDNVnDfjiYGeWCso6UpKqgZgWVEAkueT6UZGuDU9fnP+/9I04nDIV+gDG42kuu+
2cppJjvMW1/9XEZu5Zo2idH7WonKSKPr3IB5xaQFpoFwTO2F+6cdwVCqKNp8aW+P
kp5UO/06K4hWgg/6V283kQwO1CvjUeoB7nBjl2JSApcnp/9Te7Xx81yb4AET5Zto
M2QTI3aoy4xiiv8zbdCJ/sqEEaanvL3G9LhDI0WNA+ZGUFyjHYg5I4j4YFUJl79p
nHn4u99CD/ZCUcZO1ZCJ42eA5GSeByQB+bxMNYyvi7EjzIEb32QfctJuSrtaIEfX
Y3HgRlt9fjd1t0DyQBOiiAbxLN5VGe1TDDyfXmaC5r0OzkUMqF2RIwyPeCun/cPP
K0a4FixLy4G192oecKHtn04TKvjbOSWkqgVW5XN9qsDuwtPzGMy1HJIn/vCsnbEL
rI2Iz4BCC4zS1RqRE9RJoMJ1nhM571krJ1tDRcvwHgVpbNuJcYzSFmM05Vw8jhAF
OlRgmtpspHoq74sOoYuTJZgqEC56q4eVMB6ReWiZlNz8PO7mJGTnZsolctfQJDzi
RnZZ81Q0EguLOH+QTRcpIZB21SgC9J/Y/FMFqC1DLkClSZmF0tZ4+8rTcl+mUYiC
SDQGKbSh1gz3pmywl4Y7eOTCn4ccpO+rp0yiRCxumgiSAGZgNLZ0C9f3WQWw68Ww
OhpkRgY4GHyAKSEeLOxVwqVWhsiO9S51Anc+bQWrCvOLAhtQWVy4cDwkqEmFdBT1
e9UawBU8D30y2R8GISYvOUACECunX+ep4dr46VPGQA/egV4U5vBlzYzV+IDZXeeg
Ob9J7k7rLzvJonmWRwFuVv38rtn+EzfzkHvrx2Rktf6ospCckTl0875ZYg37BZZb
25NdWIlZ2aKnWXh2kpj0vrhWY14YqkzEyPrLH43lmZTph8jANbw4drUn3C0Y+/48
WZXuJ0OqpMlx7ENLTiegmtxS8CvLB8zXLs+vk7b17NT4Ey2vxccFbOHp3A8MmbcQ
niTBsM5Rj0NYQmP+v4cwgjzTrh7EPZgZc8sG+eyqodG90htPxjlVcNdQdFSwSLzj
7Bl9NLtZJg3sArNIfhnZK2Xwpu/X025KiFIdR72nPwbU64fGeFD1DTUAUaM6a84w
SAc++Z8uRFgu3eIzJiHFlUM+GsJp6sLTfBvrA+5o2fLuYJKLkKBXYf4oJI22MlCc
aHg3oCW77uQpRsYrGotMqAJnYR7qlch48lUS6Vbub7MYy8vqUlmYW+8nra9WvQmD
eoq/q6V1yuayDY5XL12DPdY2S4pp+Gsst/pJMDE3uTO9VKtvPvvllfQODoOpeLj4
CYdbdZFtLHLFuPSfXvyP6YpZ9n/HYmvU+mf0kdJQm9hB7pfY21WFyIYq0/BmKLn8
cOFZtw/Z5qMlLNEMBUBWvjojCsRfzWR6CU4BK/TNayHLaYHWDmA1U3AG+VqhOeB+
t8M18QBQhWrCZWmHuymXmBvKoCWjEz6nCVozSfTr34k6YUK1WYaZDp7ktlqeFq3D
vs8yuPe7ZcgOmrCYSRkRNfinWMluB92jd9/mttCrbVTXtsZsDE8JL9lPSUVk+6Kj
zyIim95Y+uqoy+MNv9/JsLT/2jLaq3GM+j/eI2GxVCpgx0w4YIV8wp1dGUP1UfA8
f9JvdlLZoxdIxEm2vTcsPXnt84bOj2IuaHmluXbmU+y5DvIymuLMI6l54UFdX2vg
sLTtKNwTft0kNuG1Ya8if89JnVKep8bH6Z6sOAmTz3ifGO0+wARsQh3az2ZrtoTn
zVfrX+hWhrRRokNxpTf0mNjhz1Va7+z5gszic9QTGBVD2d1SF3e8dko2pgKoky4Q
+N7pO/CoD+oOMYcvGhRhAH2ND6W/LtytJHL9J+sG50m9WZ8g81myPJngmJipLRIN
K0w5loMQ5VGv7ARTigtRwrxxIDsmZkD5Lqf9w662Am+iMiUsoozO67IXgJJfe0hA
3K3Ya6ngfMhFlDDp9YzAR4f6DVwnB2kZnsHyyCaUTp15Vde1+RdOxhVHvrzGsP+i
aa3gtUsDmi05SPekOnZtFCfb3C9jmg7vzUHVMuPhudNq4XrU8PdydVqyhwvAp/x7
dB6SVaaohOR/rO5lOSYU4ajacrvUmI/rvFfgNfKSrhVT489k7mhoTBcdoIY4NcAu
x2aaHhzoXEzkOVmI/zBhIOQucL5Y/u0lf1EIEcePceG7XyVvB5XKYVbtOW5XGDU/
YTUWI7dWeRxqU0EM5BEh2C9V7nfcRODYZj+iRcHwlVQ4+MD+Yw0PYdhpdC7Jw6wr
pXiw74VjXuxhIeyOCyUAp7DcYmDmvyZA9VenWgvTz5kORJdBACvr1cKBaDHg7bQW
CCdthmHNOBq8YorgASrWIX3CKWV4os9w7hCwC7XI5c6yWlML/adXui+HDb29dDZi
X5JlQav9fVDktD+7k+rUdwIxNNl5j5xXXI0aQy16hWzgBYVi2/EHWdI/lgyNg/ie
43o8e+eLQHg84KiJ20nyeBUGyd73kbvU47gY1wcuCKtHmmaRZXKDQpoVHLjudE29
Xaw1qnIhZRpQLF9ZLX82ehQ5rj5Q6c4PJQGlNEQzWp5h6VPV+IDKNd3+K3yUTKMk
YZm/vp5ENYR4yC7+VKgUh3ZFlpSt6cfr5/90X9jDh0ibbEIiUtnfXG9GUXYMLAjT
gFTcJYq4LSFdH5ZdTf354XCA1gsPx/JGdFg8IMhAsQa/Rs5rDNNQH21krAwgU2hN
FSf0YGEoKYzlHjzBjHNDGffux7rrNYhrryONxlB8UHisPscxprG7GFRIZ43s23aU
nOfh+dGH5U+2f4YHOlXtERYwoTzQtivonROeSGwR8zV+q0y4mCkJqJnWv9kPpIdG
WlNnQeNUVKiEkDR0dEBK0AQE3BwvcuuXU5N72S+vtKpuWqklmqPbGHABmJ2y6gBC
z5BVFEBrrTRVWQ+oqauYc8JuEbFInxA0pjnW8bSzGxz6tMb8hfbBaGxSdVr8AQ/O
xMtNpO9mkYmgN1hM/+NbL+oQ13MBo9DMzyAboGLT+OYOJ7aIqumIAwPSgIGUOjVI
jcHqa3MFZBUgFiDKcV+93FuMMyJjeqx1NrA39hA50i75IUxb5tkPLwDDfiBjGJau
I2uJd9MF9FfHAp6m1GHHHK6VI0hh/5fqj13l7LOc+rpHfl8ZynulCW8TqH0SBgN7
oy/ZOgpHoPEI8GfTA4T+FgMc3VaUjJ1GXaksyps+e9NF03Jl//0Ge/aSnkXiarsv
K8yrIoBfBzNgKmFLeROPyBgZo1oqRPWOGrlCUUFU8p4XQRMO7pt+3N64Nn70o1AY
q6yT5jTOt12N1oh7ZFBNU1TWDU/RjbKx+2RSWvV9F432kDE8Z4WwKOPnvhHwuc5M
/41VZ9B+z7WNbMd5Bh07qpFcL/Vv8r6fP1EHrf4AvHS1MLmTtxGTP1NGN0uW4Ng5
hVuWhUijK84QfRBa+Bu9Q0xwIcZOYkGS02RwGiGQWb+YG+6ohxlbyxztsvLNCuid
3+YHjt/twD1dS0mm96m9s2T9KHx2ILadD7yLvtdmOIN13ckiC8Mx4vI+xWGAdivv
eTCh3pnhh5Lf4A8lRdNjq6prVICTORxFLxDCtrNEEFhu16rHt7sLndURunKxDsfI
gl2SdB2WACi5xXeEao8i3WSLtJKW9uleD6sNIP04dBTSZsZ3DBndmn/18fm35R8r
ev4h6v717HimwluzlMkA0/1tAo+57RPd5D+AkGrCw5qbnH+k2RbkAz02MojUtuUG
E4y0q/TwX+vaq3gRpDY+ytiG2c+wrk1Fmt1WAQTbXsqPQX0oNFIWeVr6S62iczpw
XA/3w7QY7kanPomwuHOTAw/cTa3omMofDXGn7A+E405oZ+Bw57VY35jU9jq5Gghu
akhJ+6VBMrMPg4/g/ITiHwHE6iySNJlwzhptuoXuiP5JAlH8v1471MVveLDKjtf/
0g+KzxdGhRxXs9nF671dVjFdGxSEnsiIFaa/ZDkn3E18fZ6T66WNDHUbmCmx+JEJ
8FavIBPahze3G+oR6dFFJh8c5AED4l3ClpxB2b1cd+CEjrN8gTeaAcU06kDlm0EQ
w6oZcUBXDL9Xoe8hZN593YoU0PG8ORy2fByCwCFK5CKelQ/pN/jvur8uVw3bXQho
7yAd0M2rS3CZ2+/VCt3ubtczlB1XiRjmjnCtHuTRNmu/5rdEJuFrDaxjk0YeSbRV
Cbii/PEfw5q2cJk3g2Glv4R9PIbGA7EjqOeYoon8UW7lNNrwFxcEGDUHnauOznuh
uVocDf48JU+5T3wDtEe/a21Oyx0PN42zgjEkgrESt7ulfrXhrfm3C8Mq/kntJE4B
rGUEIAUNfzLcZ63d5s4WokoCVEf8VZW99XOHhSeVRo1uTVLJ6xuzyGaaRBT9DdA6
Q/tJGgp1e7E3anEz07Er3E9mdyc7sfPZ4V/TSCQurSNqPo0GBkIa8jTOdX6+k+0v
lU3BQbdt8fKUgWztLOuvXAfZfivmIyybg9Fw5kObw1alYh6HgpynbRXZyLsYlcHD
kdAJG9L9IAS3K8e9c85KsavZvsqNXOalk9keevgjEmi8WUFlRuL1yFmKBITXSPsO
CZ6pBc5hf9gRNSmjCNhQ4JBsl2iTTyldQy/e7/8D8bnAty6QBusmd3MWcoIkj8C7
jXDiW+3trOM6cKKPf7DmDq21eO4raDbUJFkyEzVtUc3JiFBoeWlB94CizpkFtiix
IRC4O4N92rISPMDG6ID9/TJYGmzC9hkn2j9HLSBq2x4Vyg2gT4wm3U+Vd7two19E
clUjG7wdiSMOW2x8VzWBHoIMug+lHOujuavUrH8lquqsmfIQAqkMbsGnmX5HuOsK
ouXymlwQxQU0uLmWlQNsdtr1ATNKasu6bHAZIA1LSwHxDptdOjP5kc5HmSsDKRJV
FrwIKdlM1063MJyyN3GcYmNJncdRgIevQdB89wP8QXw9ihREtxVREnRCyKES2pNV
gvE3w8v4bMaz/GuANGPBF3fc4XbUQgBNMZ8A3j0ySXIYwCRZluetQ4GV9qtuWRDH
3gE3b/JmSH/kKtUwPOIWGiWxs8oF6Gcw3PqrdPEgnlDnTvlJYoej7bNJ4P730gRy
NGoCH10pLPB4/lHwYwQTgpkO1a+f6PRmsOVXz6ccE5q/WPESIAp+wK6AzCDyXSEE
FW4jwjVkKgjbyCCAru8YCt4om0GDSFkSgaXYqkZmAJMGPmSbEvjeJQYG9hh07eQ2
dSDOEAXuP0vhRC/QjD3n1hfsZFns5GcdYLjP0CXJxQUrUSaG0Q61GIVxvSjN4aKt
QQA89t6Qe6oOv7u6umiPZDi5DpVRGx3GhmUGDrox1fepRq1X7s6ltCP2hbuZfM1Y
fu/zL1JfFsauoZpUeAVa+bhJ20H9VtSc6Uk3GbizzwFay2VX9mYxcyD0TUkGZ+Oi
A+KG1SRtUVC8VJWbxqNyKJEmz7fRnZiaemRIDeRanjDxa/E8+A5pxlF5SWR38wWp
tKFCFAOSAnFajR2s9x9JYIY0Yl+1rZXjASm8hvfVEHWN+H+bSN6pgJGF5FRleOKE
rAmzIPrHjdLVajvsGZJEXDeasQPv6Q3IyEB2Le7HmOjWp9IM4W9djAmEkbhACpMr
vXyXTKOxFa7/h3Si2gTbyZQoCqv40sGed6s0jYLCOWPpGXiKhYJHL1WP0dJkbncI
5YbdT5lJUOmKukookV2Rv31Z8Kfx4j8WPh7WWuB2diPscgHa2DFj4AJpuS1v1VYY
ZLeNI1X2ZktC2bCnXEwPu4v9JozcD+HwHWfOgsd2SUSO+vAXmY+HgH+Qh5MfqcN7
t5ihuxmi0VZegMiCgDWgIt05dCskhT41K/0z/0UicClNGp+ghDXY6o8bXhe+Dvwg
GJ9tzCQM/2wSD9u4UoinCS/oCcKTjVCptcroPVzwLGcBHjDcyRTf9n82pKm0mKTg
fUI98XjLlyxYgIfVKAC45B7GdQfUKcJ7i+nXqZMWWd6qjzL4k/ATgyOPTdiqBth8
AYhgxbf0b7QbbTkBbkVkqgtuxJ8eUHHcb5AevSeWzCJdhy7zFJk55QXP/1OrtgNh
dAIa2b3vfTuAcJVFFJk9OuPhITyHMSPoV19uUNyIsiOHiO4R73eYYKkKxkGVD4rk
/2GV3DXZFjCN8gF2+Hqi6VOOVuOS2LDwK3lhCdQxzizesE4/DVhegG9ddHudhZaw
1Ecm6inA0XnIFJFVMIJ9UF1qN36H9+5PEp2Ep9OEpqInOjP405jBIc79B9oXnz89
Mi5tjNOUdyUMigtK1qWZSQ9dPY9LGN5oUpXrS9pjqTrlD2krc9JMwQyUn4TqmRgs
OjNT8OcvTYHH+Li1gm+kKwQpt7P4oPQMY7mSJPPOnR+zZK2JE916gB0akEjZ+XcJ
4uakTlp5FFHJor23ryj8f9rg15ezj4uGaYUyMHbQr7Je2j5u4vnFiywmQYnSQ3WY
kchSAfcyEegOntrvBAWu+8vIxQzd/uJZxumIwfolSwEvHxPKGdLws53oK1FvMEGq
9NAz37zzhJkS5mz20JNCuW3sUOWxY/wG5zwATYiSsMi2fsV5p57qEO+2HFVgGv/8
IFyYY6oT5gC2MaT5hHt3dM/4COO01AwWOP1oOJRIu3usicOghG6BmieWHbXp8J7Y
QajYR6ct6hT2uSSaEB+W7vKFbhAUN51tkT8Obtwso9Wxw2XfLI+ur/8TnvimDyN3
yDTBZOFalzkFP6BeNRdhjoI/GXgWrMjTzzoc1om4SKxn0Do4/v3/PnnWxc7sfR2w
VqqLUcM2U3j/1CKekiMTmcBAsb1KrYDJBGF3dcV3VUGUb6XL9zCkvW3BzlOXH/vz
k73NjYlEeOjMoKz8zvoeyo1m2qhp6bKXAYuO/Tu3bxNXIZgILL12XCXazyIRTSjE
qSQtBzyCN5z3kIRZdqyHDtNgfI88tETWZs/rHF87bX9bT3to5Q8PVusg73GGgwxG
a4g67CSkG1tH1jmp+jhLcO1coIKoEjptqEXvwhte9h/eDGfL/ebySbynfLYxq57+
eLz4KWVVNAe0roL0y+l7NPjmI+pDacJlog+csVzYR4SeRr9LtHPAT6rWSd5WIZ+O
zdFg0MYIRWnko8SXaRRioEVZq7w4GqfKreo55cRjvDlzh6mdPOKmpKNzTzOvMGt+
yM5J6WCoN2rglvdnP+x+aqVmP3u0aIu2m5Yswfltj9S+Kkz5i3a9/3PjAd/Cm2yx
2q4f8LO6mN4sRwvfI3ghjYYElnloocFuvfDqmsaOn6W67PbZ9NViPYadgvgUwvsB
EDX7bDPKNQfY/RL34OwPZ320q/p+Ui7ZyOCdknCE6odMr/BT13Nq3NrFSyDlOlc6
eCzyIIjalg2zrJtgRLr5pVRLc1qpgZcHbF9WcP/kxqT0htXfyOzQ0NeAcwInb2Jn
kZcsr7j8+gKdSDa1dqKQxjwQVIXD1tNiL72X0SUf2TnrjldpoNlYCrZoFVvA1psO
sQWoMYItnDKsttUwZJPYpHQYHeMwDwtXzeSDGTL7wTmgxRD0va6213+C87Z232WV
fGH4mlFIw9OasTRD+45kQGYgQa2ZfCg2/3HgFV+7s0cqgMcdFRoc4Udp+Er7odee
XLiursUxEhQpeG7vj9ib8mWtqi7U2Ho9fhFmQHajb7TdMpb+jokCybNBzFS8Jqq6
90lgeXqOhvkvBX8HvdUxmuKdcAESHmECXkzJ3KC9/nz20vPOkrTjP/gT+3MaX8kH
lH9FqFkc05OPt4j7a/78TfU71PrWCCnxmtLUyzg16qKtGFqx6spm+dqsSl029o/z
0vvsAiuIP1BozLmcsNUx10lKQibNLVSYMEq6s67yCxKF1pcZygzKqBSi6xcJDVFv
/lQzxQ+nhvEAw91v4iUZV2TqkjtMP0VSoQf/Gg5iX/AVSvruwqf9bqdnjk7b28hg
z4bn8MBi0MKta7AqNS56mfhHEYVF61rp3SU2hfbF8hz+92TndBUtyQkbQ7o/jgpy
ZHmSNyBkDv3rkNoBWY4fmkpZEmg2Y24WJXezvn8lq8sd08kJRthcyaAZXxu4+Mb3
M2jGQoNkBkjSfGcXAFj2JNu2renj47csGu6gcBOI9a8AU9z3PD5pqdmrYcOstCMM
nufHR/tM++oPzu2eSL1bD8gkkUjfX7+CKsr0AieuAWMYBDGxPqIOluDF/lR8cG/e
zP1BDSkPRWOs7Ey+LRJ7INh/d27nAiW1OvRSxiLBuM4m3xilRO7m7p242N1Ww1fC
ZIpAGq7tjNcRgPu/gCMHLRwJZuKDYKJQEWrb7CXBDvPCQfwZdZ1xmkQAoitRR02h
snzbsM9oVFBTGEvxEu6RZij50gGpM5DP+w7qtFiTu2eui5a7D9mKMDNBkzKFit0r
XB5jrO2Xmy1fsY3QvBmgApJPpPuMGczHWYKR6YbKpQw3lRGBygk8CpIA7ssWy0h/
BFpnj+wdQ8OHj4ky2SIFB7XTD6vDu49oyOdiq1ZGeusjG8QgFiSEU9tn0waiCe8B
WoNDytMb3kMStoVkBkjUKm5Jj+5TPzQfK0cNzf6I5x1KRNySSl+qFR3vz+h1oJha
9468YnJ7VnoIN8DuJNk7fLBRaNUPQf9U3b8BVLE3k1NyFhRSOCCzY2fnbZFotsOM
DtARjDfKQdKKP6nU6lUg36kzlFhVS2GUoypYWMa6g4XcgKV9lQOK9ndMKRI9Dw4Z
o6UAx19RRhZPhbGfWjqyroO8l8q+ocrORgw6d0ANJOfAYbxdKI8haajV5k8dQlIW
cZm3jTRongNFgAqf0hqNppdPHojUfIwFtRAH5xB+9vT3wp+AlGoO3OscKr1A0TCS
mD8qkg0v6SBexlDelQG+TktRqUB1zbxrdGpOG1pL6Y1Jc8e9zSjoVORrHXiIv4NO
Srmt9MYIwRSkivEg6fhxqIThdE7ms49K+wJw1tWtXQKVvm7OdgIvFs9DlHsqyfQz
cTC4XPdtJymscJixb6Qu/SO8+2q1p3XmntNQpDPx8Uux7pyMFnBLsLReM3C/EfTz
B2UMA4m6EMqog5q19RRvFGD5pVKOULHaxH8HjbfOWGTtGxfh9QuHwqhYuEQrWpkC
dk/lWMgkWa3FQQkVtq/pxnja//xtrj+vBgRyfjgduO72YE4McPhLDyF2O6DCszxm
ReHcfHnjDb8tLGWh8Gko0thwonPK1mKJ2mwnmCpjQ1buaJL5hEFoc+vNEvpbUdzg
NqG0GOYXHwEqjRKDkTaTj5Uwk8QE92mngkAbRcHWzjAZqtbry1HeY9nhPigHuPbu
zRFNG+ryoct3Zhi8mWn9G4RLolB6j/d0PBcm8ZqS6myC9zsJd8mb7nXkoY+mxeG6
ID3oVypF20mLEInpPv62XSzcRB0f2dfO7QQ8frqZyXn7qurET1LGtOsGZ7cUVpcS
euLGU5wznN51KVhfc6FmZoucCOLlvmAi7v8z3IlloapAUk/PKxlOCMC2WnXVkXBk
VVdtkyZ0fU6hQpWV6zrHCyX6sSUQ0HPJgi105RK80/retoq71+9DLb/4i8TSQnYT
8Dd3AUpqeBtWF/d2qYXWi9xJVOD0iVKOB0Cy++ORLP6RoJ29oejxa7Vp2WWG0aOF
eeR2eyE8mQ+T/hup1RKZqQOuXQYwGV0IjebT/ba/6A6r8VHwhvlhZWkmOyldP0hF
Re7l7S61/DyTM9p4/6GDGhiGYz+Hu36MJeO/FDIan1w7rMCpEASmcN6HMY08+Flm
FqiSTa2NWnGoDP53M+LU502u3/GJs6b2A8WBPGqC/3PKXEehbv1C21ILrvNUTHPc
YpVVIkr193Zrjdg38SFEJqKlHKKzFdfGU1k9qKljWQC81gjjtleAtZ6Z5T3V8PJQ
N7i2p1OnspUZ8b9jCX/kuCiOjVzjtyDwC/xfwV8xKrUab7mkxfQN/POeNtAXJwLc
fdHgaAS8umZejOLn6xEkbrqCHHrBVY9B5WKKRGHbR+Olx+3g0Ubi8C4zIDMj2kFn
Sj+wLqR9uBD7L4DZrL7i0hu6B7tIHuTOWrMNZvdu8L5RsWTPnjD7K5IkLsclsHwm
LVr6JO0sUZk72A3pZwQb8thPK2kUYVxpW9R60pPrN5dD2lfIpCDH2dCFhnbbm/4X
aqAGG79Z8eztuVEme0Is4sRg3eeFxKCV7BclFnvabsQ627xQjOwzDGZH3Nkgeigq
83b9/ixqVaCeoF5zBRtntBVgAbT10J70xoCeD18ar5vWwIled9D+KcjYRanw9VOm
z58zJOCPLlcIeK05foTAldXeOeR38OawgUfdZ+OWSkJJ4V8QqqM7gsaf8KnuIFfW
iB6v858o2My9LmR8Q/8f/X+dWRwCvf87LcOod5MXVZpKCecZDZSnSO+85sOPM4iO
729O5MsudNjmVlxrAig6nVgu++klxKtfLNTXQR4paS4m2G3IgIAdLeBKNS7gGylX
YaTHmszFC6mgSaHGeSquzU3pu9YilNID6EMJEP0cOt+HujsS7qs2mu3jFxHvQHaJ
zywa8vEPxIGCZ6wQUsqY7z1uMZOtr4HkG9fV8kuPm3EYRL3++Qz0/Ndo8/gUeEis
Kwy1ro/WalsU1Ul19CU54MIOppwQifvXCxmNEZlIbj13N7IJrTIXcLS4EMHTgzzE
BLfs84OlRTNbQiTSZS1KatRPPC+lsZtSqkbEhNncQPYnmLHgHsb81Ylkpy3ysdX3
8y6QeP6tn3NXTlZ8WCkwq134hB+03lLnwJ7FNLoxpIJvMaJpDE3vmlHgggIkaqpr
TV8Y1Mt/TXpF2APB6qC5J4EdDcDCyQkVyYu2EREu4NqwL/PzoyZJIfXcfg58TLTo
tcP9K5HACyRY4s1Vefm9WCwDKV7mjivQwOpRtrR6C4Ouu7GXziCyVrx7QlgkWLMu
L7eFhBP7oVWwhme8v0+QDvY38lw0h7UrtkSqQn0+1d5H+tKp9zutcMNIIapy/nVe
G3heV7ki9dpSeu6ACRKsoVtgwTuyhXM3BV2/iqiyxac+1KJ0Qs7ZTeLsxoi5Ox2c
wJRUHTIdsGSZwLxxb+IpB8J0qs8A+DvizTyUIVcYiv9QlfwlonAWSx8JDlgt9vqP
ljdqCCO1a1mRkj16kWaCtNjjDiKCriNMUkZgWw8iPPj0QDhr66M/fNAMiEYpQYN/
PEl8MuW7p4JSn6vJLcyBJhSfaTUpC4ubprZp/qvzz0FS7t0Yt8C36Li6lmI6Lvxr
6gaIhWrkrqlnPU/n94m2gnIy+zjxT1vohvP9kXHW1td0ihLUVyeHygUB4MWPRMsS
yKf2OkyAjRwcdoJzT5rCIYGqB+a60vYMpmJWrufVpclbd/F0bd0y2mmASbVQZd+Q
MEFleyzjvM4y4RA/+jVl5JZ9qC31SF2Pfqnt43rGLQVIGnvTglrByzQmq2qTS8Ev
AEv3TKTTSnvnc97QYiOFeRuesRnese0GG+q4TSiUtbZo3KZn2/A5vaxusX2BZ2Ng
+nazl23Ffkf9QOhrycHJ0gM2PbAdMRu+IlzCetrEBQOywLjl9Pr7MJjx515QjjGT
i6k5/ACTRgXyBZS7KGS9+9N/2bePYZOlFbMWWEmeRXblPQYEzCuUgWxXzv1YZwK7
NY5dL2caJFhBSCDlEEbrqHprovJw581wkNH6wu/26ceARshLf/dG9b0euySQAd7Q
6P67uPCdbOXo8JUHminvWSIFBWRp3UQA/w68tvL74JNl37rbCUFescRg8v78pHki
RdVf0sfF0yuvcRvL+wkY3qzhzrxLzFHSFy1Kc3w91bnuogz885dNjaNu41FmbPpl
ELhQtt+sQJVF7b9HNiDTYZWVO+Z5CGwErXVnNQ1qSul/sWpymA+sJnxC0y5Q32b/
AT/Ad5raN+Rb9NtKL5Gz7veXsu3tHa12Xgo+nDz2dXUrv+iu14NHzJHeWJ8pe4p6
X3JKzNBruLqW+9B8ITTzPRmjZRes1BZZUvS8Hy4B6OvC7cSkB5uzB72iP8zQibtT
jdn1Z7QXxgS5Y4DgoqZo766Zn8C3n6qHea+ImF0QnzVWgDVOywVWa+wG91+1yzWC
HnEkEqzrggDD7ueOpJlwmcuAOyshjRtWqMIXOuanmUAAH82xxD6rRJNwqCb5Cl8D
i9JRQnWS7pO8Hkp4lLm1J+74ag9KR70HxPPlSNP5fErUAGHaTsmnpuAH5J/nDStK
bx0ynoWZcPf+ubizm/7s+Nm//JyFKNzL0UIuLEhTU2RlDREunZ+3xob3Rd4IbpUN
fI0WK7W6ReVroKUcZjEMr/yvV/gLX1vN4NW25y0QjSN97OaUIzE8zU6wRR2dESEG
nQjdVcOKIm6NxpwkEQBY6xmaCglX4KHjUnpQ9LdleAaQWuHVUM/z/4+Qfv8l/2xd
ldxpmpOsKkneJmENc6X1zuNZKYk97VlfcayPn+v636v66rEzgq9fQGv34ZOohkTk
7cNV73uzAOGgniJF551d/2Nb2dcJE9/d/WpROYnqPO86o+QC4o6AhiO0UGNl9/Xa
Z4WIi1j6owj/ohEYVDdOOE+5Z7zYOXo4IrJ/SUKbJ0n/rRVlxXKYMJwdo8cwyhzK
5EdbRDx39ECwD0G6UW4KC6xJo4L+yABTBCvM448BD5uUiuQeolOB3uPHr8lDnk5s
BDieHVlgx50VQ7EYZMV7etzSJ+1bLVTiNdVLPHkgZAV6muYokQldBJ1aZvDdpYrb
bwhPGUr7UxMwjjnUEoH8iaZqb3NxN/ERuDYrrSgP6qv8U+rpFCWAodSmdWFwrzAa
utpDKMZKxjwzJDc9TH6AOLpKxD2l6iYBXcevkxe5sJZrRR4mzrsuf7MUCRA9mcrQ
kbFLtZurWe7Nt9LVk+pBjm4Gi4XM+ri4jhGSt05grOtFWnQkZ6EpoV2UCMn3UVWk
hFkBzE9PRCfEwv3xFEodK+ZpWe/bTzUDJu8iquh6UbFUfB9aL9LboI3u+dQiVQs4
awKSlu1zHKyl2IYhEFQ/ipq3x8XvPRvvkTdaAYGD8Ng/qk4jdFpc893/7u2kSbj/
QCQzge9I4E9KdojduFexwfA4abgdMx94rns+U31SW9FLsqzvEPktFN8Pg3p0wSdK
6IrRzAj6hzIUl5G0IWZ2q6o8Ecl6u/7KBkfzyWuPjftLpekGLAAqlfSDx+OV+UEJ
Umg4CTdbbMVBz8dFylIIgvbyCj3+5Guxy8c8XhPMFJs19JaVuKqd4h6eaZ4sB190
aFT03ZkxK78YKuJpvWk1VkUpoSZvFFUkuzvpC3Fc8vHmQtR9Rvr6gQvFJCdBAtFg
/YHORLN3Nc9wbQ3asudAac/ymn/7D+vwB9pN7P9jCTAw9Tr/Q759DBjRkbe4JZEZ
HoqMCVU0PXU3TEm+aws4BINWfY4rq3ITXEHdNXf/FbTAhZCN/nj2wUogVt1Uj1mV
vh/KvKyymDeyQdWgGIO2033OaCZ2AeMQ8zCrysGiSf7Z5GpQNa6sLOS3oB/+MpQX
pk7OkeemuRHxL57sRk1ZVoscd/9XTrpKgHp7Jp0KxrAzow2ud0EV2s7yjCMnygP0
W61NyAlghjXbb713Wn/L5SGD3JpUHlQx3PGyv90aKVir+1lYxI0bd+Ha9vNPjTly
f/RTokVv2oZ2YNLNYZ9SXBrLdQuOx+NQ23po4JFK+rXMIOXStFtxcr9RnfqJGDXc
4f1Cq4k2ibRPj30LG6dsqe44sZ+so/X9igzOGkf/U2pj9gpjb48UC6de66erQfEl
t5FKgxFeHpwZqGzYQkcAPCLakXJm+SW1xT7yg10cNE0vMPaKdvP5TrcoVYKZaZJZ
iPI+kEcbjWY7Gt+77Oqsm/MS6oF7jjbeoVJ2gjrohpbnlSuir6EXeRLRK1+YII8Q
y7foQQD9c2cS+CHCpLRQHalabmvcK8SlDDMgkqDuePiwQXVbZlFMS2fwwMrbdmyE
0OG4K1S70Y94UeTRLUk3YX8JTDsdw1Tx67YBlUEqT6zbSuaF6CSeeGXIrBMsH/Ji
ReFo+wTl9Lqo6Z4oijgPOxOHWVzbuActRLtTJ4d8sSwBfJHbhpjYMGY9CcG3NtDd
HZjtj5TNYpR7Q0kIwYlmfQzPBrmqF5dgWbJgHpCmIgHZ7TC9zfdHUyP1O1qVKTom
/fNfFaALzkh0/r0fJpwK8Dt3193Ed5D8a5G9UuvPiwUZmzoVuigI/B43bs+qosqX
Zgk5YEC/8k/r2xwO/+e/sQyKZgnMyBksR3qv0EOXgjq0C2prXiJh2tmVJPMynpit
6nKQ16jKdmRQJHqpqLJ7rFwdOZdEM/YguQ367maSqJOKxCR7hnw7h4vy2TjW2srQ
oCuqvRNazIfdq/HKQ7aYPKtM+mIiV4/Zt3rbD5g8KBAU+E0JJdY87K0ikHZGlg+N
Jldn8ctkeDtiTCkdc3LbshJIi1+0r9SGHeV6168yb52y8MHMeOpRH76PEga61Ijt
40nRrAkvdOZeEAKqOVnfz+YYKPyY+6Du50n5fO/5M5bMZIwRZq8TRBiK6IE+Da7Q
v18EUosaz5jY+LHBy6Pws2storv1n9gwyUkrmi7fVYJ1VxYhjfG78pGzF2f03mJ1
3ZlcLo35zjlHOcCcn2/hKEIgyVzxennDJx+rlZtK7M4lzxsbbCaznLde59iZNSom
/m3OylXrz3VGG5YMEItywGtmb8ItPptUP917UiyVaUb101Vc6uvQ15RhHr9C3z/p
mM0WYJfAOQMFL5XJ2Eld+Gg7z7wVZjLKwEL4SRAEA/BO5AQrLuEflX0c238Rgscu
qf5tMn/AUItKl9MziEc3bHS+drivgaD06QdRFqKJo9EGZhw+8iFz9/Dt3JKYl8FB
4A3cDQnM8cq5x/pBgjgXbvA07Xvk4qSHM1mNO17v85DZ34pS+rYromEmRwqhev1k
ncA335xgIFibNTmzC+1bNOFV9brjp7gj0nySIgzPgA+F3MmrclU8U0TIz9dROS/B
i79dY0RoekOf1x6QMmA7huwdZgy+pIbixvFaJMnQfoGPIOgSpwns1Ja/oJAR+DRX
haG+X6Gh35f1EZIFnlyl+h285+Fz9ivvZ+3opEsZ8SgvXSGf6Qzzu7pFIntPNgM6
yBPCHJuVplqqACOSeGYuOAnHmYaFh71RFe+ybvSXma33B0vDXGX9Jdx0EQlznH//
ynNBZBH12fF6iDmH95RBZiAEZcJh2uR8IOClVI1oTtaBeKGtOxtPOFEYvn8iKd1h
v8YWZzTSFS5ux+5r/o4GBtCIETRWaSf+KVSKL3T0zbLLkA+0CULRgvbMCn5uUY9Z
NJg9VcUYLS3xhx55K+seisrJ0gAAy01d6IkM+rO5ZBXmypF6jnKuDBya5uy5xBLY
cFyMSXs3+iFBoCoXtgfX9LHdAXEuQ3REoHX1ezKiLZXES/Jr6SUlGbQi3yR5hJGW
bGOKVFlmPhcL/Pg5XSzrir2ddvgLM1tmRhA+thbxvlzdU870FviXs9kTIs2v284q
GHc0DkaV3bRaphWMPf6qk2oq6TN224xrZd85Hq91wFjrMyXCm8Z1pHqmdW5oeZK2
aVFNWT58vQjSLTGdeyOeALSnKKOBZxl4Vlhg7at4CmXboON7w/0xcCeWjZFTkmg0
WL2WlfbcjbQLZV6OxfX+x5Dj6sQNgqc4Q2ygNlsYxeAZIfT9Zqk2Rfm/Alf2zpfS
rjy74JsxFkhoK4LF5Z/gHZAe9gxGM7fBJBfdbKlHzbEhG4ViCqHu8/BvmEbgIrc5
DL9XwiXE4AAbLKG66SHGY5iINGW/1lfbZchiD0oYRwH2K9GoMlLWUmUoiVvi47QX
3wLsXRWPH19s51Tll2ytJL2EWrpXe0riqPrfFHinVac532VOZ08fjoAxJf/tGVqT
frHWjqhN9jda4/rL/D9Hg5OCvpu3QrHLeVu25J+P8jzpeBfCNi5TYuF6639z3SFn
O7OUPOP+SMrx3HEEAttj+Xg7RlUr/Bm9aOtRQgJ7uNNOIcyozbZv8tdZlXdHqExY
kFxYPSl2Ab/AKVA62ArUzcbWxrN/fdbhvpn5ZIJ4EZiPmwCdQ5lA6IS57gjn8mv7
0sWEq7XMeSABiDDTSxSeXQk6R7qAxctAQmCNEx1LL+c1n6IDnXQpaSjThAiOxmvh
4t2QdT8QvW4PhjmvztAnc5s30lK/sQuJ6rFDjlPKTbFHVbXRCAlCEccya2m9JF9I
mSstNSE1igH/Ttfp1T/NLYiyckzUgXYNPNaxQOJnMz/OUDt58Uux3r3lWCgLMyZZ
Y/vYtwv4rH8K3VobHLOsrWtAf2Ldy/uS6VK98EBahyzcLvvuQKjqxmusnasEE41R
QKiWbEuwsU3GdjwOKeDkBRx7++RHmfMUGE1wH+1aS4bgS3kN0nqRyEbmcDc5B7ET
lc40g1rvyhzV/lsexmvbTlI1R0u00c3AHr6uxtnKyOx/h4/wlveLnrVF8ekocyiU
k+zaPjE64w4OypKoGhFbPRQiNZ3yObGbmI2a6nkct9aKoqzVa2NTlFMD0bdjoa77
e8xxNKAo0afS1xaZl71HkFn9/Z0NkZxKLaeMlBsLH2FT89dfA0FbRH5ZDxW32dWo
NAh66WN2BGbpv51gbTdgyitdYKqVBdxReZ3KIuPdESfbBD9RLcdk+9VPAiPT4Qyz
LsUs/PJsN157gvJtnY1HchjuwvKGAgEeLsrXToxZKQ0vVgIEhMDOuStfcVN/U9DO
kEln4WlMj4NJoz6x6pgeetFa7ziv7KQHc+N1yjnoJKTHap9eI/0yN1nkUsTHO1Pc
LwzeTDUVFcJEkr0KQ2YoBArPUF9T/7B4HluxDJw/PJsxClBqye1FQOVG+5hpUju2
Cn1JBKcCJx+zcrITHhXHxH02pfrWb1y0esVCw5ycfCHbJAqwr6kuFJ4DTsICJ7Bz
tQVGcjsK5JGoIdqPS7gRWjB2oQnX3tBofa7BkWUasDKCdFw+8QOkNT8cHwsw4y87
DRPkjZAyEyCnlsNQ2mi+E3FYnB7uylrt+nkfJALdheUr+CHX0gtW3oSo/bGWg6te
uSZcIBbabc8O6VESSwzZon3kYOKabZkkIHYXFxVyd8TBsGV+J+qo933QWrD7Kfk4
SkqG7wIOrUcZ86gXrABp0dkrGirjZYVHRXHDjewT5bsP1cFHyA2jL8LK6ea3sIDg
lOSwHbcJikOZjaz+r4dr0iexKpjGGX5G73Eoo9h9hDlEiyXWK/NoK4wMTWeGA5a2
GWCwK/o25sJBkClkvkxwRsZ3PPV9zA5UreIXznM6M4VKcRv9aOkP/XDRo828a5ra
PWLWEcrAAOUl2KhWlnkIoZKv0UfyRPAGDhG6CNVVp6YBunwSFXBJ4LkBmox5gqUh
vzo10+ve0a9mrkEQ63/eI3KO/dl16BEoiXSJ0rHNYbrELOZ80RxBkvbRSGD/wzJ9
NwwoFi55LtDN0eu6qiaIVARfrbc5ZK031oo75tkTTePlMw43Gm3VKcQFlXTf1u/D
8nnyOEIwAnwRJCujih7YVmZGAdlsX4oI7PFfWvGvUTv7bZnlE69yK0XWHffXRbCN
MzPWjer0+HP1LF5KB0p7ti81JCqCyCnGTsdQYdY8jBRNs2bxdvxkX42yMonVtq5Q
QhFo01+gYeU8jZ4CBftQ1/wd0GO5nALgiU5PAKzbSme8Z8vG0C6qVodCAIw2CFTp
8NDS0BKKLptJ+59DJRDfZ4oHgU622wIsezJT2oqPAX4ZdCq9iu0gsjAsoVqmJaS9
+hVxVW1itvRbj7i9eAOSLZvNpjrl1hN+etedYh+eryX8FFS21/z/dgrBXgopJUOB
RR7HDYS6nUwsbIOLQFoJH+S88m3iGfC4TBtnL6SN1Y4BFi7/SfLzsxcLG8jqpPFM
bj0GTLyJrqxxch18vtYwp6bsm+cyMX9ia0qmm7GPngyRTVcDl3pMGgD26E5VFxXL
Q8SQP5NTEPOiXzSqx+OQXFnVZJA4HBA0qMmBP/Km598VorlrWubRyWHs61xqS5jX
4HVvr12yrfhW4H64nRKKEUDLbvfWg/pMS9uAE87L4745m3ICm86Xwzn9dQxLTYMd
ZX41yGipKGKfmWxtN8KpIxxCed6XEIohTHwVY1Vf+pMGj98xxfQ38CsfOkVjzfM3
A3J2zzUwM1sWNMzBVRxofB97SehqvxA17Wiqrl7Ifb08NW9cqVKgltu9HTa92ipX
yw17JETuEkbdayWJ88hZkt9qex5qg81oBzA0lFbZ6Q6UO6tLrOyhvFDufoyflsoQ
QSJNQ/QiDeJV689r8l6UyhmKPjAlkh9THn+oHRtOHrEmFBg4h6FTYbTp4qzzTqJH
kL7iwf5zqSEmgUTg0wLVPvG1Pi5GJPt0TQ0FQlE0/8nUbkX0hTcQnmsQmaEDqwTH
HOwToxiWB612b3EYcU4Tb2TKU6XTiNyALZ41ry3VtQfuewr10S2GWZYKZXQU3RWT
ZxD4//l4mrH7G5kA+Cev7g7aJ8k5mNZ8PGIwrmN/SJO2jhqcyGiwpF1TtBcIp1yX
kowE6y6JsJpuQ3ZECZF3hLYYgYc3l0GHIXqHmx4zuBs59PB1oRThWCDY40UVFRgw
1mGp9ee1kkgR2Joj/Oel2wCT5ChZuKpGPk1H11q+w7OIbNOY5/YVoF5l6B5MjGAM
UIKDW5wLXH+r9ql4kbL1ceznFup0z3l+ANQpyhIPaaZkPKvKn3g8zDHaEtPBQn1S
zAs4ruCbu/vcBjYyiHa8mPNuBdRGnc9sdl0t/rClGVoO8uUKcCUqZf8qz11Xdp/p
e5+fYgYHpOvPkSrCET739hX64qWREpyEapYBK6xFtSqKCu5orPWkcG+gnIQYGeuP
3iizwg59c1CdjcRBAMmifs+vP7F5FZwojMpBCNtktpi3KnT4bUEJ7ap53YBHjWAk
1sDbpW33uqyvR/RxFrmpUM5mpnudbF/MZynG1goU/b/zlAMM7FGKPwTGr5/HxLAW
lswsfWSWu6jc/2zhwoehL7hhtf8jp0S6XAjoundF2YHlMrsj2q9rtcKsclr9HZwU
ix4PA93Bot/sAhjAgnCSVtlyqt35Fo1Zda3k41lRhNlaYIpi+OQsRZK3fnQve5EI
3AkzXW8iE8pqQTK6y/jCKvidLST2yaZqrFIjxeMmM30wOGt+eeePW3dDEszx3JT3
J4y9H3icwu+2Fvg2XqEhf44Gagrr1ZRfnB1GkyvDQnPpTnOseipE80LYlzV3NaXr
BGxOlxRHBJSjWGZVcPAcdJzKEkEhMVWhi/fq01dlsTR40+9Lm5qwvIgGu5cHEax+
TZys+81+IXnhqDOZfV7xE6ncvy4CRi2IYozlWqZicNxVOOcrWqjhvkatPPUY/WJ4
g5Rtl2VZaB4AqSBzSEFyKQwy1qdJOAhWfCNyhjy+cp9d3myVp3PB+AFNeO55u7mo
1U8Kl5k4EMQdhkoQI2Fg1C3dYtYDgLPK6QSJwe9obFRatnjJDT221z0oC485qmop
Iov+UE+W94tCJodqazRdPZDHyTzRV0NgsU+gU86osXxGBLlrSRSpamzijLoHSDWq
qgRc4gy5sG3lC9OZTgF7hJlEjWxdUAsWndb/VVbLykQEx+m6tosxye7dH0qS8o6q
z8vztBAThdkbWDbNed53mDNCze8XphK5Zi397Qo7lUmY5VsXP0aD6gsIASpH39NQ
+llw+6yZuVPY+kh8wSgVrQdiQupMsZuFUP3M2QrrI5LDZTjSR8V/wZtIvNnWdUiQ
yp5sMH7RfIKrNmYp6SdgHy4hliwOZiBvc3DYx48T+GadGbL/WpHuVU+Ujj0X3QUB
6lLiMD63lH0XvtmemmCRVZnIluwSeMi62xuPE2/dE6dej9SDEBqUGQ7EW7F7CH9M
GXR9t/EATFOBUzl7mji1Kcyt9HcVSHaDNHmhRW3WIQy6isBLjTfftILRIGwPiWcx
0MpkbErIf3hx+4Lp1gjJbqcNlZUaV/OyepJcSYVRZ1XJcXI4SgZxO9i3fkNK+Yeu
lVIBrTwPh2xv/cnqiCCiqciUNLnDIeOM96pW8FsDfY4A61mKX79zbe5QOcmy9k/N
KBRfIFfVze5MRA0bWQfHUZIblAC4wYCBef9O8XOxbLKYZaYFXfRAAwroySuSxlXJ
TKDBNjE4qRKvoa/GHRMgLBQPbXuwSCPEKWO7EJktkd3P2TroYOSHxDDR1L8FAXAa
YwAF7PYrENzLO15uDYdYUIRLP3uRiJAGFH0qg22Tr7mxokc1HjMZKIWLRtNYa7XK
eF4+tNxwk6oKF3EIzpwDLRJ+FqLsTmWggZGO62/T9fZ2aLEKtRBihsY3m1u+NTC1
BpwDeOvYNyc6Egquh0U7lF5xH0QfiaD/uHRdVeO86GM/kDVZk7LfJIhY9fiIPXfv
kpBoEkYvcDBSTs3WAhM8mUv1YYwT3n2nseEeC5Ye+PllXeXWueq28gQ48swjjpsY
3FCQzkRIhfhw7VZV+veK1OErRIVOlHomxXMHt9ZOg/qWAlbBVUJsEHE1Qmqk6YEA
tmsucpKIXcTMMjEOFNfp2v57DM0TO1giOe2xTP5q7A5AnJavx2n1iBGsTQ0+rMmt
Voam2Kd7QDVM0Vdp6c+rqFA6MQoyUYl8hJtye0PU1E5epkTDYlJAeX9ZacSsmLxN
dhATwLILVh4rgc0TCiLUnpKP3A2YuCPEVM8rDL3+MVOohjh39LoiSYSld8a0R2f/
ev/NL9QOPYXuIORTYQRGUPt7m5NYSH6KjX7xWAwJMueaRjXyEpiDzji7vvogucDO
3h9P6aKc11HN3N0nCgNIzuJ/Ofk2FHOMVnaeTAT8kVaxcoZXxnQal8tCfEIUka21
lrMj8aihUA33pd2LtHTJWyUEst0ofef+MgR23F/Z+U/lpw9LUXF4vOKW+/n0Q5AK
ZC5QrelS6jle+f8Dabq17BRRvccQa0w3km1e/+WfUJjBixIBAbHAJDKGdr5H9SD1
TXNXj1IKQB5xrRtZ0PXHZAuEkN36Cr++E9abkmwMI9rbCRLB/lnFZTRbANzXwYJE
lQdxV3anmT5U1/dKBf9VfthQP3NcKAKwP4L/66l9i8tdE/Vs+5bodLvfE8VueCMG
vzVge4EhkOHgYgkK8TvJ9nMrkuEXq1iWKDZqiqeUemNtJn1Lx+mGl3pQK3AOKN4r
zeTVNugETSDA7WUqn5cUDJMIa1PeUKwhAs/cYBAEWJ99vBoIDUiQhsMB4ZhdvYdh
VgUaVtIs7NtYqSNrMBW1RMNzZ2ac9fyFahZY9ykmifCfAARnlRiG9EjOXBHt7ecn
3xnwcxqQMllzZ3njZk2UlPrdP55Z0e3ZSLHU14IijnKPSlgL7uOk4fMZOGyyx2fm
EQqSPwE/HP7XGYm7X1GpmCFOkuorryv/aMrXW3YUEQ2a46XkLY8B3fLS+maMPlwU
bRa5oP3pfuf6ex6G4tf+RyxMFDJYElgCV18B4Mf8BzoBxnDI5KXksMtVszEyhiBo
3h79E+Zjzu68ZvyOoMZYB2axp/g7H9Hlfxx6ImyyTwG9GPqg4S1MTwpUTtB4oywT
vNPqoHyo030GyPPwspdD32yKnoLxl8RLTxZ4M27K8f8hD/8N/88ghEkKGhPYlJID
bQDyb3l/gF730IzMk9R3I2k7wVBdzGvp6OAJaVfm5PZnMiQahTm+F1UO62qI5RPZ
CE7OtcPZsiGcTjFVgxSi+vY5mm3nnryLf7p6vcZQiCkcmSuYktdEn07jlGlyRj+T
P6UYANLkXctcZodowcrBChCmpmiJch6FZSk+olxKytdDG54Ga2/ECXflr7Qwit7s
ggjJG8w7jKhZvlgzCkmC9gY+hbJ2ocIoZ6qcJ8F0arRnVPLzcq8dP1iWfpf5+v4p
D2nrkQvYgQWd0W5JK8IQdX04NPCxVmQ/PrKldjuLlJM/zMokoXgf0gmUjoAdk3uK
PvC+L8AEQzDWu5a4KCoUmxKr27llyhevw4lJi/Y6MJC4ENjEORFDDspfnrPOWm4z
brH1Gra6PkjKDQq/oOc0do/SYJaX60NLs3kczJPWz8HJd2PBrXzF82P7gdDlZquA
vet5bOrqjwpMPHMQr3uddL/73SmUOq4f6VNxH0zqDXxMvvIMWCrkvpNNe6mxGL5S
lxcxJgGh/efVBLj1yyzA0tNcRUQFIN6xywT+6kuIgr6cNNgnmBjTgToATiN20Pbo
Isd5SdgWMW/FbsTCmnokTxclx95eyUbLn3u/HKXA/Jg6bXLe6EUFv3lLhKHuXZb3
/efukq2ZEnu2c6MnJDOTBo2p5g5NwBDwqkkchB3tYAkOPYcL0nUm2FE98tE6y28K
NfgCZ1L1D4ToNHzsDGCUr+7exNRzDxeqIqimFfkEDDIXzKtIO/u3CSwFPfkJjxOP
kuf1d2XLd24F3pogoMGYE8uja/Gu/DlHkZJArOPy71fc9PV4u8YvyB4hnyBRiVIy
GgE0fdwPYdPiLdYCqXdS4V8FdP/KQrjqkYoCYmk3ZKwd+5hZDwSiLQYHxJ0//6+2
ID/C4jQxDFhK74nT831uWmWNH8fKOAy/pi5r19bXZG/MWzW3jFC5+TU3b68NuroI
xCc6NcA+gyXZ1bNzA2qyL/tTQRm7ihabi/hfD5odCJnvDFHCne2Re2v/dC7nYytq
vRSKQjh6ob648DO1+9OAPnCSZkoJp6JLoad23tRkkiuDV4XgoO9C5P1q+gYfOuGN
TgfXsWfMgX0UtV87046q9D9FfvKrNUymPa7R0J6i2n80T/4HK9ehE89t9tA0cQ/0
HFagAESsULPYRdjhhd4tit1Uc80BOOPFrwKFxZTcSZEbeXKe2QbQl10DRb3OjcX5
gaBVnc3gIyyuRKNEKlrrEwGgGDNzaG5ezzOnTcbSYvcnD8Y+HocVOHlf3KXGPSz2
tbLgvzVO9wURhk2CTV7yDt5ywbi1taWwt90kQbkYDH1LihD2nqbKoXQ7MU61QMZr
0qZ+bKVkvNHg8vVP+vPCBhdz4KU3+icdt198FYT0OKXSnm/TyduvTrsBndU52mVw
DdcebLFQzQhJW7QTshgywFuPla0e+WGaKqx+GPPmf4IUcnryoCkUoKQPEZnnpI7q
bmmcKevq3sMo37VfYWFzCpPaVxEjC5qQeMqO4PRF5dFjkBds0h7STXbC5+Bvbk4j
Nyo2nbZEJxEoJEE0ZkLQ782ofh0+xVcVkXWBoXNJmD6se6kWXhlFdeKvi5FR55MN
8YL7FPehuZoGtWL7immBwy/6B2W8u++30/3YxeRBmF6pnqk5CCjhh1jBmTY7Uada
qr0HkyeW31UZCrKc2qWH+fOZz3/5w4SBbAp07vuTuAwVLGSrdkrrqgNBcBulhkVc
rRdrN5Xah/KhB6y0PW5vBQwb/VrPe8zaJSnfmZmzvY5w6sjUm1JiqmDo5Jwu5jdQ
OEY6fdcg4/cYpI+QQ685VGKLe0/mnAruikf6eXgn/cTR/l3v6PXnasQ5xKSlH+Hr
odnRxiaeW0Y4/P9EzOrIp3uIr2ztWC3naqen2Iwa5w7zJZmmDSNYbPjHFqXiPLDo
6fIEiS4f6tScsQTKa1yXFOM8gNV0OLFpcaJQqCWEp0O7xyyDX0hV8INEGDP8DkO6
Hje3tx9Ei7awB5VhKhGccOSBOIgt2evleeJqzIYvTaYNPZA2q6O21Mj2/1wO9StI
48xdhOA7SoSuN6b+qpJ1CZWlA0FdqnyMtN6StfEjdIRNl2WRGC/xhZ1jLFBUSqDS
VBdCwBf/CgtkUbz2FmInM7/3A+QA0yYUa1VTbo/ligcucWOCgnNma/FoZxsZgbJs
fy8ev5TBctfjrEKz3mH7Ml3Vua8xgg1P+1/hB8JtU1OKrWxAP6mkrr/oFF+4fkjC
+ODXoitOwsk85VyW08YzXGcdpQu9EKcuir/OYAlAYE3yX1TGKo4kbM90ZIYfhAk4
j0tLoQM9WuE8bQ+O5+ngGs7QuTbwoI7Rpys8MfANPKW/DViV0jL2aMrBAXzhlzr+
6oDrKsgEye0ZVbBYpnj88g9dOMWCPzS0IN3mEKrgiiams3pYYEF8nZ+UTYW8DAfd
Gp28wqxCk7KciQq8CAse6uJpRyE3e0baFoaMYcGqf0yQb2lEMi23wcGEPO8IG4s4
Ym+qHy+st4IYcdMjwNSt9tozzTvNqAnR9OddAq/F/mMnRYo5A9xkbWKxeqDjd2S8
2d0879ixm6D/+ErWrJOj7h5nXnifGZl0hmQmgHikPY8lLsrEKInY3dJn4CbqLAT7
fuU/+ngRHJXKbmRCO49T6DVmRWaI45RKRXBn9fTpgVWeSONvsJqegn3Uzv0oUWV7
FtTIvVZs0VO1vb4opQAjTaityumSuyr0firIEmPJy63S5xBjlMcYAMtV2qII+m47
4cAzp22WV5SZTxGAeNd8PQAxKLRWsnF/+j/E+7gVVY0ySKXGNMyMCvIVNrZecH33
Lu+S9nSIAZCLyJIINcRB+owtNQZPNzbDCrP//GVhDufZDf2g1nU6FKItru5PD84q
F+Msm5/0UzU54u5PGkfd0YD6QrdZJQYsaGje9r4RoNLnyu1zGCHqj+hNgL33X3Oy
+q0aLfdrWdzo4GTGI3cfmTgxZWZH8AJNk0fhVFIutQbrGiBktbA4MNdDHd1yoN62
gT+oU1uLbf5fDTb2AzXpinmnsEvA3KGmC3wGWG3MDjsuQpPIaM6QkeW/eSdR48VN
Kc2AGCy//Prd1BZt15JSffIdqu+HuB2ckg33ebqp5MS7k8ptUwz6w7WeGQkUfboO
SK8iV7tIwW2u8i2hZBa+ULG9ki32cR9kaSClEv1Yo8mykcdkkdvAY2jRXNUb6eKE
07F5nziV4AHQHk7IiA3036HAvFmmz7WJOe0KznRcbso+VCPrM95t/qw4Uuxu3nJ0
hUpb0BznAp4Ou2OaWzkLDqxqO6Aj5xa3WyvBX13FmjQtYppaixiwqNf3i6NHa67y
/pz6rBXfJEYhLqmvmxmGF7DE1o+GxcpV7MgL8lOtFNIoALCucMrrF827MPJbgUwN
uYZLZF0iG+7zVOvykqVlsenv+Rq/nAcuGsag0mLPfn4W53Q4yjBwQfZHOc+poLoB
82kcEL+6XgM2DM53qTZs1SEZ++sPnDGTMKF+K01Mw58pYfRoST8B1jC2PiwRx+c3
LF59gonnJYBialBPURDSUp9mzHeMB/A1Hafdp2o2bwj51H1W72MKeEBDev0EIpMP
pDXBDgWYaTwR/GIMF/J110kA2w4UZT0TZHAB5ZikEnT17o8ZQt1Ox1C27w02N5uk
6xuMg/j2XCJ3KOUI2eSeYY2d8mJ1Vt5UNr1GHPYOayp9HyWtl8hsnBqt1zZHrfXK
IhSh+5Xs+unYbo8bBcSjtQtInHHNxme+cwurFLpr8EiRof570iw2LFPWzLyzE8+9
2fJwbbHeUKIv6RbGAp2+xd/Z/D8ezrFRAbh37fW9C4rMXVMh3yExcXX4tM92AZAH
zNuneDhJd/j3sTPhM0FWWDIxngV/K7I/IABrUy8hqUW8xgvUymJZo2rhIZgTo9fq
QDtaGBjWr69q/9whsgUu/WO4BU3TBEyDxWN6cZUZQSdXgMXZ+4Ulg+6UHXCUnnJd
P5SEZseGs5w70uVT8SyspRhX+21LA3WxtRMpfDyM9B/zytnynUtK1bOw/BTZJ98t
dkUum02co00CGW2Zw3w+Qv6xiz0pREOsXSBUR9Kxu66ynAgauXkcY+7m/vi8WopI
3z+Bn+U9Z0suE8iAbstp8Y2DIi8XmJffqevlfG/cs3b969or426b82XcVLKrTW38
bkVHNdNm2Tlj8CdOrMUnSXmalklV85WXxsWAlkhLfD3syGb5P7xDb2E596EJyAWE
UO0yKMM3jPfxI007xVOpikpeaxYh/lMHQmWd3pkZcAb0QBUjGuNWMZWEfwTTBeP1
MRZFod4ahJpebjXDMLHvkVc//MRWqVLOP7NH5On0nChmQ64hTbNQOaG9uxTwfmcL
IBFvNUvnnwOevz9s7UPepyZupXxh5f11faBHEtx7jdb6ta6Aj87X0hzLzY4Q40z+
FRJS+CHX7ieKbUBtZT1dWATyAW23TYghcK16z7QbkHC2XZkeJRwMSbymdZpzNMZK
QaUyLHHFztfKCgX84aMYIGq3C2w3BJfS2+fCsNcZ8sHk7wZgw213o7Wv6+3q2Lb3
FzSIVnPzri3nqyXalh7Ixm8j7oCfk4IeLR7AJ/FcDidoEit1Z+yzhYVzg84VWhpT
8UK2hTBqX+Dp0GYXrSj7V9orkap//JCXDZ9pj4yUC11DU3/r+QPT2x48qNq7wRDt
eSiv8Nm9SqR57q18v734mnBEG3psTELERPmcVStlttZ4csyTGj56yysadPr0DXKx
IjpXtsrWJRoeL9DCzxp/t5AdkLVpnoRwKbBs2mnWDH3Oc6H9uV7tGE2Yw4wVwUkL
LrBy+JtoLv+iAzqSkdsUCQee4XwxlYlIcA1vW+HWSSOn2MuYwTVn/IzdXh6TCn2E
5yFGnxB5XQeKxdqf5DUpoVpeUfmBkRrEjRGD+j+5LMGpUjvnVnPE08aE72zqkNTO
9j+36C6tN1YrLcLNZ25LwwehnykCsikzGTRJ4YXZ1ajD5ijfQn8hJG8NHz3ANqv5
SKfjNZyioJTIg4+UTHi1Lqa53eILZffXmxPlSwifQj0VWwIYicYdpoEo6YZYYkET
UsnO9LTfr3RuS7LtAFzKujXzF6Dvw2+KUwuDQ29PeirReV3jWtoq3Uq7bHAMwODW
WsHZsE7nCsBH98Ir2DL8pJxf3NbtTbpofkafQqBAqEJz6C+0cw4g7rmOxAbBCzQZ
+r3xAzxgeUWaYzWZEAC3hANIRddxARv0EU8N7p3QELmTXxe9UuaQNiAhzsKZadbq
SqK2SnBoUmFlZU1t2FDPAkEnxmUVhY9KqVuNZvsVc7MjWaXym48h/ugDVPVyDAsc
Su67bYEuEQzHE2191HhFkZai6z/he7+9cHFm3o1U9f0eeNE7chV6oEg0rbH5f6KN
16WwOvPzVcgPwfPHhUY1lTTeM871YhSMvZj00sqA9MCWTRzyhBqFbtc8VDGK++SA
zTRt+BV4RZJNlH73asEjxtTwAL3QSWldjauIe0niYlZ9COEY++iQqy55lTdxaXU7
ozv/UuC87g8Ml4rc5y4V+8HOLjwXoYnIQ1iMfJGKiOAseOsPrzyXKfGZtmkHvGvM
dkLZbpn480RcsowHYpvCUnZfFSEjQ82OeTdzmkhrBd3EX/EyHrbqML3PhVr0cgTE
pD8MQ9wggmh9aqwTJmxvyxMviupEPzSvOFvT9skpZ+e/lWsK6uzvB1+ssdpJ5rz+
pQLkYGN9Wu4Ddw0A3+g84NLU9rdaalehefQcH+MPdcA7Jb5EpDx7RL4vyxHy14oQ
Dc81ms+9pKjGycYmZ2HAhYCRDHc1iUHnOjUVmVmiKNSIYgfqvu7PVmxh2l0MbfQF
Hi9lewdN2ajya78HA8lUHIAiwpzmmw/OySCIoUY1+JVNPUWMfm1XX91y+Gwcs9z/
f10z5+wQ8JhWAKKUuZyfl4JCn+EpblR0O8OjWNeI2jVyOGrsCbItWq7Npyllid4U
5VKJywTjI0rTvMVgbYwWM/D+Rg65TacIozF7KXdeQgOkFyZeMxhzCobad3yoMe1q
67VQHR2jgMUmdQdkvEzyH9yte7WIrYjPOYlwGUz54ih7VQos+1pkie4sY6JouoVD
mYfLhr4w2oKoOEpK7HA8aOKxXvdDr1YfujXwcvm8OSXzsYqSVeVEpLzdQrx7rybt
pD0jmsl5WC5/DFl6/e8IciwRYM8nC2iHqXJ3vfjzqf0rU4UHfdpqqbKpLyqiRfDu
Rl93Ma3uc6nShxOAHX7B5iFRmQlilEq8d4kdkdhSBcmHdssxo2qpyk/rf7ExtqI1
/+R/G/uKT74qx6tmfvHVdRYaOeEPYtc3DjZdoKQoU08q5CjmFdjAxKX7p01O8ojI
Igvdooh+IQkZV8nQTDpJVRKg8ASTgbrfH1tQ4H/ejK3sdQTZUwPDCR1nLbs+lGiX
sK0nvxzu1A0v2kE77cd/Ummvw2zWddrVo3hNSfIaPMYGklNIx9LzDKma1N8XMNZi
YkBuUnnl9rz0b43MAKKI16f1v4IJ1skQBLahedUMIYznNHDtxeFyzEPZOk0jBTmU
Dcf6N3/6qEvtT1aijpRUjnBZzdFWs4HJxG/oOzrrfpMZ2QmuRsGPp0u5h04MQkHZ
+yBIJxpr8gd7tQ9HmbhfZ4XyqeozFBt1rhmi3k0bsUAH4ei+mxQvsO392qBs68b/
GU76huPuxYEuFcNhhF1NeC2zRby14NZwRuLPfj++yULxayTQqOHPpIDs+sLQJ/5F
NR7AXiYQKWDk399dE2IeINyvSNdForjzS5qF5Eh2BWvQHFiug/zyqJoEUAdufZTL
AjJrHN/H464FEVhTiLbVd2WwM6Vt5C3jiUKjyQ/rIBXCgkVVUzHKtiry3pOw3AFn
si0jpKd9cpbCzdUY2TQP1K6BMYK6236yMnmBakwkU1YazC70CeCOpvLG97JSPaqX
/NBbFJ4JMK7j9BGVdyWeBgaNDFqGj/hZQI9k55IaXtjN7Ou0oweSeAGMU4UTrIh6
cUCuTnQeI3u9k8IgtC4lluq/rxaiL6w2IgHgmJArlswmC/0cPkyIj88ffv7oiAEj
2ued+m2NLnc+4pxnk0A4S1jvetewQMFMp8rhLchmyNE3PlNaPtLm/xtXfiVx/ZIJ
GPbf1KI8+RKaqNUqpicQe0GVpllNXvfWDZtGzUkOKmZbKHnh5uIAGX6wpD1LY6wA
XOsxCrDNpxI+Pzo3jO/CXBEgqt/fZK5AlZ9Ranfi3QNCZ4XWcngjO0jAwf01Lp6Z
tXKkTglWmG3gQ+QDJjqmdjipG9ujJz+BCfUFdY5+zdOqmJU0tRfpf/p9GPgyyHr3
uqxoXZHHSe6/e+GubaZxkW8B5CoYEmxOV/+mLXkyyXTZFs8yzOyK952Xkydgj4dq
+CQtxh9//go1eVMqAeZAredQsdRoOVdJm6OJR9hmAOnQ2Kmpc9keFoSTACw/KQX6
/J8QUVxUssaUOPNC3ItVjhTi0YHX/0Xhd4azhWNttR1WWVwPxF/buCgDrMbF6qwd
rwYrJf2xKEqiB/CuH3vUEpbctrkUR3zf7ZEbnBKvD3NbMZoHKpJGVDk83OpiVZ9S
Ofel/LkTueiQzaZq3xEhO+KS4kCMMoSF2NET4fbRAarMj6eq+V3fC1zqbW/0h11U
PA7j8axN2q/RVpTSI2laFvnXpYlwmO+TP9bFw/tVpQ4AG6xCC7eXVnQHBkDB7A5P
nwLsqQbUYSpraKbshYjLHF60lb5d/DKciO6I1JMK5FhNvav8HdHXlakwhqPOnd3H
u+V0TLcbIra4v5aEucNCGztpIY5xObVCbfbLTs3JuHGp4xOSyFAt0VwV1Ol6/Wai
by+VqZD5DK6gI8UJE84DXZC9/mdUaWVSpRhg1Jxaz73q7VeKVxUcD0wbeaqSBATL
uMvsR79nDRUzNOlPJBa0WColauaPR1+a9Z8etiytUca94J7a8r+7wAVAdduH9g0W
RidvqiJWYXkwFskeDs8eHOoo5uT1mDW8WCJE/Qg5RBY/T7+ST5DJr7muIp0AEzdf
yRnS1Ggs+U+dL4e3NS6ntalsAh/dn4u9JfHXAiCPY+gTJdnAer+0m0kf2wTnJ70K
m5FH0Picwl5xWhDJgXG9zILDatBp3Ygzy3NI3KWcOOxBbGRT1HWZo9nU040oVSr8
xwFUqc2xoPfkTkAil+9NX0+nR7KCtgWOHw8iHv//yVPWZqoIz/6ScBDN3udCnYxa
cbhnB6S/tCs/7ar61bETB5jKumPCL/grBvfjeACroAPD0c6h5yOqHs3uxbBPsBpr
MBJmrcbGFsLxdpoeVQM46wjtk6qqHdGd4qufLV+6G6lM/f7XcCDIwT2L0kR8OqxX
nDElVQ2co1rIZfkHOncjO/fDYWUZYaQn18nRQtST3kCuYjPie2CAdwdESTfwVrQr
xG/VMLo5CVoeIRWv7bIym775gcOIHxHzXL4ysZnNHtGQzIx8DmrrBdjLLFFzaaQn
PuZ4ZmxzGfAb2bZ5U2UopmTwWp/Th3eXL6uUx4S7Hxw0e64h3jRm0GW5tayFLYYn
nuPaWo9LgSn4d119U++cUEPAgRKb9X20gR4v4EXvyjqeJbHTVdPrzBRxN0hBDCZP
TLRUnSGrDiJd4NxHJRK9cQVXq/+HZOPJ0VnbGgP4ZCApeZQU5K0FDPfr8PiSI9S1
Ys5M77C2ovbSOrINB74DwwQgneUQKNU9EfMBiTnXk91OpJsBvIuwFLqVPu7JcKTw
iwtp1XEslFYOAe1dz5rZIUzkzH2VqLs2xFHcgqHEns+/aV1zxJwOH/JBd269jvxm
bfxz4SCQuKSJwbkSlu8O5RMZfJXE75Z84OwEYjVETnUxqabF4vv9iCfclwV+O245
2rOIhjCUM7mDvVCXj/xMoo0AAx1y9bN6sypMMW/nnnMWBu+CWJe24PJ/KqxZY2Kc
MKvZzB9xHkdJoQCQ8Qf8xVLxRiKvUFD9Bk7DVQ/Tp5081CDFH9oIceeajMVyCLEL
kSb6wR9Xj60zECRdIZitG2UayxZMnH449zRt4v3ZxB8ANFJ1cnKcteRKlc8x90+s
oCBFYRjMJSIIXszCB1dUJl2xB2b0fTR6uFVkQZlyYPUwsRbEPLauHJ43cwWw0AmH
aMclV1twAZjnX9FinRHd88a2aDTbN+kKTas02yIiNNI4TIQtJidV5RxdhFxREXSg
ZtlbUyBD2x61PlnVLWGVo4yGhMRKBvpqtceCavFtxgI1wWL0T0O837s+JUBp4Ww6
7s7RWjbYYKNx0cG/a7VSvftUkYdgxq2EEOEHYegu6bcx7TSN1Aj5iHfd/S/s+744
/XXaFEGf5s5byx+sBM5Bou3B1n7bdL5Il9WC7GCSmkaffem/3VXUvH45NU56gVhG
f0cHu7Simnnw4I0bKNEEfJFCOOvFQcQJ2HtRZ8J+OSaIPVKgl42t081j2NlAY+Ys
y7pFpTymQ1FlQAouKKNecVJMNHBppewcheN8FvtqesEzNjndVWpiz6Kc9Wtr7dBy
UA4kdZkKgPLSn6l1DluifdKWueX2ksf+HRiNa/pLEQiUkm8lr4BAf93hRIaQl2tA
ZKGJa3MKrcjMhYAKKDA8OphGYTEu8O7nC6IqL1wXlQdt0fbOC9z1OUckjWtvEgkv
5FWI+Clu4+T2zoUC1G5rmyJ9eKLc017zTYh6jNHrU++g5DfkNOua8ry4krJnEJVG
9xeeYK9x/WWMmi0jkEXB+HhkrcVwAGzexu61t3lBSB/cu+jVmSCVlTrPcrSuZ4lM
h+teex8cB/+yNXSAvjuNls4qj4EGqdTMvev4t+2XaurKL00qTUpR5fUtEgZcrf+W
wZYJl2IxdvaAajYGF/QxsOjCF45AR/AXMDtwxWbdmtJQWXlIxSErKrMlc5iucQ7p
5eeZesJYxxFIR4xh9GJ1Fqwjh0xiVNoLE518w/z0hudHd4KM4VBrnKjkwz20uN15
iOxhvAVJs7x/MCmPJD9NRCgkUyACuXwe5a97yzpH1u4NNCMcRA9DuckBHnnPYRG9
9nH6kQBYZVH7hDK2XjmxCx5fvGkH2Fyhp7D7inviAaaao3ykLZs4lEdg3MZR0GSM
sKMRX7BUsWJ1Y1cdydDJx75YlVGdY54pBmQCwfW2YtUPMNMJMpMTgwN7LwhUamQP
sG5uteST/VdYkCmDGwwKWqEMZLyP3iJ3XAbG25VPPhPci4RUoDqmtx4eyAAY4v51
e0VvL2MBWWTgNkj4ehtuUjeIReqNT75A4dMQ1nvahjW42N1BksldOfyOz/1FWV6T
0Vr5HmZPybPV2w0T1k0+JQulwRC5D1cYpLvtx5ms9dL2fAmOJOPW94ERwLig+PTn
uqddYdWQ0PluNAkHU10PUJcfkB0Cyzlc8NDbinRVDF9LV4vOV2NCoYX803r1lV4X
AzS1hori2UbFaHz7f44q/35u5DedOswsHrJoSS80IbzTmFXotIJ3eh+BzNC+kK7m
4P/wdoodZCaMiyqnnkcuHqPyDlcfvvxQek712+T5msesZcm7OnqT7NNk5r6EIwpp
XtGpKjuCA//ZkKJ1B94s7twxXhjj1AiaCZtqjykXYlUKV5mCIgQ8zS3Vq7eg5qnL
XGw/p9Wp8e1z4oDDk/BnLK5b0Kq5FFNnv34PDU4yt0xTSj5x+BiAyzURjvW0kV2u
YbmI5CBtSiuuXRhdITIe25zacWRs18RmjnYFm01JF+DBYsRughbPUh7dhMgOf9Vr
w75gCBDvmLt6H30wM1mu3geQWqXmWNOfUjVbL1ReWtsHHOa1OrjBMn+xoKKgXz2a
FgmNi53AoEmcAiGspsx0Rieqgj+DrKlF67MfiD/FFnWgrhr6WG+oXucvooL+OfSe
4E2dDSNaQ65Q2DSFW0HmBQPgVGuVLVNv1KdthV8G3cJMUmAraaB+eaAXBxK9rW/t
JgjBl8pzd1D+ZNZrPT9FE5CHCAkZZG62iLZ8TThInbDnpTsrvBl2Pr93JhQfBtLh
2e0bVlP9quj1PfL3QZXQwYF0zapdBSmbOFsbgPyAjbu/Ay7v3GoM5MxY6A1rL7UU
pblZVuzCCuCkWp7B7bBiS5QldvA6HpXl2Mn3VJ5OxIByffk8CKVUT29bcLyQ2c0l
TOwtcVmhnR60bMC6KwmydePpzWGtXFYsumdUd/bhMhiGm0QEr8N9As5JX/pOtb40
FckII1qgom+mW7ALTJVfLWkPQJ8Ok/W1Rl7MS73p94vv837IEEblkn9a8H/o9BfB
BhcU2O0zFOp3ks31C9ICOvg7iNAjMOcRQajtSPHAeSJnhBtMk+epTmNEIfNPItWk
P91jQqL9bN6uWSerI8l4f/XHCU0+XC0onlst2d550ssmVMV9GLdAzvZeNvqo+4Ih
ash6kAIrUrwaiDX1un7X86vcBWaEES/Br5MLc9KKmqjNoHoWrmqYZc1ggrL8nyjL
xWajeYZssMFwMfh3Ph3/KflV7fUXTDf7Hh4JP2cj0ry7MA0nE0uR3pyVYRPpDtNy
PMLVaYIp8S/KpTttThKWsFbMknk4ZPv4YYz5XgKv8G9nOjUkWJu8v3tMq/TA+kiO
e+k5th5NcwLqF6a5haj4M5Ky/okvcSordu6CZWVrCqHhI/5iDo/IvPU2zureNI9D
7jqmCXvDZTLPywfB1AYu9UJUnxFRgpdOBUHGx5Wu0ozUN2c0Zmlb6vtJMa/iq9R2
UJ8ZMnHbs8Gbiwg4R4PJrWm+dA2fQdAz5PbMhxy2E1g/9KYFTZ4XbOABc3SvlwZC
30g8LKXgfw22HqgKFbHM1p3DNlswgEGjqS9snCGqEiNPX5x93AGpbUni8JpV+Pmd
qecsIKnmM7Jcact3M1JDaVGovvJR0e7EqPcJZ2fxJ7D1l6PYT2/CoLP70GemzL7h
OiqFl/BswWwAN6sKrslwYThJD9Y32rnzp87Q3kt2stuqlvLthKa4Z2ayvsoN9Iqu
4Glqc6UxVV0hQJ55DZTmYX+aNGcraxwRj7X4fXXopfrBr7BLq9eL+ipumhuwD6vH
PKJ1XIdheh5oKjiUhw+t2wKmNNiGviZpruPBMPFwcbzHSpslfFFRi4UpsMCBR98Z
kmHICEQ4t9VTH1sjwnFjEcpSnZqhNX7d3hgtoVhZ+e0I0qbxT4VAvI2J3Eb5FBC6
8+0ajd7JUxYZ5GD9LawqVQ2AW4HpGN/bWskwM3ICaPl/bw/61cJJyrN8Pla/nBYl
ja5bYpB7Od/480PuLutNem+XLFlrB86P9MswnHdQdOruG+Ff57FeN4AS9LGJ1vir
5+UTiR1My2Gl+UqG94ePqjPvXwSSURMKs9S1Q/xRJlpWSaedOw1t5Mnwn8VZyNTk
8caI+iiXnp3uMusbSDRjVKbqO0Gp+OQC+deVJpt7zwbd5PoZ7e55lWacWM06n9sD
B74iDEd46Fc3MkGzc2L1V4xA5hl0Cxu8Ebp9G8VseKRovrT1coj/5xIp6i313Ijt
FE0uKbfGQAlWAn0vUCHAJpSOWcJlUACBB+Q/PvtzsPGqA5Csx4gpu8Mm5jQMfYQG
cHllTBG8TrulNcgK92EwIC5TuO4w1zFt1Z9URLNMJbEp/nI2IGJnUO86fCNBVis6
nF3NqJmBoBV5WOsWcnJapdGUz4xRKjCjFKhun+Umw8h7JF1o5kZiiGZSDYryTbkq
Imj8t6agoGnHFhYan1vMv/PYw93wO9pDjWz+rHYSrDUjikX4H5OA3TAxhJsP8Se+
XTnx5rWhHnEwYdUphu+HmOTcfer8XJdhlWIDQevBjT6caqw7lnRj0fk3aSYtjrkS
H58K8lRDYkl0OzlpoaIdhnwWGp8aMo3LxFJ4575XLcGoqzsQp3lmjI8TZzW26Qz5
0o3t6kht6ULtlE/zCMzQZ0UfiRLKZRXZxCEbkg0cQ/Y2GjR93OKe7aKEQyWW7zL3
UpX4xdkmuP+xtONOAWZacZqARtFWwRlpm89SrsR7uJB6E7RfGkoC5bB+dP9QUT9G
782MbkjQ+haXlAPd4yqCFj+yGl5Jf9W5qGGGZRYCFabYQ7ldskL+mvA12oS7bX5S
HHFh1orOmUMO68UAfT12FtWVpB11Uh8qJaDT3P4oo6zTmQopn9DhEZwo7DYbKpfO
0RUPomPpYVD7SBbE5QNdSme6wOQf/ABrB2CWIPKyCU0HbN5HcJEH0m/GvzOtjvjN
22IYagRJocWr78gWBvi5OzMCQiJJbEDmgiqx8BEjoxNVoDFSkY4yFikb1l8/0UUk
GwtBqjG5zAY59gdqO19uLN9vyDkb7FXtLRoP+n+K7ZiD87UxI40NQduj66roIjds
QbYBOxUp9pUszfGFOn3nlvQEmYakvRWOZ+nfi/WP43tjZosGBUD3zO1n4tQr3jBK
q9mQBF1fzijSvZQoezgUpi/LDcrfKRIITgLJlRmbz1AEKIYinUc5LiuCoKdC78sQ
R9sp72ubYTHRjLGRmjoHLXoUIrolC0mHh3hno/fgHnfku5ScxkvpJUtyDFefiNUT
LgBxExwmnXY6QFH9F2f4PcTiqecqbS9LagH5BsIXHCcgWmTb7lMG579N80XyOvnN
hqiXiWanBtCoIEmV/6vIJ6gGsoBbHT4NC9hI7CEIgTMv/12+hhLAalpdBPkm+1O3
XdQGbi0m8Xe8GUIujyQe+A4/0+psMca1CVOtVk8augsQLGkesoOPwxUPWxNVbHJ+
nxCO0ghtIEvW25IHuW4kKQS/bkdWdb6ZsIBK1hjv07hd4f8mIFakdQv/6IZzTx96
f+mqbEf0/3qJY+GHosW1FJmapDhFaju0iy9PKFwiYfM2vV57U9Wi/xM7P7pDJSro
FowhbYOqNJDWYR1KKIZtC+LxLc49DxLVP0/+AE2RKOgWrSV7oLi2/ItNt2HNjOY+
6mdnqv7Ngp7aGdn/uvxnBWDRx8MjGDuAEpZo/AIN9DjK6LKwSsYMrFGye4tJMGOr
CeHIh3qc9l3OuSMkVYiAP5A9F28g8W6t93MlEPl+4aA/kg5xvP9vSN2IrXY8uIWq
XO19+KaSbt9YqvRAypdCehYXe355tuXXbduS7lIL5xtiF1otnIT+xd+8dq2/Ehd7
NTMXavrHnpVqUQiedwojywQdfd7Im8GErZdklWOXdi0MumQY69WskHbOo1FJ3HYj
LxjdmJkm7RBQvCnYtsxLBj1ZyLbZiWF1n+YFfK/xiaodjbwNbItrI5XE5SxoUdhp
cpBvZsXtoqbng2ycjzi7asbgmuuHkwuiXsBx3b4MOgJZiQwO5CLuD4q3xT72d7Zo
sNLPEai3LX3Y41YzvMga7HmVFEYiKs2Cpai0EuohxQ8GcX01no92d10Npxp0MNIH
CWd7toRF8IJN49ClY3hNpmTAIwcLpyUF5FwFhbocIwiuVnlV0ehcHFnmSiC0K3vE
uVG0asAwmeftWaXumSTJLACf0s1gki1zN4idh3iWhHKEXig2+HFqntUQm1iNn7PX
qf5nZyAwrAXIeAVH5KvKrs3JbF7PFVpg4O3MBWOGIgOWqpjR2P3sPBrwH9nBPlIf
ONP9QND52WP5LCUxRoqnYVNrWIJfpzyMM87YwI0bu0xUXstZszCT0hJ4WJxH9S5h
7cxrZQgxGnCKlyv756w1PtYbW3lPPWY6T+aFJt3/KfuTXr3cXUj7m8TcSo9LmeBC
rTVKn+D2sMqeVkClEBaxJ7lHPQKMUiYmryyt/IzmBoritZii0tGTkMxC3r50BsdY
pnPffaWpIgcsP7quwCj5PmhMl1l96oHa5g/As/xgDuB1hZdtO2bB1SVax5xH8qgu
EbgAWacenG29nh5WVKxBaZyW11Fybmj+dndVb9ZETVGV0l1f5VZUpCVP5+wAkOva
mkSpR2U/CigDKSZl8ZsRFv6XtBO2ffL7z1vgf1+9gPa9nkli8fv8RQqN1LHZy9A+
/kBlLR2eZtYUwgGnLgTOp+VQ9VXvydE2uqxrG+FH70tzW2dOk177pgL0YOHzAtTj
6EVPGWNQ01HAU4/7d6Ak2nUk0DVwOXL2KzUYdYFKpmHqYNkHRZqUbdqf9g3/vjus
ifwjTISWLRclHbIbBbNzelyEAtj+pO13jn4dNTDyfPFGmhwZPmU7Syt2LCJZ+ZIt
f6Ushf+S6GAsuxWoLYPF7ZasKx8I1ijrxUKZzCHG6uDz6TA6Uq5vkxU/bjKPOEvN
xK5DXZhIGkiYxT4AxS86HbblQPQ8lu53tshppFgxv3dyh+gdXMau+Sg3n56PS6Uj
3Cx0oPJA3FrO14EtWV9/fFGTBuceq5dooMqEqH2JEjF5x00/qOP7QKFGwESPzjyV
q6J89mbGzqQIsSAYnMiOxtaFteM+aIAuxlc6xyVKZQxzkCiN/+e7E9/5LRhIiXbC
2+kv1lheeoANQTR2WnkwkOzDU9SR18XMBUMbxfojsI80Ettbb4+LjJPAenM9ySGS
r6NJvBNtg/DsZje3U8ZNYUQAIkdoPOLSFr1HQfpEBcRd3lc+lPsv8ICm15Q3s3vp
m15HSI4SFuCdqcvBr45Q4saxPiXgMtZpyeYK2JWERjZ+jjh/mOwhfsC6pj1uJ1UX
z31GBH8lQXeGR5dE1SUjGAg/VvKH/YToiald7flpZDREqile8y7Zf5ydwzC9rpKo
V9ObCgsUg+agFUuzo1BibBsis5bOm+Vo7nL9asvbPBa9RHzIZuwOE+8Svh0lmKbc
bShlCJlNohZ21eXQMWxMl7BnHR57I1qPjyOTo4I0tfHcyhwC7DRHFdtRpkFbB+7f
RtwoSckGyzv1PbsCaN2LfpRAK3hNN3Vs+liwor3f/2J4VjE+W38gBKIDmCbymNP2
P7ziCONNkalVHuBbAFQijcDh7qSk9dGPia7HCmKrFs3/qYa37OarlWYkWnQJ5UA6
XgrKFxDngImZkYWkyUVUoaWH7Vl+/iVjs+4tZvV7EcVdD8UABZK5DLu/h4Hu2oa4
0CIZL0QuRfbl/ojF75GLGtN64LsyTG9l/KbcPL/BhJxat1wgdDvxdsPBxcJ0Pkww
S6ebmDZ0pWWbE8ls8WITs+NdH+qlODh90MW1ZkGXIMzocT45ZYzwnkSiGyZXFq2n
BnIXUMdF/4P2DbsnNmOeCdpQiymbyWPMxfT+xzILNYUzmm5HesNNd/WeOQSHmbQ/
elocbxrMUo+mNQlhFu9UhVVX9hItiY35PVdOXuZQNhE6xfHP+kffR2unf5QuxVTV
ibj++Q6LmQAkAfQy3T3ifNcqGrpRhX/uGmq3wJgqx0cYU/xZLQTzsXUsxGzA+FUr
XMohKNUTppjhl+oNs0Nl5bVOespqf7hSwcnfR4bXJxomZcLgEAQ2VMRuXkRRodMz
G/Ls7umWaA1ViBF59b/rGjcgpf7YxgEXvk17ZzFmdqiB1NbdNNww14Jakkv1/j8N
Tx5KVG1fDbo+CHl5MW6fpEW85UUQCrSLCoPEjufF0yDmhAl965nnXcOsz3hOV8Hu
fUkjqSB0IfmXFK+mTjOb5FwofagftndOqLIpXy2X8A+MaoW6mty9TGo7EIsfFO1C
4mMCTmZjMx5KzOmgfRLlWeDKKfkPY7/RwAg9JF52sBxCP5KVx+qRFSSpI1Vhm+tw
jaVvqcfJwMZZCsSDjiYqFdPgd14m+Vb/fUG3TEPkD6NIkwByQ09jTO1JC/00lBKO
1QcH6Q/FFOiHRrXa7CMowi0YkE+aGAadEv5eg+QTMJyYC7N3qvvSX1Cz84LbyM7x
9LuCWCcj98dW2KdaC2mpb6yRZMi11NlronIdzsjfvEf4rJ+DDAsz820pUZEuKdPW
dA3/koPHu+V2p/dwuZa83aNxkx1AZIuLkuc4w6QB7WW7bpo8KZu00JpFLOx1D7Hv
ocSzHjjRBk9+FHElVFNPskSV4N1slc9uZY6CAB9aWV6f+r01kG1MC/BgB3yQB6Vv
+sdmCL/DHeC4RgRf9COOAFvw7DL/W0ksR0D4jatf5NpBxZkxz5r0lq+bg943SRwE
Nxer4Uk77Dy+4xANkeBdJHej9ptywIUb8KSsd5JNV5maIn0vx+DzjE7nsbBh1mNO
tp3z1SkEC5VzlS7XTOMhGtxNmegGXM7Kg6C8fguKFJGWpkpmsnlGMCgESQylATMR
f4EjAYHKQVD2L68sb3Q/lR7b5Ntu6ROAprAykZBjIkwmGKYD95Uo/Z6BztDO++og
CB0LhNLfXGApmDE7pkSLjU9Q0qbpKfPRkzYvNbuGFNgvexMCbscJwErtA3NWMhQe
+U1xR1NqSeb7nKmGN39FWDOZ48jAYY6lzqKcMVIIdIx24N+W/gPif4N2Qej0DhTE
T1sdKM4R2jFCYSjaFdRqk/nU+XHXpWMWxF8lUPciiVqJsDaJNGHnOa67Sp7FqVx1
Z2Z5m3ioqksGKJeC0WfN0/D8LypBUAtRZAY/5ofLgoFdc2mQaDUxIRPXgNXgO3Qc
IbNFdL/EcYYGuvqRRCgNnwDzYKodYeALrzgxbV9PKz7zze8jBHGGNMcPI7VPPh0n
zVLlvz8VBv7mhZfSdjPsEG4rsEgY/w2pXav+HpjR4LIt84URoGnKxnMu1ZKzpiED
qqc/nvoMpVGhWHbi8hExrxSnQ6T2aAO1qAcRvBJ0KuTVcc32QZj+DlgPRnEvuHp/
dU9vd4b4VbnqcypaodCqO1jGPByaSY3/UPVG0x0Jf5grUda3XT7qkTzT64xtk44q
/iBowiYmAvv3bN/8z7C9zGIb7OSetcnw2d4N0t3SR4oz/VSAW//E0sN5zkVA1FwR
dTMtf04twlWfqkUoGjOIU92ekH4svyr4IZFCvJHpwFtLFMcCIyAXrz3A6vEElo3U
ziobxG/o8xrt66RtyXBwCLy9qwVoOt9BrHUAbXxutwyLBGGbLjmOgsqrhbHXcN+N
vvFvwNmp307dXp2wmRKHAhAKPxoIenCHUjpSVXkJx3sIOkaxp0WCe8Ck3f4DFWOg
Ou8jc4DJ5q0EWLVpeQoKS1GI8xGSPC3kmUnfYOK+/CEpOpEfAnfeKEL0HVrc0naS
F4BjUI05JSHrmjXcQqK+EC6K0kFndeTKUNsG0lAvWPAzU8h712OBWxgc4ULG+LNn
/DimsJH0LPDFCuCyevNpHBF2DgJc4RMY8l8bt0szuXUBdbJw/Op/p6iCJ7mYYymD
AUGEjQVMFg+q/7e42H+/d1eXoiZ75ZSmXYX4a6r4+0Uto/JEIcLwTbRo7AQsHcrG
GfY2U/tzQT6HbBFs9wQTqET8wdfTsbFS02H/PJSFzBY/FBg2pDZ02vV0uVA5/AU+
iEc09kDwot3IGMQNusHVYxTMt2HzrIHIeHBIR8CmesfY4Tu5MUhevsCnzLYdVxMk
ctwMyCrJc7N7F9c8xzVd825Nu9kPFZQmz/JVncacXPe+8ocGEV3x1Ri35HUpjJer
ppUoI9RH6DJQevO3e79N81a2M7y6OkImD9Db2IW7D6g1kldHUJhVvItKcROjU+mC
nFmrkEKglzsWfENzzofQLGZj7pcy9xeYvvpHNwTS8h4PTphknM6WtPj8WNURi7rZ
kpYbBxNlo7CLgGEgsozkYjLbkoVT/Pf4xTiS+he0/6Q5Sw2OYIR7zdkYL9J486n0
mcA5lvfLBt/cy0MB5bHU4i0cXG0m2xQ4r4cEC9dyRYjdCGH0XS/yEBzAq6omvt6s
YL96s3g/awVUevodBQs/gmsU9dQ5Vrc04nJnsMgKy8w7tFWon7W1g0cXnjehdp2s
fBh0/pPpa4FgM8o7TE77qiyUOWoABaQEZNqef4X46r9bHk5MgPjDd8y3N9qt6Kwe
n5AwLLeey/4I64Q7SQY+TBNLviN21To9ifD8+tJwmsg2ifTUpAcXECnwrcbQ7iTi
cgFSdnjm2CfdNWOpHa6+C0jpRXAigvhyy8ADeA0vQKKWLCRz46Msn+QQ63F+cGaP
kuyHHqLzS6+WSn+TTHOEEy+ZTb8BtJQ0VDvPXO2F5hg9jxQX2YLGDa0XxgCHKI5+
1kK20IaeCUzQxcuiFprGWjLPnumxNOGlyGaz+evlmwS4T2qRWWrBguPXtlZobWmj
lqr2LsPCAIjuiwXtUzhgBcMoIbvEZIr41Yv5e9N8JVRhCSUvV7Bl6C9aPZx0bE2/
DJrm6LsugqbqN2jjJdm+MxzADE1HXF5UyIlL6WabHi09Lk6lzMn0FVGcB79zUUAd
7wQdkAL9T7ZP9B4CvoBGoi+PmsWme98YAdyY7EcXjBH/2b3BgmbzciE94ZFkdlma
A+812W85FXOSkFPbnuenoDMvHQLabdwUcgUAPE2nKBNbvHPQawq5soogz2wrlfnW
111/dUfIz0O7D3jlhkSvPz8SDSyZjkGMq8de/PfSBCBiDv8hmEZkwFm0AoJk0GwE
yiQ0jm3043X6EkcfbzCgvbAOnH53MGPHnVb4mAHbYTXo8l2f7sNN052lfbW3vAyX
Xk9bEPfJLwf287IRKl4RI1lgXHgvPhATM7vpNt4tyayyiGVwdVdzzXlrIE/Tr/lk
h04zVDXr0tLr9S16wP88MwUGf8m77BFLcWpjWDsIvbGdb4zrqtRkGq8GivUjY66N
DEQIJ/tU72Os9V9sjkU9WLfm0Irltgm358bzbB+Ua4/4fiFKgSiq7DEm3YhFl24Y
RnykLbaM/l0XSoNhJG3P2t31iuOG8sn7hKJmJew4YFhuZusAaGcuKeozT2dhahPF
ii1ALfyV4dFB9A+m3d0WRUxJ3te338odiiIXRXU13xvT6sy+rcieUAYEmwFyo2xj
x87tPXyNzCBd8NoT4IeONXanTZ/l8ZdyEWu9qzIQICK1u4gpXwkGHfGQMMvYV5nw
eoBgtvkybuweBmwIUu32VfpR9FB7TBMtR7+dSXAfMK8aBfoTfwpr0vKA95bCY73g
+ZRl604yoRtUSdEB6xrvBQZRs2rq+o7u5lb6sNTEFolonWcRgvq7JlKzFHLcl78u
CPrifhlP++89Ku3XQgamsq3Qjr3mC3Hke0rxOyOrbWsXZnlgy22+KNLl3ijLXFlr
gu40yKKFp85dGhdN+t0oKvS3Si6Fh8BMlRlETFmtO+VLzTeWaYQV3US8VcjgjJY+
OtgfQoynbxnU/k0+DFgSTp8IRDmIsTPtoSUobEskYFcw8GRZLJOvAQOewOjDmOnS
EU3n/UQor04IIgoKctjuPZumjzw8naPny8Dm1TAOSDVd8yeX4OcRJumE1ycxj8tE
Xoe2iaRaw5QCmyuaqd3zBqqybFYoPE1ykU3WvbZxb8bKhoLNFQL+QP0KZYLxhJyA
k8DoKWOqBIMygakIhy4BuxJSXyXjORQ4LXZN1eFYXNrZGRVlrBGGOt0VJ1zJi2kr
oYbTdVDJI4UBcDp4t0L166cL3hr1KxXVJPrDhasWwDqj49/Xr1KWMUJmJcFv0MXV
5fhjOgEIwXraL0VABzZFWFKW+ZpXcwBUqT+RawxGzO2yF8OqX8Sc7O7uWbuyltSA
boeDuRLKkMU4dipmu/MMzAQLPmEOiUruYg5RB9MWO5tcEZWpSNXCaWwU1hAjgDYE
S9OwBqmvLmTHL5qYcznWK/1sYjN51f1hR3X2xruCgX7xStZpDdtmBzGwOPyMRFVc
yy2DkaWZp1ybY47YRh+U5nJwdaQkLxUcJmELsl7MKk4iWvGNSkhn/oLwkc3YpaQB
1ct8MfnDWEvXysGb7piw4MRxS6AfTfX+noPinrSdcfb+k2BTvAwyh5CYf/T9wTxK
q9mCJzhUPJnhPD1nHY1dF4QgpgwK7vUL4cjLe3qhyjlEsUPKExjf5IyjScTFMuMr
G/7z4pW53mRZlu96mJnDyUg1n/CEQ6CYBD2NbIsltnI0JmzGkMx6YHIZTOaGBIsJ
ieN9AFoBqErDofUT2KJGMOPWIiEJHbOk+v/qwZTO3UrGxUH+SjBrJLDAGiILkmDi
Qx8gBXz5UkTWwl/5EFdZyaDznsKl0CTkcMy1vdG/BTbb+GqOT2VkeLgRTpu5XMqY
v+A25POFn2h5Ub2eEzIs42IkG51z5lSPU3tvTmy/IZesB3SAhWHJH6c072GtKxHW
UXQZHj/inmn/ZKDWGkKaugdWKmbxvrPanyvAiM5KytrhQ813acLmaTScFIqzkSZ2
GGBIM1MazRWY63VwzviQoIN//OSk/oKziwCZ9Hyp7ud9ZwgbYTyBORESgXGVj7a4
P10emqjBqhZQwDdXujJT18yALGljHM6RndAHXxVNtznTVg1YIMsbAa2V7983fo1g
ZS5rNw9p2bU64wOua06K76paPNr3638eoXe8s5VAio40L24wC1A7fZDw5RD+q/5s
cy3m0gQSxvUFLaf7miupROKANcc736RSpX3kxaSy9O9o2UKfSK4SOlFDFX7PSvCO
/hKHvQxxEgy3qp+OpEBkSbuTEepPM09Vvmj6S3zW1ROh2hignA6iUlBmaFj/x6sq
k42aV+3ELh8Iv0yRzvBIwnUx600A1QOMRFwPrdJoCdiewCh0jyDtjGUR6/IAAR36
gE0zQ5gh+FZ9HU5Xdx6lfDEPvA3lgEcltesURf2bh28zHJRpLqFD0ulZ9qR8jNVa
Zrs/VBXMql9EzcIiaqr+Qfy71xqaIhOiq8/tobPhjKMGr/aN0eoF4ecHbJefTzeL
kTro+fdoikrB5Br+b2JOyySBMNUUAxcmBpEq34ucjysqEqGBMfvjoJoq39OxT5r7
1h+x3y3rjIHxPNtL+y8Jg5GYdtUxirV5MJJIXaPd/QGBSvULW+JF/GKrxA0Djffp
VLciq3unetN48/fEFI6jOjshy/Yls4ipmHyGoqJhJo1s5LfutJRGoOP+6sfUBvY2
Gfp0FbL6j3bc0DB5UOlW6lLf5Dy0CyeEsmRmu0+tE2/cNM4IzkdU7ltAQy/Myiye
d6D4xYe/SSCNXuQSd5q6kG3C2NELEgLW5sm+oXSku6QxfZQkh1vFhB1isrdx1nN1
+NPSJ4IPizgQKHDnp070ZU9YnWWq+aCDkFfk0m7pYX9s9X5YnWHZ20HIbiWaScKH
gDA1Xmj/LCESlb8/4EPUNZ/AR4Uyy+03UBDNNMBqF+cEza9ahkwZKwnuqG481Gwo
5AbFIuILBK0gz0EDXxH0ojrmyENk4ZWaQV4eTRTbxf/97oqnWARxbFnjlUgJxfV3
qekBuSekvH/GZC6SpN+EWbkl/1QVeNsK2qbIO9PMMh2x1CokC5iwqJ4KvKaFmaUJ
DSp+9981FVDcMsAQq/QV0p6fsSdhlHfeUfCjrHpQ8JYF/HwQuf5cUKfsELT3S+oz
rKlCOvX99/Hq+6e0nJOJi2l7f00c+zUzQWRp+E0nsx5gVGvSLnAmhEiD1iD/LOHD
AZY9Vy1WgHqZaFRtvRc7m4Qn+jZxBKt8ZCBzn6lbQI2ZGMuZQ86ikINYTH/BRjGo
COCzrJ5kNwbkArhQNPBvUxu5UQKdim7dY/Mc5SeuWybhytF5KfFsPlscFy32OBPp
1IUY4hHxJZqAV3H/Ip6Ymc76r+BrwSYEte2MzORLOZsyqFIX9j6+iqnTvjF88f6z
mOPzsEl2ZcuuUPLN2tJHQ+qpsRaWWes61LoYeGgE5qTVKBv05nCibuULHmJSzbb6
EOfnVVOCqQZt7KorJ4bsaYbkk4/Me6QZiI9xal8ohKFf2Bs2Iz/SSKY+SY2L0Zyi
JtZhHV2Z7Dzyi66VqKd+JuQXGUuQbuAjeJOUWx6AmPd498HsxhZaKQdP+phk3xXr
cYp9lekp5FunASuP4uxtQAtbMn9u/tJwH5YSQw6sG4qqSsUHyU1nDHFQTHo2GQb2
DpfDCOvQbC24aQh0ydRqYwvD6Ct+GDCpOmcUuTIHYyI+ioD/Deog7V4b5SoPfOBB
xlxM4KWn+G9w1bYUaeVPEK/OZu6wL97sQj3cbQaVs7DqCvSzrD0upsZwRIxtUgrX
ZnyK/wKM1/XX3SQLIKk7JKl7b0OqG0GYwgEPyJKc0SNqHhCzr8mZEz+Ewiyy8yT8
9bBbyW63cE0nIWQlPYHW6O/LXHxjtCK92LfaJzzeoFkD6usvTrpkaclzs0SSH8eX
oRLPiS+k5IU/xVTroHkIDsmfmIXm8dYVEp+J+oxkLhxYeoLXzVVw6LytiCaKo/Qx
LLaddQnHaTr6Igdm3T4Qzj7I14Za1GTjrQLAaz2zpfewjx76PfU/9fpU6Ei1HfgS
/iDIBXJ+qxiNJi+2rt4KIzlQ1QXWm5dCa2irz47PhpjGM3eGscHfVuUlqfDdvOCc
2INX+vr0IL3r01ztQQVdrvpjvIjtAGdDwzoWxKPPaDiffnCI30tV7jIDLL3Ri8B0
iXOIvLOEGbDiA21gutXgWGXBL/HGNk3k0Pfpi01XIzmauNlBLM/u8X2HRzGzoVys
5S0wNgmyIdSPiaFys+KTJpRXzz/mC38BkF/UF7PRRMoOzGCi6LIWRjMzBHBezN8C
UW5vySlbO/3YgP6vCfL6yKd2sZx9ZIuJSXXOq3tNR+NzKjPua8JI12YsyT1Tqiyq
+c1kKwABFErypwIl0rA2MpFZjmo28iFhCLuc3iwrcWZv3aHeSv6LxS8tVrIdj1jE
bQsYnWZLLcdcD0u9KsS3j1+oYlQfEaqyx1CCWWWmQI6cNO7aEfP/Pcq4Xxgq0CUB
reeHRnsuEkDyLyxPi4uXgqhVH9KxoKWOJoLwxW85fQo6/v3rL1LcPZIXEptcjdzc
mpr11LzuyJgWzeLPjRxRsE/a1b+NFwF3ybIq1UoY3LbJaVSKUeJ7Pmum5ETHjShM
50nUDOePanW/HtGJFp4gIrKUwBAZ6SUjnHNxW3lH1kBOfXl4c26dydeh5P93AITw
6O04budPEDeDWDuxL7o3JIs8cRNVgNfpEl1kYE0ri4etr+d6P2B6tJIkJnZ9ljdc
uveQ5FH817WKE6f37dM3yHHnnn4xbPge3pNRzLhSxEE/EnUL01BVl+LNf5PrKRfB
LJY7wVVMOWwo5wbqTzFMlO9lLb8rI9rjTEpOciSI3xHuCOhy7NBACca3e5zePEJ8
QyVBK5iZ45rTy/kUu8iVGK5ECb07gtrsGo7UjCLgTaJoEjLdQxK4LVdDo5folEFn
MaT6v4w3g6Kr7NOBSfxGeg2PwybJlIoisJV6rvxfFeBwqyGcylPNAd6Yc96u4Pb0
Wug2lg9lB1JwFmuNSwXVrkN0oxlBoo1BBnbhvZQug0i+qiBUYEqCGipM6J9XaiYw
Tem4+RFMUOtIg9HVCkwikP9Tj8fpOxyVIa5dP60wi3RMytnZ6Et0/VLQ43EBe5Rq
aG2is3UL7NJB0KtVuumcH7hCc2e/4OFAfFzPZS1mBxLlNhb6kYrhl7PQmeczMO1R
5tp6LlASfEX3E9HfswbOOuFIZ1WgpHhON2LoLc7KIr/JMmlTSvyMmOKsQjwd7Lnn
6qg8spOKODhwluABbFePU9kmQlbk/ko40KX7uJwBs+cDZyb0G/4gZDDehY6BD0rG
mCo6fPd9xsE7KoLjT+k4qOu1Ug2wDxjGDD+2MLWd5UcCZTXN9QmccHJx7DBYSI8h
cp7EKT/TZDYGJkFmJHyNMVQaiuK0cKhGODT3TLDaL8khrCA/6S+naRvVevFa/+Yo
Tx0CnEzAT7rmhsbkVAjTBiBJEBStpZeyyx7QdxmuOVI/g577lLjPYz8Q6B9iWKXB
Ob0i5CVOP8CUfdN4cLWrELBlsgFqboHAhO4lb9nT1c65e0V1u4S8L1kZhW2Djq0t
jz/CA9aP8fogXx7BCcwlwBJV89uLfqz/Pyr9HLdV+/F+1AT5U+U9Slb7QvjqgCXN
YFlhlI3gxYBNVZBCmNGn89qqRLmNs4P7mb/PsCCAhrepDeZtxHJol55r2hTZe0Yz
S1jSJynQm8NgS/XI8NQ3q+ZTN9dcHmNNyRj+sCS7UXd53JIC0iDzZSVaKoxEX+G6
49Sfq3I0Edxjer/en+3husLV8hV/Rrqu+4jaJ6BZXv0qy7FmavDQkJBu+QKvd1kK
PHDmGNWRQVGPNwVOVRiCWZJaDoCAthhtWlZcgSCSfmclcDcf/Vdr6AquFjkO3Rub
sfl4lHJY15wG5270pGkNzQcF3DnBxUSL59/Yglp7Nco4p6mg/+Q4ZqbQTM5zgazD
oqMnEkdWZN0lYrOzlIp/4hF8rVEchKeH4Xdo/GFh9f52kQSWDFGPnH1vpHAzUkDK
1y3PSTM6rOqGLh89/zY/jPBDJtHEgW0hZtc22sSNGpREwamR+G1GUumkQGVQotob
CUrcGDL8XC809+HJUQnH1kyfkWVuROedD6CRN8pQD/sI9hmoowFHEguFPErP9gYp
hLS+JJWz1hs4nYBpajTjMgY/UApJoX88xcL6syyRUiBAlwwnu7mkokg5nJUcBCF7
KB+0/45PwVCsQ7aQO4Xcof36Lnbx7K9QJVsWDQouAyKZHJaFUhvlrNlB9slgoDJl
KqPAHZTtiH4XDOqLQfqnfzkavc5ENgVtifIsBkIAzO/0sq31D6KxdxRmJ2CIEjy/
bzIjoCEAqcotgU+14o5CKtD33xbEyeTzVgHAs7VAZvCns78DgNmQJfTRWo8vBzX9
THXksjG++WCy/hwSAvfgt0er+TB5mV3NlcSoNmZHtf/VEWKTUupHUcp+v0mpSVwE
jKnVQhtKG7c03p6QT45uTshwJr0RNlAAcJR09HUgIHpdFVWlpHN8DdcKskcY3XLb
PdyjQnbkQ6Q0zjXtPqBoWmZ1UsXXXGB/Pl9/yusz0jfTauKv6Xze6XW/6NogksU5
UPQ9ShXS/tYcCsz1DbvLaqPPW7F/7eTFkxOZcAaZbJrNQiiVEK3KhhkflaSOv4dM
uR50m+ZOwPRaAt/70kVkXw79OhCGvpnPbhZZqZU6/LJ4y38ta/CgJB/nMb/ernx1
D4dBpO+zyvAbOBoUsg06866gH9diE3m27fBqVOgLrZe+bDtNJrjheNWZYSb6d7av
S9DerzJdJ3bJJC/quMYeo+B7NS1ruD44rHAn3Y8N2CxcevhGLEWtX5IKI1jINIUq
Z2bXwKQ4YFQvXchSWRbUycshgwYjfYmRlbsPOIEldYp+HHRsW+CKTHQm6pEfIscQ
A+WCIGOOxfyM+wP6f8hgbLQ7VFcGV8D273o6eD1pFskZVoWKGOAgVOrGvvqFdLCG
c3f8sa38/dmyIRHKXPCU3QZyETJpepM5RemyE6p7O9jFjLk7paNJdaBYxejFIm1V
XRAIUBrYPKUS56H/Ccf3xo1ru0nzz5gufeWBQ6vpyJVWiLvMEaIpJ0adsu/IvY15
740DTW48dugPiv1p9xZxtYdkthM7SxXcygbztQKHVA6ErWosoEocc134WXT/iybT
NaTfZszq+M9cBU72lP9xaAig9uaiKcdS0aIM2y1fyvcdEwPPdvZid6SBbe72ErGb
1yqmTnJIMyNEM904LT7xWwhfaVNNUQ/5LljEW8usyPafFC/a7TcCbDE7+VovWwE4
QbrjatMNWREg0dVvYKefkg/wp8vBWFeK3cn7wh6nACMY1KYCFrTnJdwPDMTFNFhE
kAzd5fIev+yekIngdq0melH4sys0L6urPbVFmBtIrf80M22AZnhMHZq0wwAwh9+u
yXApWQlq4h981OMyGMjG00cY8zy0ysOqb47fzq3zC1/XQjjXNlRrGd4u6MQCbtLn
xVkN+hSGvyXKYLiULHBA9yFw67iJEFnkS8dSUIa0/0lgs5ZZN+9nQgc1/hTiyXNE
OxSgj7F0VFBqnKEi1U9hfm1zRnYvYkiVGy62Udg+xfg0Ud6MYzWo2FZnYJi/CHyi
EUg+1DHnIrHzuQmJzt0JXBVfRaRNLIcgnybm/6iDOGD6UX7ptOd7CMnFYjBF9zxY
tTrx5aRMZnX4v3er9igUWH1lT3PWYL44PPyzwiB03p/nz7I/pZPrX3dBFDr7MuOl
ZicHpdwbdL+l3oj44avQ2osqw2xCGp16mEMMEmJfjyH+sGagDWFn9sN/FCF4YTD5
vdGUpEBU8wKdydiskZSU+9ZsFmAqWSzFaBXB67EF4hnl0IQJcAN6ua7RRYVXZITX
dX676/vU9WDtHj34bKhX10XhKgj4fYG4xS0VEXItwzmcygXU/BZSR9YkchcHvLHK
QWl4JREZtA/tZFiBlNSYLKzrHi50GiOecG8FL1JuFPu9QSpBTns2ZKQdsC4qXE0Z
nWKJ18eqFpastrtVj3HAdUL9Dy/ZVkdqEruDKQkcfRRpsSm6FHi48ksaRsXCl8Tn
nj+8mS43ldbZk5tyoX1lqw3yos/MnSHOmVZn4fuNSoI4oqKM+65wESNXbt9Baa/4
hwP21tfr36KuohbtWBvcVrjR35BMPGKQLEiJNOKFzJRpeMxmprjI1tSGHHrJjDow
v6MzzRlE4ggpHBDo350kCC5ivtPiqUm+p5KfuqsOLjT5n5mnQGkNFJMc+h5wg6RH
KGDh71sDW9pwUIoMd2iE0DQ/gK7Z+P5uN+DkTMjdXjHalc9/lT5m2p4HCElS9Owg
+mzosk0ZNaajJ8KETDg5RBlCaTP2zUWtibKbyg+lg19H3gdJuIX+UMZrNLDcN0RB
hmgEUTVLhDdfqQVh0UzWc2uHgtr6nQ72v94bvOUgbc04eUbOOVs0Y75Vr5/1GN6L
6pU5Uc8yO6dGjR2d03NsFllgAznKBPvleDaqmombJOUM9MFhOW6r0zrKaE4odi+C
83qPrBoqFopauDCx1k18WpdcUIS7txF6fK0/adR39uxCG5ZbQMceXH8oNOdA8b+t
0SC79ZWvPps3ZQ82bgp1GRMai6aO1k8yd+De3WAYmNrFpOgvU1mmvnwF6BQgQKk/
YNNvhBve9cq3DbNOV9FsSDDleR9tokQo8iyeN/zTWE1+kl0+Z1hfTxoPzU65oMKt
AjMCOdCuD0XTjcY+/CRnIT0YPoDqLLdJfC0JL1Pz6H7BoDZDn79xzyyHJujaSdob
SzCyC+O2LcT+vX1ekhkR43h68LS3HZaYe9dEr1R3uJTPVxMJGT1doms8yA1r1+Jl
DA1QpZTXUd31rdJInc2i8kXKF7eN47w/JwMLguWG1+n/6yE03eeviX2fWGEN0zTp
svMz9ivrLOPioiknOBAIXp3jpS/JTxdVi50dEGMXk1kW4WvfHM7v4n2D5td0Qkbn
7A0gIlVEZYROlvscTvwAU/8XFxWmXbvEv5B2Ot2qRPZ3D0aGZa0XuP3dwO1/0e52
C/XAoT4BA044Lt0D7vCWli2wFvs2KQT63THyRISfCdPc0LspUepVMBVh/d5qSWTw
vw37DjsAOM9/Nd6+E8nxuGHGJRhSXONvO9TY14kjXHHlR57ATqE+SexcejjyNE7x
KzAsyOBMOmI/ndjJ0lWvtp22ITB6OfjGxKDDLfKVaD16YBtuMMhgV8X6S4RmJ6+q
BSfXVhtdciPPccLmAfvqhFtCxWkdDokbE5RDlqkBicsVjVom4CY4Etr9ZE9VM+ci
TgosjGimblUfW3WjcUtXsel0psrhFs3ofWQWLcQAKx+7zCoSfyI0kvlmBh6NRY7/
1iHmgU0YjJ+8737u/1Q4y6/NG4a1AP6DjZaOfOJ2uoLJl8NFdLeZ9HYlI7OL0j2u
y+gB8/F6KBKU4wpeSWQIG20PB4LFNuk42UO9xRX/VrNyPSrPxpNrHNjECs8EizpY
jwWLK6BSSwAaqPhVXRqKylvO5gR2IzsUKksWwfw7WjZdAhlj6DAtvESFJgBfwWME
ZVN1W76YeMuAa6e/5pa/K5tBKhrm6WDvvMNhol151m6Syf+mcukO1bdrBDJNVK8N
/auR5P79bigRqIY8qoelPtUod7aKKidOimMsTMR8FLlEDWVqOrstHPL/GvU4M0sB
EwB5F81xjy6ngzMEPt6UN2ROURDlZnmMFoEmPjHFuKz8A3H6LtBxgYAMiND6ktro
7YfgdG/xZtlbjdtyQrbGmUQE+7OgOoICoerpaVCtjWh02dhq/nI+O0vc1ukyfNog
6jIA/21XXzkswlr+C7QGNM10UHyXXNP+cHTKOILzTTxA+X05TGC31qRhluofpEHS
cLFEeO6xZUexenmZaAtk0Q2QjnaItZiWwnpnUD8lj21bXRxbH+tZBeLmifihg1je
bSkxLrd8i8HzceSxiV/rpvh0vJ10fmZq4DU/uxGKGSv/obpUN06hse46j6RLU+W7
Y8ZXF+ZxIG7LI+MoNphoGdTDjN8mbc6lw73yVdY7fGdjUnq3gGS8QqwODy3e7m2f
J1pCjQ63sw152tbo52K+yw15s8olaW+IGrPxrj+WoNogGJJ519QRKUc4yombVM1o
B83Ruwn8ibiCkNczIxLnGTly+IcLpY8Og38V4ZNXMokNvm3nqgS8qZdFNj2CxX6A
84YQJlY9H0+5SZvv4zVEfcTN1gM6RUTzB5cMOfpN+JMI8OZIPHu7qXjISsSGMNDY
rqy3U8Z33q65g8Sjol6ZINQ9XqivUd6g89li4FhUI6fsqrEci7bOlfzXi7A2h/Mj
/UX94M3mfkFdhS6kBORe74dXayPsqhUE31j9tWvl6ltkFKRWAc7GTOL5Okx4R2db
3tKkgmcUHwm0zw/Bi1WD10uaKoIzl+toGswMPguqu7UvdrR7J8+zUxoW8VvhT2pB
JLrZJGPHTYR6/Utr7IEMv1N8dgwUuOhKnh5CQ66E294GSuT94w2xzlTH01kJQwlE
ASsbJMqEAL0zWXj97LMoJLo3uiH34PngK+LNAdsYAf8kcGLf6Z5HH/HIaCsVqe6E
40kKEwcmP5+KHePRZWrjp3WGapS1dGc3ztZ/3nTsJfMdZnyKuebhmLFV6z6S1BN9
R3nLuSsaaDhI4wmLMCmMkivLAcbQR+4GOi6L+0so8KAGeTTFAyrBCgaxV7lCAeYH
QCis5RrenZOcDaZGT9b3l1wzvPjNkClVE57Es/BWvvqNKQPPkAzqytP8sH/a4xyT
/XS53OAJZQMukDsOySBKuB1znmRUT2ipAM8QHnEcNHFn8JM7WaL2y7QWn8638XhH
3hQ/8qFnMla1XcWthtJOTvNygd+RDPMlz8fiHh/NODQnobnEGp0noO5y/vnUg70q
AusRYifW62u3SQGlkLFSY6BQm5XmQxpIQot0errRxwAdZEg3khECl79+VEsQj3D8
u+qJu9SLffGQDHVH9X65pb6wFuKfiZ8ls8CbYZhs8YF3ldPli980BiJbal/v2go/
RkPaUDZHOwUjlPQRbpEdbOeqWLLZpbF2TYbzTfCzxfQh8zXRVgpyTk9oBDV8EPTv
Kb4qvXPj6RhEDceAvz42xLkYUr1a9cE318UjT+l+9dR3z8gDtxa8CcZem8Fkjav0
k368rBx2v7DExqmh2FP1U0QTgesT6rwOV1LBNfHP5ZtRxKL6j3iOhKyHGB3tmye7
3evq13A9JecuL5NHdPbpv1TSPu7NmXUlovlij5pXd/X5RjHzGqx7fERTToDiBk6E
OJOGk2lhpOa6H1XCOK4x30jgXemW/Umb2B9dQqufRcwjn/oZLA/gmATViy665tck
UjbV4JIGtaJhQ22V5mIa2avUDje/Kipw7wZA/i8Ce3JvbbF06hE8qKb0/K1fkoll
dezEQ0lgLXVM5juuf8mBjXtZJnmCHguetU7NvIpVaTUULidil3O5WZPxWET7ta0g
uYqeFWEq0AB1NnL+juNBvbrnhWY+t/Yz7ZEbhndabN+lrFa+Uurcn2iw33RhaUIW
xmHrHLliDVfGKecn6/lRd5nhNTRkb64klnEuaZh97WRJLhi7PWn8UdZgsfAq5JlW
OP5U7HKeMpNlmsIT5vqgMiyxuoObOwxaEs9lcUXG3lcsYAYBuoR9qSt0E9W/RzSt
WM7Z3OBmnPIHFG0MZ6+e1XOfIq6KvF9AEg0aJKj8U1tdfSJyX/VpBXF//9qCdMC7
B1LL7jhMyur/o/5cXJgijb5llrLBaKYBTznjqlFDIa81svtYHldCTYCKeyPpGEmQ
cTWrjTzjIoGhrPhvfV3k9/onX4IPxxJ9MDGHHssTgyZplNgkCdiTD01sScPdL6Xy
jgUrpWjUUaGjUx5BvTfcMDPD3ThxLyMhYza8GxG/qn5s3YJNTDknUzJBTkamx8io
CtwRBIHegdSge5GxVT/e4Ma80zcgukBHaLKVRhbHNrrfztrCKwkhn9p6ggecHSR3
TGe4ryUEd5gTlH6RNijUiSDsZSwBRLqKZWW2bQNDY3ZTZjI+cIRV/GLb3dDdZdQh
g54QrN8iY/Eceisw3pXclUJhhhDKqDTTuE5i7PHfgHO/vUw2GA5i06YReP2iAmBN
wJgWR3Z0Z2Xb2ixP+BuVZNYoAVurymjBU1wWxlSwrgjC9JPuu2T0zSRRLnWRSGjd
FScAQKQcJkj5STyg1diB8JKDORjkMq1ghEWhfaeY0gCpPP3Eb+K9jjsK281+Fm+z
8qdLjjrWztrV5tYnYIQg8v0x2EM+u+euwk9VqDl9sekkNgM8tPzTi+kITObrva3G
novM6mJ8aJyEIHy3JTjKUiJFxEVNqSTYyGiXNmNrGL3RQnD2U2/TEzdZyy8tv/Km
MrwfOU51UYWHg8XgOImGLzOpvFPtxzFSY5BIO6JvqkBckp83VhNzfShal+LS5E8E
BDA9imv/ZIqVF4tAB1szEWnKHbBQf2MEdZsfdPsB0+pPTyyBJxS+pbwCwNPpICBN
wAEGbbbusZpy0DJf1KZIPoG90Ft+uU0YQ33/VFMBlwYKkF3oIOCBBD0EAn/6wZNy
Q9wkLeY4rMSIU2r/s9z+sa7Mam1LYJHxasHdFUuex5IpGhcSNPFguwKKxCyl5ueE
UauZX0fnf28DOM/+RqzRIdxwwF3MaDy2Hdfi7JVWGx7ups8MkgU0h785j8NVWGiF
71xzr0iuHi6VFtnnf1CEfl6cGrRaSC4s4Ezx8RtBKupw94q2PeuwdwAoFje+gxhq
Qy6pGT0jdjGwfw9PQOdcFFE8Q/JXieWK/QLiU1KImfRvDA8NUkwwT8vU1rLS22VL
++K3CJ2KM28gpqiXYvv/2I423EOyYnaVBcI46WpRh0sBVPgKLrjjoxN14URmeTy6
g3RCou8hPoaJNPTuiiSVJmTEDPR3eSjBInOU93GIPr0aWCMd/89rgvuNe6I2gPrt
DTbbfcGnyKVKxCb3Diays7CDjRVjPy3hAG2VnVjFJTKadjFgCE4kzR8lbXHfL9qz
U/0MuD7N6J3swAfky0JcgZ5HXgl3uyJnNC6ne7KFzDg1mHC4QE2gveon88oWg1dx
NPoFHVIM92olnBfJrEeYNt0RGNvDIEKfQKude1nIsYpTrfapMaQgyPSWZ9kYm6mH
DCNR489PzpzfuOVp6kjTKxkBVDXYkegHyKm0mInb2hOomhfeuFWP8X8KMOkszWc2
BkKLPxaHUzYiUPmM/hZPSHHZz3Ddl4OivTgt07Llxz4yL29ht/iPz9pqEA7SUf97
dUZYS4E0OAB7YXzm13DC0Hla6B8kq27ZgxwMgzF8pjMrOTG3X+Axc3ZNdtFqU7wa
Ef8l6AT+jVaDVH8e0o+JZUe817oBJEtiJN6or8aEdagOF1cqdcxhdtBfh6L8pFaU
nfLln5HsRQa+tTJu/yVFjkrZqMWKKZLaGatc2AJwiY0BKIgnVnLBIao1fE79YPBf
AeakJZuCsi5HdkL1jUkzyCQLepuR8iNS3AlO7VWSn2Pytki8beziyUGw7JLIklhS
Q1m8myE0Xa2OeqPK5FGwu2rLaR9Lg70EgmeEqmUCIeITX9HV5VRiivFFc4OXSNif
NabjsprdAgCmrIu/JIcIQRpwRJIfWNef7HcNLjswiW0HlLQgtJuuF81DcejRQEtA
aRzj/4+xvUlfxtHC5iQEOQDRBdGHwjnzS/CrdbVLw1X47B2Bk9I7fpIHKK0Hzm4V
3mMoWH3Mzqx5Rg5L5Fes4HQaSMb5BPvD2NGZdHjm4gB2RbAYl6pLqidp0lAv0aMR
FYuPe8h7tVM87cbNWQhZ8C5Pj38Mw0otJ3gKYE771Yolb6aVaLwOSc+M+xz4Pq81
idguU444VvB0BRj/RNdluNT4F6Ir+TAUsDorrqXJ0LrOcRkIKC/36XDhRPG1HvJX
pb0S9WY29mSj0JA6izRuApPUbFBWXHAyA3E6O4n0DvhjEAZMTNRALwnAOHIlrGbk
CrNrKkisQqL4RyIh//24SfwmhlzfPPPc5raU7QwjxoFW1p91HCBpOsnPLpP7h68b
eJM4C7t2pfRkDgL4YoNXCDmw4OsU92FWfglj3e1k0ck7EnuIb8qd/ad4gndmZoHp
59maCJMS+RGxbCG4QZCn9O7vMjJ+fVSg4PKh4BUgrculQArpK8qstdvF4H6zsy7V
X545SUj0M01DLfo9ySAMyYVzNRxJKlzk6p/xqOZggW+nLhSEVl1IndkezkCTiW0b
CvYpVXYOP0kydv2ks27noXvnPZ0RXKVh3rPIYm5hbxRlHls6DrCARczIiOfl2lLS
KIszR2eUg1yi3KogI/Sba7Ym4k8RhxE/Q2xLc4vRPp6VTLxiAHnR9xpb5Bq/2pfn
WZfhy72GecAQCl4l5/jhe4Yfzy6zZ7eKCU/qtmedZ5/5bZAuX9HBAqlbVhH2wqG7
KC69M4Raj9qnPsIMH89a+TrcIuc4I8EfI7MY1fLPkQCZtZBxi0Xfg4KAk/5BJLWZ
5KfgED5l7IKfVof5drAe57j7yVH8RDGKfT7fGVd4HoxsWMru0JBCEclEgPBVaxmy
x11pFoc5ohKxYZVwj9f7qUDG08cEdOaxG6m4wIs/wg0ni7Ef+8CsSk/tPK8UmI5w
b6ACy4Z6jyABqa81Qx8ucMxVn6SkoTMgv4w6O2Cm1v8ZD5t4fhRZKWxhG/aM8THF
2P0E00YxHsidCyXHfdN8EChq1f0TjhOr8hE964qM08hSzZfJW0V+9yC+hoXPkpBC
NoUNW/qbRTFQOTfgw6UneIXbDhCj4CNmAox7iT56BBF9PU6dS2++oH+o/g6IsSn8
uAj3swGlAsRGsT2OTqqvW/1t5fs1MWXDqt69l0iszwn+CRguOdFDqqCqdSblcLZe
5cBe9K7zhfNZIClj+c+dftSELjzgvZS3JPle2ECDzIOvN+YRnqk5kIcvVcESgz7H
uvVuq4FLxOrDhiEk2TuLDujOgyHK99+U4nbI3JKTpPvn+il5T5454w/65T1VNxnC
nbE1IuZngV5t6EPsrNoR8pbtvWJvSeO0WyXDD1e8A9+RQNT1Tymqj7jnG2P53iyL
v0ASW/mlZEgR+d712igo2V3xffWp10aqCcZwT9yTjGcrf4ij58DejBESGF430F6M
G4GiBMyrHKOjjccCMUw5DBOmDyAM/i9SInhdRAIy3puvNPdvcB/5V6xlOOwuOC4a
sBbioqiZgyGQO4ASDITwygq3rPAcUHUBpJZesqxiHfZnQ+MllzcDxGKnachQNMdz
nX4MCU52PqhvFZtZzQK9wGi2WhkEsHvOegxJE6Z7o8clEm7YrRVDhrPVoDK/7hgN
8xshKeWueVVuhrxMosYu88hujqjxrVzetrgM1K2KVZX6DWCko8QHXByz37dZeIai
dHglatwlEzks5nOVP+SRWTiu1WB7dEtdhoq+prb0uq2eR+UIlZ4GrWq9/IY8AtNY
vWq13XWL22TKUPm64XfMPjId8cwZZX4aNNhdAnqkPwgGUHYAwnFodBXi40dqJvWL
NGvxFOrW41Yh53dQb2MYeYqnsAG6Z9EzqsDOypbcLxDXYkWjqMHcoliuQ9KW5C/G
HQ/DYP28kAReZdswgs2zaun6G/+sbUU/kdWD6qPufzTYtUTeqb2izqwvhP6ye26P
7HXqnV9Grcy4tyVO+Jr37Dx7waCglBGbr+s5VI4P+v7CEqGkB40u3Dw+92OF2Rml
2SUU/htPUIAJlYmUflgQnP7Tyb6qRETaBUpPclK7bpsn1tsQ27/ivgNyjf+pXOIp
BKTdgQAxnnyXRPCj40TALfn4XULNz5rllO2po9lq6lQCK8Nxq529KCiIY8X4hgRM
+NuRIaze2pNifsq6ZuLj+2RSlV1dWGE1h7Q9MplAEIucAS8M0kMUt/eXlR3atiL1
cesGp7p0zKviZQMqKZcAX0zOLFg+FFf4j3d58VMs6VrTOU7txBhFzPm4htVgDJeV
05TRlmCNZ+ouN6WW4u6Fw5in3IDdyYcWbW1Di0QUBb2gGqsu/PjRV7VX6BRR/DS7
ENl02c1zkc4lMmBN4+iI8YRht4cXeLmYVLpnZZEeGtLd6hp2oamibFMYALQRMwAY
F8oVBVWLxBJNuE+LpI3w8UaswQnNgdRH/IkBEEZ6fFh5EhP/7HxG07bPcmpYq3Tk
gyFBwKWhu3b+98Q5YmrJ1tFFX0qmqVKk9vbbLq1In//WEecNin/sGzX3pR7PyEvO
5r8ID47FYkMiNqTxiv2jBGZ+ha9n/cYYeVvsPWddmaJkPnsP/m/r6FXChfh9L+J+
R89J0dLxliI9mVHzSM0BWibH0C3zacwv8naSVpE2RQdGnJafphPTsAV0iA48uUPz
BpH6Ww+7JFb/F+7t1dh9I9kHBf1z+cIw8R0vMviKHHpfBsIRPBwMSlOiuNu+r0Q7
g2GOVNYo+F4FwS9rH/sQ0WPt9ZdHlAYOmnATU2Xd/bleAXy6cO6G+2+cOliBHXVj
7TEZqAW8D/SuximrzcToKijaHrKbUfBUjt+day2zNG3pynfnXpca17ZzI8vrQB4a
9OmlXY6UWiYyKI9rRxON1FIMPlMCKYYOIN3uGmB62EoFcW9Jm7WYyhQAB5mlOjS1
+QVkkQOLU/5dFC4GamyYKMnChArvw/KDZGLGql6RGt/xGrNZLPGpLGymSFXAbsZZ
rTjxMgFPjTUSwl4uV/t+6qrF42X2/juBY5SMA7i5AdPvrn4JMLVOu0fz4e8pY8DR
FyyFsN7N7QHgz13e9tzs6hrFG/NaQx3jzeOAN/5uCUFL8eU0uyoGUqHtxKheyXIT
oBMJmceSpboCaLnOQVkmyUvsrdHEJi99C32UPJLqIq7jLn2dZ9TuXU9RLy6YX/EJ
Xj4nrIBt3PnBF6Q0wAA/PggwVoBTmEBsc3Q/uO/chnn1QLzO9xKqma+2i2w5+uLW
GV6bB3gK/sVjnXSuc36HG9mwkZnFKIvggYlvX/qiDqZnjYt99HVHEKBEVNMj9uc3
cNKXaTp04ev72yvEFM05RY8/231t+fVYopH8COLm5gcKZNyP7mKgBwM4v+Q817WR
hMo9nE2lryXLRZiiNHMbcZQ8s9NnyiH+9C8y0feGiUGYCYr0QipKQBemCi6KaMqr
aRxTcTj0a1PBS0Hi0Wsr5qrQsaQCK6XPG5AcHsUqNCUCAgt5xTPGYXKSemHXl3be
BlI07yHoIg9iR0yNMD5vJCPzzlZ4tzJPfr+YuCR3QOUpqhFKVVMXBsdrModnqzCh
G/KnscR6o6D+UboJgcAcyVFKcoPscWLLAZazRs6uGkMcOoaVz8G1RwalK9o9QJ4O
6VwrEW3RED38B2G3uW1/DdnHmQO+vMGaUMz0PqELGX8K7lt5TdiFLKnbXfTigHvI
Kzqj8xkA36hNwikfZKys0QzURheIrY2jNKrHRus8+LyueDX1zam3vbz/X7AYfMHO
2zQsW+Bfjq8u7tCvlf/Z0oTY7Etthz4zDgHbzYKpQdfR7baAQ6r/Hni5n3zo3dB7
FYxi2y1EObJn//Ex+9oCytimZM5kgwR+v+OGLl0tMhsdI+iSovi3yrcHnYDmkOl9
bU0vD9dLYhKuNWjFshpNvkl5PwN7JQnTt5zD7gphVipz6KcgjH6dR26sVfhb6uMN
3y0hplGDqU+d36853Yo5ehWf7rDMMSlW2jb/0lPjqyvuAYYXkPxWihcc03fLx10c
uupcJuJnhkuBap9yps1d+LEiTSwgWM3B1ujvpw0Gu+zEpJjPyzySWDeuFgOWwX80
7fXzrQ7htoVmgkhuqj4jymW63WkMUSOhXz43E5kEd3JxQ1lDEfvLmUHGSOdGfj8V
H2TC2TsGPOqcaubT0OpOgXTELt28ah3thJWkIKyKB8WqoNzcRTz3z/O4DunPhPzz
mj65Jpi7N6JUSe/LCVhvXaqhlM/5PCzgdw4ZfZzZfCmTKdvqVtTFOQV44zTDaFbs
g7D+H1qp5hlZ/Ef2KLKaev+4Lq2SQwgR8h4zZ8QK92gzi6sQ8Zk5OC3DlSlAmyR+
Pf60t0Fl1r8qI3EBPVP3HKOiANH2Y9BKXT2vE6KMcMxfRPTk+2iqRYnUFMaTHL9I
/hyQ+KvW2XwvqJWg0pc8EhPFtJnl3VmB4A36FMmAUBrXaDbj3LnThPJ+uisNMvDt
8keECGX5b9hzWFU2F1f9oVnBcBQ1aWBhwOQ9ypQa7WUupEGeJTo8AXstGpSj3z0/
i0SyIQcyFip9YzuVANnn6JuGg23k8iZ45EEuiZ/z5F76Y0bUd15HpEVVIR0GnjVq
20IbAS8+jDVT/pyH8UvlJxlNimZ9Su3YV5WUoT6vdNeMQhTePaS8FT4Q3JvuB1Vt
5ZGp4vX19rJrs19fXgWgxDqrvQZHnUTR5jDS1mQVagQekfEjwGqcLyRhC7U6PyaC
yrDTLkly7sNUsQfdGVNQlq1bEznRMlTWT4yI80Wq0yNmRC4lGUTkFWk4m7S329w1
A70r4huYtwI71m5lcwjjc8bnzm3LRtvhyjoeJyJHsz+PalSjY8tmPSdIkINvSBiS
HOWtDdGlwua44y27VWjfVY6Ce3rJ2dq4ox7fCrlHbBLCR7gViLQrkFThWW7M+ZRj
ZejP6IausFvyeEYAT3XjvB57ww3IWQh73+I5VdVSvZE1w4VwBAol4c2xf9pVu1rB
peot+nEoxj0cRGMPg8SVkzhbPoqLElXIv9vZdGH3YTukF4jV1H82oF4N9RbCBubz
ehzDjSIB1UzOQrbUEmIhO2D7RrpFzUShF61s20/lYukiqdi1sAa9x836LtVBTKX6
7G8M8JqgrzdSRkxs814nEJRqiRviVSOEXn4z4yXWCbNSUIfwk+FYt3K8HEvfA9WZ
f0poDe0e7nMca1w+jltOsd4CTW7wVWZWVt3KxGUOS24yDkHbjeNBldABiKGToJ8W
Yb0clW5Z0mkwMzVAU8s/1YR5O3yPQU/BQYmXqx4vRONgV0xLzV0n+jDthljBim58
2BcbwAPQGGJi94WBM4ey0otCCr9//axQ9SAPrgpsjGMBlQsRbIhuucEYg1v0MV7D
V2w2Glks+2bbYj8+7ry2Yr9LOjtmLEVrcklcowqFK4WXlrf3O4NT3MXkQ819SOFG
ErQfxInaXWyrfidXvkCw6GiVrPTXVPGRTC719S19GzESgngBwTQAkbu4yvED0ZVK
sfYaskaR1TkR9Hj3MJjL2MSKuGFuyPcOLIBre1hZ+NdOUX5cnBEYK3XyIJZAP/hm
k4kVgyffoGWLSpyhakFvx0CWwbzBTZRrS+f+FaJJHgBsykHcgcoRX0b/lOgda6C0
VuwCg93UuRryEiQPdFVKLkNF7BMUsQUPtHXTZCVtyU91OZUvrZRODnXI6Mdqz+eS
WUUSEVz0KY5wySbHmL4gkdf9J1LeayJm27Jl5aRnTSYF22TkgEE0+zd+oGgv4wSi
5gbHw0uy4gy30xJmyM8JGnFZNng6ckDJMkVLeQGYRAZ69CjI0xwgrtjpQHv6kq/W
4ConIdvlqh+NukFM3JULzQ52oF/GPC72rkc4bLBoQRfVz04pxm+YmbtHZrgsbqba
8T+Bf67abE6wmtZDqTcUvmW64m/6jtNvyXi9KqL2I+JHavARHb8tLADAY3chgiEE
DcbCZjuB0eq+nilfBWOEHTqXT2YB0uOTNzMRmIQmYuQ4vSIsC/NyAwKgievNpBeE
Uqh45LqQZ/94pVPCrtE6NzX9sZg0njxya4y6MTQ7CbppBFlylapPZ/AZk6ROD1eX
XP6dy6EHwDOPeORnmkdA7W0ZyGyJ+akytcbfoL1GDKuH4OtJsqkcd8PRFGMHtMXv
f4K1elj5aPX8SRBwNH/7kkvlvLYoWS6kHPYKe/ZZVC63+loSIxbkfnYjht9Zq5qc
3pMpK67fm+/AymfZ1lAQGYZYI5YPGyVEWwC6QWkVqDtasrCToM0W/Ub+s+Dg4FVn
g9OeA3iVDb5LMlBWAHRLCv7aYI/Au8Q085/6eiqta5d+AiMFyVrP3+wQjFh6eOo0
+nxCYnP3yEenuEwlOrKzSX55W6dqzcXfdH99iMfbtiq3oRmugZS2vzZ4h61I/K0I
VMgniQQ0I1QyODjAXjVhjeOcl/5ewcQcxgOvyBVM7eL9PVh1cfqISS9OsXIzqvat
HLw2K3aXX5mxhWEYNY8+wtPGcI9qlkkO/W0+Ei7/UWjgxXoQlJJ2jJeNM4CGqjW3
lWL4TQ+0Reirm9C5yEhS2VaEkMz9IsO+n7iVeRgc7cttsj7snJrls3FTVX9/+Op1
B8Cvm/szVbK3FyKxnD+FV+Ff3Akwyni7XtW+N28ND3ePIBq80vK3HFTR12MufbRI
whl8zasxvCuvmneG8qczC/K3swp1WNBK0T1Czlmsl5e3WRLUBFg8ZNL7//ssqM6P
C+vltmf5OYqZskvly8+lsvFL7sNOWWpqtUrysuhriZKs+72NX6CCoerMYA1oF2Bc
umqKx4npwdAKX1JeV37i+wYY6JwATP24gqUp1sHnYu2g4kUvgsts1qEAo4++1CCR
cWVpMFK4hB1t6KwUlRZWxOMr9m7X4ZOH/IpkIbk8MyEKoLDiGw4vyb3cz5Isbwon
NZrxo7pz43O/56iFNsOR/sIrCrmCeyirkFIVL0G0lKG3ther9S8beyLfjyiMb830
bV5mRfoQSX6tWutL/3w222KYPifdB1RHImvQePTcgAsTLCVKdS99Us/z6493S2r3
qlPCrvlli1BzNSsUdf8bvsD27CxSpQmJkh+DMidp3j/bQcrEeQHqRzDQsGg0EJGs
r7zuEogMrEmPZqeDQPwliGz7rgQ2aADcs1bfHb92ktD1WfbeVsJbAzONE1AuEGmZ
hi7T6F4t4ccUhpsmJBnPWF8lRjIq1+D8skjvvFJIeI0k7XofvVBddI476ZdwmaqP
BMqzAhn+1BpZQlDUOGJlNp2LgP4XEnnZT7R2HSuVR7uQguVa/5/cWAswIiezyefQ
OlG3zDw8UR6PGW0yLo+VaMyrLfOr9xsTBJY5q55YA/+QtyYaZi9vXLsbRdM9uwGi
SQHpFIIinlzLkr/HZFfZ6Vn8GRrRrp83T52FyKJ4JasXMaRqVhqqMT5eails9KYA
/LtjF4fEk7x8lhh8gDNprXduCj+lDSAUAXZczWYFD/nzFIV+W6NIY+E+XlWpezk/
PEeRYkUfqWQhNvLCFO4LkiefADAADYrzpgPQoJcUKejHx/ZFAT60sHsSvimRx1yg
kBzAOS1UaoqhdV+XtkdN0MEUZYTggQVE6cvpaq4jsN6VLxxU/dA9hNhYfGerJA63
Iye1A2JrqadCE557IQg9P8SjPhz0utHYd7ho0+wqVlOohGpWzWwpSoj1uitIcI2p
g94ameFoIANFyHG22r4sGDl6cbgUl7aMGUeAonooF3tbAPYjUmPbaIi3hdmlq+nM
MQbtqWOq3X4+XIPmhfODoJuMqXrUKd6bOUquMq2hTwqxk/vQT8YS5UMgBq4Vr3aO
khKhIN6JAxtxtR5avZSTTEcz1Ri/PiaXeEgM1H5+SqJIQhOuemQLA98vnlrcYpHL
27s34lvxufjzCLJHlA2oy3MMOGArlLH/wvQQ+389krSS832kzgkv18hM5ORMUdZo
s1nEP3YnDMt7SRG1Qzd/0YcD4/8+Rw4Gl5926Qsi+VjHt7Fo//XPD6ZCB20zJKa1
ZLCyn38y93uP79MGpwhEL/L/ipqoI/o117x2l8ejbwANeS2hMRNq82+DmtFhn854
geHqaAWKr++4mFGdAXFepLs6Wt5rprJMXv2vNUPdQFPNHql/OjPnnFuAVzX4UcvB
8wvl4nGXojeeO6dIsYx2tCksq8Eh03gciDx50q3UjEOjnVSY2rE753tC5pqnPeg6
k/sMDPe31Sk1zpc7Sl/Zr9QiRUphmxh88hO9hsXEKW4dlTP3GQzV44Coxdlw5nbf
1J0B1sw6bYkQAmkhDkfgbHx6WFQlD5njiGPS3rP3+Fx0TWA4hOVjpnF0qoIOGTaR
mYBHpDyUcmIkg4nAnrZCAlKj2Lm7XvU/657i51pHos0Jj4l50tQYj7131810kMtA
p0nEjU6IZS4RDuHT1HZOy1nrhZeEgdnKVzUF5awUBD3MgAye+7TtlbFLA2GrrddR
BMlwvl+ZoWcT20vQ4sV9kr7IeNOyud3Axorc3gpnxJ5Dhx63DBax5t/VvugKMHJH
nP0s0Cqvxpb6QaYZODH9l0hvVcgRu1ufGsGBJEBgo/J3VBktXWG5OJkZcJkeW8Bu
H2Hu/AsvYhFPEe6q7/ttL4cIzJnMiTPkPoRRlKl+tlizFhhr4FgSqp/pPe6K+9Lh
kjlusHMi1nqt15VhMXlMISp4wgM4ZrZvI/Hg9u0LBI622hBylXraoK1sSCqtZiYx
LNK4T1lhUU6EYJ2IsF21u1B77l3eYVf8Oyw3/C4Hu6JPiMsf3BbAFAnAF9dfPhOI
t4Otev3oX4RD5w+igDlUoNi4B2krNTtQDBnvZ3S/PkAG10VVyGhU4F2bO3s8yAWn
6QacMzHqIZGPBUcTxfjTmcVn3U/ksZGbmZX0wkh9UX55Kt9CceSPdtMcmuG8/gmR
MBNSLQ3PH9EZ6cVi9H5iDXVceoe5ZInRaXuiRDuHTzBo46N7ohxPK8zu2ovHsJd8
yuY2mkLS5quzrcJkRi14dWcz6J+OWMaoU3Xu2YU5l0OQtav0OkH+WwtFGE+EvF9B
iFXUwYd2v/dvb4pzL9wUMsCRtMTTqVLVRV93z4cvP5xCs2GzR+LDUR2Ma2OfsSip
c1C/ZQp/4G2zJg3NtRIF5pL5dhw/ANFx1dD/nKyzRrE8kFvAPHC0UJzJL6exN0mb
mXe1W/o96fWQ4gXBTRt2rJlqubp1z82YLovHeqL33muvBUPGXLYrlub+5Scjm9r9
hnrhmNrolBjeLF1uMJ0vdkUrWXjhE+3zJI1qxmUlBcC1o4xTcyi1G7+mrfDST5LV
qPY6/oQyPboBaMUkwVxWrHo0PpvbtNSmjIFQ6f3FG0CzAJCfZ0rwfiZqtKpNXxSM
q6wZlN9MQ4GvnGN3ETg26hcX+Eak7X2qm4iXw0wPsgPx7EhmgYHR6T63bfHlktyn
31kVXihb2jRXTXxHGhbcvLKhDL65+CWzKfJbcKJFjruV8nH9kYDIfAv4bAFA3hcd
wnRDOA6scIChuuO3UD/p232jXYBry2a/9aMRKHw36+9ZdfG6YtodBQ74pKFcFUiC
Gq9bpA3xxMPB2KMW64SXiXhJKrrb1akHqvnIWZAQV5VG9UQLrmB812fNV2fmxt2M
MusVKQEwVy1eSD/bFHzxYIn9JsG/BLn5lfU7a4aJFbLTKzwWAA5Jz9NSFyKAl3l3
4FCRvQ1knfE+oQYxJxu6Kgltn4DA6snkJqgBrCnk44t8aFQ6sYrtA4NCQy7Q0aSC
R1Pvw8yZmpONpApJ6l5c3vq2YOckeBV9/3/Lr0sA6plBEDu+TMHTNSjN8IwqnAqA
eyQlU32T8d+jtEuvesEn25R0N760hGX5GK7AVxNPBjAguBRcAFDaMNPWT9lluu0E
in7dMxd5Zd2C8TEJfTLq0HoMV1ybL3MEknm+aZ3Aa3jCm2/J6avhU2OIggyrC89k
Bv8lOAgfCv0V6UVUZD+Po3MrJE9QmwG26VfFoUf4nJKvCgTpBJO0o2RmQjQ3cgK2
SZ74hwM00jidBsJs0A6k4xPAndZJL1mcKTmu7YrFTwCMhBHGS0g8ArPgtTxPpBSf
6sCZ2cjpxTnuvJcOXtfKBWzfEuXgOIumTbITBYPOiKJM3GJZuT3ByRhNpcCdS1rw
APbW9Ln5p7AcvfDqUIOAuyQI2MQZuMp+Ypxvi8cYGNL5Iidzxxc7cQEwZItvZsLa
2v54zrTKuUGw+uMQMDRD80oiuasWhLFUaA3IC861Ffds9fB7nR85q3yqwnXMc67T
A15CQ/vSmPuDNGWWm+SO5I1vQ7x37QzIh8w95oaiLhx9VI3rAw3Vk58s7foujWv8
Lo2aGKkPvyx5U7J0YeSy6rjN+8M2HClaN+L26mrh+CQlbEXpR5OywHgMffDIiUFR
yMfCekEzuTraHoliNkkuH3Qip4rMnn+k7WaRh7BN9eSmFb8Y7gOP06cHuVqqC45/
matb8PKnT17cboEkFezV3wm2kNbK4bX7YN9PAHMgodMfqtnKPQqPS62oTIklX0PQ
bEmCoJ3dR28dXyJgZGmB1XALy/yPSiuVcNxy6hSpFYCe9rD+GjGIelPvaR88iCaS
pYkutCvShRzt3JTaLRBw9iClpZTwBuDEquNzjbe5AP488qAmVQbcY8vR5cEE1xO9
2jIkZKNOPVvqhJGGKP1hPrHegvMjXr1IePDLtILlwlwvVX67Y/xq/mCEihQVCgVy
pSL/n2BNrm7L81NrHw8fUnqrPb7CgCn3377kMYqyo4Ra0LnNioav9kwY8whUZOGA
jOaX1SFqE02DD/VAw4jaxBZ6PquuDCqH59F6ZVnhEjvqhUfcbhU5M8yuLJE30kSY
ptwYkg8PH1Oq4R2s3XSL5ihgmY/9p0+m7LFRZC0CpU8DCnf3gAPvQrzK3NWhVMru
h5QIkTUSPzl2l3mSRiigBZJLPzeMfz3iCit9gWVqspUfn1+jgdrvefMkhFwS9j4I
wY2FRrBCM1AJK4Z6YVSrVWMM5fzXlhEhGY3VHdAL/TZ1TxQXxaw/Ja4XKzDZplpv
0L6vIrqYF8mn46V0euME5zq6dN65Lbw7dVhvelXG45IDLvh2mXiMM76oJF6DRQtB
L3Mg0TdwP1bmYMeJBws6V4EWo1NRgGjayP7X5waN3riYV3OU4H3bycjceQM6+azt
5GDl/4F1c+R1+FAbjRPSgLJu3IVzJW2NL9IM5z1eCS3x5osuz621dVNJdynCg/IU
EoJrKnEn8dO8wKDn6+kWzHz4tEJLDPXb+8R8nq5rgDcCpErKgKVIgCBxGsqn/922
gl5j8POSr6s2NugIHztk6PrbxyfVlACTpwACLPSbjJpT2mGnnkEZoDBBDxyZZ0cm
KANT3kiIAW90unHtaSaY1+5/qYQEr151nPTEVOCyBoGnMmiKP46gFO0JJGkhg1zQ
1FqVI8Ecvornslri7vpF5+klX+wadJ2uJPj8VkagGP7Lo7Kx6o+gFgpiP+t3zQvf
MwyIP0PXPC5QNNrF0JBQxETtVGEx7hKikZZ+PdFnjmKeaiUuG9nFY8w3m4TRPrRF
Myzo0H2xEoGSgZXybd0IX8x5jt67IMQT0Cr07CeOiLrfO37NCj6zW2EnoHW2MH4f
s16CWKt4ayRdOrm6HA/cMhtmqR5jxuZ0oWqaBf8xFp1uHfJNtte+d5bZWPlCSzjU
0B0ue1cpM1M3B6H5hE1nARIIlGalQl9LtfREUdnkdwwsvCCxwqg4V4feKybCc+cq
Tst4Z1dlDYAWHsDbGitktqmRJ6MFy80zCeOSH3yoJM9mrCINk91IEzA6XASUatNB
iH3D78f/bAaPCIYrz36Dn/H8Mgp3rzSt3KMg9lv83nSr7bBeVnktqvGEMdVW5UWD
29lE4zq1xiz5VHTyb8H6w8jGJso3KlbMzjcg6KTmOzChzLVTHnfiE1v9obDcrCxF
vIbYRND1NMHGQ2j/cI4e4rDM7UTYZN6Tt3XgNiNCIuclZyzQOMp5wwSWuJeE2lli
FDVaSdG69EPldZMntVvD9PvpZ7ZUt8HkRzqM+g847B58D2uxkXgETZl/lbXC8QBq
sUKl4DyZfiLdOTfuyyY0zasDDkmOy6GQSx3v0RHiqKSi6PN+S+26RSvX2jpLUpe0
/4FZ8Z+wq5+BT4RtSt8V/ZlFvF+/DLXg8lFj78HW1kUtkP/feqbQLaTWf2qAcMUx
45SDHQpqna+q7qliyY4V7OUmGQIX2tdZHnyXObYoU779jO492Mtkh2+x+UVIVVvn
EaDgOo7VqieF27jrUmxMdLzb0TnZ5q1WOtmQQg51gPKE7pcn0UJ41ZdAEp44p+3b
VWRvMRYJgJ4SvcicwZ6539fvRMs4SJ8YUjg6GcCTfy8OYI0mBplEqhP1EVTIIttX
SieXl1Bwo1TjuE9qg9hojXaScLXlIjvifSqJe6n/byA4zILt4SlT2Q8b62sB3wCN
v5jg9l4V9Si/52cWsrDUjtbV6cKj0K230YWEYFLl0P6i/IEnDfLd7aS/FRMcuxAh
OId8p/pEL/0/378Ql1eYIlL2kbm/VDj96JIp8ZubtcKTx5yrA0Aa6Tg/76X2/3Rg
phHM3GfFngxHUpGIZ/owYPQhPAR7uH9pT3Sl0wKn+VRk5H2OvJnB7iRtLOvKoL1k
0ZHVO8Xj2/VvIGV7KFf57b6UBt78uRdh3gn0FyEJoEim6BPjWz76TrfSfNvT/DQC
BGC2eAu9RgwXd5thu+acBNJpkKpVfa95jdAT/kpn8IRItzXRuaWMQcuvd+DN4Wyz
yOblGkttF9DH9RRXxMuxxlyUiv1tHlPMz4GR8wJFp+el1R67WkcoHt60VsD20AlQ
yCYrIuKRfV3yPnrKom5YTmIYSV9o7hPkHlnsGoDHNoU+u/ihCbvS/jmTTFgFaIiv
MozSfXk/2BYr5KtcE2ngkJ/iGi/ShRYvW9IzqQcLkB4BnOK2NnZAD2wuUp3U++kc
PQ+EW8a+NdCvDqJVjj1ZzxyxM8Grh4v0VnX/LSKxLY48Ip++FadLIjfflFyb+Pdn
QCUBRj09yNQrC359vSlzuVD7Cb3eoYNte0sZ2dVwY6uA8CAfM6OCvSrzNBcu88Bu
vRUtvzYKhG1ksV4TUUh0GoXg/6zk1tCGxtjfjFz4ACnWrjE90A1w+N/jCKpQ4q9o
SBDlt+kND+COvS7k3030RdngZefHdq0cWmtYoBoFw/LGdse0Cpk2day9I65y7ejP
gX7KOb6ECdvWjaHKlj+rrzLq7Hor0ryTI5ri5ckBrAef9jDn87xNFR4tYOxvhRl5
hGiGQ68jmwJvZMe5ctkx0vHYDuOAPpeKPDARdd+67UXWWNRy1vt02S/NhMz3eNC7
RHNpyVevyYD8MA1eqcLTRpLS7CsF9VVxfk6FIFG6a/TycU41aNMtMlDBl99orUa0
kUro79ajgSjk1naJ6ITv+bggbmSCa1tVA/nRxIIWOO1juJf/YWsGi5LQZh4k3/RE
l992yfkejKXlvuPLqrj6AHjMUuJ/sX22N2w+RO+9BF+DhoI8AWhehRYf0OV4RgUy
DQ27emzn8Pp8RlmV6/LQzGyx0+jVb6cTZhVa3KOLo/EahoO3h3TvTXCUpKtj3I8D
TxklgUjkgqCEh65yizmvFJ9/N2i27jqXvyzw5e/YzXJ8Ow3slrEVQTUB3GFl9W6F
HqD2Nzck6EnVugNzwWqhjUz32YK4nMQgaFnPuZc5riN3dZA0ZJ75NCX9ErHESGGG
NDMJnhjmZnTieEwZNJWZi/YjKbdJpOqKiTRem+Jz0S09da/Y7DIZtDgllSEGCzpg
9GnHaXpjXV0q/tLcZbwPOwHPrpk7hacTwViQC8y97tAyUGgSzqr5RaUoc68DJeRc
E3cEIF5nEz0ZF5k3Xcut5xzS/Tk43A3jjhVIW4UZxRjTAiV5+O057uPkEXjdGtmg
CqyL9NBzOvH8OLeb1gjP7D+1O33ZkqZwtsI3bCmwF7lUmVgj3vVVmusO1i4RlflM
YhtGW7dYDpWqjhXWJJUIQ41dnwWbFPWgx3+KEHo0Cl5MnBZadnSltcaS4UZs40J6
sOZshSTv20BmW7FZJFrR+8SEGoBHpH97l31/MwYYJlDgp5qNt55huQFO2JUc2GQQ
m9/XXRsDcje1QkA+8nE2Fj3K/QznsBbpLRpmoayw5lWjv7eUHnR+GPX8vLTtqi10
BMd8i1ST/9J2b+3ELjTcj+P4WLt8Qzw8o2xCjGMICXCYot1wChl4X41GOR95vPsX
OrZFqi7Duoj+LLaSzC7vZj8SVsO/+sjAU5f2hfJXriXaAMVthmToql6A3FKqotft
rFJFtOF+UlKKl3EfB4KKjx9UNpB+z7o5ipyA6loIDB5V7XDjKe8ccR8a4uVealxb
shJV3ReUyIUidoQIwpusD875mDIZKC7Bn8ArcfqdefGjIOc2wRT83GsKFfSf5Z9c
L5vFWQxqDnURuH8sRXcC9tqJdpqVdvC1OGydh35wmI2wtwNZ4aO+52g8AlY7ynGw
HwMOdFbHZ4TB6R9DzwY4v5knbDIQF7Xnpsj/QnnFlSIyb/CmpsmmFXEXYRm3i88H
J/nfXRfeCZmX3gCQcLqfAXec30lQ+9ibZVt8z816ZU+EfcLnESiicmUQrDHL7xH2
eS1tp0y+9H0W4mAbesyeEKQP++GVfKcGlSiOOClhmSXbK6JMnjKimFPQ8CykwBHm
kMyQy4/7MdkMlLJ2HOrUPF/TOXLzcrW6T3t2XkZm+aHy3fz7HkDCDFcWnH7VJSgF
zjqBWmUbw5no6e9jbs0Sg42uLp7jfX/WHvHaZRL9riKefjSQDAjaEZxG+Vp3x05z
w0tmHBTmlrequKCCyzcghHe/Kyin/wKvcgbGSA3+E8yvo1/UoucWPZrKE+FAQzvA
KVmw66P4TfRSgBM3D/Xe5qGtySLgLUxK0n+Pwn8fs6eaDydgcU1ikgB+zl8RjLqI
WmFqr8Duh04Ea61VXSB1NszZkascajZvTry8vCQJIwfWZb6MmI3gfeOx2swjILVl
DOqRTju06e1g82WBqXlS/ICLyxTIPJMDavff6fDwJ4pHPIXGbQZ7eonttKQCGsV4
/GKgA5YtsG/wnRaydFPirZEVo0JuzQbEZxLc6ifrN48tqjaOfxMCHIcccJC2bQfz
xmSYGgzxuWvuOHP37+N3iAK9C44+a0jrROWAhPPvU++vspGt3fZ/bGZvqHEHYzBK
rVqgt5rtIXtuSdcFas+hoKVyPUS0aMOyl/q8RQNvBHKXRN+0OTShXo4I6fQfCyc2
g1AIyaBaFEHNArhRufuEyhSXjXVnoAiB3kBO3P7OMQUmiL+6PkHZdGHMxYWHLuFK
PZMbpZ5iOn8O0AeDpo1coJBKqpOw7+qyVkaNHoaZcA7WrLCwAFlEmrFqC0uLcUWu
8QDeq8B9FSglV4YcbdP9LZ4kKKc9deF2UypDSHjm9XuFBocfWcUsMjZwhx1c4gTx
/vTwdIb2rHo+6hwReScBFwgusOKrv57QEclPgfSmD4bfoJv/ZN2kmlVh2DloEdCA
TXpvufZP08+nvVaOFTHD1N1VudpkagJUeK1LyXlDJqbv4BEQPNLc2FNyW+EdbSV7
hZ55F4N5rD4b4App6tqQqHzKTS6QC1Z/omkms4MGK5O1J9TwUJyFIY38Yv2RuSaB
mvYLij/r5AWc3Xd7mR6yUTbyjCu8GNHTE5qqocU4j1wMuTsrDXLvjAGE7OTf94Y0
A8aFg2GiFGG1TRNzj3PQjrnKfa7Xr5Esm4prRlNpoyTzxkGFIgngZkoGHWsIrHY/
ZUYp2R+XqdjR0CtwSYCjwSfWXTy7hrMGmjBeNZAGJsBxoRzygBc2sXXsyDEILuHM
148aUBj/UV/nko/5aAfOp8knMft95wcsspw+Cp/y1om1CX20vuRBRSqG14rY96Z8
zcyj9Qw5ETnGa9kljcxbfCpE5iO1QQ5XwE0k8m9I8SAQCv7jW1yEIDfE4B+43egB
N6FH5GaHhtHEBFN35/G63jCRZ2LgdWpDvHFndWTrDYV5wKvU7dVejds8rISekfyJ
CHvjuOgdRf5e/5xgLfYxuh0OCCL6GTgQrPDN6q7YJ6UpQ4oAFpyfcDNLpm+CaWnU
nsCcSAYPnYj4GXzx3M61KSTGkKqkYP0uMYNk31dpKsh120MTely3qk3SZOP4m+CP
J5pZUTj2pSxtJggEgjkwhQ9lgkd/LOox2Rv/27mE7S8jfdyFhc1NxCMqv24kZ+eO
CixDh7/dyeEK27zW6E/KCOGRVPBNb+uqpj1NlwQH+hGQkrk/57QRkl0O3jOqDEcT
uc846Qm0cjfPCL4+8KgZ1Jld4tymqZv8AoMZKc1EjEUa+o5p1E4nlkHTbu5VSGY2
gt9i+ouVGYUJELvRlEUyGhS0KVcdoKPA3KDrla7s5lNnpQiShGC3D60MkJxNlvd2
3J5cVkQfzEKO2SNzbG2Nryxtx+TlNIYmCYk8RdovRRPzyZdm7FrIZzDWwZQ4Uvjz
W7LtHGZagsM6wjyoD2O52+8bl5bg2TxplkDNqYh9DXHJ8eQEmqalJ6XVQqgiW+JE
4dyThAHrWjafklh8bLPTNatm2FhVwDg7duMZahoFxiFi7UqwCO/MjZsJpZrbk+XU
0qJMY0ujzfj0Isjqtx3UMHyFVX9l8dT9rGNzq29jyTE50OWcKTEDTvZ0lUlAaa4u
0QiQrLlNKO9Tefc4AQcTLPyznj/JTujUgb5WzjoBnyitdLJXZWsoB4qnBMzChSEO
B2yA8iRblSDQZpppPQ1yw5cNPnxn7VAgmYcXf0slsu0D5z3AJ2RxgDp3mtfHq3YR
glJXohOsxk62c8x9JPtUK48+L1evMawaLtYUgYV/XMFircF35nhLH/DLY70QWkk+
DrgCJ8A6tAd13YjbrgxbpBbyt/brHYhfkYV88fvuOCpBAvx/XfRguGFJSQO2iHVL
J3Xg9gNINWYA8czWMkBFp6+d8OHGG7bW+hLdr7YRdS/wBQTch1QiBzTpvIusJM49
s4oZYWY6ddE3CJX0bQUU269O4YxavRBDTFxs47ApMdUqN8asx03a8qbOk89uA+KJ
SY/zymoJWpJZoREKEBj9F2mRWybiqnAxuyNo1xuCTyHfdDptoXU+BM2/f7nQWlDA
9+vYHhUBeWZmEKZobupFUB5C/F05LsoDi+Z+em197z1p6//5kh7b7ZS0WWEm9G82
uIMd8sZRPDVxso6FGfQwZz1zUDMCdfpGlf/Pq8d4GDv1yQPUpIGUpywSzt47ncf+
/XDbqv+5N+l2NxamJ5qnVnnf5ApDPdabGqtQpbGxAwIVRgZWeKgIiXNkCxPgHxIr
RgVQBdiU9Ja7DqFpoVKbnGDjYBBCURIg7XvRVA4/wzkwpg1HtTMq78vZ/WrkOC/Z
IOq0MahSSvk/pe5ZNv7YklPyiEpJsA/IaH2wFwbsecPVgw+ckpvwxcVqsnp38U1J
mb2OHnGT1RjvK73/WJe2QQZuA7oL2MME0pqPl60quWC4Ivcoexmsb7+cE10zmWPw
3X91A9kcFZfmoUFybj62LyzOYv/vwnntfC0JAPymgLudd6skMrwu0Sdcy8m8IsVn
nmbwptPo2RatnXnLh8HaRqUHPQpNMepxKPwWmJM0WQNfOs2CV/V1sxXxWktmb53H
VmWScleQDrDETpEKIGNG3UPlrYFwl4HQ9z5dUGVKcEKQ1OrUD56de2c54/1xbuWn
HZjxhQ14SMh+IjsRQLvpuys+XWuTzwHAq1SJztlEl1vcKAV/bd3xQBBLtqHeT0bM
CjA6fKXeL6inpPGjsZ+KAGF4pfVyODcjSyRX8G/yMa2WS8tn2fd0EWsP1dcRwrEK
QXnQMCHTUzQ6EoS+3aaV2UgxOsVhq5pFT0P0K1CccaQ2cOELghzzUIqUaZev7Vh7
HonyxpqPc6cOuPnzqjSWYB7UHPX/DbQzvYELBpNMJjsrxbhsSVFwe4/9CB2dGxd+
0tTuri4XB4S3GtcZnquAE8TcbQ+ZjCzCDcMCmSa5Q5XP1Djox0t7TRDg6vLid3fY
0LRQ2B0jdezsqiDioeukfClMQ5kbPrn/oQdoXV8jqpwwudpdw3g3etDjoqjbPNgD
i7Yb97Q2MiOlnb1H4xu8PrZvfbBvmeVdvFXxsZ/f8SBlSgf3tBSfkt7f4tSzNpyk
yI4AsaKdBY+UJ7i/5exgQ3aKMDrFZFFJxHeFouKRKUIhgX4hpclb8xvvMalwNEha
FXj/23qCqp2YfTtpfzU/2q/5pWGmXG3yy4MUf/uEA/MadgeMmpIy3fIawGx6rgtI
Rpt6g/GdO3gDG8yOGJRNQxYvI7vstvW/FpL3Vj+AuCyUwqypiC0bZ+xs/+1Ip5PI
Q0VpOj2SrZwx0bpPPLfpAj3NKluGTIRgOLCcvJ1GwV1UlAiA5MZWOngVRWhVyubR
/l6BlTe2GDhXIqUqYnCGzE/z2F2yJVSkgTyL9kQG0zb9JA/vbjJVheCQfIncvTkb
yVUAbNn6zoStZymSm3XO8qGfXmRG5PAhuJBS52kK9beFSwBJXNtPVDwh8T1pEaHf
C4nxr2xcv0Qa0DT5poQtlpVv3nOx/ynjG4jf48+xl7pXkfEBTu6BDfZbqX9Hu/Rj
wKxEoSkovFP/phoNhmngK0/V7Lak3xNiZrK6B6srxOXnJuGVuQBx2L6bMQBA08u8
INZHvVB7SGxU+1i+yrfHnJBkBOyoPYth3XkBgmPFnIsuQHBxy3hadedLCsjsT7FU
w/XX/x6+tzMvmZjhyhMt07KBoo06VMEA5IT0EI2xPc/o/Tjs/pjYEWUEtaZ29BEV
ZBdyXGxcttjxwxy2vMaAWnCAvDgy4Wx2QUVrMdwfJ7RXLJIzzs40jOZEj3P6mMQS
/qvsMGuX68gx68eikXC/ayslbCTDQ9dXeE47W6MhTnlPQ/wepqxPNIuKxRPkE8bm
DK6Nzm6nX7ByfRZPOj7MijQvs7FB1OWCJXiyp/I9PvCtxyLM9gt+qNGoEjSsb4WH
GPGfUvBD5Qp2MNVPC9ovq/QJWjm1rveReHGzx9GyxCkUxYKvGrJjs9YnlCkQ35nG
Sf0gRq8sCyNfMJpyrBt/hM5oUozevnTk2+dXYkHEhPqtVGPCtUNZj7UCcsUiLrG4
repSnRgJ0yk0FEQM6DbaTNKAl0G81QL7UHjtDhR3STnU8pxRAR2WAuTncdPnlK+N
eCvrJ2nKWkPVacYJCJgNhBVUyPlMc4DuqHSsUBW7zjwodZJUK2xtzNYWxTNlR4CL
umSaO9xkf8EE/6cgF2Y2kiWRtDXkppD5qR14qqa0VfCEYajOBhlQw/UN4WnZbxG7
/7Xhfwudq2pjXwtccM5u/NRB3I7blzFxCYKCdNGGPfb3Km5ZtpJtTyFg60qLvJuF
HfpVtuODPXM9IFP3m9LMUbdNQTbcAC0MtVCtUulL2aKliGKKBdtEe2jPTe4a4qC8
Wabpi+HDM0SwMKkG2IQto0LtxUa91enOaAMcnptRhYL8Kj4gjoLng2aOYkuyk++d
pH1+SGC27hwV5n4c8rClJrHA0CbWwnqlnO8rH75vlqrIE7zFQw81750ru1GEqyxs
IuOzSgCGQy4UXffYpKILNRXgUz3DCx9m+rzR6xneH8RtxnPr2v2LOJPNdRM7RsmM
iBy+UncJMFpI3f+9zbg9m3q4i+oGUyJ2yatjb5onL7idU8+ww2LI9UxcGbLNwW0M
L77YNavnlQjb1T7lQJRU9CaX+0hS6R5/3N9bhKHn2b6wHq4sXsKoFRm6ZaGP7FFL
aN3gOrS7mwR1MDzDwdu/u3p1bo58yX39EKhqfCGaO3u6BAwzi15TG1x4M2jmXEOb
yCnYW+UdRQt2DoiUUVEE53xGrYgyAMU1m803nihaAaq6zOd69Pj5xNmqMj6KFfNn
qSh2Ap7GmSykRXhXK7QX8RTBfnbag4xrteXKHCIuHUOVhkWW8o4QxDnlKD1Zb7Vu
9rtnGiWLZU3lBJAH2eroWMhG5wWFN41kePcxoWizL6TuTTc5bGab0uiooU+ZD8BQ
gLfsjBwcWOd+1TpOztoV+hV4ZfB7ufIeWbpxQyB+pqYkhiNQLCy3yHZm8WvyTBIj
wgJAZ7e3QPNMpAGy6MxB1wD9o5edun/bP2nBIIZweLCSaojxCqO93pSsb5edhbNf
qzfnt3KUuRxNlUTljhRU5g+Cz0R/f4LBdMJJUAu+cRgLtOaFn1fenmJvNgVvUur2
8lG31bC7caKjw0ZzKgYghMKSJSTh4N2CJDCbMC8RxgZw4L/SmYKuVTPLW4AGqdeJ
81M5+AIM6hkRPe7HqeaauIUhmsPhclMmLE3SltenrZtuCz9uzxhebAHlwjnAwPuk
X+fY8x6QJnfdE9Mwspba2IEpDiIglLoHvKHp+s5gOg58tAWMjoKLUs74ejGq18JR
FSKd+l50yHCLbRBTZ5K0+39C2QIVbwGs4y7xlu5TBsQTMfeHx1YS+bbgsmfQX5Mw
gYBjWd8oMmKUFuKh/BPuKKra/TSBwIYsBIH0E9+YZlV8j1n8bnVFKAcAMnOQZmKG
mS0it5KApit+y+53+qcjiu1Ru0lL5r72++lLFhhXb6THAZd1s72j2RTJr0WXmADt
lbmTGp+7N9LuflnI0JmKDqiu5CBF87+0KFaLN2k+J0X48hU4Mvap+zZXXETQxasQ
g1LYKAbgvgfVIazEHt00tUtUNJfvbXMDh2OisTpchyDjV6avJAtHS81Xmk4CccDz
Om644ilyxXNrZacFVSaqSuZoxwkeC+23ww1l64czIHDzbeygG1ze90lcTpvcFzQ7
2tpYX0zzmeRGULebNb1kmqM8bAC2MJtyLCbVszK/Yr6SkJNfUCWrMAusvY2qxn1f
ESTJJfBJgn5IYsxxiriSKtSk1mBi3DVp+TmPjCvKVM3loZ6iZjjHhxV2MJwmObcQ
bOFACL2IfzKO+n+G5IYFd9RyiHSTFrtUKh9usJeMQesJhPCoGY0uC39TbzzgEVNG
Gz/6WPQDmJLQ9iNyZzpNVgL548Vr9EJwyBTPzB7R+r63rhGcvxTZn1djVrGWrzbV
xUuOr3DNyz4f+9uaBswuq/05sooX0qqZNdUOAOl+e3Fkijyo2JRwpaMw4l20DFIX
KKpoJTHtuADJsakJarXCStjNiHUo7KOm5CEcrUgK8iF8cOmdsb6B9CoovukrYci3
xunafuyt56SKQ/QQvJ2Bbvnotqs7JeH4GR12ahK2VU3NVZFNs5lvTFDWO3kFdhrQ
PlWVFWVNsjsAQyukj9+7PpmHYlviC6Md87qz4MECNs14e5ZJH8Mz1X30oLY5VquM
0qskSAj7eoG3vtQQ4usM3mX1QvRQXFvY4V8IRIFfr2ZPZlhIQAOOBf2c3DrZmTvl
5SyXDfVc10ULEGo72RQKfblvsvMs1W3UGwLQXklnAa2Ai3G9xsPxAohgFBxnntCx
ipdDaVue9JFNX6c2/3S3m2r6kxUvM95fudD7Qf1hlEmtR1XBKthAvzLE+Laqd8FP
382qQ2GiGEK9SkBwQgHMxF95eIAY6BG4SoiKNBr6Bqmeh/7ICFAFLln9myYiP0z5
V61iX5fISoeWoLdMsqy6UntbwUHzR7g+1NBM1d9Wv1kdJntTKrorwAW/BNI31Ear
2zY87legKFAxBrS+dpntafkpEoLh2eY4CWjNNqMG6Nc1qiqzT1b7Rh+xMLf/unWb
fSq42cC+tXLaWglAkp2s6IA2G8RRSDrFZskygjXyWPpVEh8UYNfq58xnk1nHv3Up
1SD4mSoYiYbON+GxeJkqCSwr9kJDZMBjjmN7r1nBwVtcasECmGew7HwBjmrVSXzA
/yTcQTY3n6PM6hH6gpXuv9zFwRF9V/Pe98zp8ySyn6SAYs0o0b6XEczqy4g0BdCh
wbohqMGcKFOH368k+IOqolxa/x512+B1KFP1/0DeMdXlxKUgpQf6u3WJ9uKhYPc0
KszVUBEQmvuMw+fG7P6x0dSQFNl2ak48p2fQQE2LuN05SmGDkg7i4/LXM+nuyrcO
OZsDfr6fRCmoRMJz6wiIyie2jnrV4mbsGtlp2asXxp2s47sS5wfSl3DOSEwwrDLu
ynL3/zN1dJ2drJNIascfh5VIHeT9NWwqDUAyW/HaOFH5FPa9aqPQcwykwI6t0Kmb
QpBwFF2ZZY+j6X1WKrAGAjfYxtp04jeSOOz/yYQu6QSZeDQACh+rdGU3z2um0iR/
kelX0I7FgxmF4e+qTpJ2a72UgHoN8u9EkJe2rVy9QMSvDwqv78pfG18i6XvYv9Gy
0IDxBOJQnHvgv9vfRhjwJgrKTPbez6OVkxss0rJHfEvQoOFrhR5NrlH8IFb/P86t
L1Sjqr70qidukXKhmZ41AbbcwuafuN3j5xzhAeX6YNhI34yGaibG/3KUmb5UHWjL
XtzuJgsq7EHdxAvx9SrFy222nFVCHYdLjD39nWZNDNFiS2MbqPomYPsD8HktSFPJ
/628/UQRTcWq9JzRRUF2veNvWpNB+AQ8qf7ylznhTXSA/pZhjnT8C9rorXCBxEKI
+pJSB07Lbz9WkRyHlEXOMA0vMlocwWEJod80mZVWImptpbtAWaIzHsAAe7K+aSug
232SurQcvdcMM7cND4/UdXBkpbxr4ERK3VEtobbx9ybgxq1iPL0IcdTzH9vtUsj5
3KI2PoX4jQoasMdNvu5dg1G2OXVYk8giSyiw3af9Qn8suFqv0ri8rsEyxzWovT+L
DQ4TMkIFioF+RpjGRklkLwquS+GHrN39oYEjczbNNj277Go1AZtso2ZRJ8kvlHLM
FytCB0GwpeZyJ1mG7mCY+hkU71ZebE/44PwkQxl/8G7Yo5+PkaVL+/vvS3dnTsNl
OhqDI5nOkF3OU6IN8s3m3WluUt1HQiH61uJzUWjHRUh8MF6dMVgaBJ5S/UgSi13y
ERmuXtV9vdlIlughx4v/OUPuK6+h8BCpCPtVYZWIcdzXT5+wDNaepZj5SMSIchpL
7Uval4jytwzTvWUXX13/5e9Csid9607/2tj7xl8faWg0FgipcjxngY0jtkPua7j3
GiMujXGjBianb0hD6ZuFfksoUl28ip5Hp4pufLexcXFNFFilg3ms54oVTweQoGAE
iG+RDzBQoKffB4b4GW4pnFm9Fko5QBGw72twYsetwoWwS7sIcpcsVD5TEKTP2iu6
INFGK6EAdRssdgt8XvSutUo0CXL4b+53pPc09SwD5xX00vyaz4p6GwfBEj5E9mh0
aROaGrgofTtf0/1kaCmMNhUH9RtUwpVFnRqyceyYsyeysXNmgBMoDEm5cKaF0h9Z
jC7LyZ1EVVjuWVnofADIx8vjxfqVw28u7nTyGEjKx1JniFqdB4qRbuIzGsxMI2D8
7kq+/IqAVg4wKvk4asAYUb6/hhM9TPIv4VurYhc8Q0Cwx27FxiAK3VIjrfWizGpJ
PEKcmHZvkzuNrCSmz53v72c4yMbkU/fOt57c2f2G5dwKLoyNs4u0RLQVLExyAtnE
GXJCozVs408Vt0gtgRRxPcwH0cprJZpvpT4EQlVzjgRkhFhDS4YybxAoEsmkroXV
8X+WYdQJNTFHrRvUCW5FIC7k2k+vEQ4hjKRlfhMt0JSUnDXQKgGaIN9j7WH2HOvp
+/r3CrFCYgaFcIoaMdNIfVm+RHRe4dOidVFVMFsIWEfBWjSY/0hMov6w/PwCkQnr
EzEdkAoOWzs1Zhx5NSivFtZ2nptWqiLpkU4P+NF6bWJm+W9SQiUG2tVftTEyxznU
KyYUHQpqwPkK2umJqS6cLPqTuZ88muKw1ADjNe5ppySUQUrRIexZaAjVeMUJBXra
RvKJoKoRe6OscRXn6OvLnaA3LYUYlgwZtg36H0+OjZSQxgKMHBo0/fXoYZUIWRH+
7bMJMyUiQDKOXS5o4CNuDA9pl3QdOQY2Y4CfTUQzo9jZ9rhPJw9TODsnLI1hZPvA
ijkHpfjKPZuB08d/xHkuxp2N9WknsqnauPIFtx+G3J+hkRm+oLdIuKiUUDQ4qeEP
I9e3mb9AM7qe26sPy7spVkYrwv23Q1Uo5wKL6dpCsQZQiUOqpva/PPHJbJ7DkUns
17i8bImWURUFTRNB0r+5T6i77i5aA0nGfOIeAV4N0cCEksdfgS28sw0tiYP/2OKG
hBpSAz365/9v4Y5TgXfmGUl8l1b0GSXKQyASbeKPtMeoSUwxxUrcv6yC2hc4mZVk
39Y91b2QfnRpORyGNqEv3/gRjM7MEwVei43xLDYnS1SumQNI9R1VKWwkZYCWILDH
Xb4ixikiGs6TzIenpWcnlg2UfcpeWuwaB11OsraOilWWq10lA0jBxeegGAHUhkxv
BvdW66dTW+r7JzQ9f5wSTOcKBgNBJnUnNkd5pAuUyBgyp0hv9yagQSNpgI3Zu6hB
3JLDeYT7BdMIroX2gUQYqGwefX6rNO1OaFM2wQkvCj3mKrSXqKGIKQTtF3xGjRH4
JGvhGnaXHAmjl7nE05efMNnw4XWOLONIsA99wXxG3wLizkn8Z0Ok9hORHK17Hyzu
mO6w/zJwgl8tCT0FsdawAI7dNW8vgbZAjkpJ7LkbOHsvTWv1e6Fii598XyURKJta
Te9TOHYVDmb/UkOrkz5XVu2sd1ND8Ju7Pn1yiBUYvio/BcY7QIK/ggF72zHOyq7/
aOtLH9DMxz9UX0MNMRTFf/g8Jtk43+7YKjo8OZhT/CKHU9zIAgU0jKyepED4I3Qs
e7/2g5J7oOZTkfJhKOoCcJXjDIFaJXQ6kYi7SVCUjshytdjGnrtNSdH0OMNXW+kY
Doi9BwdczAcIOb7HG8hqneU6hASJaoNAhVIt4IQYj7fRJrh27Ihck9W/jj83R/VY
Ss6TPgc722DbVj8fBMvMilF4D9Axuy0nmS/0xQRdiDYswfcI7KwWY6sBLhL3qF4/
WfDSa5e7gsgMkB5USoQu601qSrzpKdcf9yEFJDaOdDPbsKoLr+hG8A5Hy+EjjvrN
3c0JDQCSMkvZjdtV4c2sUs+BgNFD0yTvsLNJ+GPdW9b5uITFNUTuwJKKWHK0DLzo
oOvgC3/C35aVq4kN+QXu/ESahMmTioPnv/+892WwS1TuUxdQ1Cb8f3MaAAAboAIO
DKzUQNTzHMJZohJlrLXrlQMS/37pS6eqtP3Pl/4VMJo6eCXoR07BWIFCoubtwyVv
s11H9h/Q8Mxmp6OeaXP9lN/oK+AudpaFxb5N7Akr5UV+ktWTAnGJuTYBG9z3Fwo1
LBC/FS5pMxkRv1bJJPZutkYRjcy1yiPqHYqozpH939YWZD2dmmDc6TMlSUTam+kB
65c1sTqrtMwqPOr7gefmIsGrpIn4UBns3s2IcOLtU0sSt4mWWRJKEdiQRwftr4x+
De/xWRgEtwiubELixA1hRjAbuCV9UJsJQmUdrqsaS/sxSWYN+aAWdGywqP5bFcu7
QHmUC1S76YJkPYQI3pJLYFiH5ktKpwt7tr8143oqvRMvnusRuHyiY7sA6iHQSM3i
vrlyC9qdCoDrFKpon0HnRldWVfjXF9PEeDgp49rkkYCJ4uFRw5z60R1Y37iaXrHZ
T5yIo9DvreTWNrbtg8nQIo70qmgzXj7c/0DfVmLuEiZ1Q0/EIM86yEQW6tXkxJlM
ifEWoXfLARxASCSShs3GMZMG13amDbXMaThArN3Exlpnh/5x46xWFFyodhVSkzDZ
Vp8ZSpbCaX09iZ+NriVy784SqAPtsB35BKxaMzf5ZW9U0UDvOYPHQJ3CKOwbdSB3
uqgMTHEQUK2dKytnPWeAV6bMnfShhCJf1vepU0eklbHEx92krnXalKMdRnVyL6Qp
19c0xcOEZncM7H7KaBbIEZv1QvU8iUwDX4zhuwSYeUag0eXDkt/Fk25GTmWPAMXf
vF90i5taKX5gAmn41BaxNbaMWuKjOJWcvC14s+GsVQuwIMAuHwFgUCuBty7uxuqV
cuaMKRC+Mmkdig6q9Z8ZEcnLhOG7gx7VMlNu6YTIPwI3TfEvQ1PUkD0OsDIZCSNz
uRMlee7weKGXyMaRc5tFWC+ytLqY3TPuFWs8BhJMORtUwye0q2mjktoNLExPLmSL
siLZD3lDLwZ4ioJqBlGhgpNQJQqZaY2LgOaRdNpx5OhGa6nktG10r8QDXW0QSj/E
DVqzmvXjEHRzaYp5+x0xz4wMqBA2r354EWqfFfe3B3EvlqsnOPqACq/MFrQfZEFQ
+hAAATixatWJdIvuW92T5WJPI4i0Z7NNTe0EDHJH120kh5h+CMU8yEKMwixAMSwO
rUoJwnPOtL8DBqFPeAN/A3KgRNEp/47nEuG3MP7yWbhCNJm9TTje2YRd5LLDGnBp
fr1MWyuls6jW3NsT5xcOJXsv/rTdmD7hzmz2V1GZUrnBhDzYuKPzg0Uq2kcEGWZS
20l5ROEUOJjsVP4/nx1EtCHpSoDL1H7L0fmaOtylP0JAm2HMvzqrIfJx//4o9X27
OzECm9InkCsrNXt738UGQ7+lK8aehxxhuC0m55rnCLX74STk1sB/T4Wi5VK6keLK
eTU6wgYw/+MOZea7ghXxg//dSrBv8QINz31WG4q2cVPKXbsXnFjH85krDEekYuLy
3GfOXK8ilz6hS6E/cUqNjQrpHz2+BVlX/IYs9asc5lkWIwixWigfxskPyZm1KfTv
xEc7qxpixgeQSWCqzljNj4sclS7h4D7PqSr30AVmQQMswX2U4PvbZnB0iThhX2Xt
UrviemxT1L+NLjvg+A/EAOOCC8+CzB6vWEvHPofIqVpjHIM+AKMySJZ7RQklXiaC
d3mAMxy9XPTiffCuuEd8lt6LHsizc6AXF3f/8Oc5zbYiQ/omO9hO3Fb6inR+0RgP
riG7uXKh7pfKqw6LoC7unP2UxC5iA7F1BuRCRhu0+C5sFvP2t2y/LCLGS1Y4y3Hy
C2B7K9+GsBkN3fvKHbJUiLkSQkAhppo8cYznSEfMd2OyorQfQf1slw+vUI2VmmkF
4lC7jXri9kkizpIa7sgbtA0tco0ie1X/Naijr+hbtHFZ4w0CUH3ABQtiWwBh2Rrk
bOr7PyFvw+ByzMU8T/hWnUAtKLOs3wdvEHB3yVKhle1xL+OKZmkGKOyfoXPg+6Rw
4W37s5RHu0UznKKaGCoxj+cn9KzEpxv1etGsPn6LibF4disJZSdo7AjQPEQ9caHG
HU3ybsv3PqpBhoMZTGNB9H44DBzbVuP4lk2/3equC7xP++y5/SrrOoo0NNIeFbhB
TwhFN+CwB0dYyvZ0WjRIt50blN/ek9oP1vKXkifNl8y7DwHr7acGiO3MBmKwNE1n
xfu/eodng7zjCUDPFyG0W2Ks6mv5+RJPglNFdRtTQhV2zqM3VNK/H5OgcrHtvlzA
aWAWOQ2X2qglqH6vIJ0S5mgwzOWYyTTsMEt1qp0XsdT0LR/PtFJGN43QQLxVO5u/
2fIjljpqyP3cU3dHIp9SyxVK5wc9oD0PDR5unO/YN3fgGrbidSaKZlp9+VW2jU+Q
TToXlylycqWTBlvRDJlWK/+e6Fejpfgttgv8D4XwOtAoce9GtYJGzsgK7qwHx2Vo
LgqmDGGp1BohHgd7Zl7Qh7k9BpF8r90zuGk+siqiuNzbf5OUouhQ5KIDODIFSdYF
tqPLBGmLb6OkiKUSY6wRgUXLxee2Smp4RjnrQBNyyYcHfGuB/8j3C4gGBXNOj8mL
vII3N0DGKf0Uf88a8m1pxUc+tlTa7/dNweg6gYx7Pgiv2GQ5v3jDhfdt6AERTHzR
5DM+C024phiDRMyWaYMh2kBapG2xoo2VXUx1egYHDhRfcnhCnt8FnFHESHZ1TyFP
d4rXPYJQGyiaVJ6GLZHI3R7bE58H1b9pBn22s/KiHlu/SsQUtpTBa8z2EQDq9PiS
LW9YXm4LfvSb4GlXRJhumWUwORGt9l+9N3kapX7Fad7K7nQIT09SDklYJYZzbRyy
RR9cuvJa1sVPFMr4WTlzlRAQsL86l+fOlYO0mp1GVj+U8hO0O7ubGgtGFkIlBXqA
rP1KGT3sAwOIHg5hBn6BXOq+8uLhEj5KVri2lsXw5x1f8kTuRjFsUdxwaFZOF+qz
LYijWXD8XYw+sNOFUJLzBX7KmealAzeSB71/xdcEgv/9aaiNNXw+p23xE+lwcOHq
SbuM6HBLpyWwrz4/2wcQl20/TgBE6io3nmT7kqAuWlLO+uTX7lQbYDjGI0ycaSnf
cJuvszCoDHfiLfCkF1r8Oi/Z1a71CHXn61bK62PiKjCddtrjAaT4qiZ2bioLGjYH
vGyFkRWIQ+qwbToh6KQlNt7RE4qbD2tvbLtPp2QwNtI3OMLTiH9z5fNuWg28SHd+
M2OJ/k7vGwGQIuCh06kcDDGxOt4xJ5GeN1EHjStEx+4GPgB8ykbxwFUo/KiWzG3b
4xm6QCLxuJq1fCHkpwUdALG721yhmQtFz4apnPhGE+qhkr63exga4TehU2PuB0xS
24FwQO47nszgaWlDuRx0kFE5+S/GVksYJ5noe2IoGAkBk3gXrFURanCBMZLjV33M
Q4lZaI+qkPVhjTtRi3OBwklXP6NH7A2DIWQP5jEBuM6DuQDhyr6n/al8jZTmLJvO
mNZeGlY451yg53Xcd+s0/Kv9UCZENYoJpKYA8KLYZ3q+l2LIvBy/oPujMwDFC0uw
er4sHvGrAl/wfp2emya/zE07Z2eChEgY6osdmhfNlGyJjiHtXSfAS1a9TirmQs+g
o6RaEUirWVIVPUFYn1nm2Nmbwr+fWGwCzt6CP0Fi67XYrKl29nDR4+/BkeG9Ht1g
G49rUxfmnFM4YtRK+P7EDs8ea+S1YVATfUYtsKUnq5DJA5gpcOPNjEaVggIAyDS3
qIjJXaPSv++/6db3W5zRxRKEfby4DZ5aBXvLuS1GtjMSFTdCwTrWpdCYrIlH4h4A
KItuRnfUZjgZEb0s4/nUHaSe3kF5s9z0MIsA/ZCEURiCt2HdkXSmWiboHqB13/HZ
OLczmdNSTHAjZOH8jvZktFuIuZYFo42Bc4HbO/DCxQSufOb/AhrqXPBVNYYADIYt
X7MyjixW4m5E8EpfN+ZBBi3mhrf9J67tdnHPGCpoFNlfLnlKSHb3RqP13z5vfn7t
w5dzEaBsVHIdl6q3JXfcU+5tLzKbpRiBu95RL9DG7XNoOmxUzOD/4w9vBAdh37OW
saYtqmd5/p390SrUkXl/gzTYOEiAkpwC47nK2O/7PC3anmQIAmjLEGWLnf3R1tKF
FsKcQNufzYEOZLQ678MLBYGxc0c+Cw4rtIS097rgc1w5EE4Qjjf04UMCUsX7BB6D
ABbiXaXp5D7KkJNvY/tPRW1yLfhBuW/+p6j2GB1+2KaOeXFuImr3dL3DZYCGzI52
bc2rPQaPIUsE47MYzIp1ZlNYIKLOYVKZSCeBFFE8p3FDjDJcBWNb1OUtd5r3POSx
pKhdXbQZGGk1T8aD/P+inihJBWVVpOkkeVhLODYV9hD6ikL9nkxUqEbsZHEvqtGI
8uz5LDi1Vllg7GxPOjh0pMzZ6BJzcIAJHEX+swFEF8v1t2FJfdyidncEaCQLD5eO
keu0RT7aIhoR4+sNI5KwwpwNcly5mWSvkDZX8ekJDb0Gz2osL7EcBrrwXPmPL3UL
v6P9mnA+OUz+oPtnzDDZk5QkT1IDNkmWSo26bf2Bmdtcfeb242LCUwbwDeyuN8Ji
XvMoT+88ZZVkrsGKJEwmwpiHrXZ6BCqXXsJE5mqWEczT+0Y9GHSQnEalZUqqLbNI
WwCq2OeiN5jlAOt4G2rDHI8tU/r9hCGqxK+F6fgjFnOqmhDszkFDvZXQXFpP0jlH
4GCXHatoXhw9eGMnNJblruoBGbpnoaQUgLBfRJqJtTYGVpLz5NfcAGH6DNGJu6yg
2JiZWIVw8VJbfY5wkkcAVqKFTbkEgRf0L4X3nH3TVcQiv88gvcVCJ71r05PFyA69
PaEtTiLoT6PBilKR+7H+2HHxjWNjyAspTkjEAPRTKzblZb1LeX1TosIan3NqnZQ1
yrtNHd6ZsK2V4l9LuYtok490aRNkfrCc3xoXxIm+yoAJFukjc1qiqQ47qU7XKZYK
p85bZ97bLFKzZx5S9x+BzojY6H7bJOamnGt+h21sRnVySC5P02srSQMZcr2aZ3R/
gqUBWn03hbqS0CkzKnCqf6RtBsY7TsHOiaEY9ENWKuGCSd5xEIBj6YJ0ixvS5q+B
hQn2Sy9usq0k0Hhdp2yq+T7k7TmYvfHqohg07ESq76zzChVt9UwNjxrr486qdxio
ZIMeQ4vqjE3iUQ3J1/ra818iAW8vwet9nn/p9B0+v/TjLXFb9prLUB8EBhUhJZAk
5DtGvZHRJdh2+ln1l3a8Fab1NSl5nx1ImdFdR2Sfgc1JnhL90wXKXotApFO3CUVB
9GiS3RkczyDd+qJoIoMs/cElriXBidRfxWTCTAk41rKvz0NAO6Z24OBpI3setgkX
lTCARVTOQ+2/AQeSPYbU2rL95PUtMPlZcl7+mSoEcgzjlg2T1EpybOKu5XKaiiw1
Mbl8OJoHmG5Q9T2T9TDnVMTKvPKRg3xf7GozA9ByVgApVVhyHa0HIuJ5Aj+wrp0/
9V1/qKOf4fPh2lPGhKLcLBzA674PWfCoraqzEIFA6okEuCmk/iOhMjRl6hYOf1Ft
4ZkmzhzChMCtsx7rjHdjv5Qa5+kaEogotF5PSxUTjWuwNcFvOgPUvHPyZZmYwYQr
bYWlV4j7deshkzkof1/QHjOsHxlupol6XBbW7NmuP0hGSkVugeTlz+pA0IjEnRhm
rX4akUlIDl90paddN+aigyWcLWiwyVvm8TpDeue1A3djt4AGGt/Uh5pLwld4RCP/
+5Se+omjbSex5f2aJud7hqqWohEbDgFhuhDzaaH5d5vvOLW4a+F9AyVZL0LJMXZa
9jizPKkfpukYxoooIruGWiYldQBnqDO8RGxIc/Z/T2e++s0VfrlgW+QJ21TpLINK
B3sR5plLG2jdD5h5qIGI01HgpJPwnN8trsix8HZmGV05N93m6W5gFXzbdihunGbF
hERLN6ro7iQVIAPjufuRN2DggNI1tdH/HpGF4TSd0NrU+Ygk7oH8QaBw5x4bK3jm
JVs39cEjkGU2Ysax40OVw1dyfI+Nt09ewilRHREZdmJYTgyew6bz8TT32gOgb67o
KZeG6WbFbcI1J6eQALfbA3CGjD1ozZQ3JSKDKVg/JHYtqe1RKu+wnfdbgYO974jJ
ZOCcwVp9aI+ZVhDkZTdWZK/AcGlWZsVuSBZQlSQbsBspHfQqd1o+snyOBlRlHEZu
dRhZDIMvg1TPqdIB9XuvQ7Tx7sVbA1CPbe/kapFOZN02uQHSXW24ytd+MrMAbhKt
jec30DxctgFwTP5Uy//1TMAX2YeSVhGke+32cwWjty+mxBAskp/o1F5PprlZgNIz
DaC3Xcxrrgi5uJWsDP7UgUpcLIRtf0312tg5E68eay3l/iuaDFeDS86XeprHV84f
mg+43ectTevbZ+7EWb32PGQIRUQLy4GmY6ktardPeuRVTfsen+yna9CfVZ7+gxWI
zFH7bdvVH22Uw94tiEKGJUl5+NUJ1T5r8+9iYRq5h25yEtBL0of+3ARXVF/TejfE
o2jG2vSQhOaw1sbKFEEnbknay8QGOBpPjntGW1RHCeZWdOWpyTko7OcIVZgZdfhd
kpIu3iwGjxwsLC72rpoCXIlnEg3oXFb4wXPSkhf6HMqNiwVQrkoG7gtWAfGeNCEl
qFWG2XqO5ugyK/QXbTSnyTq9NiSRpOyXP0Jvdpu1dQDQrEy7OPl8Yi/LXHgje22W
gKUS/krtlnA/TZx6kvqoMdyTG4Q9R23+lfYV4+OE1kc50E+HPcR5nE9df4nJh8I7
Tcs7CONLqKN6lngoaykRt/k8wVn23b5YwoepQa7bQl6PaA/I7zDZPMUbtR+DLNJS
lJL18nA60ox+BVPxv/BT4nyF/Qqp5sHSaBYfNpnELaRZXsJTItkjpfmXQnx7aRNv
NS3q//PKolepeDsB768IYbCaCdJtwP+PYA11jdrRB/eb+ktjGtnYrrUFukes0Zjp
RMRx9qlbcSLrtkFD8N95SjKaC5KIyS/I13GaCg8qE0uK6bgKqy3pVg1a711IOohe
JREg561g93K3o+ddvGf840GmGWqar/9I28ObWG3eRwiFwD8Aqm2POtC3T3fYcQ33
BCpVSmj7mOXoe9en6ypKahfEyFS5wno1Ff/G+l9Um7djAwSHEB0IeIgmy1ebGJNA
o4jPftESU7VxFpKz5Sjx3qJVRyBTmykF6U/X1Oz4Zzw3lqhXFsNU7j7a4PvVVTsD
pU1yMUNl/TL9EvVQ6V3X1aMZ/cQbKXHI556Tfd4CFxqzRErLrxa/0RebgFVLQYjS
FWZ5jNz3KMe5wpH429+DJu50tWnruZEagpIGFpECuaSiNu9OgvvNVGaokpSm87pv
MGyH/zlJ6ZEnpzmg8PobLj/Dbh6XM9F89TZMasRD9zdriQL23zihAPduOYnY+Esy
bfl9ALUQkBJjhgiQL2qQc0eb4JVjeDHZX3T0q1zzDVGPbmtxTGPKe5J+dpBGCADK
Wettlzq65pKkqhj2kBra1PfCvv927+nbcbiZ4gijL/i1uQSvNF7T7B1qpcBPon25
SaHMwRZgD92XumKEuX7YvkH2cpuC2R+i7+hcDLRM8aom27V9z1TRFwrWaftre8BB
KBNbsv5A1/cDLH/G1tH4fR9V0wEoPK4vr3grvayA7UNsi4cqzISAoh9m6v9NObBn
LB9yzhWZClGUAkdIUCdtD6ZI20h8vHYpKZcGL2sp1zscsAGXpI7M3tzbYeYsY3hE
oR4YVWXFfWzX8T0Uzy8856hCqo6tECOrA/Tvu0ADnRAB79EeMZgnurfl2bLZf+i1
1K8fk45n1PGCm2Oj53QoAhk+KZm4o9R+hFCO+eFOp3fZkEnLK4Xx/nXtbLUI/ttn
baAiUCvfmL0ATcVQM3OA1+3n9w6QFNp1fhqwJlCrYjkfvNUWM2dNvZBMZXe4lIUs
OMksScQbDAo1WfqMTmjXb7m5XwfGxIjGfs/YonUET3NLHGwalEsGWpNddXFbt0Js
O9T5uUl+fueKKIF11R/CIvz1TIXtP/eLzo6zlseK1j3gLt4DLdnu4gOuuHI6AT+k
YLsEbdmZQ1FfmXrprhcsGY6SlyzIKZt6akwywlziknDRCREl6V6hT6ROWNx2FyQF
RDSiMghsSrqLOJTLqVAsWZZf0/AiI89yYO8CeIYYOL/+nWqWhP9zbGvvblz1g1UD
0yP5/RONhEEo/qnhEjhMc1oGof1Cxe/QiQg0lAjd6agXdSDTXWW1/bxdj79EbKRY
RntirCRiQiv9hCkzXlt6ftzcis41zKVcQCNzX7nJy6ItY/UjytxXn5fQr7pfieLB
3pJgD4ooK+4SRpAf/RoTAFJm+T+KjieRHm3iUTue6xwmZMq/ut4fF56V51OZVF2u
UF0fv7zWXmDCyoqWaglkGpFnRCGyY1Xo5RPQHFtKOBJLe30CVTyjlwvHrQUjKOuk
GclT/EatyGXH8d6wTUpqyCO9TG1e7GzbcdUYAq8Oy17OS/UnEuWjOqBTd2r3qwdo
9A272x5j811o1XSFYvaEb0ggCK2LDbyAGTkaHa8l83wdefWSvw3yj3i07dXOrdeJ
Bs1aj/i3+S5JAB5YGYvPqJjRXLVXv7fmPh0GH1PSb739TNlSKNqc4JdJRzsy8TYT
pfP8ImR4dtnI8ymod5Tp+sqIM+ZR7FknuT3asSu8yfNHQGGElT/w1pmhLQJHzdmN
kXPnZY/iErF2y79cYyLbooedL3vvGtnCfAmTZnLp4hiemuWJfNXA4Iz8nlchQ6RR
XDLyo4uQfWRLHsGQXngNlTtKJk1jqzFOQRqS0ELm7D2rkwUhuElh2GZOHnV5tJ+S
MGBTFXpyQNBu/KSWkE5G884Q1i7aosfBdHQZK6ChCcfLPnSa9Iy/TySZArvOORcw
Ii5It6UOOmYfgKo173QOJmUtnCkVcqGVk8q29ByapZhQ6PiBO/9HLJ5n3IQvNatW
hX15pfCgCKrG9rUzNxi2qYTvWu1m4M1QyhjNhcpOvFA47/bpqK5iiL+EBwNGj93t
VLBgySTNTahz2TnNMU8lPkHLl/De0zxyovSCKZciCe2R4fQJ8IWuFgtZpdB/MDtL
HFsuqv6YfZgO4XIqrl2yTf39QJTxvlCMqkPAT8EhE1a47+zThLhaUUG+DC5mktOn
FykHM8+ivFrpX2NsLAij3knGlDXk5lxkIn7FE4FU6zw7EEtmd9XyOx7cgwfKMAXb
It6gKx7CvyLTHvcT9kjuQcj2o6kIKeGmVr7cTb2LOX3rVx+bjhRFgN7noBEF5nDk
OuwGN8hWEtWT7qkI4/FpKiYmMYUGAXNwG8PsRW0DRH+IeJB1XushV51LZwDOCyif
rueFs5rGTTcoA2uzzSwb77j84b2WWSbI904ADuxTFniFWGFcZzFEeZswsqyFsv3x
u5+RXg79ZnrlZOHBcZ5cYDnW5K2v5qbDy2opp0wB2+cQSE2nyb8H5Jmel0P80195
OFAuarZEH2XZ7URJf6IJANaL48lOhJr21S3q41A1i/9yYSSR/kNfErEJrrGa052a
Upn/JIh4eKHLZoUQg+mIQ/f5iPLRPuRMAPs+oubQvxniEpu4oyArmsjVmaEi2s3p
O860+LYCa56BRe53pIqR1aXGQ7H7JwvG7EEGg948i9NyGxHz42LNSqZGPCvkTttT
xPHNr8fWReIaae4yM1cQzeKFGncZCL9VsJ8a4XPjNGU7TmNaJ9db/6WpV9iUzWGC
DjWkgKMRGtpkrhszuIVsLKU37xuNN1tXJOGGkaqiujQ1+nabukT0S7jt1tO0PuEm
SiABFw49+lqFyIGxSlVfEjBkVAMolCqDzEVGLzkENIEJmY1UOXQEpLuafkUlgwYZ
BNjF40a/vsMXS9XFKsb2GyikZH4WnVB+KZ5aw+Dh743oQe+iPc2XbZSx4yQhJZ77
2UTnIIezCUddliJDn1jc466Ga/Ej7QpBZb7QAX/UEPRfg2wxDiLt/gii6peCZpp2
rhwAgRKkECLZ0+oimYrsKvBZR6sUlveB+aiymorXbEdCIpB21OljlePmcmTt12WV
39sBTZYBtjwyyDgG8/QwB8nhELdYYhxSaVeHdzx2xXDD+20SIFUyuB27RUibJAky
z9x6if4zeNRNnMxAQJvFMuUHun6ACURnKyiF4GiKGonxYwJkiJKsHjc1bdna5UZW
GNpWgMle0/HTw/5y7E17GGQ1eC/rOjvrDiPOytLcfIJPu6Iv9hqhak6a4xwXI5gh
fJg4yvGj0wNJ+JAezNZRaQ9Fnj6nl+clhlr47yy44PL+9nUYdW1nyQwBlojAlfNf
1cT7XVm3fe2n5ncFSd4NHEhY5T4jjrCzfEAGYS4eGqPbZEpBTux7FMMRdQDNunwJ
G6Ua7RAFvrafI5VSFf2fl5plt1M8Pq52Scnkb3KXidY5VRI/xTRC/RTVzaccWJ9E
3bI9PmBMkUU7Pp9Sif+GsJ9m2+sHMOVRynzhU2P8IHNjo+Pu/aqsNkUxxyNshkUj
waTksYI5Ep4JUaPbPkkLf8PSHz7m9IW79xZfylLnlmzk3zQlLFWX4vBkzzYXlRqE
AMXAWvzFdZWpNabByL+hsqSbJ8gEg7REt9MdIGAU0Jwc+gxnOK4zD40WDTAU47nC
gfaqc8UXuyXZSY/JSxxo2hFMfht1El589mnxRUS7F0cYuXpxU06jr6WFxhwvpTRE
hC0OGtbdnfAbY2ep8MP9zlW2G1WvqC6MEmWRV2d116JfEKRoHgNIz2Mgsg/tyMQG
0dPoEedLoO2ie+Ni2DqOLUsYg5/ViyMZOFzXs38d7QFWjl8fgw/lIA2ONDS1H7+M
fOS3wx0Ytpimvq/EPFPemk4QeYBh9lTIS7hyeAv7mw1wcEYVFBsAkejVda5+VNG3
/V0PRWqhbymnKwzar0bCscXawM2GsMtpKhlxQZOqhO7MzpNr1RhSXShQXAHx9KFe
9QQTu7sCi/cpIwtRzuiRyqpzhR2jciNCobeqjUD0D/IDOh5nxJ8/7m0Qou10iIL0
idgwxz1i77SInDBcAMtJPkey0oPju/yM1lhAD2CF7wPxmcPEj+rm51qekAQNEMnS
LIzm3xz8/QuXjceK2xJ03FzXs5ibfnk+r/L4ULr2adNJEv1KNd1u9UQG5pX96qZp
dPzVLnX/7C6hjQXsG6/wWBxGDm/j8GiyWTEdAAHHmT4y6JTqbJAofRO07xCoGpoA
3oO7pcmO2FQSmQi3BkDxa7OLughsIZyo9UQgpbuxWJY/DMrZBW1MecN3QsQ/4C7r
WcAbLmxzf4O/TBSe8JCYKtZpjpJdq3XVbD8qguhQIOCoqqEj72m5elho4OGzf7IJ
vazl0kBjsolma4v7RcDmaezaQPvi4xGFcTlFlXmnXSsj4UPUHs2cSY22sVWocQBh
m0DNoaqTugOWtBfbTfZfU25Nnm0unK84ec40eCdUPcwsrHClJ17KVzk1qLZxDQHD
/LKredfucX/nZmNyn03fR7d0BiZtFqtwrwyQmePEqfya0AFCQ6M5uhK4SaJhXHxD
jCsrGd4Ol7tVf51wkxRV0HbdDggb9WtltbAUbFUyCxEBzuKRz3XpCjwTm1hs0Mb+
+b4AEYsLKEGJ87nvKzpowmKpmd7MLLtgUX0hzEbHuMLBnZkdtftycPLKtBL4CaZP
wqudGOuCWtx98lwVlQzd0rZW5OAQnoT2JZK83/Golo/AXtbKtdHnRQvE5QbkZBv3
Dkr3ZhYANp9c/m0l733TKxzqpto94zNhbR/u+DU1gzaaf6xyO/5KyPhe7kHVmshM
qMlka763XEWVLhDYbVDOgNtBB/W5YgSxKDvzCpJ2lLTw+4EjsqSfVl4Wp7Dt0uf2
4u2kfO/WT9is34lNaZuG8qUtn4knAxSYgyai4d537PNchYA0Bt/hnpkwBO5gWdON
Nb90aXJ7Z7o+rfRWzNm91JOc9x1GFwDtFZ6/h/OoY9jSgN7/HRBsjRJYOfw7OJyE
MuyEjFrnWZdh/7DPSCBJfljBRNcWOLFUzx6ORH0oyzUKWWwEMvSPNcp+l3XfoheA
gtJzDa1vQalzccTv70Z7AYBjFPTepP/LfNvxOQ6d2a3uyXmZiJavCtsXe9wxKAoo
1WGZ+xuSJ3xnZMkieoeZQa3MPfP2EdZS/vmh6NnGXTi5FKQzGJt15XIdf1p9wMMz
F8G90+xsO17zb+BS85K+CanJx8ggNKKZSdP9shodS0KQV2L5qu6KV2YX3Xbmab32
CsgTD+Tgc45NQDEID7y+V5ctgq6Xod8d79McAk9PXUv3WaheImtmx9o52LqY3dT3
StIJhP9czR2o/N6qI8YR4LB/J32Pj0pXxeqGu5FWbPezDobpobbfHEKjGaFKF8Sr
Ly1wJFuRI/jupykBq5x7lRUEOm+au30OnGQ3/IPy6WSvkIF/BGfDLxNURbUKJPOd
V0rtP5Tl7YiEBw1xW+C70k8qDsW1cNb5Y6NiaXx00oEeLLrvIePkF5Q+4cDBR1RT
zZjNN6DgwNZnJAROvvXyarOu0mDzzsV1J2mFLxm+4DtNIuAYzaFvU88ZWJUld/0Q
v4+SpUFQ/h2z3rKyX2GElWaZgQ8PeZfYDl79jjTX+BCkQud6na8p8S8XDoth8xHD
Wt4fdWjpSUPRNO0iuohxAEv5ngeL5t0+IsINgrM4cOwuAlIgDpR8rYwlTurfrqr9
zY+zeATvthMuesejdv2ALwK21UPPwZkiHd8IrRKIrAXLmeCy4WVtXtYEf/35OQh5
TnmXZQn9LSdVTtUQihKxqg9E/rl4pwBdrELQ/+fOUS5QXRtIjwCrJSoul6Csm6O0
B6qrSijEHWDcdHnYlO3bEKR6Om3DHZNiGR2lLaqnWQ8Ez7Fz5GHo42caBN2APsm9
mD0woE7b1zeJXh03ZFb9TfpGU3z8dXIFpRp1xe4Rwk4OtvBtL4QRcmQxA9zKpcbs
WuiScnvBXW1guzprdv1QO15xhQ+ycZERV/X11mvaaoheeoVXwxKml/pTg7zzvjfq
zN1Vxg522bsOcGFnAHkHGMq2I75HtUQvUtiCLCdqU1xcDAVy3Ub3H3vaSCnimM4d
kpVQxxz1Lk/viqJpBUF2gOagyHY2ve4tSslIIQfWUcfISJAoARM2LiUyubjJZbtK
TFUjZ+Y++sA9TfMeoLJH1JbdJpLRwZ18EMEFRIqw/+x7KRjZixb6sCAhVFDmzyEY
9AQ9SyMjrLatBpAxRxBPjauVndfvmLvxk08lwQJV1hucUDLjbxGqcxHgWda+AhoL
eLxMfVsHEtX68XGdedzu9XAzz+OxyWx/6PFmQXhHbUneFiKYTN5tIiF7gVAu8YZG
FZ0D5URdd1vaZZthfKuUVnU0Jc/MUmGxLb0xOo+pw3CUNy5VNQ6IBSaPFWKaGVJh
m2pyXgDam7993dLZhzPBlwqKodeTXtALqKEv6HvIM3wwYsUk+XfvLK1iZcCAG6xL
OdH/26IjpdYinb7De+/sxbYy6zdU53RhNe7OXkTqB/ctg3U2HPkkC5pSmGT0dWaj
NVX9WnElwLNFowFBjvXFCX4D14vkMDKsji+jQF+PdLIn+JJQHA/QG+NoaqBq5BuZ
9PeAIAD2Yj+cUFwZAZEoTwm2TvyryP4Ye0FYCuboHy6fBxyct1/dY8GtL1Jo1XV9
6trm1M7I50SHgCBZTM0f1tqHNq/mHC486dKfsDOgnmLfNVkGs8/sAZKbYmOy22JP
WlKKPISPbTKu21BwaZW+69xLDJC2Jub7bh8CQOG6E5pxfqibWKBp8EPnVzMx+BxF
+0jMaU4Mh/IGw4t5FwERp3JvYNzEW0VO8PKbEO0FtYUNEoqV7RZJnYkZhkECQlg2
Soc5i+1SLmoUpdQxpM/WamxRNfkg7luOVlQGjvmVH2Oe6IgTQXyCfTfU/5vqCELm
T84EpIWE3Ce+SoxMca05sLPVBmPIp1zpMa4Z/V03pqbwEwa1iE/YzhdVAkyTirGG
8VNtUWnElfCdahYclohen4rRLD0SZ8aYcUCoSVR20XSrvopjqnFZqS2TfGFeq8ei
/WywXj3xs9blUNP4NcaZ7LjRaIJKbSEe36Z9RHMXFLz9Wv6awXup4L3da22AUBxv
/kSVL5XKdwo5wZelJjNu5IX04vcFHndC+jHcdLJrArToKxlCifg5aV5jNxcrWHDn
iAd4NrKMLtKTbN7vf/qTEidz8uNGj+byP2YtBJCcm9H+RvIERXSfmwzyfOOYtHu2
vz6T0P+o0tO9r7UZ3kJLSIc6PeNzS7KrfEPbNUzTea1btA7lIbCgdvbXhmIlb/mw
HXbIuXZUKaN/6U8vKYg5TWKKqNzADY/xrPRxHFZbuieiRQYsodLPambJutD+AMkX
ek0SetACr1ZckZu6PIxg1AkL+60pwp+JlPemKOPFuS67p3pwTHSBmJH9mSR+vNN6
PZqztUK4p9a2SqXNqgI6J+gfGwHIk1F6Jl5Prt7LFQVwo1v54Fb+QOwV6MCB06BR
ihAb7Od1ADiyWzTa78olnQlRI42CFiLhfepWQ76D2/Gry9zk07Vg9P8B+GhHtmkE
1IA8Jt7F4uzZ3zbRE6yqH7oLw81E7RlMRNjJWNBPD1TTj+7JU7sFSl8EY1DVZGvy
4oom7Z/OG/IVYXiwStKqDS8clFH+B/YoUEjA3ZsH6aht3Ha1+O0xu9YFbaKdVCil
S7R5AvMa6+8CpcFz4+F3DxPfnJfo+HF86zWn6zQW90xMTlxYrI8iUCoYg8R6o0i5
22UYZYgGpitVq6uFXIwZYH8kHM5hqFKQYFK4/WjYnilf1uAOgd1kN5bMoC8NX3SM
BCqnYZ5kjwoibkwyWGVRfXdhIJu3/+l7/Hefko/bUIbVB74FEtceT5OLPPAWApCy
U6jgDRwb/sBkAFzDEiYWXJWjzihvZMkCMMKtMhZ9jQcGasv3ft1GLN0gIi1EJe1K
pUsucqKicrnDDFfQ1S90XduO/BrNU0xqSJdfz42FxGP1W6AwfiFdRkWPpNw+t+Hd
EnHSSc5FLhxIBPTrEPzk915M82HnFpa6/eiPH6+LmIVSRdNrvQBZwVnLuSrxFb5N
qrni5aS3vkIcVyV9qSoD5ZTd651HuyFsHe8x+L6v0KmHyJeBDpRQa+orC1KPSkEE
5jXYSmXniEn5NmSvJr/Z2imiLIWcPoX1c/FXhV3MUX8jQUsleWcAOVyN4yliymUB
iWDUjAI7GVF9Ei3kCIAuJQipXOw8myWjBVhR76MW5OqFov/Zwksddqv7d0w5SgG3
6/8yj7qTs1m7PqqsqYrjfSiAJhI4M35REAfzpQqHaKOxiVSMa5tqPBLRtRFL47c6
cnAQ8SE+Q6PN54gQgGt6AbGta2EgU3/WzvYJWg4ULgDcZzdXaKLB0RSS4kQPi9N0
r6pnDBcCoNXJx/VroSjxfKnOMGp+y94zPfH7PnDGJ7NZE0LhHw07KGyAKkw2Mmwa
fmgTZNIWfVkXjo7bgigcsnL1VLVpJYUrJAFdQ9Ohq4nROO3V6lRjkcCcq6+KqXg6
SKNZwBY9mWgKoFUxOAPPdrJmoXKcbWxMm4XvRjNHn1ltONPS5M3uq4ea5/FL4Yul
6ndEpaYtP29mKfmFfV36RSewzjct6RBXNThlcUqUf6j2IfJBmgpjMf/YGxcv+niN
lelvpQkva1QNSqNIE14VdbFkOGpT1rGOBnaZUYkfb6UOO8z/Zcv7LMDCqASa56ot
IjB4yzfOzmUAyKlJ6Gl+hxVc9N0KU5zyaP8HLzcfys8WDdzvvEKimbnbSxxZM5XV
VbI324i9OHdEk9jyMmRNuaMmaNjtlUFIxEGi4zAJP7M4YUqTVWhik39ftqrkkg9/
jLoAORoXXWi/K765/ZQeSsRtWmxSfD8OPjbFVlJxY3IijDwX98NRNex1HKOrDnBy
Bn1hnK5lgrxeKIjzCCtsAj5RBMxyNaBBpDAu+nxEUoiR9Vc2N7+7QV3JXNYgFIgA
J4q1oYg3esCCjrzeXh5YFCWq7eJpDY1wsA+eWq/wBjzh7m4qdrbPsfWZlLUpYJth
JgwOuxUlqeORH9lst1jqMJHxWizB91sT6B0lyP6kqre2L01eQ+VjdAAYcySRYPdM
WdTtUvRNsArPrcXxnnELicDI/SmvPmneXDwogLvz/LFHO7qxtpz+jqmypPsm3qM5
Je5gURulpqjWL6goXuAYariGAz4DSWGnOEVLb3umVthY039izSYMreyjGUgjYTx8
T/V481CyTCaRnwdQPpxkmP9vWsTd4I4e6VtwHN0mKZiHFxNMS5hkyWq3xBsLajAW
7d/4w6p9gL9VylCqGk75fvm6uxPCi4/EbZd2tCKyxAOFWrJM9QVnlgxhA6Lbnodr
8qgHbOTSQ7EPbFr0nvCX5fvG+RxOPWrDABmzLerBktus9zqM7c4khYIPkmTJ/mW9
WKYAkaibaf1NgcAGZSEhA8EhdbRAX0SQMph75T+GXnXdrovQVpAx0Z3Pjbh2upE+
qAns9t11rIvKrD03SHWf1+AJhrBCwMW7/AXRsOWp+tcCNpMqxx1/Sb7K75NkAGWR
/Zu+8KbjFApkKLpfwyMuzaNxUNrGTESyNP7+0Nb6uiiLeFB8KgzI4jSV3oDvNPeK
TpNA9C0OcL9UXt/ya3bRnNsk6U7zjJrLgT2zF0c0bIXa8sBEojVDE0Ee8CgeH/71
kBTS+Xg5nTMOmi2I0wL9ZSYcuWv2bCOXPydfc0gJHdPFnu72pCnkENQ3Lxezqa43
9PHyeNeyU2jOIrf1PcMcZ52Spp9mkgz5vIoUtxJ1XFHvX1H4jx0kxhQtjD2hp2Ab
4CZvf1joR+XuiaBblf9GlKwAXqxFPgNQHSNMcdqdx9lvMN7w5Rh9LXhwoqxNKYBR
1oW/dJUNWVaCoLsRsw8r+gHaSpWWFu9oAV/JtcSnQ4VJUK6EQc9RScPUKOylnEAQ
cxmhFqfh+JYN6Eg3MRsleKRxWOdKP/6nY3sNS3SLeKpU9DT6dCP1DuDspMVv5I1T
qhe2QZS1Pa9Xopn1YeBIlqzOsObctDgo8URN8xcGAOZDXw3APIq1gU/0UHwQLAD1
iwgX1qwSkS/gJ33yil/AYYfFwN3mKpdrxv7qBwHaH2hCDGFvH1Y0knmF/1sjD5ub
xlYQH+rH0Nwcjoiri1M2lN6XmmwstFMrQqcejFtUlNlKQx4z+cBQc6qa6estHHUP
akjr18jfk7BTyMC3cDQ3NPQ5Fyk0N3cex6HjqrpjJBdyqbBUw8lNGxH1ps8JCjv5
4RmMnQN2L5FULgw2znHLnVCX69cZQav/e+WiA0cRkCQ+KbDUnoH7AAcaqlmI1Bqy
+ek9tpZYQ66RvT27lhrVx8dA+SzrTpUk0oeHFwXPKvMuhgg4iXK5XETkTjId/XKc
b7oESk4lZA9f3snprttllStBNKXMuQrfRVh4w7rqBC/jGslSXzSJdwfgX2dJmXWr
HFKPydtiySZHto+kDp39jx1vYWyIvkTgzvisMl7d0a49cgJx6SZM83iRDpj+bcOL
Y2R5jB+MUyqvpZ11+Oywti7WFGXTNsND7JKar8IvJDAbK1MDaL3Wt38VOAaS37UX
0xkL1Kt7I3E2NF0wna7Xfd58IBFKnmkhxJ7HJRxvUE495ALvzLQJEHM0fN0LVUad
hJyHpYOZVG7+An5rXoeMCPkxYq9awoASjFV/klA8iwr5aNnJRDJ54RG4ruvCFA1A
JKeoK5wjuFc67sdUGDPq8U/U9Oot1oh5pulLHQhcTpO0cbdmGEmnFr9w4pD5k8y1
S/2wJpMmldVn/IRhQJ9DmcydQ3BtpOocnqGf8NfC0YmquC+86ZiCjYwyuYbdcOZU
+T5GrpeyfZTjAkz6vaQu9yS6JHLpQSuJgsmVJYH8MKX6ve/Dyx1Il3tNVrsTgfK5
U+p1MVmGfXdqFG5BLC6St/gjNOCO5PRRnLIuLq7prcDgr9AfSnxaUXO+YgSdkCoW
mAsLTYc8nFU+kqrxHHXpXjICxCs0hX57k1py0kH1q1EajNSvCEO2sBLB4rDf1DJM
suGRA89LGaG4tOFBHcrduVj3tq05rC9eRPPtkZUurbKoMRNBydCP9phiW/KDlHSr
W6C8oT80G9SkIZY4ksyt4l7nW2a2+zUdqu2HSMh44OYwMGo4J9ok4mv2xRQRUskT
nd6Kuplc1e7REoMXIv2lRsFwEj2QUYFa0SOEPFSZxC5uX2iyVxFHxbrYgutsfYN1
XFyZBkcrc7zkJzj/fBE1w/inj7tY6iXIoKbtXlUYVX1SQV0LTv3ooYkfDUyqUCtn
PXpOsUbj4wMUXEGULDAJTjjCR/SWPctvNo8ahg8GHVeQb3B6E5Fmj0xOkOMi9c4f
xwjm2Xg+/WASq8kxdu1Ipt8kOVWOsxyUdAaEPNSeRd5DYDPWDwrJpprgMIXLlJBy
2z46A3xjXhgWFt/Kfd2E3FZoBglcoGgQmc+4LGywnXCGH9cjiaXsxE89T6dNTQpP
siBGaP4FObFCUIhzBAOV3iUb9GHXpBBpwYPEnqTtr9D91sq3cOMcCFDBmlpfDawN
+ShO3Fe7ezkJDLlvrA8gzTghVv03FNLB5bnR11yXbB+M6sltJdT4kd1DIwMeYBgg
0iuKV+eZvUpVzeF4hy8x7sdAeiFuqqGaaIn+S1LJcR4PPYzLnS+8ehIdRZCcCHBh
p3Ozx6JwYONqRrMNK8YBsee5Qfi/eeh+snfLpeDnL4nUj5Iv3IEijY4olfGoWvcu
WmC2gjnjf8QUA/C+FQACZ4SFVNp93FXKRa25K4Cmzzg2png4vzb1YabivfHJMqtS
gA0i0LN25hJiiYd4qBuqJ3bjrFXCknEhkUa82RA9a8bu9JXFTaixtD1aY0ps1u7L
8zh1E7uZacMgXHAs+8qhirO2VLAZVf1ho9XjY9wx1Ko+09kDPk1m5hmyTMg5nJOW
f57jX2nYuaqvqDnZQj2yJTF6IkVWEDpDWvI7P+U81NddkBimziTjPvFLa+8Z/AG2
7htO08rohiuFpBQy1rXlrH+e1FnUqt9uVVSBD1RKTObGv3aJCAoroJwxrHFO7r2n
qWklsGoBCAGGqQhAuDSZPhKmpbJT+IKSLYhjKNCAc6IPf9gl0kk/F+d/YPJWc8Us
BPvfgc8uNm52lGp7pflUOgQ5IFPlwlP7t0QYa6u9M9qR69TZZ+Ieq2k2XYZsKhQs
3Qvq06NeyMogQ0uNvmhnp44DQwA7z9Jvm7CZmvbu73w6SKRUN1Kobq2VgRR560MD
12biYPwYTHUxX5hSrrs3QFm/fq/qgGtpBwHWoU9W4QBmqUyy21Fz7Jw8HOdDksU1
oPQI4bUN0+BAXw0b5gH1L8IPXnRA0vwUMcIR7mDJrEOyHg98yS014SjOYJfwTCZY
5i6oaLcuqzaJxKNhm7oIcWvDXMgUh/nwhuKgCQnyGsNKI5B3loAeRQPFOmmjTSoh
c6B5GVdjSLQcYIctBnCMeU0KThSpL3ZEWlubzJygrNLmIhxfmeTghHAJGfdU3Cxr
2KiUH2Vfj4L3Or23/XXwSCso+YKbLY6PMW0wDRQc4+GvDNtDdm8s3EXfyPNghzYF
WB+xFCcc0wqDYVIGfAbFnZAKGJWROHmT1F8L0QZL2PzXmxE+pM/dcU/P4OGOvh2g
y2PnfkBb/AwBaIbUgZrFf5uFHd9QMfXfd9qNcavmszEfWkOwzdxNR2q2m1ASKSe4
iEBE5GNGvHtQanXDsBLTohBA1L8cpEr03NYapwqZ6fdMHXik0MVa+aCVyR/WKn6n
1TZb5qHd8nig1J0ulzMZroI2Qh97oMqHL+RHHME1Ime44NiIoyyngnJolnoEPd+k
WAwDPCqmrvRz7wlJeOShxWZAn1ZPyIA93sLhnB0ZHzornqGRn+EOmM9b+uozN8ti
DT79Wzp4FLMAv5xwhmboL4D5IcNJSmf7FUxwESd8cMjKKOFZ3sVgH/XpuceTMNe0
b5AcDHA324SxUVycw85k5vSkTBfLS8XDoiL4EDU7oarLXQLrT3+NCfFCCj71+3D9
FJU1h8mF0du4AqHDFdME/cnJrsVVhhiFVkVOJTI57E5LOilLykQ1vhi+CHTN0que
LsQW7qa8dnkUog4oDzNRVUVYGCsX6zAFvKBLSr8XaPuKNqXDaHaD3j+PBYkKwBc8
lXOAx7jAP3SnnnMfG7c4sGTyo3Bnxd8SWQaq0AomNZmsmcKfqt/IHxEr+RC5t1he
keUrtNsxLfp036xb3AG7lmXRJmaCL3poELTWJVGsQDx/Tp7t5Wncvp6NbDgv+Bj0
BYdHCEj+GybhhqarzaIpEOG1GXhWT8GE5UxTaB4D9NDfyKQlUQsxBWFyT6ssf6bW
cwz8kLNMnW/Z1eN20MHUT1FDg5DEv0RP/IKqDyLRs6FGDZbrX5lKkYzxMvvM+eBa
mufF/Rj55BEom8Gt52pXQViBpl8If6kjEHsrughZ0HVxwHU062n9NzrntvkvbO+J
RQ27aA1PUIlCwc73Gu38LuKIxKDzWNzzgjPgKiSjWAPcNFICVWHoFYNNb3BLm64F
PE42OT0P3wznLoTff3u+G35EdSWpJS8Yt38EzqYaE60qxmjxzIvNkZPv9W8mtq6z
cOmKItYPTnmV5eOLUtRUhKTf9WiTPqeU0N2kPeiVQXR3M76ky0xwe9ozeWhnhwm9
37WDetiV0UI7l6vNE80wjvtpWirjf8ZhH4MUrDJ6g4j0AgHVeBenKn2xMqePakxS
xKThJ/wz4WPYk0J8BbfOVgli0jkSleR5jqv1NyRBOsNx/osrBxyghIUMZUGCJLZy
WjGi/hnXCPoqXLjO3Tn0FGMKTB74O+pXgJPNPbxQeFTfewscwioty5rRHMmeiZWQ
Q3YjCLL61zlMr/Tt3hGZNIi3r2HJ8Oj4FxlO14emCqPrP1prsH/+47T+cBv8Scd+
XyELNaJkV7INpNSbzEJROuCCGNJYr79tYdmfzJO7Sr0Z7dYxux+rt+ARR8pdGb7n
OkAgTcRagQT+FbB6+88JKfYDniP2xI3tEJUQzOzp8IIPvN1UM6IM6rbUWZ+eLyC/
R+qS1uyXerNMLoUS4CWxBe158MtYhTTExiA1c/zrOF2GC10rlWjPQyLXZ86yBUQq
k9A2UeUCsC19i5nGlqvN9Vy9BL396hn3COEH0D1RMQ66JJPZCOogdB+IuBNNiD2o
rhzph5ByWd1vWKat2lr1AnqvcGczrnXSrs1Xx8fFYgw7fjQhiuomz0Eacaz3dfSb
b2zbDjzVVo54FR1+4Y6n+Co9jnvTwCsybu7CpgtDP2MWUNtsrL335jU5HyUFnE5h
z6hcq431jGboXvXOpecoEuScfjLMcQlqTpCInnsUidBeY3qh61VRJkkMHgU5SJ0Q
QDLmQvy8j8/1dsyzGM5wTNqiz977MG37G/I8w8P9mco/YX/YufBi4XtSSxaHj9nZ
sKgmbgmttXDQtdac//sCoP8OuRjQKYqWHWqAVRwy6wOF7CpoxFhnD/9V9po9a6SO
BqX+1hABGB19cg6p+itx/XMEmQaEkWJ/1mFfXN6CwEJPkfs3gQEEssAXMZcO9FQh
0t9/r3FfCTqvjhfz4m2qygJWPzbWIEE/dMI8NScnUVbMKPKg9/TrbkXs4+9TlgL6
lqExTyFjnBTJtB8kM6N22Ka4bqxo58nVRbBxO2mVl4oE1MZaIIjJasSmnHCwd5W5
Pd4qjcv5uz2GCjsD+6pTr1JNixSeRP2H+B9J/Em9V9WM25B1/iwwWRt8R2Uz8Pk+
lwnNyt4oxa7jjF5BPGRAv9ZyuOj8FWyikegFu/3TieBw3Mop2U9C9+egAnUa7/zC
XbmiA9c/HLaxhxONY7jf9t5US+vnk6SW51lYTUgzcVcwz4xUGavQJHET/ObLUglt
oOYKLpUrgbSoK2nxVxPtgCj9/QfbImUMXwe/XK04SO4FlltRFRgTFfE2qDy5/0yZ
Ai04mrH6y6SXMu0ucE+VU3r68eucQFpoJ7n+nfubV21YGblnrZM8ugtLHoG2UyVE
GVWtxEEb0DWyrPNX8uswXbNADL0yfhluf0NKPSaho1XGesYFJZ1aN/KujdaecGEC
fZumzEcEvp92PvZKrhREN72ICWLUurV+uGu44fvZm9Y1FDd1Syqc4AhDKf0mQpG1
3JytAXhA7s9z6eCJmsZI5ARVDgwYPv5H6yKBSjpKbvAFUySk22fDN1I7KD3s3YQG
EwyVXXWlgwdts/FPJWl7iTgZvCwi7LiisPTnMhYJ4t3cJpgudzxFjV4SHU+nizSL
DI+ToqIJ0vRJKMr04vxCPJ/fVU1yr3mV3Fk2ZJ1rRTw7bCPminoei4PjT1vFo+Q2
h1JfPqixODgunCXqIzLpz4yvfAFL8BZA5egkT4zE433jq2QeDI3SvL8ifu8U2Jwm
3VIOeuYI83wx8AgMv8IkW9dab4jbzM74Ozm/MJJnSI0+3OqNBselz0D9mYrR5ipd
tyOG6ne39QK/n95YZaCLdd20KlNvJpfnodLrD1UTDaAEp8+XZekXZbJNsO2/LJjK
ujNkP5qAt33LWtZFMYOvx6Q/lolBgXHAlMVoyJe7SUNpZWpVfXnj/2T+Y2u8eWlS
U+SBlG+X+/WiwdLe+6HvPqFVYe/5JsHF1sjwoDF9pELHAc7UBl8uaoJgTeXAoeTa
uPYv8mDeC+Xl1sJL4GjPr1C3xDu+HbYQwVDTcjr0H1uQYN6WIQSI/RVO2GCZi56o
gVxa4GbYTYJsn1oQ1ftYr8AkeAuz1+ToE/dnvyKS6+0S899tjxUjXT9lN2e/elHK
APekyBxir5W9pVjIFhHqu0w79ysGohQlMvPeWOxS6saFnqWO8Ixa2CtcE7HWDoGZ
8tteuGW0co7tTXrpYDZboSIjFn0cWV4hcPWb7mFpV1nS0uB066MbSpzW9L18s9a/
c6KSbbmilovDw6qBb8NjytB1PyuOid2Ot0x11xZbto0SDZZyqAB0vC73aGyoOB0g
7hcILjz6Ne8Z5vBuZqPovR7rvdGPOo1o8hKs2lg+t/fyQS769xv8QsbfbutnvDZ1
HbGQs6BIuNvbIaFg8aYlGGYmarnbYtaPC/VQ3MGjs2sUV5diw4gTGyww0bwEouq+
j3r/3TBN5o1RaiC/ywQRXVl9TtvvsEY5D0EUtGzKP10eW1H8R9n2EGXo68rE+3/3
8sdNhCjVIDuX6md3JOaxJuIPZKSrHBSl8RbZekNizEd+DcUFyxf+D0DUyHhCDjVI
bt4x2UokkhlKBtZbXVmUibjmESrUIMsLCRpo1aMfHyrH8FUU/ubOVbqzLDicxgAE
zPDcPxq24SW69JiaXb8nac7WmUR8SSBb92w0Y/xoael+opzT0zvAUzk2+gbzd+Oa
SD1vpmrOKakE9lZbXB+rquKkic40X43o7rkOm/lv6B4bOsQNqd3nl4A+77jEbZuK
REJA1271rN0zUbOx0LJ2sl38ZgxoV1qukCVLdK3vcVWiD86/+8Xm7SBjWs5b/IRt
6jH+VhFP79w+4miOnd9tjgZDcY3lrpCJtOUiJX/B+o2CeBd+QfRJnsGqYTzyE1Mv
T2ihGgf09AabhhuYbvt78w4AQ3tsT5n1zju3MmnNNdAaTS2E6OdAv5Bpy7jFzqfA
J+a8POHE08VQxADKuMPlkFOFTSNXq2oW2F6sQOoGMNAAlCmX+Yzglas84bL9zBO3
cOdKc8fjDhpow9OgXYSlccbKvY+tg1yMkCQ87Bze9IP3OaqIzz4jkJSq0Omr1Ns3
VzJfgeb8TtaWAeE5j9bbQ27KRf/wVv1klx7pdiXr7fYGHw1NIQ8RBTAu9kYLcZGt
OcsbDGVplNiZC8GDcfxqMFJddX8aC49mD2H19cx9+ZdZqbipoGUFkQpNVEsDCsgd
CbPKNsavne3mz2Nr+2KVPZpH+UC6og8ohzh1APy4mAxOU5BrzmlLj8iCEeO/z5PY
LHmy8otQvR1kRc60CRNBHC3VFwduf1CsuP25lStDxxU0degt2u+cGRLdbN6IQI8p
dEkyiIOhAFtMYDqKCtlOLb7/+GxRWTUBx/4qc3iRWGnJ6Dv/EU7oLiZ8QiJtzCcl
R7y8egbcfzmW7+/jj4AQX14RGPvgBu0k/gLwPOU7aFit0G5namKwQEM07XT+WWut
B+7K8bGsiLPJLNv64oNJ3shYrzpJBbzY+0rqKt7BVFApcUKHLSkd32UPC1lydM9+
JOYQhTZI6ncQjDduwdd6iCyg+l5Dz3NNVPGwPSyY5wCPDGMHLWaWnmRrSDK0NGNA
KkU7M7y/oJ/bDO84QVp0Ub6AFCmQZ4f8H7kB2CXo4IRzeCIN5EY/vDkj0js6RsCI
hVnHFmgCobllwprMjNbjLzLfU+H8wOFPFscQAbXO0ovimFyPHY9azodi8TJ9DtNv
ni3QsLqrt3Ab3DyrC553BVdF7EEv6Om+zJD2a6Owyz0xg/j0Srq9Mr2yPge7k0Zl
SkYjRdHwI7B7HAcJozqb5OnIpSobGC4QOSa9v69wfPps6kh2fKDwGIJaqQJLG0Ol
gIx1kwEsOPoNpJ35fG1MmlR+zwkp6w1ru2DYkwt7iX+PaHz+IpX13lzdBKHsyDYq
cRf9pZOeLg8RP1lOQL5mo+BPYtDHnG32FavgW3jYfyFPKNXA+LoyrcpFxqyYB8Ny
0VpPYxWkQQzQnr+gy9u6vKdWCLEIfgXgc+8HrukhHqS4cUjY/7/1ij5f29pbxe48
VAk+N/3mdEvh6U56pi3T5LH2BsZSVxbeolvEa2VCEkoo6J+IJNFlldAEFYkBnAMc
ObJuo6S6PghNl+ac1yCulF5K4v5JEdNC7uwVQ6SfsHyWFphN+igYG7MNTl3S8vWP
81A20KdMEwCAZOpib7cGJV2N4wERNr/zoY7TMM6xnPkHhGND9+w9u3PcWTjlfg9n
2wN6NuHyOuJbcsMnoCW4W/6xfBLrLzSjKWBds9hjEdT/rK+jwK7jtNDOTtSbCeET
feAaQgXTQwF/kz33iCDbxLgDjIXmfeNwGJhQeATxzm+sCvdO8VC+5ybs0lxIh5VR
e/I0TN7iBhnK4CDsRj21KB/d8/7ykrfORLPUodKUMeYbkf6SXWo5uLx7AZMkO871
PkLImkwRJNplOENTmCtrKTzeJ4p/JkKtAIRxxjP4cCDXJS1lHstLPnL1vsifngHi
Vxqt92PPHTGIpKJ+X9skBoO3POu7G33Zz7uxJK9d1tSIUUtfrhoJGlyBVZYQu+t4
8iK5mbpYXcFmKsFajbIOQYqkNMCo7qZnsP0cHxlJxznCJfJJE/g0oqYzQWk3bI/3
k+ErQoHDGRZZ0mHEBgKOojB4yvWVu2nnJs6JScxv8ukmvnXZ9XYriVuxHn7cMAax
UGZH20LHOhxPhGwXiPQtg/+rqSpUeBaTXahoBYZcy5u2/k6lzdJmQVrwbHxFgThg
e+ngOBT6jb0h8EP4Eh0Kpd136HEEfmw0+0twBFFijPYDf+6XF6oqg7zpbFSbD9uc
v/Asdj/CYMkhX7yMneq5A7oaHUhDhpLx5zkOhkQIr8+FwasjDoKmcxoQTmL12pnf
HPLWbIq1OJiW07kkrDbrU1yqmEFiaJCjDd8j+hMaiuOkRNTPwIvLGZPXo66RwF1j
XfFwSPDZIjSLZwea95Yn4GI1wlV0MBjISjmsHDax7xwXbpLSw9XB30JGnJS2/Va0
7pfI6a9nJD5ooIVvEFC3DsO1mZ6b7mACCm4lbmgXyvT+4Jk8Inq4CvW5Fpvoeyaz
SO+yy4m7WbtjX52jggC68gHB1PcfpZDfBeMveB3QiDlzsMX0roQcIx7vRJFxQNE3
dHWoabtPte8o8gKW8UAO68WMHHBDs2jixtRBQoSippdjGvsz5Stu5C5l9DXR5H+O
pBq9sSrKCOJRhVELVzlRAVUBTKTcV51n7pOtRv4WUEjgavICuBiKgea+/sLMYArs
vhkdFRR74xcJpcQY4CEJVRzvMJjxp89D+SZAWf/gldk8vy+KjgFrh3RqkOMTsrbp
ATflrLdy2mw5f+tZfD4WiXOYayqVIs2AcI2GL/AvTtF64hVjis+KUBJR3zNs+y84
aSxQ6knpcEkwSE1EIkEIi9xHVr4W8+ceJN1e0gPud6J/6OY66mBicAa8xtx6iiXS
pTV2CrES+ZwpGf6v1eHSW/+p+/TzQXCU1kSHAfxSKdZOfJGhEEkFieHYLrNdOZ2y
XvUEUNQWE6G16r3YTwtx7XdUbqwPDZYRuus64bQBF4IsDvxwxPLofX9+lPCbvgKN
qT0nNoKNaa1RMs51/enf/gypMQrp5I9Vjp5VYjBsBgziFq++8EDgZT82/j9Fox3X
mQ+MHX58E+wt0ody8F5RMs/BCzRBTHlVgB7iQinieuZGud7qQVz3n6Q40slxK4Hw
GyGlrH1x2kkWfJephE7zOCGyTMX7KSRNgyOsmWoFtG4N3W1pQaqvcQk63PLrqyFY
Gb+o295dDGMZJWdaiVz3ccq3uQLiLi3/qES8pWtCDJIQEc+5hW6iesMnc4nSrjBN
bP4QXtEz4t/4TmXeN9PQXgjuohTw4VMgOf0dlORywUgS9nnVcOnMX+UGKJvBxJRS
bpfD2UVI8k7ihDgQ9VyIIL6m/EpcbJhmGq/dDBShUh8vDCb1JESbefmvQ2x/Y2Se
qOqxEM/oIQvz1EClrZfdICPX+VB2AKdLA3diZ6+LNX3CUBEyNOhkBS3WOZSYaci5
db3vA8NXpl8YzhuSS9gLEfDHjA5ISwMbtnX1h8lCtvb8adxcRphjK4ZtM/BIs2t1
xguZBwRNwNfMDlV6ySR4YYYclEFJOmSIFdNRykdjUnhmV43ycQmpWKoExZT5W5FB
9JsxYX06gCT1GYoQLSGWHpg8x1TBcvdoERBH86wVfhCWsDc7iKo0psRvfegGPgb4
NCuwVjx3+uy5uI5SfsJyvJlA53gupPx7lbWWU1bYeV4I1i1tZ17X0uJjq/aqCxZh
peOwik3nSyPN1/APaIQpts5RrNU0tQnsMrNrI0rzpX7gHbsuq8fjHmQZusLHA0yy
dlb1ntjsfSPfIZBEw7FnQUhh2GqW+RLMYN+myAtzWQ5ELmIXHv+yk8mMpmYOt3Q5
bGUpFgzJSY3PLlgdJf7G8MNZZGWKKD5GoFUxy2VNnw0WK9YyNsfF0/el4a428wnM
9iDC9VGgLX3dOGWp28IUs68FeoxsdVXSgkPq/2S+Jf0FmF3d7lyahkhep69FEojO
mIG/zJciUABf9H5a9U2PO1GGIhfVQ02YcTjJvVNpTMm8LwWRpfit6KW3l9Gkz2L9
BwIAyTVV9dRknSTVGtNhMPM/EsWA2p+HUkTC6NdjuB5Y/uygiOt8xHrh5me02k7C
XXwqnvgcZSDUXJGWoNvUEKbV1S8T2Gp1m2krkwUo6Cu+u3cCOagIz74DCYCBlUV/
Gl4tdo7ab4KoEW7uMfeNF6yEbMgtBpXQNhzZzjaUy0PysNQQhV3GYPLeHV8zQtHx
uuwjas7FgPLwGmseXBmkaZlVM+moydRMP8xt9vcGj8GYLTrYNeFSWvLg55XUBv7C
hBL3r9IIha18fQMbgJAn+jMmOtEBkwWF1EE+HAcQZ81/xZx52/Q2aXwwyRb5OAcw
pljLBd8tpj4hxlTl2FsEgjs30CXiNpgl3sITOGY/lna0yBud/5tbbUyP+NpfJINf
DjYbLZlhfRVLMpifq+PXCLZdVhs58GFsCB1L9egS+RAFR+3KSStiRJCYuUwVLeoe
hYeF0WTgRSKAAG7rEb8iloMBmUpGwRLzlyP0oQE7CNbu5qWL2dQTo7Kx9UqvShE4
o+vx691F9npmzD+6O30BqTKLSM6wwxDWv6rLQ/WCllOXFP/TtV7Kkv7GdO/it33p
z9ZiKZ6QIlJG7GQnJFuDbr+3z9i39ZVX7vPj+58C3w0FTQ6lkY7o3/QB0eyq6mAb
QcPXaTg+GEgdMUEKhzvQpWF/k0osCFsEMaDOPbgFAL2SChm6SnZ0ggQwzsji5meR
cll4kcGXD+8eS/28/hwhrsGr7mJTOFZkjFnjryTdsPA/bOZMOgy6x8gevcvL9cR5
m3/ND4r6sYPJU+3h6aQ/Yclw2PxGynNXUfc/K/Hoatwly3zdGjUZblQOURFtaaWC
lt32XxctoPRhfVtRD1kGtTKiP4DEWW6gXdBHPzmXB+e1SrVEVt/SmWY4pyx6XzCA
wI8xJqY3yy3NW18ZTWjpdAqmQSE0XYXZL5C1g69kVC6RAnwlJmLKP8Nc306chTD+
L0mwxrKjJKP/UnRMDwP8ztvPMcro4Sp03vdIU/HP80Z50fQhMAXdHYiXkOsVP8PO
Jxebbn94HMEvqsQRWH3bsJQ11Qkm2iKLcWWlJqQ5xQgg+ezpo33JikX9d3HnrqvR
x7geKCuDHetPnhxbL93EdwkKh2mM1oaBmTau7kSQaSNrznWHbef6v8ndXna+VlSr
fAROiiNZcedibFgw9G7szkaCy+j0tQwwY7NjiFlxP3uQ5c4fJOvC2doxiXsLQk1c
GxOCoc0FVGw89SwzqiVYSEkD5Ro1vHFeReh+JOs+nwWBBHbjJfJkIKXcApctTWdj
iqwB5JkInaFQnncL5Js5mukczYOibHo37MTBo8n3Cl1OaZpqBHsxe8Lkp21Mf75r
LT+WoQBknX8z362AHJJ1s91HKbWkk0tcn+xRPGZLWtibhYH8wkPardIjWByK2VOv
i3Epq1dxO+53ewb0Q680E2dktZ+D89ptLrXv71nO3iSXF0I3oicReJXDfekJm+6w
njmeZJ/iaGf98Iq4J7WIqIbqUa+KbDoAVdGvHXxYL8ciFrRETiGnMPDoNgKqDhN5
jumy+0ej+CBoiFSY7M16R8U69XN1aP+lySMbQpA6ssDxi8zjy9OCj8W+ilvGsvAj
m6Xoerj6dE6VlhN+ymLRZ+e+P7+kJnW842ZloOneId23ih0LZioE0vq9Av6BkuDE
yoREaVWuom7DbIaCZ0yPK6JQu7J/r0pVSJ92mxwplmDYoKm13O33jiqqCgrgtD1v
IHDzboShzPcsA9a+T+EAvgrjW2tPFEufzTxN8q9TAGkg0TSMzRbUPHB7d+ux6xSH
7DKr/NraSf1kiIBrUEcysQpyR9B55baeBi71fa6WhQh+GFIhWlL0JRpi7FU8dr4A
c/W38pGdJ5J70o17emuN67axp00IFBdlNEw6gX6EauP5aU3IFtRA+U7WuzAk403o
+r5wg3FSH6aPeYmpVDfSW7kJO9kc2GGRPy7pPAmDQe+67x3Xpzld/elStvk9XY+s
PxJP/5Nee2rcYzWYHKXYm5gF6dQ3Cl2HB+tUfDCv586SsPO1k7lsqrw1RwaAQmZW
gcIgLTbHyIx4GxRvlEgxudXcYfQ7jQhgoUDnEP/fxUsdqj7O6gM2yWjGk08wux4m
uhB9fXhHl0WHKgdpgMaM0q8uyq6KP1N+t+IwL7vklDWSC0/Lydy8PwW7DHn4To6s
rPxt7ZmS7IGMKpgrHySQ+JDLUTG7ChUiPnu7W5Mps+yZXOlBPzo8JAuiwuKqXvVi
8YX49p/K7DX4vaV8Z3qH1Uyqxnz9kEZUDnnNIaNHwTYTKnVg66dZAxZFB8kXwkHH
20WsscSD75NyuCzw3I5oeERNkhetzPSxi4j+qfcMd3/YGV1E2aKF2bGf8rL4u91A
zbdgrymsFAqkFPgSBmdX48toEVbLKWLYHOxluMKqKWjGbH9+8nTHIrknxHhY6BLA
xuHph0grqcZFSTI6TWXbsjNFnF266S1GSMDzDuYgpD0VdtlGSXZrEn29eqFM07fY
Im3HgDfi71W4UzXy5IEFZjqufmLX4hzW6rDeGaEWPmhg/7UGEW/4b7sub+aU3piq
a4PJOB4EFBA8KCyalM9ou/Fk+E8ur+lzLfVwYXwbFhTj1SlFhzT8H6izRf/y/Qel
OrKWaBS1YUeH6pfyBvFz6iQQK41XYI3dI4jeFZV15b0Ta+jYTYfIsR/sLRsg9tEq
dnpY48qEgJDg97ejk6L9iR5UHjuV4UPfVT0FER9QxhimMJw0UYR0L4WaRz9GOY/T
FyFPASfM9XtKrZQfbjEVTr61dXJmlnyCwJGzKFE84mhemwgmoiPsabfn1QZ8YzM0
uJJFr/jPWmNVKCNdx4YryYXl5itKPwwM5hVoWoPk0z4O12+96iwX6k4apkk25vXP
uzhvdYyFctcrcoZsD5AobXsfQ1o2ShCdST5E8yOsDNHYoar5Nr/UIc8Vz5QrXJ6B
Bd17nDAr/pxnyhLw/bGyHMRI/DETI3M7eqODIGrSfXgNWBa8QBfPSaVhbR3WnoZM
CE1xG69QHANJ0X397w41j8VGQfVH37B9WFsKRrStPFL6hhttkyapHHsJkV0FW6gc
tv+Ik+NKMuvZbQ8K4j7XdbjdO5Aej6OykoqX3uBuh7Owuyfh3571nuQzEcTkysqj
FHKri5kIlMx//kizNqnujEySSOSNux1sWKom9RWjaBrOK3O+xnd5IwGukT6pashn
cgr2fz2YNK0AdO14XNNZmZbe6z4j0wJ/R/eu0xZKZUe07BDKpaK45umdkU/HJCCj
WsqQoKTI+8qGaZP9pR9vyVmbjloJjpsqPEKsP03IR/fvskk7ls2Pz1BUsGVtcdKE
VFsRKx4Ass7DlcPP2VhkG/YNfU8sn1QhJMjEni9z4oYs6M0Kus32eFVSIcR9Hzkn
LbFOY54cfdNdayGgL9PbO4tO81otKtzy71drXErJ1sN//jjAQvVRzDWvaO3fGB5p
QQM9DZHkmP8KzZX97w5mqF4tODlBtDQaTb2BMzDD0U8cXdjYxr7JDutMyTIwoeJ1
O1f8nxwSNJWsgp/xSeLg2GMdiMw/mB9HpfHP/RxEXS9QmejWzYiy/EHGb51br7K8
R+ANiSSbFyNcjXk5Ytg1ESSgLAztudduZvAQ5BhzIEi7iopc4GOilY2d1Axethrb
YnAMFcaR1vI7IzKHg7De0EPJP8v7Onx2ZyBWTC3e51s7bMLfvwUGu9J7N1FmGa+v
pKgMrlNmS7Gmd9GfAHiKIaAcZCW0QUgGKYZkMkLviyc6IiOcwubCKyZJ7X/JYHey
cT2MYXLLZo9kXNliOH2yUXLEgrQe7DMVMQIY2g2DAoUIzN8uDHmfPB3lHB+wr0EF
VpW2TsByD1oqAZke2Scp/JSR5j7yncenvDtB6HPZVkPJjguqcy4De/xWhxhmMljm
4h1GSwj0Q5UO1LFQDot4BtYCaDkxH/XqdlropC2T+Tupv+Sg30fgwD0ftY2XrMF/
hb5soP6ChqYSyTBuvprCBMxGTWXh/QsBO48XYRyCIc0h7bHskfsN2JKBZPPorKS2
dNXL1c8btofGMONS9nyN8CbKhvkMzkqwBUq8NDy0ZhkKb6EFnPm/OgyTSJt2aFdk
52ASPYF+jUjHm8lwqyRR/iK33gtB78cVwLcIQ3v3GSMoSPZxG/TzJ1z2tQgXj4xp
XQYO1TG4MuWsCqcfFy0N/342PG+73KFYcVAJ137GRkJGhR91WFJQZzBN2XVuWzoY
LuT+msKwlUdVa++gBaAi3GFADfQkMUe6gvMuDphLjZnByx4XOMJdot6iq1oCII9W
6Od2J9lOHgSBsV0MLKvu9EmHvVRiN1s3k14N1OKyyQZsmP2NfisnY1C7COwotSLB
J15niUw0/aF7eAA4JCQnCZaea9yc9hj0p+RzqsQaTSn9wSziBpx3IfQExNS9PM4b
Bk5q4G3n3xkTLpuh0WR00CBelIejXzf1fFz5LBDBh4MKF9wmZi6TmPNbmjcRgZ1W
ez5/5GC5uSZj/4nvVYgDSk7VV8nZjjY70P7rMxtxz/ceOml5iRemdMsj96IOt1xx
YCsFceR3tfh/v0jgNgcwreWwMA9RhbdHDGsseH1tA38I9kNAX6ROkFif/vWdgLWv
J0RyQ26SMSpi/ffB9RBmIQIgzQ0dA0tmMtyyNIOd+Ina6xEsRB5YgfYrsyXLTzgf
emjnMBP+sAykLM1q1BpC7NTX7TgmrURPYWo4VHRJl38wDtdtjAxraF2Zn0rtfbCW
MAWIX6ONfKCTgeHfW99FQUKiDP8tZmo6DNT7hHFwD9yIuKAClguhO0/S02pg+pJf
CzTv+rktbtSM6xXrF/HK6DCZis8lEQjmdOZTMm8hdIrnOPxs4ZNMLOSKuQzCMTHK
rrFVI4ou2hGEsCi5VJYIbgeQADDhSl+1Sq4rkenMju3hE40X5pk4de904D45kioF
AjkqaHelsH2wtXcbjSMv00MwaqsC8TvxHv5rFvKZ79jV7HpQOBbR3DwXq6tBAIT0
O0h851o9eqv3hLfZRrjUU5Wx9F2N5rPI0hvmHhQABBXtoFfAuswJZbq7UYkl4Fn4
ldyHiJ/sjCHCaOrAeaAm9Ey1hogU01hNUpNCZF39SbMWlb5GaopqP+J5288ZNHEE
hIa3A0hkioNXCsEXiX/Z147y1GCMksYnGgZT40OOaqwVNHQ249GUUhnra64Y+hbl
+8QUX415/DmbGk4iACKGO54yu8EDOI1d1vwr3jnit6YXETzUWz4cNnVr5nh6Hw6y
/MiqwWXyssPS7g7PStBk/TaLIX+D/BN76GejOIpT/Tesngw7GPjz69aTjFzrlK/D
2DsFEuRsSN89GuNOIQ+mP8suedqfd9wjQ0q+lCGBojaWssnwpjp57YD/D5mRIkPQ
CwS3uCVvCgma+EWry20wnmlix3Ar/NGHusPe0BmeNN0O2RnFvNnKCgYc0CC4pGem
cSs9+CwF49RntAYK0YGGEOWAoIPGAbkKK5j95B7EJq6aFsgPb8u8iWsgf3hQ+Lmt
aqYUd8Z433lcvY0hj0VfUsN5VKDro7gAIeeaxjsHV/3Lx9XqtNnvazE9PunmuePV
ENCKJ0Mvb8NGbjD7Mag70/cQTUGHxMPrNtPbszcbdc7LzOEklkPhzkX9H2xEtzRi
Jm6cciZ8LUxsO5Z/aMq1YsZ9SXyvLcj9nx0hRSfg5Ntt0UnJoCrofeGS82N7rpZe
vjuttMFB1WkUGm0bjZyJLAkhBIQKUArjuFMJ45YAgfH6qmggJnAOoUs8GPNChY2h
Gq0EMRyTP4+RRRHXV3NOoDp+4Yh8q+7U5T3h6sK/uWIpjPpEw7fmMFJIzUL8+A17
kYItYeFsxefUreLhwRYsWt40khkuAnVAaP0suBHuLTmNyHbTUXBYUKAcDd0AK7/G
8gdFf2FSwqYc0q9aD6w/fKJeP6hTLwRY8f/W3rcGx2J6eZkOW9JHnoLT6Xtdz/5Q
UIaGVCNmTj7A6bHtB2huVQVGPViUaJjnf7W3jXKTy7joOd+1LTTXl7FbbxcjLz40
PqG0Cxsw5N+J0z0vkg2/wRf3+10BHtLHDgIoAuChRLvJqOEN4ToRljd1nMBEPvtX
W8zBiM/9lPCo7mdpJYzycYQoUulQTrLYe3mW6suVumfljE6Ei2WVaEUGffh7sE4R
rdrVgl3pBj+OwfDbUFFi6GK4iBNIXqwz85ChT+5dZrxjkx0jnN+Kqu/Lc3d1zUBL
V+JqEO7zgzMmfMn3VVpMRMIbUoMHuVoJa1tL9vRR7tn14+JB+uo/H29vQEspPwk9
iqhTC2MGPDnqQA5InwMqE1lqHLw8TbLv8P1yfEM1H6+iX6ns6d9ljvk5O4qqO+Sp
lCigdQyFJz5fy6SfimvWVx4ftaSk7H2SWhiEa2TsIsZw+Vw1JYSY9wUJIR1EK8kD
58ocnd9ZKnHlq+L62FkIQQxRZQ0bnDvK1cpCzCP/Kaip4289UEN7CogegxeLdrdR
FubhSvH95VVrtlBhZECwkGtnjmIMtI1tjK23ypV6drvChhCVmlNUp8BEL4fFlJ+y
IQyfK1zKQ5GH8HcDYglS/PW5AXegA/JDlWxTuFq0ZfQI1DqpQcL/uDzR9yvbQykv
KDvYlPTgotKlE3SZZ8cxTOcODRNMe0ggESnNeN45YzqiSUolEjlTQGG4OTSBtTGK
jE1eLCN57PaG/Tn41thKAgFjV9XPqhSQOcmQ6lb7MA25fvxG1OYKFbGk4t56h9T9
KZRyDYuyBTMQ01nC3nVIrnByGPIAIvbhzH+LjtCff4e5z71dzp+zBViIf+cySr/B
SdmYZ6ZtH0374KbW6w61ivEotISnUQe/kmknMTwVIuYr/WKOQIdmyU7kFrHmLfam
99Z9FPKP1tcfoIoEMKQWhudkojE20n36WLCLFjWSGWLQfnJKtPunVjEWPTGOXCBd
MwuQ3iNeG1mZyAg6+0G7uFrP0uPW13ThTbyi4KbgUtwMK1qgHAe0LuMf8f9QWd5v
EOhfY07OInFHR4xclDvF9bBjzBB30svkvpEkZy+O2Ayj//TQv7bY1rJcSMFwJp+/
LwhJD8Acf7gY7TRsI/TMwiesYkm6uyWSZvfLp/1QGfl49R82jWu5NrHCH98hPWhG
1DlJGkSCWUhMro9FrgTFoBcvSzg3tzYaEK7wYeLgCRPWJT3uxyeMqvY6jdc6sFQB
DuFbdvJYS0s4Sx4Q1/TK1oDdaiqwjI2MmFGzI1JpM4+Pdw+VxgDZzYRNuEMucOWE
TvkmKuSyl+qVGDufLqFPABOxIhpTBBtAOoizu1PzPOIVAczvrcprNXsyh/dWt65l
NmFWSaGdTEeISWVfgwVGyFkQPeZPmKQbEYOnP01mgGn19eTw06rmmhC7pj9l+HW+
TJuduj3w4KZfbRBRBqXoh+/RBNsvEGKyyFr40pXL1UWhBRsamVWqe5fxubJEDdYx
IMviMYMLKi2aBpOucfthxFl6GonEB4so6sDxatOswD0KgwhgH7MgV0t2PmXE/+YM
ylHksxEJnyQ36sjcFLSEEvIcHP/jT5baMNkesNqqsJ7CqFzH3aTC67/JlZc7z9H4
3QgCEFh+PVRox2N+25y8aK0K5io2c2qFZgUYqc0jk9qRR3XwQNobp/fG61AcdvdW
HSMC7WWzRRs36rcNSlbXKgPny9itsQjVXLTtznjP7XgN1KJstyp24ILW/UUvZOOz
c27SreA1VoZNuyPexXL9+9frq/qg3tLyv1HZBvoW9cd3DXnSRmvBTygIAhAoueZY
J2A+BO2xVN6IGO1PYtE9u20WyuZl5pmglJD2IaA43fKSOOtDUo6bR5fjNRzoOAG6
9wfepS/MSz6MZG03nHyrY/t4Iadk4ngdVVuo0EAhPGlo7WQZXZ2jhlClGRHlRA0F
o1vNZMarLFyzmz4ljqReYZ3fWXqOC9kO6tE/WqZ7c/xzGxHoyK/YlHqCj23y2rIu
zLSsjEBN6P+obpvUNZI8jDRA1mJbi2Nnv8cykPa19Zzy5jnqkzfsUnx7WltIxJqg
SIIZ4dy5XQ2Ea+KFKrpkQEltGnQFLup4QJX5ZonqTqqqjJvRA80/6klWw84fzs/W
jSPoX4Fh5Ec/JIRrHFrSI2kFCoXLrGi1hqzNLhnzuH0h7yFvzyB+FmATYw2dCnBj
FR0Cn7LqMCmSsfG/65jfAPeef9oBQEBaQWBisnkY/sb2ZqHE/rQeeAjlUKOSJgpD
mrMV6TfN4VdrNG6WJM/qTp0ZQHOKao3nO/Szl4yntqxoNiE30Odl/QHx1igdOimB
CJX19VDOZzDZHoX6MWruMuKbUZESLscngUjo1QdhB8Vzc8eQNTseB71uSYq+tETn
KYPmVkQ8PbpLamIwGwJSZzGlxYBzOv63xuuC5r6tE6idkwyByoMMqMvrmx4vix8v
o7mosTrWsleczJmlsEQ3MvjMc9N03KNUXWsSMqghIjJE31y27JHHyKMnQGwCGtsN
7Dz2ODWHZhSWDglzyIiQBJ7eWNLxRmn/IJw7eHUGwb3RlLL2o5BptXak+mP5nAfV
8KjMbdMgctqAkcBZ0JSz8OT1yyTTKU6w3ZFO9WxnzphMaG65iixp1GIxIY7pyJq7
T033JtRLaVmNQXRfJX3O8udBZXvLpkwrQ8f9QJXi3LE88SB8+LkAbKGPm722nA85
a18wNm06aRv4p34eGEtu8XisKuF9wSY5cgxKBGbmxwofvZ4qLXzToNuuL5Dz0Oma
kJmaLvoIjl3Wk0qZDNPPTjhr5k+JITCEY9KFy8WSi5uKVKmdYwEqCXwPXIMcy+Z3
6MFAWrn7EhRe9uXuXQpGW0pR2mk6K+2r1+5/15aEKti49KxFG30qPdRRBDjzjQrV
yDeZEp2TFW/9M+QLKjQFJNCLXCIZPQ/7eQfdOpF4MC4uTeyuOe4dvjro+KtcgmnY
ggmi6sC2vqaHFchvp1d92V0WHgcXU/HyfellfOwspkUtCuSJm5mm+HQw3o/J3hDw
d/HUcusoce1R40r92k+5ZgrLlujrBdt7gFzWPmb7urMv3wxpRRfjsj2gTaNtfgwf
Lr8NlBK7lLSYZ5SI11AdbbL7s/JwzrXMPPGwUYpRzKz29Sxt50sygDYy77jFuG9r
rHUszMoIrB4wdWUNexrRH1A+/v0ISacOncwTSzDuhByEOurRfLwOUKyNfZncTOCU
1XvZc8xGU58qIJ6sp818niBt8OloPISHYRVqzX8lf++pqdweAkz3tOPouDinzcpJ
x7RblfAPdfl73+82jvJA9W+MYHL4RihABPKllAy1IwGVyyodrXBKgK5k0lvn4APq
asjKAA2ed3OxjQX3Wu65e9KkXK+pk3laZnboELKX+8qpNtCSkv+VpDMN09X7wArb
x4iAe+m/4cl4h7lIb8FVYSXJIVLMySlujJPlGW/gFgLhongTlAJeKhMXcTcqZu3K
nHgkHBYYqBjdE0IdVp+TVBPTnY+b/Fd6RadQ41qSQDDCSgAIkirKzPEC3EVZ/tUa
yrvAsTQtd7634NKLa3HwAutFpYGMoE3dMI2VCqW+VrMYv5xA5cX6zqd6GtD9m8eS
eFfe+lhZAHz8f//s+2QnGdqqNf75uSThY9D/X8O98WcS1faMC2XOVrcQXwXvD216
AFiSaqxK2p+iczhRqyPafk8C8e81jEbm1MzM74nACM5CJ3rHom0kl4CHBLOCOoDn
X9ZHS/OtXkb5hETjm11Lid3WXncAYwtJoQotqXQ4okbtsIGplwbN4dmdgMSbpg80
VvQxu1x+LQc2E9Vbqsfo9hCx8OrZCuEFh+goDOUiw577yxpeYyjMmGTT+ZHh33HY
mMD0NV8xXhatPptpV8aCFgybUcPCYQ1vRTzj5mI6xgZl9Y3bBNcnHddgZ2G3n12k
IcUiRH6RGwHs50K/YlWh39ChIc8NkGXbGrjDQA4u6SvTr/OpzjROkQNC1M1PC/MO
KLN72RASz6+mBeIecYJPgB4KXDpzDe2KZSQwP9CQ5fXmSpNjfQXxv+DbVopG7M80
sNN2mQCPEyu5C3fHPK04FWWvzT6GA+bLFVcP2xiiz6hjcsGHzYUreaJVBwKkbkY8
gDTfoTpf+mMLcKvmUxb8/TdpATqSzHfZDNJ9qQASY+mk8msOkwwKytYTPD4ckaDr
5gVrleh7zTz9LhiVWm1slQ3tk3CgtiZamPf2Oqbol3uZTE2EVpQmrBc+lfmoTWt3
AboBt+gyKnR3m7ujnqVpNgs/BLbbA4jsrKfyJ7gvRqeKUClPft+W72ijcp0/TqUC
+ARi4dz0MWeOgB24vo94tQ/oFstX/EreHxMFWo4vSQNk/PJAGLf9NeQxfiYvRm8K
CKn2huo9CKWWPN6FPNFgo/eL5oAlr1vAftMqQSLqopvMZIvNBwwaqEFdFJNcKMMB
IPwzNamspDZDni2d2ftwgg3wXINF+boMkQGBc5dVBkYmJRFA5UmrY0TYuwpDm206
663v5mvxytqH+DAPu74KhMfu7E2p47IRfe9QnDe5cXa5S/ZKefb3b1ZWunzZgxa8
Hk8pH5rxKiTXpoD1DWRtBg9skelB0HmP708YQ0P3Wk9+LQ0Yy1W1Nt10CK6sdTd/
nUp/TLfzQOY6HoxeRBYqnGOz0jarKsWq3v1w5rQaOr9oxdsm4Z2IH5xwXUfoI4mg
IqZrly5zqF2yeEQxt+VyoelHava8FuEdadQkckkLBbQB16MqeM/4pu2QzASF0pzP
VLO/uWQD8xrDfUU9nqMhyQCPU1vTA17v+DXlTiERUEKoscP07vOrrG6JB5wJ3Sby
rIWt/dMdomoRnaRGLh0Su58Xyq3XNOZ+YrfDztRyoHHehAu2At8OnYWJQaaLxU6/
44jvwm52T7Trg+egoU6siO2tMWGtbegNgIgr8bPEDdUDRBvbgSLhbMiZEOnDfFPD
TsymxR2iw152dnEMf/xB+RJBatRh3iPwe560EB0i6JjC0NVe0joOJkVhXc3W+hVR
g2qdxbWXVCbuvNg1BzZuaiVBAOQndn0DErs9Y8t3QctnwrVDHytnF87H+dNzRd+7
O4jU+kWeJ7p4L6+aPw9Bd+VHWoPVxGIvhp6w+qaA7x6ZRUy9j3nlFSmtRoIzA+b4
LG3lg8SsA3WjM2mMUF8f1tkO/uhvCCvfTnSc0cXGKeofyWq4QYQ9IRu/h5tdBB0H
/WxusfOftweGffmijcvL9To+20bhtDo7kuY3yCcEnYVDmv7ZrpuTEAz58t9lr4fb
wktZANJ0mwpy4suerlOgCQjB0VhWH5SXDIrUL/X/5CMjpvP2zyL93rPilvvpl5W0
a7PBw07IQNOjMNDEvJqytrNEQeRG4xNVPYtE0todgxHpl+AbsgR24JoBaaa7/UXN
7gCiXbEunQL9MIYaPmSFNLPRwMkcGLYcN4SMQXFSqzs+runt4fyk9PepgEp5CNYF
u9d2nuIzYfxHWankkKM1qmjR41GSKUrCz3P+YMFAvst0OaEVPSQ6UWEZpn1FCJ97
3k3aDhvP7NenOTie+qN5S5m4nZrS0CJRuEDHGKEUvV8w714zjZGCSMneArOrkKIb
0BwOcrcQjZNYFe62SMSc/jlowp0MS7GgP1bZy3b6NFMkGybTTDYKwZcT+s8bSi7l
JINMBxUeGPx+RJFTtpCOSF9NzFW+/JkIuOwspmnXC5G0dfi6ZGDGpA0fmdYPyIcG
DT4xNBVB8fethS1WbMxh8w+37ieitAqFc59X/6SByuft77A7RxMEu7O2ntyZa2gf
UXQukd6fLqhAJTzw+EJSDZ3nkxQi7Z92DMhdIhcRa6qs5We6NLhNdcGa6FC8kgPE
8wCDvrYkmiW4TU9uqZqkJFolzemE2lg0EM2x63gJMO5JJAmuvfu7oyluuaPOGWWA
Fux3ABe9AvOQMdY6G69JBsNBQEvJ7YvBS33GkaWti1XVbSyFFwzevk4VQOwompS8
jSa9QQq5XubWv2XuKmsiqcVkm0boFfnzLdYbLZWk6MvHgQLJTF2xHfgKxQSubnui
ORkfxYjOIuFF0cnSCu97VGHFJXQV17s+IUwOp85dn+CQxVJCEjhN0KpGev2KRPQJ
lUpmj8C0+7m208fklyIBBMix3xZBIMDZTolBTQLOwxX+4VJKMSDkSmolKEprxi5g
YUQhiKKkUaZWbgLIOhSQv2qtf8KNJpvAO3swoURyDIfPpJlo20CyZdxgxzvIibJm
KCA3mqPOuOxiVgx0PMwsdKzRvylskiOoqwKfGR7Nn4OLoXF7Pl4e4gqghq8aYTJn
PVXL9hRI67fnFVtz9bos2idygYCaCpUjFAlT3ukVFSn3FwPQS0YrvMuGO94llLEg
Roddt4y/OrS0j+n2+kU8zTTUQ2lKZ7raVbpONj/00VZ2EmbbZ2T8Qx+12nXrhbbg
QroRhaQnOOzfApjfIdh32C24E0o7pfu1zrzdn/RcSYq/AT5a+qRPrQFHePWbHj68
zFwsdVuiIiHXBOHrXkHAGQXbELmG4TATlPmv5gtcR+EUx/e2OIfcgldivVPb5oH3
6stbxYBL1ETQkN+PlNI9IBH8C/J7OM0WsBJdo8GgDYgryaIJj4CowiFxk/UuqfVv
ldksuxON3ykSaesq3ijfNTUP9D0ae2e9DzLmkYTruevnvlbro7A8c4iPQ32kwGQJ
enStT88y1LkK415eM+6BMjd6EoIVslqQtj/CYrcwAA3OKwMrzF580edRxPy9lMQz
pJgdZyAq5zYgVAhzhwrsjF6GVAY0z/0lpM71oCNqT+Q0KfGvmhTgqNR+E1dO5gyC
L+ZoBDgR4cppNB9xYeRX7Yb1r49UdfpDUqVh2Vcy+wuHfNEaI1Nc3Het2W8kOJDy
qGqwmThOhYDKNigwdn3jGeXbfGONDOqzvZcoAH8046n5Q3nEL3glEK3HRDZ3SId3
8cdH1Vhpfk7bH3CSEdy6+p9o7fDEQKZt4NmC1ggmqYUZtT2iAj868xzxhPNxI64Q
t/UsB18YX5uFR4J6Z701xHdvFs1VZRoMroFUm3sIBy0RbRZ/QTjTW2NzBAaL4/Wz
KMYm4IVjgpsJcKsMXNDxAWBnMJEswfAHZjqOkr/2s8c86dMKvGZR+HEo09ofmqGo
hQAmg9Y2gW8nzo9p7u7h7lssolFtMW3iQD+49RhF5iTrL1Bo8J856DReApY5BR0d
3QXl4LJkABPnDaCeVQ2M9TlgsjJYmigyrs1FKs9k3X7Je9R8E1mIfn1P7bhzlwDd
GUelh43U0bCQ3bDztpbk6zS/hTfrvdCWPQRmveUjUCQhYqsaANYZQ77v7iCNj74/
8Dq9eZhBpi/Yb6EWVb2MHZt/YVl7WQYf96wmZ4yXXRvN5ITDh83tvPCs16SGNkRL
+fAUyz1D/qfVKlPLdLm+PGSVgLNK664vmOg+2ZEZbQt1AvcAWmtfkvQZzebDuRTp
TvnotxVJj0KVmtThNkdSr9lZd3NvyEKC9XfRyEpRKZmEE7lUlx220Dh732DlcjVA
xOFL4dzSrxI2hHDxBKwT2PrzJiHJo0n0iKb2tcFQEhvVjHM64N69PBYVYpwgh6JO
PN7VAsccY9cWH6LIqRwPuUO+cwxKZbDKWvNyXmwYF+OaqUrrR5J+PJUUFsuptbH7
de04S+DOG+FiR6Ko1T/lgw+2T+GUOPh5o1fxmeRWQkqfqOhJjYXxU+R7Olxo2DGv
R3qcLUeXQrN1UM4JZTUNaTw079CYIF1/yAy/WgyAGAjQd1AtSgdd/DXP0/ytr5Of
VtzCOBDVNlhDilTcTtxrXqiSZmYBLMU7ncHuMvkSGDMjIpsNWzjR4HJqDKTQcuY+
FvWmKTQgBwLtixbl1RqDNuLvjgcrcDEbRgH/yq1y/+f35Qtwc6T5DfBP8u3QjMgf
xCGZiEKzJlupPbBeM4iWMHWm56CZMqdhWt5UMOwLEN3pV/p1E2EeUgkrnNytBiJQ
IkyRVYPCTw4WgyxmrDbDsXp+67d70UxhejCIDQhELV3xGryH4LztVbNAyaXyjuFq
SNVWAzfmqIKIPQ0XmhxPhV99QBgUJ54VZZd9+F/2hDg24/1Tv9rEdSzUwmAEoYgm
seKmBdcSSXwYyFH6RBIcdPeufXQdD4ODfY2jFFKKeA7ZZV5OqlDmpDI5PW696X0Y
/BV3BTcvzMgyC4LMSsalSxHKWxQOEDzZESoPXKxlKAwGQx+92Qlj0WIEYPNlXsSt
uvZe89iRTcfkWvmgGmaWOIiOI3Sg3vU+fdbcTJ1yPBr7mkHUCRHT5+2aB5p05r/T
6PxhM3mkbtchRqDb5cKTnNCxVhJa+0nKge3elKDInsi0i2Y0I1WOgg3lw/4lowsc
x39TNqtjq1KoHBqcwh4izwEfQYN4WEGEz2rLSTDMxhEenaP64KcOyOpsw9j5L/R0
uXMDvrX+qaqsW2RJMxFCZb3tMCr0goeclt6WQ+8adX18hXpupUTwYs+LMuDrzodQ
24H/2oa4MaFVidl0P4liKVVI3wMM75DOrEfe4gNdureWgRLGly0IjLt3uqyEXvy9
mgyUkDTgkkjcUkJECdKfO60Wnqw0n0PdA7ws4UqJrrCCZourX2MCajqYm+pLntJL
Z+cAsNZG43V13FK4my1zA5stLTP5bUskeXANqWjQqu5hXCpUVPwpvyf5w8yW2EGz
v82zZE5EHWdrBl81LuN+rRTFwbUhrj5HwFaAjHGVlbKW7yEeudDddB7XaZDFpFSI
qNmHEknK7baG2EFlMlV/Nlq6sneTc9G6ZbV0Gmwb9JbiHIm86VqAkb/zZ5pqUx20
W4snNvVvaPUlM5hKYYr7ESp9fkYD7f65FUvRnMtqaKb4ssfxoRARbwF36SORJdyu
gPjRmrLSsJQSo2HOitPFMvfIknTWwpjtU6ZU3N9yQPybgwb7IecU6q5aHCKT6y8s
8FL8qQurCcFovMF4cAPY28ZBBMRkilVS/FhUgZnLL4Z8VP7Lh+9jtkK8030F4qUs
2Bc4rEBQ3Ja0Qmnsk4IRFxr5izNP55nqXypVMoVK+pb+KyGX5X1dwX0reJm7OQIC
JkcengW8/17IF2/5ExSNMza36QxT9zdkbvXQsfXA2BWYbsbfFGHH146eeUrmCNmz
GDZLsqelMQfOyb4CsYK13JpNI/2DtvpKtzlLc51KLGr9p3py6ddVTLH8wnlni/0e
bA2vozGj44ws00stRYOS1ji/Iev0oeecwwWPI4k/cQfO0+bGJsZmLYqqVNALHCOK
63iOyWqEAoS+mTiNdU8XQmIvZoWpsb5nfysThr4DDRe9s7a5KWRANN6ezRkONr2J
S2+WOQh/mq9p5FrSsHBWnTw/XbafxctKDjDJBALMXk5/ga8ZliMHBC64TrYmhTA7
CscUwRWTtowg0FbPKzhrTGrkuIcp86ZwLDVW+pKBoCMjkm8yqKhVCC3WAF2cxj7X
Y4I+W+plRdBYytCMSqbIbvm2PuPQYmQuBS0VxoU0SGKpXXpk18qvntOuoOZWHclR
jlMcQpMP28+SsHDvapydRkK0PTUujLJB7TkTFl5yTkyFz1T1HCXg6Q23deIvGqhb
BjvP+EwMIWujOTJoHaOm7DRfMxKUKnJdrwS+u6iz1Z99xDVsX2UvygP9xMh6SdWb
mUz2t1xT9MNGQMb06q85fUdVY6gzNie4aN1m799W0oxZqcos2/eH2PRNsIZy7sWf
83PVrXj3cuj32hmiYURmxG+GY8EL9scnCGI8Gov8vHGr+cMBjc4Rh5SyzzI5+jbd
wZ4RATAiLIiHjh4li5+hySA3GzGnr3z9EFFaVsaLthQOlE0Na04e0Uk1exWhTM5c
0WwVGPL4Siafoc1ds+YgphjHykjNskEo40LB/xPRsmLZX6rnlK+29aM7q9z4X0T/
V7WIxaa2pUxoBF4yelt03ljqbL+2dIVMWPdiAB5xtFmPM3m/gwqU8Kxuetx5I1yl
AWSOHyuSto3/nyMapeSMae4/YMvquqTAxrd0XwTdhMZoteFAk+1v3BhpMNCiKjyl
RhLQkdxyUjNsvT9TEIdQeflWCOQZy7GwUwWtMGKB0gVcxQdnZLs4Ld5N+15SPcDn
W/1bSkSIBcc8jrcrg8O0po7OUYQOW7d9CeLbdcMDmTiU2vZOR2cSfxyLKxQwXMyH
mCwIweaXSINIZRGkPw1jNPK6yT2FW4PhfR3pr6VcQoBQ/2GLMzrFjreNdxJrhcxx
XaH5KAj0VGoGxrY2K3OCM45ZWG+JwqJe5PdhJ69UBjJ3e0Nqzpu+ZYhMsszdanLf
KoqYfUfwd5oZXLT8lwn47YPEuJfmwqSrWPefwNXhbA2nrp7ZUxg7Iq60UweVL4uW
URHN1u4Jlifhmwb1zjLtYhhz5TPflRV4q4DuBk6SM/lBuQU22VhAm+S9+lqK+2L+
wOeJ7rTQZ8dg719xO8MgYnb/X6YReZbOCiF9e2EgNRdFDCJ/wj7CuvOY8HFqVHap
eouhbREdqLVBqT2ZrMw9epWNTAVU4KKA1LTtu2/QB+B914hvM4Gy+TNuNgY124oj
lZKN0ww0Lg8UYkJzR2AZM4z/agCHfucWHwHq7Z2GylYkoL7jeROSZ8bWlsuniVs6
G6fNXsPwMS2iB+VFZzLiWtOSkQybAuK4kJTo8d21iEvHBR3+3cCdWfD1nUlwveGA
IUul8x4hS7urNIIggBjNJYcjrU7r6uI5xKFlw9YuEyLBW9bSGirhHNynOboNPJ6V
wPkfShKvxX6NyHCaR/uSGZTqecosG2irZUEqCX3kfFr5M29h8NeXRfPgJoGhSH+l
gVbGSL1+G1UAAd0AISpdV+Npz82WRFpAd537YYBSiZv81tXgNjr3oAi9eVcF8Jxs
8eylraTprFFMFa7fG6reikdp8HdpddGKUeJMyG7WXkrF1HavydVFR0TKXPM9zOe1
sIRJrq7224j7QBCk/8rYjfH1yKi3B8/jOJ4vZ6AXqPH/5+F7fN2pyNB48/cHcegY
e9Lw8e2tabrDKSlnX5dkYGzh2609q78BEyjGIwF4N9y6ni3JxExLCB9h3p2YX7t5
ssGtxIzGV5ZBKXvO1KEQ+xqXC90VRgsC+BkGRhSnjOuP4ZMiKqjwsJdXqfsrSQle
FHyGLuQMTLzKE3el5wkeNbDQ2Ivk6DiQO+NZqs9CnI0B/Y2yorkAgnJ4l9CO6e12
RDa/gmUP/osih0K5rrQpmPRGqokcryIiFmUcq6WkqRQ9s2ajSTjacodiLoKho6Nb
yZqZublpGNey9KuBDF0O5/jWJbzYEuPn5Z0MlGdvXKpktFanmoEoyflXYBqHfZHi
Zp15CprsGRZVYJMAjPJEsg7UXa1WbcmC16EcIuE0zLJgST2hxDsTJBAUTjYUPxkG
kr7XWMLfVrCEO/sa+vRYIHXPP1eyOaP741pc7pGORlIFjDSTEAW0J1acNHBEBErN
a/9RrwnSlbB+BxvEdPgBVcbxSIyLM7aT9oS+bEw8qig6dKfqEZLdAt0m7N9jCcXf
splFhAsyRMqCxF9aLKVnyPCuBw82+dvJjAJwUkJ/1kn9DK8o0IEQt3EBCxHW/eu7
PkAJqTo+nx6QC3xyhWBOKR4LNZPfoo8XQUSQ2zqxcgjTUoBduL+XA7qVk4SLA/Yg
EecPYtSirkOSvn0EbF7ZD8xyUC1AaWfa2Dz9/1L6ptwK71tMWY689Bkcn/dmZhBg
CtbxweCpwPZQJHAqZ3fT3k7QM73RBcJOfqNtj5nP0UIBa7YxSF46aodoLJD5DlSn
Iv0aqZ+QyGXClP0SbjNedCVBc/TbnWA6nIzqOMjCMhr2/9Yh5xHDC0cFzrKNd91o
wD1N5P2ETtlAdFGiptLtCAuWijN8iPx3iZ5mjXNrzo7ElrUmEAY8eV0QhxMImgd0
l2f333KOdPJzgq8HRJnzBS/TqYkCo+3DRQZGwoIwuRzz9grFMffE4BeAcHMU3sQE
P4OR6DCBf6W0R89aoyoRiRRKiwV1HmXzQL9e/863VeK99OG+cxWN/fdB2tDSMdC+
NAJI1JJX1DSUNcelA8no6aUVj39X18oi8ZN1FUw00elbB9RD5Xu/b0XL51/eby69
UQ5zGbmfLWoMPrd4ZbKUTaKF2cckO0FJRx9iPP9/3+Hd1w/0U5OEdunBfQ/czi2B
cDsfZDrvpzWhZ2Gi+vWpn0NzBhdDFODpXwy0KDR7WnYSM5mFk2yjrzeUPs5QMD60
pL5Esfv7dTyWzYFvMuWcnO9VwPasYq9uk6RQH8lhyZUL6xcpNu5wFBKvvawj10Sq
5V+L/KykPUSmtqemI5ChKWG+y9G44/Y+VpmxQD4kgBWg+VZLdEr9VGmqnDKw1DoI
5xUlID5LXEm7B5c6AdgJ7ns+BG3Rz0zutaW5j1ana9jCeXuLFu9SknfZwDiFzfCf
CVswRLIH/HatHchOvue6Wj+5hFejooQgHR8y16Ku4fkAhXUhktW4JC00MI7b/3aH
uLYK7tHuJHY4Vzebl1tqddB2jqgngDL+NPTdynUTbwZ8aU3djTPIMLZKZJRxYaLO
Qe8ljb0JC9PVINvvsmWUOzbyw7wfwTVWlIgBnR5QgvNjJNheABPduW6LD95/JOP3
+UEXkFF0EvuBjXwVGnqlse4n68Yein3Gl1W6drw8c4RW6HfjW+DNM/Yk/1s38tSl
4yBqmf+5eI1GtAubwH+TKcf0+BxViQlkobHLmdAC7+7eFi8NWTk5Wfj/9RPK+jhE
138TyDPFtZqyIriZQhoSnhylic/ppeMfMM8u3Vm0IukxMlvmGl8L94Q2qCpMYZcg
6woCaoK291qDIXANfVWNyNg2fdR9zfyeMOWcdBEbIYPs2q6BfAjcgfmYIV8ZsxAQ
QTDHoSVlRf4ZTdJqjZjTb1Sst7sYXSK5yjP4nUAHivL06G7OAfX3HoDOTLV6uZpq
krswEXWCvhucIPhl0cxf0wtQZj2EgU0/NU86CKhDUMPECNrF/jzxyO0/X2E077zU
C/RXAZncuZabH6ELgyoIAkn+essy1g1xzbJZHXGvGvQdAZ4IwPKu1fFWGrpy93PO
dn6Zcj8+r3x1dYke/KstBEnsMJYrmKyjuy7pdztS5YUW3UVVuKK28oQKD6la/LfC
zeWwjwnDqKzDnYKXx436ahMfIghISk/8B2L5zga4H1V0xG/wnLgV2MCBo+9fUALJ
BgrIvexXd3Tt/vmB2MYopTdgt1xyJ7CTZQoK86qPxU3hcuIQ4viCEz+s3LUlpNP8
5gWg2ACvY6WUWgJf9hjB6WA/CiFRf8DAKSGmohb2ABA180O7c6hyEGt+l040q9Uv
NPQIaB7Q0OLS/daVeKrM0BHbslqteIECFD463XeU8GwMX8HpXqxfEvSUwa90qqch
KbTXv3wpapZsMoCbhN7lHeenGLQLfyDpofx3vi0kxHYUNxz/xZevoOtFeoYGouuZ
hl+QDr41tikkFJhKvrbORyPRxtT6JI8NMLN+kEjIr9dsv82Nkj5La4tGEVbP3y2O
RO0HBCB9KXy+cMo4K4Iha774tm5ivOS7dXgqVyhklfESdFnHP2EjmPry5mjrOoWP
hBX28Wa+myluxD4OOhOmfn9BZuL75TCbaxxnMcVn+MSVzqMAo0dPUNM6Oa+fekmq
Ey59MM02/zGftY6qB5qYO2aBwN54o5thJYbsBNmMfKDA0oC2MbR2qY9ExvE/MNOS
d/3ibFI7voeFDC0wjHF9/ANN1fpeWhHHcRRShQ8sZUmuslHeKRsV9f7yXfIDle/Q
4sk7OVS3EB830kZ7siTX72XpedRqZRqNjZiskr9xaXIeGN21KnM2FVFbgow0VBXY
3TneWhQYBzxlS4uJzbw46Sl/dF2S4jBL5947PG0Xs3ivLxz8ioAAieeriL9et+8B
y9cqlk8pqh+/VjllGyNRx11wNWa1jKCfbYMGW7JTClqYNvvx+45YwDfm+3T42oPm
cmOmwBfG6+QKehEB8bAZsKfy0tZVgsDNILa39DtUmqBIe7JP6f9JZ+1sveZ00NyV
7sV6umAFO/HT/ZxLbIJKEVhC5L8AEiEAElfNCGb2TLJpZXtCMe1rpmqXVXh151+d
/QRdh7fXyzV1g1vNX/+sIf24B5IzpYYaNXeVkuvDZjb48Cohq/OQJY6WPENS65Jq
3t+EjGyeN3SkeKd1lVgt8X6nAVz4tV5vA6mT4Ix86yIznIJX17ARvu1NrOb9wZKM
kHqzGbNFaZsl+wiN7pK8aksjvuIUHC0SG/th8BOVDkVlDb6EwSwhgVAHlHbFkXG8
sDOCFmYKyLGerx3imMM0vwjOe0Q6kFBlFbujcRHUuu4c6dFITGl/POE6iErltV0w
76hy2JqfkqOJVBjuxoMcLx79bYqprvSUEMh/c4PkY5R9J+AaiytJ1kv8kLik5xEf
8maRV6O/iCnf25qdg8RVJvt2n/P+WA3c+E5VP+hG2GBR3SZEeM1TqPklm9bK/JDw
z07TXlHFSiY6xkpV0QAy2FzC4RJcH/djnescmLLoKVfaaXD4DPdfHJrjdxJZVZXg
ovYa3lKLEwxMUngmcb2vTjszQ360L04ZXSAMnAXIs8c2oQ8ufhajMStXqxOV8Byh
FLtSjbe1/55gRidcaVCp89bScLNi0ksyB2fp5aAx6VgAGXYPCjSs7e9BlPODfoRR
rMoUrg/uMYLGUO93Z38JSLsuNFGf8CuCrTHcEfD9eHd1Yy8Q0Ct4q0ks+m6RnIzW
MlNUlMwsps6vMShRRhyVXldltGZKdFBtlbkXLSHYCzD6C80wd639Vb/NkuxF6DW4
yYUtuxSWUrTsBdt62YFgmf7qriKmQrzMsPdlPXDvEAm1hApmbV26x6aSdHn2mEQo
LVDGO4rzKYoB9v6qIdkOa3Qstql/uscvhOZFZ4/Ca7s9djSm2oS4Xnk9AWICfOph
3jWsYciiJNi4W4BQnG8FrVPKecS6PSPh0QxwwhLBtPJRszVY8C8L3638Pf+19o+z
Ilku3PiaHD41HS2JXV+QhUbuln8bVOYyOh4BHR3e8dIJN+3sy5ygPsHXsPdq6asL
GI16INaP8k8VMfBoi62eR7RbpvqYKi3YqmW6jDhuIVYKZ+8l+O5somhiWKtJwjzv
ZMdqJy8PvgEtR70w0L2EMCQAqjvCxzsylKXtLz0M9kFwBwCyH4fF3MmylcXiftBK
TdJSPJn6fHTxeo2iAuuyAGgzEKsgAhjlSROxLQWul1Tgzge+PyhVpBSt7fMRvnj5
v2mNqnNiTxsstD6eNB6stGg6JzZAGfWQEmD/zXm2U8xc9pzjLytrtduDYr5ajJzD
b/dRhkixGUT5vUIBpXIE81sVynCXxe36i5vOB86WkAn/SamY8Q3tmK7BfbkNeybE
yVef+KKcjBzM7dACDVR0CFwT976dAdGwYMbyfnbhCC275XIPJMofv0uEBLvucqvw
YXQbGL66bDLMJEWdisf4Ex+QA9t5ZBZHl9TM6LhcwPlG4uSKS3cbxl5WyFq4Rnt1
iDzXlS/ptdKZef4N9LHMfyuj6RQCkWHgSagArdi4BwFHym35sgigX8hNlx+z44NS
ZlkWPwS6HY1QfL7QA6I6Sh/tuVUddRX2ROn8Fa+PAhh0k7ug0Xm2SRjcjbWwmBb8
V8K2A8vppTtS2n2W/20o/IheUIJFOFO05LsSvhYgORfsuYOFbYr8pSTGcbp5m6Vi
RfvIMoqrcpE6k9ya03GLl3+d/F4fIyVkSGb4M8YLEkFn63N/DJoO0czn0UpRgCmb
s5+7GDAtDL6udePTtK8nie4JODnkG1QEtocnQlpUygiBN6lC0FL8pB0ybnlOOGOx
9r3y8IzGho3RTmN4h2bphRZRocvsyEJ2XHoDMX1NIe2IUpH2l9YJAXTumKKPCvul
mcMtcVks91UfUXVK+fnpvpOyht8MAUkblsIvabrZi+6OqiKZgY0NMd2vMHYsIoAn
lckFltAvErYlomdCGY4PLBTz8b5RcvItMJqDX6bNcFGSd8Nc8A0JoyOVcjCrtxE0
vf0mOsYTd5sGodwNWPHD21mKKQNYbwyIDX0fGLMZo1ZKQwaYWAY0NmZcJEq1ql+Q
neS9C+v/5rv3qydiQZgKWXStMQaNsXY/R8kuZRKeNewFsuHkisSiCqVM/m+PgbE7
izVI3hnezdV33Urh64/fzJZoMbLr7cRXYqjLEFpailsc4835zsQ9BVSITYChriPs
V1ozE+2X4tZqlriSw11E4yFTVUXv8kYfLCdbZb9zV4U+q3Pq3TJFXQM5nEnZa/Ga
/XOC0Rh7yfkYokTRXOUw3dmPEIuOaCRahAMCKRVMdBIpUe5wBBSKi/N5hJ4Mssq5
0PgeU/WbTtYpkg+kmfkjsdndWR6Afd+kmuckOlDszeylY4P+XABwmR17mbpylvM1
rHThFt1V0nAA55/d0/KQnsVMQyyF7BNnSGsPax8MoZFrTRr9B5YvxJ8EHN5iwAtw
5mEHBSs3niPzAbLD0apF0EcpHjgBEtKWto1gmo3PrlvXLx4wGaFBoZpNdk4FppxF
h7mrdMcfoyY+Wn+wUlzgPLrjpyxmG80RQ2w2keqX1F3LYQSAvE3n9R/GpvdKrmNn
qo+OaKgiPXaKedHn69QbeEco2Q7iBwEPctm8dubCY5H42rp1FDiTa/qSFP1EooG/
mvIeP2EIXenuyGaaQRw5rIx4Nt3sH0S3OtdhzVtw8ejkCVAO7e+WoXmhqo6uv/Pq
zRsQK7M2W0+OBGsnS6yMXmYwCWdYywJX33FCkaR6EQSXbKKPxKroBL8tPRYj6SgQ
M/1uTHj/EW0en+q/dBLdWtnDRbx4kZe32VCvwEbsQVE14NMTmmCA7D9Ssnq6lm9E
6+WuW1bm/twM66qk2WT6DiAAbLyBHXpeCE+XR4O0K6kHwU1NNt8IyWtb0xx9LExI
5Loy212V5/SvVgUz/iXgmHP/5OjSZSrQtYgiJsli09t8D/P+/1mP3nO4gQL1BnU2
bUQDNKQhbJKMAeXWf1MVKqOUGuI6m9a7iMKrRbu2fsCnC0Q7Sz35AQfAt8BJA3XJ
w6dzmA8FKqzIe8ZPlTg2w6uF6Bnf5jS3/9mOMQruHdcYZmk4twdJVBHEmq7CGuyU
hDuyGA5GacCJOwFU9WmuWlEi8RsnOKblGJ48SJqjxf2r0KJVdLiHDinEaVA0Rz0I
3lRH0OyPJ2kIfYQAFgaioWeQuFNdUBwRBxFqTx3R7nJOofRRnrS35Ej52G0mYG/r
TU9xGVUAtb6oCUQBsSMuZnLoO7EoXAqmGMyvIfKDIOvS5mXYz6IsUNpm7ZcjLFD2
dBhJtadBpT1haIc4d1KaE3odPGjxzlbaFjyJWvCCkpWMWl+THnPyji5eCCtCJTO7
v6aCHuhca2Ke6uEjCG3eIGiT6vEuRlJso1MtRkt+BhDpxr7iWpS/JGBSDM/d2zcn
2o4IkhKk6/eqPT1Vgj6PUGmVcjuoHKcMJUyrj98p/+li+C9MPGGNbr+iFCKmFUhQ
qy6TU+d3If0cFamb577ZY30Ozv5csIJ1Yoig5cgW1AgnPHNkAxQdzihEHqHKnNNS
+UqKD139LcGBeoDObzZ+AfrAjDaOsQLWc6/0D9Q448Olw8ZGvvXA+peBSw3iz038
xjZXZnrHGlARlkcooNl5hYK9ZhqU2GxMBOuThHBnI7UvIF39jQRt0wAj2Gt1uigF
OaunSUSoz2j5iYelOrAI0lxmO8ds8wjOagn0zRUcxSE4ax5iJgsC+H0HgVOYM857
IN7b63czqyRcacagZtQwksCook7VO3klSg2me/f5FwL8KnUxISSnnKnHOJKSXa3U
0lu28oOVLX3rFQsn3NQD7zZRzsdaAWQ0qY3eLOdktAfXRHqBrf/jCCIxN/XGrF/V
90WB+JXnJtMGFR8TwLLNYK6L5DstMIoAV61U/Dyml7xQ2As5N5Jd61e3A5fgVLK0
7iBUuyNTcycPvg1OH7FZpfmQOjEl/KFaMQ+VFq96+0musH0gFnA/WETSh68qEo3L
NxxcqUFgzi9gq1SlltOIqaSHbgSqsQJZd0qKS8OtuAx6QNjy8F9wV1w3M++FwHaD
QbD2xVyZpAZo5ydrt+bXhXNKXqPMWJYS64oIpoG4nwsQN2n7N60KvmTnha3iisI3
l+G4xYSonccIgr/ubJjz3uGSR/EIpMJnk1cYHpQbg54h43Frphj11Vx+ehZJ1ki+
gUEKCoYpbWj06yplOFtKWA0ffmPwMdKVWvm0jkPwS6uhQRlw21jIxnogyX+Af2Z7
OWx0Ne22jlkZ9iyYLTmMXz1AJik3GlkHCWkFN+ktHa2ukisb/xdMDlWe0uRiRHaV
KXnHWIXKo3YDCVmJ/sMnPOPMbbf+vOdsfy2Si4VAtezNs6VJYQ1Hp+K7lqE7fNHg
3YimD2/TdH/tFYWC0xYWSONN+EiTfuWzztDsBAWTYOUiXwzqql1i60QzZZLVB3CR
p7XLwRS3pxCJEenOTeoJEIeQYP+7EPCw3Y7tsRU0VuWcVqlEzxgyW+WDsK5H+lPG
BqLCR65qaKUI83h9J7/omoT2sxj2J0BjbBb/ALNa2IRzO2SCwKFPR4q1Fz8/W6Ih
TmmEOOmpKUxHuQDbFovgTpiTp+IvsOMtWEi8+EKzqm1fnXIFBPWAT4wwV2c2F7Nk
XLEgqNRYbDxdKvH3o5EtRku89mY5/M6wpXj2T/meeIIC9w+lbvVWbSZoOA8pnixv
qVF0ZTUs04CaGscF/sn+gIk/0k4AenkvIxx5Wxu9rp8FGHLcZFEi5vBDYSWgZKoi
Ic1uDyBNVoWcJrMNv2c0NCq2BU80cQYJNA6nnT4DWVorfJ/e9WksFHfwpGBacLm/
JeJyj8kY6hDU6hIujTmj5NlkBOUJxQuUo6QXOUYMXq31tHlfA5QgcG8g6wSYTK/T
U6k6MksR71UopoCaA3hjxNofvhRn/Ji/IXRZrZtOWflYrgM9Gz4szWA9Q5XJcF/w
I1lp+DGxbUFPBZ2jewyGSEiARjZbil43qRfkJEHzNzbh+ir0uFuGWYVB4z47+43E
S4nfKXB7thIwrHGtu32hQK9Ie+o6AVpOqVhJD1acIotOuP1d/93KSoqSyPcxF6VI
JH0iT7oG0jXNGvc8/Dkjy0nMwwvM48Pw9qLZfwa9gcNz39m82xt0JKS4jdKmKYFO
roQFgcrJc3KcWpVFU0TgSDeZnZgOmdZoR8cA//ivxr8yhHjFBY+fzLg5aOVtGz35
t4e0umQZeNrXjx9t9PuEOONspCYu7WnFdYTKLYtTXn0cc/G28e9tPJvdsz+/DRML
jKIAqKmuVFxoJA+czpSxVD8+nIrGzgSdbdOUb8ux4nTkBGmC24qj+3Pyr7Bpokir
OodC3H81baB2TXmE0ND57HkSjxdePfjrMrtYpzamXGixWFIlMIomWG4WEGdRbGpM
yuz97mwHeeYllfFxZMiO9gFmChfD3NCzadVHbWAYBnfJoowdZfDrky19f1ApNtAl
86LlBuNcNSw++tfA9VeEIPagZidp2/fpucQqhy9mU0Vf/N1JPKXCDvWNloFawXNK
rpVMohpplxAXI28YuTsytO3xzquV0w1f7fUkrJIUjoQuUyYuLOtC9RyNX7VM7s94
zp/1CI73rEmRzatm6JkerJko9H/qirYvDLwfGWWegCmPbgbFiHsP61c6un3jL0Cu
8hsZIGyJnuX1hS6ANDper95ivu2D91ISznBMhzzzscN5uzW6iyUns+YVkrBeJGii
YDbIvUmNKTvE7SIH+ygiBYzDnrp1LGb8CvRgXG2QHbkrK5egLW9TuGfF7uQ0qAyt
MOz6U8OSeDL+BRD5uZemm3jq8gdWpPYUdqnZq6p/5VsUD8RAkNjpipXzzeUE+hBv
vEN69CjFzLRbyzGr2+cUMEMS1DqTTrpKaBVlG06IYVgsPhgmWxA9qRUokKQEtkqg
CDGCSLpR5HeGTUqrrzmPmtDpv0ZBak1BQoceR7nrD+oEw7YrUfQ3IOMHD/KiluZT
H7DNWvDHMc50TWspNdYlmck8UxlYDJqxJzA4mFHB1kHPAVHa8R4loiN5CaeEtIQ8
p2ULPRz/e1bJuF5heH4CIvvhHm1ZAM2RIlDlzYWJ93CYNRnG4vKTV0mxTXUeQs2h
Fpc+Al4NE44d2ySbjVHYk9onAxmBIFlVQB+6jOIax9Eo9vkF4cxW+MNdmdTl+UR8
3VssAmVZuWfnkDTCqNgOrfC7JuvYj4k+9ja6Iz1PvDTVSH1AlXo1ANpFnpUq/TGg
4ZfwevpI2qOUu1GyP3WdbNbpqppKfZkMwfWTmCwr31Z0t0ISpKMKQvYRfUB8Yrx3
zwMVqHxOsIgOiIKA8Z41xo5MNOfXnMJKiWzQt84M0MlBofQMehcn2shambUbSrX6
MPIBwL5sUBtvkKbW7ZJXJRjR9u+ILTDD12f6G9pKONkzhPEHW2lnQCaNfG5cU9Gz
TMC0TfVxXvPvQ6DxOpBuAJIVjiN/NRlhW1RFYc99ZZD6OqWWqhdUutAz64Nhkd8I
jZMSTyOOnOtWUcoZXoFzAHxcyjjeCTO6SdGSH4/W+bRbycDp7OetaqnZoCgCrKea
q1srgEMR8G8aaBrbLLCNC+YGNAjMUv4fU0iu9e0icvPYEIkzF9jZPWii5NzAIn0n
JfcERS4wh1SVQYsJzvj/P5J1VVQbubhcRcXvLEDSCNr74b3B9iAuIt1NfA6SVOiV
jGAHmdT3rpolkUaJvmWpU3q95hwHWV18JgwAfIfoNyETFKPAEMfhCQPexLsTy3Pp
jgrlPz6ZSroV+u9sngSY2SO4EzeuJvURrUTALxSbd7KQtV7PHq7YGBxfV72QMuGB
/N9AVwEbLGYeEId6U6nh6Vot9Rh39w2xqgXoOUyX/0pA0TcaUK9F7knX4ObKFiox
ZxhZSLQjtKJvtEum4sRbTTNa4UiwLpyBJioc6IxA9c1FrcP04BkjWropZYfxllUc
9elYyZiddcHFo5ar4EeLAd9v8Y+q5bQlbK8kDbKwOO+EZrtimyoixsYmF75bTPiU
H9/aVNRPlOcOoM7p1Mg2G2qbyQRB0bXmWFLwwlrxr6E0JqQyMOVZeUt1v+zCWwmG
puoPfJBs/6Rq8Z9H2PmwFLt8NtOxhAOYVCfAz44TtD47v2QZhQq4G61++8v7v052
6Ezuca0lQyREjQCCyB3LpsuPOL0owig4LZEoxg8GUGxrUPc0M339A0eV5ACuHksh
EqTtatidSPpRCwS05aqnZe69hJUP6iBtCQR8tkoyd0MPtlCSV/T8fto9dUQzgMXW
XPxS6uOC/bbEgZ3CO4OkOuDhMgLbsziYHCi/13A/61nARuBg00BCBnVCo0ci7ObX
mqZSAfsd866jIze4GTkslMPnbAwl6McIFWr/S/8KUINovUci5RxWECmSyvQWJ7JQ
ECc3BMB0g9qa8UKrIvnnPMvIAwMquumoJaAF1+ic8fYJRMEFE8rxAM57iBfJrV/8
Q5UvZLwov8dx8VY3pNP2+v/f+xO/Sew49Tk95Sflajcs0Uz/wEr1ZtYnoup7aRgd
Cbt6HlWA6+Y2/kjXYms7cEtYj4FRzBfhSy068GYocqgbvQWSun+HmT7LnQ5x6p0U
l50hZnC3PGe0sk8QyfEav/boIo/751Ov3u1t9Enm8NlVj2sDYZ7i6Xga0rZXufw4
btxyccn8Em+F9TE1p6CX3G4LHjVbBbi8YMRc7zcU0QCsO35iLBUVovj3z3egmIh6
IwKCWgzXS2Fq2fi/Z0Kw6gOocCDevxkwQQyS60Yjz2GNtfFIaDsWj4fdP2D2i3wd
wOa9OIXahZTO1dIJE4ejtNLCiki3z8vGbofSNr18PVTgw6YVXWcmBBxOaVqCltsw
PU/Lkd2a5JODhdwWLP9//KWie8XYlmXDAubnAHzwT/YC0otlLxU6OsEse/0mTdJp
VK9VSCvjaHhD87X/3c7B34/ZE+JFkddrg8ZqsI95rcDvHGSfWKf3Qooo4T4djrCP
SnxGMF1vFEXHn7TIYImR1L9gZSuUAF6MqoMBalb9GhdZ30hCkOYuAtEZrvFIrb2H
y5xikmrlMkRIyQ/DbSTDMBvr2JXTRklGsEyHrW4AfRwk1Afqcfgw+nDa1qUajkZ5
Q54CtVUewweQsCzKx0c/8cMwQmRH2xlU4aTnlrxww+VWggU3i0NZfq6N4XYisl9b
zdID5nA4lvGMlUxoyErqXaiZbUwtrCHqpFrUPIiTBuT7LU7MTWOThS2txxxS2U3Z
eGyazDU3wEXKIXHsY0vflzwyply/3THIAvMZ2KoT488okIB089SK+1e+JdxAxtJN
QRD7ClcqbMT9gZ2DY3m7x1bpMFdJmqczRwOHoVXkaUIzzULoCMDqFt9KtUSBd/fw
yqHKFM9HioSKIRAXjVfALEzMAIHoTVaIMJGTxzFaOBaTAAphFq1x7Rhy+RlxxrpJ
fYwbXfokxSTV8ZeQN9wy+6yq2NDVka5zIMf6YmCcwj3Ho6w4b0oAtgxiKaQXDYLh
lCYwjF4Bu9BhHPqfbiMCYV/wpJDH5RSGk265IM6CfTbgduSChVuj5xbFrtJsJQOe
eGZz7+bo+AXYeB/ibDe8j0ySP3bpkmE01vsPHEaKS9wiVg7EHqUhdJk7LH6Zx8HQ
/KPrgN0/RXbbpaZ8jZQxgKf6SsNm8dh8RVnLj7rm15LIekkPdmCGkROi4bUrdamC
ap8+M3RBAvilhCWx08n9WATnsyz/R7inst7aLlEdB0mwdlKMasBQ/0NVEuwV7jK8
w1xSPZYqlvhtMX8YpDVdnJmBuDHd7xZfNIily2QUMrMvcbO3M/i9/tLdLAiGSCiC
Y773raVbx/g7nxDxtC/OihvZYMV72qlWgwhnEozmmymlwM0CyUajO6eq64MXHbav
lIu1/lrJBMp0z4gf2UySXt7NVkDhaM9u9EUW2hFObrBAImm/i0gI3dfb0IVov5Tx
E1x0an89uBx4pCAlhdbpw9ck9NdGonJ3OuHuMOBPcTjw8PSrVY/J75eNQrhuF4EB
M1sDxhiJEYmnmKgJg+0OwhplHYt5W1txhYcz7sg9wQcQv9eHKRi+d/oO/rCKExzW
4jsb7wV5GdTNnQbCUHeubgIEo6w/QmbIIqYOWVTqke1MOq3Yc2fkRWBnrnFLB/DO
jLVxXt5KcOQpAaLqRQvCltoXywWwsa3hBaiT9JcEyeW1HfSvVIPL/4ggZLSZqIVf
sMIdKfFucbnYGGGk6vLV4lc94dLgnV9qpLBT3Th0s6WEgDKz+kVeE5J/l8MkVjMm
o30P+qL2ABMmxy7nWMnP6ogu6y6IsekUXZp6IiIRSIpVy3i/9vMrgje7vagCozWO
yp9Jvbyrk0sHWXN8lPmnuRkyKHJtsfHoSkwutPd8NIQg6NL8UhwyQp6EzrCvKssn
a0lEDh3ZY+ebjwY6YB0/b5kLok0oAa1QeV0wLsOhKurzU3uAbdXOAB3XEwOfJtyu
unnzyrTM6+gXlGulPX0oCCQmpXHe+oREIgTKN0Lja7x8oVy5pNzeNGSE90xeo11b
pEdXYL3fjUZ136qNzbpxfNxrCF0nsPwKCJZV3ANPrmVRLA3kiumE12f1cwuyedPM
LsbtUwhXOkCaA7kTS4Sij5nLwPzfbpLzd1awD75C4wapuX9FuIUdMd2noP3KD2ZY
Z+ogsL05hmfM1YUHG9O5DbGqneM/WVEt5qCukH1jCBZChoLHnnnmJokGg6IasPit
7bTNLqdkwsFYvh9asxJhZ2FrpSPDL3ceCdC2Ohd68+UVZAd5hI6/3tLGpQKUPZL3
a0mF3277kWSN9dZC585r0w5/BZfd+pAADHrAbdGWs1sW2eAIg142LZVRFLjR77Yi
2THsvX6B1BfqbQRlydhq0XtOypUptmLtpDdes1T0fl9yXb+EmZQJCljrTR8xuiq0
AiMpohaWfG8zxPQB6YmTm0qOw305BQACSrOx5lANowTBwLa3JF8LHN1n6OPaSIMF
8EYWDX6t+1R9Rbrp49pfsQj+SpVxO17uDY4Fn/jo7j+69CMPf6Mvj1bjccnyE6AY
K14Ki5fIsZZS99b4wDmxRk5ybkZUm5NkdnGSwBT1OpgkN9SKqPlhmdqwvWSmLPY9
pWN1H/dsWwbxdLiqwg0EPqtS23ccNvmQ1HfNYX/rU0jPoGEiKQJq3m+ZoFAiJrUc
3ClZiP0wUqkYGJfek0Y/U8rnph+khvdRS3yG+lnKuPJlHkybQcs4+ZsXHPaW3W6Y
RWAas9EsbR9cX6uMuinaVuJxvQKWsc0NgZt8RosnycpJ/eIauT73dIRQVm1Q67cY
A2frhuAvnTvmuMm5x4EOv97JJbwwE19H8tplAgYQLanXoBkqn2TXhQCwo2vL5gEv
lTk2fVfQg9Yk57CJAA+se7aR3i7I4cvGgTzoKHY8Femf2/buCyDtJP38gqYqhCmS
Bx8oBBKabiKPQzwW6x2MPlS1Ow+UbwuM8eJZtg2Z2pJUnObGTB2Y8ZGaWXJ9jl/F
2x7pkxSHGdRPJAemqd61KiZvmEFTt/BSiSjEKsNdf6fpb1JqOU+Pf3GujyVfbIIT
777tkxHLZV8pgzfFhKyHmU+Tvg/VF+WypdjgbhUOewxCr6cKFVfNM+YDyMSivce3
zMZm6l2ZcVQf6L0wM8Z8OAstUI5xN20OEUauHb0cLGXJxQAPB36pju7Sro4KHtl/
wfTxStoxuFZAo6wyMAgd6YBujVkFyxEJpwtn/s0gPynLaI3YVBzCR7XesArdacRw
j3SNO3Bu+LjIOgL5dQZ1dDJi7FpLdHuymuPxnZOJ4/qD1z1gTjmn8n3zeqx8aNm8
H8HzAWTsbFjkrLwiqyuFbDGgONLed0NmBIbE7ZbloG44GFljzEjoAXkmvicCutgJ
c/5VKDNPcyKFDnz5WH00BaJu+Gvsn8MbBJ9aCvrGd8gIVcX+0/CoK3TlKjLOznyg
4uFTte/4kaYj3vncqr9sU1oDUMoNP/HKY1YUeWrPLmCjOZ9YNgJ5m0hD3R6PQHRZ
r80ZYYaaGtHk/2Q0exKiI0QR5yOx53lHfbu4efn7eAdz9gmXs5+o2MzY9QX9kKix
C28dvYsvIEuuDfKdOR82glH1/VYUpXMVQP6SAqBtUK2OcFPKfuZz/944tiyDjpoB
PYDca0+ag/0XURbOfE6cfwfEQcUJGve5XeyGXJCpKXS6AzdWsuI+wR9oCyhdeZcJ
Qr2RxyW8jkGcxFWp46x6K4dcz7eu2iVvqjbFloFkI0EkSmyfWKF36ZkWNZYc5bGQ
kB4/kaOsZeV4jSVd3z9WYOd734Rphr9u1k5KQjQayhBxJ6lMD8ssDS5dkeBn4XEw
YfFyc325trwEc+YdjCzpm3yY9IANFjVA3gHSLlR75+bZ6ZCWydpC69+tf7e3GvgO
woLsiYXLDwajBToT1OURdeUd+7o7RIikbump9lZgefpGt3DgUXTx7cxSdw4kwMft
424Jk4EBx4tkSeSiHRZ1y0e9oW4PuQ/XAl0Q8lV8pEEWfj9rWldVx5Iq5+goBmFp
x8rwdp1h41I94/DVLGR5D25XFSLGhDby2V1aV0y5JCw9X1thIl80AIsU3pVgtCjf
NA5UQ3RfzF+sRonOyFGgY6kQnARWuKHKyeiJl5uFzVGhZsM1vJuQrmUlaALMS8wH
z9RDLnMxPsqxX/1pHohUkfc44GVQ7Susjd+XMh2dzz3cWJULuJwOKAXFjA46Mfbs
pNK6S7Lm7JoohG6HECwrEJWNPvoDKAz4xDax7AhreO0/6librp0f38JlwWfAG5BL
iMLGPUGndOWELIbS/8hXgy29sFYB0FGyZr7aYONjggOLau4eFPZn8/dxkZvArldH
x7YR+vixwhqM4X6yPBfHUEzjWrJzn3FOwyzz/9eL0y/0RCjobGQyG6yOfDwMePFj
jwwpjds5mkhSdo8rK5EfDNfE7NgCSDi5BCd5/qCUOGmvvmNwHx2/s1TK3FTzgN69
1t/di7Vn6uSG3Tyl/MaG3kq7tR6T/vRbDvdJKwW2maOA0jbmD+eIk1Gvnxn8t6Br
RGY4RjRyPPc5Vjap0qkEttoGIh1jIjCvOOwmClFTkSedcjwg1XvI2/T0AQBibtiD
r4lL6A6ggrWSLTm+DVQ0+9v7QraEAHGaN7bov0bX7obVTwe36bru5KqaHX9QcGK9
/zzKgnvs+XsNWOxXeUxL4W1lzu2kkkW+cWxPuQLyufuC3cKn6efWgfBFMn/w9O/O
ySYiSYQKXgeE0+jnQRFmUW1PhFnjsurJTsVcJxKS9t2Dzbng+b3aaW8gT6GC+Toq
ex7DPc8e3f25OUh1CyApVB9LxyJHwkmOd0j4nTPjznqXY0exCcwaTaZlHEyWuhdN
3F5z9O5B1tqGK2xN2ypjIeRNW5w1vhBu/YL99CXeeH3kc39U/ZJsPAQ7wdYH4SaA
2/pZ6zCrWZ5IaxKswpdlSVn9rircdreNl1lyslHegdFII4WVy/QRLmoZw7CIWkfL
tJC2h1CpvHiH6jmUqknX7p9MxIBYy7dyYVZt3fTqoSXRX3fwUX0372gstpqA+YKM
PMMXa7KBvtDezo6gTIOKPsuIpkyOU2CBlReZoNC/svP/IvZqvMK/FAunYKeMn82f
zbsGEbjRyPZCxnBFBK4E0E9Rt6NI7CfqA1umxRV2Hm5o28jI+yyDxrkIcL7lx0S3
oAO+EldjL3nh1L6CAcEsEZoSwvEgQod2hbmfNos+x5PWkbTABqlZRcEIj8Smtqdi
Na9b/g36tnAM/7NVcfzc/7BFmaG2kd1o2b+y3HHVJZvQaWzyQ/Z1HrnIA0YDOXjn
e8H6KnLJg2HuXGjvodagjVtZBmMkSOjroB7EkCQ1eM+UvG/hT1M8hlM5FIqkSyAC
cvjP63FAJbFfmFEhoZV+zLkfC2jkIFlOEpx62Mr4cOoHlVSeZgQajBTrXV9R9+I1
QC/J/hWGhbpzadTE1q+P1Ofe93RvYPwcxwu+OzTFAorU7Lb8juOgwl3ToEYImh5W
c/XxtYa3PbBey1pi4QluJq44XF843N4/TU4f+QynkFLi9hVkhHz9kQvZM8Oj0khH
BT4vEbLeMztNzs0CR6u/EhI5f1u1DVolmkWfomemgJsRvXn48TYTCZH7DSb0qyqb
idHYMhOyTwzbiEK9KXBo32/qjyi34q5uI/w3YkItMKKmGND8RHbpzNqI0bTH3h3j
g6KpuxsoYqE+FCMS9lJ7YXMujqRRRvft7cdZGY3BoJNeR5cjuAYlj6IYuQCbnFQH
KTgLMjkTFbfwvMIsVvGloZaC1846/30jheJfYRpLqUq6bg0EIikWTrSGDRa9s5Hc
LW3xvz07tfUVmnq0wdvE/qS21VT3OtdW/EorTgB2n1aPeYkH3kw/m1HT/JhbaXzz
KHY4cHJrjfHh5C16KrAfABwpC2IN9v6ePsJrkhq+g01JGpHyXv6cD8VRKHBn1u2V
10EiDpFbvj6lon3DdvEqMgvMy6iFWrPhAe08dZJhOtClXE83YbZB2kDk4sbyqn3W
+BuMSn+QNoOolBEe5vmHU14PJiHtv+/+f6tLIKY5wEwdZJB1ZdD4GSLwL0XkTfFM
RcqY3Sti+eCP/OH3i0fw2pYeXRshXXUmqslqpqzmv2LemT/SNBa22vHrtjhBVbCX
7P0lw466K1Yp3gxWd4Pp6ePXrXArtDVkvNMESNWPVYcz3QW00qLD6QwH50o3vBPv
GEMua8bkg15Ym3oQKeymNh+9HhydcJjokFt8mdTmS7mtj5CB+x+xVHfsDtByPr2s
cC+B0/xqUo5u/ZqRDXsLPjtUBTZ/da2WJCPnHL7Hs9+NzNdirq9vGyPJ2rawqAsq
wcvFJooinEJR3L2SW9viWUXT7/55K8cltRA0hcFrrXjJOR4LkQSIBi7bMTACeatA
Xlx5LzPBDOCHoFMa9UJlBr+WAteiBE+qpLiAkjmcjJAJ1DFmRf9AwdwBXpp+NxnW
NAsQkjcaSQWw1QDcxrv6dSLQra7HfM8bEWPIAQmDLl1AcKQbTWmGxRv8856JfKJy
chAT9zg0nvLPW5VOYdZRQhKlinbNQEiLadqwJV/kns5vGnCu0VpuRUt7US9rMFH1
+iGW8ia/pD4Xz0e2MBJevBvi1DtEJryOWhKFzVi52t+9HZmADEafmOSJpGfQJau2
kZK5gTjgSeSVGIYYibYVQJWZ+RPMejVSRX0smA7PhheEo74R6SRQTP1suXFp1FxJ
67OpQSfu16bCx4lPvaD5gFgyelZegpuhEHSFTPenb5VTz2prdP1okXOSEO9UD89j
aZy4ekGqVG1JthtjN3z38zNGh402NI/UcwDDnfwiqcPHYr54lVGd7W8vr7B3uLIr
dI6sa4CK2ZDG4PABSD8gq4VHBK0P/D6wwsx3ha5YfXyHbSRlhp5Oqptz52AbiI6J
T4zbtMXr8IRnNIHjNnA3Aa5a/MPZnVehHh/MIOFvQ5MG+ybexZZuXLnvs+lcaHCN
7bpx1WXM/g5lLvkuww2jK3xutkaCxsBF2BHkHeZVVAv8YPduhBdJq2hIvwF69DXn
Q18y8lMDDjgmo3PpXUHzJxFsK7PYtB+/taNKzO9PnBrtXuD4IIXBftoICHrOfvdC
vaGBXpZ8ENLhr7i649Vf/LF5xZLJOFdZC6woNg3G49kBjUZVqQdJNG9WH6VX+jCM
caf7xaxNHvC2og2CbqV39N6eN8oajiBwyMwM0Ern41+Chs8AeUgg3l+jIQ68rORn
1MP7XCUsHOqj9NVVL17CyY2FYFtgNnV9jhfozpN4AYZMcDWt8H0iR5Gx12/UmQQC
7DdbO0/5wqoAfdQzG2rCtBySpAg2LADjdcni/OTYBQ9G+Tql+Yb/VA+jB7Dz8WRy
NJN7q4d+t+cGBqUdH1SftLo2y5fvgqzswICICvU61DXEOSSiER01I8SoipfcrVVe
ATfXxp9wJJ0F363XMco/Fl3GBGbSMQ1dAh2lJ/660P88B6sUtYpIxCgpllJ8ZwBh
uMyezal65jD38DGb7WSJi2UuMV+w6TulT7sM1/XLHX779ONuwJLVEm/YkaqivH/V
g3efabA8CvzdeOvqA0+Q4X3BnnntsqV7LWTZA7jDk76rO5CezjdiUFyCZ8/mpZGd
fH3oCKJA5M1LU8iFN/Tmz9D6EP9Qwzo7TcfGniR2zgimLj3elPBgazqmNWGDG6jW
kHWZuHeFe5kipEPlK0Kq7ntVA9Z/8B9lq4d2nvSrmyunI7at5uBPNuP16RICM1UC
423v3uaXtvCoPTCDQsS0fp4z0T8VP8pbQylwU6gnZyE3/TzHSxPag4EsutGex2AH
VMub9fFrFu9s3sq0jWNDHe9B9uad9rJ7aQ4lVNegTFP/vJH8F7Yw85axPyfEQz27
f3deDAglPCbWcTFlKIZx7RUofPrgiL28bmdND35F5D3s6w+ixSV4qjckHSSfa1q1
3CQqOOrzi0EsI3BymOF+YYP0h3fw5HTV1H7+NODG3l53jKNqexsdZGhfAUTkFx+2
nRxQwnAPyUMnQf8wtrx4rt3pp+lfoAyY+b4vFK3M2VmKz4H4HZCjFNHtZbNlahLw
a1iLxOEzNSiynNk/fs08gzXdLK8uCLLNj2GsQ766O/YFyVt5n0V7Qujw/UFtg0DE
D0QRj5TBeKBGVWFSvoUxuf8ZIPWG7CLMJ8G1EKcf++Nc9rBrOIRv4TBfazxOuAUP
gbBHzTjVniPH3PODcve03ARGipAUbn0dfPbJA+Yuj3uyCLiot9oZzxS+cxzFvfaq
z9TpzuaT4QftSjO/+Z7ZGOZRygH06IJVa6a8QMXfKkAQKsu0MroKoHu/+iFT89VI
AzBedXRhxMYrfq2PhHFnUiN4UlSlXTWjgq4ijVqsQpnVBrkiLMvvUmbYPu1GLq46
E1L95vpc1Bz3/lg0ydIdOnKKMiZGsJWFrJ+ugBzdMbbnnGz5p2nnvbGtykdNMr9j
lK8NEcfARG0x5N2utyWu1+UbA46qP8rIT5m0ImeOpRGBPk/Pkb/jGVmdfTHBDYyb
7qkH4Zx6bxPFhCLuWwpPPVZli73Bf+dspah9EarJsBFxKxdDSbJq5aiC0w5i5Yyy
A+/+EK9MTMjLSCYmdtfUcc6KXIhqn65eQoYc+eqKoTX4/4EdOy/1cZop2H2qZsDC
mTNKLuyfjk790reFrUjMY9TBk+4VHj6IOcqUgExbf9jRFACLH1L1gfE13QVNFDch
bLxbo/YYNvdajOHXPr1cNu/29zuZGJCplK3iCftoT3OUWSY23DV0VfzRn7rzIKJe
9ZirUTehLOFzqRTHfPQmlQvjD7mImjkkD3kcE6j/SlO7KJuI3mQ1fYnUTeF2oyRd
b5kCu9i2wHCcykocBxYvvTmuRKqTpWn62sVl91QfG3HZLM1CkxeaYdpHcC/B6Kpi
fyRtJms1GRgSN+L1v9jk3bB1qjjaFp9K9h7iQNMtteD1z3ySNUsHLZDkfZrvK75H
j4/PRapxuDjRgA/6PZDiqkdXceX5lE+U9fHqT310aAltCoRcqHDwgI8RvApMpwf7
lkScQunfJ1gLBJs+c1ATSCrYBG3Z3aKd458C82UqpWYdWi4YMN8wegm3UymsIYXL
pTmJ1vBCSxq4Z/CO+LLHqVq8vAstsBzRA5sQohtXKypl2ZUt6i3ZBFzl6pF/VesV
AXsp3fErh6/0mTuPNrYRmxYh9n1jMjI1d2rLQyJBbHg/8/pSzjznawp1BfSQqVOg
dcFtBncrQioDLQAvjDZvLCuOGwhzTFQrhBDp1RBQ6ktFSVbGBCkqQ9gqFUwH7Erl
AxzYWQEPyUeDAWWGQuZjRZuaUjvxrw3TMWIM+5wMGOBWV9UEa7+18oiCZ2gbthkZ
QrNY8fUar6S2UsLjYQGPurye8af2c0RAPE9nOVwz220zC5hSLvzxMQgPYBuwlAxG
8wjkg9LId57ubpP9tbTeQzMX6/ZtL/lRMTW8vkM+11/U0/p5cNqlyKqEKevXwPE3
a7BUOcII5wg7A7Tk9TngCmveOg8iNZSQW6dY4HHkUSwzAc0nuyBTBF8HfMHVwwHU
oi8ZeYmannrKzXDqdGb0t56RD6IUYzR57iqBGvhVe9lUfXTzrxNFG9DYf6X9LTkO
MB880kW09gDQwyimYw+cRdEuC+ews5oBIstzkhsGcqWeCYSq96M21hAJabO4BYdS
NKWJnbi6xVj27RFdt7wcFLjwrslZdUGdOXv+o6l6H/RJb0KdxbQjrUT1OUi1hD7R
7zFA3k5z2vim1GR8LPV6oPYapzSSR32+26N1jFWuPjofEH5zCOGckmtGNTjhl6Wi
Z5VgW7dzHunCSvuiosRuk0h/9UD/AmpFEAuvAMq29UxFFY1sKVkxuU17m+dopkjA
coX0Ts2ebaezHT08xtjYeyekjOO79OTHLpqOUZezH0e8eNU0bG/qlUZyP9F6NQ6Y
x5wvU0sirPeWzN/B5uG7C59DaEjOYEYc9rI8b9UDSg49l9WUoNbxLbOdttt0gEFE
OF7n01QmkHcd39SJIqm2peuYhgJ2coISC6KExPLvI9e4r1nKScMKfMhd8NuFJf6a
4QFia5IPbbRtS6xDWDxhPlv+rUbeIyYca7Eik99cyUB7M6JHFd0MD6MBbzubYv9W
KWzRrWjJw4P7iaYMX70giyWtKPZJyAQFW0OJVTjVFE1w0QXSk3cY7TOOhz/2dPX/
isBZ7pQk5x39z49Uzl3UDqEF11PBB1vAypToOqw/EWQdh6TxCkuWyRKzs6KXx8iu
XrBu8wm/FrVWX2lX22JsFJFBRUX8rCZjLKxrD5OPUmpJU+VeUbnFiOXrV8zudxDo
k7+L+fQluWkjFOOxPE93IhGJSnV3Ytp9uWjOOgkBuwFUaXsm9nU6awon7sMk6Nqn
i46NwLZWSn3gwTnYbn4RlqahkBzKVSKnFGmaHhn3gwfn5z6y0pRQoEJJsGcJwVOK
qnO0YKlEc65kGujs9B1STDsIG7cx/UqO9vxLcz2n4NUP1qu+CevPN+B9Mr8PlaG2
OFfMt92UoAfEpU2F29G8Ukq1FArv4PfD6Et5ME1CEh8vJHryPuDdEx/5bjSxI8A3
a1sLqxUnEFUWhwPLj47eVcz2LpTY1FtI9zsIUHKQCnrsegt9NiRiLmibgIGfCFjN
9TAukcolnLtvU7kp/8E+AOfYWF7wZ8GxWw+KzPFs4SYpBdkoOGWcjcPvH5pQr+Ux
ctD+BIK/REck7qGi0x3rAqizXeUViluCOZI+EnrzThhw8S1nhSZm/CgMXRS/nVw9
nxDR2UXS5wf1HSd+YsdjtB/TPz+Rg/oQG+jJHtoEaJpPr/tMqZVF4q5uKjz3ZoU+
84XbtMAH2GfzHxB2P0IJA2ALkArYVfp80zfb1pYE9kNDHLTX2W4Mvmg5Rq2j/EUs
ExTTENAoXWGzWxuK84ArH1S1sZTlG2Z6Ta0ZCBe0nNGS8hepK4EduwymzDlWu2yP
jDSmad6k/GTCZsQxk5I+KbmjIPgxop/IADea44vJc+MOxfyj28VdoSlEyZ14FA52
VqMF7R+/1RU7kijmpLcqhLhqX7j+v+H81iMXkKRUwIjCepKCQgjRhU8MlXurRZJM
vwe0XKW1aUd20cYMwl38QGmDnEgq8u2dYAVq+z+JjmvcPYw3mqxqf3bUW/UI/nxS
m+tMmJ1E4geUAOFZbuuLRzBvsbzHUh0MPuCmeqQuJl1kyPoxE8nj9GXfA11+m+mi
uW6zGB5N2S7ipH+hRr1hl/fLjMe7ZXgjedNe9k/iFp7zzS/XJUo7ayIbV19CJfJC
qe+kIghGU/Vr1NNsW82ppY5wEdTymmnchRjyKLnW4udLu7Xn4D3csBzS7MXcObMc
P2mFGIGU/t/PVIBjYz790Rm6Vos3EN1jOWmJlnedy2DEW8ZpFaaQaEy0QK3u9BOI
iP0CwjPep3/Uer5PUByA4vK0Lesqsa3WBnSMHxjMt7zxSiaPWrZgt/KNoKCdoHTd
2hkcNW4XaWz1dGdEKHAF+6AwHslhXnhSD2apZkrSI70hfZHT3XNWcldubTAKNxdT
bRLj6PZ93y1PnD9u5IV1mQ68PNpoNBdHSRROhQFgI+kfN4Tku2hEgRnWdq/oY+9A
NhV+4P59BRMUjCm1x7fN1Lc7/B5TEERGBOgFNjwCzhW1k8Zbif1OPpNL6Mx8Hpu9
791tm1ZW5OxWXtAM3aT/Bl5IOD76L1xS4nTAct0T/o1pSPI6ZFqTieasH6H2mNfg
Oj+sfAKst6l8XqDVIIZYB9Uu/emgZJkpnrD9hRHobS7Rl/oC5PGsgoCdakCdB+nl
VbBbQb8X6cN8oijEffxAIB/uVGJrmHZ2zPCxfDK2i8aSptygrOoNWO8gowmefW3o
q4ZpIwUdysgUIUQnZp7M+oViykXZdPD+g84t9An6hIwCB+MtOrBD/rLRYHTR0i8C
ldcPKtJhwSlwFZZj475ygUa4Ktwft+uOXeCTANijfPXeywAA/M6Lpm44o+l597CA
hkbZraHD14mUN6mBWo9NGuKoWFbFShnoMYuWh2z9nUPOBoARnJjAokwp1k5j824X
BIAfHcyPFWBI6ZlLvJQRAlpz3tZ35/rj5aQ56NEVvTPNIknqK2xeNxZ2DPKssUXM
IWxm+FKF3ShxUqsSCsLGOg4yDgKL+1aoXzM6Ifvc5QxsETKqxMfKiTnp2Q1MEuuY
Wv6jPCAVnGdop1YhBa5mVsRR2zv1nhZwY2I2DLTmdOx86eWYVODMJgN05dtE0CWk
DuSJi2qeq51oI7IZtJgYH6MHiv5+HLVdhzYxub0fCYNmsuAB2Q9SzJ1SEFJ7r7Gg
8Tehr8xLciDWYgUs3e3sPb0smhmvgNT1GHsdZuN18zwgSussb8pVx649ONwjH0es
Q4A9+Wo4RSLRzhYG5f37jLJD2ct2aWlDWievO46NIURJCoodwVj50Sl8DDnE1hzr
GW5lmsXhq/860T0IN760wj7IB+DjbMU47GMgb3Z+R7Vo2aPlg1aWq2m2A6/ubT3+
8akwlTUBJkrKaBXVofVL+OWodcXXOwRCpfkWm4zLce3U/L5JHSEd5Dd8nJIg12su
iefGeZTrjYSVA4WmKDrX5ZUbZpJGGX/vV1dIM1f/V5SBJxP1oKEQBAopRftof2i7
ZP5DMD29ZxKsA2VR6/IIfLtKIz0OjTvMv3HUdG6IuXCJ+tvwrfyGe92rSP3l5KVW
LgvAixg8JpYil2GF+FZLIeqgmHrR560ukSXFIl1S3KVKf0TFCmXe9PX36caOZ9f3
rVxcY6Y3vrIQlPRsXqmj9avMN3XqeS/RQd5dfVGBOJr4i4pg4wjyyqo6E1h1MaJR
PoKxtGjJW/ugcvs/VSDq7bFpZsi2T0mC+RjyDF8/D3qjMDLi5JZKW42kaLNjhmCg
3l1CmSsLpJpCoF0jGvamBctatRjh5rWgy62t4QYTfHWZmzZH05z6sxRlWQamP4Ul
oTJSyix07NjIAmz3pkJA7ud7+qDkBAmAOLQ7/TZNXBTqMM9H4njb0baYNUCipXwK
6474lx4ubPJqzpOGfecEE58vUTLFuf8LSLv2yWyq9OkFfyl3wvA+LpXDm5KHDAQ9
PJN6J6eFxq+dCh1H5ks2PvK72PZfd5PL2S7c3x16wC/xfcRWS8Oop7kfyNczGyuP
EmBYKjqpFCjbOV23Ki9W3OzrnOgLhVYEjDnt2GqI2PlbwPFBGyjpci3APhvoA+HU
b9ehQzAGNFK2UF0ihbmISximP4NErUtzYa44IvR6Q2KhudIahMqEvLskwbgkpts6
DO8BmP6p5eVJs1Bxl864MJcX7lCGiGDi3Fh1wmJoipIONcmuZ941znPaxe2AKjp7
FRdj/G2QFLSZsyqiV5mzW41yLbO5qcT3go/Jyusnupb4pVaNFIWcoo7dsXIMZfss
TRi7tWR7NKS54ARxE56YX41HIGPWlUW5p01Ju3ur1yBtu5owhCx4X/N2PzSuu0O0
xjnkA6m445yJIF9WeD6Fz+/yr8uah0tJ6JsYqURyl6klfkH2G8Gh7iYxEw+9ixDl
ofvOwUxznJjoq96q1TNXACR+2/8j40yymX3j21W5oRKLZzxt9jQR1hQBg5iOe6Hq
moKDxvRdnVd1r3+oboKHtISw83F/+EKO6mzhPGYQv0SCmHQa/82vjcxAH1pgVKf6
ONO6ATeC1wspZadPvmWj9epsCTKm1VvxKWynVS45J5LfQy7fw43C6zmg6aidraIm
uC5syrZgt8/RTOtEk75DNrPMBMrph575fikAByKWt0sXM9/f4uILk0lv3BJ/Z89v
2SJ6M7nZaSJiXzSkm/SbNiVihnO7ySqpQA9wEep4wT3dSNvQ8EFtoztx9fvgiaCt
doHPs1+1MtYKHs8vIWTre80YbY2bJMO621fuLtEOELitxsAwazA58GEWOIuhMnN2
ZCnZD6EQZoMdWv/2vX7+V+DiIWzVtaCJvdvReMLHU2KGtFT+gYYsxfNkBQKKC95J
BqsuqtXNYcyKeLB27G40N1a2GxhthSB8gqs8fWVlQ8MyM3RNfvFztFCTm/LBOvjS
q2qsL0INIjM2Q6COQCrPOzrbdIKuaY7uJyQsezS1QY6wHVfKOinDYBV7YWpUaoSA
Fh3DaWyxgkgx3h2UdHUGTKpn1eu/YsSBZ7jFytt1Ndm+/fXskcWcZSernUtToQB5
bghByMvAZAq79rZWt1uH8dCTd2xAJyXlWBgDoWwkp5nh4Y8B7izlPkC9MSXjjlfA
HmCNRuwUc+iYNuUC3TrQAgYVEsoE83i+QLCfxs9EP942salrHHxpV+HSDOBerR9s
p6qITfC+PNTTOQfGyfy17ldTsWmHihlvRxQ+eg96M0hvTEtqNefOz+P8jOuzExqv
LR2pRezvAgo6XSUdJ3iGTv3pKaRBZzZSj+aNZadlXoBVELzyQwewKYnF0Wg6HHn1
pEg/iJG2kD/Xc8aSiB9OGxjA1iYnoA+yD2cXLRvK8i/blzOU7Nq2nAXv4iNXyOVC
LfCCEydSDvbqCBlgze1XVKZRRExYIMq7KlfhCDa0nc20tQB3xP4o0BGoMgB7e66/
MqFdAdpakP7Dwl1Nckfmg80iblQrg3rdwsfas6JOB9JNR7MkPqdX3eIJE5GqaCWn
8b+Rt9LZZWcRLwF18eW0Y0j+24QAVo+n0GRcPw7wBeizetLm/GeeYZneRqGmYW0z
7e0LMNBA8JdYFhOGamZFwYy00LgUyL9oiSxKlZhn/cIHIrZjWlsJPP2iHdRhzOtU
jdxnXLHQRMtjXhwwF62T8GCTn2gxPgLpzMp/uqjjlw8/DlxkX4GCY7x/d/emYc2L
SAUfVf93Xq2YZkpr5TpoSausePnHCWOaSoRY8kVWzPReTuVS80p/BQY7N4c520eF
BosyYhmRdhcX/JfCxbD6HXCkWdQBB8QH7pr6KGQLABvZRzdwICk/1bFUIaBRgcRX
WZNqg8t+Ft5JxAMTtzSUyo8yn5xS6ZkZ9XTc0oTk980uDpJGKfRrdCdqWeO2CuRp
uBVOmeno/Hqa2wBY8/8+MQh0/+bf5tYp1pSuQEaqDN4hxezRDTaxMVW0DLYnd2hZ
FLwLAB1rvI0IHR4q1gYlpJ94aqF+B//09iqItAqfSv5M7OUzTS2JxxJTgl/s3oJQ
2qgf3X+TJ/kRu1WuZPWISSMljwzzhro/EZ6s/4edZHqBnjHqiGpeXb8t4JKCbipg
BgNy00CU6k53wPWrMKq0tWQRv6GLefaUHeBzwQ4vS8mQpJ6olNX1tKjjDS/JUQ70
o1ku0ObGWoAgZasQH3uphssbybfSB8JweW/HFuvOyRi4CM/9EEbUafZNBF5ZuaJ2
JkFVC+EjM6bbVHocUKh+5FW0UH7bw+z3ncMrXcugG6Lgmsjhmo/BLDYwXVWovwUc
i+e2k3dCtoYnlzbJpN251R4KiFLn7cOxn9laRUSJ1vq7inWfAwi/PbIsLNSYQC6U
hvyCcaWQ82gy67IlyYRX/gKPdOQQXmUdyN29085WNto43P50hESyD4SybVMwi4fa
I0t45sWbPPtrtflA9K+Wq79g3Wu5ZdTQyao1Gmm8lvy2qdtH2tljMf3JEqPDPyAX
uwI6HfbiQBd0m26ic/uj3SoorBinyTHA5/Fbwd6nq8adAwwIz184dznR+K0xAJgY
jkPDelx07cBNwH4u21pwV4LirrvbgnhLdo7Rc/8Inkae2rIQjor8h9r7izHgZD2W
/RfSMXZO1hdTi3TeGtJdw14iTWHuPix8wm58gDp0l5i/FDFnnhoSgDiS4/DewPCD
JZOZDIhkljHrCSaJXbSQp+6g3V5ooOIB3pvh11rDdjoHbzmT5VemOi+QRFFXxlc8
LJ84urHGqi7/l4r1DkMpkUwv4c3SufnV+xP54ngt0Rpj3WMhvRTYeuzGCelU9OUJ
e/PP6RCngG+GAgJALPVAtFmi42IB99W2xIS0DKRRl2dDQPuS88Guylfz/b+Cr/Mh
XP2I6rzwP4HBCkLqWlFWjwR1Ul4ZtamdCdSuA1brxD9lZZOaQnMaIFBczOan9XT5
0jDmoEoQF48Um0+4nh53ovrbQiTdHHvQ/drq32aTLSp5ecqWjB5ttg0sD2pPSofW
XYkpquEnmco4HB32+zXatHKclqWiNQjoSa02B5FaA6DSAKlScOfAhvFl310w1ggy
dcf3zshil7uaKbWmtXPLp8E6fURdjObWfKDwBvpEFNIzJJ0gypJQKGX1h4s08p1R
kLKUiAEIEICdLUREAmAct+KmET15GjNJm4RuIoOjDrHxY6KrhCwR38YGNZh5gAjx
inFL7/FPQNU2DdyKPuto1nEd5pvz7TyMqhPQyRM8UCXE0ZGsrOPbbCFyW8kl7v0b
004G8p47FE8xKVp2JYsHbygilZCALskn+X18irdb8WvLqbBdCRf0IRGc9mqOTQQ8
gqX6yUUhevfKd5ZfDuAAFj+r0cFU1pKAwctoailkerJWW8konC+OMegXMx8oR3cB
wRYXK0ermkuZ9QhQnGtuuejdv7m5khOwCXlhJLmZ7tobkNjRDvObLJI2AHXUoV9Z
nKXwvwI+EmZSIkbx5UxX61HSd/54Zzs5yaEi00U1VEd1330i249eGQ6Gm8PCpFE5
tdGCdQCCzMINg2twnJh+wo6geoTjtvlc+rjDawWkbMW4HU9w0LFZcUFg/oPWefEJ
G924lPla9l4H0r/CWsGlFn8KNFTwsn/b3d29CKe94RizcX20L4IobvepsOIs0npm
OsTPfHvYtsfg12kkRcT750o/8Y+LzASpAm5uKz/xSAqj2aqNWgLHqa+rn2l1iqx4
tGnZMYIyHKlq44O1meXwqeFeHeWt/7wvOqeFCFMi/yc/vko6KvxpLHCb2ByB57il
1hbRpbxma+OR73lVfF9cDgjSHzWczm9tcp0QUjYUqgiVZpbDgPsnwz26x/8f76WI
IPCM8SPxHoW2urs54242X2Ou1YYZ+n5dxB5oQvh7OLlPwnxduVNK3u3VnRDpsV6g
numpd5O/yuFU3rdsG7dsVl5ovIcSdZaNHeCDwuparssst6x4cEVioyNn8ePMUtFK
2IxfU1bdUdE/K0luOHi3YkUEAQm9y+lG/h7zsQJVFWzlPJl9xgYV7svCgGltUY1E
lqou8Nk7pFcpqVquBZvAo5vgAetp7hJDHjgRQOaZcGCZBjX7Pz00qQMEKws/xTih
/3dQX1nMd9Q1FBp7WHvBFd1BAii2IXo5iJujEZ/OZEc4NS+3QCfD0mZngVOKzjiO
l6BjGJBDINcz9ig9GUQ9XpqScv9xSvFNGy/rtW00T+EHrxRWbtfuqHe8sfYF+Opd
hgwhJP7DsWXQSK9tA461gBuMEuKiPXzBJkUB1mQPBZYnEbUfxymwtK/9j3uE+FRp
FhOGO3f636AVQk9PssZowcAA38j1L14Gy4lH/6SO3Fu3JmR0v02lYKOtJ2lR5axo
Zge4X0MIqH0ftHTO3puwFnD9RoipcPeFRc605nSG/IoAL7JHDMrt7WA4ePAtcB/l
t8yugJ1TAeafDPGZEBpRgwSg9wG8R1IOGYirfoaT6d4pcxoCEaEyOdnIpXyNGZh9
ZPAJIkXZ6WNyWid49Sb2wojA25Etwy+H5y1AnlN8lsau7ISQS5uMziC4alsKhg24
LzWiss133AtiEgjnJEDXXnizuwjUqG7QPuwZN9AtxpCEjvwrEXjg3cVXwOAsJJI6
cpwRAMNlYdfUUPSgSAvmha8MET5eIWdrni3iCSa/L/hGGxQOijJygm9YdnpPzGKp
tt1wTsPCwvCsslAuqIxg6QPVoZarmhclQv+BTanteRBdw3vq8YNIl3mXM6exjFHa
Knyl27+UM1zficBxbQuY+o6GJ8nPyM6MRY5cT6wqvo/WBuTQufEG9J3nEaaZHwY2
VDUhz8ot4kwotnArEvufUCurZTDn5GrEUzqPn+jdq527iHDwSHnKxM6/vs0rV0y4
mUvnbb28YlK5jHDKnoFsEI0tVK+NUOkWXl6fZfAA3kO9mrf5mA34rlKcdp/Xe0rq
vT4ndWcBmsv2WmCbT/Hf0KJ/ycya9T5hpI4+0LdB3mj4HghXX8y8M4e6wwu4y1N9
/ZNXUSakNJx1CpgRRYppk9GI2R8V5x+5p7VlstaPQXKf/NAakqqrmgdKzkscJXnu
rX4qP91PnzT5zfIOL33hcE7QF49qtGLkhzR6gHb7tHnup2Th29dkybKYeoZAifMW
XWf9uCEvwSmO4sJBmqqVYEsrpTXBbLRq6SL8Z/9ldFOD07h0BVPXGBCwHnZgBabA
fMN4ecPuvoqkonz4cgksyW6JPwWnX1n6XIpKyjiuhmz41Z4uob2HRN4ur1KqK4W9
n+YeBKB9U/qkC0sr8tDKEi8W8KycNhmmUYNDYTGaCaYqet1rBshyjUrugalLpn+z
z5NmJkSpNObIj5FrVfHzd1KYCByxwhxAlCnC2l47Qm85ipHVMWwRAa7eIj0j+RLw
bni/JR2a6fdId/r0dw60xMfgUv1KVt/w2ydMxgJF5IyiBi5KzgOceDh9O5WNYcGH
CfLKKD2M1HX4FxayO8hz2okWvpKBnciwmwmnivSCIG3nvN367UOUO8YzoDkyj6qG
+ZhR8Ad+4taNAP3i5rIvw/5MuG4Fx7fuEOV123M9Cv2PgnXgaIKPhfl9mR/GzzP8
JMWpdZVt7rzw1HvdB+ckht98wuaGtV93SGaDpYpL3IjCqpSRGkoH1eB8m8N9Eg7z
hPjCx2ZIiOkCPbDErmt0zPgrEOdsax9jjLq4SdhdIn7m+1/D0tglrZIIiSj2QxOG
ezc6jHroc1tFd+lqJL2D2wGzlU9/pjJpoDS/t2cs7ETFzHRDLVCOiVBCoj4Rp5RQ
C4es2v7ASCl3c/GD6IKPZbEHS/2XLpjmsUVXIcLF3JLew2cdVw0GFLzzs/Qog56i
02ljiSiUvD09hQ2vTtWFqHM5pVlWdpkr1s4aqwJE0EKQURDG1Yt8dImzjP0/VKpy
1A5VIa7cHlFyUjgmMYa2TcUTEBisZ0k0kRSh/a99nOyqK6Q/vm7GvIZSSqivd6Mg
Uy0l5dHeAIGB1hMdn3hUz7rZ54dsLhhYDS15Ds2vEn+VEqsWX/j/ppdDoGC1X6oT
wPPld0/FL3UQTa1Y238E6Ce4i/BMp1ShNNJ1bQkvAIrTRRtcZcoSODCifprH3dD7
sQ1pq8BhX4HiAcap6NNq9XOG/UWJjuuVkkIsa+bBicecb4yZO43jFCBpjWDxLDt8
xr0ELTdt++wFpAuM7cvCAOQLdP9wwcHQtqfaJ2jRYGNztzNEn8w/m1pwrcjSuu9u
9tUThbolMab09eKd7DjXHrXu6wvoru78jGUzQhRuP1CGg0m5jKbe+F/397nEDnuI
s4+T4n6JNNuRF+Sw0HlrwkFv04DLc7r+BwxIGgNPA9QAlbZSC/oqP11YwWHPd1x0
ANoUFJgHOQlLDaPD19U1kB6bcRYQV6QczGCDS7KPp86URhXhOqBcrvW33LXlcfed
UFmYGaLR3kJix7SInUYf5IYOVMAZdcajluBeJhkyfV6Sp3kmu0w1NDNK4YaDcASz
S2HRwlEUqDcazkmWPN4x0qsI19qkapkVRVBstekdongElEy0HVK9tzsx8ULwEAdr
ypD3X1B1VGAODkqz2cyMUE8paiq7f9E5+fa9rm6oh80tfGvnj+FQ8tqkZcek0gO/
aZNG8O5oI+yDE+VlSDC62PcCjuGHyK92lzZU8kJcJr+cYMuClh/JPxgbBz98uR6s
jPi7CEbEdCGsIJ8hEuFJMJEiu0aJsQ2ZatiDE5Pfni2N9QuyB0HizrHnVFVJ0LP4
7z5AFgKhXCnoJl0Q3N7HQYgYFjR8d8VW0Z20ceA4jJydnHzo7XmEA/rnroCF6ZoA
eWZzzQ84TCiEi98tgseAApz2M9JMVzsNp2xnyQI8pgwIcgsRjnRCpaQrud+Bqnp3
fKbu1SYia3N3FlErfXj14iDoeWz3y2oALiBk+hLwR/6Pft3HQ/IhSrUxWK7VT7+m
DV83j5APjOK/GLwaeqEy/+PFZ33d3AKdjHY0GfMqMe+kVsPr07ZsFDQ/ZWaWS/N4
p9FIHJeqDFXmI69Ap/Neg/N7wjLMn8VOvuOSHq+DLFSFrBYITsXDfXl70hMjoV37
zf/Fqr3qjS25N1vUfWlOWsGdVqoQXJfFd4xHn7d8D8WmLAXRB77DJpfYT4XWIzBz
7MfEtwgFZVvtS+4EjdN8hfjVQZjpdn56QOOOsyhJk6VzLJzaoTpzy3XTjmqBWCIF
2CxSp4KC/kcwUSgMoCw4zl7SR8n3wWW9935/fCGKX3b4pm9NCrRdy4b4MWrjqXj+
ZoKhhpJXWvHmpyw1Uy0KesbAElgEnl1EO32QdHdfU52qhvTag2IVlysiIshi3DHR
DtFeSnyc+PLZVntvTHmZGKUSMLDABrE4fN7IEBk7gcYIbqrcyFF3ppR4TQTLeGQd
y58Uyo6g7vdst60PFYBfypF9D+/bSSNIp5wBCI1MDocFjrDWra+/t0dfhtlK5d0A
M9kNUDb8k0fDMjN8ZL6DUtrZlLZDsJllpjRwnq86XMIZ4v3cL5ZrpI2j7GTefbG8
aUL4v37mumKh+YD//UbHCewQ8JaWx9Qyq0n6Oby/sbOkDZlA4qTvB4PaHvR8/t9h
cQHZjY2Bdcm+MSjRDikOx7ote87E47ZuWeifMHno/CcP1CMMDuj+8QnrbU/VPCVz
ED2NAQ5xF6i4SCbhPNrGKhYDbufUUj8UFJz5nGfaQQbpMgA4iLxohJBq+iddFM7H
W/qR1R7TfHPpYbE7adUdLaxhnpMSLlPyWNwBPRG4wEPqVjpuBoHpDPETmrZqnWkb
fuOt6/CQKjo/dvrXJvQWBDDLwlQCaJIQfeKaoaASZ9wNiNgHEBnVVS4/obNXNmJj
UQv0xcXP4DIoVNTXJwE6Y0C/SlQL47NGEKSj7S3AI0MsXupEbKeJykG4uUTG0q8W
EhWaKOQ07UW0j6/VEyhZqgEctf4PyslCIeBTUArNt/ZtL8vtFRf3gosNE/5ykO4v
QaI06DX8S77kzre3/4z7gLP+Cl3TrcuxbY7usx+rBX5XIjXlG2aA3ux3klEFYuxh
vlciSsPl1zYQLaBkJw4fMq5Coasoe7fRbXhPQz8Q0MeLCD010x8yT8b4Cr/arw6R
TMfqhgVaYjnzamMOIPEApCMPJpQ7G96kJtSOi4dK9hhuqmiwsYxhEhs+06o7bsD9
5IBkh/M46VXMuXveV3s0qKZZy3t/PHmk3qnmm7ydVvmxVpldmSk7nOhZ5yKIq5cZ
DeE/xSi4GLaHSZLLi62WMrUfsFnSXF3Ss4InywD0VFzW0KkeScQqNrjTyCHBn5+e
uKWvtEGxZtJiIAmRQDBIAXMqG4jmUrS/B5sCeHZXEH0Cq91lPAR9/8zz6NZQp1Yw
T6f7UV7a4LhoG+0V+M+dMo1UIA6zBVDOoDaKsp+5HsFkZuNkddPcY8wSb6x9ErMo
eFVfPLgOMsLaeTEMIpTauGDTZGMeQn+7sLqVRDbbj6vtU3AGGoszdfW9h0TLbZ0g
UnjFVM5Agx7jT0B8zu1TNpcUEmpjvkVBpwcWVituAdZb3CzTzkIFT1i5RmVHkr3N
VFzwj2FEONl1w6lmgNi0++lILJpgcZFfHQchVh0/RKu2H4C0ku1mD14hgMs73Rk9
68S75cK+uTqirGq75VkPnWJJHoBxPS3E/UZ++tXosBKCJRsrcFUlNf+xeq+eW180
pzZDfe8Ha//L0eudLnmYc3USZ++3TazG0JTVNnYbAvoQ3k6sp3LJZYEHqq9E9aoN
wvw9egTUjcPnar1m3giGY9I9+MmcwVgSEG5kaielwzs6kFTo1dNU2fm0AQy8sOA2
ezsBEwDOS9VexW/GyKYZFhv2wBrigre/EIvdV2Lgjd7/08dO4JtV6Q8Yr3/9wGIO
k/75XcGBFCpaihMO5+OW9kFPP/DrtMNQpE/NS4UPm7ZQveJCW63TUUKGx59Gh5Vk
GPcmw121g+HpZ3vHSq3kfbTdMunx9Z299unBsHdyxSHDMUi4hhkM+TTWJ02PhIYR
dlM418JR6G2tDWssIbMPeqEE1FneYdOkVE17ZqIoRKZ60DXmYG1WX3nR0u2BYKhj
+E4rehk7SVb1+nAzId1Uns9EZNz66R0movHYtoXDsjIcZ/jVsnoNkOyYd8uCadfR
6TvB6J53NXRCVBqQoHqTIym7sSScNrhiAtVmxqKRjW93eaiaMpEqq3YTdm0BGIHT
YAvNWSiNb7QRJGOajn5nFV6rM5dxDpf+8jbwGBGTjIEPqmO5vx4Y2jwkh3/opI8G
loBiTS0Czp1a4ZIP3swBeVVzv54dQ5ZPNl3sr+5TVEUnPW67YNuk6+4ENBW19S83
obbnf9KAtShXKyHxsjsWfkoMtB85u7ziK6MKlofSBngrHWSTIjsiCvjsKd16qG1+
YJCfls5YKZerirjkcCdVF2Jhww/IiiuJpPIV+BCW2JGkvqx0bms4+MTyVYuSp04z
VV/ZY2CtQUwkxN2l2tcgYwiJvUIvBxJNH82tn7jE/22mzNAZKnNKjfWEbryC1nsX
tlLaxk9fAfhNA+VpZtwvyQ+NwwA6O2I5iXAbkcfNf+dxHKgz8RJxBMXO/k9GEZL4
GkPTrmrGHEKPLpt4X34Q7HzMkYadvpFEhpB7YFQjRys4qiEjqfZA57EahhXguSPB
e2VEkdArHRIqDLIw37cobpF7sfaVlkOzmZQ0E8CuwLwqG+wME1ij5WHCvUh1ls4j
dXUC3sIbmeI/DJL2Lgg0EJKPxlyr01XeIY+FKl9JM9gf6B9XA6NQVu8e/d0p7Ir/
N6BmPYtFIQgnM6aQOVQkv8dUFz0aL7ZDolNTBh9Cosj+I2i/aNJcM5BQgf6idt2g
uvzLK7+tN6GHmpl42n/9ADyojNV6cyvy5myAL6SeQniQgKI4uu2fyvR3NbmI/iY2
4FXk5oRh+eSbUljTlSPwDQoT3WnKpXo265te5zhv0RGsiwXMIBH8u+uucHwxxnz2
+xsXY+wNbb/3nhon+fmClS7/uk/yAEIz3dh34TZNhA73eHMXL5rPigy/zRjWz4P/
syngnqc6QQ90raI3nWr/osWI7sGWWgUB7YfL928vumEUQVLpoAt2KKdTzb3NhZEE
x4Hd1PomxCOCmk7q0ez5iRkvbsavzvVDvEO48TGKwzec9IOWaL7oDgOfBSeEZ4Um
z0EGXrjdmXGd6KsThvetjsafodPSk9AynWEFdQt9tpi0nq2KOttrPlUhWD4eojXA
UCNIbWoGsupU/P5G5ENW/N5RynqkRP0+T8yu4OL0by/+G3jbp+OqDQdweaFgGfQm
oa5IrqQMVFKy8Hc7lI7/+NVce1L6XS3U+QS6N4DHaEWtwdoXuASc+4d1VmfPcPm5
FlTzZsGRvRvCxA96W3t6NAK2syEB09PuS8bvp0J8Fy/yRzQahsQthtuk1a0nVvT7
RPSl8a31BVCRfBJ17CUgcq3QuGY6cGppH1P+dD8JpUKD1gtQyp+mTFX8K652CI2m
MWFms/ypibxX19eCD8TwNR/AUQcWOMEZylBr+0nCcrpgRxwJ/fpRQ5le91efzEoB
1th4iz8LJbhLanrM9rofcphL/jP45lQDngZbyE3byiN6tS+gpNxhw+icTXvGidCe
QoD6hcxS5vLAdyMo3h1gm6CwQkFNeiepoFGtbW2kLhKxjZbxQb1tX+fkKYDIfpIB
f3iocckvC5wSOM9uqvVuGgzwMFb6RDpD23yBwDBumhU3AP/CEtPFJqSnXEBSA0HK
RxbbJA9FB8nqxRokl9KHNuQlTGPhmy8n2jdWebty49WTFOxDnzaCHjFOOshQWC0w
jPn3uq0cwhpGPf6yicyMnco/XnXKaSLL0A+KnmCPau2VUz55vqAn+eh0Ahtf6IBJ
C2mpNJnCV30f83i2vm7madymTrmssuvZYlSvdhofuXEbNeODVuFJU12PP99MXp3+
0BN744aWTVQ5rIa+O1+Y2vCukyTf5Ib8jjxhHqRJCgCOvUtT5gVWa7n3eHSD0hPN
EXxdDHUduN6DYv7nqxXGT9wuG30vM3gDL6EO4WsQLJaT6PqE8zSvCuke26ZBe9jD
G95IDVj+K2FWhQANthlMSMY/wOvJ/ZDEogD8LsETHmJ9ouy09yjm6nO/KmB9Js0W
wXm0Ur4V/PklFEVXfeWitdrD2/DTBUSFec7q9xIcCYDBP9f0kaO+fHNlwgIZK9jp
reZAmEg3nziihipO1iuzL/NMH6Sn7BbWxhcn1jy2UR5HOg+0ZPXjnB4XqMc63EIF
+I6yAVe9WDhJKkh2kCl4Iz9FU0n1g97GCcoNQRy3tbiHs4pTToB3TDvJtTzQuScQ
mWJZhQC4/sEANytMiUVvTssuTe7wxjwy+DbPpCSyYUYdzgJlDxRya9EujlbOSwMD
NHL+cjaAl9O1CCHcu3HakPaPwcZpPBqH7RlxeWEJk0rb8wfE0t3l9S9EHPOdd5u3
ESqDE5Vhv0qZA4yyQO0IJ9gS2zjLSpe4WtFUw7z8xE8GsUrQfJJq7iWd27qi4T6C
hfmEcQxgE27Uyz/YPh5WLXJ3k49n/BV8j/L0BUxBGhwTiJ11aTKUD3P2JCnqCA9/
Lt0avaF52V9unzD4DEhJ294R88XgSDQFC1qzFlybu2Fycl6U29U+QFlJ7poggrin
dsIarp46zzOagd7nFKCxAIr42CMPKzflWTqU+OLd1XVBhGNzADYJfzOK4DeYoPcE
u/sGn1GSzI0KQxbazJxF7ngGvl42QzpKPcoDxAV2PAHqLjbxf3P8eK3e5KHmP5FX
5G6/HJbQwEDscFabu2ANfMrlldXHKeoH4JGJjJbDgpdAY4dYt68kfG61Nv57RuVm
C6tkR232Qe/1kOFDafolLBAo1ysaW8hNu0RolMCq+eai//FCaeRUO4wdCmkZYkcl
+RN+sfjgo1VGQgiWXqCNtioK5iZqvdR3UqyhIef/UxSmrUYfgJJM4/WxJZ2f/xmv
iP0J8hEN/vKYPLpXSpE/OpoQujU4FJ0kaR14gOLZg0gGV+BCHAaEBRCLYzuEb/nt
gjZ1zYcacndzfQEspY/litjALhJt99Idi3R1bjreIpj86Cfk/4x5xXTzjExadxvo
qq8N0yPd7navqvUOn6s61F5kBgggyzuRbyhc5MQkwh+Lc2FEXcpa73fg0BhlV/Nk
qqooEzXIq1th8bnKO8WA1WSbPS2JQ4TAlNXnJpQR4tW9Wi+B7bJDny5uPVzDRDbo
gcXFebQIbosPfcmXsmT+Drqj1qCvc97TEgh4yBvr90ihH4f5PoPS0DhtAYwXjJQM
+IRovf69ca9lHP58DuDrd9xeVOK5/bSk3jZaXkOvJfIP1h1KRzmbDtat5f7rx3xl
KyrQzB7kzhi1+Nus6AMKUra6pTk9vnGx84UJ+T3ujuMjWlaEo0UpeTvXyjRIout0
OfjfLyLSKR9Di4kgwVxN3pGPLEYgkDWxrlNYtAl5A+7/HSMsGe1t5qqh8covjfRu
I/FheHjp+IAnK3HXow2EUMCqnnie5Uha/IBDjngiQhJNcLFYVdauxjkc+vxzgqPF
rPetgR8f5rQ2nGs6USkj+oxjzz5ZoAkB8KmU1a6Yz22SJYL09J8k76AJGsjbK51q
BdbRYfQtGTWx4hDyXoHoPa3GfYU1Co6f6E4RLwp73JiIqIioBJL+zvwvG0rPwXuZ
wiZ7QmfjBkjlEXmPB9wdD2KNK73NVOlThwk4JBCVIJJaEX2Q9sMlrGwa2m6IccRf
mYRFyacxqo6Rr+jKfF1p3BpPpdr6pJQ/pN3lS8Pkljltv/edQcSQb6d+j5jtQ82Y
QzxR+8byZaTvJJ2pR9KFJ5D/I3X5whmcn10sMlbiZdNme3AIM8fGEalM8QL2dwvj
SEfR5JJVJ07/g4xo1pM8W4dDtz6GGSHJCZja25yz2v6eQTEvYLB0YCGjQngSq6AJ
e0Ou7d9fL6mKhZ15G0lMWolxghi7MGJF4VAtQPwQiykv0z8DM0wkTzDF9tOZxU3z
rRAlOXOTQniwQtWwMqCAMXGfT8HOH3Nk/8O5ZHJJrRfh9ta2I5aWVVRy4fDU37tf
UnC1WLjyUbzxkXIbuW1WU8ZP3VjGLdQ6oC+E/rmKD6OBUO5ktI82Tt5Ki+sVAFHm
lwSnlWEMZz7ziSi9OCN8GTQYbCVs9/q5lysXVOsnryzMXKfnWsxpCxLJQHHPAR0n
VQ5wW7mWVZa0UbD9yXaJS9gnZihS+056OBneP/iLDogsGLWEyNHqoQNAekodK50V
o2wSybcIRFhkfS5/jsk6wgYoaRxLDloN8fSzWieyzg96Ct7IEOt/SZrn3QmMfhmH
AY0lyZ1yNViq7Ih3vxEzvMZCsaB0U/bVLKyHKJOqNIRDAWfv2Y0dqEdG5g0PJSuc
POoIp24UfKJUGHWnetK/CTrGP7leaDXCpoF8TQMlv4yuE2Od8yMDM4m8botIslUq
TiIoMP/iUdoptXqbL8gBVpksQMA1LMRlVjCtb1RJImFi3VEaou6VsS31Kb9OWWOe
MaOw9Jo03Pippjm/iPRRbtE1rj0OtlzLWHFMQ2ha7Fz+XoncPiM2YKVvvjaCL14M
l+I8KiJrZWTznyLh7s/nSb4DTanutzR9ZtQWdV/bcD4bve1VyVvcRJCUpquy6Ih9
n09sg5RDTBJoAiqZaX4gCrCV6dvm4y+RzHS33PRvUpzsliQypny5f7Z1bJlmlMME
YavSoT9PU/GarfCTJd1eqwEJXjSxuKjuFpb/e6FG6VGwUTq+P7kb0BK+iAS/h/ch
ICtNLeVBhOdu7k88zAgB+6PeL7sifIKWJGSVWsX2P4InUPLY0eW+1ZRWqAKhC3gu
d925aXZS52VxR4K2ZWuMqAEKfLFCymqmapI/bcX3Ks0oj1qwLlVCo5h+DLKOQfcx
JpGUUOoPQf1EJc+45AVQ5QmXETT1kAcm/Wu0wuKAZo3jUKk3gkUAiXYfANoxeJSh
r7jUTxWAfxHxx/fNpoHYyy/Si2dt1IBe8kTJdecYYz4GV1uhDpa4ulxT74pZoHGp
FZbJHaPbEXtUhClNxPVyRqkxm9ekKzLwi65k9WbWwD7+tU3dlUsvVCxNXYtwy7FQ
45rJfTMls8db78iNwvxhOipcgoFvdDuWjsaiLNy/D8dlIB6eFJxGVo67QMqJEhoj
0UCudXaaA+dBlRkhZ1kteid4k1zrYFjNNUYaQdVN0Y7UKMawahrcgZRqpMWViVoK
LR7YJ9cDGuZLCUELJ7UBjsfrhBrKVrq+Qb7TZjbPTESuRxQLo8rmyX2a4CYzCZCG
ef5UlByIO/XTsfd4jYmRZTgSvpaHpGvVtsTgUbXh9vU+v7MET2P8xCQRVbJr2q45
M8uGTzfZf8HKL0hsNZg3oid05s/bey49gCPkoD0ogFDfiFus9zmLleMKwr+WqmLR
WFblBIXp438OKa89CuXe4HHKRjWmVpy6/tCWKbOf/RDdanWAkQqdgcxL4HrowDaq
iiz7iOEzqHz+4+We52oRSdsNu2MS+V1tp9SBxEYq8I+rh6FxZccfue0iF+lr9dXq
+3q7D8kvuoK0kgWvV9/TAfziBL2ICxoW6LbXE4AIGGeCjeZiVitORjD4+N1MvVcQ
93fvpegoOTXfTuD0vM/1PTplE5O4rYSnqZ2r6siRcyRjwjEwRYa1YMlaOml5dvx4
OG//w7i3OCdg8O0VP0igTGTl4sTu1jRzobif8o1dN33dYXInk5+j6n2roI1ONH45
SlvWTEF2TVkzFIovPXQmt/v2DcJhx43Aa4FV0AKPBVMZUUuS/bFHJ+UV7LVwFbHi
3m3wJtGdCFAkpfCqkasD/5pfmW+w+X6P9nd9doYu2Tpm5ieMz+HcYLvN1PWb4CMV
OQJo9Q9FLXEkPUgaal1jTNqbU4ALg/HFRj8uGjwPOcSiKqqh3tcbXVB9q253W37x
oJflw+Nq/AIYnbI6VDUrA4cOGvzA8QXEe13GmABQZJoWa669bdJpP+fPXwDgzYjo
wU2u2pa6RZ1/9S7tnN+O95Bfrk0HEAObeEbzFuOuzfe24MRq6IBlK1yt4+xopsnt
Gf4uHnZXGvteTN5cVjem6HlcTIBkspdyhXDcGjqT3tqmOR31JxhZ40Utbzqy3dUJ
NPEfhzWrUagqySwKvpM9fNEF/nuoJX/7QQXKeRRo+DXetv1NUVKPL4YxIGYXzzZs
gYS3kU7IiyLbddwHbPwiTP1RsA4Ac4XLTVo54LJHWUO+A4nvED/5VmnNQ526DDV5
DVDibwKz4VtJ7hc2ycJNIfkYJerS5zVjYsUTG/bqmkE1fTpdOZZ9sZUYOAlSvRNY
TrXLaeqhXim6mrB5t+RgsjiM1GkP9+C8TMC0yKYtzKnh6MgWR+NRAs46+OBiAI5b
bX7lVIIuEePY8WMKzMFHyXu6X42o/YjW6YsWyh1N6Z0pQFVOxxG8SetspW5f2Mmn
xgy/OprpDkqwb9EHRdYQx3SC947a2b7nJn7jVxoc//8JdNa1Utc5yGMgSdb9yZsv
qOVAoJekUbDwaRKythe1hexQbIsUnqlMz/3s4zby43XIvklGQDDFQz3c6uavBvzV
T4wrnr5oL+xWhuyr5Gf7fnsJWmcTbf9X4WcZD8qGm9x6Aie8Cyz6rj0CQI+6V3z6
mahLs/asg2GQCfofb9KgpMoX8mtCM7xu1t1VBRqQQ5qKjhEQe6X3nspE4RERjU8Y
UijojuSP8ERx4mnM71feddIhKJWTXJCwZ6Nn3QRXI1ChpLm2SAC2Z1y/0Ytq9au4
I1cmBkfXNAF9iLHYS7p++HoBb6GByiV62RiHF/355Ad7LtFDibG8HEPBX6aaTOzb
iTzcrQKOWmMgxFolA4PwtJzX7f87aZEPop0zcwDerBKu5/pwU9JNtTEhiarvoxRl
RtzdsIrLWg8JP+jw6Mmer+1jwD3ZkMQ4aFJwZIjf0GESnlWYrsr5XKq8BZO+iCzw
iq7R2eWgI35a3l7XI0tLnFu5kY+ebwPZt9LppqxjeiBfEH8J+e54MZ1n8tKOrlWP
HNQxQehhXsUZ90R2UZI5ahIZ/bptaksIlGZ6rHHJRaqCQsiPhCOv8gnXQMhrlT+v
w6KfF7qMi/MmayoRZ6XTTg7QzP+wP6c4Y52lG1PXtid/th7DIWG5mf+9q/gRphrm
Y6CnHpClXoLxSJAJwKfxktuxlxY1X9TcYautOy+PO84B6lmAsSuZocuvIakgcLw3
liFTul8kyNEDwNHylYf5tYzOG9WOtJD8mRAsBTGnI9sPH9tRDP5a8n923zCP/Lha
SjqW9MhffR47TqpQZLE2hfjY/fs4eUrMCzlgkMIGqFMX+EB6qCo3Wk85YaljGghV
bp/gb+7iI+vOR6KJm039OPPOawdEsKm7CAzFnmGEQLJD0urfqyGmo9CimNqAW5Zg
9Rjmina3gWif50WNVoKu9jAWozSF6uAmcGJ/PbhhO9CBVn4jfRtEpf70dOd++wC5
MNKe9AkqoT5Gz5KdLOJdqAZP2zo2YPQhfKGlSS42iBc1PKRz126kythAR6IM+HEc
gGQ1PLo2/C0mqdwZaypd5MkdBOq+sKAxVZpTgVqtuZe04MxVcqbXf076MbVvlRo+
jRIRUJxyUMUOekzmJMgspNy4pEhBrZ7r2T8+vrhN5QDQYuQEUpQ82D5cCK8DTVR5
LLMaldPlb2rUCSFA+SCHpdfsZjR9B9q7oEmqKwLttY2IOzy7xByulL4peRaQG/Sj
IxfuLXeR5Jk2AjuBobBspLB3g2jwVVBpjeln2tTVebqnwBK7aeZEnl5E3kUrscU7
hoADqSXBpKECnZp3qOB4ZW2+6+GW2sKHMcJvwwTx7jqikbodzCJW9l0WNVrzDxwL
vvk3eo9BORba65cHku6u02ClYq0Cx5T1q02pJ3I6MgNJA2f7TTc4dmJ3BNf5OE0I
tUk+9xlC8+WrZdV54b9odJ3+sni7pLdDhsxBWVd2p20YQEkk59VeJ39CHiGw6hML
QvO6u2/9gOzwwPIPESz1DI1otfE0qEyq7YUuiDLdpS6V0oCmZLGSrPueizNEjqye
n4YTUQNTNakDYwKhigHtuuLTyAe7dwo8P/Oo7MgAyQ+KjmX9Prw+I05yyjzJk2yP
FiEvyUnqkp+hkiSYKoqA9kAHRjBQJL5MxSqdga4xKs/kOAAt9+I1dnLkEFdndavl
2yTmHCwzLa/4Bx7l6Jmn8JeSFq3CC4qX04G98EbWWDEPWZtUTGIkkDpcCI75vEZv
binLMfLup9D6+2Wh+9To1tFpbL07hDrCo5pRmXj2lS6Ezrhw1dgWAStifKCbj3W7
T43RJtvjDWOw++jqi7LruCeM5IptUPVjnGj+QzJSH+5KmftF9XpMyZbkjobK8bFQ
/TRankHaps+mv9Ic3yf+S/GHLWHUWmQuzQmhKF/YrS7dAjMsY+E+GkYEMnqGyUh0
tEjmejd9vzl/U9W5oJZe1JyNfBQJm1fLasoaA5totbXXJXZ4AasfJrCbYd7lBoF3
m10i5CClu7tARI2G5Ek1LEhiNUCnq3+dnvTyE8VkyfMgTGME8ChYyqzui1IA7M5e
qY/H19wM3x3vMB9ibeGln04fQiqMs4AzZHGQK14jgveBzjrLuaaxRpH9eDc74Ydw
ym0/cKaPloX8BO2eNV9OGkgC2n/XhR78HB7bHomWjY94ep1FNIB7FeFdDyph49Jq
qiMQq/gMvJ13a72gH109cK8ztl93HuSxtgYrIeN6egyDVZ9AMhMkdQU4tuJdUi+F
5otu7ATu9gggPNWCe5NeJ5T8wL2vw2C7LbGdYVq+FH54McnRwXwfu+rXdQHGqbn8
SElV7GAAtv6OgMkZHbV1XUSVq5bPiGtteo43iTIYywsXUOAv07DWxINFH3GLK0bX
5oPo/Dizk0cBV/qm79y902t1hAcP7fBW7pxHXiCcp4Xbw+hFAU9enk4orjNprnFj
pLekvR2J86a72LLO2QqrDc7cgvNBL0jjJJclBw2ZPBC2zCv/ytjGT0fxWPynKEuj
kY21VKIM53kIGtcZ/33CJ4zaEo8MSod61MfdjQy/SevlzjzO0ZpyLs6ZLKwgDE3d
VtriEgFqJfe5oFr2CeZ3slBe/0PJN5hTgl8sK9Cwjfea9DzI5GFoCVyyxGlNVJj7
iYfbAmbX+G+2IQ0zl5tcNS++SLaCicvswE59guRI/Lz0ZgpcFtsu/83YUjnxvO3N
mxcZfaAFScSKeXpUiW2PEr1pWLyS5ftqTYNv7flUPDEzwt2wRcot8ckFvNIkluCU
MKBA/lKRIwF/BPlWFAPHkA9d7OHr9Uf7pA4i2/mqnMA1xxEmkkkcJ5gLfdRd6ob3
er46kQ8N8gbEkexDhBLVyfr44GWtKmIF5fe4LihVSksHgcfyuZHe/hXxzdwoVigQ
pN9cC78arusMjLquxhitf1jJurEsK0JKYRru3nM62DJVQgY5mYKD38YprDEsc9JF
lNi1TnBuli2m9ZG5aVx/fzH9kFv+Z0MpsMmXrmyf5abVWjVmFsXek5hYDkTN29/R
jUGnktoRhIFgBr7kX5Vs0rl3PKaVV/6Xb0oqmJRi5niVaaoDRjBRi1N82ubDrXdj
pXDqJFJ+AuRMhLDedt8d6wxtyNfhwP3JqLaJW+Hx4yTdNzUidJNhk8BKfJ7nxZAe
/ot5Mw/XJEKw1e1YajdddhLicMRPoEJQEq6RYuk/q9C6PDtdjAYcEYwV6hD7U3JY
lbV7zWxBj7H2pg/4y3HGDNUakMgDS5rO0VjS1szdJTqzqWReVrF7WsRNNBeXljfM
qMw6TazV3E8HEJ2Xf9gshszBwP92jwkCprVJn4HdZy5LgGxS2JgqCe6kGD5dDygD
QCGWM3K9AsySNPlIIbN2Gp1iSXLXuUmuCmxvQkt1WD0q7TSw2ZQqPDDcvgudMHMM
40TYI2OQ2QX+l2uLyksyx26RJdlaOi98EzoLm+Izj6txHanxYq/9E8aYCe2Vezgo
DcRlbIVcDSJP4NafT112B8AfsDzbuQF0q6hieQuFZ9DCMvgNAjOOnu3+Q/i0VDH4
PuZiSsx78818vsFGrKidI9n1Re6Ew+ZYmlOpXnEJNHO3kXg7clBSCSp8Jc3gopbl
VC3En9oaWcQugkyKGj1UBskUdlRZhsrn4S7kpuC+6scYbXs87/cuhEOeUnLhSX6F
6cuI4wiiItCQrpJLt+DGGHx1SSKaj7sVPl/kEjxXDOYwjGii3B8vyNBUJvBfrGbw
sa7uFH0OTdFfPSwsdmaWuhlm48L8iA5CqOVgEoTepE2AzRfipHAPgeT2ZPFibUw/
pgk8jAVtL3ui0ftFFpQoH3nW+wJzaVoDGPZs0Def1CsJtQLRKvEYnDVb++21rzkb
l7SoZCp2HGpHLiDoWGj41RKssRfC01bhTxemK7p5/VKghgAjX85T54XKZOl8rjEV
bSqiJuwmNB0XvcICbn1oLll0ErY8yMbzADH7VHtv+a7bH4lcE7KZLpSrNRT9Jrly
LfMncu4CmKPHTFnOBcJ5Lz/+wbuDYQgd5pMqXToLa1cYxda3yxtbpPUlbbz5Wysw
E2jeM8Lg4+bMoFc6TzowLJFeBTwPxQ0gaMpCfK3d9rMC+tobKZheKyUlKpHUui6L
6AIASGeHZkHog5t7Kwpv9cn/VSKyLQpqWgc2UJn0YS1Pn35PIWNolXJywcYeUqo8
SbuzH5lw2XItGRCv2D28DYMl89OAQU4n6Wk3NPm+8iS3Ol/Qf5xthATrx2RNixUU
AkvSYQDyjisxj7X8nVFle0Oq7XE/huPJ1i3GaQN2j9+jQP7RdjAfRWRhwhyEBZZe
XRTPHqg0vBXh5dIjR43jFoY5hNrFuXF/osA1/5LOQhp/9es74wNgCG42/lnd9P0x
tt8FfTo0x2XhGTdEr9HTgwTfNTnReOPG1e2rU48vSSrtW0YV8IycLwmcFIrXoXxW
lXHiM/S2GBVxnNgKtYqKfA7rCufXsQPgulJkMp6GJjoFNsjxa0zDCpactB7GSduv
sM77obVHM+/TgEPQ0Ks/Nb6e5MitB+BSuMezgWw65hPFGZ7nA4sbu6PGgCylFOq4
FXCXXShwXYP1Z6DFKKcL0RBhGyH5U2hxtkYU0K1TCH41BoAYNHoJm4fQlzVevSNc
uxW08VA/b3r7eh06uVCkQYTVHNKq+wkH0rBdpw7hAvQyAyU7nHMIuiwJC3gzf5Q1
FvJBeJT/jLOWyuOhEWJXi73RyjRacI5CbvPGW7nsMyUIpMol7UoyGvo4DkBk+Jd2
Z51T5TX+igzHVMW9DBI0Cs+NmW5LWrPabH9CFuaWTngRP5lO90eofnacMLB5F2+B
b9IO8u5TlukE2W6y699fyqxIgv1WQYcd3WrX1wLk0aGqQwXZ1/hV6DrPQKY1b3N1
Aqg5LJY/NsPl4DX1PiOWP98iSAmg6VXZiZhUgZfrCciN2q0gWP3O8F/0D3mfbk5E
i1+Mhn9WojB08vRa6gPR9W18ZkCYdDA8Wp3ZH9n9JMZocNedU0Kkjk6AvqFl3FMh
25+JFXPsZ3XCJNSiTeMJovcgmXD8nyyZXuVrXAExzRckRgenI2au1QiH0m4mT2RG
ErdTuIRJFS79irE5UPkIebS59AMbCCBg2dQKlMR6C+RkHzDl7RrUa3bzHdDL7Vmo
O9sA/3RZZodmVkftYVNa1cXhZpNCATj7psdx064mTzk9keJmLj6KZrTbviTSlgZm
mUK4gBkma4fGj2JGw1m38vPROh/xpXoRJUBtIbbjOSCRABrGT+M2Yn+NU2/fuUIH
aoOy8Zopd3kmuEuCWE+SKiwM6RM8HPQQHLwD0hvll2QvRQ3/zMjOxhPr9csKwPm0
5Y9kb/iVT/Wgc5+GL/G9M5vYa4NYe4gLNj97TkKo+Tw3rOJw1zawMmgrSOJ93xHE
LbTSvx8hiJVkcG5M2Le756qY8QLAqfe+PpyRX678aRYQraEL1IDeouHiCXC+ItF2
wCLl+8UNhtt14R5UWOCTqzpOzfPCb2pLawBtKjI4Gf12/wNhIuCTXphTuB9GKsuQ
bXecyG9ubWgc8eBF0LekFIO/LMP3to7MkpIoNuZM5e9ZIH1kG7fOuMefo6L/5uC5
en2A+XDczg/rESwjrp+S4ZDyXOT5Qh4Q66JVoyYniNGSkHezciX/d6u1NZ5/mFVI
qd37mPTeR2ismkVgWeJHUJ6BwnZA9eQ0sr1zSJA+jCsGJvoSJGubEDvbznjwTwlT
0Vz5aCQ4tdE8rwIXn9WInss2YGKHdk5c0v3qOw8Z106OX/bIxGyxxlbtc+I55K1b
u8Uq3UKQbFxAmeZWwhORutRy0psw/pqTebTqASemJuYRImJ9XL+rrr2JJzZb1JpW
S7OpkE2a9raFzWqkHw8FNSe0lZlP2gio4y+qJO14AnZMls0VB/I9pP7So+7RtGLb
XxCclmyNxi3SpHGS60yEnUJWp2NRQx+0udVQ3MXosIKeeJRkRYhjSqdLggwD5CDe
Q9deg88rpDQlc4P5KVX/9snA2I3btd9RJEimR64kJHc7v7ZGSgVXHdVtv/Y/Zeeb
YP4gStx+6qqeLcd8fMU390bUgUJDrztr8+AacCJNrj08og+PKW8xzRtJN9jU60s7
Hsh9Zo+HZPxxqhbwb1Od0j0+u59sFfmLizw/+ba004sos0Xzu4B8J7uNkPK/B8fQ
nCwu04tAEZtHaOWEMdpa6CCjELCbbWj9sg4VzydvZToweueDsbMEL8JwmgD91a4+
alXZaAvC6ACmC/SXlPbFkDCep3yPGcUeJW7HgG9Xs2o58buwrpliCPKOd8bwsmc9
IVVe8MmstdgelOSHLSaJgAjIclQBeJ4Hk72OiIONStTlNYvywE/mhIMktLPJp5Wz
p6nbUxmwyC755M3GDvBC5BmT9JYdMfrvuCBaX2HYGTLyZBB/I+4sw9/U34oSdjvQ
oS7L2bthfDkPy38pSr+1yX8SZ3Br+BGoRxJ3leS0CtzXwktkaEeckvj9KxP6lBwZ
jhGqZ8uK7OoEWWWW47QWL97AvL3EWaroU45eMeiQrFbNKvGryttmzN8AqrgDGd+X
Rsxs49Cr2aDpLslVTYXqI10N/+z5B/d5HDeZgPmIlYdL5FsT1f5LsDTTz3wNLR/j
CXRV/+rAZYoK0aMazQRvsROcdiZau43mkX2thsxw6sa9tpSMG67o+TTQN1xyo7L8
+RtxK2LoB5R/jtkdX4cghN/bMqgRmmqTFGbJt+GMlL2vY22+LgcCMSHAYun+xb/X
OndN7bUMtfI80q0SKiC9cBluODgzBhwwz2JlTBe7BG5nJsuwrghAS/xjwgbx4gbU
ydtyBdNlh5t745AYWDCjQOD6aRolBKulazUg53qBRrHvpURNRLQIQ+Xr03dcuxvW
fHlU3uun9uQfjc/mH/IU4GifJmY19CGbgO8M0911hldANnISzJ5sQP+dYUeVVQ9a
XhT9jjNy/L/LCGP+Yvk/bJPMKMLDEg5/6QD55dxDYlTEBlypzCIVyzb6mUmtTg1F
ievxynyO3Wry6fKakgSI6wYlXBAe9UO7uiAaMvCcroa1QyK69+FOb7TmT5Hm1VwQ
wRowe3D77qCknkitDfbyBU7hSllEIJ29WFW+LMvh04enekEIYpi4QTdOgTJ8cN77
lDrE2gTkP2pb4QEoiEDsm3ZNQSmJ6CVDnueS9vtXyQ+TBCzqVVJ1H0zev9ltg+wK
AfCLS9nUehSrec+6I3uTrzdKP8LAeG8Pn0cLMcLUjLsuBaP2luurxav6a1R0dj7c
i1yJpJKC720iQ3CliWRh55YCsDBUUBsml13nvb7qea8s1+9IVNnVnX/uQhYh5VOQ
YxZ1SBcHx0lH6a1NQEZl3/t6hXmKKXLQ2pEG3lLNEkxPpI3JjbiIFm1AymyLBi8N
H1Vnxov7kycHfJE+XKBykFv3ZaqB8YVb9YxqLzotR0IM0QaSxy72q03iaoolhhO9
VpKjdeMRWx3EevJO8y9UZ/v+VELYLUA88dxBoiNOCVlcjoy5AZ/1rVEXe+sR9dIM
3cjy+7BCFS1Ftlh5lPHeokVWXJ+RTeEI7slWgvbo8HB9cQiBH1ZvayNv8kgpxdMI
g1hp/GRoENTmcvGYBVUNuQbHyCZ6QulLDE5heiUcb0Y5kZFZn0ukng3h1DYC9QpA
QOcNcobNswALKg+vWDFAWioUjN8RSOZwqkKR1+Ak6qtU/B185azbwLfkwh1l1vyS
L2QkeSOU4+5cqziRkXdtsVbNHRywPmIV8obI2H0b/dYBFc22fRjlX6JGJ1FsrnNp
nXC81PeszPLQpktCW0Y1KatC1tIGYMl37Nx3g35hCw6QLN1qvbsmtBAaWIDhIqms
6CkqJWFuuDIP4R9sFR6ydPr79UScAX66FUQI+0kixOxXrZXL9dzJ1b7APmuAZ/Ry
A351xMjx3V/1TW4QsxrwxuDYMXpaZu4RHD7+1quHhf0eIEuu/MhsOYJqr+qhJkxn
3X80R15AQ562mJ5d/aojE5Bx5GJdk7WDjB51nwqwpcSGn3K5+NzsbKYIJPEsYZL3
A+FCoEz8NqSnFJaK3M+tVtb2owpFiJOA2xmfH+ySdnOHguV+1sbT2lnOxoCc/fSV
9sBgEBIlg+SHdjbWH37RmCNG3uFKQbG9yCGfjGZmpKdHBuZyTIGxWcapY5F/Hgeo
5SHlHj3nWh7X0CgcZHQhxNom7/KLfjoCwdi3BeLnPO5rybjDLEMPZZTOOvNgL13c
jU5WvD6u4pkzsPkqxv/J2kEo7JF73XPOMU20Php34+SM9dN7qumINveBB65zPI5y
DWmOzrUjhiWkkFBlZJIvZSOBTz94pZFVyYVdhRMG6hwOfK5i3BnO6ShsoKQ4mvd6
VXVrggo58YtieMgUeax6R17qs3Ipksgm8Ilg88bvwXg4nwwBs032FgjI8J5Q95qP
GpTps0XXklSUNdmM2z3b2y9psxZclAWNGuUn+iHbfVRC9a+QeojZZx6IAP2H/PX7
270VXUBCBSGs2P2B8cKjGLDknrFPx94OBnaGlUycKqPrirspFc9doL7Ii1elWok/
vaJBb+TBXIV45EfuGDv9sNefFrNSM4yxaXtoWpDSnF5CwSvOOeedxmDRikimcqBX
8OMkfFE58Vl0yDom5BltkKLuoinCgmZQQ1zlDrU6XSKFQZTXAVf2aWZDgusjdFLT
8y48hWOWk1182Xw06HBuZb4/gC9r0dRfAYRp23jkE5nLYXjeNGDslN0s8oqwXf2X
DZEXCPAEdANVglFFhOh9srsRTAgjs49zok8n8M6ZYeLqszvHUcaLqpeM6Bu6wxk4
vhWgEHkLpwVBfwjgGe94QlwTxfVRjthOeWzMbRsIm8TaoyxQbrFCPXZxyHhvl3Ze
K0QSAjSrlCBYdmc+T/v7yLyf29Mf+yT8l1oKd6EuZjL9sVqdCkx+Tb83X0Gy8Whd
2eyusa6loiwNxDS1Is06T6VhTTO9idTEZq4U7Tv6lJ91A6uu4v6YMyOOMz6WMvZZ
rpAaIP2vKfU0s03E9pHH32D8HeEGCpcwAbirL90VYmCNhDt7UbvBAusoZTssGHjC
r7EXmCR+kWHXWGQfPjOKX/CuhpQ/dc4qMHFIL6f6fUO93Nt041cI7Wgvtu2Z3znZ
BvnEFjnlrpQdcgreMjfFdzfP3dtgVnSWhsqBYDv1xREjL9wFgw2Jietv6ZIbGN/3
MPPFf8zZimIXGB5eojv4egi2whQY32gV7ChgpJdOayaM+BPiyd6nZyRUA7S1nNu1
8mKjaf51ltfwfYl3ovCNE/+lCgroTlEPhkAYG5/FXqWdwLG0dll0XH4HMNy/w2Yw
+jV9hdQGss8y1MpFT2/S+jFbznCp2claiDPKtceIkRSUEQ5cmwoGCxnStMsb3lzs
H6xblL/OzSeocFc6zVZNgl+wMqG9WYKG3CoC7645tpl3Oztl6vTbNLMLBf2NuNQq
XJ+/CG4SPK7TtrUzuEVhHIRauK79Mrl9QC9NQlN780Fi7oWP6tQSHk/ouqLEQAuQ
EJyNDJGpddhstzN3Jq8aDrOUKxvjRWNOr5F4h7swUuwkH9aqoTTfJQUwYPShuDQK
rZxX0uf++QQsY/gAO/lgyNTJZDw9TlDlJwTnpSqHRXC4GHwOZkq4WVgdjPHY7wFv
vYkrVtiGWAgyJpPxUWGqpbxye4X4qBkaIgubHgznJ6yBS1ZpIb+ZtfDghTkKxLn5
G5fk1cHtvcvpVmZBc2rE6wPV85VGIg/af35iIWnFNwaBk6Cpk+0L8O1jJhKRNYoW
FNVgLTGuywqLrKn2NbVyxhPt1pV/YGaR6dWrT6+wIk9fUnMrWw4eb83FRkjG1Gdw
sQYQpZkrIW+ycdvBnLCXL4TKj3rmbXsjC4Igoz38krCYJ9sRVCeBgRLSjtaQJ8kN
qyK5c0/im0R0Rld3DQdokXm3GKquOayPvLgLgr4UK7DxE5MgTZQmpuyMa9Gpsn3I
cpgsfERh6P/ybLRhQvDyQE83Xww2qzQAqUzc+JxruTD7pScHbRtVsFbUaWpHFruN
9UZiEUm5a478E3wIr85iJ2mpgd0IkoizvqdSplTV7DGPkcLyyoLhq9WsRApp7AgN
pGxrkoTf/4Ei3U2w4XXIdEnEVhSI3kBS8wITZ6eZ/fwNVnZbCFt5AQ0vPDdFivP1
1omWuxeqbB+pf4XZEJat9TPa39t/hHLogqnK2dwb9SgyzptR+kZ1kAYovWUK5XgN
dqjgVstYHrIJICiYFuJ8Z31328TIoIsLzEM9bCuZNtrhhndoso7uMZqWkixjwv9V
uLIC2/j1CMsaosc5XOT9QsB/kBTxjk6JO0QtjGm92Kc5WWu3gThTGfjLDcT8H7Tc
HCNpiOz1MQmIosdmqY+GQIWzBhF3/JROcfyUtDQXdPhIBfOZLj6IpoyWlYlPLo9G
PSLlk2gXF2mz39hmbDVptrHGaM88SH4jQLfxNE/6gCU2/ng2swHUecATeVOVBekP
VcM6ZgPEUffVvFHv9PIyrfIzI3d/qBCwo8BNqTu1IhQXJ2QHL9p/jWewaaZ06p0q
Mose3Wo4HToiq+RgQU9aE9enbngBrcqNh/vE659qa87pMAtwvdKRWQlI4KRnIP6n
coO6bCYvN1b6ITy+/lGLxJTZUPte6e8ajegl4yARELG3oZxLZsaHQVriZQ3CRXZI
GIdE10cIQGuzOE/Y4+ma9rpbLztcw3rN+TVg18Fuwzd3+dlHRfLvAFURP/RG+7Uc
r1t8jpk+mvkCncQbcg6e1l6JGu8CcGW2B65bq5wUWITs+Lrqq70Js1UE7oKED0OM
l6nvQlCWCYZ4VYUSpFGMJixqSDBLvNr15wU5lasehe5gZA0/qYZjvimmq/m9GYF6
Pftm1GXRT4r20cCphLKV5crrhMOhWyaSbhnA7PujP8X+A8TA+r9CvX1CQ7nCzzpq
IzRUixieJY8lldgUXpSG9SGwXdkdEhLfdoS8rG4FLnQhwOoiBbx1T+vd49KLknJ4
KOJFiC7nGnDw65spZZ7GU+U+11AZthbTM7d5hAJqUz7MKFYNmngKES4tu2eEzKZT
4dOviq6vGNmYsqKcOQ5b8n9WXl/ht/yLm9BSoSY6Midkl4Ql0twerftV7QnUs5sv
o0pnw/G2inxX5gJfYWu+dgbunZWJSL2B0KgEMxU2gZIayj0IUWGei1iI2kLK17UV
plRX1L0He4uEYQ9ugM2pdNGr06yJJ7pRcE5UKRtwAxkPmOGduxxTlLULF94mdmKO
dvcDBqAhYNaqD6RjaR704eGjd9gmvSq4o2+rR3jmfkgfe6KziRJbM6cffewcVzH7
SZraGb2wJriZUM1/L3gGgYfH33K3HGJfXUU8waOYtjN3jYp3N+/byVzwKWBTDAGA
ej4ozhWlE21TSLfPDXJOjoJuaShEkl9EVrfodFGcpmqbfcDUdRQoKOknpmNEWi3Q
6b7aIgagOtVS6Emp4opjW1Qwqy7i7bvtEYARgZGHV1xxmeZ3slcfduQFioUpuzai
0s8/qh+QYCSJyVlEXBjS1D22tsPzSCDDHvv2OIehRVjS5RvSk5uTIdolzajIUXpt
DHZ9abZB4LBlF332E1oUVCUFB2KcYErqaimRW1y5Qc4AJTHqbQN+RGhoaSrAdMI3
u8O4eKpDARg+97nPT262BPLqnsJJwVxOFSItaaMkol5Xun7d+k7vbT+bOR+lnJZk
cA5LDd9PSOXGgBH1fGiWu44aE5gK+3KCtGKgLotVLYD2AYu7euniu8l8Ek82j/9t
sz8N72uu4IJjA0uODBpMsE2xJtm+77qL5CJ8I5ZFty+ikk3UdeatTJmDfmvgYaaT
yBoA0LyPD+CG0IF7ZUksoc/2AXIdXdxooTCdfqO9W7SH6iDqRu2Ks+v12WZNaXcQ
Y6YS6QrXIvEdZtLiwc/Sst+ZgzJFZpyRF1aZY3Gevd5+wXDh/d2pld76HTxFOa1U
f1daZ3r1J3wcybBR8+ByzDV4Vjom5/1kW4JXIvwJGYr9ZBGDU8CSUWdSsaC2mc2i
X/pJwj6Jfc6ZZJugq2MCwkOLby3PdAGqmZ5d1t1RlWsn4vkM62RXF9hzlrodsR18
8q6ooQmUMbjOLGN+Bbb+xkbpZStpHMw3zH8fZzBSf7jcFAGo0tSvomSa/mfG6czb
mlHk5k6SNv3dw4050IxiQuxQ4PjUVpvkDW0N7gb0eiq8/Piv8SxInWMxvfLPsrhO
Q+IhD3Iq1nhcquvgJmINVRRiE81MxdSQfvFWayIVP3lLR9EgDBr9QtSZ0cpgkl9P
FYQ2OrgMFr0F1zTFyZzsWtZ+LYFQ33INn66fQGtO5LJs/SNb+Um88JQz2RWUvcDT
l1p7E6ysty17slSRdfzBWQd3Q0L9CazqV8I3PPfT3bVmKRmdsB0eyMBHe0B0sDgn
dFRqvmmkPEkXkuKwpVY0NcrxUAqnTSVvTFyFRNo6VAFfmmcVO8qzwyDBC76Wqf/C
zErxUb+6q/ZZ+dP1ccduaaorcE9L2QXArlMOL/Aap9YGCcAAaVCE3cYTO9oO8kNJ
RqZhWe3oTR/PjDn50nP0e5Dm+n6aiYA6nG8ylS/6M3mOlCoWU9d8FNd6G27fsohm
YAIIJWX9wibgSx7pTyQLhfcKOi9AbqOMtcjTcbJyGbGzJZvXLAyIdi1WiNV/Ueh0
NXpx2MS5Qc8KCZlO5CMLVEdWP/EXaD1o+s9NC8pBEL3RYzAlxjwVt9J0Q9aYTcew
ZV022Z06rJdYTv80cBYcrmlYn++i0CqaRp6rUZyJfZZtQbd/MIeYzctae7b+upnF
F8O7czgIyn5jfQXcgVV4wx8XBgh4puVtZp70kuDQFdYHBGjOwasFeQhYy1uFnGFJ
qqsJN9YGhZIlYswovz8ru0EMG8P3yQdpIjnqQP1Ofh+hAQfGvYJ4pCgFNm9eN0T3
4E4xklttvBOdEihIT/ORtLzfXFYyUBYUu13bEUdSoQSsifEHKUXDI8+ahbB/CnYB
G4c/Y1FZBqMPqCW2qmaDEx5h4vrw3hCn5aTDYGdW/zMpyEZaBW+hSNlLACariHUn
+FEG7TeVmTA5o6M1FoQAEub8CWw1ymbLdjNBCic0t+mXiKS3XZWsUNIcWqN3gOzj
qTRXAJ2i/6rHfQzV66fCNkR/8X7A6+1aqxM9RJyoQsMhPe/TuykZUyRikoQpClmz
C/uQu0/MtuRL4pMm5O1gVWEi4qF8qI8xKAG5kQ5Dt7RST0VNTnSO+I0XnTyKV0eG
b+3j/DR38fNhMn+kgL84kqgTCPVVQtNnmgEt6znwrI2HNzFXcCrSphR+Mzl3zATu
lMZII8j5pkq/FAjBCql2Yfcf8fmp7xDeNGmzeNJyvOi+mg1Jb8xV0Z65QHi4+E5w
RFeAhxgNmI26jRqjcZjx31m6hWgbsrvqmA8H5BXItOjSqMF1jfYfR33B1AWM0kN3
g07AkZE74mmlNSrcp9vKfWyfAu1erOqLIbLV3m1MPNF06D9dMiwHpopDtibpswSC
TWK7z4HkcdiV0w0wZ0hekGjAWfzJcpEt8whQRs15/+70bDH6pIR9PFoQ4M6ERxeK
FpQVNcsKH3v+hbdIp5/hoOQ2f7adPblXZZHsU1sX47uqXH8eo8dCCuA5n4hzlMbS
e+q1L9OHOhL5Ix0EzF7CYIJ8H0CIJIkxw7lwmVN7ZREJb+Oh3OopkpgIZUn0H7VH
yxWSckXwjyMx4BFTwuDniG95LxyraTOEb8ErjnDknUrxYcyIKarHMwXm+6vWSCiy
GilD7WifFYj+pFi3Gf0IAmTt4Yk5FtIKUyKz3PGQXBNpK/pU1m32m/IUo5sMarEk
5c5dQwawRv2Tid4UUAWAbjaOqCHaT9i3qaonKKLLjzYndrLM9RI+xUTc58z/p/oh
oG0DdwXJenaqP/O8EbvMPOpDB7N0OqyTjXOXBCePMnRdMIr2+JKJdIppQz86GR9q
U139438DEZS4oQzAW7359NQlhPDee5yDf47M0hvVWQ3VUilIstE9cSGGptGVBcl7
CG9UIEOfFZXGhEdVHmnvoGt+Gn2Nq4XLSZD5aECXl2VCWeXlQi3Ti4eU+SWI1Tjh
Em3bRwozs171BW1JyFOMQ8coKO/kPf8Xs4hkov/9YVL91o6XQLnwrFwjYEpxLBUu
+i8FAATn+wXfmzvdoYghBWq2/zhFSK05scROlp6DPCTUydDBhiXXN0ca1+2Cg2Dd
qr0nQfBKXGpklJFilW6PDLCsv6UfkYC5payVORb9G3XhZRTTnGrFzfB/LFCGCYme
26mr8Dt8Fot+6vrjeoJKq5KQPARhNDpSsLFdeBFJeycsqUedLQ160pV/aJbqasFD
aXroh2yKpjWDE9SUyd19rSS3QhyUYhs+6jTmsogY5Bvl1+NtX3jHl17R045fkelq
cbAAdAuv+Zi7ZLRLRAq6jUYsPrhyAcEJSnINAAMWkbpaQAC4olSb+rxIhrL3D27v
y5D8dUnyMBUrbrAR44NJDYZ5ugq3PA0WXkTI/TOWQkq7Nu1JPyOGZ7v2FLfuTjWs
BJN30fiMy/A9s4F0LBgSOa2DmLxL8Lkt0EKoGjIAzp7nZkMlAL+ZHHnylm8mfxSF
tFsKR0dwD5J/8jKn8/ycteQSO45LMWw1KuTGI8NiwPMOvHTyZStIH07UlDyUVCDa
hFe2jgJQSQpnHRnCiN5pbkOByjoZR8iPV7ZIG91IyMHiOm2Ks4oHNYVOL3NUqysI
asBJJK6wUjDzt7xCWCyEvu3DM3vy5tQMNcqMw1eXU+4eAofoyj9aX+a57wY6Rffb
qVIPpVg+w6JgIb0DZh4KNeLmTc3ujU5/aYXxS4t41L43cNK0r+6oWjCtXvjYLZpp
t9/+VroA54aq+r+TCsjo12F5fLzvEfb0MLQ0Gy97ReFtKDLR9iLLjDp95mbjo5P6
l+XeZaEx0EQbbUjHQMVXx+r/0WWaaXHTBfQ2CIH/EWomVjw6KAfp6YWeDKhqBkRH
4qR4/26IZh5xHRzmoTtwwq3dJNBSlqKS/qcGhZCugZBeXY3G5u0G2vpNbY2De/i4
6ni28qy3wuV6gofx6zrJPhGTlukaqO6CFKbkSFX1HmPGg3WEGQKFdaAAKYgP9zgW
4+UR6BlnoCec/tiO1fofiJlL05ZHA+eoPSDhDlEu4Q4dyTsmtNr2roEgFUYLNiB9
NL3QdRA0QO7fAVY8kvmEFS/0lMrcwGZlRbos8Xq+3KztMubOG9CcI0AeXTOu7jqT
EhsaPG4v2dWniu2rhEw/nQBlbsL0oRl8wA+YUIbA32i1iGIBiEmxAqG7cJOsmSjz
yj2EQM7tLrpDpgDZN5F27kZyc9kKbVnz3A8tisTJr8oM9OT++K1IpX0HwqRRbMfC
gjYzYUdqzo8/5/p0kP+o5qJtPABelzJkPuLiDKakh5sWI8yWy2X0Xqlg6CPJW0Tc
OC5D7/xAx2mex1tnpUizeEYbNJziCD1UCBZjJFUdbbrCAqUICGkm8GwbPzKDLRHl
5ADx3hbxKhjHvW5TjsMiIPipc5qiyZp8AV+qZw3Y1IqyVzG+7uE2Ne6JP3GYDc/O
vKkKTXxORwc3DMr8RGyiFZz3KT+csyva+WuKNCSi5nihX8z2Jh1k3k8+EGjV0IA5
hNBXzkLKt/BB77jkxGzbQ8xhYx6pkJPyyhJFWodDiPC1sCZ1gfXCABc/JHRi0B36
iOnbTmX29LBe4715qBbVQN6DHV8eyii1uJisbgRbPxEm85ZnExCB2Rf94Oi4bGA1
fDuMG+AakMHbRKCPP0ham3VFZO1OwBZJzhVjvYJV+iHGT3LlbIWsKWQmwHS32J7S
6/hdk5Kh89NWmaOWFJeWrW15wf3+mxPEkDXvLrrzEOhfItSCDxfnl2sU/3+8apAx
9+BgCZ0IB8y3T+PYNS0U6RNp9Rbrlk4GL9ErcZ0cGHPWq5mTyy+1U4Gr1OTr7me1
PY6YHi4cK8WDMqX8xl2j1A1EBkvVj1s1H+sBEBeEj7Zsj6TrjVna0BoXojhRUeol
oWalg12tV7LxfYu//9br7KIaIdUrASm09NVc4EMTq1LC7AMUXXQhTnsYo9lA/jga
YNWORfZCDZOdVTwRZ25DC8+sz+zR0QALgd7xGaj5NgVOjL5rFk/3DNU4JVSDP+LC
Pnk2tOfx64ajz+eCpruZNguWK6e7tgOKd6uyyEWx3eYskLrchvbuDATVsrmeCv8t
nDDD0fUXVBYD89dX6ayQxswokn7hKKi25R3tanPlDGJfeyTez0lCPA4SXw4q3Chv
AWX4+VpGvh/0qkkr566MhKVe1wtngRftjAR/QNBiOqXObucqJ8Lim2/uIxvLudGG
CdtBDCRmb/PUd5itfKTtJDkkBH2AStk43aB3IkXmED2cneHAg9pxJ908W/KlqxJK
yguwGVLyCWw3Nl/1XnGdBMCL3yLCM7yrf7iId0aKJkxvtJGFoP88/2c4OP+mnlj/
FCPtnpzPYBpU6PCkuIg/sHZlE5avBmV+HGbiAP/AbbgnlVjWrR++nS7S0TWNp7e1
XfTYLjtr8z3eLHRirS1WFdLFdfI3TAwG4jdxhZJbAF6EQd9puwh0Y2fGWacTgIL9
POHuS3tfPN7WLuH2vKADA/GoVXVWqo07IYaLzSuZGb8BKnX2pZNYghZWNo8o/08v
6wF2I22Homu5bMoTYWJ+aoqxN27d60xSrTivVKwi2c3beW1qcZdk7y/WOW51F03h
N5F//Y5tZGSsSnuVxvxcTsYQFfImRO4MZ8fX9CG4fmeeaeIz3TOi0Oya5+HmkXN0
iNiEDYRLwKOr3FjhGFJJCL0qea1SEOfqoWQWfLw9HlF2UwtWizlxMlTdMbUz65J0
0fdPy8km8sjXUXR3Hm7CYA8fus/z3DEPhOlndb61PTQBDl2u67idJp6TkD789bNk
NmnITOEpj8Sw+8Aoatpolc0pmbAGcG+2MPiAkc5vUjglpIiLawKVOUXiHbLUsZg6
rIrkMuqJcwLr7d3Wkh8F+33BKcETPjKZOTH+2FD19ZdvAwDZgmn1urap/M/sr+8Q
t9l3h74u0GlcV7TfQy1YmlRwH9lB2A/1axbKKJk14S7iRXPC87gnV+GYwLxKrZTa
wdmwLMSobG3fMGV0kO7RSbI9bUxS4YoSVbG4TXMNtYQI+LfdMG7Dmhm6PHrB+3EJ
lXIBDbwPBEPNqBIHJSzUEDszSR33dpdSu3+rA097eg1vvhELdyWcIMpdm/42BV3o
00Ncu4dLgFzwcJ2zNLZMFn2HiP0sbX23UFquHYaZI2wAYjEqOn8c2/z0dv1W/wrY
GxGY8Ii5xZZc6sUEb4aY1kwire32v0eRVdo+AqbqqA2EOPtw3mzsHdZQEf7xEA7T
4qt1QrK/Ey0P5qyc/CjhY3MEGNU0dHt1V+NFwLVeP3gSf92vqxLibq7SP4aEV+O8
fUWO1xIw1OVUrYk5tExsbL8cx5PbjtACugFzN9zJc+NrApEOY+oAO3yjRIHDEcIy
SgVmPMLz0BR2BnmD58mtxqC9RIriUH+zo8sIy65wGtH86XIeggtrFiGhqZC+UTuL
XpBs+gUNN4tuVHpF7TvbrMKAHVjWRUsQvmXVHW7JLBzZ+n9on0C53noL/Wm0CKTi
GTmRM26pEiTqkX7nRASCbYgywMxvsEkf4+627KZJlUTpVcTxHuVBQAMYZ1gkIrJg
MfjH12e0QH8TMS675gyJbJHs4N20I+THe+TL4e4NyOZfztRCdBUyWoJTkcDeUNMU
+p4VSzjWTK8TgGC/9yxZNQKMYdF9qIbpRuGNH+OPA5C0wALq9OZj0oWT4VneTT2H
c3poNvsjeYh2ncMHvDyclLNESd2jjRY8ODzV28Vq8IDqLrSS5SvVsiJNhQl1zth4
RKoPuIjBD7ZHUxr2y0vTRTUzJBcRz3E97KGSoWEhq8T2q+3Gn6DjBhGsMXg4zid8
+WE2fjNU8bCKw6yCziayurRTHNimBPGFfm0EciPmTXKQE0bDYWC/kQQpC3gU8Mnq
NpqgK+Kc0PyU8KZ0i1RRBTVaN16TI70fSozza00oBRgu4/orT/pnXBI9mxH8G+Qh
TE3nqMMx/hfaP92TADxP5hiMafcRNosTU4R6jLxa0g9Hb5NRUMNFu+2CnV67ne5z
GtultZq5DU/lwF0dDW/+UBDIH6TNB7TYpHbwIlwnFdM+XpX0xLXeEQLRlHB53F9a
HWSv4lsdO5Zv4ZscWSC6eIMdNuajbNSDMrHhEi/oxF/SdyTXD3R+nrcwTsBGjymU
amzkiUrTsTegxTjoL1ewAzzDzLXia2cq9LxUID8S5fSi+cQc3yk14vnEnlPT/H31
GOU/IlD96bIpJoLjF60/uAk1H5NUUtBiNi3Mlubu4NfLt6UsZBHHfvQYB8lLr5/I
f1J5qALUJSXIQ+SMva9BscMy5CVwGnPk/eG8MbMs1Q0JG6m+Rblh5agKN/lHUJYS
SY/YHa7LZKL09o3f5c5VEFeSpbf44oILzNI5ZPtan7c92eviy9iJCX7xJeKF3q5A
1mIYriBkyRhUCJ0kRoEhimQlVLISmqV786wtTk/Eha3LcB4drDleN5AleKjtZZ6X
r6DSwyB06YSICVEQcyH5KbXk+Li9Yir0KDJvmd39Kudl7LadijFtAX3QKMeMS4U1
EQ9zlNqA3xWK85AHG3J4x8JUgzFz1Xwpap4Y2L/To4hhk3PaB5PaqdNxXhd2FdrO
5EcL0TNz7hAHBipvdE0WauOYFbtN3nuysa5ie0a/8OVTejpwOSQlBpwino3XmK1i
e3N0BgbpX3TqtuYc27VQGBZO0XNFq0gaN+3x/4Slca8Jaz53nP6tk8I+2YCjF2Ou
9RIC//Z/HpI//W+UgCHiJDC+5yfHH4h/oNAYvYAkMYnaeynzhUPRACLJ35Q1uKr0
AlEPDxKzjOtu9SthpUCtk4nsNamJjSHt4kb1N+5FRrxzv9B35e3xwXmXzJ0xi3Ye
rP9BbJxccot0aA2l/mhW8NM4dyRZ8ZkHUqYjnshTBRsOyt/0jRw5fiQQpDnxShjL
gEBGhc554BMRfyAKKI3xL20AfqaocVomVQVC16B4gWt2bM3M5ZM0qmAwZtEK635E
20zm3ZlvtVozBY5D7rD6k6qrMNajKAX1298gGZY+Ma0wocSaHCvtL+pMbbG/LBQP
SMS3wDb2BSRoOlRqU56DOdzZUjQFfc9ZM64oVJCJZ51OCnEEc8KrsKe5jhvcPcI5
m3Ja6aMrA2Qcr5KdFdXSpFXuY/IKXRHRdpUFx8rJbjFKjl0RfWG1pIUaW3yZWBH6
08oVnwnTyqcykIpmmhOd4Dw2RXqRu4qbvtgpVwZdBAB5k9gxoaAqSNazkerzo974
76bUMQhAUhorCFBsgmSdosr1m9mGxWS3Nk/1wEash+c85VmsIzHHRgr9OQXvZ8CQ
Bdl4ok0OTocONPGa1PX99IKTCNz9nHwaGoHCfKHXYdD4ORSav3EX9cdUYjV6NbG9
ijPy3PpZhFOkNSuo9/feerIvmodF4NDsRAxTI/95jBau5kDalariWInphcZNqxz0
2w1HdrQsKTRUcu8Lm6OMjSFWbTiWuxkvLKO7yfJELNp7icusbxPJMl3poGm7ohKP
bWHsD0iEJjmSsdw31yQPg29uIs8QqTEWnbbOASQJvG/wny/VzGSIp6OlDYYMxmo0
5oT2ErTg96GTWkD/ISf9bL+TVUB6C1SwPsJk7MlEZPPqtBO7ML86/MGR8KS4QbGf
GTBBs0O8/EL6Fs+LKRNDTmLtvtf3zxiQ0Dx9qj91T4Tt2/4BVLodrPAAjfSr9lQ3
5dRFJMqkxFTFkMpKHm+cv+YLkADVEVg7mxyRguqmfJfqIVz5CCAnYWcGvX84xih/
2UQliZHXUHEcVQ0keb0MVGsS5nvEkmQkxdE7W92G5mBXGAZH9VjQNDyK40ekL9rl
O2Q3Inw2FTUPlGqM5RNy31t0UCGt9EDXVMcr1itso8nNllgyAw4NInEbPaVRbBtr
nUjZm4eEbURv00bYm3MzPjpwmOJF32VAjPqcc4/2WNj1ykSstFEsoz5sxqDXlD1E
3XKD44ZtNKTKirs6BbV0TBDUKjV8xFHtqwF9moIl2tJnlRbR4hu00i3ZZuUnjSNu
FhGmTmUA6y9FcyEi9gGP1LpCPQgLKXPDG+T7iDAtL4QkwyxOm4EKlDhYkWr1wRAa
ZLcHQK4B1SpqfYQYaACSs6QO9mXF9QBxDchODwzPVJQ0EN1r7lix1QzJS2z5qoMc
HADcN2okor6ru9dlP6kI9qoU0/uAh3vmqc9FKdtV5gUbCNUpT4HjqOr5RuMmzj/i
EAYn8lqal/cAkXhkjSkTUxWDbJflya72hvLxgUlgDhX418KqTnLz3rOf/l4xuLh2
wCwOWMO+z+RuTSz/6mu/Px+TcbaqJ+06k8EzDgPs8k07baJRwIGGtwSHz4CENzlB
PPUdC5NMnclC1e3UZU6kItPMrV0qIvsKAlf2XIbwJtYxAG9Pd3uGHYXeHHBPCfSg
UzG2b9Z411MKrzCwQtmvYe0TEDmcHRGqKaXwAvXR57tQmCo2Y/P6Bn/Vsh8FXkne
4zimzjTh+JWL1ffR/wout9O81EHVB+woAcLIF4MwXjQpZZ4FTHB+OSGYZh96Bly9
YrWozqJW9SHkUsSZCW6mpD4jn1+Hs90/I3daipQ2QH2Ol/dVfMa2EF1n/R2i6Xo8
84/9l3AHUDo7IKrypVGcPNMo5C+mlxNhi48QfDJS+xAIJkwO1P5ptYDOCHvAc0oH
lkx87Pqc5Khaxli8rF9/08UVPJWEB4C601ePblTuR9Bt5zbzDp+mFYiQsbv9IaNh
B0lKJ/2bf0adguQja2pvVE1t5c+WmqCb+BocLrkowya2A74hOkmpZHeTjBTE7xTg
hGUGRCrXQUAEljsAPzycEINHmSK5Ko6ZxLh60QJ9545/C7kre+wnGANIoS3zXa50
oPZmrBWJpOtVaIpZCjKrS0yGg7q0M+rYygNc9qHjO0+eZ//IKeoIT3SwavahTxAD
OshQDnHrzbPq512EoUDZk3MSbTqxagBrdlIGK3b3/naz8kVeZovLcBbBXTRMk+ba
6M8JZCYuYp7U7dPl/nIVfNAVIVwapLooaGKsm6BufeivJpM82yIOSTarlKQig8z9
crvzTxJnZLdPbkQpvHTmmKEv4nSQbDHoKHwuAsqocTJfgxc8RGsgK18d5WGfG9TD
lkthNdlo+9kDSb3qbgfrYNa2qVaKLYfQvqaF/dpzaiVmlb8g9KRkZpgj8UymDtyo
upWEi+hHHQVGLBCA+9rSY3ccU7KtOTS0LmkxlnsSBXCCdfK4JaJ9w998wHTRqUoh
wxmMpvIOQLV07AZeop8WDZ38I3TEe7pwNRcpTWNZw5NoyMzzV1q1d7HrAvqDNRJC
d3WwD9hGET6ripwbe98/hgUOHLjPup9o4loRHs0Ik4hP3cQ37uJhkMHohKPWtG1v
Vb+AJ3qKy6vcxc+qospqTUGuM/aZPB5WztzDYg9VpHMSWMydBZQvB3wN1g7NLc6v
xPuHqpC7I+bLg8NvT1e3qaU3KC+psoi/aiI93tpL5nxR+xgoNH+0abY/r6ybGq3G
3x8UO45vUP1eB58sp3ZKnI6WcgIZk9ZpgGx/v/5qGurI4nBc2/yFA4QnJcWvp5vX
m6knTJTgubxttU0jh8boh6zDMDWoYp/ARQj2xHik6XKg/AESQm4lqYy1mhjT8AeZ
Ofv3/3yW/X7qCuDrUTk+meumsIAmG+toQe8eFEvSR9UKt7FVzX2HUKiVL/tZyUK9
XrXoTZJEdm/8dsaKbpeo+VQfuu82Oz9Hg+x9CQ9oJFTs1EHhf9sqi/X5k4VNPqzi
xMc1CJCZxErnhJoFU3i1lfvnQtJfIDwaO31FMTKrKXt1Q30JUjMO6rAAah5ZVe5v
ItARG3OswhdqdkbGDej0sntR4tQjA5pS5B5AoQf3tOlBErxxUOHJP3eqOrE1lM0R
MxisD2Xpr1jU2EFSx4U64V90KzB7+g4cZNMxLqq/Po3HAxsRBZS5a2wbJTyvu8yE
EkSf50BaoqvNj2oRGNtQAUI/Wdw+rzMpejDv2r+ZcN14l/RbArx9ajWoxjGjg6q8
m4hYim0ljMbsK6Xt5zLYq7RoARDudjciqo9uL/JE9tguQg7Yopg/EYR/AMxnVnUN
FyykSfCSW1r2u3VbPqm8cyJOhMnNO1bUeItKBwsPcsPlcKs8g0gYZtlM8z0jXV4N
kqbwzxg9QraZLPYJm0UN+1puv7aAz7O4PW2j6hsWgMDqhh4g1GM7Y2uH+802cAl9
VeLnjCCQ3SMavhqUvxCjH4K8sHgnPGesoUsgTj1vigiHGFh8aiQiFx/NwrbvvMv1
iTlbYQ47KRBy+31wmOMXBGvCbwekdduqi7JEIVzWXYqCZ1MaLFYjmsWVm56P5JEX
sH+0S8wOmC6osZqYNLgrPhSO3xjk6OV3WAOqzvQ4rZu6AeWdIiBRcV9dAu6ntAhK
PRWFAvFI9aci8iAobm2/q96HggkTT3uzqtf0iizo0BvsyKzZmcKrEX3e7oxcGbwh
jHE0vy+EcojWrMtruez1XibTijg7lMjScYF0/KS2iODmUNWyv4pgCw0o1tSH/HEQ
Dvgy7r32+k2ocYLIK7G0M0hphKeHca9bXmB0Z86Aafvh4szO1/c7vY1Xq8P5SKrZ
CnQI6YuvahZAdwEI77za0aYFX5+81sr2uhasSZwIr//uqF4rADMaeu/XkUOnWvWt
ywLoM1rQxKb5K26L7ep8uNekC5yX9Csxw2xKUrXDFZk7OZkx0pqKYVETSJYX1IEX
/uVt9x6VgZSHWjau3EGEMMM/9xRp4mk/WutlCC0tNFkDRo6bSFK3Gv8vJzgFoYzx
iovlPBoT402+TcJ/du/1Dw46pmR/GtL8AuGMe4M0QG6k7/4I6YRBf/hOlqEv8EtE
B9T/EQ23vFk0I3ib4ObBtDs/HSLR/fW1RC7q3av5wn3RmFLrg+4n73vnipb/7h1x
L1wBTw/exUHPoj9RZA+hvCBMOtUVa/Kqky3dMep8mdWS9+cLMvmER4EZiuO/G4mT
PgLw7gIjtT6QVACWNU3e9hpAgXjKGkVZ2JhlmzDclYF6dHaujN5tdUAH2TE5pfuB
EM80JTedWFXTYMupg54tYtUArhiRu4GPYfOezgHOot891ga55/RJbtlvqEMHR2Ed
RTchYVsiFWCxz9hSyPX3aznyDiyA7A6DtOTEMwnkQsKokpNx1ILQAPOn8O/7X9b3
ohgWCPnQ5LDLNYdl9rdRrxofBbH1d/UNtDA4BH0TQDdQawE+9hfp11UZGYydb432
Drc4refEqm55eZ1tax44N7WzK+zEsIyMINTBpnpGiKzujTwyRz0ubxqaMrx066Wj
4vBSIOeaUu36LxJ5l7e98p+ujD83Q7ec5t2HBq7GQQPyRL5kEdsQq7W5rdXOSbTD
7IOPahM1pyeqSppOI/pDNUNmwjQKrwr/Op50JY0ZsASTjFlT9E90ZaPU9C+77mCB
WjNCOU+Ym2RDy/vVgDW6xZAQhAQUvRS7fnleSkg0zC2KrFMFGKi7buw8ywP9MxWM
8hxa+CzfREToBEmixCVwBKlLyGOPDTGX1hPbJ6+ROr6ImlqWLORf7+9T2SeV/blp
GLeV3+5Jbcl6HFiGSWU2WcuZWy81k2SWwLBCqwvKV2Gyv1Js2mSKFhCCGzJ9tXvu
jyLM5budw7OnUDI9tnOQW/NmaC+6flMwuoVP6XSW5W9Db7kS1TTPaktgTBb0+3eu
GY9PDy+wwkrkv4dZJI5MQiKy+3VijWsV5SPW2GqqmNouyWDMNlzMeNX3NKTCQzBN
kLUd8t8olhB4CZxFfbmpi1WDDuqLQYlnSL9Uh6TVx2amT9TmQrnpIiQKUIexQeI0
c6f/MijCtff1yBw/pgb7Wb1XQRSEFmdsFRxQ26oux0JnD6rMuvnPCCbMFT2gZ6Ax
ZwFDLvnGMMbyGK0zoEsmkNdcVyUCjPl12hj5oAiVLe02OVvJwPCLA7WQRekbZGvu
ekOVA2nXu3DSFO2xY7ss6KwKdYCKTUW4T3j5It/28zO+Cb6nJrYuhrK7y7kD5fjL
QzwjBV4eefJSQD/ArNQVpti5kHpIGSns9r+uAXiz7Eu1Po7+EOWEpH0miTi40opf
/0JO11ZmwCPHsaPLmLd7tiUqM/uW9QU9L7O8EsHz1QWAZaFF9HkiNFBXZPeP5k5N
SF0akv7vP/qTxrlnlRClZYZWMnf5RS8jFcdVg7AeiuhhCxkumulsXSj0eCbrGjtJ
25CAw+NiUZ9eONW7olDlhIOP4LjKp4Yq9jxS71Zf+8kUjF/Ygdl7adHnoD4iVd4A
iqtfhRcHN8qTkInoAoMYj/9wGW2ympjgP+Hl6oWz3fUPuFas2LtsfLKaftNchfqs
tWTD6T9DGTXS4DzPAfNSezzikDaBIUEPf9LXrd+iESuCzGPiDCw06XkEXysHKeP1
NEtag96u85go1EK0l5Ed/oV5+eo+Uecg7sybeFDkbvnZU13T9IVi5NZMsyrXXhLb
+BPma423cNr2rz51TLesCoFoR5y722bHxpbglcn+Hi3GX6H1qwBVlkapanoJT1bX
Bpmptm/gOEbFokQatD0HcJeOXWyamXut6h/+nmey3MOJRR3NNrdN/IKf1QwWnZfL
Ztakf2YIvVflhldvLxBF/o7Wm4ZRmbEItDkyXsWvlcBGv9axGq6KDh2CwoFKst58
sS7cMfPjkBk3LoMrIH53RN6fEyo9Ea4n4pF5xJUfW6HrX12X+VfVMAjOISVC/Hqg
lnWN+eIC9sp61uWVzneIXmLZY0tZv9ARI7T9E8kO3b+NgCisCXSFPgndVj0ryPRx
6+xc0iL4bicCWJiA8lRAXiuo04h0uH7KdN6nc7YP58xG648MaY0We41MDce3fgmG
9cSqqbenDSJ+5zaEF5OA8NlAg4swyASH9USsnfYvmB4VIZYUHhObXdVPlT7QcH3t
n7oup0w/3aBys0XTCjhBLrsImLuq8AqnAlbuP7z/kEqW19enaNg0hSt7RdK+4gvJ
p5HN9jbdkccD6SOjFF+A+UHBzUw44Bh8U8IZiclFXHoMwM3k8XkqWndubtUzg8h9
0MU5PngU6XAXZwzKsOkGXvCyePmwQi6+lDGSRhHXPJLJQeYoSUVtbjjCYJGZ8ECe
MKgPyQWirxZzf+6SdLDXTSJszHSWzR9F93sw1sJn+pdYaV44CJYoVGsD7IB9/zmi
ZujmqKvB6YFzQZk9ME3Zc1DgNvTEqASNVgHumrMW8x3CT5r5pWkAcmk30wLOfbxW
WNNqNNoGuD/UJLI/J/jzrjoSVGxW24Uoz/HAhLn7u8ntBh1Ac1ZVGk6NTMf90leL
jN1Pq4oTC4MhsNU3WchUb4bQaMo20vq7AHk6LSYNcJxJy9Nd4bAlU+qxP84o6tQ6
X0xHr6PXkqhwaDIB0GOYVFewbsyoe4zMV5R2rJWHI51hRRXi0tAZ/IwS9bJNEVWk
LAsAzL2gDcA/DQFPKrBuV9gY7Om/n2rxbVQLAw+cJ86zHu6F6l/JeVo9UfJOFm9x
JAl63n5hszVxGsdaBMU/KyKm2G+IQfmYhnLQZMRD52lusCjleSlQles3CW2rwPY/
1NBV7L0F77g3KS/QJ370pJdtBcjTlePpkX4X1cWgZLfHfuOuVTENaHoXgsRpe/uu
yJtPruTrLoLPVwS9BwlQbe9uNuBS1VYelksEAKpSIneyls7EQOlwnYKROrplb0IX
2o4aNQSEUjKbEKnF/Rcy+ioLCYCy5UUg4t5PLE1T/Tv6HyyZzCyKNZ84OFo/lVhH
0rxS4fWLrQyts6HPpn2qbCZKt5co4wr/qMKqx8SA1LNLTXB8+dHp2D9N3jSmQS8C
8YDACQCxTkR7eWqh7B4f71BBigZ+6JWhOJPTzNFSBouaTPzlCc2eRPoRkz7dOT7R
LMGCi3xvtbERdisIaP+keTKFigXsS8jZpf96OLWbdGumrY52fBsk3akXTvF9Gs78
RK+66A0jm7zMITdnsiHSOjzXzLyLPsNMGWVqLShMNr2CO6H6LV0vtoWCglOEfHmd
Y/c762VCzct73Gw8g8XWctlSrt48zTvXdJypVie5oDxdgqooabw06qAGsZXcfJFm
Wt9+/PRjRj3tswMQEFd1dKHGOj6ikqY6xDY/IM4XPRMsJARY1kWtHirKitzm0ysG
2tHUA798OBlO9RNWnrjqGcs0OBw+BV9KWovZ6W2vw6Dvi7V/6mqsrdzqiegw9R5c
SknsfCrANoGn4jhVng8qLqtFlPe6VGOAEPJwPkb6Q03IOgHHeLlzchUCRJuGu4Rm
aC8yyMVlNNx+wXvOoNiEi54Cr6cCvgBzTT7IgPAKcXvssQrqEl6Djs83cCtHZ9iX
MBMuKtkDVqe0weLiSGEmFSd8UbwCazBoHzBLlAd7fnCUR0i2o3r4ivoTR4I/n3dK
HXiH/tnI0Xx2NsGeRsCET37mi2k6e6W4HFmuS3DFwVmwjNIQlD531S5EZAaQjCie
z/5qwxWRCjxMFtvZ2KHt7jdsoRogr8/19ptfGEF3+khjSj/lVNJ8T3WZL/W6qMLm
2zBO0AVOj9D+Z56osPJJIEqa4qzD8Omezdno0ahgfe/XpQF5B/8rH6SRK3RxoSf+
5/f6G6bIVwaYGDzykaO5PPO0SFZPtnS3v3Ez413mBNuW76SCa4lPCyV/nvEU5hhC
A5nYOXWAdtVSm1FopKw41/JwzfieZqa03HXENw6N0NA+0E1/JXOvDmPlM6LlXGeT
yOw7LPTnK9gwbRhkLbsYg9EAd5dkhIFWoM+yB7jTYTV1vxxkqDuTBQiuXaHrHgEv
YI7oMooVvcZhDi+uG5tb6vk8Gl2xwWvAI0OqOrgvDq7HeywAy/lZ/P6RENdkRKf/
5m08b5jLK7uVDxUKHk+Mf5BuDJ3k37m3tf+ORxWHPZBJSXGYMj4Y7msoFVoKlvK6
YhAJ7fT4dZ9fU388Kk6mS4vtoH51VfWx5RQWruiSfdVpCjer9dKXM6UBhPRuxCVS
aPy5rULboRTgBKJA80rvbjwiLFaFaRF08c0kLMjmVZBKUo1xnhxpbOWn8LaUd17S
Bjklzy654qoThHaVnfveXLYw6MKEUAtF3kqQDPB2G2Yyb2ZbhxxKb2o8SrU1KQj0
SoGBMmV+4cAJ09yhfLeiJnbqPBuD2UD9CxRKLaYT6xrW1og5BFQivYVlbqcgiv4B
27oZn1dg/Bnuh1AsOpz1HYgWf03aOmInDhHJ9wJuoN+oFvS02JJjlDmaw3pUKdoA
L0KocTcwRkdA1ajAJNcxIvi5/ENQq32eqlB9LAGNVACRobn/BbiJVRA9D6lQLTip
Pz4mj5mzNtvxVyIfJGsdRtjqvRCcmpxgRewstqK+azwa42EsohqXHzg3DivOqt33
dURtb/fA/7+UDtDQCE7w0/G+6KAlNSzjgMrrutJQRqGeXPmnOIrvAyucAoO+TFCp
RyT8CCjWwguoY6mees8qmEDjdJ4+IAlxfc3xuKNr/0b0t3jRHyRo79sOwXg6eraq
HNHtCW8w3IANavlDbfyPeDhGzywmkoUuwLrHj82WYpMHxsk2FTOU9hPSAEl2A4QC
gV0/AqxH9iJ6sp2f53IH4VIQZRZ4bfWfLhhmNTM17d/w0J5eRtYgJqAw2xTggG8I
ZD+rDe4dn+1BDNO+5nzRpeehZQO64p2uGsB59plapLOuptgfsMxuMhTPQptaL8x5
UidSuGO6Mg+toEBaXyLNqIkhsxE/UJRy92pWrovDifippqzNc1VUrqelaq329TTL
9hKxaArNxm5tuamVU0X6FO4vL7UDdzyIs3/R2lzrF6x2NNlZGRkJwKu3TYgpaB1B
qVlT5ca9I/It50dncCeFRldz/P4maLhdjZudzCwYwJf/4WqL8CJ5IJ+vscz/itdV
LMTB7Si4Ks98N5UlsSn8W38BDZYI6sH0zkySr6Yppd35ElJaCankr8tF8eSH9sbA
3EAGsBl+E9fryUhAq7FSdu9ESF+REIwcJW+x5/vWWLWrA3mB3SsQzqbnBhWmBonA
O7XeJLiKJz60XeYC0JadGWkTlX1EyGkJtsEvmeDkXmXc4Hk05vvKfX3dulAuKe11
3zbljkzZITfVmmAtqAF+WAzi88RLTfKb+iMoYWiggzvGh2J7ROQGIQ/k316D35nD
ehrlxAYBnIMjqKRreClZ5ReMdAk125iqZQQIQ4LmoKeQ4SknTy+2O1v5GEDXhSr+
HxktDoG/aMoftZVHpQFyPJNq76XaaZbkBIy3mP1Aian+qg4y7TYcfViw+5gdCTN9
Wkpgfa54/etVK4to8F4lTbLIsTzdwtrVjnN5pM1cT8NVjLqSo5kKONKY15OFLtuR
hT0on4mtabBUXlV2/ElsGdyWcfoAKcFLM0CW30ZLSGP9xKcXtpOrTJ04PNiFJ1yT
GFD6RTlLiT8cp619WvHSx6hc1wcsIrbQ4gq+k8KRtK3I8eV/6grzrCIuwfmpBPJe
e1hRMJRoafvZOkYzAN8U8I+zOTBPRUi3rCWWFzBOddXScup10jywW2JwLOICJDkb
q9bk35TQ6VKWP7k6I2hZb+qOrLSqGvO73EkD1Pc5uhq4PQuH3a6WVFT6TH2k1pLm
Euo2WNg2uXgGQzwlP9wtvCIZtIXu6S76DKO1XQdoupgitkAph4O+x068VQoc5Fug
7u3TNJpRUuFM2dxpDhTtO9lX7XxmrPDBKo45L+5xxINoM0xW6C4V4Xk/vjrDlRKA
pEhGA0NuSgHdJV+bI4CsKPyB5cs0AJWs6bV2R2U/MWobyI+SV9pIF2XVR6Jkgw2D
dW/8uTQh9ya4SxP9OZA0m/ywLNoCELmPN9VzPb6TAP6CSIBl80WO82lgWCmAff2W
Xt6DKINECRUtXDVPsfQlCazqmwnrXRHlyQKSpP3/b2v+WRLL7hM/sbvROmgaG7yp
0FLyKXn/cLWy5tBV7+EcEec2AAZ3QHl5XVPI48jpb7mf28MziT8MJPq+xdTfM/oM
oat88Py6u1QTfqDDhIppXo3xktNU20Z/YPT/5244OwAgu0Jb/AxAg9pssjqTEezL
hf/S885QnmftBzRdEHe94Ut2OShzkl/np39oOsSpkO7rwb4cyYX0MiWfcVdVe1UM
g8M6+y5VJra2j+zwkAT8hfn6nZqMjnXlkOUAIM10qgjVFUVGaUvkPhpfpp+CcS4f
ArPUDyi1uahrqzIDqN5abzq/oyTyg+xdAkdKrR8fvGGLuOZjPkD/yigOs2HWvH4q
seNt6L+In0jqVlmuVkhIJ4vw8jc5dO3C2HbQ1wr4/vgw/EKUsjvFcTh04BaNTryk
66h8KABHiFANuaBaU7x+0lBG/ImnteoKw9xDJkAbvD4IS7yrJKIHiV6OO/S9TJjo
UNp7jToyBrpToOvfuEi21YM9Tj6u9DCnZK31LsK68qDU/3bR1cVvwTovPxXUtvfD
fdG5ChCtnzPupzpA9CFcbjnoB4+h70y9lthrJZPeUgJs3rMc6bb1j3hlGjaJfLLm
E2aYubOdiWpojunH8xzmqKBEjh7chyCwXn8FyEae80zHDxn7Oh7cvpBV31q8PCga
zCv2ovavNd7cQ6Shs//dAyimbRe0+oO/dyWIihs10clCzjLWmSoTSsaIKGkeu7I7
kzIVuSCOwUfmPfh/99RdzBdtYhY9ZX7OTjpsU2DWQKwE5qMVc9LUqyoqB2Yyg6xv
mN2KLWChfUwTWxoBEFQsM9mIyx1E5/SCZG1zWFHQ+gOeNoMtQGxWo1GOLHQt4FII
CvBjftyng7ukkGAv5bQacl6GiaGALDkurWrGr6maPFgzn+fWScG9tipUl3H8lDuC
1PxlCOHi3JnUIUa1CSywBgH2/1tA0TsqdNWIGgFv3zb0j3IQtXZ1M0L3+OVqCUQ5
DZUkPjRtqMVOkz5iif12yXE7OjhSopfvzOYv2Kj5ncDtfsB5jxkbJMmQjoguY7Ad
VsNjNVBCePl6afwDMI9n5i0qwPmiTKjoT1MOhbKgclnW48oWyQlZ1ft3sKzX2bjd
9wemnlytRJFCd4MT8+Fyku+PJ/EqmXfkLHuY34lVRdm8Ug5dsxTxNrUpxXfoAAaM
zvFe9uJ/HT26HmWe2tyYYN0xjHqTb4c6tro6i6c8I4FpJ7MnbHP2EUpNE/dju6qt
rX1sJtS8xL82temYX1loUCSS+ypfa9SMZO1bq819GFvwWp6IKlg2JD7OG8lmw3Gb
NvJLxgpdTxq5J9mbLIivV3htdN1roRoJft87WqnjpC+RhlCRnFGUOqKT0QS5ptyQ
fWP/hwJ1l1ZagkJ9AliuA+r7guaTuY5/udEBexwnVI4HsdLpM0jEFmoc1QZ41GpM
+aLhfplVkWXCa3qftWVAfLwyinE8de87izYbEsVJN8DUl4HgCgufdPukbPobTGdQ
C1oc3qe34uhCO2uAkDLbhu52BBv9nPZ3aCsDrILK368Xe+tcU67FUyRFvNMUdcDD
JXDMX4Zv0RJyn1PR4YmZLZCsfYVWc9mf3EZ234i7TxlM1YmsjCt8sHAjbx39VAYA
YPL5dnnSmm05fhDGLjm2YF6Yi73j+C2e0JIZQL7Et5IITmU4xQb3ReRJgjlGoRVu
hazmHHSrczKC4HEVYiXT2ZRb9WYiW3hpfVcylpyMub/j3mrE1c0uinYA5fHkwOEM
Q+bzsQjIqjiXib3btiyp0SjRD1ihiD86cbKBjdn/k6grYX5t7O4yStnfejK1eR4n
Thjqu/xDnRx/I27l6gjbMiQ4cXCAX26DniCAextr51GukZKcER9T3WkpWnHVOt1f
3o2EIqNhYM1ydwxCErmynG9toR5rce2sJ4RUjo5h6w4OqS9XBaDKzCle55/xAFRQ
JWxH88iVAfKuLaQ3dd1a5K3BYw9V1Rn093xfM1YopdrTbWLdLoSHY5733k1j89x4
i/7Q/KM94u/9x6SfPJ2FF1c5Z7nTSuMyINmEQJ+CVV2HfR3JXTYFBNGNFw3eHAVH
FC/nLnKDufyAUKE63jRvS5L0WhMszYey2qv9/eaXfTrD+LKJKdXm8o+/794+M7Vo
Set6u4FIliDpG8rEexQruG3/NHBZjMO4RMsEgtoocl+5lm4CCGUMTh3UFmUIxKK9
yhklLsU/2pBTnd2iaexgcGagPYDYuxqnqxoGsEETTVOOPvN9kJiAswpYIySdm8C0
6Dy9MMVWA+7pBpGMgYZv3IXzIt88ngt0SONtNeU3xhVcy9C0Vh1tJFQZQHytIxRV
Yb6NzytzvoNkQSBhTf6NAA0RzQOHhrgtVxACud22Wz2msSgOX/eXv92cHx/yToKb
aKrK4hgG5nemb+YgZfBVuKc7rl6diOO3ThJpgVXTvf5HfUC1M5WXFlAXI478OuYj
tWG8PoEttdX33cuUh2lBqkRPLFP7cUIb/y/sE9qR1SHXMyK2jAyQrPOH+fAGoHqX
2biRpcxvQlEJR/o5RlmCRi8/Bwc3hKTfidFt3ASot6mI+rQedy4/I6UdKfHWRgjD
AglpEAuA8Jv2M9VBc9bdWizXvtYwPaqUqdntRy2z8xRPa5MdWnGEsBGD2LLSvRnu
lXUk8itPdKRB7MwWEYrjuiJRoYgwjeWvb4oWnigDeb+Wm370FguH5SLrquKlgCx4
RAuxlQLj3aWiZlf8Q/ACiiWI1kIo4vc6eVv3agIzny8xzBwMUYWrQX0eqA3+qSqW
rowEO1tzR79RQrior2i7mUOCidygJOj5DxwvHxzM4VkgVGs4eXeLDnEfJxMvLLf9
wRxTQzO4Xe4S18di8ZSIgltIyCHBwuB94UKyeLDs2DkNjEtj0YtEehcplcP6c6W9
csP9cfcuO0Lsl8F/y+yPvy+sndU5zWd87v27QOghofpxLNfjxF7HAX1UoQphK5Y8
4rTjG+AdJcUIHGeby7PW66PGtv4Vx8j0K4TCFSdInrS1G8XUMuYxR9YhfbBVCOeU
q2A3dyTeZtXRauq4UA0nbXAcKQLbdMxyx0pgXLBHxIYmSKouACFmsaggWc45G+Mp
wSrhnIm3zDNMnZAskcYpjVhSASLdjBHYbHb1eg6D0X1hrnRYBNTBx45RcYAOhxS8
+YyA/fy6eUQHbR2E00CY12YhYvmwZ2Sd3rZOUa2eivp4iJi5cVsCtOMxHV3SJeUY
7Rl5OzZ9eVQsL+bea99e6NXYG19T9kdhYQKpbq5vvH3YHtXH4uEMdFvuXSuILRfC
kOMbdac2aXQK1ysgAZ0KOwInNtd1IolJpczTkLzLCuhz1TIA85q5ZEmBuQZ4hivO
AAcnoGInb9j84hgbZJ4r7LwuHiX19UjBBgRzKJ8RmVpDdF/pU9m+PTWdwL/X6IAR
6Tnp9sD7pe4b+tNKOzH7nTj9JrzElB+2lcBvNrR3TJtztAEdUlYEgoHikXLqEvo9
kt3D7O617NVU1qZPZubYGYDok3XKTEGklK3+AJykZuSB9vVs8nTJkthu8vc2keV1
EotMUWg/UUluWOQrlXNhFuoNi6HYbiFEfmGhHcMXbv6z61BxHwzt3WXv8vWm4s6x
kygzEh9Pm6JNzxAZmlFk2P8F0UO3DVjzqkVgyAuA8rTjvm5odzYEplRKNWa2Lv3D
0EAUK4vTsXaAO/IwUeXoLA4bz5dKj1wvoJxCdKYC2p6YOav9Zut07jYbc7ilGYOE
M6PqK+7x0REMC5jGcp+gN1dgj4pALtAL4piC1DATQS2e9iE1rxRfzw3Ejj5JtRdj
IvnirjP5DNVhjH3GLi9P6s/LuUyLiY+GOST5Noml+jYj3xCRUwaTSRYjfoWUvvMR
BOQi748L4vRlJt3uK7xvEoy3xzFdJZH8i5hV2wyxtX7asnsDWYRrZ7W1Vg0fAqDU
0lv9KXVQkrOBLjlS+Kvjw+/jOW+0GxXaakRWRK6oEQsP56P6MvRx0Ws4QjkZADs4
psh7plUUQV9FEkYoDFYG0yekWmHyG7wAfQUhQW9pXQuSCww2AyAkAyBjmzguS65D
b0y7qlH6kYJIxf2vkUjsHPkJZDWhlh2Vn9OOz0qTkhrpLsJM1EGrIW9ZpXYapAcC
2VVTrJQh7OFuY4jZcfErggudb7JaPaNwxoE7Bp+hPdUu0yUdgpj0fYn08hSejd4A
KCe4LuP/sF0ai/nydMm1emBkndXasUOw70NPSxQ2LlzMPBYvI43VNsR/OU/5gaK+
dvUQSuroa6YgNez3BJBIno3/nVZz6kNTxDC7weckk8f6bRGq43DRftkkrRt014J/
cGWuZg7JGpq6a8bziGeP3mAWAAKUKO+E0NXitgO+xnpwVUXFl7m8KvMq0xzXCwjJ
dAUF3WZMEJLGUxBAm8turNj18kuuWq1UE4ZrhEwZuVWgACg/xPUpqoPlWBzhMbc4
aAsOAsz+oIqpTHB3jt5cFPVuecEZkATNzChAIJDnum4jw2WnZs1MiiUCJiPQOYEm
AL39MWCGm4lj/BV8fWnqz14VGCDBkrq1HdCWZNNVnQWXyjlRWXhbu/HMmUjq4crh
yyhUeiy3yuVI54vCk+lcc24z74IgSOcnUCOGiqaGU/rmjNnuVXskhHeR7TZvzuzq
9cdrid7A8XX58Z/1uiRTHOSorTwe/mu0peZQCLXKJk+vXMLsCzWtj4KmitMbLiQN
/a3hOWcDCCyQvUAvRtOW1PXXhkQ13tyGj8HUmIakW+8R6afKXtGW+B1xw+EZV3f6
mO8hqONlzTcwvVkLRPnKSpStHvy1VtLmpLqhwD7oEeVdGzrHmmiy5ycZSj4MiwrT
M2StO4GuKExhFWsOrcXfOEkQtXYjIxuVk0DE9DHjksb3DoD7mPiW+m1nroG4yIBj
g7qw1UIe5vxncbDnT1cN7i9woNu+hfvbCxe+xFNx3oKnT6Iqa6utSf3Nfl9taHg7
vuIKvkwh2Dwh2toAfM5KGf/SdVD328wI86FIzrpPO6i76cJXNu3kInpmfB3RId0f
K7wR3D3F7LYhLFtUrE4TCXSnaLcLnru263yMNb/AA/VJVRYwvGyC3BZpxmpkFA1z
NO3Kt9XI0v0dS991BG77ShUPmX8cCfQxDoHDBNFJol3DO1tA/8ZPdYsrcMZdjzA4
IBNdjzEr/BwQ3VGjlg4Sx7QVNEIJ3H3eSrNsebQ+Lmk9P2C3RY3knr6Jpadcz0Wr
j007etDjEkq+8vcdkTTkieI1t+qCpY9ABpgEjO3t7q2sc5GzCbMm3z4jsPwA60Lq
tJv65ZG7udnEd9UDo14gQY8qw0BAzkGMELRjkoylmiuRf5T3Q5metAy1v8kEfN/n
ie8fMYJQ45vpXxou0JaA6KJlFT105ZL8j3zBC15XIqll4lA4G0dQ0oZ+QahNRlop
Kb8naRZDQWbArsIqzk2YUgwCsnGxiCpa1MYYfEgbwjMMz32rSXuKq2VgLYW4HXEG
XuyCBHl3MUlrvBNmwdoigs/e71mrYf/1B9kI+LtSjsR89VpBGYVsQi2fkYJB/l0g
4Hi3Qlv4N9ULgY3MJGWQrUwZfMbE/TGOT6Lh9xtS+REfjfEUHBUEFidQr6RRFTWz
Ew58mLfP8FP328FodpEvzysm7DCtRXuhSKodwJQeHfXShEO4O1mXO+cj1pqX3hCI
CSGj83Fbq4t7vcsKtDdjdpMZ2F3GoqFGdRMV0kBQVgvlfLHh5VpV7U0t7AvpS6a6
oZF8vIg2sz1ngZ4oevijsvSQ3tzSkdG57PoFXphiaJn5bxhhJvn9B1oWc88RJ07X
gVdoLG0wlUi0h+xHwsW6pNctuN6pxAAFN6gpg3vdZB/YHcMvRClDzpwunGtnyDlH
82Ifw3XMaYHJusRch07OZzycS0gufQH3SmBd1aPj75jEnHRIAT8VukVM4Sx8W9aT
QZpREhz/X80DS3KSBmYYcQdaIPyh3IxiMS5ak5zMgM1Hnm2mCROXaCaufWUtWUXe
EkgH3iKmYzJajm9jlbAsRe/aCQ1NS2s9+K019P5uP/1YDmPAjhPAwP+pBgoBvhIy
jtd5iv2jq7eIqZ07qxwAQa+XCuRcLcHEjzu7sDeFyXDEcPwBeC+NvpyMIBjIO5BB
vxQS/ujJOCsQwaZ9BgvfyoiSToYPuSohGtUHRV64lFx8iBGzyvWmF6YLsfTPlCp/
nSstRFvm5sUIFPqXyormqzkexT+dytVuJl7WWVmgeelIkdjb5AlTisxIs3Ls6iY+
bEvS1H0qTlP/MoVYFpT25nzYiCFmzkWbBK4hKP9RFMSQCyPI6pLQNsrB1ICl/gjQ
m38d9zphd5LfufmgOsVQTqF05nDBpnjHA2KwK3w6xhcMYUH2GX5bshxUVIuVwEgy
FGEA7iwNFDvO2JGKG6761ubSjy/2MHwa88bdCsFQbk/aYB+Hed/xhrA6ene4FCur
daHQTHUifrCgv+7HdcQx7/NCDfPzGw6nA+6+TWhgYDbZr3FEDFdjqXUsn7MOHACe
zpijakynATtYuJKzxF1Euz0G/34UYmOyeoihaiUjN4LwSfQPs0f5ssmLJ4JW2RDh
0HWrakQiQTiue5H8PvysXUT2nI5iNFIdg9Q0TF5sefwSbv/SNayNBqmXv2W5p9b4
5oz/PtIO/3a1v5x9of1wY7+KPnWsflVG42Qgcgwq0Qxux3aoclZJsnRs5DyNEvcp
/FQ8Np56J19ttzausEAbKr4pvn33CClMCpXDqgeOWx2DodBNAuV/JzgtBdMjv4sG
PopukVWxfjNSL/jwXXNQLbefrZnAdA0ttWMp+XsAJMixyipe0xqr44rUFgz556Sw
S01EvKRz7x0EyUGyaDJGpiAFAkgcAGq5xvjNwN+7YlGw8F0s/Le05xrfnDiuVVpm
HZA+hhNpontBZWzp6T1UJLcnvvSdWZxKX6b8POWY9B5wnpaK1/pN5Lkt23Ye2QmO
0KTx7Sn+hNaWP4WGeAe/VnybOnWelUt/vDUPmCqAQ4yh7rh/3rAEawtLiS8N6lof
ncWBxZBfytpJrzlI23ADNpm6hRduhhltASrsnmAT+h/v+EosU06L4xIUjlbFq//u
wAzUPZ/P25WsxfV6pvOdpDcexv33XbucSBk0V2g80h1CGcpkro2axWIyuHoyfRi+
afQMYgXCUHaVixfAKdiVo3P+GmvtaLgV7Fd5RMrhZ+EHu3X6M8pCklQ8QfUv5oty
bUL8p70FdikYz8aY5eW6vLZIHfRik0IfBe3vViXd+s/RD3HsRhgpfWdfZyCN8X1c
13i96HE1yEq0G1kPRFUV2rl3AUtjmX5X/aJQbRhbmt9wZcSqq1Vrab01EkxX8qSj
10Rz7jCI9EXuKuUzwC8UMKgJAW3eqUC560sKb2kC4TjnqpBjpdZQBDBF/J7GhNrS
hv3s8VUnXKiCB5LFarVrXMekF3dEGmicAohE7ePbgmVjMwIe2WWQPpLDrqNLMNaj
1s9uaSQJ0q9LaJCxZ+4MG+0z26H3g3i+iVHalgoJhSuGWStxeo2VdRnieZ+BSvgW
egpsIfzCizfB+xXvEK9ck7WloCg5Pp3qtsbi4oS4iiG0ivvGviq+lfVOr6EaX17O
ru6YCIlRJA9BKHuo+/y+FGcCVNx+mKbuL6/HVGOi70Jl+O/gmwNqVykuUQX9W6Ux
0GYN65mz+2m13u5s09N/K8T2Tx/uKD+Ghhm/hucEUhDx92pG98f12XZR9u2rV45i
PPuOGjh+Bf7hS1ejrAwV/7xK0N5pl3Qnrp1UOHRw4J/tevfLanejd1B5N0KWrwBj
a2kIj+nWne/a6g/QgW313m8Nhc/gT0cSwZsauygT5FKBCMwmq34SJcHGw17MNJEr
4b2Alcxq19uI6LpkR9rKVtGZ3HDkH3EsNQ53raMMXHzKkdbsjD26yS8FlSNhjC/1
+RMj1A41a3kZBQLPu1WVM3KDILYewMkGIaYkWRF0A1LPRdWuxbrBfAR01FgGBNeS
+2/1DscNI2h006ndP4Y4xP40f4CX/3o6IcfjSV2KaPK3l8jqOadSJviqlVZV5JvQ
3ZDTQslSS6eW7f4m6bE2QVZ/JdrdNu34H5U2Pr8a9xP1fdRIvyhXPi37EocHHH4X
4QxfQiU5/4BTizb8ZrL34erMpzU/SGEMkiqJHMLj5gP4S8MmasL7uYAb7ymL4OKX
KYZnzDk1P8nDOb5nHc1+GRwjV5eaRA52NF9SHi5jVvqMeiPN/v2tj/9D0esvZsjq
8iQtdE2vKi2gd2vreS4jUnGkc0BKCBxNazeBL0ZyrgpkINCH2yHMHeinLV90O4Ng
tmXmfuu6Tj1DAXcRfsHmmB4I4hDmW/o/h9GeI6butTBhiNo+BPRwLtuBGF9b74E7
tKe9Cmdm1LzVF7jD2PoltmFoHpVZ/yEkk+FjcXaQqNcRsSRI1X34SiuOCvmpGquR
eECfu7IsUv0w8SoQ+oEM8l5SmLPtKISsgHJxFYqn6StOJxwig7ey+gndt40W9Yeo
qZ6z2v5smijW5qva88EJjj6ytpj4BgZzbnRWsGnzTA7OhIt4S2AAfdRTW6pMl9Hm
+v9dY34e+xMzlBXCLYXoVreg1kQ6kDt2or45mKPaOmqygf+Tq/2PmWe5v0uz9u0H
Vm5eEgGFHwVHqX45wGTAQHhinYfTmMqSpdMjmVy91i574UAQP0UdVZt90J5EOWFq
EsDi5niaSM3Shs6cfUkVdn98+gQjmbSx0bY+EQMdI2AbZamh5qAS3LZSmGZecGd0
gGwpAGJPsxP6dp4IsPhh9uFvzLQB3cwBD1QwnEBRf8SYXkQfqkyGZ/t++NFH7yeI
xO+lhfKqFc48ZMjn3uwBA4PJgEXr85JiwMAyVRdTtN9Qn4llHlGWGzB3QnF3+eIv
yYdM1uiBtSDlvITr8Rgk9GtgZd2wbkEtrILobujDCOPz7c95E0nOsW3V5D0X46L0
06Vj31GTVIyWe3FrpwPZE/jV6qEYOP8aDCQ6LXEqL8XUPlaBgRwwN9ak/jjXSy/i
BX9WsiZ0+Odu4G5sST3/twZA8SrRfMHqft6UDOGl/WepI5LEy/brAdEPqKU2pGCh
DActiFVc0Soud5283LbHyKtXJfzGTyY8CrSG9DJ65sLf5Yw+XHbjHbFjyxms554h
iJyj9PlEf0TIMB5zzQc0BKTkD9ONaDQwvErIz8ulscMMdipKbcOQux6RyQy//PEh
d+eYqXTGPh2X5FqV/Ev2sHoSF2G9CrAj6s5tsedbbUNDR8d6gGkdVdgkoQ171wpz
o+x8jUxwROfEJS7/p5V/fPyUxPLuReaF4nw+v+nJ99FCF/pDGEvPnRS98S96kPgO
TXftiH2BOHwOYvnxaMfj1aiG2+vVI/VYkSTxjIZdTDoXjf2xsaKA8CzYzbSrcrcd
kIUVKSQtsGeMTxGraeUMox6XaUYeV/HBfQ8e9ep2G6oqIl56XYihpGkXzX1q60VU
OjcC08HIgSUishIxmahCXkPVrSlwPXHGzg2PFIyKjqTUPKiU4CkE6TGFwa4O8DbD
f5wv2bII5x75DmBEyefLzMqUKihFRjzmz3qvPUTaS7L44IGCvJS6BD+Uo6vn/zAU
Goy0Isfvzv2kNXMSu3yC4E7LLca2ccfOzPaktW8nEOlKqJQs9rrctqV9kuNa6R5v
z3k0jAxyH/X1+8Iwp9AMTNcmD0MZRRkaF2XCU8A/pwDaXQmb7nV++kEg7YAv7nqI
axI7OwmTidrhwW4B1IAt2vO0t2620XtCAy81ciphamO7kTepkKw0b4dsrAJRlBTS
ylJHYTobzznrc0iNJPqFPGJs0OfUZ8bC6EP5CV+klMZfZYqEKxCMPuOxgeKeh1A+
OBXQf3lLQ2fDa2w4y546aJZqrHK3UAEab9wsB29IcrrnIEov7c93QNLFbdksv89Z
0n/zTWw9FmdO+f/naa9gkwX4+ptIO1+5KhLaWJMo5pIxA/nNb+2OYSO0rExziCUO
YpH9NE2RolO9QFbxeeVsLvi6V6m2K3s+22+yujwbaYr29G0ShpAr38HyeWCY7aD6
4ZaZ41FBkk6zimf3iMu/8go5ApIdOFvC03o4+oeRtfdP3eJ83Bx6A/YUpEK3qrqU
I02Gu56N5DEpnyPujgYGS3vfsTzkNG4NgMM9+rRSq0OlmDxJZwavZNemC/vxghe4
x5DkkHD4i90HVshcwvoMkfAJ6dxkaW5cPd+rL7iwUoh8pWkLqlkKNHCL5aNS1CWU
djrhL9bR9Fb8b1x0EMzbPQGN9Evnjhc7XgI5+cPbGPkFbT1mpOM/TgP/f5WwCmdl
jEuDDTfz4xF+JKreFret6JyJbHP7pFfUu6aIQC1ZcVng0/59ikGES4Dn1GIyu2Nl
/T08FXo+0xd+JQdr3m5/CXCFoFUkKPRnTOzn6kPnkNUd3zS+LrTh5ghKJAhZEkTr
MywDeY20taznehDVoy4lqONu+JqgqUZSBHNqjJHGPLgZ1UrBGbLBhtHy+mX0x0nT
00M8IQtloIkdWSK9LJkryNzSav1KCvy2BqDC/FsyfsKmpqeMHXL22mu/h3slKtLE
fzFnvAenry6Uk0WK5PmpbS9UBHAAL1h7UTkXvE836h8ZjXQIU9D8BeppsffxPhn9
MEuHMEw0g8YhFe3nVbVfYFMa/ZJCw4kBScL4AUTPFN5xEa/8ugFR84apx2sQXLzr
0KA3KtiUT+Kl8J358lpqO40y6X+NMr4d1V7FZzyCw1/vERVafitNTBh2Ue4/Joc0
bZKtY9Lrcnjc0o1kd7LLzCUdC1ks5R/qTwFOxzldCLhiJ/CwsyOsZjFSsZCPA95g
B30Nw4lNYQmMytmPGA5G7x0kkoT9eaV9SPHdapBc0aurDuWTWZDJRpS/8ujT9sGu
xIdP1XdfpFzLdOKvGx545T+6ExOfxcYmoJvtrW6ZsdxtCLwqR1dwf46d8TrVGJC/
3vbiGiynk7NGmSPSSpqBHLWzZpRUFjScrCH5RS9WdjGIWMfVzaeYkN6IECK2pKZI
A+wTQ84IaYiZZ8KA7GRCebdiHvwoH6zhQ+QBhABAaRJGVhlFxhohcH00l4/sdkZZ
DVsBsF/6w2W0/y/h1ImknrTgEkP61etN2q8DMO+q29s+CKiVER5vOJIj5m6sytQC
cMyE2oBJLM7FOP7HRy7AI08T6l04bBkqHaV1y3VLsYnSLnOkQc5fqfSmVgjP/WsY
9ze+gCF6qd3eV9qKlhZ57Iwji/HrHVrItbyohNsl4nFQOVJqqhuhJ4F342cMZZAO
tlqG9uVNiD0KtUKe6BK+FB90Xg2vG7k9yWf6Si9OHe0DwBN1RWr0w7ppA7feSAl6
Yg22U6sJS/ueMJ7ZZXUkxcVYV0LhxrBGHZmx2CmvVHk952HgoaMWp8zxDiKQSidc
bIoPdLwiCNZOKXhAUuP2LGUel24cdRn7C1Rn8iEwx9IUelSd7AAbkRfcks69JY+k
gCdy7GBQDRGNEogtEBLAn1Uixq0CrSgWLcwWWEzuWAwWw3XJrn6/M9cywL+RDEDd
VFAK39oHAomaB8QBqNFehB4ReMBTka9yc770oBlObZVm3tHJvocAY7nkKGZU7UkT
4IZgAhDBMpxDA6I+8GdnUART/jywPWlKWKmUGIHmbhm07iX7CWWFM6dXqF3VNs7Y
EjIFGkgos3mqCdOnuc41WnAKZ1D+uja0kGR+4lnFrosTEKT2uZog1uA5XXc9+F2y
o9jyicuSehoaJFxZ6MtbatUZdobj30SqHybyd8YAJHrZjESuFTIuOAMfc/N3swvJ
Hvj5YGimpf7174gBkjaPadA9mNUAqsGuSUqcnqQI38ih95/9lTrnwmp/yetCs3OS
Xwc6c98wLz+c4+ZvGUluD7zk+lXUkERomjuRvtmFF1JwdDWOSAxU4TKc96g/kFfk
YLlYN0vnrRRha5Up1b6aDlQrwSQUPGGkXlJENk3CVijKaFUZxuXiHmuaYw3hIY/L
QiCb60bA7/DzhzRNz6mH1jD2UMmJWHabi2sYRiUyG8i8VZddsCjUHbOskGbuXk6J
nnn0hfQ8zvv496xhe5VDdrT1d4hD46drHE1WxNMW5DG+cUjZPPncCXrlTRYn2w/t
TjmWXvBTt5qaCYNfdHg76gwLcLnGhzjfXCrUrY4fsISvn4qoFXYwDUMqUO0X0TfM
mkicJoERlkxnUrOWbzEVKeuRW5qu94kul+Nzpcn8fg7TsONQfqz8tQEdrkAaoaOb
2bhRSpIWkkJjlAoCBpyVB1BE//USt6uTTyihL2iGsmq3bNrhhcs8v38EFUk2HvDs
gGEG/kpkhn8hEJy+vhwj75IuakcgCPhJ9bPFFEL6s1FY9ELaoNoDIM6RVTxIxawv
n2rM5bHtG0B54RB/tPJRr9F4iX35gBsEJGcTXmtWTOJTsyNCbw0TxgAV50ulZt+o
qav5DFkFhCD156NVAnPW57ciplFW/Ox0yZq5sEUK2xT7HRZHuQzDnd8OXFsPqX4p
C4amQqqUfEo5oPWLpsfcWV+lMetdzWpTMmjIFnGa3qZBwMWXTgZIs8hdiHSkvp7I
bTR3ScN1yg+s5443uy2UM/AMQqmfMe+PdrQK0h/TtdvufeklzNARF//ktUgq0j7D
bCD4MJSesbcz5xBUhxRfI5jcuYck8MjEbRyckCfX8tIiSVd2EDfA4bqzPS0Tkaiz
1YlkQjUIE4Kiv2zwyANsdzgFAEjmRZhzUrUu5YkVKphZM5aRjpaKnfUKME8iQptZ
Wdo1rFa1CxGanLapBV2TiGxqoIa08vkUJ5wsFhvPhyu5O6bsm0OP76d4bZaePO7b
sVRKfIT2EWjyW8YLVZmcSt25XBWDC0IIPqA6u5DYi8MYQk1YWaQF4LFXG0iVg6WV
sWOOkCUYe7KRHj1ZMVcdGgGFIrvMiSzbRucrFahB808IteCezmoKh0NS4L7dzb0K
vFtlVoWqqpZ0seV1RPrqk6Ad1uNWYew4p0VFor+g/bq6sQw8EAgjnbksfyPdu1wv
k6vrfyc3GPZxBuuhNrLtQ6Y5Fx/aKSuevefsrpFIbR+sju71OFP5gaTw4xdCFSuv
Hlr87Q9EMvGYRcTuTW4avhUnYNcFc0rIHqPMYERKKM2ovZmnVeU2dWwSOuBnoQ6j
KbTdA+kAQ6RXAbraZpWQSCdUwvolmydA84HH1YOhsgi0/6lPG/TQnYF/13feRD8J
+ioIYgIoAydBK/aS/8f91I0wxPVuRxZotxs00y9adhmV0MKhgMInzjT59E/Vq46r
8TvtOzR+amKdSdCKuELnSr0iiPpyA0Kc1muIKqoLct2tIUtuLbYnwWZsHAvTAQbI
6q8Laxx7nM+FbYwxi3gSWOFCqOjZUg1fTZyHEo8Dau91zWcRRCI/bpLcHSdM5buT
I2cSAkvQCyjWLfmvvpax1/wMimIOaPStXDruvpKAjrLt3Ii3++g1SGDNN/9eBevd
ylkTxI6q3N9bAAMyK/1fU8HNzYUF+C81CCvjptCjWXTD2i+Lx8hRzhG88zJoCG4W
73Y6xl6opZ8ITYL2Fs8XM95RlGncQOCeTvAzAh7oYbUMHPFYhL+fTzQX9Zf50I1B
M8Q6Yal4lP1SsMwz62VA0j4oo3rAu0dXElHrAmpHVmCAWP9kvYeq4FPcubQWautt
hZIVRLzcwTrVqQPyaPSWWcnOfgHZMP9VMSNyKwrhVwPThUd72MqglaguewNDJch0
SznZXri9SObC0eUrP7o+iWJGy660R1oF1UkYVz4SI3W/SgHymQ5/Tq5aQLTKHDXZ
HeftfMN51MhC9iNEvvnExKSl9VQR87hAPAFNHQ/TP6O6LkZLz0i4t5CohJXM3yVE
cg5PaJJRosfnnfiZc6tSogRqggIH+H3qM3M9+/osTpRwF01bgUtY8n5D856oTbQ1
WYYqz+Iox0Fe+mundCWkX9tylPySvU9fBSyM84tRQECiAZ8JX9SpxR+i/+rRFZD2
vab1nlCpD8QOIVZ7cVCwSLGoLuwENOQL93kF2RlkJGemf630PZI0t88CwFRxzLgs
0rzKvHEkfv+GFJSRmlzt5rG7wxg4UIpeSaPu3AdwnHeJfuVSxtVX+VWeq2yciLEa
qZDUBUGBUZdbTPyx4BhiUeLCk2TErSyej+VkTPNIMinRcvizEkW3kOblJA0xWClh
pQ44qYa+lFUtreUoAXheyS82kIxxwpgEkCuZRIZBaQkT5Jjjl+mGXuc28Vyf4v4G
xIqIOTGRThlso2G1X3JFqfVkgNJxJNlaEHiY1Vjy1GeXU1oBrANMGkuow4hKx2NQ
RD8ZpHgwzLuU3jJjjq/6lI+wZUFPjoUpHyymLQfMwkX81seTHF4RcOc2m0/q5CFG
wOKiWFa//sDxTMKEZtILICDQfpxzSb2irxK/UGnzWLaHAdtEAEKfWmZffIc2Hv5q
w1V7m9t+7PQRUG8MbxKaWUl+PPDzKbXsB2Q8MPuf4EKoal5XkDgRqQ5lQmkr3ZSi
6tae05OzVbZaPLuHETyM38SrSme5am5MWQfKd2OePlJPapffaxMHv4JUDLslofNy
EwRnAbU3HAV+Qd92BCnoXCuW36We/4fo0iqbfJbWurtGdfHU6BUT6D1zy6Nj/svD
oOkwaiwsxHK7MPVHqmANmmfqqwP4ffqzsmoOCAOsR4j4k9hwe2plsJsNT1UAQsNZ
Biyxa+Vk+bSBIXk+qi0B1OiLHPwbrBmMsvwguHrwfJVhD69T74tvK/6JpPNOg/eh
oY62Jr7ZhrOhHRFZ6uk7hjZvYTuOrzJxHwrNH4P0jiuYLkWBMdhLLeRcVkXX0g1O
IYMd6TkTQ13n5v2gATwV1zZDukRbpsjPQZcoIyVb4tTY04GgNqPExxpRysDXNXjJ
Ov8OPUnLZoRZpM4vFOnU/RdrGyXrudM1LJuNcgF4sy1kx+cZZvQxC5SRLopAQh7y
hP3wsAWOmQtB0jmIoR6pqv/Wxq4ZjD3oLYbhb1/GRsKWTNX3+mN664vfoKtOG/r7
kh8TCSuPlWYqU1PIJkzna2mW8HwtrtYPsvuotyG9pr/Og6qieUsel9VgFRf6zqbr
5nmev9899XzjXWlHmZ0DczwNhg7IupLlkTbsEN9Gp+ftIsQnvNf6tF9MpS2jzHOw
pt3YDoTk2s3NKC6DuZQYoJSfo8c0Cv9pcuFJRCbDJgsHkj3QTBBhMSb4BxPKNAaZ
RFZ4GeeUKPRNVP6GEwaK5yee6hin2Ua6jmpQAidjjcQPVijaCxnGiyQrMVmHt2Af
yOJGmORxWmGzlWkUqqiZy6JA0CgmmKmurqVNctOf4brx6Vztfw2TU7IOpmaASwka
s1JsCXZgjE/FHVFTNYU344kRKITrA09/+lO5TRYLJw27BUo3nXr7OiHcFhftjT+J
hMw+ENTvRC70BKlAjJuRd/UYMtuffHm2zJY35rap8k0Fafyn5jV997dhkqbzuLcp
i7p71qZoDIGc5+Zd2PlacGLtjbMC0d4SzqkBzkFF15dEGf6srZPJ73Ijr4MQDyUZ
3vJuxM8J0sO2oNMU+MWYEEZvD3NggKZlAOg1/n86pDOrp7L8apNFgxx5ijaqAcAY
REX9X5bv0Hx5ZkgmM7ue1lio9wdNtRXbcqJlqnU0Na6442Y5rrZd6ZHKJUMJ7Dzx
gcBzkxLObyQnSY1/r+ifaGajBR+vyyX+N5xU86xA/LinlcQAls63FzlgYojpH526
4TNxmoxgCjZQdsAnm6toWIFoqQl3ElFLcEScyijRmi3SkgYeNdlNXxTWJIGeh/in
IENUH6ll0g5mbpVrIjWYr6HCn82sBPxlV729lnOUUwTYyD5NgYP+3+UsWO7kgcYs
3u39PxrBi1zCF98puh00WGsvmLYV9oFkDgSz8CXlAAKvSKCFmMi3DScN2CN7JLqU
jBzepSJ83bnbhcPdbfVQR/r/f1SQOQemCNopWqqNfVnLCZSltzOnhT3nC2O9ERUL
YDDS8KWMJxK4qWlp4w9n6XU2j7QB5Q9oyk8ZKOooEE4fJc4Fl/nAi3rFwUt0W71h
csQmi/i96o4Go1dtGVRog5zIkLFT1ylwNqYJsCqJu8nMYPeezvnxADFony7clgkL
cdAJ1YFg/zND1pUaA1MFsTvMTfEEhFAhNSTeE4xwGv3YZRP7AUXUIqua++r1S/rg
jFbJUm00Mx6jOYVKVmw1Xh7N9llyxZUw1wjw27l8H513srF7PLWkHuiX9ol2VOB2
zP4KIB57SBkj6KjdiH/eF/J+ofw2hRuPzbdzDulYc2Im7LEn5yISiSNXDKjRQlkW
a+zcdv5Gn4nMaVbavzl+ssQHsElLm4+uHIvSQycpEPczEorHi8Lez40KlYotDEKM
aF7TTeJXQIb2oFjoqkQ4fcyvEd+wanJuM7E725G2eVMFHaOezVFV7/uwXD/CPvGO
a3zZDvhXhry8l0JocVjXs8emi6QSRuNHg/ReM1pyIOs7fk9to1RqHiNrnSL8rmHM
GmP08MOWgl/MpTCN9IN8ghh1KfHKfLoj2pFORiDkPM3wa3UBsr+ToS+/znMq2EmH
abDlkt9bU6M15JGxksRvNINPaN1uzz6vRGb8NdEMuIzhljm5APaHXxEw02ZYBHaC
csuuwNiM+iAyMpan7BaQqB1nFOCjNQF6lFBJqRUP9xxdYtOBG57obEN+UTNa9pJZ
mVwCmVN8lsPdw1shMVmc0m80/W3aC2/siSR+iB8wxP7eDLpbwrj43N+00sc1fm3H
v5RjmNPmUmjp+HtI2G2yIqeU6v51ylkAznVV/jaKqg3OXesgmQ9zIPC7JlzUR7lb
cIMONPROw6XyH2/L2U/Nf+kVm10zOaOfllJpxuoYhZD55OA4JIFn8ecGY1e10mdu
veR9DqMU9kGMEY4IHlDomazbBv6AhtQcTnR6TFuCr54M+TLUKKOBTELhKuFw86kF
m9JvZT2RICYchVfaWlI/MnE5QYI2JQYPXNP0uGA6hqpzeDtREwHHd1l+ztDxs23a
UHZx0DmAwBDSzAMegtAp836K1tjVZfrsxcusW6Nxoh42/XVY8msje40rmHKuGsU2
N9cpUWinNa1m5M22kUte0ZWDagiGeskLxCHvXf0s05EBUySM2HlAr+FgYauArBTM
TusEmHdXvYb4KbIAy5mOBb/LVplSeJ6mrvRqom0wqFtlXiZeDzk8K1LxCu+dAhUh
NpdVZJfHvYiAdqi2l91PuM1wQTpt8H7ECXkGTIWOOv2sVJflkrxOHb30VjWEcZn+
qc9bIK3Y36xKTAblRja1f5sMCGk0Nx+pGej6fn6nF+PywCDPDpUuVce+AEW43pN4
3pURuf/s6QoJBCWmKDcWec0lIjL2F83JTJPQMeAUPGD9PDAygCTZGek27SLqhpMa
DNnjFIfupoTTUOXj558fZCUV76M2Th+ovT8xsDgUCk35wGPuMU9hi+4zX13y/8ct
5J+e0lUW97Mctq3kOt1bBVmo4cXRa6oBu/U+fbrkuwtyeO/9jXMEPLI5Dw+UVpEj
KtvJuXeJt/Dzz6WAnlg6+P9bqoLyrutDbcGtxU/L3GgCUaE3f1qQZManwqogSx/v
ukpjAfvrSLOnMiouuagPGDB0qTkW6VqM7sRjkyVtp42szc+oKGwPibvNDGfAyUai
4dDka88eM5SysasiUjPGTxAIQOxbbhHiwezA+PjaAI7CScyNtI30QqFP6NnOuRFw
jUBliirwvcO/TRPdlp/Bptqoux9vVr27yGMWi25RA9yc7ZbsFa/Mxf9tpImbNsr2
NPtzgFugWa7TTk83/zqN8bZAvao3B4v0gRFTCdMz+bl4tkF4or3sCvJqObeWzMBQ
s2vwXOIX6T8x6GIY58Hx/XBEvJGjD3W325B41wbhSffWf5XJrWbdQ0kHfZrzY2KX
7hqDPLhSmplJI9njtwFvuIm7IagsYcsQki99jgTvqqDA9cI/WsnXVtTEeqdqVuli
eXQvAAqaw8Kkak0YCZx4B4RrJsUaWbgHREvCa2yrySySP6tKsvmC97d2kfJSVn2J
PLN+EmdE6o4q6GVHZo40W862cbVj9VUJBxNC3wLDPTlQx5UNn/pNUjUX6NhS9/id
Ir3xFsBcLW0gsPdnQi3r6hsZn+b+1GIFKzO70AaT+lDNOIbaNTbLl3l++xbygJn3
jKTrdIW7k0VS3IIFHTFUI2WW01EKNkeOch9w58oeUOyaQWEdUJo8uyT5ZGE8qhmG
l9pxINExcTCDzvafmY1NE+MFBA9dmXelNPJqoShZUX2Q+Ek4TUEBhFoKy11qXKr4
yDR2SMb+ResZ9SlXD73Ifr0f4MuMcTwstBQCVBFYfNrbwT8HCLXgX17Nqa1bDJht
HLLZu5h8OpB3WrCfNB0Tg2X4Hf2OxlvSJkzt/EmXQvdQGLyzdm7dQv62Gl4CdgbR
ryb7341PAmuOpgaLVWgTbSDBhIEEvpuOVp1e2bfUmH5M06II8QzWWirZzt0N0Anq
cPq4XLnwZiYwBroiCIeFi4PB+NsDN6UyQh2qnC6wc3JhOZMqHmZsAiu1DhAUgmet
qXZgyrFQi/Lq8tbfzviHvq+6nSxPhPKOHKj5PUlKHGzZX2htLnd9lAKDiTcQEll2
PTE9pDVxo+XiA2z7YO+46/7+mdv2r6Uv4rMPck9BYcLKbxR45tNPYL+E3moBsUql
E4Fu0BrBwcAAF6qcswByW947BSwpoAVbMYJg96wNtwmSLs7GPvpedLcwcdKIYRg3
iFo2iX0RVKQpSPd5U1J6Lot4Oj+GCy9Y5tq7KYWygcrQ0O0H1VnJ+mAW127Z9K5G
cqy8dhnqaZkar5gtXNBZnufWCvflrviP5tLCx2xMRWS7D9PXzfmyi2HUFaD9EgKI
RZsd+xsg78MshVtY98Dr1eV4sNjimP7b/m7t1v2N3InmXpPvcUbdBWpd+mZRzNrw
rf6vdGJH1zNQP68yX0NpQ0HnsU2G+8JhayZ2xgcnu94AfwmBLn4Ec+YRfzO2u9CX
yFv2hLSOySkqlRIfk3ZptEPD9pxjSnVrc1vYPgeDrYhcfLV9/nGMECSZ/OR5GZ3J
Es+9FCygOvgW7h5KZXTP6zcFGdwML9mcmso8OIOY7wY0NsIQb7bEbLEVMgS9BJer
49D42SJRJh1ApR+ZbAtNFTDdILr+GqJPnaLeFasMQQTrr4WF9BbQforLV6Z5JuuM
ckGqpj28uofXBw5vOsPwQHDVxQ6wQqgD5+s6hRfEE4D4KJdwwMIYH8aKOwUDitq0
w/Hle78gzBB7cNpViWTXgpxyK8IT37WwqVXHNgbjqdxFiH1gUEsiNEfyHyKyeKYr
wrKjEIoisyp5EU2DjRNFlMHRb6BHoI5Gyer1cjwD0rScXO5zB84T7wKdK5fu8Se6
0KNJEVk8Oqm2O+SUG+G9d1o5E4vGKny3YZDjiQ2BE7yYdNtH10Pjn0eEBsDlJfBe
wqUEFRoyXdb7hQMdgV6CCKYJPwgCTqzlkdoXvGauKBvW5frp+HcJtUjV3Ilz1Ies
DJYL/4HKZeV1Vg6Al0hWFYtf7g+sner1qgfv89Jey5/vcb1dEjM9uWWSNJ0nBprf
e6P4w1PVsdQU9FOcpALEVYfNaxRNEnFx0Z631hlbblEbnMvP8JWGRYUZY0qCWG2h
89J+Z6jEuHU4ueeZWzX1+Hqi9OhMcNURMHAraEwZxZtXFpmUEyQvh8yF6midVXoP
7dx21TiTQxdMc3hOZ+bUTbuxS1iipOFv9n3nEvV9D37zjLSrtFXqc6t9bzve8hZA
IkZ26H64z6PTHhHTuI3Cph+emevXJSonpP1wP5w7iYKqRd5RAwx1WTMJhlZrAMiZ
j3PgqIh1QYtIfXC5r+Afv3k6uvCyX7grsr9XB7YcrZWHuZJTMqw2fGohqneg1dpT
wa7+KdFa+0l8hEdYuw/OImN/S7rusVKpu+abU2eEIPKYWxzjAfVsF0fvrKdy1rXx
WKoK2L9REcSQhqP+pPHZnaBSRjLB2ieQjn8Rfii6qkhO5iaBmMsv4a7UmPNE0GQv
NSJY1t7zFBVLoEjybPGv1RBL/4qjTPU40OYwI0pgTmo3uwPdMAzO/Y6Wlv6QD5uN
Gn1amCMgyX4KEan/YWniDU6ILIEaIIM63MPTjW1YzpKm+LzwOLCHclhrywYXnC4D
69k6I1adF3nebIbBU3lGBvCKaiJr865Bkyy8VfBPIedw2GsL8hSv5ueaKdjA4LEB
hgbA5oFYxE4GAXrT+Q1WknQtUfK18EojOnyEevFJz+gpB2bQaIRGHHb9gaLYZPth
WSfFrMHm9cj2zAd+2t8u1FslziDPEV7ppOZZO93hlr3txjnmF63kMX3oLIK0cC9j
YHCUI6aV9E24Wnh4H3jTouyOWIhz4oHfn+kLf1yQK95pD2TIpDtPI2iZrTjR9cOS
ci0Jxwc+fmROFmkEWDp74J7oOUkDXGarsmreBFT3UulOUgAMgZ0Fro+IUQ59bu1L
vNpmqLODQ+iATGiZrz2sVsNKzNFYZGL3v97B301RR7yUaIiNV6uAPUzPWZB7ZSG0
QinXC3W3pwI2WtPL/0YCwg4X6tgOUb6EN5D/dDKzfEFYVCkSOzvyt6TP5AJf2D+D
tLy5J5UsXYfTWjkxSxFmINW72xWUKYYUoTDjNl8JcxQGK+3IiGAjELRDGMvXtPAX
HX8ibQ+R9VuSkuCCGUk8KzrNxM/dn8nGBN99BVwnGlzj0xaa8/AlVQCZGTo//3ym
gfagYHAiRvzzUevrFlpBE9H5RQy0n7Qpa4J/+F7WJCuuMOXp7NPd2zAuoaO+yRvi
jy1vhj4NMUYJHN+xCcp2a5hgvWPorBgWhq4/ORPt0t7Ws2UuyTTP4/1JI8noY3Op
XPVsOtucoRUdl0G00mymV1lKUIp1HCCi87eenHdu3aKqrbp4YN/mT31OKYCZaGGU
dr0JREfSRPHWzFs+WNdZH2/i7EZbtAPRANMnzpfMHF+sc8ZrD+AWUnbKrbC1gNjL
ISNFXO3T12mYtl3W/NW6CjwsmccNeDG0sjH+6edt13ER0am+maspLzUBWzlJ1H1s
ZV4tKzrVqPUchYnId5ENhOt0Bi3oGktD1q5rDuVjFlRXH4aWjRbCSjX0A/vzOE3+
Nff4uP8OFVIo4DTs9SA2woh+aq91aufXpS0GQnMccU3TVEhs/F96gUfnIa2uxwRH
GGioz1dtEmaJ3MK5SisnxuGSgH4d4f+dz7lwKvsEIRt78W2rvdfOjhhC2MUmntzT
pvoh7/t+h/UYxMfbliI4rFbenjLu+LJNpVbH24PA2ubsJTJ+rLozxuiPPw1I51FO
CkP6CHFcakm7SMBvE83zID7JlwSZPTAxgKEv0GsNvrDb+bejfE5k5Zk5VL4DGX6K
KOxn1FuJiNZFI57T2roXyA/TyfmWrbb1mCDFTeqKGwN3EhwwnjI1A6V9ySLHzJkD
hYDyvNBabR/XWYwEfP2QwJnOTc0S720nJZ51z6DiQOLv6IPxmxabN/VlnEGfKQV2
ntBL8VMmb+Wd7uAPbVMffsC2mVsqv3WbKOAJOvKj7tslyhv5SKLgUb+2qu5A5FhU
ZbRcHgKTIX6Io2/k0Hy215xTeOod082VqG8hQnsFAaTNQIG5EJfDMSPVVmKQr+M0
+QYfzA/kDC2F5tNKlTetCtOYk/YjX2MmTghKWxyT5V1ij5MmlULN88toYu5egFwJ
WPm74/vgeB7PNRcedps3da6JtuPootCBpTAjE7sH+W4m4yznUU+Oe4lZYxQFmR0y
oFMK0k4OjU1+6VebE+WW+rM37LeCnmdMKGie5DYsZ+CGnV2O+XLInQSGxBlLQV3l
1LqqTvnC9wiGbWfnbaeXBs3TJNrSVQQ4H7sgyJ55cA9T86F7nInL+kgun0J/AAmz
/HVTQ4jqQLh4s2APtQbj7QX5Y7q8RS1QQT7FpxsRFe/JuyR/I5K0g886NGxPRH6Q
yjGGb9WB8KnWpfutRr/zAF2ze2aHxJlymBXtRWOkJBVVDAuGO20eWF+wmlUIf4M5
TaHCh0dIoyYKtNPEbB+OCyUwKjLJaqs1gfOPQW36e1S7dRA3W4rdaTbEAvaJ7qmC
3cyi8TN6evWQi8olBAFiU22B0dhg8ilZKaFef8CYvjusqnR3/QyR/FY0IdRr3CPf
DlG6ebSBV6gy2LtlapQifmsip6SW5kI1Kd8MfcHowo2ivxA4t5b86Qz61cLVWyMW
gpdXmZK4suVkOQA07O78llpGZjzi8FFobRM5JsZOrXR8Qu63ltUChQbK4aE5Kikj
2dgodqL/LNR4f16KApeBXlbsW+HIPcxmcPnweGGC8nr5DkZYTa7Su8ooS02abzzN
wFoMJeRLLA+FykelfD7+8WoCm30+ek+NgfYdl1T94lPNbzDG0r7/lBVgf6jhj/5W
oRjTaeyR6aU36DkbqPctvOPiSPWTUD45CP3K0yYxElFVLiGsbHX8C6ys4eeZ6ZpI
r3IvqyPDGOF9412CnHV28VBqWhgxhrxOFTVtx+AatOXQ2MJW34dFMhifpOGWNABf
p1pUC2+1Akyt/UMD5YgwgXsvAhjWQXNm/oRjzVkQj3QLaQmMJBoSHduEs0qmWMwt
9GLSmYR92rlGAVw9FJCWbFSzHHddOJiLH35iDJuzAaqQnyWRUnRJr5kveeJV+GDB
IrTu3RrX2riewk7U9+ncX6SYOquywn98GXJBHqAk1Wlguo/NO33bXYyvxSTKPseL
pK8e5arYpD03+dZZ8pY4t5hotm2xjj6pwDefcNLfgqi9CZ4gb3XR7Fl02TcOzqU2
F3QqSbTAamfs8PPTPJSH5lMOHJsjR7FXO+xuWCiWGLHZ1ltQL4IB6x/14EsoEDTZ
IbyvPPtKIJIuLAoQe8hJ/1Vh+1X6r07yPYSh5LtOO5huvtgWfkePNkivlUqRANa/
x/zTvWFtXLSYSAFQkcIQJyJUZD7qmXOMQoolX1/w6cyDe1kA0fBGfZM7QFTRqovZ
pYyYdg/be8d2FCfqHXnrjK3+1XBW29ubXcYafyFsrl6TNOYmIAFa/U2MwgLG/uZA
71RxdY3BLPCOhBqxCnBb32Za75yuc98iYCAznqlQoZZm1qhdhFZHAO842WCEKY7d
ub3L09TH7o/kYmN1xCPfETtb7AtKQMvY8HdYXjObTwBcf3ptxzr4xX9rDYopvO8Q
04OH/sl3r6G50lhgq1ZXkkoIliKAdMxYAP81M5X/P/5G64fLo1aX/lcmke/Z7DY5
nEmmZOOPFvW612t3emupDUN/CAd8XCQRMntLQb/eVuKbWZY+3fGYwgrsF/srWIvJ
IH5uAtL9/Jnkhc3DjOKPGwP5m6YEROsWXcLc2I/1zE1R5DAeXgWj6pHrhEJwfP8i
HvoRlh9Ek6tP8LwObM7LVs1xlIrvHZg0jUCem+aA95Pxc+PQEaIP/eznFfa0+IH4
a/TdQIUi4Ns7Tk1dOQr7s+fjUpoEIkZnkjH88k2bFcjuR04J59Glzx8TYw3k9G4o
jyTd3NnNQGHakxTyTONYWh5HOWhaDjPGAE1+TmtyK7+OXPdBxdn28drP2p82GF7C
QeQiZA+kARZWZErIxTRR9MS51LC2twdj987l0gA6YsMuXFP7IqYBnskYNbkYD5Zi
Xp+ocL91nzxuaXVDufSIH+TLt/4oFHDGXWt73kzTuSHcghScBAHjjD+tbpS4LubP
utWkTT7W73WJw1NBJl0wccS/DQ0ReNtShbtCASexDSork0oSkTEK73RhWjR2aZ25
qTkceOHco872v+OOPwiJR9cIsrTIR7BOZ5EhkVwZ5by2sIQVgU2lxrNI9SwQsDnr
Uiq5xwY2lrzQDlK3v59ZgMQ4/QTL91SD691qtaaFcvLaHaIaqkX44YJuriBW3V7G
PjyUFCzn981M/1h0GjQulD1dMYNqWX7bSe+55fmFif9o++EAZvipSqbkFLNY6n7B
wovFewlnbjUaEUkKrZmNjJ1dHkVdux44nQDMTT3XQs53rhGYeucZ8ZfvImnA4/fS
v35ZM+GEemCZDfg5dbh9P2mT8OUygyB96l64DAqhhu39e0kD55xiLWhvdrCM32dv
AgnQGzFxx3nt3JzUzGbOxz0WAjQ+ap6wOafk7ssKqsNp7T0F9UzCcHqbcsGlPQiL
zsTTxis1TixWILTYjPIRs9MvtJfX9deJpjFIcbUTz5SN4bnM9j0MJA9OHYCy0FhC
+2OlkgQYnZ7/pxGkJulXfwI1aphtGjahH/XHQGLPWc/ONdU7zHXQDPTnQ3ivQnSs
nwF51CRNVEt6E+E6sJX5mkIFp15DG3nM6xfSuL5HxIc4lEc7cW3f9uA8HMLn6ynz
9j2RBV1pVhIL9AOzl1UhFMNoiXwUflgJ37Sg/axLgsOQvj7vRQzERYVcZC2//Dm5
wH7dmgPsa2ooy+Zr/WQvU8uKMepU4NAYlJwXtWi9qgyADgNci1Rl+nTiGFmOhU+H
k5CFXjBudImA5L+01GgplsHpmCUGvVQS2mj1Tz4Rj/p/8BeB3u/WXwi7hwSC/m0r
XxAEGwbp1TvuSP1zWuBsHnwo71AD2MXw5cKEbuAkowFmZt3dWKte14BbSeAdpc9Y
x+dKwiyPIMMMxggequvE6Rqm0SvyPw/Tkw9mWtVM9jWAR7RignZ7n2lUnBFtjEYk
9OxWp1fc7IIui6qDmwRK+PWWN1HcZUR2VmKZhPd8IaghOiybaknfjNyhFXwZygRw
IBcanQrmw/bvDCMOjOISQo88UEahFU5jB3Hfcxuahsmy6IVQC06oEtNv19RKicFm
xIRH7RskL6iD+piSCgEdZrhyWqDFEFIroWA5NV4p+gWQIXaUZov5KfaUP9xQig2T
fySD0YVcXCkYWNdotaz2/776oHnneWmaYtJg/YuVzVUyvC4w8FOXZmMpP8J+tJiO
lWL8W95l9IeAvms8S38ZSjoe9ygDi/gx9dLnVp2drEpZiVSMwOIKe2qwlvf5RGT7
l1CSyEmrjEFLOTiwD7/PGk2dbeYo+C+AySg6TKFS78TSPbRnJu4G49u53+2N+/Z4
mt4rFsvE1dPKcmwdlfPaGlBlFO51uhOQDrxuoq9xEvRFPvmKUixGgYDMixPOeThH
PoUrm2+OdgCFz9WKL2FencX+UN1KGAUsvf1CdIjnxIM9t/XRnN8FTuiNohp+is9p
627ylcxYOh/PFJ3mGO+JVC11PVfcmuPB2R2nZUB1GEjXx8lrjz7VekMCSTUuktfb
PWfBnBKCR3N98/jpQuuZppiIHFO2agXn4R1YIFWtaSMmXeOPMxMvDfrBKQtwwmuh
bE7b5vYA0DohMqHO8RA2ZO5ShxEIjV+Vnu7fzHgspwfydl/pUwVgpgWND4+jShKX
oELE9VHE845YIt48xMgUWqHoYvUJzkxcVkWmgfHFa+wK0kFbiIqR5LsHpjzpPSPi
OwL0rCvF2bnhEUD0tjuretagLJWpEDZR3KYKK8gpvPtLRrh1APyAfXqpMv980OeW
M20QhbUhsa3PS3tT6XTxDp4tO5E8RchEAsh6zVYqMFAUQJ/INl53Drj7ZYWGkGwf
+FcU+CgiX1fFTcsQyx0R5aikfzcOx/xX3YQ8HPKOGhdTvjBurXqvF3xxJk5RG2gs
kCgJknONZSKOdRBYjTAV26lsCBhwapnZ0sgh74NKKNCXEanIbsEp8ypzl2XRLnoo
XuPlHkuFGjwJ1DnAgGwFCIJbXiLrBi918RuaG4GfH5fu7nU+OMPXyYoE7tOIoXFJ
PnCsYyIQN8yNYRFUBloKb+gTjYXIDaTqhld/3+SYauMOMEyn7lAIXRlh5lEynqnu
4H6zqSZWcb617nIdLCgTdpYtnCzqxdo/FXIktx8s16mKf8ZWX8cg+fk81mfr6H4Z
de2cXTe1itzMaoWMGSp5ZGoPvzIAkbA2VjTLLm0bSMV35q6xChYy4EAKnHLfQ19O
PaKDD6aoqn4T9oIfwKtxyB7KSd38wka24TAFl4K1S5JYSsr1HFJkv85FJAL+12BM
TuySLJe1eHcZvJhroDKJYQ3m24BRIGWQSH/AYqZZTqYevviGx8k5YI0hXuQgIFyz
e47vpjs5/V5iLTljByfRojPf1z0rOUrz8IRNmWhSMOepTeNqZlzCbZAOEvhZ2gOX
r98mlCH+NO4KKFctMEPvGsH+rzy8dp8WtDQDdpuolFRFLipnRsDfXomOKCBx1VXx
JM53bAx9ujrmH5jyhGYc6DZ3jCiFTrUCKFvDP4EhUR1jblFmNyHORruT3QHeQd7X
N/LgiC11QGDt0AhL2YoPadEvZel3BD1CMwWW2yIZRGvo1QPR7Ud2uG/Ce9Lk7YaB
ih8qhsHE7GuBlx/QU/uEOYXGlm/MtJYmGVnBhckA/oSO/6z/u7pxZeFQhhPT+y2L
5Wb9ePxVpo/rDhZivkvSxUZMwTiLn1JD900S9/IkASv2XOFwS5AwMpUxeEbX2Rq0
553iZTZw4k7n3W0JivA6/PE3gTte22juYPl0aUdEXbhQm4GUG2T8LRhg+3wJ9//O
JrX4/lI0KxDx+qpYxeQgrMX+8+/9oGuqJI2sRLnkhFX36v3kcqUzTzE9i4nF6hEY
NtZtwZnGVvvHN0fvYALFKrwuSw+vyH6AxTQ2lB/0xGXY2fdhdoFg68rMDJTdKOKw
uC1aZ3d2xyk0LLO8slIcjrITZoyCOushzwI6KrzsXbLuCMRW2edI2eP4DLjXEzyN
NpZQmJ4WEK89pzEnJMFmWjpKMekEebgtRsiBj1uLRtAwD5M/A8YSBpe51zQym7Qq
wqLcQLu42VPh7ZesWuytd7wtIJC6M54p1QHbNC3IPnaMTj1ldQcC9KQavxwLRuRn
welqqzUqjQdAJihpc7KNs+DgeTJpV5yfTlGXPc7GeIeS86kk2AXLEezcvbZqYLHy
0Saa2VRzZwgiRK5B/dvH7xZDSZeZ4WEuCNF8PA7oWrh0mbJoM8nYiSzaI6bixJ+u
m7tFpS7+/PTU1akJ7FX7CyBtchH4xzTRNYHl2IahuKYPNSeu3HL2+1+azk4CKUKj
CvehyNFAY7F1XsVr1qbR+IGIR7NGAT6svnZ6Xu0xrl9wsivXN1LzohZf46h/FeVn
LgT7u6oRr0vOpMD3/pFLDLaTUBRLchy0XGNDWBQcQaR8qXK0Wj7aGbpHXzjAtWyH
ZwuCG/rUESKUt1Qd2L/eiM7MrX0Mk8+OLM4gVSneYOOMA1uyaBCjykWYBF6tM5qS
kY29QJthkGvupD/SPE78Ba9hmbZPmCi3KB29VergoO4rXmTWUdal7LFeuBLyq6pU
tU2d3L2dRE64V8n6nAksCZKALOf125Elydm7s4yokKvB7tR37GAiKWy6GfwfGWT9
6or/lmBtGh1lKGp6BNhvrVPUSVjlCd7GaM0MrNjzJUZcqpacpJw2oXdBEApM9hmu
3xrwuxdfYA01kw9Mj8ocVuWpqmNftq7Latcjcx9yuXPuVZAAQW31FZXwVv42rWgF
raMBhFyIUzrY4vcd8XMPmVkMugB+5iKjMk4wwXDKdWGJBBOS0xXFBgCw+L+wNgIz
mTdpxV4U/12mySq08chVYE9EcoQEJBVPCipq+3rv+YbgCOX6WVFjC82QVjhOkaqk
1o2fp9Q6MliFaz23T1K23/SoqWrgsq2F7itsAjIjAVOgwwZFEQOBpnGDwU54OY6a
w/YfVyEoraZmo6IULy/ldkPgeK72crKbM4E8c/tlvtmqvJrBSkv2zDVJXT2YXA+9
2pF3p9MzT+ggfOIJsYmc+ydGCaJEewZVpQheJ9p4lfOGyM9ej12C38ZcYIQwGLpk
J2wQJ9AcbVBSd1ZLv182gXGZjkJ+dAO3sVwNYbYP6wkEpFleWXnzIOgWzgmeb4VC
Zg29D5U9mBuInHdhWVujpFfpF2j+diBiTS6vshQ7O8pQWPo2M2z8mUVEQYlVuWGo
ufaKU0x5dD25L5+a4TBOu9cBnmfuGGnYPciLJfdAUIRKiBxgaInOgJEYLSDd0Kkl
I8visnwyuUROkUA7YUcCXV1AC9TQrdLgHYh78Sq5OjAA5+vgXFe5UeUKyKK5jCcf
zzRJmvB+P3YIWdMZcgxwqgA1qvsPsw81ogJlvrYTEUS2L/I8QXL3s9jVe8gyjjsh
0rLgEFDGoXodkWCXLdj9QLRbiydt9A8o49TybQ9JxTQdv5KtWDGeDjao8Df91Z11
lieh2Dcfb/mCe3sd/M/m8Mag1/p26JvRPVH3JKNZ0y4eipuMaYgVtEzXYwg8W+YM
v683WCFn1OEpE106oX1J7dmZGYgvy7ThYb5u2Mu/09ivjDb0KSyaYsEDE1DE4G9r
hxxuvOiI52rNxmEkcP9uK6t0P1jnQiq9Yb+2/269o2lqoFJ4QSal1YP0oT2bVnfK
0RHMtR7o8Ko365IxcLEavbqcU/akzG3moizkoPwuq6pBXJMfHfBs317biuHDNXXe
DC2RfmO9S7JDi6b4DLXzhFd0jwMFAJs1UpG7DCCB7dmupM+fFawed6kPzKZ/rzL4
UKrwOEjaFsUlhpGG2+jFiTKwnJB6/jFLt8/f484xZYhn40pQdfGlGYvbyc4vID9P
x3PNrU2sgBQiqvLM0WMa8bizJk28NXBLxIYgFDC2GxgStvTH5zr1XaHfxamYKU5L
IHvWDpnhYCCpRjlyFH6lwiv23TnQ3j0E469eUlr16aON8Mf8edohIpT4rDQmkLP8
uoBpAzCoBL7MoTjRPe1nrcRDKvSeuU3F5cMmEzMkLg9/dMAzf+15Pea/VYq+Te9Q
2U0FTWS9WQECETwy5dFcTv6YrajvlXOERvR9o8VGvr8gxtyvqFTqOpzVX8a2wTbL
2v4yjq9yX6xl+BGGTwmbQnuXa2749plkiynMfcctcp3SGfQ7NRNLO3T/UeH8kyvL
zIWJ8jFB0bWHdrofFL/nrSNX9kOYTakt+w/3tpPftm8Jw9wWfxYDnHSbYLkBkRDl
+bzwCMPgL+JyKA1KEj5Su0/MfebflPCVtAZW4u+soiw1eiRyupy6TlZKYMUv2Dxd
yAqflPF/G0Tesrwi+RCIm6oHmfPusE2X1KkLjU8Mi+t6b2KQTAs0b3LCf73z4Ik8
ZM6ql7FmnrWJes8lmeI7GXCP5RDW/HEKsLzEiYnDziO/efIotwue99Bt2CD7vIXh
MCnwtLNFuYxtESeBflRAzTRBiqCtyqbC3pM4SlEppXiBlOEvj5Sq16cQsx/eSxqc
QwQqYX+TDqRxGkIbJMqPQBl901z9E3rkshY+DhsIaQ9SJbpF+Fj2Mfqv7YWndP/2
dxUTEZyGA6Y86PFwAvxkbxwvBXM6uy/XtxHjJBwmloRN3IDp85Y/M19KhuzOM0MB
sU8koCmnwKDE2Tp67dMZQ/D1iPKcFyp5JS+WxWLKinmIwaTPHBKAg5ljLEL59Ppa
tjjf07f/+FAOk7aU8Wy4k/kjpqa1It097JnK4WlXLzcHrHIv/47a2kXx6OJ7pInr
HAiD9HEUK2XB7RNImagWvbrw0/45jrM6BGG3E6zUslmUtPrpFDl1O6xS7tbQnpOl
un3To5I+aMnz5uFGGsY0pi9WJtJmtdb/e+uNIE2uBUn5rrr5M0hnNM2WK16rO3yH
lO5pbAJzEE9DWljDQTUY4BZJnGGvv2OAONrrI6sNKErQnwN5DOJVcMJoUJoIhoyi
fiZt0y3R6FNvgEoYTXldQ3pZS83F8oPwXJYsqs+qhgxNurwnNYZ3aFcrvzWnSNG8
biv5vC6QrpcyyBrBurFcohmdg61d9U4ZCJmzQthZhDCTrYZ5Ro1e8e3cOkEUdOPo
RCQAk7AV0GP91xThM9NyeIPX1SdueRMhx39kujlMXEHwnZdKhsnqBMfSr/s2L8Oy
H2OHyenIc/tcxuyMv7h5Mj6CoK7IXHRvfDGw+JJ1NcrKSA3r074ZojDLT4I8SfyN
TzJl4xrvXndqlCWvFzgNDtkBGpewh7Hzpgp2LMpI596pwf5Ih6ewrrU+9CGzCnXN
JVhwOKyOJTMf8m3mJlCTeY+sdmg+AIM15uwyrk9lPkAQGphEZ3pMHZm16DSr0DZb
71k44RwuAkDlJ39ULGKvHkOICpRKwQFgTvUZuhKlJgLjzu37KsUwAzsVugxgyCyo
NbDORcyIYbngUhuBZ4yw33wBEzwCdH/4aMkJ8wkFH3pBuezazWYjQ0lWiupBND2Z
UEs1kTljz0i+yN5LTcuz6oTv5N+uJGVJZwcTcqTzxhGuFA2YqiNk5ZjZCUczgXu1
EQe3wpOoel9UUR0RrRyA5AU+54Y7AJYxNb3DR3OpNW81QfBNxswOdeuo6j9JPZAI
AEUN+D2qbKX/kj3DkLP4U2Wi9FBPWU0k7SZUcW9DTqDZ5EC2mz4E/hV5er9W/Lv2
BnAMrfIJd1jSiA0tFykHYQTwghz5QMLf4vGcMEWZnPe/RMINV1z4k2+AKcIQJ+km
kJEneESpA8GvhFPL1RMFupJyOPhEN2SfF60fCburL4lrx1ztXtTUKrnJfBkOnfks
1ZPFHnyfA2n9rcc/2NKreOsx+UCQ7G/mqb/TkJEg9brlSRRtchudV2WlZhmlBw7d
xA2RTJvt8UaPVeMNfaJQHtCjYJE+CB3PGIqiDt9NDsqTtOtYZmbVZtw6HG/HBTZm
7LUybe66mqSWSUQkw848xj3QTu28DSYpS7+u/ruaZgx4L/PUHR5HbZmFVg3JnX4f
GHK2ThDPhDhpaTpfl/CIid53SQYTfah3FTIAnOTvhLaFZsDk83KUDeCu9uYiawSV
+UPko0W+esWuz0kL9iSaiBMQPblgjTYfrHu2vhLqePm5u6ZG352HspnsZAUP10Gf
JT/R2QgHXM/QfY2VCzBXknoBea+ZicUNg0GPughJiKB1obPZltCKkRsSIwszE/gh
i1UFZ4vQB23wm7wdOxJCpBL12rxqrXGvP/RROZO3E2rpAz1Tczv4SJS5CN7Pw0XT
fwvtaJUiOhjAMPj+hbJy8kdyDHxB/PBPyAT9+Cby+uhX2G7jVQ1mkLJPDEIgPL8f
AIIpykuB5X98f4f21Y+biVZyaLejM73+csVP9anipIcAcI1NfPSAnDWwMrw2aj4A
hnfx/hFgUqZU5IjpmM0hJd5XNV3bMRC88CGQlf62qotMUliP/RcrFZsVesmsbfXy
IajUr87iOv9ME4UAAAcMogk4IqPnWK+ohhkf/MyDRCKSBGrFelP+ZCGykmyx09+D
svlSg+pACKUV3DYtktcZ9yn4nndvg50YY4hEOqmJvFMIgaAtXPcR0vkp/UR7N5K6
Ww7t/OTarYCh/FRBJf0ZgkEue6d4kohwFRShZ6UiXN2pOXHiw91O0qgGskrLG0tZ
K+l9FDHTyJBTY4uo7IgL4uoGVStIa+FrqjmhMRTB1T/Pj78Wb6XFAQwRwturDUkH
5BW4wfkETjwYPewej/X0EdBdbPJkR9WvClfihK7UvHo+byhvS1qsZJMqeHm6e439
mvitAGyG0YmJtq8T/RhvJTeXx70MDQ3LwIBR6nqEtSucwm+eNIlGHKpRyICytDkI
RAEEZdB+DWwIom6FjNvOII7Vd0SW6+gB9/CGy0qzYg3Rzsxwmyf+WTH8Ipbnjh8z
kE8mHXTMZ/Y3LiSJxc5g8PsQkB8VhI0Ap7tK9MZaenMQbTcsB7h/RVwabZQ3Tjxo
wDhX8SPt3wh3uKn/0n3CrHI3FwCgTSeD5bY+u2fw3ETmJ/PSyelUCpnBqFv7aKuX
Vili4l2Vz5GUzOSt+l3UFrlGkqOys6LKxddRiai/5VBdxayqqmi29wsFWGZKUqBM
caqs9dqyICPRpt3PUalJ6fDgh369Dg4YkOLkrEJbip8/zZDph2QErPJwNjS9uI7e
A5/yFXE5zR1EjyXrEnBybuNn9XntxZpnctEjQJMpVMr9mruFzbIfoM22Mehak+z9
QlLGwySksSToWEeVEVAfuS2TGiH5ghNGNIass3f5hgpd7V26xCMRk9rNrltNS4cW
xVuyZ2tc4pcX5M7Z7XzO3hGHEG1W3hgQmCiHp08ezcFN1Lh0DNeAJRDTGdiT/L5w
2iVWLFP7QaQDfukpdoODfa3o7NlhyPemU92XAlKsR8JJtTcYiC3rVfzklfvC0hmd
hLT9zszawzV1RZz9+ktXG1U5XSYSu4Mr/3Pt0Y8qwfnQtfjuF5SjarAK3UnJmvMx
Is/34XfkBOyDgRvNXqIThZqS+1hDMGJMvq+pWDQ+xJ/ro44V/zgDr+jJ4xQhQDXs
esBWIRUu9vvXJ55vCMZSSrf06NHO9MH7GnXydipHdhIBz/SOGjhTUiuyFDEFBz2B
jJfNKXHA3UxqUK+kzkAKJFMQl5aW5zVv1e3Ru75T0XRzujlhH2HdYKgicUKVmxfC
vbpXzJR7HBPc9lwOmhOM3QdqVdXBwwX7kr/lF7zCir1hlID7jQFvA2u0v0FtPimf
0aXhJgnEf6AdTsWyqh2tb510GfsnNkD8VIiFRjcbossgWxR+Q4VtpEVWl9hj3Rtb
XHH1eQr0AfLiOL3a8q3XicoMC7Zw5dEMH7L6r4EmwPnxUHFRZMEfwnXlBmi6SIF8
4+Q6AKDjgd0FusCfrf9alKWRpavtKflymT+f9A52uzk7bVpxckUkhZ1xAPZvzfDX
tm/40xdMHfMAxIvUxD5yRp8ZZDLm3SqQk85dIl31cTO7iO4YSMp1GjRnrZujM/5I
bFQRriG5wPSu3nswBAOKJrhkposUoDLoqPTRh9k5qiE4IF/ncz1QV2jL+pRu3wkT
HjVqj651jOyhXo8Bo/v5GVAtkXe7pkO8j2758WH0CfiDkyULDZjsuAuqT5O4UJev
MRvkcxbxmetOnpJ2Jpd01g3pbpCK1RIlqOcISDud0GYsEf2Qj2LR+/s1uAX3LwIh
QxtZDoiKsjBGo381p/4ohb2cKkZK5AoF4oaCsh52FvMCoM2aDZMniwhgA7nIyLmG
mZ+Rr8INW3aFVkOj98ghtKOuMy4X0ORFg+Ff/vMchLHCRE0bV16vY811BLaHojqe
SSacH60CYJIFasgkQmiaZzkw6UcXrA+bphfixoNldqLautTh6RkIM42b2aTVImgO
pEBeo1drRv1tg7kWzHdPQqMt7Za4ILQT2Sc2sclLDeadXZf+E8UlV/bQTd+H8qz1
P7nDrfOTB0cMyCjYnigFfgdAHACHoFFo5uFAZ4AwzULZT5jnbkewpmPF4fe7iah1
6lPtOSZN1DwNZjlfBjB/B4z0cbfM7W/JOJ0CjfuhDrETZz0+Yhno/lVSlBGr6fh6
qPKQO9ixcIEliEkGVXz69tNRyrvkq0Umh9MfOdwoBEnh4N34H0bjgclYkjGnCrKz
ghK3B7fU/a0aaxpyMw0yTboDE3Thkn23Q2CWVIZ03fGLoGZyEgcOcGO4sT12JjBn
zgz4nlLUWFtwmVF6yZlNlWtHBjQV+mPJAIr2o8cNV6DiBSl0pvJgibSTaGd/IL6b
TnHoABo6vSs+zh2H696L5XP/d/TDSEyMur/YDx28jZL0K5n6M7PDsma9d2d4zq3a
l8T/S21tQwaTttT8O/ukUt9gqyIyQ1atk4TVJ5f8n42WM59cP7VCGSzfwyLa8Cd8
M19aKwIaHUdCv3S0XoBqBh/sEXzhdeQtjnS0/tsRT+ep/MjCe5okTVY6urlq72r5
h6i9eRoqx9+4dhVfsRnkXcP1idXF3Ufok695m2s5AxnAbhGLFxuE2sMOy8QJeoEa
t8bvPsNphFBRgAe6INvSCYBt+N5/hspLyVmY32rNdzcHf84jy4WDT7CZTE6vW6aW
RpRcjvIKb9weFDHhF6ZMzsxbCGO+E2lTuVcMNu1zbnUcEo9zwi8gTwPnZjqMfOVx
6XEChMuNmqfqsLYz86E1Dh8TiFUnz9GJFRDJ4vJ3+lGkoYiceGAYFTJyg2eogcHP
XLNGf+DduWz8RjNpdeHHQulh9APd4ahJPxujxy6y6Py4T90O88N411eCL2ZjjA2g
DgDI6PxBiVf1DfzPYAHuV+xSLPr0p8O+fgk517tQeuJRN5/6j7r+tD1QcCm25edx
VPLoX7sofuoeEtMnShylcTMN42Oz4cdMQdim3sS7/V2GIZpvqq7xC6/D++q1j0Kb
cHGKtjOgJtLdoAfX33O+W0PnJ99Nh33NTzsFcUZc2fgbWFXJG7hgOuJJQ/26/CwV
QI4clZNsumHGLRmObbfebswelpIK5BGLOIcm4y6YO5KaXPAn5w9usO+4ih28Mmcv
ThdUhMZLQ/xtF9zT3MGbC1adElskJdioUSbvU4BUKziHMTGglWZK/e2AJO9h/oSN
8TBgfvTzr61LaaTq/SGQtoteqZ3AKUzDVCqjya3Hdem0T4y+k/ax0z84LMqlc9Kj
wxMm/ldHSnZR8f3O0FIdVGNHG2K7MxBrRuTvPVh3btnX1d/82dqQYlTR30QwBm78
LlUZ+x0+uG0uFyQwhkDDoFMdGPsJnnjF3VXpyMBlBvsGIIxAFtwx8/DtffU15AUa
XhtnlUojlC4f6aKBNo/ayjIuWkyuJ/jDNAvuEuTUq9OacO1WtsMVpgv9aaC868Td
QTm+LXlmqBjcJL//u6LAuYgQjxw09IBi4gMyBTXM+bWEji7+5Lf/1z/NbpUHjtOM
vOPNlxFKxrp4m0seQH86I2/yz/cBkovnu4AFMXHI9uxeC+VMo977Q1HdfFc10SGV
rSXs7tscrmaSVmOizzP8Sz8rX9Nh14rKXLNO0dEpPZssi/obwnS3CdLVtEHxUWx6
QzdzB/r/1I3XditgfYBTn6bTJecZEt/mw+GcZvcXEOmuo2XmJ6y5bZA/2t10ct/b
lRM4PCImMBSbFo5odcqW8UamB9Vij28syiOd4Iiz1mWVbvp5INxg5VCX21G4+ydq
2UJKL4wrLSi0a1J/Un/L5b907OxbOQKG7oXy/mR+8V813fc/aPokHIDVQ/I170U6
X4JjqMwnHiP2hEBfEfflKQcX1cSdBg2hLHe1oVUg0L8l4ymm78aiDjv+DbDy+e6D
p4h/Z+SP3pHtG5Ua7joM7zjsEVfkVMCZr52iTm4PzmIqciE1m42Ry/sdRxxQphCN
qSWhkuSU0fSzyqDCdSlkD309TeyWVM7MWG+00mRedySNgDU3yKNSIfZ8+vmPW0mA
asrrCvCvd025DZndLqxv6e/otAlDw4MLhX+XiIJ5JES9/VnVRw/uaj6aubga8e/c
TdwuDz9vSmHzkHDXK+NJl1RRGOyz1IR2zuqJD7edSn3gWeJubGnsDT9ANsVBMhnf
5AHM6gpcYOWdakl9mGb91+6UpDuYTbEQsFi4zc45mex6bU5c0Vztch9D3UaECFf8
C5wqtx45/l7vUqGzLqHaM2AdXNqGqF4plmpgJO+TDzf7FSuvEiDErSK8GZ9G/zwK
iPU39dVFPqsYHU88xDhviCzQMKXaxFCbC6nOHNQnHzCfNjVDPwg8/CI2w2HKAf7M
l+sRAwZXW3p+752+80dmfq2XeFpoUn/MAa7Ji3yWHPtxIEAWd8m6rGP37fGikGjw
mnbKi1cFdziru9L5IiM0N/5M8mnaijf1XVB4GnmqTaloH/AI6G9y0l9oSGnDNe/q
huAzqgELuL/35QRArzNS9PIP5r0lQ9lXGXW3HOYKl4MaUwmc7l9dvNBMQPzzGv83
JZAksHw/n//DXWXlonSOWVVGB5fpeSYaiIj/DdgcRZeQv9nLSq4/gdqmrFVFefcu
5M//mxZOo6lrH4+X25/ZjSWEWzQu3XqH7+Zb1EtnYE2Ka/SzkHJ0Lg2jJ+TL96eU
vdQsIAcobpanwDWbbVLgrPGprZ3IMeGvklIMLmSNaWcro45wpDw+4bp+epAFUU6n
r9yRiU1LtDVUw8qonAzU4F/lKLUi+bJy/+OyhYwO7fTyfAgPeWSlh5Zsj8HlQt0x
2VRqZNFarJYMnc8DYeAK0bzTtBkAzFIHsWKcDHsUijpGxUODkOKyZCnRA5TXfCVT
D4cCqdf97A/JZImHB8EWPhGE7LrtyuQeMDGiIQIi6C5B2Zr6/X40v7iGB4G1Nsjv
d79qPI62CnlcdaQxj1KFzM1TGY1wYRZAz4avkCM3EB52tywdZ87Ajo60bFrzfQcD
PRb8iGNwPrbw6fkhPepg2ID1AOQrp4MPHHmqautnXTNKJaWCRUiYZebmhfRQmqcQ
tYQMdx6C7T4JwgmdT3cCDk76QKsqeMe2Tp+fxLmZ8ejKBj3hdxkLyL7JOGnHi1dw
9Y1QhaSWyCsecJfjnoCNtgg1hXk1XytmMx/PxK1iNOTVkd2V990E/gfO8XfS1tR6
y+fZHzMaRppwzCxSdy8VtKPcLG39bJ7Fioff0GQc1ARQTW0puYQjUcaSvhI26rOm
TE3NhoPJuLMUV7w5OXEnxiCR/vnYNS6fLqjc47nMK2wVkyFbOlSrz5prrFPMR1Vq
w8OWZP5nYGNGDCXsv4Q7Dfc0IEcahqRRF7SilmoNTQQUc6tkxGWqbGi1shkSpxzF
2hmg/uOqDtj/KUQ+oOeB044bS6u7e9AmnzheH4Ix/jMJGbXuRfX8lVKv9LsDDeln
CnSXcoMHsV4l5RL0FpoHT3HEvlnRaE11DNm0+V3GpveT8YbJlxmZbYF6480BYshW
UCrd15o72d2n82I0SngdP1rxrXrXe7lajFVNezruI/83osuvuo1o+bMAfkiCjNvI
F+wg/nm2nX0VzzFn2loHSd30lFSTrheEIpKhZps5HuSOUSfYa1WXXgF2oK9g1JNd
nm4H7CzDRrWvWYbssdvaqwsGbPdaPHyUj6h1HjqAL0en5LoiTHp0ASEJf1c4oZWj
6IZZGau6cU0LCBKiN0zuoHv9SNcbndSC0sNlGhP5rL1uV9v2Qxbq1LpoMhJ4W5Vr
HiFVF2g98CLPvI1ktHitBphMWW9vEmegJ4AtyRnshy+kNC7Td3LqIOjRXhja7ByW
Hh7hSIstVZOv93/SzfmQRHz8ZvDj6Uwwd7gA5aYgHe6Md4rD/rGZ+BVKzAe8ZFek
4Lzi/QBTtL/FFIRI1Leagtf8tYWX7FlYC9sFzMjwXhDo+efRdJ3OqG/+bLjEcUti
57CGpZTbQUW9sM54mJ2prbh9UJ1pz2CjjXxsJrTvuM5hTQbUH2W7jsikRtKX2aIJ
mTuWEbl1OlKV4IsY1igZOcTGAYBBe88YGzc+VItU69vwbaKpzQvSmK6RGtgUXbnP
aFkRZ3QTfVcUMpEvILp9g8AxyOEG+8jSCKj8dRlq7TSnf4koD9KtsUbT0zk5DRAH
8pTQ+WX4xYfonCqx13xAGBUjxxGwtoW5KG4NUycK1Et1vbqXlcHhaPQiWEOgF8hn
rcQMX5gSdfpsVM6KC46vpEFCbdhveZedy/Qom49mDBRl6p4/RiawAuCLEkyin4kw
WiTYQf8ZHg5LQXWvQe079s58yXNnycHCRYgYLya1UNLC745TQI8NzJx9BzMZtKyr
zG2BBdH+wRK0f6D5Wzxql1bcfQP12sl0/nQLN65E/2+MtaTP2DlfM1sbK2jIzQtg
3vG2S4MgIJdSBFj/lW9mcpMBl7tr08DYLGe8TqIOmauDCMOgWWoOWQSQrbRaGgKm
7Jtf13ZuCRq90RhPJsOvGVDYT8E8bNo9oEm1XUYfR+UfpeX1AnxAhJZj5MR662e0
pAF9NkRx4lE8SFl2ayunGO5nB6yzhlmtyJvbTsViXqkAGJzcGZzLoglY7iGeXG0v
G5aqRasrL8lb41zf9WyAMYHbNKC4WwXr1STpHGZOiqys9rG+JZrtMY6709GNzh/U
tOKOL/65NoKs3oU5lGcE2UrlLr8DG+G7/vfhcHfTZ18eLEtndR/6CpgIoBKWCihC
ZJ4481ti4zdKYqKb6U/gzPmABz1jxGrEF/clvKK0gO2XH1eFFoNro5z4AzC41E9X
zW0KHVVJudQPHWLUZYa/+E4sMy0CbJAVIzTQgJLzmm9YyJRnYYhQxflAUsMfkKau
4M6kwX6kkpieJobkg0JKnTKxIfrpL50Rze/9eQRgUFcBAruvb6l/mkbSV26UIot1
VyFMVBDTxvg5UMemo2CKBs+ICatVAyXbhSTHGSLPr5G3DVxWZTA0uU7BhaeSTKcG
11NuoJABRD8GsyKd3oKTA3IAXZ8PMbfCB0z1t+VaNHI4qkq0VZyKiFsJPSW737bV
hUXFn+ivZrG+F3Y5zCHNS8Tg9pvQR1g2lzLqCzDpj9rrVkFYPb6khdHIRWwJCAOB
n8mXkvjIW/q58FQLYW+XpFVpLRwZkKmPitPFKPY1To1oJrMcVuLjBMt7wp8L5+CH
W74r2GP+VZ7CjA7hBDdlpHnOKIb0DjKVp5Suzg2GobmL5tE7Bdn0cTl18D911ecb
rFZ6wkgoxi8AkVvx0EGvAjktmGlpQ7VE2+mdwAM+A4MJPSjMkAW5ggKeVO8D2TfR
FHDHf/XgpQAgue4oBpGE6xomUE4bLqfC9CEJenY6bFNfGK5tiVUIP7WPQ1gFM9Ju
wThmeScWJvoh9UfZPYfRB1aZUKXnp4CWgr80xNELvyhXct4DizZtAJsORX5unqiq
Vy38BXMtofRwOBDBgRm0hj8vhzLUXijQWJQS9SPIW5n7c52cNlwtay5UnEaISZdX
G0wCft3eOQ5Dn12xtbPWfgeWuy7kcC30nJio4COxcfYC93a0TKOETW/6+TEQiPRU
A//LNPJZ2x/GotFOi5RA0v73ZbfMYzl961d6rbiq2zPa81SSf2e7c+NYMGf4PtjS
brHW7kI8uFBOueIwSGMXpL1FSeRe7bG/yLAWrb6Qus/I/vh2XwsErSpHQYdGVO2M
Blne/28Qf8LI8clfsQIVK4MlgXiyP5Nuyx9lLbfVvqon1q9OTN5aDu8NhEAlSgmc
yvUiUSwGQ6/wAQpnY8iaa+vH8G6H4b6f/2hTPlNLQPgkuIJsu52ZZ2BFlF99H6pP
13YD7/4x4SIk9rih21Fh0TPyI9AvKDCRQkojm1m+Xe5GzI3A044xMjES80odP6ec
xygxTdtD9EjrcDmLrmZOTaza8688M7ZRlHHl6XSpUoHj/Gi9DK0yphW1VdXMU/2k
5v0GF+4VT/Kw4iTHuiI1OVcr2uo0NaAv4MNx1MuulOG+1dpcq+63LFG1/67YbEPF
03vqAIFYWR24nIA4UqwLrVo/uIxqmDNVuVTFEUIcBIClrE1qsiWbKDj1RDc6ayBF
7bZ9SLDk3ZXnQvigopr7IP04ZkqgogSGNBUrfSscNaooyg34mjiWitUBLoGQ1enh
xA8obFDgpRsCyOpwmYbRly/BneLSraSJB4Gp+rApRg8MyjWK5QovnrIfJcFVLxE9
xsBAj5JS1EI719XUsA23ukYvLqCPDhslcdUy4n87CYg3JYYRJccLGfRzisfK08C4
9yw4v2ZD11SgmmzMbNVZldY3iRebeSthNVFWaqJOJRM2MeIkM6gYcpcViDduRybu
4LdvSb+SKr6aJmoyAePMgnwyVsWQFM2Ae1FvlC7KnXn7csdwf8shjlviMQ8e5oNu
r0neGH2RLlU1pfsluvaY2cGgS+QuLV8BfL7uIdC/IiH5KRPnbZ8MeKB40Dmg6yI8
IeDPxJRkQW7/4oPDeTpgCJJLbBlF0OnhD6EFD5RBqS9FLVv7FDOBb1hsff9FbvLe
eQatgkOPQimBt+o+x4xmnDm2CUQf0aaehRE0N2A4Zk+A4LETaFpFUCyyOo6Gc3hS
Z9jhm/zSpABEJwZve9Sl0dGRxKNLxdJWMJLfK2vygYi51ONyEQUedS+fk+2FjkAi
X3fhR5Np5WrXYUuue47IJjrl4ighq/ivhwY9sZ51LsYQd3r20i6Pf4CoDBx0+RSM
7WoZTJzrZG5/ToEAKbliVRyBfSaSLXNmnJva/BvzWrI5ClYzFXe/VuGP3NsMSHQW
/m5z1fkkG8uQ8SWFeC6uy0+K6myorWhJaL+am2K9ZLQQhW0MXZorvQqAMpuO+FTp
IGy4wQxidgyiD92K+5GpuVEDrrm4nxss1g0BBCsldpvylGuz+3WmdKmPIbqGlY/F
+ythoctBDzWm0Nt7aNgC0JV55b3JJp9rt2Maacx0rSyBC7IM5Kzm84mvmC3cv4p9
cxyqgUG/1yP6S6ZB2Mnc/9qvFwMKcXYJH370MfgCUGbIS6DPHDWV6XT1o7uyqQHH
wO3FAgoCjZkOQ6rr1mQLZTkLU0psCxmn7LvnEFyeblevJSpF1MesTRfjpf6NNZxa
NAN4HzyVmDL3EPBUYEME19Ao0KtH2aoL4mWkp+hQeAUfOI3sWcLvzf0crca1nU1C
ipQp9bvbTkUtcGF6WISomfPcVyf3r3Dj98+SRVFQ1issFXrL9ALgmdeMpfnIsaAu
ApXG28rMhS7Xq5fPuKD7NHcH+SZHjCiBQEoAsGKY6/qylgn4QDUKvCC08mRFTa47
hB96kdN60YAJEU5GaY7o5ZEZncnRbk8TuaI2gCKhCAe5AMb6lN+OBT7k8fkSTCSq
7uSscwUKVzos2BIDN+dtOcAWzx86xMA3D9hf/UyzR16r8RR6CUeiN5nOfGhie7Lw
WxxY50XEvJ6hptccic/gAMJ4jXg1e+MS06VwBm4870WuIX5qTkjgcC3DonUqsMoz
CgJfVemQI1I5qkh7Y40v8LqXc+DKWW0b8nSkqecpWxdFS/0ixDZcAklr36CKiZFz
WQ655Vejr9oA1AZUktLGK/Cjahso44Mw1BfSnyUbHs/XGJ9wgniJ2mzC0VtAJBf2
w0fxhj9+tTj++b4E/wAUm/bDhGsya4uBS5HwoY95P8y+X2lhkqFRWQjt4jNun6OL
zt26jaHKdHJHXqzVyH4B9daU8ZAOsBobw/KOpDWH5OfWGyPAqkQ1etONxjhfM7yI
Zl+Qe3dKrbgi7+7O3NapoY2xuo3c2UnVKE2PjLc+HZ4kr20VyHT+oQ1TEwqbMPeI
CnCallsnEkTcBlSV6Ae/0PLqTqoVECDwvQNEF2POzhM8c2emJkpCbV7bICfrmdSh
aBRH/9Q58nm4QsPvblPKbzbpP4A06BfLtHUjBOcR/BAAIsCnq1W6rbs7dLbVbrZn
ojwOEdpAkXcLzAWCO8cgv0hJ01gOoFwf9Xblvyi6skpiqEBT6A9aVagVxBJe7jMr
8CXG0PNxnA+wYryxC6cAQ+oc5vQi01P1HTj44PG+eqZTAHgke0MBroDJsrm9HrgT
K/0fqkdB+hQuEvyE4mtevLlmgaNH83BMlRsNklKUdbuQfPPnvyeo1c+URAxRw/Hj
bkfzR5EOeo4Foe4AqQ4EqnuRBvtwZMrR5ZxWOHvoyfo5gUX23LvqTmUW2DRCXDWa
VqU5SqIQTO4IDGAeE88cBFxrGWTXVPNc6NLPv5dK1XKP45DtGE1MszK6EjYt/YfF
TNVhwla0Xh4j5e1JgV5rxH3ptBA9pbZ/9ekW6S3IFs6M+d0Tp1d8iTz3DWJ78pAv
yPq+4izif39cBBmvL17XOeyGEC5r66+2HkD5ZxM9AzKtNFcSIGLR6wYx/qESuD0h
CKByfntpGgXgQLwX9SNsJtzVFFI3HqU8jVUPE0Y/0aT7+9J0zD2f+awa4jhYJka7
NjOIppscHWbtXyfFpk0+zDmCV3Lw+uTWiTsV52cqaDHyNDXj40GSKv0hVNbQnH7R
6el490Dn0JkopENNryLhWIWt6fFIMNcqTrUFjjiMpJLNweszWcEa3NhDYKbgR8ER
2UEXcScteFJ+MVO/4E4bg1FE/eYFNeUGWc5QaaT/YoQcDZXGokuZrfB2UArudI94
QRm70VUSzuNmQnnai48BHLWxqRtmdXJZex2MEoDZGoHQQPiT/d+HHu7DlutsNNde
fHELfdExXgOKkXGaZcor0fJCcY+JVPjUMHH/wH0vhKTzEXYTmxJ7r7rLTaKlvire
kV38snuZlGXRMGwf3b6XVcszY4d9pAiw5W3PgtTEJEj5RDXa4LgKpGMHR+a2hXi/
2yLCpnELcTwNtxUnIznbWB+Y0XorpYfedqjAEN89GRuiXUlwXcFy19GxxRLlmM2R
SRiRNDgfrbPAbuKhpdbZvFu6b74cczi0HMkciOQQO9zq5K1pRbqDbOrW7Yb0YoOq
GVr299tDge1IOfzXWsYrgGmb++3cDetVZQgxxXA47rmIl7JG4VhO0tCp93dKlpzL
043B+2T3qqTIRgrQiHSAaOS5U82z3E8S+wDpvD2NW96c/qbAuwgiA5412C8OqQt+
A4VXVsgnhnOrNoMDwgmxa7JjRxXuG9BxezwZXQ3CFeIoT6ZJ3WkKd0oFT1Pcq13y
iio7MUcbYc0e32Td8acIG7ttyJ2ubrrt4Jsdui3g+wCvDIWKgEU0mFefphOjGegv
eac1va0I7F7rC4VPD36/q6DGckI0DP3zAfB/5Y714cScUhNEB8mQSpj7oxCP64Fg
t1O00NOo8p8tEGCSfBVa/XyhhtXDZbN7QO4TVLR7ZMLXIg+f7p1K1OG8526KC55K
3LnHjpHmHicpKN23agoLV70Jf6oUDC8O+0cNRGohB98VGI2RjSzgpFv2fDxVip5U
3YAJJvVekB2rmcMHGcYpHENJNiOCQ9ZFVT7T4q1yYyv/rSDcSDb2+F6E4E2mCW6g
+JQ/xDgLIbo1LdmSUNhYzwRXgf31CaY8P9PRHZZZ6eukSVLQB4xI29MonD8SKOou
kni5YjXxnOw9u23Z51T4b4UKIY/eEzy6jmd1MUQR3+ZawhTW+4whQfSyIUZ1/8gB
l8ZRH62hCxGMcgz++y4wPMNhcAMi8cqCTCseu1GRlZ1Gt+soKSfXPkLGlSSJyG4S
Lzrr6UIXc4PVDTxy9nFengb45gW7v3RA0G6X/1xfzePDJP3gnQsy1jkHUyX85stS
nOEAckMjfAnq13UAXTXOKLhgVMBcgZj21ye34sb2lWW+/5TP+cLzynUHQt3XtIfM
igl/6OWf910tatmu2I2OovG3IHsKMYbuTxf1rXjQwF9506uRlm97UMLQUoWUK892
CBdMkZDQ4lwy1jNJ/RTAAI4ddBtPYkwhm3wvTV2vnWsyucA3jT+pLPJWaQlyDOP2
/2rEEvdLcrzDRGq6abmZYKd3Qxa0RQOsuObJgbAVFqUr6FEuN0vD8fZpLjOPbWM5
fG4iceCIltKd8P4MjqWcyr2lgjBhmRBhgNW/gmVOGjpD+OM/2wyP98+V1LHkFhBm
Ls/yfKrF5wNicU/rwKFMYQ5Y/rbVc2owyvhq15ZMY+TzU9wq75NILLAVfXXIb5md
ybyZamQpz8td8auR7tkNadXUUnsSL/ynXjrLzrpsP1xccP3H2l7c3FTRhgY/S7DD
KQU022xO8sKvoug4Kh3jWElaUkt+RZeBFrcrySoB2sUVDsqgFneE15EHHDCwl2V6
Rh9GoF05Cgey3sRZjSSKsGiQqFtOsmgmzn3QNbh+Bip2IQpbs9QgA1mge1HKGi2W
P4K8+/u4ej8rhK8rnGFJMWgJg69DBZpL6Z75f3fWAl1VPY3ByTj63Ervz0Z2rQsB
LyYfbLrrPeam828fNuqNKX4TffshG3edNCiAMg+E2BvnGUTX8XBIi/yqonFb4cGp
hcx+/nCM8qPFiYCmd5FYXA7FAneczDP97UT41JyWuofDDieG5iXvWkBk4YsJbY1P
RSD9zvkwn05SytOSsTH023P+6eCM3aYba1t9fGWLz2Uy5owZIXWJ5AHXxpG5Aptf
HCyqDRh1zimQnf5taU/tdi2LD8y4xUyzEKFlGcYCFUASNBriAvR8tYUu7YgB63Dp
ZGCBaCvVwmwOAjR7qrDzqgnDD3wDQU55u54Gjo+2KwVuGl/NoKwfwB/TktHi3ghe
vvZSYLLx8fixSAXaZ6QN1T+5bc5pkbu9d5u7VhSha+joLn+BowUb6C2+ldVN4qe6
p+6hTf08vFbf5gj3uDDsg+VrS2se7AFC5aSVNONwcfRW+VT2a4US19LeBzaQARm5
k6CfFLBmk2oO7E/kHn79oRkcmzlxmnAY4eSuVRFuWrC+eBoIq0oiPRGjFlG7Bhbl
hpsaASW024TlgZw4Nq4nP94EypGz4lGsdCRQIsa62slJhF+dH25W/T55EBDlK3IP
CfBHA4Ss8IF/nKmYVVZVsAyxORP99SVgZ91JxwLp1XyKiZYH/qITTq88ZrxYilld
zBC0yr/oii3fVOlLeNx5viHlz/s9kUNlS7h7JudkfYl4juXkPhePCm+FZB+2B2A3
F3gTWI68ndC0hU7v3CzM01W9YJY4DHrVw0kfGLMNVCqIcCxtUqyfIYbOCplmwLNU
y4vzHzmTyM2lef9iA+zjS0Dfrx14YeB08NoNv0hyCWL9Vdd0tc/gQKgPXRYinaUm
9IM41SJg1lQRoTv5VTT+T/yfnsI1smEV6i8OaYvBnh11BFesOagnyDHnNRM1YhpI
tMym5EqwGEH+aKGQRcgREs2Bm8SlFSse7/DDKySLNuZxeq//kGhqODCN6rpTGV3/
kn8Q0EvuVTudN7V1uEiaTG5CRNm59Lwbz6pyQz4cpACDxEMAADIphkFKBJGI8PmV
+MkZChmAae6NvbZ5uFnEF5pI8pKsiFKjDLCb0j9C+ueLkgnAmMlrHW2I651NGnwc
CADb/RsGZQ/Bsv+1kGf0kD+0lVhVqhmg4dvhX8YswvHZf0KighieEB/tueAa2Esx
bJmlqwkBMtVIKzlauWqsFFuSFR/Qeq4jQCiyYr1UhCg3ED6jKYh1UmIBxPV51yTX
ANYg2jPu+Ko8xvWmH/+dsSAb8SOZyXR2Y6mFcTtq/boXphcl1FhV0m0bmwoKqiOe
iaJmL9mSRNq5tHizINk+MidyvHYoktLl/Y45gRXObP21l1oPIgD2cvdAzGOZxLPA
JlwPSV6KXZyS/HaDAItsJgwsCOcxZGXIjLQdNFmViVDB5FKxI0/qNTIHq02uHgo8
zCwYdUFn/v7cIqlUSl6iLh+rAcrem2/bja0ovnVTOx5FDll5KJ9GkJ7/GxLsoWze
MzOCipbWCzKweCwWkedWkchC0HTIRjDlTOjACGEDaPrTV0GB2JnWIleE2sxMi7sz
nvOJTsjBX9wPYS31f9nkIhHg7bbcMfg/VstpGNb9YHA7/yZ1XLu7M3OXsGcDXkGp
vDTFib1Uces3mIEnTlVRCXqJN94OVHbK1HzjALRozVBfCkjHBokN1Bt51tprHVSV
hJomI+M5qEzWje0kv3C1sbm+tbZP9KxMAUPIRZ2OryRRAyZvcQgK4g9cS6LMR/BQ
OVpU9pm6kHelwMFnVKwufaQnN1u9W7OMn+hCYMK3lp9FamC87433eow0eqM8nJYX
6yRIuD2KzfyCU6JZJzPRVvj64HPu2EMLxnLXFnIQyuVZg+I3HnBWvN4rj1f6LUOU
kdXQPX4F3Z4Q04Y1Lti072b+vF+mk7/xWSY2R9/Apc8z9/a5RMDOQ7bbet0NNgCU
tIQIlh2aGpyzGRn6NvAAvPFZoF1B4PuYioGBX5M4jtLZe+qyy4MTUq5y3153/2Yn
RWuKoPeh0P1+rjA4zpCspM0jC2o/s8kdM1ZqFfDpIuZjevSMuTb+tosbLSKGCEwG
AebS1UZQ/ZC2wV5MERnpp6a3I5p9lKgm8QMR7tsD2xyOwotUYD4gt6FMuASlo3UL
xG8PtNHNfgzrvZ6lYLnhpci2SUfdRFGYeuOHMA5ddJ+ACe9ZU7HZMg6DiOn7J6Sd
DR9CIoDloAlI+xqg+KnFrFtg8yY+PjF+FfUCJb40wkWXCh9F4t3Qvs2PmLNo/yCy
qv7X3TS7zNUNlB68TjmWuYhLtwmn5FtTRnemrpmgOd/LwKliP1FhP/9DeWqPT0d7
upSTH4xksVxHr/krFagupJeHiMH4sRzX8aZ2CBVcddkFlw6oWm8fIMy0OJtMqU4m
HmFuW9J4Szw3s6uQSUZA4QKkc1tYTo6XJHruYcW6XvWlQ0xxRFq2q/oIwARRUyiq
P0NfznAIA/9w/EFVWzuYMOZ3rVcKykTAPAJne1F1WRBF3jtsbj82+C7dcRBLT16T
FNOIjzm6qwVJPzGHgNf01omnCoGQSkrXGMsU+Fmq4tY28SGHB9JjDO1pPpfbsKnq
En1+ElgDQtyzym3+EjOd7/KGfp42uuXBje+B3ve9kQQUTrPGUfbfE+DuP7CGn7wO
XN7T1Z/GRLW3RPbVE0Vphs4Zcft1HU1ncjewgIQ7wh2pYN6V8nvw3SsgPiEYeW6C
4AClG84tzXHsLSeHzpJiutVXzjX4xm+MLoc1vpMTsMfL+IWiBSSRcDvCyIA8WDSV
s6vt9KY90W9kQaYT8e+6cjBruHXRUIt9nR125k2MqT1BUlgyLh03z3xrFE8o7uPm
3uj6OD3Xt6rFd67r4DMIWHDWSU4bT22QHVSmK7qJgaASMrxq/axxgkHQ4Ud5Qwql
F5cl6btB2PAxTbv3/F3RIQT4NONwHvAc4kwKITEhqD7MoBIn041cpF637gZ0i05T
Wg4C7gtuqT9A2G3U5WBmqwwZ3UM3Q3lI8n7xzBU+oYAJ3l6IQiv6uUleUfwCg77I
EoAimx85cR7ToguExp+rnkhQxlwvKfqYioqwLjmTFLc1pX5RyexbAUvVjg5c8qnP
tQIrJoj37jOMAiutVEtNZ/HbwMXX6OMLqsoWSCncxD5serkU4zCRkpaKWQ72lu83
4vD1YbpnrWAAg/VMsfcPjd41iHcHx+6BUVL/vsJACDOK8sL1miH82aiYD0gkmXmS
XP6whWA5YJW+LZQF3yM5Tpc19cTxZXj+hPzVFhgelXj0jXghKEovqIBX09yK1QmC
B2JaTAmhpvSXjHbtK4n5hv0OUDvmhL4qyMs+WmqRrhTBuXvITi9UF0g/ozDq+5jw
SBv9pJ1Nm542hyJ+Ww1Abtd25txjTiZhof/ExypiFXqNyVHLflEFEOtcrmpyuU5y
SVuG8siyOb9BotE189OnUKt09zDaL72EhrTejMDDjycY+tgulwbS8+BsFaRwYaWr
pG18g/UnvGknW+RbnNstvVTj6ZjBRMKJFBkS7e0/R4gKpKYd3If0rC/B6SWaeadt
RmyS8NIDNN8d9Zj84MqK5IXlsal8VC/H4XnN/OIiADyFxS8kHFm8HzO07W5q/444
pUnWP/SSX4QD/Sccc8VE83G4o6s9alre4HJmCLIet75w5Lc36b5fE1kpOZJT4qwO
tfuMAsqmUP+z7LJTN9SJ3o6wXCkqtXpm+KILyuhxrN0dcEdiBajhnzc8eYDhJc6f
EXKjjXEi+D6TlSdLfTx6pe/Ztg/11PdYuII071phTA44Fz2NInNffsiOJWMCwlBr
/KSgRBQu6vj5Xta5PKSU2NCeTsVQ963RF1PBh6icXj1fOfufqjkdW364ZT/SiDLX
eSEGbQzpn7TlxeMrwHwkllp7ln5nFMaQky6P721MISfEAWgxcppVOpgsUjeAWJuz
uk2thg/61TwUZd5hnWK5Q6e8hw2t8juiK/UXLVvAQkq35ZDVcqn8N9Bw4zOO64r7
MOfrWVXOGlDh4O2afp0Zny0zyukietI07WCGyqvdPQp/XBOiS579LuBwijLpDXiZ
IrpzkiA8iAFUYRiAF2IeCrF+yfAr3BDcxQE7bj4xZcPO16i6YYT59hZTfd+Xoox4
LyNkuBMS6MFrDvK38ewvjdzj2jnerbZ84GMF5W56uRU08JdsxRrzJu4ASzCjSIGy
EGEUe8GYrYttNIClLsXXwn0cKjyBvRb62WXuVRuuLlZQnz7vY7GEjwypTSX31Fhd
nit/7FF1R9f2zND+PYTBCFJvGRKcS5t+dLMpuf95mrugzQh79YIo/zFuzZx8w7gB
cQKGyrkyCYzH7BlpjyS4OBU4W8qRLaI15/ZB392s2g+fuudRD5OAZCUMOBkKPqmE
fQotBhnam9ovmSdKVTGpY90wmQVuA7dxUAWPGEu2LOZa50b2epFWSfJe82iiS8HK
KcR/WZNAy+WAABjJf1fIxhlh7Hs/Z65nnaFo8Y1ZqnWj+bxNEpRc+zCW9fToUWpg
xNjslghrS4EXnTYK70fEUiDbkpMdVtndfMURzxVdHWRgCaKZwjDk+W4zwb713zcV
uWsk/BCaRSFKkq0wafQX9HeNeLBnhN0nhoaK1RWoYZuyENm0DeqJQUBeFFGweOoq
t9F88PZ/rPDiALMv9uRra7O6sC2ij+xYVkcyf4GtBXzN5eMPvwIbC8EHG+JMyyD+
BKpe6FplK32JNuBLI4kTEwFnHr3uYDqvT3GV3eragu4bqnzI/3M/egwW/K6qTAiJ
Q8OyzUwj0JN+QtUgRsLhzQO/Y8tuO6BvyMkarpwj285aWnGpnzk7+3mmq52jMiZh
RlhJVIKyiXKgtapPq0Zk0wRT8lh17tYbVxTOW6hTTL+9FL3+O7GL9wwNVDdZXoEv
ZNGISo/8pB5QpJf//oZY5IBWHVUWYeyOoGhxbfsoeSV9qVv0XH2aTgJ5oKjyPlXa
W9iKu4Pq5F0Xaosekwb1vMHiMIZaRXKoE0xjMDUq20Op1D/d0b/ar3vszzckvjjd
/ip2RPexe6I/PN/nQY1Tt3mVo6EC58/gV16rTjlpx80Y6cGIDVqGUEsQ1v8TzGZ1
3INK5PeYGdQFQ4OkMhInDZcjiuHOqRFu5+v1W9AS1+NIdKVnRqBafb1sKzrAmc1C
0IXoSbnfl34uqyhM44zGRWr3BLFy/CSOsWSrSKr+6PV3Yk0bdLPkkJOWUcOEy+Gx
shvVrjJDYNrgghy0uaiYkMlxUTectlvoyBDsuqQwOBNGp22BA1GAoLaxVV3UqNg5
xS4Eod3jZbOeL5LjeAT+ZDrbkvGqgpINqwUb0XxQM5V7VOVE5Jzmk0/YebDfy+50
p8VW5YzFP8th2pMsjmUxR4jipRrxWqc1JprDi2m0dJG7rKZtPZscM0gO6Vj+c22P
udbT0Y4eS/0WlFGmnENf9UAaIhhjrfMBvrZfPO3YEkrc4IxfyjTix/Odka8MKPsx
SL3JydTneK8+YZBU5PuY7veRgg7Zgo/S1b5uAxdrT2iavcYv8bON/oqqQUEsu26w
9n0nCiM6GE6DNVFdi4s/UpcFI3sUtRn9y6WglIp62x0iURF1t64rJy+Uz55DrqKe
Nyvo0G3W49UCNDAdMhA5JaUlcTo5B5v49b1dDliPOQZhpHFzT0KkwMMNsBfWUsru
98rUvU7uM9DPnqUHvHWYTLBrzwTPPHzyE3cVHpaiJ/X+m0l2iNq6Xjlq+jgwG8fd
sAahU4/ERfnAZZ0VbWXalUB0f3HEL5u3esghhx08JKVO4EwBQskdGBUyJdOSmz6A
WYVTLoxExGE0S2DOLuHHIaQL4b8oru9IFeZjgxUlROE5yTnG6qiTxp6ygbMzWE1Z
JDK7smKpxUGrUHtshP354OjpyxDL+A0haqIKFYV6pmMiJZA8nikUMgOhNKPTTLA2
+7RQVFzoA3rtBOM3kcVleYt/EZfUCF04PkT3f7QnhNN6Cm4luVORLIRSBejntnqt
QRdaqSO+cBdLyIM0bX6iORDDTTrDOEnY+3liYDIsxAymBuOxTzkcAFOVVONLX70E
VTqyiJNBxMa6sW1NzycPzM5JJ+Q/KvxMhG7omBIFjxyBMKORTMawVb7Myh8fIHCE
oE0fqtqWEmEjYzprw5C+Na+pGx6DSppf3OZpWTMkyBpFBpm+/CbFb30YkeFiY8dE
6TRTjMnIqAx5X9HQeCdn41MY4fyt+W6UTCcraTC/WQ5X02uUMf4Y7xZKgfB0HV54
V5PBYepuiKdLlhIBIj73FjnY82xpJ/Xo3o+IziC4ITaIt5vV2pKpbw+8vP3iQcEJ
lQhafGRgWvE5lPiAYx+dJQrOJluYdFwpbGIsDdBEGgIn7Brg6FtdMJYirpDhd8fU
cYL2WjniN7yVMZgaFfOcEHakh+khIGam1VnQbFlNCGUj+mZyk9aYWs/ra+NCK0u7
mh3DawkatGTK7PD9YxeAYFlPZOdwocAhyaSI3EGX9OnPCfKIBeAFr6R7ooypOTD2
TY2tVVs1F3jOaiuQ23ja+ZY+Er9vPpY/t+ZrnEwRaqI0nDJzTT7HGlwi4RbY3UTW
jlnCNGrM8DMWWOfnH/9wYAzlEuMM8rEWcKvGezQjBfUq2bo6enwuGPi67ASrSyzV
H2UQSwxndHyRWyNgyOMXU0MoK+tBFbjWrimydslV2D8C93OaIR/PdXSgx0XryAP/
sYy54ZrkKuFBc7IbInnW4LSb8nMCWjLKcxGIzijG5S2amJvZDjIx/CFOJ0TXmaaU
sp6LV4wfZ2w3cb7s2BJmdwQn8nl5zXVQRBL907vtuwvMJDcWvzXTu8FqijU/e4Sd
aP19CKi0Gteexyu9mz/d0Pp/21Cnn44wwyp0iD3fSWbvQ2kcgplHLbk4TOXzjcnA
GpN5S3ZcJvVXclyvcetPBRQNz6qzIUcR5+HVD1f5MDHS1KamjRR6pwX2Fl0npP7P
PwwC6I1fiCLPkJuq893200X/ChilYUbYRCfKrE3z7hogOUti5XNuUBwQMbJ2oE3h
nKT0UZBMz6jsg755TebXszzcVA8gRtslydtoM9Y/D5KtvZ9XwLvuGp2qGfcO4Q9b
gezk9tyjnztlzuVQMrlMtZ8qjZTAZZs/ODmsF7mFCdXlEMv6YAFMSN8W6dikl7+v
NioezwpHfHlHBqS1emYfwBW8l+j1Ya67u4a69J03M3zxboQW3G3aUizZZurstxKq
i9vMD+0igKw/BY3d+WDnDf6WUb5mfR5aL66I1//Br9cQYKBDdvhG0InYObmovNFk
f/F82EvAGVqnReuNheOMgqBSsv/lWdEhy02n/zZWqsZWRDDnhKW2zZMp6VYoSMmZ
2uLLHdH/yWb9gOy9V5lDpwvkRlAWUa+FCEIB+dztG5ZOZEB27OJane+THgpuxOe9
d+KOAE15JgF4VZUXTH9Y91Ok4OsthnNYgZHHnArSe0ImX6a9HkGBWl/yXVavZjRD
hjw2G8g0Lk3oIQuUaVB4GKh3UVj65K6Q84OlNHD8/fTVE6wO7v0rmAKhGGKl56db
c6CxPWFbBp4l49sd8cwsaVS4UKoaUAUqeghx2fnEDlDrNYSy8khsNQRfeZiCbPLo
Tyu+ybou9MCTlXOeXQyX6anshcx51LFz3auAajQG2Fdts34VllcqxuuB7gVhuJYK
ehervJRG+hnYSdWh9+halRtfE3DzYHqe+2JPt04NwrjzpWvUh8eHtwyBD70ZOXpV
TxG4Frq27qlo17JjpTMs1+FDsO8TEsZ6DcvaJrZ1BcGafi9U7ng3/SKelFNDQh/2
tU/egjrKXfcseMhb3Sr1gdK+ztRwHSxMD1nCtWta7UfmOejq60pv1M9oYGMYGFMH
FPX8HWWyJa0DrmUtiF4xuowwsdQjX73XUF9OhIR+ZjH0haRYo6UIenS7jvkOY3s+
luSHzxb+XEYSoBBz0reQv85F9f0lcoVqZ3H9opjbpuXx8QAWOo6kC86U4bIt17mf
kQAsgFX/gSxvaVT8F3JT/o6DIQpiUQioGWk3WzEmJgv1Uvlqfa4XyIebKfF0EwUe
8XwhDUUYWKxlthUqumVNM34NQg7Vwk+rtS5/DZ0M1rMycmo2dQWu3r36otYLT8YJ
LzeiMuxtxLCDuP3IWwKvicXvCAcY+ZFESzGiVBDxdglYLwULs5tlPR8Nj/iH6+9i
Md3DvwSCFlftCiI30vXBLLG+rckifWmZ0EFYnnTag2AknEY8x54Pl6JS94gfkAUK
H3dRlvcAQX41pCJQzPdsiXOSTVBPoghtgqiSYKy2f+dhDLbPgZpWcq+XssRpqrS8
8PJSRK8U2oIFfWKCOXmdY5mWoewzElx4MCxnHCiNlF3cC20kfK5kv+o34oDdLKns
3ZVEmH1kpWCQnS2IKOxku34j53W57DU/D6QsmmsomAujU+qdD8Vkv2G8YL2j0aJc
jcu19UGzOUVuXRGn/dnyd3uJKb7Dve12Ig54lhEYhyEWjIb9ZqRfZh5UVzruSxcp
lgNQqW7zVtan5FNTil6ZbglhaY0oJ9IbNo70whH0fVxqKTgCBngMeXKi5QlfTS0d
oItkHs85yJV5aUSH3GeQfFdOVwxUwBt2S3vZkRxnH242tyzHGZ6q1Vt/zDbwyRfJ
6CaoPqSbxbaVgpgAKGK4IuiCwFZHh8p0k3GbfUOFZoYM8IoBIUr/LX5GdvOx96eV
Gy8ZIthPQmzlfQzCJo76ORydeYncz9Dk6IQ5Hrw/xnzL/9JuESqNHglODYjjG5iE
SVHsVXT5nEWgKrcEM/8yv3TNrLNN7ll5ucE96qb2GMPRaX28rhvl6GIoBVeOeYvB
dcSUXrjnGMEK96h4EuxpcxHU+eIveem/mwydlQH8pT/GOXoV1qTK5Qx99da0uHz3
n2TOXYTVSbtnSP+WLAvBTmRa2iW8pgabjFUAFr1O+5Ai4AjH5xDT/v5b1am7tcW1
SWVHNJI1YWQ26R/js2KzjcGgSRDH6jzgIWMg0VDns/FF1qICLJB9Y8kOjcCTpf12
3UZG4zNo72Dn4fyZ/sHhHh9hQJLIMTEkyGs4OxgspQWiWJrKUKnbvDdP/7F6TICB
iaeOrtnbYC09MkbQiOR52XoMzKYWmSCWu6HuY5UOCNzxeoAK/KeL166AAj12NC8l
8GMjpCK7vri11gtC5Tgd7i4Tlayfdkui8OdFqP93qRdNzG66CqKSA2GqA7+A2zRy
FfaAMJEs+BGFatfqauB7w4sUVbzP2UgZr0uilNRTvCHAx/hDI786s0TQfwJSanbx
qMcQkEHisoM27UoYAGXzxYzKTDfJ/xDdwqnb5rwA5WDhrkWXUjr2HNq1l92qATpY
chsgLKtUjRuAwfLCcYNRakf8CyPIQX89JriSQqKKctBeNYugDuQCcKOfs0AElivd
rOg1S+FdbDK7+VGmIxgLHNmT7JIt8dc2ZSNfXe9iCEQhlOGwkfz7R6xOva0LnRxh
Q2BUeabfT10EobAsrH2RdKjvZ6ot3/q/LaXL1IPsS5k2VRe5fpsKj9f5x8SQO9vW
+OIOtKn532boZ55yt9r93dqJXWh2GDd5mTXjSmT2WUW/V/fLqjm3PFHAxkUce1HF
0AAyOyAALE+/7NmVJFf04eUNEhTvn9DreAaC+HDjkSwynNKKQCoAXM9NDVOY66pp
pqzxqPv3fkC52ObAAmn5UWVGWJh2dWtA+GXZhU+zJ6zL9JWO70GzL4en33Rt1RPZ
goCRUkj/CK4AVObB5kIlmcZn2JzdvtHXhb/bBpfSIckRRQ/jhI/HhwNkVvd1lYCp
sFggYhoxfcCwD9cqJXC2aTkFQepL19Nr0nBCZ1GjQEsOpwamLYU6RiVeVVOIc/Ly
i7JIiYEHJMVXdYx84y8G5pP5kAKFbMLF9TpO2V3GE1lCPWKvugpOhXVBl0C5iCIA
UkoQGbLlSIYjdJpei10f0/LrwaQFSiVgskIGgrzOHLd3v1duPxKMribf8h9j+P/w
6o+S3UixSTmVPh8Hq6CTBL+1d/5ePYX9Eiq5TRQCAoctr5in/A24qwNIIqGnnHJy
4PRqlnt6EfSx0OsM/bwgpYUp6t1TiC5GNW2qmX2lMRAn6+6t2LUEuJqOSKrQ0zMf
zhyGfniauBgrBPMW4whsNql/krfxnitIX9ga30itPbK+x1z1JV0wjc7pjnpz2/ze
Tz67scpCqH602iqxlVqaD6V1jxJwAdM7ptIjZQHH5z7Ov/SNdMyCZEv6wOa1t/qE
70ZZcPcqFBgyCVUOjm9cBUPN8MNZN5xml/vxpuBEW7O5N6h9GMlceHYJ2EFkGw2+
MGH2Pu9gKHGUdYAVyawkmezHZSmK26iSFCSdfe+M2+QYodQjbC7zS1ZPobaYEDWk
/sFhW/fDkxU6otgqjkb0VO+KJgzTXK13/rWPayhFYXVaOp7pdt3HJIWrokmpnvok
ZPldfLjXYrk5yyZ+zHLDt2jJG2kxxRQ3Di19o7ghLxIHDiqxJGu6jhPI7dKgPpwt
YiZa//KUQy66PGiWtkV/l7xwC5sDafha1LEnmPzO7US48jZBO3bZlocrJYxyoQqP
TOlRYU7J4iZrDoOwFTPy9AP/TZehUebkNrTM3UPE+3OqigmSNWqJEffM1JZRcyEX
nsoJ0+hmuHOndCRdfQQnrVI05XolB+WCFnCoXVU8zdqQUDCbXEseoqqm9d12iRZN
z1JaKkyNVlr6pIrJVhSU7C8nvkzkeOxci2+kGLM66h/7kbmqkRtuh5uE/z7MU+ni
5yyd8N9rx5tAcmdHqbkM3DRoV6OLrHfda5Zc9UW0xD3KcttdS20wwb0jdfgE2nE+
2ugYHzeTwIYSxwTI/P+Ky3LtQR+beIqGjUZmggpGRCUtKkAGjK+ciedTpyt31fSq
YnpDiPjSJRhNnDCvDsiTCxLuECMOgrSFV/+NV5VDu1qF/gFgbledELxc1GioXSBc
56JIwbLWhVuyYgy2zCUDa8xJvQhMtzrPRtd5bthPxxvy7snuMl/ks6tw95DS+wqf
DejMfdlG7/u84Jbl+nJvFLAOsAqgeAoqZhP89J+ky4EHvtdEs1n+7VI1rfeVY9n0
VANx6+1zSZjAK25qpR3N8yv6LAIJ4GI9INeSU6zP7SpRX/GDldF3XXC4ApUQg526
+QUWXIeTt7VuhbqYqBn06qAOqOvqeiZ0vjiNYiRgG18pGxYzN1SjMTE00p3NCaB+
p+W2lJlSpu05NtQsf/gxCrvJWBV/FSVCXTGbhI+BeQRegQRyRsgFH0AKCdcfmIkO
27MqDLv4msKE/wWusNhioOhXLAjVu3+dOJdCJs1zyxYVecBLX9kdGgMemXJl3LvG
UoAcC4DDPdAVAv5JFA8n+3Aye7aWA+550+772g3AntWuxu0nh4dbiUyaVSuTE/pa
y4rTicctVt30A6MlwOmrRx1+tdHm5UQNVrZQC8rJXwTOUu0WaUYPnPHNv03OFyNe
EJ4ZMkq+chLDieyo9663LPP6o8kfhDNT3GF6hL+tIAm6GzJeN8tUgVkmmCgbsPQp
RCUrSqcGD4IAb8PvgSB8qVRvemW13UyJDftpsLv0sJGImVeAXl8hELYDM+Z8cKZ7
JfAMqb1irXewxehfMxcJbNX0z3y3DDodzN/5QukmStRIjEMwx0hF2i6JTYCwM7hm
RvSD/JMH6xN8mA0XuFjvLDUKX6DfxHzB0ArM7k1Z1djhMy5XSgYZsnELcl5+HlKF
fReSI8gvoYGQXVPE/fbuFVMX2ONNoeTclCbiIyoiYccu0LKBhfGTPAnGIF+yykcS
m9bdqfsmvYZbQ6NJSimp5vVVqbZLQ/Yo0dbODbJOs0oDQth1XhjLcZSVDFbPeDmF
PeFD1I+vERv3KvDAlcChHioHFjjcQjSpy4cXGE0sc7jf/xwRNKtzZFJK7b7oX2Ye
KJeHcVxsnG7cjNrdwimMaxUyPdubvrOa/LmyBLeilZ3i5DgNbn/HViU2nb6TNhDW
NSdpH2BBGfq8gwSgUg+u8rhCPE0uDLAwAej74pPfDn6kN7+hi4gNJDOjK35YhvfZ
5UUTPTfK1tkHL1jnLTEB+dzOgteWm6y1dP0W3CMs9fEXKaWD1vKzGUvdLN632JCb
xwFfeKUEUlMgVNjnfnBgMhYOuMxcgBX83ofeceVkZ54kpSMsOHk33oClvpzJDUt5
5lBczNI1uwkhPfuctEPemRPHmvGLL1rppvCZLAaY5UkYERoWvjJWEuN6rQIavukw
9c2zm7vwrXF7bSF0XmP9Je3vpedBYZVAma723CEZWTuFABZCawiswzXPOg+DgnNO
M+Pdh/ajUmJoVbwoW6n7T62CJEBtBDusuxw78lox4suoNaB3brDXkQ88m09SVtD4
LjqzUVZA2oy6g8ATOUhVB8zDp0GoU2j7R/HxDWgu1MlXrrMUpXysGF8d79lUOocu
jklkKupM/bvBTyYGV4t/8FqeBOmnyw8rv70CftPqmRE8YwYN1EnRc+SakKbo3Vmz
fDthMeTLJOvmqg7coiV1Kiv0xj1Y/sWD6i2RKafEv3+wXWGCVU1nEVXmytCxjKJ8
jNX9MflDWA1lw1ghVH4Yfj0GNosboTZ05BMcV9HjBb4K6AFDdqNhE652gOO9uj+a
yBNiGm6K/LXswJYf0hWbHno+Hv1x/pisaL54djIW6/rT7Hp5Qsty3NnwQFYz/XiY
tF3+MdawQODTPjEvfE2kGTGtDvklxILCDF8ICzWKUpj/LvfEkAwq49xVGvBZXoBC
4i8JQ/Wq02p97Sab+vxfURAwxBt60/iqJbBvnKWjdHCAE2Q+bdY+kslX0muGTsbU
/a2vnG9PbFvlbNRaUTYCQgZtjgvrO7FoVIp80iQCvfpkPI8KbQw+y1Umyv9AxyYL
BUmn6DtUjI7qrjgeDbmEMhjYInlC24wSwmiEUTwJJvDZnyPIW/izm8crb6RgXKPp
mcTbZe9lgDyjgzbuOG8evDqNpEJq9Ao0yTCMU5BH35stEn4bLfl03IblsgvQFEjf
BhMbGAgkqzmMyXtfIgq+0SX6gRp9vGXE0p00UPi4o5UJNz9+aodW2HFAFpKaEJ1s
Gx3BkNuh+6/dcB5JRTAo8sO0Xjq2bt5eQYKhTMrDUsyP8a0tqUA8o4YnqxFa6hl3
5NDHV0uJ3/TcDexoILCrVS7PvUGWVdsOGOu7dFavbN5swgw2MFqD0k+1EoJhc0bZ
Dn7cCP5z7T1hk0E+Oc2yGfJmD4pj/O8y0/8R41MJT37t1GjQ3K4JvvzDKyecnDdI
NM1/iw+4+jxc4Y+SryVUpv8MT8n2wvzw4CQt9X7YmA8+vxheTgPnT7ME96ntfZ2r
mywB8K7CHUL8FRY9QOkRJZ3B5YmXywGYp/HJ30ljy/R2JmXXr8vOxETci71BAikb
ExSEpHwKEcCH/dW76rRBxoYTn8IkEsska9q3B81QduC+OEO8QuFMiqPxB1PbONrI
tHI0uxpj1SVJyTo7wfUVo8b3oySuiotA7zGaJOgAedBEcc8ji7aRybtb/aPJEC0/
65QpXILEMMcuRhtSEokTVMVDLNKTfuk+/iipA60ytEKVom2dDGQ5zPEVf1xNARrc
JnLOboxSOqs9Fb95zsk3RaUYp7eLj1fYmoPfkbYC+kLMQlJNaMYpR8QJ++qJzcxI
hS0ZWafLGFxNE9MUBx8P+uMOTkh7bFpBpkYnoO9J94h20NGBkKJ0WTh78Jzn+NjM
A523Og04OgQi6Y4cBb3b8NFZoAh3S/BONm19eOnTyBzc0nnzrM8B2rx/bAANzTnj
FMdvmi5aMokSU5hPkKNK5BbKLSJcMqAdYX+opwVw6MX9N8pSbVhk45p1ZDCjQ0Rq
Gvi6vzt0a71MXnGlPLaqD7+mIxHuQXbGGu2rw3h7IHfTIon1UXTGcGL7nW7HxwjM
UPBZMp5NZN22+i7dAwSmiEYWPC6BOyr9+Lu2Kzu6dlSnOjyugejTB/kEGWb+pQHS
AnIX9ddqFAYc9WNtSbHJQU0OEn8+yuBECw/5FXyJiiK80bkKkCtiy1KEYP7hAMRk
ddD+Kmi71VOBsNix3yfC1h2LAqZVOhZKhQuzRYVJAZ0ODF7Z01cUNQ5jyyOFjlOG
+p0KL6/aGa6wqXY3pTrqpbRdKk8PDxr33XZ9M9idK/1JMwNSzswGzVT3jGwxKQVk
tCYTf60zBPXrLYKQE3pQBNvKr8PRnqun+4FdY3Cx802H+0mZqQvaQu11rWJ0CxuY
RilQI0zP38BsOKTNfMaWDaXtGvk8X17VnEOUyd5Zx52NZHq2n7ATzo4RUkhlZrc+
Q8o1A25Dp/hskZL3ZodcYeJNJ6CbO4JCfO3WLXAO9XcV8w76VbmwQ31eUSIqog5G
13TV4feZh3UjlqwI101ZRhSQr/xKmtiY3rkRc8gNH3pSmqEstGiVbpc7kWgCsSGh
oPwkKy0qTGF3vpUSKMBAFP3NK4zGyKL83g78Omv3wnvpvPs39lo/pltlON/FCp/X
7VDxFBomMfo1oKWYF/yK7HFXzQW1q9+dIEn1x6wjAFcfXH7ZbuR4NCw3jEkV3qbU
i4cERXIZE2P7P8mZ4oFMQuAv3UbJ0EbEplTgZD3rKbUgV5i3JJh+XE89pJwvEtGz
zjoGuHkOiL6HxXiRWZN323Am2IYImq90P8jjVy7+T+pwy3W/ikVmGBhGwLv8lwRN
icoMTyf84mFxotWtdcZAxAqflEk+fCUkoupeyAMhyWhpoQB74cdIwKFUnGabo3vF
kiYE6YlnF6au+xceWMQekpE6d2wR79B0vokSgFEGbWBHuMC+0OXYgcK7Chzb6mUB
da1o6dwiC+Xx2DxOIMynlyiRroaNJz8XUhC0/MBD1nMGaWVaiieKiwViAFbshkw+
G0EWAsYFhwrstBosD0lH+/2OxTsDbD8BzOttIVQ41WxSWylOgrwl1Jl4YbRR0GCI
ZJYQ1ZUv3cKZIYfSmY816kIpcfohc/gqoyE3ewN69QX4qgPZvoyEMHSXHSLBIPNH
CYEyDZB/53f2ritTQI1p9X5DdUCMHNXgXAMen/un2nH21ErXr6R4rZZ6o7N5eUyd
pBvWeDjQ2zBeDTfz46yc55Q+XL+2ta0i/uTCjv10aIsuUR0WzrN2ht1DC9ahfXZa
Q0s/FGaSewwzApRGr25q9nn6Ujcjp3DuwdVprsdzQLm0QrGVDC/RXhZVtIp0x+BA
vo6CJxc+bWVr68vKdo+fxlhBkL4ZvfA3f/8i4fSWKYwjYzuqfwF3ggBN7wnkDHVL
t26Bkjo85J3EZDNOHnrSeaWOeIxUT8LCl5NHlZgjlSyUA/qYQA1RtSgKbcOSjAEc
7I73xbRCsYl7IdwNUGh3VyRRD1JAORKrTcfZa3ebzpOCD73jMkRNTC9Va1hd+WG3
ceD9qerCZB9BzVyJ8X8UswCukLIDcYGPTELjBXLwhxmpE4mAEVMdIB/VdlrfPwOD
LSbQ3BWSxPleCsP0BTiZqxXRsLIBnkxRPbzOWkLuqJ75FIOF6GD4pAfPqFviuctd
vvrQ2s/LMUIVOt7GlSI4k7fmEggFo7uOLWHSwA07TuqRErO0ua0XjRM98EGiYDkA
oh76nNnucQtpBzCbkkHFP+tklvikRQpXnRNv4lvXQpkvDZQF6y0KP7suD2eAJRJZ
gMHzhoGqU7VlPkIf91bJfEJCPYOs22cN+BSdnj+NUO9pOtB6HPUcSSQceLVt4Xhs
xuy6/fNaP+aEaTlG/1GuBlySvGgC3DyAwffjWhoRG3Hnu58I4lSbBofLprKyYjbR
85Jq7XgCH1IOMIXm5bsu1uEZlfJ6DyOcgY72YYIANqRp/Z+8tf2rCg89wb8Dwkca
7t2tXRchRYUxaF7gm5Gi0MgBOnh510G1bYgQ0/22Xm5gij9VM0BFTM5ISINJtqMe
m+zetq5T7JKtC64+wMtTv6RNhWxshFB6/wzMQmbSkK8UvkWAJVq0rmum0/J2SPTp
7TsAJi2NeU/NLUl4ssW1lTHPY2Nnt4yezu5MUNpTl5UN7BfSBlJ0qxpi8H2YiZuV
E3EUQqa6FflYemPNoHGTZU7oxbPH/4BRBANwoCO2iVhaMPmhwAII0k2+/8HOV84p
gKg90tzE7f8ESV+sBSpkYFza0HZufmegB6Ui0y+qs+9Z2mBcRiqYLhMSV6/7k/0V
9Vjnmv60Pfw2R+NMLRBROzvVz94slwV7oXUVWYW94aCABEFqvC+fXd38anlYzL36
pkMtAIvvf2gyBEUuk+TvqUpwRIHUQqBiFE3VU6OmTx2amF9PiefU2ZQg2vvtvmd6
MbUzaabrST2CPfbDoeWVD70GZIwswYhSJf22zlzaibusA0x8ZEfgfOezayREnBBp
vCt24l+S+N67VGeQbfFe152Y893CynE7aatQODOHkQvzSbz3xRJ1ChpgOGWH8Cp2
nlldE6/L+2PyTf2d6eAXk1N89WIFtSXvCvylzgFqLZgFtbHQYNpCB0v9uu2zFSdc
7l6Q6s1Q1q7YuUHseP7n1yReVFpZAhXEfgVclfdeJgeQFMZ1UvO1Wln4ycAAhyN6
RtaoIc7vk+l/m7Qh8Q0/KWcyGMQR0KWlwDRE+a27RkVMmGK9/1SqNFzwWmFxofkg
M/M5R/k5lpj+j/pfztyNABnDE7vyYNb/MEi2idPpiwZILKLyX8kfeCWvU8SrYMVN
8xeHJlbqb/yPc2mI2nd9oS8JcTJlEOBrdqUgzvlvfXMNQ50W4Ik36UG18xfR4POA
vbA+pa6sqIvQ1ErQpWMrb2a+dcXcK9Qiy1vlEvjKs/332YZix8SYPNkKxC3oRL38
7JVUiyxEB1J8ZAvfmLpqZdTInPohB2u4RyzEBJfBvOJucjBRUaAy1nX4ptGUpAuA
ArTUOq3nkBafzkEiNRkBGkFzd8QAVPp+PY3yIwydUpEcBHuDQN50h2l+obkWuC2a
ZC0EApfK7qCxKvElUPEdvnQeyxoXilQ01fe9CmpaDAYXFVlkX8mbqqeJ4qRXQxiM
a6PKar9VAgaSDuPKK+XO01/YFoKKY8c+B1XPrbsMNKcZ/FQhvC9hKmMx84t9dTBK
vvYRT/Msv4A31ycGLFskJ3H73dwksiYdHuvvFjFyZIhuHdM0bA76DLefGVcsmO+9
RfcshESRS9gscb7C1aleofAQ58B++JFRR2TU2kSCRWWWYcbI8N/6CufICFpGuX2r
BpQba6nbof4bARVrIuw7MjaMMy2bWiGOrdZQ9GJ3fUTD1JUgYEQkD1QS62tzim10
nrCDG6kM2dtxkV5BXgD3PMxCz30Uf6MIz29cVwWGiiiY9FAK4R5cYnfWSc0sDJOc
14t8wMRzbOE75TAu2hRwrYvOfULYA8fPTgezsbVAdSjljSMMSeZjdo+cUBxMvOjS
9YjOiDi30eypn9BjywmL6qjE1gEQpGXub+KGkVodlQ0TDUDCsm94BXY4UtaiVZ0x
Bf11N0EGkftpbAMwVaCGQz1o23J9SM2DVi1kIHuD2E3Z1QD1Z3RPHIWcjGNPjTPk
UIXkijoKQT/7gdAsxaRvS6FSFPAgsfaqrqBaOL3JsxP6h7a8Y3MOAZ7pI6+fMs9+
ZKzWrCdrp/n+rQ7UDSYEJ9Ov69TiGBW6PUM+VO9okGHWzrfyHsmYv2COXXnNkNHt
kXmhay6G6pHR6bhZDTo5yOThDdMcU3W8MB4ySZfwnIhgmyDcbfZ3g3Him3Y5x+nS
3CJ8oPv/RZE2nfQw19hal0pqtBpaKNdLC2yzjx72GWvef1y/0pRMGzHuYXDv6klx
wZZCPLlhtEYggyqZCHZzzIu/yk8TRrFijqVgMlaKvO8lB0/dF7EobhHVzFuHECvr
HsRAqQKW1mMFbsuIZPxvnbp9rlUTsfBSHfxnggKh/qGnK8/eY+gL8CIz83SBfVwB
PV1vPd9oULTgM5dGP3jFlkrBGHRymkuKSvGOyV2eBvcCMmUXlH4YZDpVyO6xrjN2
RGVwRdytPNv1chBGLy0rutUQl7jm5L46GKKkvmQyd8OvheUkhWRlo10rjKJPNFBa
wPpXwHRWgO6SV4nuwdtm2eB0rYhaAcoXrRYU2uI720Wl9bFMrjGaxKTs8lKOvRRN
xt4oyDHOlH+HH434NcXsHKQ7Plh+A0dY5vOF6t0WLYuJC2Tsvx5iBaZBiwnt33uL
tAK6IPP6G++nq9JLT10rkWDlpkdu/v+RdQw/WzNhnSx0/Y9F6Ez8Uu6AaFX6ZTm6
lP1a9d4GDPIg0hd9EwImiRKi5JOsV43006MzHTipvXBniLyFjAUvFxfXhw7oj2x6
N/FEW5PnGeVzKJgBqyQr/qp/2L1wO9hIY9imVK+W1arMYRaOJrpG48by14yn2Skx
yyNTjbwF020aqyKFLfz7XM66bheNeneWTyCnZtiK8di7C8a4cBXhI9vyJT2J0Qpo
U5RJp1y7d0PLVbdLMmiK+4qcfl9P/2UmcugN+Lz5MDxZLAHdXNm6byaomK0k0M7g
9Ttq6AFpJluKnLVyPR0YXfzg4FN/ZpVjXA/qrSva7W6BJlPvBJSbfb3Tqm8eD+SB
9IxUewI5Re+qTfHdz6KVK+RAGA2oVVAv9TJ/W8f+ayMLTFQq6mpCoDOyy5gbiK3a
G32pQ8QPAtYPRx6qjMD5IMGqU0GgGUVDZCoc49g3QgEFU+2HwxHVb04INfR4yf/b
8X7xFSeqazaxdLAIc8kOcEbrHx+PAbBhAMVLfbiszyno3P2qiDoQHjGO4Hn7/bru
uOYlBiF2+gFJ4Z+BluCy5stE0UwBwnutVE02VOh4oGIINl4vTqWJSJLOXFbKRG4/
IZub0USDGME0OYDopdKYZrgcpzHYjfppamH2KaW1goIkUGPP0WV1kiou7ISbtw1T
L5z8D6Eu6ZokML9n1cfxx64iJ/zOJIlqrHAB8TooHElszXBXWI6t/jNun40e/r+y
x3S7F4JVF6cV03mrdXOmVBqKmGuifddM7VUCiNhdUi1hpiokGB6Y31rTPURC+Z2/
B0u5ST/NBlvdzPZwsES1Z3W32OITWF7LVaysdNSLN0ABdT/YNHug6SEB+3G4tcDE
/6roaaGofznSi+HV93WXlJ15Ulu7wRxSZwoppBErqsCeyPFJXvm/ehpVzgY+gSRX
l0w0/UhQydjmsoQEq0vsKguH0Yz38gp4Dn12jnzBTpQ/Vo4Ybqf9kwqoLJ2gR+x0
QpMGEWsErO2x6ztuDJvEubvoDZdbuKU2ohVOyn+ZNX+U3qYOSRjUAvhTORNwZ6Hf
cinHG+yhWxdizr29mbTBo6H2tfZI/2cFNYoVVYVsDz55mAV96VdUjSAFkbGoRtnR
5MlwVIADD2SqWUK+KEZ04ngWnHTBzG2XaiQvLSI0GhuBtPoWfnQTVrVpupw67RCo
t3w5ajGOaBVIDFJStVPG8H5R0PisfaT4G2CfON5F3zgcGxUADwCWALFfmuM0GGcB
mnOmfsrlLwL/EWXisacxSTe0h9HdJH8F3pjHRNaaDiVoUyqth/2xupHFnCXADrds
YzAE7/1VPzrEeeh2ST/GsLXVvKEvJNRXtLvuWr5vi6/8+I/EjKQ2bpzO//zkXTbg
4Y6Eu9Q+LJmPayeyZaJwqW+tZAO8uZCKe/GyHNH4nWNT/qpaGuPSO+4exlLqFX0L
oEsKsMr2aYUtL50o2dvhq5bgDrfDjPNPD8DDFbmIuUpUeJhkPoYDfrDBZa6d2v1E
BH0Lfq3NilypVGZvaxy2sg+fpGJzgvDS6zCPKiyfgZdCjsQiX510g+p4jdLcIgg0
MgyS0+ur1MUXn1vu3n9TAtQxQEBq3cSrlCGz09fbTeZjUAqoR0hJUsSkSiQmOiHJ
a0hzSgvXCLgaVwrs186OCW96kFiFtIQ8auDY4IATaEOlxFuzH+bfEnBFXUhoeVhy
lngqDZKC/crFqYpVOENbgr3VYZqAKIAY50xgkzD1iq2IyJhwe1DsLPZFLf+Sh5+F
FBvRUWtG7DKZviooacFpzu6e7tvZhaReqSR438ZSfqIRUMJZkeeLRbN0qb16k0JB
+nrwDRcZn3MLqg3YogskFJpnOpHALyLs0wUHHG9wbSDhYq0EOiLO8lwUCCjWaxRh
fhE5J7CgzaiYvGUCpSSivd88zP0QY/Xilm0EBp9kE8ZnApOVSBqE2en1s0fxE7R1
0SqrcVyFa18pw9MAqUrQCepA8PhcRBp/GZCHspRfTbUVVaWD6FjbVeWsC/jyUmUn
59C9WRcqhxVfUldgv2YCWqMZ4DRWQs6lR4QmJwoK3AmNWa00Ng2eClfk8iEfdiex
S5g0WItFmHJhHTDZyH99WHHe0k0T8Fk8ZZqaMT+a3nhKxSHdKOTAuDWeyUq2la0T
rmtEeDxDKeD4uhVoga3miUho0SKmWcRPOal+0UxfkUuUJ5+CmUxzX8v2azVSLO54
OGeYFa1qyGIwSI/JRIxtRwdQcq5zEnpEbcmOOQ64RB7VAr4XIjkUpJbeslvKwGYd
nbzT1/UN/rNbc/+eS33owhBwb9s4hKEPGHfmNW1SfNjyx0TLVHQH75t/d38b4N/Z
d3xFXWy4PHDrBzqg4927WjCbCb1LHWL/RwXvY06sYpu2YWhmkyfS3HkF1U/CP4LX
W9tJ6eHfYGY/S8rERrdCt91MrMni4iUfpeUHW3pjPkparzSAcO/It17y4vrhqKVA
rXj5D8fjq0ytBacKXx1vHShYLsys2Eqrm+UiQ/Lj0ENEokUTfDOnuMcd/L6vJtuG
lizK3RzE31i3RRQoPyJAauMCETVois180mPHs5Qc3O+/nAcAnouofl6L/6po0/F3
1rL+37pdGhoH7slIMZcKy8aeRu8j1U3JwbVvS2NJ5nxL3K25RZ0jq9eoAazV2DUN
h3Aky0tXRL6Y3ETh+cgPM82EChGxpit0VMF2YrRm2BRPJI5BaOzpyedSrsgoOLE3
Fuw87Pz5ifDr+9zXxOs6imgQGH0j/Xq1KAa9myyYbv/J8B8+FPZbiw6AoR4hJXle
VvLs3gec1xphUM+0aZpOESjzi8+SbXlGCtVah7TUVP1DpKzVulJdSGzc39iXMYs9
eBJqQ4vzpBRfs0V0iNTRHEhMROxEXmgjEgZnu4MfMpnaYsowH4nZxsV1cTyY8HqA
MefLCGgqeddreFupmQNQCSx1fKpoDECN7z1r41+dMUrVlfuWKaiSRIzzqYf+bOW8
Lj8aPr1H7SRHUna+7BilX75czKWT0CgDbeAwh9BK//ZUawgGRNAkIBSHF5dGDRyp
WrHQ/kSyL/IX1RJMcedzglWdteuKvikk6lahwghqTEGlSFvZvNvq6M8MDGcX4P/K
DGMVVYEcGeGcX1VYcwStVlgyNzHHRJj6jmTnWVnxlFJR76+zqroqIqGKqi46XpO7
fJHqKsA4ws5mem6CcmXfRYgNocbvGgjNskdIiAzQm2vmrlyg1qqGNzeC7S7cVqxq
59l5Y/eleNlmC6UFtl3N2hGFnRkopWBd/sun9GIXvGTlC4ZadXDDAnvLm+MbCYdK
OTRK5Icu/DLsXbFsLfrisQc0Tg+jnV8qtEdz+BzUHqs14+e93RV9L5bblp37lk2n
hwZ+jYkTJEAEx2yMk1HLcwbW2PX2z1a26SQ1kUKTuOS3Nh6gvOUtybnTi3NEvWCE
hM/yKCOLSyAqLRq/6LFJ1kIZEE7OlD0NqRBk+iiqOgLo9YZH0jtKzcHKeBKvpMoh
YdYy+1roT60GcoY8SHBc4Khowi0tE1ezKw7aX5Uoku7bkBiKjIVEkm6+FhQIIYKz
59KE17L5fgrJw+QpLt47sQurM4UrMmoIZ6rLlH0+f61QXI8KsFbxl8dJK9EzUhaB
TmXdR2tABYovF3Xmj+sYymYxi7pdjD7icrnune3uCCPfpOLkcfdCi5hHokAi8YMl
W9s3TbvkH4LUj+oxDJspSMghcwssvMA+3IqHWyL6SwA6UAmNf0fFt2dKLth9q49D
7TPqJjEStrly0EcOobk4JzQYcs0UHGuA1kEHk+TWOzM7AkxVQSmK9KP6EgMhrJZF
ifMF4ka277Czjtx6XkFoHGkf/FpQtXpk1bxV/5y1mKMGHbwFJ2AxlfBEDQ9HDXPI
cvi+dr3YbF085NiJB4k9hQ5mFM6HdisCx2owtVZdD9WDZEoMnLWyVygBlqdLNV8s
xjvByMytBw/XLHOk6lJH1qS3xDOFhUahOpzdPvqSOv7ZyJU/CnXpTBknMYPJDEaM
hIZKNp547rh/UDpFBRrxo7m6/ggn1ot54StoLTGBosDsFFO1FDTUf1ae5o+6l2jq
oUGRTA3B7NwdHyx2qJGONzOV3fntHkb0qPcjBU07hOofnkW/BKJhooYF9ibULm5l
XgsQvV5r7qAXe6O2qVIKIjuvvcQtsq23llEvLv7vDQ+/MRArswC/CASM2iQztGT2
omydjV47TppFRdt291jfjlwf+nudxV8T+yNcRIJvR5bzgEFuQcy+Qds4VJYS+BQI
wxQcYQw4Jq3axaRAFwQNL5VmCeMKC/OuOSol7xhdYLwGrq9l/SfKje21jDo1xUUq
n4puG8N4gga7lseQBpqPxSrVtOrJPSSLIVBV8cHFeIRyjUSRuozefvkTVceJc3f8
+yN05jvucS/GH7i3xGnr22NRGzZ4hDKeRXGJRjbZ2WVz49BCjqjJa4EyKChKsdHV
ZEWqDBw+x83xUN6bAjwGlWYA5gf6K8VH8gI7v0iIydEci2UzxMefGWN026hPuDII
B2FSZ2oOxsXh4WwM1rYZetw6u7KbyMVszvuJIdDeEamOW93yTNJnZnjCM0nOhufc
9HauuWAp7Y+T5wgPGtUpik0Mv1HwYljk+ghVDP9qjARPzVuhrK+SdYcDZIYnzEo2
GzEPI3HyxYv0FEnmONRj+GX8J30g2xa9nytQ+IPVagKnskxUItBjRvoF98rES/8f
314lDRGxiv/leEcvTiehJ/2maxikMLz+wP8H7jJ0whPNIw7yQ0UsNWOF0zjAhWEv
yRKwou7Jl6nzF5AlSKNUaYdMOunKieZtjhVFvEdci4DTmj8kXC87mdFomOl0Yhg2
yRcnkhR3+zomGNP2OLdk6qgy51f9VeJuqfovaOkhPc6kCULfXlbdcD7/43UxxUNJ
sO3ipbu4+efK3tBO3sEKLQo8tO4og9yzHRCSaHJKIKe2ZOI2cM9uF34/1Jb8VG/G
ZchS+DGgryC16/T0PUUmwcD1ByGlCo3bX1RM6voT3gcbthG2QrNrAFkSOBMvPXKZ
8GpMwbz8xd3YWTk9zzO0DC22x9ZHmFZ59BTs7jXJto5Jjqs6Z3rt96TCi/D/fgvi
Gu7uDB89t3aPZUBleTGPRHzcrBpk9Sg+2XlQkCk+OcgimEfTFlUarHYLbLbJGkNx
FoQcFydSywxOHoLnwsoNJ5AHPugKvdYY9HnzFXZyHjgEzoBti47BaxnogXREom36
IQvPaBuZ0uzeK5M+Ibn27e9pFoqBEH1rd8FWzxtWYeRN95GV7DAdOJ/WmcjsfBXx
PpG28xOw8PWGoesOcSbcXZ/jWKI//TgKoAnt/inzQxs9HWtRoIUOTwFB7eUuvpuW
Iv9nTjWGYab+EUNgRcNvhhCsZH7PCzMunyqV8yOzphgkao1bzSieCwcVsaOGDYt3
k6MzL5g/6sxsUnNun/TWlrTASoz1aQ+R/0ExyjKHp7Tu2rkc44+OiNKYzZVrY+TR
776vIsqtQryCnkqsJOYvPci5JtglNz0ZsmzQp4qCFsuHZUJ//wVgK0dZyQEf4Kur
g42nyP8SvsZGaqhDw/i7P2nD1D3pLMHqpQ4OHqNGTzee9FyiJDY/IDI/WO5YMsWo
SLBYewi7A/GnyVmwWuIRbvtdaQ9EnA7bN33r4ogAjrgsjZ5t7T6UkxxC/3+9GSHz
d5GQEzszQw0M3S8RySPsiRy55DTNoOeFaHspItU4lbErGpO079lzPJklwBD4oIAA
QprRjJAeuK6WWrg2+tPh9gc8U05iiTiMhwHpL8NLZ8kW7512kYR/lS3DlXLPYs1q
qYZoK3wuCtxbM0qJatZjuLh3q/pJso6R3NE4Ifugp96EMT7jg2C3w4skKHonDgRA
uPhLpFug6c43D3y/N4xqevICWk0gDIQHi49iWPbTVNMf5AG1lRcsYWIT3e1X6Ugl
05XrRFSUdLW33eFn4a1crPyOCpMXYf+PsBqudtd9J3KCflUK6QM9bWbcd84qU9K1
COOtUlvIa8ZOipA+0NAa9tC3FIHRnStYGzCcM4O9WM0nuWdwXeBDTtqjnSETwzaY
qLcT5CGnFT0+8GhyIOUG5d1amqb1xjoWsSZrHxXHw4coZ6KdQLyWAAJVi5sC114D
HbW1ThcOtqEk6DAMoUqxsTYb/EsaW+w7g6XRjHtKdfkp7VlazY/voRoIWjI5oq34
xttHARIXWMzskWHaxWHw0W9hbxZHBgAQyUtaAevkD82FiLjhZrTVbW1FNOuZNwQH
sGSrPPXXL25ocJnRwBMxnkBBE2Ez1PWeL/TTIlWDSupSDtHU1MWO4kKs5zD4Rq0b
Q9P1FvIKlUcFo9GU28pDQ8/9uYkkrU71lHsaqeahT/CLuxSesqDfmJj6mj5ZJpCZ
aMcThgBBvXWRnm2bF+V/x9s5KmdFkmJcwnCech9FMTzm5BCpwVH55AfwzI2dFoi4
3qdiQjnoWQUkEszfBRFJv/kJfv3JagD3QxGL8uXQG+vCQLiHYpQFl6L5acy/VfwH
w3iVUsKchSVnzMLj0xf9FZqtgO2nBVOQo01u6KGlpYReBP/MLbZHNkZMy5C2S/x9
eolmNBBNBBuhn5bImCx97nBAYLp3OiZpCc5+mQzCGL0+cpJHKn8f9dMOrABh4VgM
oQqX4sl2GE4TLE6gI+nqe/hb2rGU+v3euHEaYMyx04RiXu3X4Uh4DQ4DMgmoGo7h
WldVyRiBYK5Ws4XiaJ0pdMEfiplkx4+iEmGJfGqW7tM9obLebxS1jdSQiNctLpVH
ILnorpGKE8B9y9Q1DVJ/MHhIWOGYeIoH15tkqr5VUooTD7l8LaIGiIfLNNoYh2hE
s2Fcfjae/EIfjKCc/hmmhwO2QkolcWpVU0aYm1C+yH+e1aUOffLDTcTujHgbS4xi
xuA+JJQJ303+t+bzt9BwJa6NN16eCd6+wZa9a0XmNGwDhIGZB8CvdmfCPCfFbcJZ
FwWK0ZlGpn0jAbJPJXIVx2YEgvWB5z8RX5H1FvhFU6z/gFr3s0gL3HlywAVGyGx/
+Nuw0ZGjL3L9DzSZDLgwy3ZUheNrzKsUDczECRPxpZVyBBN2NCtwdUFQgWzWUpAi
lmHpu06uVf/BZxXLrgMYo8iQmregbchGIPcPiH7fUpheJ1YEa1n0zGBVc5bMxnQY
IYjZ2LD74yYHmUO1nuDTUPyzAlThKBxgQ/LcH90l9Gb8LBbs7WzRlWb5ay2hB85d
1Gr3NQS41hDh15iUKSBRCBa8xPKRdA2baJIKwRE4YD74OY5KgadX995tu6T/Nhnp
pqRImxyy+d1JRacOGOhjGbRhT82q5lC1Lf0HMb5wAzGoWMH5P5Md7Ov36eZZhWBQ
+Futf6GLADpQVyn6HuQRHfyI68jp2yPH80nJ9Yb6Dlan2vwhBjq0q9RzmxiXFX14
9vbkJNol8WqsFXfjzqYfvr/ice0ra4bef208kfy1YlWNtxGdwnsZqcUO2QnJDMIz
0TZA2HqsNgMI/M9I13JOZMJolkE19q3sM5Ar7auaejxK2rzwobQDXcB6Mp9o9zGj
AS0eon+RQ4rARDMLey1BfsnnZ1VuxdE0c6uqyezS3njKflkQ0ZFPJN6dcDJJhtcE
lmNymf4Ekq6gpW5vKWnF9dNyF95LF8AclZiaeTtpfH/9zplucjzhEghPWjUz8Mcs
0rW6R1o82iEnOuVT4mMjD9zWVEg06mVM1MA9zpmYcruCbenu8j0A2wqpGt6nrK8I
X4gUofAbqSRA/niCoI2cKJ7GgslCwjwk11NaiV+yd9uQ4XN4drKLu314zzJ8oyIh
Ck/lVKStw7d3uOxnfHY/hIVTw409c2dis9PorzIbLK6x4+DPEsMhfKY1heoH34UT
vx0xSv7VfjNtaEjJ37D7OR84hENXxFAe8J2SAjfAjsN0ckwMK4liOKAzj2gMGjVz
XbVuB0/vrex9mJ1VSCpvEn3nkL7/abOQ+NJIU836TVSzyP0qI/hLZBPp1uBRJ5dk
HkcDr8zV0/c3LhddGcx3p6ZWE8zu5ib8UVT8sMBNMfx0Ixg2cSk9AffHNxVCsSYP
hiOQUzO11kZPTCTkrbvtjTiqYRqhfzaEXGO5zE0euFHeywPZqryGNfrugXjipRe0
HlLb2YAqcBqBjt+yGkj6VRakekDnRfGAzK/2In5OVf6vjrLDCpbDAJxeXXEdaihp
Y669FRrPP4V73ifLu/xKouOJ9diNLnr4Ol/1yly2ppx9PVjrDCifLf4I3Ys/Z4sB
wPnwgaqnxk8ZGrmfKJy8yKZlVvOCv0euFXRFuv0OFZFQoybXgobZxz7wVO787v5+
s97BPlAlci8BxvZUn4G4HaYp+aRloMYierWiKhooAWrujJXIhpUCFoO9uAMU3ObO
BtvdtaHg/fBoljJzMCsZu4s5NG0yhMEByu1+25kxxqWOi3HdnzkWfaecaYaekCMH
vFp8BlG+Gcu5DoJYTDFQErJJEnZOERPTPs3SPJBHRrM4Cyc0+5ADmWp5D5RnMsuN
EjC8rRiVVUMRTLgmjH4L7Hz0LipmTWS6AnfJ0TQFAVch6efvjT5sWnQ54zYcCFoH
CwCKFRrzDWFjWoIfLk29hZ7WzKzL6w/KLwKoG2L48l5Nqv225Oe9+GwIuhlTqub/
cKx6ox75ug3Qy5QdM1vFz7NKG/pS2bt1p+MRdVzOUozZNs9R5QiNql471un/M0vD
Svt+eUi8BBPIFd/0IQJGGHYIqZGTxgwggJ+BR2GI281D/TTvZXLJAC3YjE0dVYOy
wMSSjf/cifpK0d9cVCc0AMQDL2oNoAmfHi8NYuhljU8Vo/Hnp4NLaBGfU5x4vIIC
KEEU2/Q5sLHEF/vaWF7t9XhF5jtoKFDswsbuR0ui7ZE/vlxMMnAcIqkSt2Uvl4GC
DyZ+ObCi2Yn2Xv/SzbYCo+W5N1Ij+LQebSkMjvx7uFK9b/cXoR0LTmgV+h9KXkUp
rgCR3I1FNu05O3cl+g0GIsQDcrzTvkyACfi5/ew5fRxE7VuNB+iLVckVRk+WfWQK
vB7jMGLsXWiCRqxDqZ+D2CjScMkKPVG2houBQX33+ByLr68MaJBBrWAsR5hsOGNv
IqZRWUYqXOjVMBjfcIzGtbDjUrDMo4gk3gCFtFMTsHxlbea63QUSuO7osvSDMb4P
JP8skFASyC93+7ixSnWzijnWGL3VQEt8eHmKM2Tuo71rO5dTJ0wUKYzuWCaII8Cc
H6HVWRCO8B5zAvScaEzozDFCo1EHCVjY8aQl1QghluVcburFwH/V7pkdIVmKsuM7
iNZztymtfUJdEPDIkZpwUTbE7o0KW/X3lcYD1XdE1n69SW5MX0tf/C/7gII8FrFu
+0VRaZ8LUM8kAZADfOJtZoRcFv8R1dDavJiHzOhXgLrCupRFPilIiTQkjNYB96Sk
HiusbZI06m2F0OUl3tUaTSexcyTJa+Lt1sKaLGArg5spgK96dG9B/9mSXEXdM05R
2gdaztV4atno1ldoyZkqe3XBzLrZLmnBGdpY4FY9qSCYUny+2JBEBbdAtxCmkqyU
KNSv/k2+fO7hUjndieLKXwPCtintnyZdhm9v25qMq9fOcuaR7mqlDf/v4jp0Z+Az
HYgIoezTGck+gAXoZeCVKk9m2pJoaj9uciCQ8uGmzyx5Ff/ixFNPiw/fjhi6wm4V
IULw66oRLFV5nIoFYBG9fTjWd73Npp3UKCOB18dA5dqh05iiOWlHYf97aseeZsMq
eUSomjTy6ytr6aQ7tnG3Y8nMx0uNvDlKMkj3RWlngCZg8wqVK4Xk8jPFSvFzRcBo
gPTORV2xclTJePX7Iqd6PVger7L7PW267gWQCyPKXPwxBtFzKCvp/H1GmpXvyDKC
GY3ndbORKp1BCMl6aOdDuMUq+0tfpxc9NDdgeOO+w96diGiFcX4g9I3RWCCMWKc2
uQ2hvOOpPGyvNNTvablbgW0FP+AFzyVCGEQOCGTkZ/Dr79rlX0cFOEbkjFr495bZ
f1wikYFz0lTKXyZlNY8PkzUIaiTybSzfICG72BRjl7sY8hVw4dwB0ZBDu2DxSudV
Hs+ICopDECmVEQ74cRvJ50k3+jd+6Cc5METnLVh3TLsAonjMYdoOoK/4xw9UmvA3
UX2PC55WuImOZWUAkh0ogaKTTKoGE2evsRQoUMWmICK1x+BdTOP540SAg4PpM0jy
ITTVwSmfRNe2wVPlFbb9ATl1FaK5uWLC8nAEpVeFk8qsipcrCjcILTj5eE+ldKhV
yP0fOv9GRa6RJHtGIYwhNEw7A63l91xOF87XHtld+mMcIC5g9Stf2GBLkXxbJNI8
8v3jN34f73+9isUqzGrzVf4bto83AvnIZLFYmxlKERcT+gd3qqnhd816qy11ukb5
UZrwdoz20dAmnW6RGuaZ2fMmGxZWGsPH7+RWd2iZeeAQQfNjwODY4klCwJ4cCu2d
bj1jxb8kZXoZ2+p+mnbrcXJMXG4BhO3Trb6/Zt0GCrkMPd4/LMTDm/bYOweAijNV
564Tbx/HT5wm9PYwuQt/UEdwSqLDZzN+LVGi21Kcp1BA5wGwFqUSqG63tVi3ePHe
lggFZWN/XKbx3mifBOH0+Cqoh0ks9i6rdpteBbC4PrNIizA9eaax6EFu63Sz0zwr
pQKVRU2+cBTt7tn8U/VUUG/eHnXtmlHfRD2gjghV3P2/rw4TooGbbsAD/AlfgHc7
Q1RIpQrJtWlqG32G7T4dxEjt6yv8gOTbyS4Zs+vM6jcoUi1Xt5ebmOa/rHRK0xED
GtVQU341uh92l4Q7cDeHxVgzcS66L1d6550UwZsBeLmoe40lAiZJ9lU492umtW7O
FZQbeImKcB9i9Jwb6xDgH1MoEarCal3rtEoKZVg6MMPqhP2nWpJz/CLT7MKB0Hzs
E0Ps4ter1y4ZchiaUdYE7CXqPE20RLwQDWsYvzu+JzFO6t0rKYropnsd3/F0kjcJ
PSyojSHM52+pBtrOwDvemOWrUzmUKu8yCt7vWCYt5JNcQ2GK22ytgJRvK+N4oMXu
G8H2DyGM66bfF/WM/+192w8ovJzrDKnphQeVqy4vwIUvUQJVJ0Xx/DyEYsWx7Lct
mwXbVicsIzZeSs5si2y9ZQmHRn0PYKl5ba91y5l7KgRcz23ITXq1BCbGq88JBILN
EoO1rVPtsAHad04NPEAoH4Yc4mGbfHYBNz1qsgqUxEoXJsJODMp9qZeV/1CpTlKy
2KL+RFXX/8Bnm+euS+bn4B6Z0FwqgsLMiPTL0DYMLg6eRCE8sJqno/Yvq83pV+sw
rdZ2G8FjIRQRpO4trg3r9wK1RaOkMHySrPePW53vbQO45UPc5zOj22P3DfeNWf59
4XZFYjKdI24MGrEtqVj4wfJ/S/2wyBxCNSgwXPzFHz0c+0ab7jbBIK/ZBZ8NyNYo
+13f4409HWWopadXRUn726uAGVINQu472i35dcvUG9e1kFcLj8B+PD4b9Xu6YKRP
1Vq4U00luTeOVIUI2vHUujPbUhdg7WOJwik9JkaAB9AofrFsfoPZejF2dS8h8w3f
5lgXqxG5ZjH0n2xux43U94n06NE4x6N0MJWUk9sIIvOmY5wWyNCAppFxhP9YTat2
rPBE+Nn/2xZU99oyOS2TQ8K0fFCChrHqlSsM/NIORQN/UzKh1z0vvHh5nZp3BOVJ
xHN3+JSlARQVkTX/etDtgSmAk5g0FNAy3zdKexni3aRi/CZKAeiTFLpWw0q9hHTm
GK5gV4TnG+Y2JpKbwiffdlVNBnDrfgUfshu6hdhLL18otIoh1yJ3tSO8jvgX+Rj9
FfV/eCP+EwwCXswBvsYIbJIBDdZvaMBJQ7lzpydnpA9NnzyWFw6NZPQ9aXUY/4nV
E/EZftrWuvQW6d5QjzuhzcheUOM/0as0IaxQMfClAz2p2aX8NJVHPprxvxJEM7Ca
JpzxfRtXV+jiPtyBryQdVFNbk3WibqQv7tlx4x4Zc3XS79yLGdK+X3+rbuxyPVKt
57MT+eS97tjeyR0EUyR6hIjXRI5Xzy4w714SNqg8ZHDLg8DnT1Oi1oOCjXi8MLFR
pKd9icmGjEnSMLaumTsn3SW5fQ0Z2Gr2mEiq1qrj7aLHY+OiIOrJAbBcVtYFph2t
+ugVaFgIKfEr8TwknWEY7HHid21q565GDJCcGHpUnZv2/xKSKG5bYUSmGos9u79V
7jKaF/PPrq2Xq8spPL2S0zE1dRV/dVBo/89wzEFQei2fetGV/mn51KYV0KoBh6rW
uxAdPbVHM1NxeB2Bs4SbXEo1rqpglm98ZHNWKuIYZwydigk9ab0GN+MjFUZKOCn2
kEEZvSO2fLMQaKcAgTe841/n+78KYL922DFxgGsdcC4JD4Wdwlln/vrSk1VoS+ii
qUtxt0bouiIw1nrpL75LWLI2MX/3BcjgdYso0RcFZNMKqxmoeQmX95nddtM450zk
192+/YdCXr3qeQF7I0h/3uK3AOoJ7I9l/plxx2KBuVPnew8FJOFNiNKTqc8SBXDK
RERtsQL83SUECNgpuuUg/PegBESxXXQliG8kISYQDOfOkT9ATJGQFneJl5hz38CD
HyyyT8I6mk9GF6fPrtcmzWtSA6nzqnUxFDeazFgMA51jpf5B/PpX+tQEOA272gTJ
PyQVkAK2/4UIVX0XZrKj/CSZmRFdnC76FKq1Qy9uP9sieK+7dHR7OOvDm0dJwqlJ
B4ntKJZBSK1o6V6Vmx4rsxGANlMNtmJsOEWs7rzrapp2mZsxyV2O/rf9iQeCRjCW
yQuoNhZvh/bHxVu/96K2u7WCl+BR8ducyJWVVvylGgK8wn/qte+vy5i8SqwW3xWY
kZmw7ogZUWORCrn1n0ioiXj6RpxHo83w6tmbsh354+01vYsu84juCy8d7hm1daJC
myzQ0U3fycHvxYpEbg0bGfmgKZdVhzOU8F4yFuqCEOoiiPNNaXugOWbOzngB3/s7
Dn3BDSyvKP8FT5mgWkAOQxKRkRVuYFt4036emaVo2n3HFLJeku/zxf/q2fzoVOo/
6Qhz9qyVEYf1v+ECf9YYcNYJDuQwZiT7JNHchhKj2SfBnI+1m/NAtLGhJu8RHvHe
8OFTMiXmOh3vDF053V3fuJEYP29aAOWn+nU0ZC+P9gRyJlaXtNK8BC2+qOAUHDtn
/3e6KsouCcjkQOFDX1o0HSB0X0d6T4VsWvHTnO+ikjtFxCesZt/eDy6bWP3bqWoW
1ttNYR60Ve9JG3ItzJQZB99PeSl5iAhnFkp9uIoQlU7jSurzaKZujNPyOPWp/00U
03zMWm1tvxOIt0YeX36zsCcC6m3B4IwuyhSfcKxkg/1atdp6VCBXyfA+ons914z5
YsQsWfYenaZhyTUM/ZsuLC1osWRfLOD8qpE52+krndeUZOXB0bNczuzMDHivJtXE
BXy+jWtLU+aTk9Q8yRVea2t3DEAUv9es2ysH0z3+q0PvStPeLsev7DHVi+o48vQx
UgJxgDtVZeVshykqMGORFVG1XD1IiKCMPhK3leqQAFMkQ1I2YPSHckgB818UbACk
GMcmKNI4/k0N70cnYAi2PAyzVIuevkKGaGRAJ66JyuAk6ZmHyzXNub2EGAnMXdxr
JNWHt79TTH+1H4/FGzkUA/jED/oXtKN4iqtopzZpxq5xdt8ah/KsmfKQe2AJ20ee
1OC/Mxbl91SGDf+YLBEPausFD9+sxdfkpKG6VbY9ndsiKJejlpYR5UpjNomwaX3o
VTo4/vkOrDSrrB2J5ldoeL4rqnN/ssoUQFOUhqSjJwLhrZWlwe7gSPhjxMRxUd+1
L8/1O7SZTOEjnT+DL1yT7Qp/EN/ogdl5CJOzvyLYzEK1FHn9tC1bP5cAZEdZ8MQl
Ibl3jhdDNYgkCc1SjzQam6/hhE/qE1gQmFW/BUPO2WvZ89yvcCpTVhy6jOUth0zK
LI9srjxTBvZeBTHC5YJMbGQJvitRvHl870H9K8fx9S850nkCf1TWGY6HNaX043JO
rM1mxqFJDxcZF9PhMU2UzgRQMx9He+Bbr/VQ1S9JvHx54VyFIdRad8TXNoPdJUTX
Llh/OgbK/L4Rc6xQoHTUqf+YcPwKGZWSZ+tYbySlf0RuYWrlW5jCGJ6rWrzyfplz
6Q7H5pnxmTuDbVglMlxrBFfE0V93DK8yuDYKfZxOdTdXdHzksaJ/EtRX2Uk5Bwpl
YAQqf1obc3sa73ilyXaiH6L1fpszbGzoU+j6DfFSKPiqQZ1p2DfzugW6NCP4BGCR
Mq8Vtuk0bk3sh9hzHD4tuNvaahG1lK0bhMWihH/gf5phEbzqBk+XACo7i/W6iWtN
HRWFUVA7iUnsdduw5jfLIrAM1OQLamlCCfXD28XrUoc+p9rL5KqUH9rJBotU98+h
MOYz7HDP1q0cpkoI7qmB3OWP4zoBl5/81hcCkpXZzqlhcClZJHeXD03gHMwtcMAZ
DSDlDlzq2R/HQOWFRcHY8+HcfI+sxX1cCyXf5KA91p/Df3mfek823tz2iVzhXqLv
UIE9e5AQrHIJzza55H+AF+kc6tae80AruqfyeOiBQky6poOEifqJzD/pe7Ugsuvf
TSny10JZrSJPR7MtWAPrB9xBciB9oRfK5mzzQ1JOdH9VYu51oNR2Ydt3SCrFBS62
xXTtUACBlXL8FB0OhMshHdD06Lnj9x/UiJvD0VHvkCefU8CLs0EXqRDFxdCGWR3m
U7xLX2TPJRmP5dAmfYkejT8jNXL4pYidlODmX21pQSj8GZ6ahUdTKteZrhdOrZcU
VJHrl1UuOsTWIOZr7EPk+OS5SzYqf3XMDQKbGFbcIYeRcwNrX3hx8m06lGnkmn9k
xkKPiYOuAe61FW4dC62HYNGD+3PDYxRhN5IpJaXL6+F2Pti+GK+Yw7q7uKyLMkYn
PK2Y/oQLV3/SUXmIldOOPfoj/BrhtGdtYFGXWVKRe5zPMYG4SRXf4U1P9hSjEQ/l
+dccUNw6BOQSXIjA/FJY++hHxSuOaNpAS71rltt2zlbFW+uXtLpN4pMCsOuucVes
8Ce9/dS+GmD1r0dzMoXQx4opIHczzhC7mdgsNzAsvTq4m18hpzG43z9m2wcTbKUR
ovb6+vzghBMxbhFSqHZEGP8wlEJwlha6DpPtyin/oWKnoXU6R0XrJYfSdelrB9Bk
MoS+s++Z+QJ06cRvxg7O7lQ9EjRgxVgIYDO8FqIyQszv07BD03yWst0NIfbb3aej
Vr/oBjt+RSTU9AIDcocHs6dSKeBQIsaUeV8ZKVYvUqOtRud/lA2xxQZ8tedP96yT
CNUmOoFKecxxDxzCC5fAnHhsZ0zH/ZQQYNKP4JM4hVfST5fvwMn/e433Q5z6lFGd
Ete5r5bIvMsnU3/CTvTS9x1BRtzAPtr4/p/j/8vT5fnCtFNhUBZRdiTbrPMQdzEC
YQyZd/dD/9F7dMiJABSjM7FO4MaKuuF7Q5ewACifsroy4qqNiUCZZqblPGJd+REd
KKlBb7/7FrnRk/60LDKMXrqZ1A75eP3qOCBx37mdKr8qNIeC9ACAmmdgbaalVyz1
drdzI9a10BWU29VO6lqi4BunBwxjeiV9a40kmaI9nLQgxkdrq+oitkvSlc1B5QDX
X4Z8nUHlVRTPUal/5ibXLE5KMICph0FbxT8lhiJdpTsnpA+QiLBX4unLTyExdnxK
CX51ufx7D0K2/Wi5juTsqK507/WSpz/7bCFJJsjaj20ezvborRH7n2SiLPQemHgE
xD9rz/G3n6DG6MRCLs1FhkPGerUZiF0fvcrnTLZhtMHkbHBwNMhxf5pb4kj84CE7
oeq/XYDgMJ0OxKaQH3dqYD4KYPONPGHx2Gm9qYWRmNfQ1ac1tf5mCaQf1R3H0A3B
y5WvEENP0KnVdCl1B4yUNTYeCfc2euvwalMTrIEyDgoikTnkB9Yo+LzoC41NGaNJ
FJ55rAMiyAAKZeTXhInMQ7UizAPm/qryD7ENnMT6fffGKxliPs7sbnIWCi4hBIX+
AJy1q6SyPFLugXeykHx6g+HzVqx2pCy4EWoiiGEi7aA0Ocdug7V0ZNyau58UGQbd
jfTN7jcW5MjKuSZXNs32Kqk2xy0K558xqGkQPiTmWlLIDz1HVu41htWhv6Lzscl9
hR34igaOy0SH7pnGmv+fre/r65LPM69Ymg02Ie3SXlCBPxeOoYNv8qt75Xt5ExOQ
5k8AYQvXfL0J6QFFEMDAuV89P/M3o/ZUYFkrXWmg6iKQGf7JMkcD+pDqQhZpSs38
QnVVEsabACD6zQkois+fm2vde9xasvD8E8Ro7fNzlUO3Y49yY2lVE9cubeZi+U2h
rEB+NoABHmRSTQx0XwoebOglOMEzBqaPc6lqTgD+tygNQFl7gDgNF2qXY1LnmemO
fKMFpW9EoXDaQMmgK94kK8gHvTvcCAzz+PCrX7uzUEM3/Y2rgZMewP+736N8ObAd
XXXMpJfpR7Fy5xT3wSzEnL81vi8rbF7uPjR5qHZO/IeFbu7ExRdlouA+RjibKLiu
JHNh7ANjdX7aDP89FFzlApMMkSriwohEQ5N++l0a+T2o45ShWh6ptW6fQ2HGk8Mg
SVmadrDaUCPdBxVkzJDWZX1xoMOa2hKDovcVOIkSN+RuY/RqXHm6tWHqbinG5jIX
TifUkzaUmJKx6Zr+zIK89wMfCngRmhuqfjoYSOSPt14RGe8dRZABOflpIsqLpj5H
oWqXURDu6+qQbv4vHVXWQeH/B6LtOtBSZhBNiL90eP5vqlIq84Q4HJSgDVumRzZS
NyqkDnQdAYCP/zb6CkswVaRHXSHroVWJoc4/8nbL4Y32Gc/dUX7NU9CfF3+JlAU+
lQM7A9paYt2tB0VBuowIT244d+eVTzI3pwIlzSyqpMc44RDKw5Ym/DyTQ/ThU/Te
bz7ofbKSZDn9Nw5uv64dDWj0oYM4kSIZQ8Q/l7ncpKcomNpprIv2Ibn2vjEfxSDR
PewYwe5Ol9i4qO1htEQIWIBY5SzQreMASjziPCn+lmdl2PxJvfe+D0GVwKcK7lZX
JhzbEwLPh7LwMdaapOywQqlUD17e8yzfdRJpREUlk76Ed3SJdu/JYSvbCh0NxeBw
40MIHMrmeWLCsI2d+U20byzaMWI94h/FYW+Nso7o+2yQpKtHO0PMCQ5ZrydYdp3R
HeM3bFjHuFizt15Ac7zsw4HDuOKuOSkrU6MkS8ytuih9zWVHHZYt2dCatNmmEMJw
4gRcFnaWUbUKu2uiiZ6rGK+XPmsBv8pj5MB5lHahIjrHFpcMLkMFmGlgIUtkEGQx
JJrB2dAC0M24YdQJxgmSxmspjK+NnZLtoLryR5trPp6ASJcSiw2XJQG2GhAfE1ge
s0pGc1OIT1x80tuwM211drs3h2rgpIFZWizHUUzPyDG0HN5VJxEot6GGC7jrqKch
ZyvlFhqc4+L3kV6PrRFlO/fNPs/np3yHs1qxrrT580XG4bos1D5LHvALPtwNZw5j
fHTjslFW0LMlKFLkqdNJJUsrY6YbV8zhW2fy+STj84KVs2h0zwmVkJADqKghfCqD
pKfe8+Ske40SPIG2H8YIHePgxjIcDge8Dk50ZS+Huk+MO01oWW/gVazabyTwMRGH
MuIBEi/YS+57Z5AyIWK0SfcAiOF/7EHe1it1INGa5PYHvHkaWc1Dn22Up/zdW3Wk
GV0Wo1mdr7HjsUKbrYxtb5o7bbPbqwGs2Lu7qujKWYHgRr+VNhF00QZGErE/1utb
65rFDND65g07JcKjY6X6rNOo54+6kgCRbVJujHkk7gvozxogbPyGCoZE41AMb0BB
htCK9j13j32Hb1la5kCpDov+QuiC2dvm2Y1QNS1Hkv5WYXMe7aQ7m0qozYWmq49f
xktj74KEDNzqAwVeKPdCnW/pgFQiSneYq5Z2pDCOLpFAEE4H0ansVErDsew1OwS4
luEN5f1FG8VZsgC3BaqSrcB3mLCaJ70cCOolKvfD1R/3HsR02f8Tzp1t13GUzWFM
n9y0J44tN5ZvvKS3PdkwhfXrClWg5IUmwUF60LNG6/U0olxiMv+LkR3+VVWtaBVt
8Sq+LjAri8Cit7gNAseTnNkpA+cGiwHBrGTnStr9RIw0epwcm91MCWPxo43a3t/4
5FhUJz30IwaepoTACCj0/f2d+sCofnX1OcT+dNlJ2/9yA0dKTdergNIPzgaY/Eu5
v+qu/1CoWrJBpI34mKsBfDi0FRygvwV92kkaeQzbfiXBuOdKSXpul408iBGhzCgz
TkFsmbd7wRXZAJMlYoHQpq1/kp09/gFagDXJvbA+NVKbseSHFDwNGmskxRV5pNl3
VROGQB2aK9XLTO+Uxr1unM+WyZLXMWvnOkmzVDsD0Nqw4jDUzRPHddhy5e8Fg8+b
dJRH4CYTxH44Gg6GQs5HKsb4Usrglp/AIQDskJnc9N6MdBRndrlmGpuJQW1sxm+l
z7Jc+OJ+AohA5nmqFhsnlcJH1TtNpEnlNPrZLQs+tBb5SH427Rxj12BtrLWndqL0
z9R54XdL+o7S7EqTES+SfJmIamf/03Zq5zNeXW9JARPdLgc3LOxN4SVR6pHcB8Nl
DUnZO8cUWiZpPvRERk1LYZ40uuNPTPc+KRkyQOuVy3a9RCC10UHzUlJitc2sYT12
YSiY2AScaRPKBAltPXfC3hUOLkwtTk12iu1JuTTqMl5SS30wlMCyLeTYA5C2T5S+
FGZOHcWy7iOJamnUOZQDPq5AeYAEUG2vZBy6t45GzOr/gGNUOe+aXwLqfECv4KVb
jWrnyMU2BCaWiDvo0Wg9jyvsfuRsKCIlKTQPtLK8vSlea5USheTEERnLSJ79HECR
bhbMMBBv7c40G1MaUL8BA0DDUnUTg7OgX9OiBxChmtskbEh/n05w6xE43SNXl/D7
HU7M+4vcZmqmyP6AdHebBcp+FLD1erS0YO8cDhHU9l2FqCSgtKe5hXqIJZkvMw7k
Trymr2VlvRBNUu7VdCogaTwqTs/P6623f1+Doe2TdEefQ11+Tj5DOT/j1/Edmlt5
Set+k5Czw0tyxSR4rctPXiCln9PxQ9lMOyDBKrCMS+5QPNp4V6AvBLfwNCtEhQei
IrsfhIuDXsLe3PTS/tfiix1oL46NhjFpoO6/efKRgtTQ1HF+4VF+O/yeIHXDf8MR
WDSOxA2mMUishmEjuDuH5wrgP9XMEHmJO1DVgt65rVRWXWQ9LqNIpgndxmLJ4HnY
AVsfoLKs0VBcjYI6P/kK3B7F0/iEjgaCRg6NMKODtrguZAv6Z/AXR6hRnvO6SrqY
n7goP4VpSJR6ZRtRkh/h0mdZbyHlrruuZUcnDJN50exK7jxy26ms9TQbADvMuTty
klp5/hWVIWID/xE5cU9ic2j+3wUmG/2I6JeIT/Moir+tmVgiBuK8+WVw7WnEHyfc
fBBX+5Q3Rmqud4A2BRoYLA5/zRX+ArPTitChDcKD6BsQWd+xsOh8FBEFRc2FDN/5
8c2bTYOdgX8mjEYP+8iTJITLis5IeD/WZ8wAsiUQwx6aNF0/HC6DVtN6geuohADV
S8mvPVHDvE4E8iLvLQ5+fC5srF67d6u6OPBO0MA7WlZSd4w5td3Y+c06JutTiSDX
OpwGSadRv2wjGkoXZpwoDk6pKbs/jggXbC5X3bnQHU70A8JQEN7LRWZ3i8yHDg+m
klnyubkeh3ZIUZGm2OFbEGZMoKgFHDmhlywIrh6dJ/anLMO5iGNNTOe9BA8ibgQw
6ptpVvFgY3sqgefxPvfC1T1ZZXadY66pZsd69zMqipoI8mONRQbi9TarK6aDnwuK
Ljms+3uJbDzBVbNikwYUCC/CVvu3jG26kPYGqyW2KDJwbsJ7pL2dwZ+FEj37Pumk
uDRwlc+2PChQ+ezlM9owiw5Y/SoPFI+gOn30sUuq78RNrETRQDQRUrI8jd6JHzhf
HMWjRSFK2aLcDltgF9N1RyZFZ/jOOKUVOPPe5j/mLR4QCyq0JsVDEfToZqC5ziIX
0VbPt/4F1+IeDBPADDirmQLJ+P8ZKeIKAYgIZH6BxZAe8QUE5B9nXF2fduoxzRxR
hYJ27Yq23/xT6f2jwA4FrayZelLTD595S9vKMDJm6XuruTo6YkfixFaIeMSGXEX7
QF23XuKFqQu/WYfW1Qc7G1AHA7VarBa/qn2ePeuxvskSOGYnwRrBFpy7dCkxB0L9
VZAAKJ/lKcHNN3pCHWSw21to5J1JztSzl0cM1AkJO3STPYmY9K8b22gykK5G8NT7
WlF0bDIsijge7ZpYmCBFvSGtfWxAZ+2Kdsi3AHyhUisBCdnQTYNWW1NQg6I7glF/
VLCxixRAT5bZ+HnZEUbyZDZJ3qNmg4j7XQ87i5UizgQQkplLLTFx6VWqrqFDfDG5
idEgHiafS061FtZF6QLGRD7Tho84r2As6E574qseiYRrlElMv+I8FLXXVYf/z70i
XVmCbmuayJ3vKfqFKJ/py0Zodx3fq90P/upZUKIlNIjb4j7u4dPzl/1J1OD3v5qo
fs93Lr9INyH0/atSw/cYy7m3S4O60yJ0Je6l/iKK/a0OE+lxN1iYJYXoDkBtoMcW
hTa3QCMbtc9zZdo1V/UzVmZrBPbRbAxhR/hE6RPJIeGjsV7FKZY3ieWyy1OlCU7J
mNwdEWHojZRau1P2K0HUUDiqA3ENVkvCx5t+AmmPqEkuS8AesKGEOFc5Psi3rPRi
uy1MZ6NpbWxsxJ7lfUm2tZL/87I8gk1TwSd/iL9YxNjp8W+nlgOcbWYGugjofJk6
Y0O8joms4cMMYzWjtItM4w203wBOcrWtgDEb4qzNijPhWVZmoEHQJscU20DMPy1o
Mti/eUncY0U1uP/WVp74GpV1ek3OROx2PN08FG5UsBJ0a1dl6RRsl9p+RJoC2rbE
KkPyNhVE9eP01QbkdKmUUp8bMAE8frDEqDcHR8VUDLdk8ByAEZeYQWyOyyoyVuWz
bNtEp2XhXiSeUdALHZWpW1/vb3YXOukB54yu7M7GJdVsQ+zUsxz+puM+u6CQLYVp
YtjNgxpv2VjnPow8hnDJBqFvBq0rL4hSmqErPti68dsWTwTvV1/BoigesLpeGwJ/
aIUaFFO+PQfRV0up4QBnkL/CO2eKLXT9DLNNqPFUzoWVT3NSSHHlzLxvHHhJXolI
+mgDJuQ658yTIpJ52w69twstMPslljkt+ApAPyzgen2mHfuVUiw9Lp0l14DoXWaI
4TgRKebOMk6poOA8bFYFQemqheWRH97OPzvcMAHronXac0d8+GtoiEhsDAVUEcuC
kpr/GR3Ry6Hm3CX4YDwH9sCrgGhkww4xpDSMGlbC+UqUkMwNflQODutM1dfaiRSz
BRqQwp3LsOLD3koQGgPddjetsz3Jfq+vA4UsfDLuI6r2t63Zw+iKoQHpISqoFrGs
nWhQn3R7lc8gucJ6N40gpFjPC/VZWmmKhn1LcCgl5+/TdQBzbj5U4FgoG9Sydt5F
FZepH82VNrYZIkq3tg6AS1MSR/xuRmDAWpiP527EcQQQjvN8d2fKvcl/gumeofCG
P+wVuCxoC1pLHGIZBq4ob3N+gAEYyJ/ORkf2sKGnCpZ6mLDT2VuFRrfvQPT+B//M
WtZpEnngLkB89wIihfmZoVJj1cv6CUY1yAcyMo7/chXWcoedBEFH9pc4z2MrNMoE
KqkUC3Ld9LQ4l7quwjRvbNWdN53sGe8oTQZnbryMcOoLm/xqHe/USC2smIx1Tydf
Afk/WOu8Hb0ufOICwR7ByQrPpTIEQ++rPnItwlc2mlO5r9Z7+KTtY+/dXZm+ah4q
WX/sBN/m3FHimOIfHLKVmIgJYxahFfyeTc7t6OqeQRhY8RjJPDeTbEAWynLDGKud
Hlda1SBkttxgWJAOu/BmrjGjF+8UJbnqRpf5RGcPnPBEBbOKlfgcj5XX7uwXWQ6e
JgWkvqnNZ3sIYxlvQBo59hTCBE+QvJrIs0wjNwMPn8wjLIA8UX9jGq1BRAmHPgba
qEQUAtZgR8227tTmfEScsww4kws0Vn1depj+/8X6OGfpm/+Cjv2poPAFd2p9JHIk
Whue1gZqaCFm0kuRPh5c7ZvVurPZEBbrx9evMY6jzb6CQ2QcuvIs/gup3eUwB6hD
NeQBbFEq51bBNjHO407Ii0DPlRgfYrcqfi2Evy/Ub5D1QQmjNpAGBUBiBbFX2ZCV
HtIaBkni5/Dz1TPE0w/ej6se22/Zh6QeXYEvrI0DcMZHZh7oSzIRYtd3Q+EsP2ti
a23HESiMw5D7de51Yb1ZV3/QSpvupY7eYap3YuPgF0rSpn++s3FsLVkhBugNFR0D
iO3OA3n2PL3u1yj4NuWtqYIC41BYzU3Dn+wwyd1TG1jAIL5iCvc1ps6hfeC84jno
V58B6VU92ps9s3sxptiaiK9lkfcxDw1msYkqX4u+pKMeZ5zem+OIOi9QkSZ6JF42
4Rnt4BKoH78lQG7qAKH4Aadsh5JynQjjfJPn+dLg5RmtNFyb+scktKzxxHboOdJs
QMxmluyWC+dBrNzI5XUBHpyw9/EnMQxD/AYS0nQZ68eS66FSInVyeJcz37Ee12bF
5gM12ndwUM1QVTV7oV7B0EKlftTuRXyCf+GhbDWUP4ki9CND/uKNH8t6EK66uH+9
cNlf9VsvppoITRKgPHzd0qo0stf0qm4CAlh4NISSHMTw0RWZqr9hj2Ev+u5jySl6
SF+9DwVanFllP6WS5dJk+khBSzab+QabMz/TtdL/p/5whghTw3O6COUS7gnPa6Tl
ypra7lWRY0KMsIQR6R6l0QTzUL1GbRMGlvSnNgwSgpxvSsQmioVj2Ec2MEUzH7WT
LbSLtYeAMWtRIBDx+X4CT0RYUWp+7tZ6cjbrLxtufmvBbrgkIMPPK1vYRAhgfr2O
R3QjJrmk2KaYSX/VYusGTRaQ0E/JVJnrXWn56iVaHRs/wZlGsWNK0rxaa1WPPyrC
oYb2/ScS5npWcyr0ClI4Qsn6tM3hVlIKY40WdSVGcs8yn7gs1Xzq31KMBpry4K1m
W+PMjZInItQ28cz4Evwof70LUiDqwzRj6W0IaoKn2bpRqbB9zOIGDUerc2eU1i2Q
xaS/JDOifgA8swYJioMRNEhG6VO7kdJ8D/XvXUJwRBWy1gM6RCMOdb9QAynTGFgY
9qsteW4xyxPc5lxLqNMJDVBRaSEa2nyod5Al4PWvhfmx3+kVaCjpsX61xZ/LVoYm
JRuJrZ/6X7O1+jqexGHreVvi5aizRTaFdXLHqeib443fB+4Kya2VuYrOC0QeYJd/
xphoVCPM+vbOVlbvDV25t8KfWi1/iILR+lA00Daw+NefvbThLUmxPvVn56rhYRDk
mbfOCLUSGPKDuqjbTcGA6WI8qLx0mDCJdmsrnnjFGV1qDwmb8x47gDomQylhGHuL
m5MU+zBiCquJrtIpA0zcoRn68ehDvmJZuyVF0Ht+livaNVtHS1dH84wKqMMcuGCJ
F71Mw2brj8tHZmpRNlnHbMZrpRIRvoqOkJq3oef5MkiW2e0jSUi0xVbSHwR520T6
b6xepKSkiqOFQyAUVs7NEIUcms//BgMMhLJboV1UEbAaEfCO2rKK0gsZgQznJKIf
R23sv0f6XpTRh3C8fbNKKzVq5y0q1uFG0kGKhAlGGVkgfTEdtlW7sLhLE8IFYfEt
CAhMmg2f3MIVZwPInd85uHyMkjbHBO/eGtOafgaiBYuuW9VwWHpaJW+/ldzC3VMz
UR7ms1zq2y5apzhS3BxzNTLWOjpGVW1d9lludW8378oYjnDYrjoUalHV6cvaSg8Q
HrajFE46EzWTBl9QYlk8c97kTzb1P6uCzBlY+ilXQ2vwiLUHcQvRHvDHtHAykkTX
Avo5YJ1ZVcavTJE31DHVFggNuAcRjJIKlug5O0dZ4JD4FrhRfHmV5dfJQ0ERcVqo
vk/Y7funPGFKz/2q0htMJA8P1uN2KZkSola9fBS7+syVm33w0d/s5Wsq8yampnNW
KaDQgLQzYJBcphhoBaYcInzU9RZfulWnFGM6iIwSY6Gz38FZ90SYAwMfGM17MwqY
TIWrZcfpxqlMnbQ4nv+mjdGczL0cUI90hiAvUIj8MDjRzJ6gbQe3wZkuvoFNlHMB
Gefa3Da+fZFXLGV+75W5HRA6ynGEQU5LtXnq+HfoQee9xNIxkeIViqHulFXAvpK7
NtipfxuKjQGvfHXM6lvtVcaMnsaYpVHdr4hklrHnzgWnpXPGOrL9BOfG102qe8Cy
33c1hJriGAPa87HZ7D0U6lBmH9PVnnaO0UlTsjoLfZXSr3e1nrccUHowFfRXeXIV
j7TBg6UKUpN+5oEJn2LC+Lkf4LLhrgWI6/hUc45pQmUcQ8EcSTv86I0FMBWe9tLs
NNyNGvzHE+C4oI678GrZkGmY2NB8wRIqWw/GH8K8MksTUEJPCpmnVn2Nr4o1dOt/
o3um4phNHkfMBEAw1PZao12CbOIfsDcis1atSt5Xsouexg4sIlh3sDio7yjHBG9g
8pjU8TVJg0hBNdbClRbTtZ7znEN6Lc7xrMnG91oTelFUcIHmxRSnMnoe1oJznWM4
+nqZ4T+UxWdh2rIpaOMuYwjRqrCKPTpn/jFOePQ4n0qiCT9uWzixOaBibV62NE2H
LmfioMDMQUU5FRQEp+4QToBMSNwb6+9dlEkZVVmlGtAWcbWKE6i4I3Odm4PYxkTU
zkI+UZXh1jmUftxnGCXtAvZBMZqoczZl/L5MNFO1cwbinZMiW03G36xNxUI5SpsX
SbOi23aO6VEvJPu0ishkbgV1VjJXwYsrq0BCzpTtBH80FMhwnfxS3j+iuX5AiQ9r
o/7XsWbUSspZW6jBCnI02iEhzoZRrmoEXPnKoi9MaYsiAVszS2ykSRf1ceYG9Jc+
jCL71TPo+tQ2r+LBL4cVFPI9ENOG2j1ddhsqnQGTR+r0c59/IZe10U8gpeqSy3Oe
0ObiNzxlSimaHL2uFu+xBrQDTFOtcHWRvhU3pM7ycwV5FlYgoOeBjSxvz5kwvUXU
ULwxH4VKHI0iNfSxjBFIX22svsd27uduTvf/lDmC54cGJGGvt9SMBls8ZXQDF+JS
FIM1CZbQI9EKnxMfMKL9HM6x4PQEzwYTK2iM2US/RhMgwNe2kZBrpkwdrVct8O9C
lH7je2b8K1gBfCxLkkidRk6wyPn0S7uhhmTDPFF/6fv1PW4ltFTsJiBu3WEsE3rZ
S0lDQ5jgr29cpFVtHuqM55R1KBuaJXOjObidaXUlP4CEQRIIob97HCbypJmaBAa9
dBy68P/4lDA2z4P2813Fi/nGG3C75+aPqtlP31vg8KmEiPb7pOphI5zde2Goxb/f
odzl+KnT9eEWBjRmuzpcMCxE0TDJl9DrNtqkAxoU0o6k+2F4m0qCScZDfhBGk38P
Y9qS1DZs2wH58pOE/X1uz5hwdYkrI1f2I5BAG+aByZiO8vzaYtAgLVNO1+4JqS5Q
/qZongVpicWIp11Oxg8W+qWbOQWtEhU5Id8Ec3Vbq7ABalx3yfg3nmX4Bcsqiume
8g+Juo2L0Xwz/sSmRSq5pXGMguJdq025+Z8c0iPzl7orL9BuMp/htUq8spMK1tdd
PKZnAt1oOOXMH2MPi4imZnVfCJr3IWrdFFpsQn0e8fqaQO34hVaD+Hhl80Vcmnm5
g4rDC1V7+YkyNJQDqS8gYj8xzs7bkRWsqBt3DmQW4u1Ndmf0e9MfhSseuL7VxHWc
9FAY4QmGryTb1pBdeBli9Bj6UQOgvtUUG7J7DX2IEbcH32c9Pzv1LvIanFNKZrAn
/IQtTOyo1I4wE5aiOIwW7InX/KYsYhaDDggMNawaJZOmlEyRBiztclo8s45KkQ3d
lQXGJ3BKIivycuB6IkmoFE5PNtANqV5gc1X4irI5cC2qSP191/YXUz4D5XuHHLQL
2Dk2Rt1LzncH0nBmTeTY41VSXp93Alcd0mPhaJBOztBqOpoHN8XUA4xmI2GIQHtP
8uViYdme+oh0vHJUZVSU3iIr+7Tf3SyQJV4qfbal23aEik3yJ1mpghcXzCxYgLS6
OU6mlLvOxwNGrorNostmOWT8MbEli5AdneZkPOLvC0QmPiRAS71Y1Xt19V/U+1U5
yFRSFESfpos6xS134W4vdhvnIrniBpGaH9aFUA3Kr9gOPRMijk1nmC2Nlv+xyDxH
tXXG6ZbkRsly/klGfMI5ZBYmEy0VNjYujOKj9zGSKjU37+J7JDPpw1quybPK76nu
w4EnJ6olCoON5otPMoVZAw8usFRm/egfP/uIR1Sarh91XN+BksTlkVWTrU/cW9IN
uMkmMOAOrmlvpJafRskFNoSWqa2zwhN/Uiw79zqsewrksZy0U2jxKe4czRv8V9XJ
LKlRJUjK8enwSAnjRQlzFdk/fTjqx3m+5N3DB3ZHTgNNIav+Pd+sZawIhmv1XF+8
EEYjt73hPzf0AbJvViE+uUxZVIlIOAe4RdbBVU0NS3k3eLe4IvCclymDCnThcn9r
VVQ9RtP5jhZnuNh26ZLfs+d9auI/tjXRbwBrMcv3px3xr1JX4rzYa2VZpFmerXk1
R81D97MOvJY8YQY2T5qi1ohSyyvyxQwYookhBZB7U0B1v/kwQvtdqL4yGsE2kaUO
+UMzHsqBVorIOTSYvULP/suFTjmcKxdnuRVAxz3g9oWp8l2PKmbMIzvz8JX7ALIA
VoXmV7W3akHvoDWKH3nWcY9qD0AJxuB44+ZK/TbewEVG575FJIRMLPjJyUBpnKyY
At7uGoWKjuIjLIJuWqJP6IQzJ7PjcFekuIYRqqQFeHoQ+Vcq36J3v0sDVXLbwaPS
suZbPnnmbKFn/4FD7FU5TbzbyNEYkb05V4XOJXU53BLb7r8QEf2mRfpatk6Y3Cu3
6h2XuZC94pv+LKXQRMY+GRNMJdYdvy64n6mx6peGHYJUbSgR+EG275t6BuKSdvyh
h8LUqxwwspVJtV1VzusX0dzT9ECweWrL3W46Vtz0n+CcU8XDgKoiJwnvrvAXQ5II
GFHYuh796vPd54XiCV5vu41ioFkJSf6u1McwlqHRCQXlKwelFQckan/U5zZu2RtW
ng3g8D+z7WsVAm786/qmtyWSqiK4l+wdP4/XyN/BauvNQFNid+56CyA2yYbPt7Ky
LrfsGu2WOvOkZt2h9reTcDuDvkRk6Gbrc/abXMSEGSzvby6ryfJ/rieCeakafdlU
SydHySAIBwfM2yjNuTeXYbP5fAVHgre9vdXnLm7uDjz9+MtirlwAhBWW/+FxRuEx
LG51D1gWj+B8Po3HKZ5n9rgDwXVn0487MvtSo23IItDv8pMkFRQauz7KarfFJxRZ
zjJiPqbLZsuVd5opKNyx9PAGwCOI13E3l/xRBoAzoLUzKONqwbHAd4+3R1t8EuWi
e4rpOt+HrWMarjgSkQi1l3V1+6UyDP3z3lh2sMHl24bxjviSAI1XViFpd98bpzo8
V/GP+V5u+eZW8Fed6Ono5qzgCme1AOlUZaKZbh8wBJnPv7YWQ+GVe5xNeGSrbKJR
gc0+J+f9wqCLNVY0ab8T7MM4LaYmo77QKortyo85QvPnBMwYVx22o8cxQpIllQxE
xH/z3r5vUujPvFhBwVOZf4t404CiqNzZiD+JMCUYpjP7mtFBmejI+P5h6fimkA6P
q/VQH5crtwy8Bz9rLlmX6f/SH0UsKvStScCVXnRvjdKYVt5VSDj0tvNl13E/8jmo
lhLoMbkaQ9eLd8WaIsx0cAl8e+KiUxfSBQKUxqAjs6L5lDtNnzdgpFDjRncxiOPb
chde/Y0IG0p/Ui0/3cWzKhtLheD/o7T9pld/kEwdh0gqstlTjERoFU2ioR8IL0bG
ip62Vcp3SybzXZn0Yulc/bDcsCWYAs+wrL4HHk7YJQlKkXuAF5rN4NPNsFXOvZJ0
KlxSj74qe5oXEevZl6Dr9gIpsmPKSR8Q9/cxOiRl3D7zPqTP8c87iZB8g6TiCqUi
dAIzcVHS2tTcgzftqiycN4WN7elGJJlZS7fBfqEi/zFttvrW+EJn3F2LF5sttyex
UmOUfIV3nezOyf+B3zLau/wZdX6CpaFQrWZiJ1HS8l51Dotrp//JdfG9VBK8ksP/
LXymCXtTVO6NzaLIuEi6ovDmCpCOTqdbWfFhdb3gg50ZE6REIjuduCOW5YhOZhDB
KmLxBzfbiqIazTQqy6NUioAis3JMszNXp4CSZDeSdkGPnTltBYlMX8X3Bw+EQ86y
Y1uRa6iIZlQ4+5mOAjYDzeN87vJ2WiFByHeSfmzNUvGlqHatdSY1jA0eSgiA6Pi8
Ab6Tez0rWdPjFI5uMX8lA6161/lP4LgLw4wVztX01w8Vn+aGVTZNteSPxw0vACv2
ypjH9dEBqkOrCkv+iYXqLuboZWh8HGgUS5QC9dnP4A30nRVH45Z0oSOLc4ueHueC
WOyV5T+5LHLUdU0z54phvipzXhwC3gmpFcVqrNZBcdyGL0HSo07wTWTD9Yw22+dQ
+jicsolpPOSeX0srK7YE7DMRPrgUr3MCXLkZzxzRozCA8eS74af9cj1Hr/Vi7c5i
2fb1urs7FvzTCmWvSKYGT308n71yvvkVK3clOw8eSDJRBdSnsd7VLORPB4BBuiGQ
Wv08ypapT8oHL+9mwdxC7zKpGRDnZ7mjCNAvVZO/cInOgISeAXdhmR6U7H64D88q
CZHJk2FlXogo+t19ROX5tGzFSWFP8MKX5nowTD7Ov9Ay6XZTrBS40gWJn+nOotL4
ytvj6DMUYW5+9Mesa7vooPF5jcCtf/ehyER8Xxq5B8ycCjPJhZUOX47ESdGyx2IF
KIYRzFTVImiCcyaCJdDGmeUGKhuXuBmAdOZDp85oVIFiOg+DHltOrkQGjj8Z3yLb
6RvuhWQafl1BEOAWTV22zXYvniRD8MbLFg3otcL9S+KcVTfjNWdmCj2aRewOSJBo
e8RO5y3QGbTA6ch6vYxW8FTBKoGWVpM9Wi1vxZQAjtd7ER31gN6JHA/MRwhCJOJT
K4C2R/xIqCShO19XxZIH92XFCXD8BKpAlDKGhmUKLltSnVpZTiw8khLAr0O4HW+6
cF6SlhdCHHVzANUQh/bUqQJPQtCOLfJNBZe7sAeJpr4zxuW22dgxvJrTH+NX3AjL
Ys23fZ+fL7ErDNCnKewzW7p/FsczkqbY+Q7CrlLuRbPAVxXo07z/K9tDWMMjpIm3
MzBpYMPNj7bCpXMn0oR2hXHsNnyL/KVhgbDIxzuYLEt1nG70G/sBdBugCpv0lW4Y
NaBAvNbEg6cqUkVTLxhSy1vlZPkftCLQP3RYA94dEuQlYbwcmVc1FGCxswT0bVsr
UQGV4Y7RHf4Uo3/oFIVEqlAsWJEiqcUa5+W+PobM8NoLwTGX40mBJ/fDweMIn1Dm
NX8PeLAODPVYcA13Qh9NRypUdvvO7UIUEq01EQ5QM8pkAgvBczyC2HuayHdulLpU
jTDuJOlp+j7B21rK/SjDPnmNDSZj+LdHH07VQfjOyAV3qn2RIBnCavW9R+lEA0Oz
Amrpuab8L9JAW5pH/XvqiD72FsDlsqKYa9W5fb3OflCQVGrGdlXpLvIZ63PCAkJ5
CcTtl+ppf7eYy3cBUwE2ThW5EHI3EXKDQXSZECJbNCkPICtwRnH9OoQt4NbiedOq
6bkUlrwr/PjSw/uJkBj1ZrW2N542zT4ptGAzJUHWb9NQAiWzbg0/ITabKF69OC4o
Yaf7yIOXkRTNaWrKciWnlrLLPnAlqIKJ2ktgSA87R7ii+UcsH1+LJWt78lHAo+Zh
CJhBKceOCrT6pjZurbMO6Vz2W8cFJfLvxKhXoV02E4y79hK+rtmec9crmxbQ23Gu
xrJA+hInYvXEaoKvejBGFjCP/Vu6MtEEOFSoohEGiIYqEBLtrkIq3HhLE34ZhoQ7
RdiVsm8vOeLsLsryBKLprPS8YBsd1OxFEP0agxjtQ7fgkGIkVQN47Iz07s9bcrDt
Tf3uSWXBjQoGAs0P7q4cGPOCpwzaCJXblxifjJsn7jU4CQW2zEzgT50xt/FpG2+k
652nOgqo6MxRtR45jgYV/a35hbP30iS8xAT+Nm+tBAOzluYY2Oj8p42u8yRc+eB3
Pouh3Fgsw0+dBAriwHIIFxX2qIFNtSqk74jGTq91SUi0WBtxGaoCbg6bRHdTHFAk
rkxAQXLY0iVgdIrCXvsn0KsQ3uqLnx5l1qFIUemZlbRixTkV+XCNWdoq6ufnI77v
2pNKME2upgGePcQqRK248xX6E/8Z0hGGsz3o3l3K59683zZ/GVGa6CKHWx7WO6Dt
FVBTYT9kFJ5TslaEs8pmudJ/+kjG6iQubdFJvKWFeGCOnwcgreSab979zU4z7xQ0
/PT/B7hodZ5WfRev3Q8Of4zK8sEmDFSWw30vM98k1i1C8gbu3yj2FeadcXK3Q1Rf
nPIpe3wVjD6uF9ut5lZFKBxVWhQ8CVr/q5DnCI8iq89CFqAKyk4PC9AH8oLZ3FGq
Ke5ETF+JsZSe7yuB6eM7T2hoqH7glh1uIda0KPMRZbo1emuwKY+YEmgInX/L0SGt
i7mbfD6LLx3hwxR/xNYduVY2gxkX6kIog3OjQg4XaFPU9mcXmQ/cPCb7J3nBNAOG
86uJdQwkNb4H+U0aCBOmt5Hg89ov8T91Pl2ej5Ti1caXR5ZJNofLbRP+y9AifSrm
jaAuEhf/shYOu/PJSmBeo/WGx9vE1M0oRKzwwJcidKKYCkVfeIZOZT7iBF8U3qnV
b+mHxVUXOoqIc2bHS1tz8cj61rpg1he2JZyd7ObabYbCdMO+E0GMFuvPukVjpSjc
PwnIZOl2ZUEjby/Fnqx3U5N8bEBcLtwH356dRdZhdzenET6KtJUYaDHzK3cf8NuE
zxzZ3rIwo8BomCEMkimTv4njbw4VhON1FEgp6zPClQhl17sJ9YnbeIXsDHK77YYN
44KrjmWnNGClLJC+T/mpm5xVPhS48LKPq4rriDqILAYgERszUtqqUl2fNx1V2yDR
AxkudgccGsXpGdoUoAH4WpxMQp6E4y+ubbqw+qymyrfHR7q2XO4VaXe34mzaTO1j
eF5l3e0XWZTatYa+Q2lWYRqx0LiedPCjj+uyikypx8loxd8j7/q4BQiSpFoPqBFM
5OYEdr6oc/CqrGF5guW92ebkHQGMO9loulB8xcHaFBHINAF9fh6uN33ww0e9oCn1
JPDlahnzr14sLdhOxJSVvhOYeyLRMxR43MPILB0/Z6xQNQnLdKdTFrzLMDE/LTnW
D1iz3LpOFHG4dQwJXXzWJTJeznWabI1XNoCRKXEMKRrZKVsJyj6aOTxqrPHEybUG
5hdPP8ctnYVbRZSBN1cN3/2sSS5vrvEdRtgSgXXd3pu1qA5toj/7+Aisa/A9uT9A
3dpNz+hgAC4X+rcnPwV8hqgc43/5RHkKmhCJTNYip3hXj1+vicJw/BU5rKnYFrfs
nYcNH1E/7Cg01P8qKOK5cLCk0fzjMMJGxYIplesJ27XpmtNW1fCGynXv1gBiJC8h
m7iErjb9C9zkGXoApHVqBCBheCULsQPlzD+TbL9Hav6DGtR3M8MAZFVAez07kM2w
SWiiBlqoHeYtd5P0VpUYVTW2yhNGlY1l4gTyjccqRTPzdzsRsWBvYG20ejoLrKj6
bed5wl33IqR2qCGoiHOfSrvsCxeCn4CtnYlZw3pyFGTfgdJyIrmlqv8GEfF5Q1hy
HHeReqN/NKaOjUPLZFmfa4CYKMjDvC7OF0K6eScAWhZGswYVAi4GtkUfpnW1wmMO
tz+iFlRDwe4BxKWPGgTx6vU7ARVGbmO86/IdKIWQVy+tbUFEzIuIioZcDUgu+hQ8
/EaJFi5s50UDR685YrlHxseCHfNkTaSNm6Sa4NXJwAAmlB4zN49SMMOtfBqMKpxs
3taN6e0Sfhs17LlXvfEQN34JHsL/qij1E+eKGHxvTGaGjBkl9l1bxU3fjX62pGQT
+HS54ARmof/UJnXZDYSe7qBYxtNRCmr+LhTi6vZR3BhLtUJxFEBAGJhydJDxOMiI
d0rK/VWuO2zVLp60NpP3bqnyQpGcl+jnPAiUk/KawYXSUtp9Lt+wFxmVbZTI3FHf
IqP7Wy0CnJoWHXrwQCpCASMJH9fqGC1htc5jPjoTOyltxOz8gw3VEQrm2nhmtf3r
MiFpNc5FXXCJsEdj9Hjgds8gq7yjIq4CCZiXvbanwvGskzrarbvbBg33GAYDHYFg
kaQ2ZtSQAHrKRIp4EUIgjD8Sh+DjOdW9IkoAYW+1R93YzoJFmtMi1Bh5qv4B7/dQ
0ZyN9lZaccp16kG7rXE9KPTll2StG6LiaiUVPvkzRwAGiW5BkItnHUfoP+Mr3MJb
xyOlI52148m8fqFL7L7sftmp09IjpbggrpERf8G0uIDUbmhlA471GQW5eh7vPh88
OZfImJdtOjC2WuPxvRSifAe7OdydM0N7JaMDA1iUb/gEw775uTyx3pRot3BLaHjW
3I1UUF8G7eGuj7dVXdwZoDpWKVfL3GJF2Unmb1fRulcLl3ggZsCWYAFCyxYHQvZc
G4GHA6mJkrKya54m9kenqqzRE7+/T1BxsXhNbZ0qsguFt3JHBZ9DCHTqP8FcaazD
OQwppRAVIbWc5mylpApFkQ0JH0lhPLBXKDAFKrCzQ4TgAZqatWlQedeE/NLiHFGr
6QULn5YmXNWtI/53bqGEwywn4IVL4ZVnpDOmFS/TArAZZBZz/SzkZ/Uxmi3sWXi8
1zgl4EVxcBqoFGJx13b+Uxgn1Xn9IcOxj/rOk8RAOkUVwGBYjeofYO8XM0atATSf
e27yWDxpgpTURu1FuEPJNQJUjBT1Bmsb8a25+dzu1qHExhxzAo5XoJy719L9CHE0
Jz5IQ8zHFcvAAyj05Ywxzat9rTU1nsW+5THPSMwWVbU5IpWtZazlzVzVLUGt8T6F
35FOulNy+5A10t7VYqh00G2ywIBm0BSjHbDQ25r1iyFi+F/s6PV++YRQQ+TEMkaW
HF+xMjVzB2Ev+H14vPugcVpdYFPvffpBN8OgF68czbuV0aZitFGDP3KyfyD5vwJj
2yBSdA9nezKZxWFk/sB8+xLvT8urUKtgMnbZ1/N0RdiN5wVDWUbEXHKO8YMUPFbZ
kRVs0XoTDsMsIENiHwftdNxOHvinpF4EbFtrce3eTWwr0kJopS2cCMQy+unWNLkc
kAuTucznLhlqwaN7U21liHfqCpGZ8GphCEjLa1Le0ft4iHmw9Lm6ferqbXywB9B+
r7vtfCr0uOzjwsRKr8ddik/KZWYSjcTeqpDI1oo2iz0kFrXvzzULO28sbuPx2nbi
a3WvzpRAc3ZBWewNTtIeiZHnHdT6VUNzefz8yAPn4czLZUFHubwhJuIEbLr6sS5k
3rNW8IAhlFzUxZyvABYj6cuo0PX6FyzZMXhkjw3jJbNehwwZ40z8LHuxK4gzjUc4
xRkulYIH8N6C5nuGnElFt+9SW7i2lVOZwndFTAwiJ+yFFEkid+Qx1az7+/bEbq9P
SGMwaAMX/Z8Ebs8jWDtpQelW1MLswe3Ze1h2uDOdgIepV32SGztpm8cx6+TOTxwH
8MhjqDyEOoS4mp4d5ca83RXEpWI+Nd02AZqo4g4g1BQBIPpYIQqkbDZbd3TksjFh
HKbSgQs4/r5upG+o2J8/5gT1U4ba+pjyR84jcv8z7GJ45SXQouPLtaJZu/1PyZtK
yR0cTspnARziAjabvCeBqdWDF0aEs69kMZu3nDT6PhPGcMSgAlDq+XQhf/hZ8ojI
zaqeqOcXha+p52JR7M/h4cdDKcclDFsecOs4vbdx9Q8qk4UYksaf5ECXRxudC9+r
6od8n5f7+OxgVqudKl/bpzk5Yd9N8FFJZkO+WJh46jWE9jrXDgsdjNy/AXZXEXAx
LV+ypbfC4kne9WpY+qwWHS/rCYedTDmane8X4JM6zR5pwdLAbP1ORyNMiZ/s71eX
Ed+22hSLiN3UZUlcy4Fngprc3DLg/NreG0hrL7DtICrS2PHXpNKN2GmdKId8Fs/p
jTLBP5kTXCV+ycgIFO7m2gIdfNmKZEFWUdAIS974gsdSToV3eXXfnJnHqbeWOyOy
K4o3qXyG2MYD0rK/EngsYSJlMieBVuxZ/DSSnJdHDAXcYGYsFS1GncNCXuTeb8Kf
jSZCPnyWLyiQsawkbAM6Q+60DOT14GgDGeFryMrGmz9Hr9MfdUgSM8dr7YZ8U5Bw
vG+gSoFXFNeHBERThmUJQaHPZ2ZKCSgXOXwddjq1wD9vXOWjrdOGv2W2GfDQNkue
rcQAAHyhkNmuDa1ZDK8r8uA2XFfwk6o2/s41wQw7fvz60YAEuhePwRLZ6Nszp5S8
G9D0Wh5XmCEW2VFHiv+Qd8tHAb6d07fHP8WaHVyhPeTDU0x8a27rNwqr4WwqoVzj
IMjMjqLaxr1EtEUUcmoX/Po/26RVatEinnh+BFkwTjd0LfwYwwDCHPRWhFu4CGMt
ti2QUBZ7AnF/Lklgn2mCEl2O1nrvtzH+eonOpKcO20FWgH/Ym+pM3eq9DzGto8Jn
GSQaUO8ljb5JmAwp8aY1CqhlEzcX4HUDsltdVRiRUnvHazhhnDzYNN3oDjceJQx0
TC4Osq1piYlHJTBIGBNrgqQ2HF9gm7HSskgXCqv3nCj1YgOE+TyY1YIbq75xk1jV
B9iPw576JgQxvSeSIEJoMRiyrzuHuvARXxOMVI9bOx47abLu2G3vSlR5lewlUpAI
RXf5r+zOR8F5oOphQ9LmQdIoGOOPr4uHVoJwxJx2474wbqwAArAJTlcfcmN2PdRv
rNXcfI3uyNdY+8XWsAZydAsK/g6DI+nvQTQXdNutBjptVGzt88Dv39kJesBVLTuD
AUbhPCv5VmzuhLNK49QeMKgmxLi1KuQKzCec6XFxiILya/1nfY9XOBfuDoUolmbS
H/9y9ztXREsN6W2UaVTOemGs+S8OMKlOeqPuvTFA+xVNRqGtqejxLPOt2j6qT4Wm
OOLGL5Nc0UiJC1pT3V3tEQBA7ErrUX8TYfD2Ahk3QtwLERPr/1BbAlX2cr9cv/ZW
EpCkMT3587c6Y73JN2QoLGrbgb5K+ClD0KIgecUTjvh2ibNMd6i3TrL308QXN6Ln
z4+OlYNaz5akvsVcOGVYKhSxY/e8TGoYzPYAwc7nBNNUYFRPN2as0yS7cU5UaT1B
4UtVt0LKf7R+L4+pvY8ajFlM4elMpeoKiNzmfurq8OhVIvRVtQFZWLl1MXUL3as4
8WvvSvOP1vWRWNgbZIDuS9tYetMlW8kH8LZbEPGzM4ZZ1QSAArqwPM9RXz/+oEdp
cltXzEQgNHpSszgfbNHNOFMDKUZUhkSXj717vWjJn9VUNMrh41oVyWiWP5n91rwX
fkpo2UkNMVpuRK7h6AevPfNWQvWpVYkMMFzQ44r+oTXZp/Zo1aVLRBOt6qzEJh06
FWnnBZ8Y32ONPdSGTLKE5ST8o1dbjyKxeHe+GYz6oKnAIdeO4/9RyZWZH3HkE8g5
fk8faucB5CZz1JLRwonmM89yd2QD2REtXi1+Mu14UdkUom7Vh6BI7QKpFztbcx9B
YLLfRui9XmDtM0Faanl69qyq8Xlj9cY/ivhybdtPcfXmdv+h9EvnkSxo33Fpwcy5
fBMnlb6DeOMpt0t6mRzKD580tDiQLe4NBCDE+tONW3GdQevnpsUYn1Tm7bkpKzFV
KbbWhoz1sV60Gf8MW2y3HlCvkZtrU25dnLQWNIZlQ7zt0m2S9dSfej6QgXP2kKYD
eABi/85LQJVhzP9e5uy8/vD/9Ppshr8y5CU1/T33oL2Jixw2HlMLOJu70iWVhCiC
RchbKuzaVQ3t+JKeZhckNEPq8oLoo65ayedQyUlH1rZ6wH2TC0DZ+d94lyBl+daS
HggT+LBJ4HtbsB3y6KqEg4vtS3WK6Wz+U38ZwP9Ae+itJtDfbsRunWH0F1G1fkPB
6h5Cu4ZnTlxgeHwrFmKKkeanha3X/4QQOX8jEw0daohSAOZmVoXnc70CMpq+pvcv
hSWzEJ00KrtAQWNrDvfExGwwetHSYGvT29ItCB/bS7QRw4X1uBC1+3VP37k2w/dP
S5X+pAl0W2z0ODMWovmyRa+7ltsx5tNx9JJXIaCqbLSVB9PZ97vRQ7JdASJRopok
3zj5BltqTizMR5MKhPq1tzfq9rvgUbleExTv04GkI+40NL6aqrz/U0K1gliz65Jf
B5yWWBsKs9CPzNSXO0FE7KnZhRCMssc+Y7QCGu+NCUA4RZGty8RNsOsuo0HbdHpn
XEn2imENV14N3700b3YHo25D/KrInOfK+ff29qgQYplPkbLcvyiH53e9vjEAha7H
E9eRMsLy7N5H6z/HR1NZvvzaLdAPOcDvhTHwgm8AquheSCGSmbf66xAAfWlZ1vnm
JI0lkrK6jgEIWZk88gA/Fb+UeKTrElW3Jey0xIXE56YxMBMqOh83lOoBfVArBPm5
+n9fPxSgM0Qex5GrgPY5MIpWjan+eEj/Q5DOi3H84gMUYO8pVUrwv7KaH7beVyVa
zN4gv3NdYPjNpTQkK8mQY3UqpqvCWuh2hUqkMfICHaGV186GwxCxyandu7pNebVY
MEHstE0ljaGX33DoG4bNJtFPcj81M267saPXUf28jdawa2eOoUEKRZcXLIFpyo/J
T4LAuV4RanVHNJcoTmWjCSc6Snzch2K0X7rmFEhRvhLeWFAbY3F0wA1FUI/z1qeC
esx0D310OuUtECW+JfIpKnRb9D0EjIXJZPLK9ilymsBVxHS3TVwNNwhIin6nGLlM
WJkAtZ3LoRBoFQLJdHgyXqu1tnP3Wc/Wg1Ca48nhOi1TtIJW5iKcoccPnwyZJh4K
rcgEsdb3rtyIcRHyR/okxb15x9gDetDzKKUuTuods3gWu4hL98LN+WC27w8zeH1m
3tHmDXfH7t7lXzrmgAl4/ondxfErDajZwcNVG+qJRyRXuElRSleKXFx04SrVcbbm
bQznYtJ013xrjPKbUwJg55SDzM5YXqnO8hgn3xMVm5cfQIayJWm5P8aQQ+nbiTD8
cNvEb+6XvQzZ777qkLcIlbAauNV5ZElDoBifE+IAXBm4E/5sgYhZMTCqD8rlJJdv
adPV6CIYwGmWoGfobKnj1HfkABx4ZqlrTaiL+1Ytdm9rQftX2HIzVSWU8DY2lreN
MeBd4b4T4seMuLZTN5rTGRCxCTGWeqIyh+pRcCj0jQLr6UyE1T2hF8Lh9cZqW7Ak
6lkOscKuorphqMr+zp3KJxY/fxBSwqY0yYf/M8PNU3F2U47IU2Nw9hZPtMZK+suu
XOQ4+6wXAP3lOwDt1rNNMUeX40rt0lT4AwnsC2RKwQ2kwn4OYzoXs8jYyHe6ZgbN
HH0utAwWeb4KgHhONvEj2ZKNZcfscZoKVM1vo/el/Ncc6ukhvvsZUUNvJVg0T7A/
NKaUV4vieiZTB9evl5MJNKpPMBU/5qfDUW5OwyTjH2k2KJGBGY4FhbAybCM7Ebp3
pITrjRHoefjN2Pn4NIEQrt8eyj0Gehtr6puiPg9UPZQLAFOxBwzR9+DB/OnBh7HP
sqDk6ubvmMwT56VzVgaUCu48wWPOHNcExXIJWxMRgSLOoSKC3eH4TmnO08xD0rSt
OGR4RqTpgh23bI1ygZwUWowuq63aqjL+bw7SQDRijIvHgjY3ltRL3NHnrgxQcIuk
Z6czQFUAZuSR/ad67g95EvzxtIQF3HLOkb3W0ou8zmEm6D2RRcUDgxoZMpFvWAqM
MzIkZsDyw2I+zG/QcxZrOf0RkWhYX+nxb6XTqnLOqINbqilYhzkhDOyru42Y2VWh
L1Qtd9ZEZCWI44U6MBNnRX1SSSju5Hmgg3lJdUkEff6FPNh8qGmxbqgwpjs6nIeQ
TH0yjgaagh0GIw4WRLlT8JnfmvBxQs0GaP+6BskGl+Wrx6pBV/PeT3omKOKkc67P
xjHcRqxTVJtJBdvZrG2tAYAiKQWKbLVhbk9wdf5oLND1Vj7JDChK3fydui+6vK36
QeFmBrzync5aJ5jQj9CufTkFLine8bwoKNZEwpvefPdyjQlLQYDk8J+mXIvM1Tyl
aDUvZnSRLm38VPU97jswZPg0Qhyw/UnfrbhpbqZ0CIHzyn8J0zU6GTVz2hzMGrAV
JrTWIh8tn+Js6jYESJX6lITcjE6NSKJVDttrOs/3eOhViAe95oKA9cnsoEJotoHt
JI1flbvHomrpbEn4hKuOrtitF/mGjUn1YnBpMaiiFu4ofRIolwiUER0vwhsFrXmf
tCyjoHnj3ZAIjZZA7f/3Lp+wC2kjVBRdhmzV58qvQaTN6uoP8iucMWXxkEaWTh76
SZjRROHj9p4Id5Fg6clids1O0HEi70+QVlUzPhmxyhowLdmVzMtn0k1Hxgj+1u0u
MrbVrvlTsQaRD3DEZSf+ufnfDrejh+GOBTqesaGClgimxL02Xemabuy/zNiKbJGN
jvy7x/9jojgKZItiKXKnqOaF9psrZBsiYxcu/7Nc/2yiFHoUtOl0KQXZRz9I2ZR6
hv3s7lWycMWb1qoHv6LzGpsDovT+O3O+7lh/OvK48248TPkfqzBhpk4Xvt6C4fP1
gqzFA6Rp70DTmXu7dEM1QXnVM+2RSg7NrpD2YSy60FFI7TVZ/lhdS21Lc6to4SpU
X69fChqGcugRGBZTWU8o2tPqS6zZw3NC2uc1fPgR3bHPu0gDpMDXwyJu5lB+/S1m
mI+77hMsi0h5SK80noX/XA7bKSOQj2CvpqNu/a4i5GTg0TXf22z3bww0pfnEKqVx
8+OFwau2VkznPmnyHbd35hARwrtjUjWkkw+iKWTKGQuxTIb0J0OvWvvVWLj3eXJ8
57CLo9m5Vt4W+ngmu0IRtsfdwYPMVnfwbFxjEjFnBWWiSvYqv9Q+wRqkce2xvxhp
dlxbmDaD/7GC/uvS8hGry2YfSI6M9tHHemLRG/vEFIA9VuuM1yEeEpcuf51Z82U7
KbmeCmYS6i70yFNqnp+2jY0fzkBs/o7gosbV4tb/saulXHTfuepMFCSj2U859dGz
V8anHzJy7mEOPyLyJ9EuDgVvKBQ7DIEYlwqN2Mc1DNhxgo8v+derRLM7JewoTOk+
m1xSVHzS3MVigCfRbjLCpN0fW2SW5Q5VJU10E+iCJG089yF/CO52g3n1wvFvy9Zy
dgdzzt3OmP9agjikQjsi5hrbSebyGAhH51JFTD8zQ7MU6OpxwYYJCrFdX1L0jeGA
V4C7c3wHt2t2ECtlcxOSaWgVcR+g2st1qk/YMDIA+4ltt4Qyw/dG45U2w876bf11
EDU5vGP2IG1bsCxNbdaF0/AAM+WRdo0ccbBdAVfLkoJFBRpQd14jCFtpZuUIdVVH
GYnE/aiPfBwIaR9/3aMs8shRlhRXmzi7t7iS/PiwOG0mQyZcGSk1/JagxjFsDHzm
0vNzIjMRR5vWlb/ABvLzULEykFl3Hxc//fq/DT/66+++3JHJ5qHlKxdvHQIsO21G
wfzXF1ZYZRJuWTh4mbuOrxpz7P3HfMcGWp0jpi77VIs/SilfpAFju88r97xk8smy
F2F6FRURYkWFcxbUGFuVNqT5QN+fuBKkf1X2Z7R6VTUPbz6/6MzHXIZBJEJ2+JG0
OtoSGxjuP8LWyB69z34Itys2uzmk2/80ftGRDwzRcC9i6lj1J6FdZ7aXtD0OxiFq
jB4u7BoMhd1O1TNmLIXw04lIPMHFDydpU91VsaXFIdKE6iPZOuIDRZM1rN7f1EoK
2x+vDZNBo39tniadlt6AU0pTnvBHOzGOgstRyAXshsDZisjVEY7qI9g4CPwoYrea
IoYL0eEblCmBeibe6+Gd6HJtdrrMT1jxxiF6Bf3MR8ZOclPB7xA7LP7wOmvOWsNH
Lj6DO7AKht9LSWkK8HUnouluARJcGjINNo2SpQbhxCicZALTjO1h6VOFCcYKfqhb
H+KFAXz3NLXE23yZP4G5CtqE+8H2hbEYARBhkrjoyP/yeigLSIegIX7p+xioMeGI
D/Ut8wVh2XV6kkLs4uM5hvxmAKa1B2Rkpph1z3vupd1daCNuU4bIqmDFhzOE1nLX
4g+R4XKJFCD6mkg0hKAPuctMqZyP+MTZdFABbMolmduU7XsnkyxDMcMfBTc+zJYN
nE/Bwk1AFWm2URSgw5ZbCMvEErSPupK+ZqHqUYWQh6SFEgaZRsiBnW5JlaqVS75k
QAR2jj/iZrH9dRDRFpVh/7aMeve+OWVxCDovEy3m6MAEZhY5NmY+Y/hNJ9CFH3dI
X4m90HyNlxKOYMk4rmvIzNWLHWdhFx2t9J48nUUtq+d7m8A2n3WUcLYXhgp0usYw
cI7vEPoy3z1uQ4iUsoT480w1QWyPcGdp3bQ33vljXj+VQOv0l+zDs4Gwh6MDSYde
POkULTwF15+Iw7OWuP1JCPgtz1k2NfJTOpn/6DRBJlXuXf1/Kn6fBf57PyjOU7j9
4WwedfsVZZMY188E13XUYP0EGDEIwfoqculzv9LMnA/D0H2HlNkVDE26X06YiLBJ
6XT8FxjrJIbGnl4rMo7y0E9VFH0kGVKC6ywMiDsJ1kt3J+ick3QVbhgKtQ+LDQuh
CRNv8PgInTzC9o2t5uUzk5liuBTAnrUuMQA+YZ/xdMZHBsuDK5QkVQvfDDBO8OgQ
VFzmCSziXNklwns15KcqyfbVMmM5GKqbkwAhTApJA4q884N89CWFvLTB8LFFesmr
bIrRGhs2Ihzt9bsWVjBNPvLCecDE/8/vq5dT6LmeGrSC8GaiebNdY4zN4xjVUj/v
Nh5oXRGy2CYjl0cmCaZ6c/FlgsjCZ4HbHqmm98WN49Jfh8qIwF3v1yNGijYpoX4B
NumCVIA/USyWQ1TWQbVT/ShFlK6OqtcyebIzCZk5/HUtM1rQgx6WGZN1lNsrqT//
OwPQ1Z/pV9j5V16Q9v9w6BlbrNmpy5Cnu1oScJlSsY6toATvoSYqo3+XneTxzg1d
PRmdVjWbPEOSvm0D0gKEcMD0PgS7jaiRQc4Kxb7pEnYTbO4LgSLB7paOIQAUMW4g
QlwMTWqhd8JOd8kph/lzpvp49L85HUV4wu295ubQRuF2U7yXHxOan4ak2ufhurFH
jOtv99dDScQ1BcwPhmsztpFEXxPR+agS+/bmjJgcd8YHIpkf485CQ1vwVlwpvZcg
PdaPl60J9xAo+LXU6SBCupWAptbZgm6R/vE91XpTJyiCLldIa3AVqZJ1yfjkTyU2
O9ct96LzJ0Kn2elxus9I7gtRXbQ3RrluGdBDRuJIm8wjeP68CPJXeSl6dPcRI3PI
U1SEzVk9cNJsidyDFZtn9VbfMqkeMsIt38NZfSUCYfMgE8RpByoxUlCDd9i4+lBH
SCw2Iqamenw05NS4hN5Kt16Homz2Nq4/ht7YbMjtNj6FdeEJAbzqeScbNjJ+FQnp
ZfkOuNgRfBObKbCX/T2qezlFX63eKJErei1ptsGYBmKXSMlbaR9dwNesXZxz2Kf1
V3D3PFaJTQEaBwHS4l4rn12bFUC6TDt+A+CQrzm0ttx4v1R9mJNKvcjq0lTh+NAq
qnTzXayjGX4yU3er+xPQ7uiL9Drl2QZp5wHStC7E3E5PK1j0rgo5Tia9Xdz1D37O
8zYwEfsGXkmrWyaaSieLKlBAEp3Gxk6JcOOPZjlPulGWbghF2KJ+Sffjks1DS+mN
QmfhPYGSfATkFonII/t8onJEXZDsaDnK6JE0YGenjh4xchCssZbafZ9A5+e1QSkF
PX7t8BQmCJpGCgmwhDECKqb0+SeHOdIjekBI3CnazUFtIYWkZV4ikgI1L3iCQNqo
+qVdOtWA0o7jF7RBaGoORXpxQZ+T3JykCmJ+GDvzYd/ion62aPEax4CWOYAp6b+o
4uDQX9kHs/YRa/Sq0ceUkHJafE2GXMvk2xQ2EJjrQjRo8oGOadZLZAdWN48yVCx/
j2HQyqy4OTqAsFraVlXYk2EwJj5A2NVeIY9Y3JZd6uHlwaPvPclMlfD9RWsP2sXE
Y1b/rkINtD8Wfg0sunH6o5nceobswUdHMxMSh/zduEXw/w7mM1Ro82gYUC4vLKiK
u4F/TlOke1xZMqfW1T1WULImJ0t570+xiX88TQaV52BwuIWfvS6nWIOpTcyCmDYf
wp5+L/LNzttXQJ6hPwOa0MrVJwjlQPbmhp2uClc2NknSyGRRhCK8UgGyritnfxgj
KelQKxOsDKXXT+j8vHKuCp99VPRYmFml364/WabkKIEAaCX0+LZauUqVM0Harbik
4qLWMzwRxPtxpiKgQagjyS7hgsZgwWPoslMFs4A+KntBhtLLHxQb8wiBk9WFxJjx
ul75p5N8SaqEhbTaorOmfyGlZDMCi74QVRvy98caoOQEWRXy2xI15b2+2r9NwNk3
fWhsDuqtmfB3Mvahv7PcZ3dvY1PQXipWjVAGcDSOt4cWR5clv49xag3TgJUeiTt+
EjQgu1SltDms8kG/v5JXMuJ6bmiJjERkKikdJyYOyqTKgtKQOs/vu0TgePkFC9BP
aDWTNMa7ToU2S1lfHe7Z3o8zSWgViQMAOGbTYOlBbWD9SAasxzRLNxE9XXA5pVG6
JmhQwY5IjzPTvJHSVRPQXDQe4ehCM1jXC6QbjQ2M9KHkM4PCZ99AIa+IUccSJqR4
h5+mO8+eroBa1qdMTgAkLSbO1QkUI6Cr8NMjyUSrW/n1n9YUS+lEbHkvE/YLAQm7
eZeaa6n2xrcnJjm1hY90aZWjrpogk7dwEqktmvHJzT33ehFuag8TGHFo+vZ0+a/L
7jqGaB3BzALff+qpRGd03thQOHgoLxWIHSpyi3Kqt0lbqrhXCpjnmkZNAiugpI6t
ZxlkdGfBc7ZgypgIfdKZKFRWVlwsNEnahNuumY/SBr4yL64hrA88lowuy6PWaVdR
WE6zULfW8F5pirHwkR8DdD5OMykokDg8xiekoCOPvTTOeQcud4/v//ErfbIl1DsK
ITgkD07zw3U6nLwCfyFSyU1nzYzyOAmBeXvHfQ2D9sjQhPadCD4+uQ4JclvuATZA
FpN5nTF9/OqUkiLKFUwnUSBANF5TdLHYChxyaKhqe77c9tckefRQTvQDXiapGp+W
1at4Gky/XnPniXJisH3Uv7tNoB+RjYS3nMbqwiBiP6f2ZIbuWnfK8WxPzmiqHU5I
ZcGw93Nmf2ufi0p99hSd6ghnxZULsCPxYcm9L571azznORHOSFPlR+NZIiAgGrqt
qL8djb9mxYZUNM7GqjsFoDjUSGDZdY6K/oPP20rHxOUoVZVsemw8wJxgKOA3r93L
mSVYEJGdVtch7VMQxqUAqZZim+Tpo2lfTIYs4bwvAUvIGWwMIsQVqPF+iVsn/cZ/
boqpDOezWtt9OqCgjKZFqlTpvN3fg+xM3dpZmf9jZOj6cfoZFBj3bxr16EbxyFGD
cL8L88Nq8QAJt0DEImh1GLVzhBeBioAcUg+X3ptZS3QDErAzlXaGpgpqQ1Y8oT6K
lyLHkiQRpKiLd+mEf+PgDlfrEQiukEXUCG1sJhSmlfDC/iQzyW8wQ6rfb8sx/iou
BCNRdAv8MrTiFqxpfs+uw3rcRUX1V8+VRdGhlepnADd/pjS7zmYwLmRUogZUlonp
ksiF+VnN6+D6xp3A7qDTkTaheVgF56DMSTe0UDmZTm5MjQocRsvgB8kxOu50UC5D
A5HZx431QdUEp5hWFsAm9fUh3wKGh+K4xgFdPgDzZB4g9b8DUN1BUmvMmuoMnf1B
Pbd1p5WSp4BkDsGBDtfh1cooXxuEBHCP2T1n+A15HGjH2hoehm16/U4adslX4ORW
Qf+2843m/XjJmWy0wtxVxe7euSOIkvVUpbCOqfO3yVgkwyZuKY3ebfxjEsDPOGF+
1IOyp9m65reasc4erTcHQW8CG7NKqroKqfoAUvvsl5C1ozS/NIIwWgB5zvmtjAsI
DzADkrX2LihUemJkI3PIFCcUnbaxrJrFbH2DYkxBRlAkOcCeAmF4Q3rHe3JLJF+G
/yP1Mb5Jo98eS/huIpNOx7C32KXGwIf2rO/Jrj9Bon1cpfHNFcbW7/rNzmmOBsCg
FcxoFPYEh0VY/4fj9YFQTnia12esiDJtkMaPqzl5SoB5iXF3sEedHQCi5Z0QjH9e
cwlb4TSwT06YtHaiX9BNKeZhjvjqkHLtLVOQNz8/4m4Vno9Ym86C4ADokNH78Zpb
3TGnIVocUiFNiT6rgIzV5bnMiN+1PlHyqmabYA77W7h6MPKz2rhf6H1DFDDJIB3H
aDx9P2rzWrQ7yrA9LnQ4axTxVno9UqOanB3GrxNYsa16rx6wNsPxeP6SfsRActo5
kAckZez7XeE2D4UzA78Vv1fi6kCOIeJiUgQLuK72IOWv7A/LfHNdXBOWB59XGF62
GCLzOEt9Qy3WcmrbtcZEje9nE8N/ZPr2wohR1I5SeHV7NumXrKgHgN9e35zmrTHG
U4GoeDJGCK+eckkoCGfhW+OhtxvhWnLupmoi+nzV5WEoag+PJpAWTU49XrAJqJ92
+GO1w09X6jWZi2ZV4Tym0t5LZiPctq1O0+eN7A3lmEl1fPz/TvFu7xR9W11pMtvk
M7Hwa+kCw5jBP30Ep8n+vx/uv72w9DtMg4nJGXgXCKOYtK33O/jtAxyscxms8Gxz
+ZIqje6ygQp1saJOYK/uft+TKo6yVKBsvztOr1YHhMgv90EOMyXDommSv+2dxLO4
lZzxY437a9xDhsoMhw2qVCZ+SgUlIsowi0/85dWIuYuAc6esdb/ZbCm5WSANHXvL
8T487pufm7V61BDl3GwSx+LVxSlnLUMw9pDlwwoQg15NEJBXfYk42h7rNdvJ/tRH
uHA1LTW9qRTCxmayrWqRH+VaJT/nQz/nBC3qeN7WRLGno+E295PhBTKSHc3Uf0mt
iTNQNSCc1Q+KKdyx8Zi6eGsBfarmm0f9ory9bsCzSk4mnvoJfTIUdr/sR/LKuxRX
rPRIfj8FKsOL1K5F0+fxghCj2DH7G9MFPx80Pl0r0cVkSy6n7XP1n3TcDmJxgxF4
N0CDgLSp8VSAJMmyFvY9CrKCJ8e7o/zpuA0NnDwIuUbxW84IxJWEdRielVDrJ9Vc
XadUz6/X3d5CFtM0adIY7wyCsm7vIUuvtMLitqWf9b6RVqxUTajwLesZG7n9oBjI
GXz/ozD+XzFAFK8XSjgMNJG67ToD2WVCbYiBHkaOucEcMZlD326CsVvhHPihaqBK
z/5K3y/4mWTywvo3438k/dY0+swenXU7M7a3v36pB1/puFc7w4p2qSqMrZbbOwQs
0UyCG/3uMeDE9WIJYi5MQ8KcoC3mIsttZcX4oxgEfpr6XTGoS1gEhDJVgXzmQkfK
yaQUnMTksPb3CJ8zKDNadxaV/BM+IeKlXilp5q//Ahuk5jbvLYscF9ybuN0/4HD8
C/ZHV/hEvZ/Vz81XyOrKGDRI1nsiJ+v4i8681D4c1xWdurRZUT5+Kg9O+gLweyo1
iR4FQk5zI6ijjBwkvb5062VhLVXmu3PBTFUAvPe7ILvmUBmvg/XdkY9IxWGezZlE
Of0s2YW22aF/L5upYXD4Q9YNWtw9owrrQH5ggU5bDixzEYs3ocl8ldFrYdA97bI5
3FBi61bg0NgCqR7oYrpkf6hkwgNszgvCyQp55WMOs2zNf3qbssep+HmVirULRAlC
ptpNGvt3p5aw6W8RwHdugsC6CvtaycQjkYb8g3+jYCTxzwq0sXQ29ACJUdUECHMb
4lQUCU1dczwdM7xPyr8LZKjFvffhJAqpIifVCPtP+4waDcJMBGlTyG+K2YlV0TYc
eY/1FWMAORiyTkwIrIUus8ikvySYZ2jL3nJ5OwwSRS8qKkIrYMK95b3ADxzILu5n
H4unmikaIRM6WUeIUFxdKaFHRbR21Hg0+5vyhB5mT4U1EnqaakuH8y0OBVMyzF66
jBlzN/tkSx26nuZfcrRGD7rBaR0AUY4uVZ+5YdjMjZO3qBeKqp2rPCLG09p5MRnK
auKNltB7ZNPDMGXOgAYCtyaj1J4gR/fwdGM1Foj91HpnyYDicEfEyX4tebYgZuXV
4hbJC4xLc3oivVDMaMFtabZMe+S9RuDteRmzhXGsvRJEp37q9o7cOa8S6FtFATrX
4hhVin4W0bCeqRfwTYNyisE1hL+Fbi8JhFnmm/5AbffsAJOeSWE0RpzqVZImksGT
0qzILn6Z+4g1Uo8D5QEdjqOmKNxta67FFKlETWheta8vaqWckh1Pv3DsgDcO4CYM
ygxBBu35yF2Kd9k+ulveUcdop08Cb8Lesr9JURZxgnlDBvfgBjBm3lNSGu2/7UfA
oQcNrFN9vHGSNiwnJ9BmNZAurRVIyQo9YlDull0ZjfrZeaCxJJa6G/C2AVxtV5zT
MnB/m4rTjUrqgM8H7qE99JIz242H/DaR5AZ8DTeyRPB5NQhE5/CGO2SnibNVa6AF
absVI3a0OP1075N+bPewohybvqAEfzTXfo3HXcHx6f18/z+TMv9e9Xhe/qJaZ2mD
AK7I1hin2GsV9jgUIt+frrPdG+jeGNcqXROCy1dsGHTcl4z+ImHfVPKLSS4wLZwn
SDoQT/9See8pnIX2uoY11RhI6GNVvICm1JLt+pJgQ4xjECFXM8dmKnZA5IVQ5q+a
o3edxwQEbAp/zE0b7dq+QRay3Tt/h6SEPlG2dhBULNjPONxsZfc67bI6iielYjxz
eiBk4fmdy5MzBGkUneuJdTl3ilmeji30alodfXouKnV6zo73uuRjvOXqUZNB4TiT
A7Xfwk+CjciO7dUu3vDSYbiSIfVWeiKapo+vLLHr3mqJmBaL/ZECsHO+mwmny+0J
4oDO7eJrqaisAjO89FI3razWfSb5kL2C15vLIzoe076My+1+Lbpqc8bqsBDzcn0+
5dmL/Xzr9rAjFF11DASRn0UyJtfnCpfXbODSxm4VW3awfQ344QWNp6l672KteHaO
9bmop6ZUsgSrIE/6qISkEyISJl6zPX2i+qQTyemZVZO0wktBXB3NQBDxXWz7j5J+
sYaw97M4bRp6MO34zjC/lVtjCiQiEP51SgAVZ66EoOF48tDgSpolN1bN4TBhQSfB
SIx5sPX7ZsQ1H2I8V3wbDSL4Mx7DNQeVIk/GP3P9zBjvFj7HKv+9VsS/FcQE96RW
nZiL8m/Ic/6dPV5omZkCavk2DBGR9LFvZq7xlOeJElvh9xl9UFGX5F09m11Co+Nv
fQNnCTqScCD6kfVrQjbeP0Pb4PXChyGErUS0HzkFvSEWMrFaPmD56dLRZv02Ah5t
un3eG5+xIwnLKaJbWUVuAzZADw3XgnQPp5tETZlgl4Jm5ZlFALs2lFXAlezGwny4
JjfBdls5XuVbyPnHjPzk5k/qjOUE6VmKiDtG/eZWOB/T1XBFO+sLZfk7P/KDDJIT
Lr386o8WivdTNK4vlbwjeYmogHo2PxbRCJXaLfZiBpazW6sbmd81MbGr4DK7rnRr
6gbHib9GnKLbpKy2X5d+vBcDAK5ZiX/mE2RYIZOd1taFN3y5CtB1e/v1L5jQElqb
baums0nOYu3LWTDP1oKFbpQmudjn5C88qxlaxcgGrLzBPwFHf2oR6dWE6wM7PuCh
drbyJ/YGohZLhp6OPM2+QnfRCDOb9/Zr/iYi+ax80l6RtCCprJikjnvB/T3J0y0r
VyyMEkrsvEl1qea8GNlQIGmj3kDJlaBgLSjOcxNoXsqHiOacc+mgm8IO9Q5QTl55
F0A4jij+jDoybrL7CxgFmD5ypVK8b4QhlO6BArI7uWN7wkWPvcsZ5o2AXdSpWl8c
ieBurxBlv1n1p1otvFJHEE40dLuDJv/yr6P8xCQ3qOVSu2/VnC9Qlucfb8YzSjLb
RGdrIU0i6MD9BDa+nyQOV7wJG4wsTjZOsRAiRP8CumsUGS05rZ6hI5vuvXkdFHLq
gaxq/g0ft2Usn5MgveLkc5a14dVkEVmSXkyXmgXE4Xnih+V7BD5pOZnN32i/bpzF
m3a34lD/Qzex3IxSCt2nDlJE/0UC7FOplmGzfwviaAJbtX4yFq+2H1h2CJWuL77I
kz0wmclecP0IuTQ8wuXaS8iUTNv85ZpuNSGCOLX+uDIHdmrLO3E10K0Zx/HDY0lO
zLMJ+I/YgU4AaaXjlyjpRzMrquTb1lVonJuOqh+rIaOxSEjyJTXnGOMh40vdBjPT
JKqDmzlcEhufaU0NhSwlI06Ro98oLAFD7d02/js7Exd+9rcwS3B4KPn9nCYWvrNg
FLlUX+wK2nhjNovsF7o9EgBDC8Owlrv/SPGA69XQn2FrfGAZT3O8IAGQNAshJhp/
UrZ6NqGFW0mtPqCHHz5fq3tzTDhSoLfRngxzqZfEDAQIBRT6lhrjF53fB5Iq0gzz
Nh8+DNY3rJmZplpQyjqZwQrD8xnR20p8y+WsoGKooP8rJHGh+p6IuexuZ386T7oh
r3kvuYAvguVHHUSh++yOIlK4LOtVGnx1cj+dU5TV8BoIBxYjjgLM5O6FmQhf0ONC
LeuOoIzmfxtNUYb3SVvpCJV9gxxx19I6l0dnxjOv+j2KmDJWaqPYzg8zb4fhwcVu
DOVOYPsdaMPuQAl1MjTWwEdKfKJVgcq+ZXZFfuMTF0YgL+dZ2LjaviG0YGfigCas
T5HkAoOLVcJUckhjDcha5ivjcBEEKcOMckxPFDla3B/psTD2VU6UAzVOpUUJ6l6+
1uNdE88wvTXAnnWjQpjW9TG0FkT8I8UQeQGzxDl0NMJO6kbtxcmcCQomTgO5qGnv
n78mxqRPExcT9wqCfj0K861gZ3Tcek703oVTf35V49TjlHJQxxuOLBYlkISQjhCJ
WIDolpR7jJLceUVDo6CgLa2wkaRFpK1DK7vIV8wzobRYTMn0/YevayC79U7Zst4h
9+gCnvof7XG/P00jxtK9aOOdABobSqwLWvpg6Q15Sc1MNMByXoBao4weC7b83yBW
HbFe99g97f4zIumd6BJlE0+bAGCTeoB3Z/UeKhGLl5YJ+ubEVyCMewEo4K62jtGl
/tlMbQiFBhd1EuqrKA0ph3fCanu/+VO7Ut+G6eDnWPC7vJZmdrnr+IFOCr781yBX
WWIAmWx19QT5//6eq6mFN3klGi7//CSuIHQ6lTNQMnpoqxq6VSN3AmPnbgIQKlYq
kxUitQtWQeTC2gz9j+4QcNqQt9UbYKHiHwdAlbaskLHbR/4pRPjf1PKN50rIgmqv
Dp53pXKmzAvrQmMWepCmlBq3TWPSk9HPfbcIH/2FPv5OFfPOoINSLeJWj9QIuqri
9kJIdAHZ42KxvUijzjSlTJdZUH4RifWxoRmzZyEKguEq8qnTNrtW1t4DMmsQ8yjB
pHFAhGw0hbIsejk7KrIh5yzVGTikQdS0ZVVObLhxpJp8ec8Ecz5suxTLI7V2eHON
VPNY4XrfRe7CcwjtArlprhG87JpCBgUxIKgTYQ/+/VpeDULtZO+BEWSDepUDZBRo
GuWcbSx5uwDmeeNjRrpRMmURwH66QAOsGCdIr62z5PpjOrs+ejeQCsjEvshcqeeF
FqSmRT3d5FqyChTcOKED6xWKWqN6zetPpNaDUdaSIExpm/emGfZ4oTQRZ8eCoNgt
zVN/KxcgDyfqdKr9wyuBi+r2aqN+b7jNcDeHCxOafVYqPZjjFBWvLA1rq3NdX1EQ
8idDCRe6GsbsbmK8BZ1rOoRu74LLMWG1L9Z/5SCH6CYJNKXKoqDDVo0EkhSql6TX
AQgpKwYY7zYj7mpd6RPxI9hGt76sFN4KMx8RQvZNLcKwCbqVWq1SKS95vH/Hy8li
JxZSvtLDk+JsY7wkf0fEF897+1Kygg+XI+3XA/S0GJaTqjsXvIPKLzVemMnURe+6
ssxChvtIIS7j2xZWKpa3WsFWRQpWTPimQjtVmbgbzYvgpY9JPu8M4TY5JOB0MLTJ
Q/GOkvYCrPuVp6CMB4D2jkT0oA10lGIIG1VJazxwd7EAz5h4lWM55Wf2ytyaLhaZ
p0KLTG1cEe632qopseyz5ZW0adqajHg/pn605n/lJ5Cfv74B9OPTm2LmUh7PRti1
P/AHa51pYfshhtTdsSUPZkeeeTorbx9cKtWXsZQ7wcBX6pJn5hveiVJhJn0f6+rI
192BmG42gmnX7FveAIIZU+/BgF5EpQo0/Q0BE+8XHNWsEJVTVC9oF8Lpnx2BA6EY
LCLtMu5BrhiPCgK7SFGEqEf3KVJJ687+NdXPqjfXq9zPNeZ9AUeQG0Tv0jPpXfwK
lfeGg8YpYbk86fTYGX7Lb4QB02ILzspqU+/3NEIvW0EtsrUf68u2KXgD3Xs79P/u
zFyrKngOsHd0I4zz0aa0aYZJH7Iup8loRB0YW7NeK9yCXcfXwfYCEsM5mrwSlZs5
979Hf+zc+QmoUcwktzXcaRqp7Bw2g7GEbacfbUTPc961BccN5Ci8Ukv6M/m33nCo
4m2NLO7m3fBRsEckiG7eWJZyCZFDT+8W2IWMn5rrWiwv54X2THZeya2Kj/kSRyBC
nAgMxO7GIUOIlak2h+DQL4riN05r1spjkdCP6Hjg7SCQIe/8mryXsHmq+hERsrMO
VChxFsMNNKK/TM1S555JI9oTQAYdc64MkMz8WA7yFgIROV51NisXN4kLcFowGZvT
Wo9bzlztdYUw0Wz+TKOgxpOVmIXScxX+qu64V+D607qA+rc+7JQiDp+ttvZnvNCM
EkOtc090RbsobOl655o1l82lMRujUZJcCRSaGtqghymK/lL+AwBbSwt+vwrk3KmD
CLryvgi9MakOkwm2iOCgTaG3dTJIn4fZVu6poyDe7HxUuTNBFD4V6TkRKBLLWtD7
LpY90VlUzWytaJehBZX83EN3WeRK05kt70E/0uM0HbnQoHND8ugrGjlyr2XOqvxA
f/sfcd669h/5SfMz1G18fhHgJsPwWxe6wUKh83dektTWsh0OtDlztMHQKyepGKFB
YOADyFCWqQReJnFfM59uXItcTv8yixoijlq2L2oixZEpoGyL01H/vUHb3/JYADCD
qQirinU3+IfqkzQFHDf5zMUs+uGDardlvLdOrP+8VmPPgtrowrz96oErWraHmtB7
Msp1eLs8TIh6kXIc1zpvpqctF1T2sactE+d/fOGesERxNJFn2/bOZ3I7XR0HD4y1
/ZiNhfwAZ3vUAGZ9tC70XeOxcyGSkWkyeMEX/LEl3D8XnKQEgDWzJMyX7cRuLD//
iG/7Ar2cCx7bIfx6RPTtvn46t9Mbah8Pyzof6DVaZOLPusRKmvYfZrwItwkoKxNy
AoNngkbwZljG628eXyO1G9Bx8W5Y5ReHq7BaH/B94K3sJTH75RDhsPn9DhkxxaO9
GyYkj/ZL0NnTA/Ig54N9EuA8zM1/ixNZajnM2kIaJn/k4bUGbmhHah8CW4Icv8WC
SrpaU4Hqy9Tdu4zbkZ7MkSmyAFH+SNQOi19lMbWMDEq5vDkmzdnEBFEtOab2vc5x
gYdipLRUvVY/41uzKWQagY2zfmEcZVcPoRpchzbJQhWwV0WxO+MtbIWeDudrt+gA
2yfrDYrbYPec0I3zZdfZrkP3Z5SItJYPWGgwpy0rPG+j9Se+gJXFqnqagjKy8Ogu
kch0TBBGhjt5OsVnmKw6jQNyJ44PZnswLOcPcmZGafHXBv3XLhNq8VVNqKBMz02U
RN4knfanQ58Z+HsT02TGGnevn5XV0+5PUZVZs6i6M2Zswcpsc/s1n1OIWduhfkp9
Lv1svDG1YVzgZ3IsFm4GTA5eZvjnyokUgYi1RUfB6cUep4dkzPEslnjHphEQNb5o
74q2nuwReN/D92YyEShgFQl7nXxNkP8hTP93roBmZVzPCkfYPeosEHAZxSLfOLl6
0kGybFQeLtUM0L1KNCs7hNTWHDNYLzx/9HuUMVW5eFjPVaR/d6a8y0GJIdy2s4p0
3A6Pe60eR5Dt6YOr4oPAvST6GbsvE7TRMT5HEvP8B99oX2FADLgXJeY/tRCCEAVG
c724ox8vOtlzD4lrjls0v94tRb0S+hOzLl9lTdQBAxa+zJjEHtD/xKp4vzWq7/Qu
FSg2EQjiMfh4nXsaRQQOff2tLX25WwJJleHIVzbAMcEZSM/Xsr4M1NiP0hyLRqOP
yLjjCsOA4vt/SeV7bNZyGAampYtPhtGGIWf3Fe3t1Xh9fFa0ncwxWQZ1tF0Y0jow
3CmBFrIMoJstSCLyy44CyGckFXTa8K6ZNPAaNOoWB9TF90AoZqT3N+NI5kjPw9Qm
HUyTI6KKzOjfoKAArWRMLFQyob0f1cLdujzs2UdHHi/gv8QvMGzcp4/bHI+ZQd4k
HShEibq03O1PUPwyJg0/4qFarlfA5Jw2IdI01JJmOdftcholCPicNmE/XkhsXF0G
2GK0Si/buGS0It2bPaY4rgbFwXxo8vat9IiVV8er68rYrimCRBBDYHGNxXmBfwhN
1MNykJpQfOEH8oFDGaGZu6r67b+X5YxZPUTLLJNbTDEBsg0RHi9WlqQjpAGWufDz
uCZg1ezhfrAJl2FO9bzAQae/lKi2+ICjWfDikY2uOx7sseY0PKxKatg3zjCPipa/
Sw8xM0StWBH6nFz+n820z27wRwuPlC+jSlw7q6ThQZHZB+oZoR4TpHQ6sC9dCFrM
zQM5Yo5CyEDBlwVGWcltspTVkp70HZEh00Lt12BsYl6hppYxkcOkeT7OSFBx5LA2
3fwNIhGxs1wjBvhW7H635c42AFMYKbaT2Q/6U9krsYZpUIeNk6QGmk0Idfy8po+I
yIN7IFcmALPkRkkt+EXyoYyuobntIw5UxEzcl419d22/3ORdgDnDE1cRLaHTE9r3
U5KJA/8cIJ71eklzBGxqKtsC0k9SfaYSIzRpFUCMkUBN+fgLKcv3R5wkxS5DZpO/
ASwxWt7BDI+UKnutmhk9Gr6zECAQjSCE/QZZ/vZzg3bbj5LpF7z9UVd4QzUpGEVw
2KsUHjn/gckRMwX2fZ6wx3kGSL4yKS1Xx4Da/+JlOj/Mt+s+dcH497My4+EDkQy8
pdQIXkAfx7w39aQkE7nfTHVvyAGBEguq6BubJOncuJudU1GWZmbsTD8nVYqqfrfb
Bj1ignBsGEtDs5QLBCX9/vlJltmGyXRI9fCr1TC7abtTiZSPh8eHAulXZTpqxrGw
P++EUynFkJ3N7ZGsBLU1cDS/UAleDEYEeK/O/tSD1pxe06pTwkApDRf81w7197Ti
wdGaQF6Ul9UnOaHm7du5oZyO5guuKUdIbh5zQxM1w+kpLb7IAG4JdKmDCmjv9qrF
8KBMzf8BL3h+IqmKpwzhXKpNd2ocUIH85YLZiVWrPIptdW9UlfRineTurUQQmQZL
WMsdNQ+4aMerXAECkPSe4e/cxJPWofn4lVmBejh/xt/1xW3Oz11b2D2QEv81hFHB
grsfCWE6ADvtGSWP+zJpq8CXSi5TdJR7nMYCjv8JDFTb83xvVKn3BDcbQ4PRc2vA
aFunhi8EKPGAThw2zpUhgZfFPf/AjksqXkNceAnI9yMFKM8dyLgOCnirQn7ZYpaH
n7QUMopY5UcpdXy2d5N9MR5cn4ztgQ/7FJWDuLpeB7xUPWDZjWEGK67fICc3QNHZ
RSnWgm2lcgmgwoBnVFDCYlovqUpsJ4pJdrDSgG5JkFBJpjXEy8ZfiWCIgQtmFHla
e8Gq7+I9Jbd0m0AJXYhv9ttFFFD3E/DDHg8kwYGhPn9L2aFsX1KnuRcSNT35rEd8
vUKc+QiDcPRbBRsLm/mLDwTqvDV6GYuigH36QkVjsk4G+UI9Sro/HqsFfWBWWUuA
RlVxSfrYoe7sjZ0rKdplEPyMSrqw3jTTFWFLvvOYH/XbyGtxLZhy4fZfmLDt/KYi
h60rKAJzm7UNDhYEGf8FM4iazKRCUIAgr6o9gLkaMOB3pWeVFC1GJBWRNBYH7ebm
tjAYY9E0HXMg5eRYoG3k6PjOSlUzOCWqHFLFqmrQ2VIUoVFYhMN5/jtS/gh49g13
cSg3xpBzIzQ+A9w6m+XlGGl3Rn/eRgDj0LF8RSTHabBFLy80N0tvzdXuQHLs7yum
myxWt637HMGpN4TmgOSiBw13B6KHLdFQwUpNjW0+taymNJBNn6DByYyNt+OSFxNO
0wzSnH5mQoi3wEawRe4aOj1lrtWcucUjnUe93fbZEU6P8GdvUuyEs/rBLh3eV2F6
0+MbYu34hNRBItp2XIfvLq4RdDH6LX465453K4KfFcY5Nxe+N+pYkfwX9zSImiEn
RGnSvdagtsNMDQd9mXrY6+8+tftlTINAiUK9+nLs4AMPVpyDJ712UZLcQJpCCM+y
UdAaFBY5Q6p0QLtCBjdOPl2fSuOwYVf5J+eQTZ0XOqYrbZ/jiJ2BID80eLJMN64R
7h2RhhQoBf7uH7e8rBRS/MS+ngOTUeBYvMQKQzoRLodg1gNNAZISEKPkd2VUy4Rk
ruH7Z/VRckMAoLDaeC6SXiFcTuAPRs4AL1SI3UTNwWF9VsQhCJz74v8usH0Hoqze
B/VoZlk0ic3f3gB8QPzwhLJx637KSsIN4bSamg3Jed3fjkmiXGqnTGyr6B4Vx56W
yC3pfTYTH+SGCdCcTIYV4h4suAutNjHfQdJbIvzLQAru1ElD5L7QZXyKOpTjfKj5
TUbFcnzWdY5TfdG0dTqea5TtHJYCkewUX1DFhLxWpUxI22WvoZ+AQHHh85OYw02E
UC+sN4hDGQukwOjCeRgjOiwqSzZKF+9Mtyr5km0OoSecZsohyIPFKlhRFJ8G6/WK
ppD/ALg4FYW8LVNuHERTJp7NM++CxF0zO4fGMQo+0nDqgvNhrZDoU0GBu55+PDYP
AIn7LB/SnhXLlh+Yx6GmJ7gW/S6lwsRREFkxho9RnyBk1T6NUnrpqyudq1vtgdXz
nIxqfcejaWnyu1wYj6knGrqDSg7RCHN+IRs7ISMyvB+E/O1mbRVZh+1+QD4/nCgH
N+Z2e5XY7/Q3LEg6WkYvFoau48Ks4K7btPTRND9rabrzqlaSOtvNXbG2nb7Mz955
qqobuWc0hn1zrQbv+rn6lgUlKuLBupLRxRR9R2r0En9yhUkSmreuYdutwzjRD849
++eIcfW0AkCcXcwsowGuMq9k/JnoCr4z5vxXYbCOYBWm9nJIl+S+Dt4LxoikW9+5
AvCw9Wax6YpJO1q8OZIEBvFLG4hbRBxviwcQ31j6Jq/45bT3nI/gxq657bcNh0LW
z0Seiz8YRNiiRKtO7su8326W30tNPaEi9w28zhiK2M0lwUDZRwSAWaitm5/hyUt+
U25DlHQeo9knPYOVyAFAw28cMefsgoSmLKKbknhyhQS8FJUelGV1uSN114GMflwb
nf5lSXkHcTZwSAoz/Af1V0rzWoKemgGQo/DKqsQbL27NYG6yPz+tPb579iw8YpzO
cwIwj7Mi1korBZxpY6yo3bPgLNWthkDhxhC5EENb6htiQtK1L5fsS7QC9tFhM/Lo
eXAe03f/2sL6VsEjDce70MhC9TBLlP8OVlrp2l8KrQhEJlpL1EfUsr9Sf5No1SxF
M8CnFLY1PrX+tm1y3YUjYN4WOvLu3Y6hiJ6pJzrFh5eKO0v0nnuKrBYAbQgPyQ1/
CVfrZUZGCML7B0ou1QjkL7b53ixC47167Z0MyTPfb605Qh5KRinf7vMWSSOjchLl
njIGcoUfBMQFkfIHgVAf1hD6/Wnwupr8weS8pmr8A6bvo9aLV+wZoGYQe/aBWkOR
a0/TTyFVh+qHWlQySF/9Ar2QevCSU1tDCAMBl1mMGp+RegPqgbdmRwhtzMwwd1iV
WBqjgjTDfFaSV62Rrj/LMC7fAnje5jeg8YBmcUHVQMX8dvLX5V6qx8XCsTzgKEBY
auegG6qGy/0GPAQP0v0KMQDYRtEKRKf5UcgMQ6Xq7trnHHHdZaoXiKL6fq0YV9Y3
xTlM1VBznPZkOUt6Tzm19lMskDRoIM79Gx7Srpw0iJB9c+IUoCzPxvBdBdvmpsOH
SQCO/gfA3Bqb1STjcaNQfuDaYzuGoYHvDFvpwfhDG52cJNqLukarnUz7GMOcGs9f
gcdRJYzBontMtuuRLAFM/Q5HNABq9yXaEj8u2zOnAfZOBOFuF8FroqtSYziTza7f
9hXDnEnpwdqLXbL4JXO7V19iz4QRNXv/4IonWxq/Q+RbmZzcBj5fhJh00knVIiH2
MH2sU+7z6kvzUnjJElv5knbkPB9t5SiNrG7qESK+0lXHwha36Uwsv4z/1BDA/JzL
xfIBF2jPPCGzU9B+RnIn1f9cPuT+qxoxJU4eSXhTUacdV1RBPuCTKFMQ5ro9IGDg
90lieaB7+xcTKoxGvtqCfA7g7I0ERII4OQh2g2Hf/hrul00d3xkoqoQ1l9ENi2Ic
r4ZlH7HVRjyxukxgIUWuaIMindcZEFac2boT3b6gmVU3i+DRq+Bzg1GH43ksuGtE
anhX/yq95hp8mv+xQd+/pg2NMYee5gxWVa+aT1Y1TJ7GobhM7tJKY8loyUJ0+z2o
OmOisbBOEUI0ZYkKKKaMhxyPI4Ull05baza3fzsSneTCnkYHywycrLzkZacRHdJf
5X6LrgD7yjrT2UFzYbXzROJfpeRJE5TjU3DdXfl3FlMuqoMrMKVDlLGNdNCiMbtc
IEnopVc5gyns4yniTSd0rps+GfIwQCX0VDhbzdX2VsLDksX4XFlALK+QxJTw10QQ
1LhDMIIFWAAvp9GrKkd98bIDHREYJ2Sc3jt8wUY/UlzkewXxt+So8nHhG+sFs2W+
bdhrrCtzjWYTmJpokFewjrZz0Menu/mUWixF+0cfw4kc27hju8rH/dpN6CJGahpu
VP2za8eibexPWxjiRNw4pE49hhckzavD13Pjz+cGfHvrzlKbAy6fCgXuneF8hL1K
2bS2hh4fg2ae4VJWoCRi7Zw8UR0O+DxnVzRbZAAiLXEUBlQzBM3RbETRes+yxPY5
WSbZa1FFmuW8COWMENnmCSLWTLKw8MNCEPOYRMnHlZCWELVie/SBWkHRNdvWrHjc
hysVQvbyB3jXGkCJmp4b0OBSL7qFeRb/sx/mla/tBjncptuxWNyd3bWSQPLV5Tgh
UsD9fjy5u2dTyJIYekIkgP0ZPJZHJwKNuuBWKGwZ+DjZn8CJjk/XaLcdp5ntW9I0
Bn2nc6K1I523sMGMI3iZbyDZEtabwaH3lXEzTj6ypdVswZUKhV4Gdv9tqxpp+4c/
KzZvVdpTeGfdomAJu14XXX8/kTsz6u6SRgdarudluh65F973mmlMCvPcCcQ2/+zB
payxK0nXm6e9JIlHc5FZ6nBbyt9jD/12WmtUWuX1KDsBGZE9gkXvbZ4B4RuZ3ytD
v+6fD9KOJdoiA3dtFrYca4iRnn0h5h91UOp+NX1hFc2pWbtw+b58335hmSAAVqF6
szOdEhXHFxBfDh2hdt30EbGCJHemlp8llJgjin6IMBYFQeXR/L20DfV3OtAx/SvP
pAiLPKdJdNV4aP2yvBb8+YdSYosIEtRzAuWPferVCw9B5AwK4bJaDfEx2wD4HMwJ
7WeBuRDEmHQTQfF7l6LSBN96j1VSUkL7t/6b+dfjz1C0aq6oV/Az4FY+NZeTHLP8
rW5t+/2QjZecU6Wu3cULuAknwfaSWdMnLfYZ76zjC1183OXnnzauNnDxK/MyqNr3
duOCAKhQJ9gE5VrsL7BdDX6xC8YvWCfCUot5EQbbfvCWbJmIwx6M6Dsx6vd/IEhl
bPcJysZTtIi7xgxjKkTlbrB/S9pm8tt3ZEgJXYgIoTM5D6ZcFkhYVwQreGrFa5uL
rnijQnfBjx69sXLC6reEkTmlGC0MSZNNme4CxpiIs2hQsamxHZpnCeLAdYOTPlkZ
3L2csaUUZvKkXsOvpHwq+m/OBdaVmHvG3WkzIWVdRCMqS1BZg/5++MD+f97gHE/K
4x5L8cv2wDHLPeZk6+Cu1V0vtKrX0FEVaJ7HsIbEcgh09sd29B5ssOFpOBNGkRFa
AGtd3LweWOynxxCoiXpiod+ncmp18AdDl8qZ6Ae+kpwqUgj6Pw8YteM02ZAqfJJA
wdTRUfNgHPiSqlEleQsCOSSUPlI5bII22cB/LUIU3vN0yWtnErfpfxnqygDEswmP
gVz9h7B5mSIDSU4E7nb1XpKWG6IMKep2GRJB3cWgCQTd+p/Ps+XtZzK37KndG10S
lEF6Zc47aKaR8kLzuHLkxVqZEArS/WhVhVlESu0ow3LHIimSpfTlsbiprkF0c3O2
aBfuZ2qxLGWAO/D9DoSh0YLkFv7GeBGaR/epoRxL9oZ1gY+PSC//Zt0y++d1vC+o
5S4d1+b9dMOYyHg/1HX72IAkoLAtDshag2SO7fU5E6qbaEmNqqdp6vHdEjcX82KY
LWEIZOrV9mGix4iMC7QhJzVb0qbiS4V1DfJxzdBTVwRtXJ5X5FbY85E6xLIGpJ3z
1KjyghRGNkvdIQ3iTTnJKFPioEC1uNGtQW/jxlgjMN8VYXCUVJ3oIPhDU94EC+iV
pfOJJyCNW6ozmVYWjk/C3NTfJxhZezLtQRsgY0iWBlCCexAACbvMcAwhB+E1Zc7e
bZnpzU+TEeww+nUm+FjfHdW5jXK52oMv7wcmeYIynpDoOrWJ7EY5H5TKGmNOqhnq
/M+Q4wYWN4TXsFuXGRHu7YcazaX3pFSVlD44B3ZClIFgW/0VGK+r7cH1cGRF3XbQ
yCG0yIyHyoygoqIQt6664LMFMMdDxdBfBLJvwFDZ6hk4iBse58Un3KHhmPYhQEfh
0Guw4n+UMHqrGATe5Y4pEo2wHMmhn5b0z4yk0/0TjB1CZBq1/KYTI8+D22mVkgyp
2Scj6QC5jU1ZwLdZrkf0lfSHNf7bsU3+rOK7Q1ryGu0oYCyf+SM8sN4zLubLn4fH
ZorE9AGNHff/KAEfP+ilWMc3kw/yWtFGssjr2a+7nqx/B5enXx3iGG/i4jTESnrK
HZsDfbrrWs02IShpqVfDw3Qdd/s3sS+1JsXtuYVj8/hmLOzPgNGeRQO+c9SBbZRv
rWUNiFP9wihmLA3HaBVP5Ad2RW/F5DkV3BF3fWvJp2NUky2A6GluJ4dBobgXilfX
RBYjfDAL66aMELKXRexo+40xnGp/SQXVAdT4vQ7ZvbezFry8bgJvivBN2uwKfvqF
Aze4BFyHktftodUbwUCiC4iJ8RY0Uew0NmDQ3hLRvZ6ZTlnr45VM4OuhSgoHEcFP
y0iz7AQowaIOOJCLvdZi1W+WF1z+wQJoebvCLNeyZ0BKK7DtxJ6n+OPKHROhlemy
A7xMCc10yQfHvlFVeHFWA8mzrPrjcIBXaEFbUdtqlsc0UvtUBvmeAX4jub5Ybwcq
nVPmX2dV7T3z/1kxJMDVaSWSxRoPEYhsxIGhUYihAEAm7OBcIbHv1jgEmW+q/XSp
F1ROvydXMMFXFmlqoZIvlndP4nkbpCmDcuWGIS6rm/pe0dfCQt7tFYZNCsw1FyBq
6WamQjgUS4Txyb2mAaXhtMiFN3G6omcXFYYWJFfpLmKYvHxbbMGt9qmrHzKvCQPH
Z+hZ6SVd/E0frWZfoTRc2dyPq/766NWa/rLVRld2qqut33MwhV7eeXOS6wIoRGaG
9C9AT6VWAChfzxAUs5fUot6rpVn0t2GU66cpl59AzuznozNfXCxCn1U3riscsHKk
KXWOmvXGQfltxSmfgkyly/MvpKjlPH6RS+mS8le+gFyG6UYN28OQwRx5RLXSOsRs
+KRDmoc9NaGg7dJ/Iu3Sq1q+lpHNzhRBODQcF0muuuIbq7Nhnwxfm0Qqr6oa/ZF+
xZABAfysBftWGkwNvVgf9kYbIbPy+7CuNdjvo1lmIL1MwR6R36e6WkCTBXIkr+41
Wok+QIDaFIXO4zlwHbk4jpj7zY5+QQlBbpswbeRc7HQP/eRn4fG+WtH7kTNSeOat
dPiv/kUIRPeSYxZWnUnCVaOHLHGg+ecRGpvTxkMKHUyBk5LqVdjntRKq0AA1y/Vj
/E8r0jhBZ03/EP4fCPqIryHa0qBDhQO5a010wf3Mco2NZt81F+vbbuF8yC/scvvh
Sp2sw7CqEythPhvUyuibO9L/x3GgXzDOP1HHRCHJ3VzhFOd637byMR3r2RLGqLYP
74Z3gKDZn6+RhMUBD7U3qjMPH/mxbyuXQRhQ8GK2hZP2TvDjLyzJvlIbRhPZpfDl
IOCxzSokCrEpC/VT2GvIHT0VXOjcvAMlrq5KZEKRZWG1mlwn/1/b+2V6wLv3KHTg
RiTvaPWQ+m09nqmhji8erDaZezKGPQjoh3TT7P5emQ9OSeSx/zKJELmfKsKQFNTk
N2rCTWyIZmen4l2lopjprynHMmxger8f//xKfzpeJMQ42xNEodBFAwtC+fUxtHXE
se5yvxu9Hc6HlliwrJ2Fee5YmjqWYo19kRyZEAf7NhzSjs2D0iJR0KFBOhu/Gk6f
gAFNJCheRgkxIdUd4MF9HXRQfmJUya6cSWtQUtIMg6my/lSpj0VliAuFTFritEHc
+2WxJmYRoelsjI0SsMPXv1PEPO3aForyOEkhEU/KgTZs2GWdLvvBPEzJU6PHt15o
YNrlGS+mgS64qk6ndEo9eCARxD7dWy7r+GkoN6Qk/g6yoo/VQNlBZrDxUalea1fh
mu0UfwxaQ/tOCkhLuU68/jATMzRa92xCvIy5kzI+FfItkqYsn4O2KO833ryW+D5t
J+NuFhY2bQcgcg0wvz1QdmboPyAjpmrY2mNzGQDExFcox9VIkcIJGRXqM2FqhPzl
eRMiA7NFHyzNxyJfaCHCMkr/GFrUw/njqGLXkWAff9Xw+U18potBP6+2Chc/xPLQ
zdAt/x+CBWCnxRLRoNquO7LRQnptkMNgpVsiL6K84tvX+eIR97yIvD5nyip7d+Mj
3sAGTRkv9C3Q/zHBY6NC22u4xWZmHW4FVplwmGebC8WNvjq2yH5x4C+9Pf0jE3H0
328BkpC/jpn3xA9cR6LlkvLYwh4t+iMuAJpi2N/85r/3o+UMW30JNezxynE8pGuY
ii2Y5tbrxoD8YgfhyhOkfrM2uaRlNm9aY9gsQGC+65sq3jfsgDOmZNdFVXdtCmEf
Z6eeiTTUNGIOll5EsZOAZ3rMetWhOMcKpCQwE4yguKSW7I5eLsnZFgnGll9XP1rI
izVaDWlampOicZcdG/gZBpmJHYWQUJ7kWIR8IGIyVUSMH9rIYe7DQpYI+IqaZHb7
lcdW2J1sYdF9D6SShLVhLbhsNu9c+Uotmuzim+0vH2iMoh7PpzjNUqwcuMr4SKPL
nd6lqnkQN3BQ4AbmoaoO65eUkwSjKMlwM7SUms8+hRCw639Dpg4yU+/ao3IRn1Yx
jrEXuethBPhrEfZUYztwdWr+VbdzQqLeDXqL9bT+aRfKt2H8k1kgz7AR+ysuMcXL
52y/e011gOhJFO7z1b3pF+kt+k4AExFr2ADmhy1N4i5sQB/4LoqY/J6448LJTSMb
2Kmj4pMNHDJE6UR1bOg/KQce7ooMpQHS07gJBEqvkxpRZLTytUJnykYX+pvp6IlC
tc5CwutcbZYEduGmsP8cklQJWTHcYt2IkIinRG4IAwKy1NWeGCwkF0384H03Nuim
lRT8gYrgv96WLo62MAVT1T+LP05EL38JAitRa5V5cqCbqm5FwpMCS+WF/PmSFq7w
YV3ZUr/mKR5qOjHorRFtyOcYLw/5T+N5G2eHV6zyKIayqZYK1YfBuAqD/l4GzCM5
SFc/FbFG3Qu9rdWRDLMJ2/rTQx6IJRLffVbYCYVAymPppOW7YxgRXqg1wWkQ+Kld
qQNVGDNXWmiId7aJrQXxoGsJU7KAiF0ReVmjOfYE2W9fOB+4vLRm3wQieZmCgmmD
tiOqBL5g9cgdtByqSVwm4vJnlgxxQiOQuVpZhybRnQlF2kx6Tc90VBMeacxyQbRw
pggFO/iLzwPiKt6G0CThvMrfuwPfl0zYbbbQnDkxh5lzpOSVvwQ1ZJwmvVIWqhYg
rS6VkFiJmpeTEv3XIbKH+zygljcfVlbGHbHqzGnKn4jVaDwNRmAQwSRozvy0dWBs
CRif8XwFKsDsAPV7Wny11Qib+A4gByvCVmCBC91WhuE0rRmjLDmmSO6Li5PP3yFF
LiwJdFP2pxUyWouGFfXZgETntX0GcqnO+nBW+zlFaAvgzqus3ch5iXeEtK8pV1uR
r+hKRw0DPJ9eyP1AqYNihaosWjdFCiMt56HOp1g8SQgVNOeJG48A+YRn9MkQBO+Y
Jk2HhJ7bImE8Ddjg3446sWHSg8UbTbVapGktWtxcnCghouJxj5BlM0cO1zKCVXkM
ENVO2uhjzxjtiSmUYAQdLlqoT/P78ChbYu9foHUfYtbBctxXfUFmzc8hhnxKaPw5
AdDpU2vAQPbPCpp4qbzXo8DYjGJZQvgHOBRK7YoAwrx3fspTbPauae+ufRb2pdYI
OOWKfcA5DQtskj9eUAlIC8nArijJY1t4PS2Fgw8XcldjgPCxRS5jA9wOkZG5kqTs
qrznvk4HHpbI5wR85OtJkGRODNzNPJ34JgkWJyVf/TpWb97Rfwov9YjCy90NqKwG
9OYrB+p+4L8u4TF3w+AVxS2/PPfs1AobwBZzoxaNqgupUqvJL+gLVLZczoO3jkPy
1dDM+rUNYgyQYYyUgORTg15k21Cit22ayCUxRCZkcSa/iI0hCO1x+BWeA1OAXsAi
H/2jh45sLr5ilcNjEf15yYV1y63RKEaHOLG2oqUUzzJSDn2+bmZ87mbHfHIBVy3C
dnZRskf5K8pe/NFSGhbhGNHh7k1+osREkfmE4vYAj4PH77KgMhrymDnhE6ZqOGff
40VqvPghT1Vf4WTY8Gt0OzLNtT29o6YaDQmicqb3uTZZFcctjWgVd7vMs8RVS8Qb
Y2y1LR1HLR63OwcLG2DvKGbCBAZliqHzVH6hlAb4r6Y9vZr0j1f2lzJsXNnHpZVU
edspxrJcnwOcRCuhcE0UvSkEU0VrjFF4SH9HrkLSGgLStWPsEJtca+8yhdI/h8yF
X+CBZgColMKGm5R/bAX52qTMabIeOHfZ1vJDgctPaOOPJtS8t5XbhgpO7vsIGEEp
BWns1AC+2fbMjpgJ5nCv/j1pTD4JJojCw7599hOuu9uu9j/bWCIpwroRvJDxS775
N9akAuoLHR5z8pwf/6tccrvxoj6mFk7EqiS1B566DCoUccyZGGlaCCn2N7S285ks
Fen4+lBYcqXS855luj9/86b/VE4Hi4B8m6mnMMoZj0nQZP6FNO2mHqtbvQTLoz3d
JzGQAFjXQlza04D1iR0IvsYEPb4MSfek0DDv5xH/E5FPfYozTyK8mEiLNNOS4zwX
ZvmaNabOsXnZpQEHCSmROjKEjBX/tKtizL/nHZERc+SzbNV6VA/vuLsBUOj+0N4R
c25Pc+DLqeHGrv+6Kywh2qeBVsknK07F6LjlWeqqmP94mMCT/8lkaVooR1fzLeDI
IOPm/PQ/5Zh/vAZBJRrhVCibZhq/0ZyZFWAcqFGiJapS9lLEAcPPjpqjk02/B7y4
6CuazV4lczNcY/BQAF4wMFMoKvuXZ4D/0nv/74TPVSM9LktwyGL1NQ+5/aGOwhhk
+pL61LwvQQcj9BkCC/U7J5FqG/LfnSCpKjNWBc2giNkfucZ6YbYjVE2O89q2ROzT
fricRsl4rGlwGi8VPEAWyShb8aJz3ng2DhXXYnE8eqqzKraWZcucLgaBNSG1kEli
+Tbm9hZ239Goqg3PrBEffKB/nCrHHiUqiFaH+XgASLhfnYQE2IXwv8OLe9ycVN+E
Y+uBiP55M/BJzLr9WXUGrnB5gMRKTBFeL7FdnYY8KTJxrcy3ahEXGNfAwfZvXtUR
3pg2/fFgyXSEyIeSCOA9ju9kCQuaiUvQwVa2wagnUg0ZpYcOKKcHxHqn6+cpeE8n
GwtlGnNKrTCMrXs6C0oDGDho9gLl2vg2bz+bwEy0f0vJJp2mEjiDynRjotOxAlU0
HELkQF2uBOWC96gCufVMBcKvKuFo61dK5eoV0JDT14tujPuxI1VTicYuHDmfcQ9V
1JvCpmclRcg676WnOHifuEnuA4bEzSDlQrdJyRSii/EIin989rx2W+SxaMoKwUlz
E5oMjSZYEYF47AKcV+o7cdau/rE2OuKMtv807keDts/Isy0p2SPrcdCtr8itKRlO
TFj2JyVzVGKNdOM8DLnOdR6VovOGiQLYU3fsULUr+wzp2WFx0qItmAIzNgHkrc09
hsfgDAylYc11J7JGmVSKLxHzncm394TYd4NPgJTfAqxvFNWN/jWl/tDwTbB0tm2b
R9Pu8FDwhb/LGmty85+MH5OCXRD2VxVSjPGhKvyoq25w56Ryaxm7NBet6w61upwx
yd1vUOy8sUlp+2n0pRVy4MSgNyF2ctyffuYWlnRVzvD6klyufkb7GpbcYpnfhc9P
2zvkY61f0Qmhw1dLB14iXTEM8SLRziR14NJuP/rXNf2c/6Uu6iRsYNuqc5B/XPI9
CF5zQgh6M0DTFZnp1+PdVfkLfkJbXBn6WM16py+t3AAeXZdkULdejSXp7NZ2Dm8I
3vfRMUhaQEGOHOOn3PIiJSjBTSOa22Hw+B2ZSOAaYtNuiLSVTWjM1BXEQjdmTIoA
EXhO1OD8AGOuq7wzY8V22g7NxlQ2bnPG7k6/7x9qP7vXQoGoh31O9L235ypZ66cG
CQF4TtABJcjGhnB5/nscCaTp67E1LKVAABEbJXfIhuqdRNi+uBkjY4rHRVoQE25d
p2ONiR8swjmsmuQPVO3FR37WT528kTHaqIdWV8TMqQ9XgvMTkXPPFRp1pbP1UMSl
7KEyPN8uZ6VjIbWAKjuDs1q2/EVwx3eGIxOhPNOicik3pf7UBY5s5khe1+QOw4hX
Vv02OjnBZIeN1eH8ESNOMpy0V2pm7A2y1NI/v+b/HFL5LcgNDAie5cBmco035mbs
oAAUlgtQ1BiDz7WzjtH3Ikwr48rWEr2mhVqq2tkeQfp88yDwrVWDeWBIV/Ts2W4K
hBtrie7CpN51UXoz/frVSS4n/7jxFPsryFbPpMVOlCbhZo9A0jopJwiJ5PVcOVaV
6VQ1+MJnUS2mVWEeR0+tdImbJNJi8ChVu2xtEENvzFC7yaSpiVzaR1d2Q0csfY5j
w6rRdEuy3q1aBhslnyoYNWDyoFMgl/Sltlwvm/RHUOVbUFfjBVFR4HY7jT4sd5ZN
mSmjnV4mSoJssEL/3Y9uUDRKH3mdCYWe78+SAEEcZ/seaqZSVCu8KaXA3XtY3Tum
S6k0ZoJVRMMp8kbyVtUQKtxbrhtGxeZvfxt8nv1Scu1C3Gg7O7FhLWNPwGdHGbVY
79lgvMls9Qfl3nuVbV6LNaOD3HbE1WkL7edvj+c3NBzEjsyXaGKTcvbYF/sPp7HS
YjcyPZFfR39nH4m4xWZuDPz9kyP3YhJ+SjKnxzJo6UY/TPdrG2HQdyGgUbJhfxHF
7Sy5si4l1HVNgoQgzkCFdpQeAb/fZMA9v2ZSZBmiQtlP/UFhJ/0xARC1KZWs4hiM
T8Xtq/uHwrOFAmwBN7Spkdo4QyaW7prJNSezsF+rt6e81pDCFvnSTd+zFgKmB+cg
2FEEM73WL6odCaUkoWaBU3cNVhkeAH0NV0e/lswpjMqA/2s/C9WUMkQ1cy31ZHDb
/iHi+loA+K+NcrnIPgQ3dxpAZTVFRnbwQ1kns3nHRzdgICYOwfaWD+h7Zk4VchNq
HZsaiZd2957MEDC1SU9yeKQtVic6DH0Qu03X+1UojOC04ubASv1edlgDVcHaXSqy
f3cODXWqcMpLArqmi44SbcWCXptD9MHAWcTQY50brLs/ORBkvzf3G3yWhlYKBnlv
SGdhAbsEfbdnBtRsGZZU6rTfLPlc8g6rcZbuQ2ltztqXhKz1b8JGoMr/quyVzYSk
vO8k7ArMRf1TcbiB71Z+xMArGaLKN8zkiry5C52yTbT88nwxveXmV9gIQJP4haVK
XysKV7MRjpBjqiOWS0s5oLhE0YHZxi+JpUI1jy3jDGBLzuOZKyrVV9Fe1g3BXoc7
rmNQpbKmJ/QAGx3yy0PjfONFpr9FjFzX9U8K4GYPc/xvTf4irYF6Oj8OYVMKddY5
jTLiidVo3Kp0hl204OdqCzwjdeLj/L0GCHNj3VmsU0c2HH+Amp6pGMzAhsUDmpVA
pDW1Ajl97R6JdreeN5vCL97Fn+oWaPWffhP0uRKKDZU6fuZ33a11kDLYBLDuaaCu
/WfTv+VZ2xEg6Fenl1nhLLFqz9Sp1lgJEyglxLNQ8Qh53zVKvG90ytkUP5GIf7Im
mE74ky5cX0FuUxVUjfC2tbyDGCUz0E2FmqXVheKrCkz8U/DahbH/O4ByjiuvtnxK
nyXXASsgDLSkglaJrD7ZC03u2izWSl9NnvQ7eMw6gglPs8FP+n3qz51JSVOENA4o
ENv8ZM5Why6wxiseeqbAe16h7CepA8RmapvcU57rI3htdsc/nKd/iZ4xShA0UVTN
+IO+WVW6+bPl/IFOM6H8AumvA4RkYYmHyIjhQyWeF3klOyA05WOwr1KktVWDNLPW
aD3iTB7j+9Z/6sFwW8/Chro5SOiz1eseMrVaOMEFt4mzVzUQJHd4PMSFOmt6gC6A
UBzRzhV7IRvwbZLQoggMfb9G6GLqYzACkDuHI8JzK9ByUVh/PRl7GZGQIFNh21NN
7tJybmfN6Nr59LhZ2/WUtGPfeHQ2J3J6w46jSVkdKeloydP0rpY2dZzoD4FPm3jA
kYeI5//KRsQupVxlmrTafYgsAuqkvpWdJw6k9Mkie8X1JKR+nNbZKzvE9LWyLwlo
IA4X2nfCU1FUIRy5qV+2FbXCyACKLdE65WmuusGoAmPk4wXzNPV2tB+g7+abG2pf
68lvEmeqWvn71IvUFvry9NwBDM7pI6W2hV59SgDGtRCQNTjYLvRgGQI0roeVp/gT
MYB3BgTChRXEWTNdKsvPUJRDQT7U0bg+mvEC+dfv2SPq640eqCSmup7vI2EMrZWs
zSBI3Dyio0Zt6IRTeqxtRYA8gY7fW+/xAotSqu+m4CB0+fbjeolNFDjfGTJP9ZcJ
+lWv54jldH1Tsa2AcU+K82tnfUm1lVswzxtSxKxpP/X9CakotkN+LFYJ9cgA/uQv
7N3N9ClpPULeIVgM+Vnja2qLI2eMdOSh+mspxJ7sGBz0NBl8hsg8SwVlHE/xK3VP
7pqztyFXZ6vCSnz8bFRQ+S/PKJ+TXlFbhiGW5QTh4ACktECUG+rMMSWok3hmkO5m
8WhGSLI+XnAGkVlL1kz3IwAL16smsh/j8e/KyiIGH1cL9iBtoysG52HaZthmy7ao
5E7sEl+vkYdgJoq0XireLuRP8HndzJMiJIVUekkgroDdud8XdHK/ZD7R/tTNmJdo
6ZZ83ESxAeSsY9sOTJtHie/hb9B3a1evRkmhSDw2T6xnOjyGXJOAMe+wZrmuvfVI
9wbEjo93txyQjR168IsmXNtXPF2fF/LIs6gaiM1iuzF6eS0DxdEHoNTLDBlVhezz
7jbvTXDUz7I9syL2KnZxqqMD88DtDmW9R3Nt4GOwZTvaxNhgzmannjkEVFUGlq1m
VbiM7jlkjcHLMssIMZQJ9gyi2IaLgj6QU8c0LTHDAo7lJYxB0zv7Fgzv2pfNNHw+
ANK75J2ClICmRvVUdE0XItEJivWfmhoohpQrGNgqL1Qj2edgoZC9rUMi2PO6DBgR
H+D8iJGsxDuDRWR8C3i6ccLPdBCoyR01cxDhHHr18E+nvs0ReDUdlLBSjVfrKcV3
7K/nZmZWUkoIoCVfsKismJVGJyki7waP771nYv70sHegDPDDBHtVsEiesmVoAbWl
n/lPM23WK9nK4bFXDVAbI6cNsWsZIipmf+ZwadE4RjQCq2+hvUNMOstT9A+Na/2B
8xaiburrNqfnsrkKI5c3l+DEm5nY7WkDXMMwYSqIDBIGgFy8htb0GZNIcCSzZNep
yCiHPVsq5DuRjvlGD26lfrME5C9yn16F9zY4/YpGiLUKlwg6aX5hOshaaG/RNnym
GqEMnvUNjrSLAxSqvpyiaFacsmbnSlItvSisnqcEhmZLkY1LcmiD9C0ZjjXfsuqK
CG4Ek3WuNilllfA1r4rv92dX37l6v9qvwxquPjVJcQVLunry62kbgHxxX4A7Qwii
cni9dw2dEgzx36tWjqzYd1pU66U/GM7Upk5GublF5IGdNjvDkACzlYLwyKNqAkam
efjrQlG8e0fpugs+PiLE4L3bsiQK6oVUDT/zLezCN65gPnMF94DTphH1jxRlBuDl
jona5RH7Qk05BxFBDLt4xmKwmm1w15gxlxEEpCpTRPc9zei0i6YH+hfEETxPZmLF
4bKpQ5bigbUYYXYFUgN0Q6JlCmTZQOJFDpTEhi22V5wr9KfQVGlXa1xxBMEv0oDV
`pragma protect end_protected
