module pll2 (
		output wire  locked,   //  locked.export
		output wire  outclk_0, // outclk0.clk
		input  wire  refclk,   //  refclk.clk
		input  wire  rst       //   reset.reset
	);
endmodule

