////////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2012  Bluespec, Inc.  ALL RIGHTS RESERVED.
// $Revision$
// $Date$
////////////////////////////////////////////////////////////////////////////////
//  Filename      : XilinxDDR3.bsv
//  Description   : 
////////////////////////////////////////////////////////////////////////////////
package XilinxDDR3;

// Notes :

////////////////////////////////////////////////////////////////////////////////
/// Imports
////////////////////////////////////////////////////////////////////////////////
import DDR3                ::*;
import XilinxB2000TDDR3    ::*;
import XilinxDNV7F2ADDR3   ::*;
import XilinxVC707DDR3     ::*;
import XilinxVC709DDR3     ::*;
import XilinxDN10GK7LLDDR3 ::*;
import XilinxKC705DDR3     ::*;
import XilinxML605DDR3     ::*;

////////////////////////////////////////////////////////////////////////////////
/// Exports
////////////////////////////////////////////////////////////////////////////////
export DDR3                ::*;
export XilinxB2000TDDR3    ::*;
export XilinxDNV7F2ADDR3   ::*;
export XilinxVC707DDR3     ::*;
export XilinxVC709DDR3     ::*;
export XilinxDN10GK7LLDDR3 ::*;
export XilinxKC705DDR3     ::*;
export XilinxML605DDR3     ::*;

endpackage: XilinxDDR3

