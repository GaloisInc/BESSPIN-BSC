// Copyright (c) 2012 Bluespec, Inc.  All rights reserved.
// $Revision$
// $Date$

package Math;

import Complex::*;
import FixedPoint::*;
import NumberTypes::*;
import Divide::*;
import SquareRoot::*;
import FloatingPoint::*;

endpackage
