// Copyright (c) 2007--2009 Bluespec, Inc.  All rights reserved.
// $Revision$
// $Date$

package TLM;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

import TLMCBusAdapter::*;
import TLMDefines::*;
import TLMRam::*;
import TLMReadWriteRam::*;
import TLMReduce::*;
import TLMUtils::*;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

export TLMCBusAdapter::*;
export TLMDefines::*;
export TLMRam::*;
export TLMReadWriteRam::*;
export TLMReduce::*;
export TLMUtils::*;

endpackage
