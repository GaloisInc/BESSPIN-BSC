////////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2008 - 2009  Bluespec, Inc.   ALL RIGHTS RESERVED.
// $Revision$
// $Date$
////////////////////////////////////////////////////////////////////////////////
//  Filename      : XilinxUtils.bsv
//  Description   : Xilinx evaluation board utilities
////////////////////////////////////////////////////////////////////////////////
package XilinxUtils;

////////////////////////////////////////////////////////////////////////////////
/// Imports
////////////////////////////////////////////////////////////////////////////////
import DIPSwitch        ::*;
import ButtonController ::*;
import LEDController    ::*;
import LCDController    ::*;
import DVIController    ::*;
import GPIOController   ::*;
import HDMIController   ::*;

////////////////////////////////////////////////////////////////////////////////
/// Exports
////////////////////////////////////////////////////////////////////////////////
export DIPSwitch        ::*;
export ButtonController ::*;
export LEDController    ::*;
export LCDController    ::*;
export DVIController    ::*;
export GPIOController   ::*;
export HDMIController   ::*;

endpackage: XilinxUtils
