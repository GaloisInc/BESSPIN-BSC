// Copyright (c) 2013 Bluespec, Inc.  All rights reserved.
// $Revision$
// $Date$

package Xactors;

import XactorsDefines :: *;
import XactorsCommon :: *;

import XactorsAhb   :: *;
import XactorsApb   :: *;
import XactorsAxi   :: *;
import XactorsAxi4  :: *;
import XactorsAxi4L :: *;
import XactorsFlow  :: *;

export XactorsDefines :: *;
export XactorsAhb   :: *;
export XactorsApb   :: *;
export XactorsAxi   :: *;
export XactorsAxi4  :: *;
export XactorsAxi4L :: *;
export XactorsFlow  :: *;


import XactorsAhbSceMi :: *;
import XactorsApbSceMi :: *;
import XactorsAxiSceMi :: *;
import XactorsAxi4SceMi :: *;
import XactorsAxi4LSceMi :: *;

export XactorsAhbSceMi :: *;
export XactorsApbSceMi :: *;
export XactorsAxiSceMi :: *;
export XactorsAxi4SceMi :: *;
export XactorsAxi4LSceMi :: *;

endpackage
