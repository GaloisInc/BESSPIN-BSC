// Copyright 2009-2010 Bluespec, Inc.  All rights reserved.
// $Revision$
// $Date$

package DDR2;

import DDR2Types::*;
import DDR2FakeBurst::*;
import ML507_DDR2::*;
import ML507_mig_33_wrapper::*;

export DDR2Types::*;
export DDR2FakeBurst::*;
export ML507_DDR2::*;
export ML507_mig_33_wrapper::*;

endpackage
