////////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2008 - 2009  Bluespec, Inc.   ALL RIGHTS RESERVED.
// $Revision$
// $Date$
////////////////////////////////////////////////////////////////////////////////
//  Filename      : Altera.bsv
//  Description   : Altera specific libraries
////////////////////////////////////////////////////////////////////////////////
package Altera;

// Notes :

////////////////////////////////////////////////////////////////////////////////
/// Imports
////////////////////////////////////////////////////////////////////////////////
import AlteraCells       ::*;

////////////////////////////////////////////////////////////////////////////////
/// Exports
////////////////////////////////////////////////////////////////////////////////
export AlteraCells       ::*;

endpackage: Altera
