////////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2008 - 2009  Bluespec, Inc.   ALL RIGHTS RESERVED.
// $Revision$
// $Date$
////////////////////////////////////////////////////////////////////////////////
//  Filename      : Dini.bsv
//  Description   : Dini board specific libraries
////////////////////////////////////////////////////////////////////////////////
package Dini;

// Notes :

////////////////////////////////////////////////////////////////////////////////
/// Imports
////////////////////////////////////////////////////////////////////////////////
import DiniPCIE   :: *;
import DiniRS232  :: *;
import DiniSODIMM :: *;
import Dini7002   :: *;
import Dini7006   :: *;
import Dini7406   :: *;

////////////////////////////////////////////////////////////////////////////////
/// Exports
////////////////////////////////////////////////////////////////////////////////
export DiniPCIE   :: *;
export DiniRS232  :: *;
export DiniSODIMM :: *;
export Dini7002   :: *;
export Dini7006   :: *;
export Dini7406   :: *;

endpackage: Dini
