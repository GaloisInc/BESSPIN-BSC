// Copyright 2000--2003 Bluespec, Inc.  All rights reserved.

// $Id$

package RWire ;

// The entire contents of this package have been moved to the PreludeBSV package.

endpackage

