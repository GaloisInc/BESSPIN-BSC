`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oduZ3dZfsOUYq8ffh6KfIcVZSEJbypyQ8CAq5n/AM6tgoXzPLfIWkt2pk+ofPN7m
ZpBteAtaW3AAM5kmn3KA+UHNe+52B/EweygnRhlKf6EcY+zu+LynUqSk6hQghFSb
yrhtWe836ZvulRezPpvs2Seee43TyzM6AhExiw4rN3s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4080)
+q1puak1DXybbr7ddwAtFKCRUf+/sIKSIzZcWKyfXgbyihy6Ag4va4/DMxfi5Bee
TzrRkvNmmfDBEEaVJJ4ymOu5Lof55jJEFDLYDnU2o4eh4LUJFT51E2+miSV/9CR6
sWDI6H4uTo68qWbDAoC9pJLI9Poa/Ow554s5NZXwf+sUJJOBGHnuq6FCZtXyvHgu
NnRA+ae7IkxvgGZdeSk6d6LAptn+1KPEcozhzHKVjZWfs3n1/qVFfPQrobw57dqv
yzX5c/QDVeqmMiDYLe6vHgBy/iwUJBUcMTY+xrqov6XUwFo/uXAq4ZI6KhezCb3j
l7EZDYhpCLKmd4Fy5n4dTBmDarvVeURIWjFrMU4/gDQ0E7OyaIZfQIR+ri87P361
Bqg12ClgpJkKjhPZ3NPQz/DKKqLSR5CtSB/ouipIF309oOcGQivT3nU4AVlbV9X5
3P/YCUIETzlFQvsaTOjJy5LXFfHx5nNpmqvcaxTOTDWEgIgWevPlO2GUCDj26oAm
/Pz037dkOYDsQFMxZ+5R8jLQnGgbPuTOqnij0lTSHcdpmH0bNvyWkMAENk4Avfh0
dJFozcuzWb5kQ7GC3UclBKtOvUR48ZLUBia9gsilDmfbWi/rBha22jR3+91mMmCH
UPcA0PpxIXFCY77D9yQeyAcJNwA9n1Yu4z2VoBBeQigmnmj9PPtDDVShvQULki4r
NcM1KXQ6bNLrCBNiNrX40H++M1+V1Lm2w2ee0nhn5/H3j76C58VEJ4Meywvse+0h
JzrMCVLe+lPQLz9RDb3peIlbWcSY/BUHeNA6PeVYlovC86QBAzcl2SHfUw8sJmFO
2xFJOadqBE5M+h1LohTpyQA5WxNDac6YuEXNA1UrBM1Uv2YCzzrQv992t4ZxMUKT
IRXaWbnPH/3zm+kB5xM2Y9t8PnSEykzZAmlGp3IvH77eFrrfVZAElh0UcahLh0vs
+vRW679uRn6Ti+VCvmEMJl96OVROypJBfbfYCRlaLuOr3CANwZxqxJmp3CkjUXWz
BpEyVXQmfFu6uCNdiswIH5u6wtD7NgjZCQWd2hEWRtXpkZwVaxTPp5x3xxhtQS4N
1aCC1M1faE49VPzm4yAKur6MJtNIPm+q/gf7sr4QdPQJqzWRxnP/O8bktEBmQ90P
SoBNRU2ym7oan1KDCCGqJgn67q+f2LH6V+dAec3xHHBZNawzs0SraHn2FnCWWlYa
gfaVF2lJZ9ueZGVWaslBPvBaGJQncygPyv5+RM7qL7C4oUt11l2kNiWOSu8jhjm2
mgFdhVL5lGiitasVtPIcLKd49U9ZndWKRl8UjScpitjoXH0Dl54RcPH3bt53z2Tg
0MQXwoLXup5WGjM9rExluhuZuG9x+jpJjBBzwhQYv813bTXBCc2BOHYdr/j/Gp85
h5b2TBoBtV2nrb/kP2mbOX6UEV8oWPhcQqwe0DnafsqqccteW/i44o8COan68LzY
jJ2Wt5JJEnYCH9NTyqj9BawqmH+j6cJoFpru1yr/U5AoEgjfM2GmPW7HbF0o5EMp
EqlU0D5owemgJVtYT2puA2efp4xBidtkW51y8UJa1zyyJ/9twNZ1dpEVycAJelHb
ujiDULPZmCgveXgNa01qxb1KZwBUAxvt1R0viRnIAQsJAt5qWDdE2q1ydVo0swHl
pvtqQFIu36Ybjdhl5NLApJKQpUk1++LQ/lp5v1BO1IkPXZDZmw1iyLt6QPhIGUle
DH73s4REIfEfbEF2/6V8852K+i8Gua7GgYF9bP++sMjHqDe2z6EjBggr/RNZcuM0
+WtID4frSYLulGHJLGOy4+MzmVbysF83Lqo0GX6ANolYLoaEg7GyQ+s23a3Fhtg5
kftZR5Mt6ZabFB0Z19qc18W4nS1vS8Py8wcxI6Io9v4HMxD1WUQxPDKWJLo+6bus
CIiUr/nSvTLv4w9hmkDeQ2HocOl3MAF5SAhLjSFop1AeE2GCFn4qA8LwLjcBZTY9
IVezANlwp6aDPlhavlqhp71XvVLpibCd3R3RJJoijvvtCUCxSEcoXlZKiJt7/doH
GItkbmfMiYvE0uIkLDyvQZR/N6VlahnC09FcxWq1RDh3Wtfgc8xZ5c73Ep8o/Z2Y
Pxp0xaDGk7b049B4xQSS0LoROwPn0MzNrp9bxUmQuq9YbVv68706cg/QwyDwWdNj
vydrHwB/FoqO3VqlrCuiW8jMgRKfGrfquPe7XeH6m5/LnIIK+9es3RLqWsAnZjT9
QBBOQYI00cLoYJ0ShIwo5F5FxrVzp0oWkbsN/mXMSkB+JCuHJylvDcXrpB8QKM2F
5WhMX4hTEC/RmMZCPKTlLOOamKdV2D0jhLCbsqssnXg6E3Z0IwGdwmj4RQCZydz8
O1n6ciiFQKkovaduX/sMgMTzvJ+mSLWTnsYPjjYRSsRrm8fbGfc7x2B0IBdwgCGt
ykdyR55B6D8fzRLP8Rax+K4GqMAOk++Bx9q8UCOSN7BTHdmYHCAn9CCuQyqKYKLk
Nd302R5K2B73OvE+hvNgWaDzuawqjfrXsCEVyoIIhfWDdTqBWndjqdp7aoynyQLQ
w8pae+aycFrYe70P5/u5iNw8qp4q4Znmz9ARtjq6cJFGm5o4YIdBhROnQ8k+Tnk7
mRayUYJnNHgmvUwUg4hqjV8dQJuywzLDBI0TAvxTFiCdluMvwM59317mc6Jwk8vM
Eb0b57+WwvxR1U+2b4rcC7iQzj+Il2/beU/ZHPGhWpNLXePpeoG/F7C4nS5fy97z
sfvOPeAmh3gwQczPp2VQWlR5Px8Rr0GHI7hWu8K2Jn83f06lMF/uf2+b6etmoHZT
oTON8QA9ZjyyWnZIrTDOs/jnVCgm/66UYIbQwwEsyIUZ/CkW/C+LF9odt1p7REZp
kkODj/2Rs1/rN3rAxQReQ3CGI3y9rTBi9/gP1EL4oqvRQSn+frL/4WmGvui9koIN
VzZ0Joyu47iGQF9CPv40MYdxv0LODAr3Gjb0TuW8W1MPZNzFndJ98taCf7aAMWwX
bi6YrBNLGNszkfredDf9O40tW6vV0nYqsQKglMTpzT+ty6lHYtJDGy+FfrBsth8B
FUhdVe3HnUIqohp3tQoVjtqcz7pI+EKzrUOLxv1fROrZuOrSCYOr0upNFsFBEfGM
xOE1W7Q2rrUCYSysqYzIvEYO8oTwio7/VT5lvG+J9KCkrlkG5TYnUufvqj3ZwMKo
2aEUFegzLeG1ncvA9zERjgRu0+lIrwhylte+lqMXrZNReyPv7m0SNXyZel+5+UA+
wxvY/lR4qAolEh85XJHRxxy/61e+Ij2Aui28qC2cn6S6xScHduR530FxPSkSGtf/
z/3iRsWyaCY0u572bEk88luoFQIM9WGP5a8zWB6L5ZXPcG4iar1iFrEWUBX1LGr4
e4bvW2u5cD3lftDJUZM46OxI7IFBsBDAknxyIR+mPLcyCPAQ9hT+CGWPGIFiYW3e
rLgdIccT4QZwZ6vmxUo5UAn7zpVgG6nFmVSf6WvzrHi899Kcewh4MIRIxyRJ3LH8
2C0tilFfGIMUv/6QTu5GZWA7SiPoEoFQshLCkRyznhB6I0zBjhg86Vr7v8bRrq1F
FY3tjtyHatCh57StBDx5T0rRwnqUy3/HU+a2fZH87QAhqdd5V9JtNsqslR9r1MXG
u0sQsAhNOcOL+z7I1bCzMXP3E6ajMwns4I3RTvelpn/OKwqJwoKVpE8Ew8t2Ve0M
8RotG1vX2Rb2+jJ40h3Xtb1DcU1dGpJI3qsinnPm4b1u749M5PsL0jil0UEEYc45
ez/+wf9YBao5uVMQDPM+aghEIDN5gbLLyHgDitA6ZwJCpuntCjxZ4jrRPTo6/Cpf
/YVszL+muOYraDdT3uZZFSx7HG78l6MQ1p3ucpVKvo+cLIfu3mKsk5OfcUrdNeob
kBKDlzIXbscBH9WfHk+7ZE7dgr1a5UfVz/OR4xoZWZgKnNPTcRcO2gQmkLnvcDt4
qKU4klPupNp7aegF1LzabexTpmOpBRsIz+H7LDaXWeVVUiv8mORe60oMPm9il0nC
r1tIHa4/0FiEEP2Js0O7r2PhlCSIRN6rPCHmIQw8iOnByZ1O8rZSp0KI5xs0IDVj
7RlFYpDMiEiKqTp+LQ7xmWeZNoP3IqM0hG3/Ifdj4vch3KnmD83ua65fmjlWao5v
YiNermIiI/isqRVLzNeeC08ZlwccQ39t0k22CnX/4zS95JILM9KsrUGlxatLQ3pg
3VHFat1PhL9qWmgzWtF92qdHSqmAdhhu5ukA4obhqGgWzvw3Nmj3Rzp9XTNy2iFd
JpZqghLej4ehlw+ATXQjw/bMRYKlG/xsSIsBL2DEgFSrnXZv62fWz064LAX66qIM
oeo/0fEApINF66yRmHHMH1wmyh0pKfRR1pROfoJ2GB86ECkLZEQiD8TACcZvhVJn
Mt2Y7lMO5UkNm5blkIkMx22yfCmcsm3L2WoErr3KOSXPhCqp/2CbVm29UX3ymumk
1qa7gvcRP8LjSkCUZmuQE1tKQXdViq33KUSkvhP+ldVfRM2yie6A85STJa3FUh8f
dnK89WKuaOu+q5GpNI2Gtw+fwtWLC6LRsbZQMuylrgngIP4GVK1lMdS7k6/V7OI1
0endow7Hys1ObEwpM9oB++ib/WcQSxyqahKTYLVb+bjr6SCidO2vcFeYbQzpDTlf
6rJskP60b93QCt3hiov4y+YJYVikwg6KeT4F4eOzZrbedKy1wip+3nBM+9Qs6IbP
cb5YvPwAHIgq3ldnWHgYRFdK1+o9mU9WbRdwDGjRYY6pXSPmjCHefqYCDGKyMtW4
5YimbvjGfgF8iMYbGTJiNomaa3SU1H9s5Pcc1GPiJYjiK07n9tVLn2mgIxBHIAAr
c1LSOSizxiUR3yCVh9q7ENP3/Gg7ZNlck9QfJ5Kmey2w34lBFu733SfzmGFb41Kq
cOkHkc0QOnUFzAilJj3FtEghJS1gu4QDPHSbM72b6utHMohCIZ/vr1Gp1MQ229Aw
XBNCJEDSnUIhxNri6zHWIpWmykMjduSYrt24WrdfTtNyALdA+bqgFlJZJXtf5LWT
2kw1VshjAyGLQJEJZRQXdMri+T5W6R4tkG9ZvW2LUuvgKvgOEDYCVwqhAursPczd
w8N/J2m2zuFd44i3vhhlEZ9Mq1CCO7GtHpNLPnHJ9YmImfGRgkUwqeZGglhZibDb
8AImNYnM5A52TxSduUU4l/+xcWPKcAmEFbP/L55l4z1/LVYuDAX/BLVzt7RJGEAT
dIGCm29QB0d/vdhrkEQh0YMYAhRr7PhADoSw686gPiCDYZMqLFQIB3k/Jl+HnrkV
y25bAFlnFx0dl6kQEOBGGCEa9wObAdfqo3jv02ETSeWdO7F4c7K5545iXY6omFA3
fkpLqqu6ory93fDw4UytpHyuYULYKeZ1NYMCbMjjk7ycFFmV4GQVq02yfXZtzppV
`pragma protect end_protected
