`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
K7d1/dsetrW/25dxr/DYJwMXi4I3RBN2GUZeq8uYtJulfTcYT8ronVZr+clVQpqQ
Jco1G/qDD/HfdLkC7z9DrxFgMHhJaG8X0Eg7jqw/21Enhzb9Dw2UhHXXeVzTym5V
l1rVzwntUJyXFbCFCiqyMgCEmpxQfxjj/SCFEt0jLf8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 70480)
WQi7xdDfiAJzwaJTYv8n5WpD4Hie/sH9PnaImt2EvoqcdC1Im4ZlccttK2Z59meO
AviU68YutX7C7ncjGrbxwUTIZoQXa13c9I7MLWOPweEcnTV+UKLYC4iQdqlaHKDS
xjRkTV1IYoSjiwEib9bWBILFWP7e1XbuD7+Hqna1b/b6MOTJkFvG6P1YzrLKgSW0
rYoYTJKk1cXxCYorCty2/pmg9LR8mc4g2fPWxjEmDexAgXf1+86qvOfEsd1piDXa
jGSD3+2Us7HaQ5sUhVBe8JdXEPUFTaifX2c8fNVQ7tJgmT/02QZAgqhoz1T+ES23
V10tuLfR/mk6ExA8HlRlpyvUfSFQFSuVwhqvJzjRCL2ybZFf3vZZzxCrc57Ey+2v
TD8WQmSLWpfFEoqDGihJ62OJ2UYaUw4SIFWeUsTDx3/JYSGsErPT/ECAk9Eb5RMH
BZ22CNjVT14C9qpqgjrD31dYKctWRELHW+wUzXZ7HpzhrjyF5/+7+G3qDYgSxpoz
rY8fqx7rD/PrkWp16/CcxD1c/YopkpT+aT518GcLrbdCEVFVH/TD/Vqa7OuPbFag
TSBYsHLOWBWvyrZPs2eWkW5T1gemFdQRQlTw6zqtkrjzSwYJpkP6Xs2uruFrHBOF
Wv0tALy3XUw6inzI48yt66hWWxXGmqNmGrlfa5rlBUA4s2dZH2IFmXcgQ2G/FqSz
zB9NCap3iQKmhF9OFSbKHSd5Cm+h8w81GqJGolK9kVggFso0BA1d3vhLNkkU3Xzf
x4zviv+76aj47Sp+YXUbjbYmMmeQdRoiw2xNReNoYsyzorBreATtTJ3VX8WqldQh
Q2Twwmv9eS4Ib5qkJdGcDSj4GNKXQCBMmzLPgwsYZuzA8VUFu3bzMiaP9EPGRbh+
bUs+gk4PJcrvM3348HztZICjOHo6DAf9Mmy2ZjRCrvtfVC3r122xhAYkwDfQ6mDo
LcfCTLsIq2ll3Cp6TIOwWDCnhWQOUJDsSiwuYutCQxwyWjO9ZwHWfoxp31j13gSr
mq8PxfMGe83IPpZM8alFjNj27ET0CSMK/Bsp1yBV69SrvC/IuczaqxZp13jngsYy
6SNevlH5L2ue6UBHAEaQT+JrvVF9VEH+3RoKx5RRe6cU30gl/J7lVPcUz6bK3475
7DN8Cd1SPJqUS9bVaTzksLA/qxYWGpv0yugr/7+2pBRRdsST8GCaXjaCp8HhLeG5
w4pKygsVsrwB3c0ML8rLyYEDABmqqQuuDizgUkEVXpvOVP0gjAJMUD5mSGRTvpPp
YXnXJ3In7nDgd3IhGdcUW/MKW/n6kTLVz8k5QGQtb+ZMvZr+iiJ8UdgeS3rsomh0
edzgHXfaemhJSAxKkdSs0/Qdod8/TCXAlvqTZaXOdtCiGJXENbc7mzYXGQcjTOXL
0G4+woRf0TeXicwnjsTJ+ZmDAIfM9+eczeOZOl1IyXZqJU5V2iIlpSRQAmYB5dhn
9q2g5L8n+Q5gXqO+y6qRXQD9588qnSP+6niY3t/4DaB3xFZ+crysjhic58+AmMLA
3zXL58cg1O3pWjllP4WHQnyNJE/54Dv1wkRunqE6mxTOXUiP5Byxwg8doUarHawP
muxc5VLAGuraw8rzD8ppPwg/yQyN5gqAsZwdlbGQKysK/pceoGnXOJbQmAL6F6zO
badF7dEsS7LIOuOuPHSTDf281laM9nz8g3RdXwRgA+WP6zw34lOiuBRYcUfLCUFw
bontPWwAagBjfg0OGFA8G9xQyshgExI7fgK2zTtRHGlUjEK3U7ruM31t2UB7T+l6
wh36D4iXsxbbYxf2WDXTk2QYB1nb8CdK5OSN4tH4xCkudgqDNgUekIngFAXMeUjw
zxHoi5vQkZ2LOUe18hAiOMFWI9g0AicOap64+V4KptUinpjiuXc3xFbjPVUuJJ4w
viR2mq28UjfgEx6uCJkxVKeJewOrKRZSPn/FnDHLCLy2L7baefLexYZ3HHr8Wvtw
ob7k53OO7BP4bZxAzD0TdXWymQPILmPsCwQs1lY9DUnI3CkYuE2zqxRLoO+eqaqJ
nw9fMOkf9SRdhqTP/upD5Fe4eoLbKuStzl0++AB0eWm7UfmUBMY2NSeL/06MNXSX
ICWLTv34X8cjXt/XuiEjlCZW7f/HONOjghOPZpbH3m28zyNVHVVWDwx2EzK23+lS
HS1BA9+RUDXpvPeM0vJf4TshJJqWUvPsEMGnfDxjd6ABMk9LTDrnykuh2DwVddN+
6K6GYvKUg0nrVY1zFpCPW47Dzrvq3JMfpJkJEy5lshC3YBH2qR9F3IuzkVevCoeS
EW12BtBCvO9CRNC3Xq5l+Vsz4xyclu+u8TXWDT6gmMS3J/oITmBERohZnfjUqgmS
mRimAro/O8of1VOy5KCRY/Jeera9ysChAgQrQrNYB/s87nuNAVbMWwmapVIYwDAn
pRD/UtTb+p8+2g6Vk8yj0ykIJgwFtKxR7IkDI0jirbmYToJZdhBYBZXl/j0u9ink
jiMg2H3X9DvsNlQccmGtus6pKCJb1LGzXw4nZSvQIkwD+5gc3Kf1Jb6hHEv8J58J
LYtdl3nHAFQWoKGEgIRiZ4PebKn9glb8BZ8Ed2kQqRTcLHMyrenTNLiqO66pQaRu
D9FqQ2AL8kPtDTl1RWaANh6O7E5oM0Kegk718aFSt5ePWPsnHRdhJezCsIuHsxmR
cRe7YCO+o0xUDAtnh3cPMIoLAzf1QBc3LLgzTYvt5a9JML8CP5xwJuk8GCYzSiMQ
5+rJ+ZOSf720WZXMuMrmClsGP60ezqm1SaDLt8pZoNvABcYJfuTnnua787lssKgi
6Bvj0yD/5+hvQKzovSHKlE2+PCyLfZt9mDSbm/8HPJip03a/OKgNmHoWF86n4gAC
EnPtflh937LEowamyuD2Vxxo8ve9Pp5eFatVuli7FvjHW5CY+K08XoMtEDzcGrsC
9B9ALf89HbkSwbR7JXdgjdAgatVmps/Ac5erUfAn26I0LlaAGKFQSNW2im6I+YpF
KE58LY5t1OaJ0j+UzIO6SsT+v/uw17QxKip4Mejb2DjmZgNi7Mb8TbxMzp6OHLPH
Gtzolu+AhfKqeuwyxdpcTr+x4z8qhx7H2/3KoxG62MsNr7LBmNoWmvGTyqLmpNxv
hhHncjKx7ulXyl1vSgV/4ab6j6PXKqS8Dj3k2DzFxXMqGsFRHkJrNu9fwlWa8va9
VHi7SA+JguWkKLEE7LCbLMviNDsRxGCajsVDP9iy3tlhwnld+RZPPb1mJ0jHdACC
PdojhqHZYqYTBXkDdF4I2tlGVko6t1zbm/BfkPHNSJ8Lill/YVZCVxi8oXJ07p9k
f7roJsj8/1ErD1Btwi+7wg6ECy/465PF5MPtulfB2qE1tK+lu/XJwbpv3RZZjUcH
DMnmnTSuoPJ5V0SfZz5Ok0V3cE1Rj/EM//RHQ8Y7elo7unIjN3QvdJRAseK2pOzb
RHTwuoDcXAqRUJxvAu3XNix4Uupcqsz3kpeMxI5UfKacDWKDPSnoDCInz+VDBfnr
siahMjEy7bKjmE4Gq4Wf5US9ruWt2A/54boTmRi3+niDrp2tSAYG3k3VmIRhCHUy
nms5PrNBOX1o+Afzju8cZ/VoJcpGTG9Z0EigraPIE3alOfhlUE7WxJYKRMI5j9gf
c0hvo7AGGfScJiwP26b3jiHJfsXk9DZoAlYihyk6GVm4lJdKKtpd/Pze3aO2J2MJ
CQbXdAHN+UYj0OxJ50lNGG7SkKt74KkVqna+lp33HK1Oq23x6zCQKHmmIq3cjaBc
prCmhmdpuZFfPS6oAOMWLGkRQlpGs8PKbtxjOpOmVjpAZSUq0TFiWx8wI5FxRFue
7pQmHrLhyS6VS5i1KKpvovhIzRUAxy6X1SfA8CHLoPmEVv9sw81JUAhQJhCBUvvq
MgoFjpCeu1k2M/gJu3NNlfc+j/kRD1EUjrsmuOKuV3BOtTgvxyOfGdoc11p39j5/
5dXsdJlVb07KCEWrfcuoO/EYgqUddzZQp80iJuykwwQRiNRptFBSsVy93e9VTQX/
Nsj2N6jQgKLdQP4b98+0b9XdDEytM8QJeEcBxPZ5uQEoDRPMYmKpX9FgiEnqmcUe
DzAM1ex04AdnOmAv/CTNSjrv7yHmjrGWszcmzyRKlCjSdypJE0opYWkOwGtfEkYW
6OWWuUUkuBOCeBRNSYPnv0AB9d0lTDtPt+Eu4DR7/YNm1isCY6H1Lf2blunqFOju
4iQSThsea2I5cImXW12GGM8UnRJdDYsfWO+5RbLg1bt3Qz+DWt2JHu4Neq6etFis
g8BjHzL7Y5x9nJOju+MYHJupHO7gSeIVlj6BepUssTxRvx+zImZV6dRd95n/wu9l
FB00wnKlVtNojzigfTTxzYVnk4QgkWxb+vKlNIZqDuaraCjpP2JOZqvSXhp4xPAj
c76LANnehWzCBQqUzlEj2oFMjuHEH8ZJdvNnQ7586Zsys467OZCqae3g/R0o+dGQ
pdByqJHqqQ8xxCyQrKJwRPt7xxRwiJI59dLfikqASEOk4GqH4woW6jziZEz0SrHN
kgiP2gnPmfcvsNPHb7focO+YexzQTPcpNc4NYq1BG+Ia67zFezMSK5oyjOCtTfbz
ZI964C8oDpoZqSKhYCGK6tMaSgfd0UPdcBOAab8y2J3tLoqUgd4qgKdRedKWY0CE
/ot8z8oVhxSanqfAEmXE8Uu59QhE+ZEIE25yiJZjmau049eOQxX+l6zNOxVeNS66
GRslPrEbcDuAph50qorELsUZQZ7VXk9GN/P3eV49FUFNZzAoUPyeddduTXTF1ev1
VaJ63BXRs/xUgJwLAH//IPSKAz/U+/734bw0pE2Th2MlG4elENFE3PPOI6ETF5HS
L/MwUpw+Ac5jmQ3uQqq9Rzs8lbHaerU5V9xgGPvKFjHXWm8DXnlGtqWxdsgbMtwt
DtZZBy+j7OnqFCUhrHzF6A/Cjdrc8uUtINJhohfaGcH6SKfPv1q/vuTT6Ohi2S2j
xIbZh3PBfPywVf7rhShFhZzJLpfnOVT9ypKd0DP0kuwl4jnD9Dbf9oT+MaOAnYwq
C9jQp1p9s3Okz6QB3H79YyXvKkoBGshKDMs0PMnIR6PHyHt5lTjtJLMGj+xDuJQT
Dpl2PC1Hmsa+dqq3OcT94tsrYjU+Kw+LpxvVvDKgUq5hG8M/pUD3UH+GpoYuuNGR
aMyZhQ6fhSZmtNNIFln/0KK/EjDK9AXQ+UUy6mp0B4lPjQLroqlboME/Ck6GcIYZ
VFBrkgu1LQuyd6iphygwiSKJ8HSveqIfJeDAr2b2n4KVZlq3kC62SbFirHd3AQ22
vyOcYAGCKL7X1Pkak98pMPeZf1ChD06B6zzsuJM/ZWzlyvgjrPRR9wOUkwmvhzBq
IhFWBpNsxgtlPZ7XTNgA0fpYMxlQQmL1kvbg26/Sh2w+yYdyBRzOV1iThf85PKTH
UMJQmNPVKYAASLJoBRIwmLArx5xKAskpdiE4w5uhLLTeUAKGOvM72WrtSO5xE1PW
uHbWhb7Niv80yfF+BoLJZOdmISZSaUVOWFqHw7+3EQ3LrvXf96KZ2Vx/U1r39KQr
+2nQqh6dob+L3eIbTSsmyk1pNDWwGm3R7wwpAPy87g1VPis9XPSBRgDLRqj+Xyuj
ynbhVMyCHjaEolyQEcUViEImEd0ved1xANF8sWnWYneXY40wP5XrVqKZaiJIj2gF
uZOdrEQQtxK/pZl6g8HleopGBzM5Y/QQAi7Q1Ub8qxZ9OnKCaagL9xhB4J4yaL9k
Kb15d/PVl9285xqTCsNh/pLWdYTbHAIwfeIkQNvE29ZbKhik1RoF6vxVhwZoqDJi
NUT23dWOpJMyyVYLFdMYChcmRqj6deHqepGZwhZQiOridpjempkru9bFZkGT23r5
lKNn96KzirFqsiuOUX1tS+AL/jMkvsZq7MMtGGDSfEi7ggQlD/cJXCe/5y7kHufJ
8e5b9Erxy1vqn4bcNBlonOuAOtAUQxxANpPvXousTKMe72XOfJ1LG9Uj2sHggoht
+4FCggcXpIoHkvMly3EIaVVScDNJyjDQEAAkFORp9KJOwdVWqNBIiGSVMlwJuLIb
stXGEyjQ8c/yVHBN/LBsDuwPQBMoxQc7Q8kC2LBRh0RAIYMJPvyllQLTnyqWfYFx
IAOdrgpo9m3/U/CheMLmCGvwKLCw8+PT2XilM/KwyqO3wlG9bvueRJhrjxuDECWL
nHhtDJ6Y2idUBT3ZSZYA1cB2ntuZ40BhJmN22Cc5sES8k8rUFOSCJfsGjdKXVUGu
ScQhI7/i2GRj50CDjtJs0yi01tCOIWJ24mHG65KYMB3WNp7GdwhcfetoR90Q/bUD
7cqrPB9fqH1Ub0iK+rTLZS+xzfcIMiRoHia6b+ZGriqVRTMx3ppqX7ByeEwuW5kv
E+4XBUA56X03iUDJyexsOo1XwZ1Vj41olNADAJKP4Ac9MSo/OHjDlmi0lP2IlJwx
dQG+ElLyAB/DO+tysDQqT9Nuv3FvlosUzoWnPxne5FnR+91VHRZgdoOLhcodfFlx
wxVRo/n7rxMhWjYfC67gYz+G+09cCp+2aHYrRylhlbcgelDCY63VxUPG+1JVVQmp
afbjsTc65sIQNoRCOOfaPOWtkmx9VV5hyWPKXqmQqDiyYBWWWvjJnNKBKVYu7GYI
PLcQeoZmNAX1Sj1AJvvjMRdAlf397lgq1XQIZmAiRWiGqxV0HvEwVBqRljk+5+ud
4uuXd0XFk9Ue5y4y1pVRsiyaKKGuHZmytX3ESg2WT87vNit0NlWpp1AXIU2bL446
jmr8k/c/OtPWrKedHNrrfEEdSaPMUgHO3ut/liMNJMfzUGMTflwvWB0zMXAine1E
BD3bsg+7XwDcZORHT5qO7dsFYO1yHwzM7VBgjQWlqgvosphUZbQFm1or7n0fAeFH
3I6eUqEWvn6qYph2kFqyVp739arjH0rXT89c7+43QEgYjCRF04mFSXOf+acAXuuC
ahk/sUZMOURoO0lre80YXdMrnL9OqI7VVoK3g3pZEbbTVBxAtt4Ret3ZbgI5+9gy
j7avXmTbHskbXQg4+yH14REm0p+47rPt/LmDoVDnG0ftap6hQC2mWAAqBRKjiqpZ
vANTmUiI1T58S8ppF9EbuMYSZYGXLPP9+CCKbA17T6id2U20HSToHE8QJ7mY5HP4
jkeka0nbA3zWEUH6F/Rj3nlXJC0+tVvl74V4uSfCXmXH8thN1r2pIiMZqTiHsJB+
CZlqPBhdabHDz9KzmZLylzUc0rL/dGWk0nk0pl/B/4mvpb8jsURgylTlsWVq4kGf
9tEWVqZ4MnvaB5J6nv3DzfDIEj1qTWf7BhgWHNT92XoyfF47cY25XLsFnfUJt1of
udUj5WJtSR5rkZfw+xAMlZ2Leqlw7IYx5siBY+9IuuEsVDkhbqjzQG5GD5Goza/P
T9d8LKXWKVnnQeHqAWtvZWoiusrB9040A/Dd7M2o+WpLEqhntAkqM5ygE1TxgJyI
k7103kAA5I7WYfwv59E/Uobf9Bp//usQe5u1azGJxuLuRNTtO8eA6PLHhXOIGiAt
5z/9PWly3+95WJuK0/KcxmW6YQZsz4TieoQCzeI++QC4TYDbURHNPmFROPkHs+vU
e/Y7GlvaNIhieRqdChMqONiLbP+RoFLwtd2BxB411bOXe1hlSv3qUHd9G/YcMzIR
M7+J/0dxSzrt2f9zadH9KI0Kr6i2i2KuCtOu2ttbwRX55CqA4jvsZg2fwz30H43+
juPg2EHH0B4A7BmJx+UFG/eOs/L5EuglPQdV8ymb39wj7zULiPRP9Qps1n8exb6y
G0t376WnMGk5AtAjVHFBnczxbZRb7eUqPbacfE4qr6PyEy7tn5uhb9eyAAir5hoH
Qo0Li28YJehh1pqHaqen5+Rhf+581Wp/Qd757Lwis6x/xA5LrgJ03Uq1iN6ck6T6
YrbaEeJiVPdBHkwhFoYAkBbJHwxti9tbMLxAf9KULABQgD0IO/pMq3tucpnryzRM
gZb4zP7Znr6vjArhogIXlhyy1jb2QRgz2TOTIJaOkqkT2gURmvZ+29m6ojDHgeXM
Sm6/LmfnR4Go8Qmm3DO7Zg6GERlwmQxr8NBMaspYIZSJDPWmRPBFyb6D6ZrlV5Pr
fwUQNZFoWUlXuKE0qSjm7mbZ0JoQnhwX9U0NN+wPqKbgqOqZDXf3KTl+5kSiqdF5
4yBM3NjvBUZwZTO9WfsjoHfrPTs8f9wYwLAL85peLAh2V/X/VurhfGrc7kDFCYqM
FPrOox8er0J+7K8e89mn64lBoRdawLJVDKXjp6oBHbLxJgonfoLsNnwZOmFFveRc
qg+HLpctEW9/3+R61TMNnz5rAlAh60vA1cvO86aompNgWiyZ51mQbsHFfRbZWUAk
iN58WJpWrVYrvp1lWsHjD4YxE2rBv8URxtuRAVPoVM7K4hEzqou2glWFntGQWEkc
yTWNLvTCqV3dLdJZwQehWWLwcLLpnK7W9izAt8UB+8pbK8uodHR4xH34XRTqB66p
9AbQTraQmrF8aYgLn29cPX1uGnL8YjOW20q2oRhCBaI8HBDCRmwKMFyIArO0+DXZ
ROTLIZR7vDm6p94fvwsw4hg0wBY1kSObQT50k6RFGIuFPQ8WG81obCJWGtaiW9aK
1KmC1LD9YBxgpui4W7snMBed0zTQENe1jTqM2rC0F8ckl6j91yfmjW0jawc0z137
QpMwieht9U2AZk7pU1olMNWZzTwj2Toa+F4JeyiBe2mspIWjLjWwYNEbUgwpFDhL
gwwEw9JNlS0nCkrsj+eXACEqgg0NwLdktmb4aBZFkA+byI3MQH7IJonpxDIHBarm
33esVol0CWExSSNi6EYJ5y8ToT/3eCdxdW/VLA9E4l9QZi4vm7DecdT2NuA8oHCp
XruvZo/E0CMT6yKEoMMkYqk0z+8l+0rIY0RqOgLx3ndys6G96PA9E0IQmucE3AXh
7YqNpdRPffy9z0GQY5uUWLbAZr7rJ6nEwg0Kf7p7f3oR2/v5ZpyhR3tl4YR1GskQ
JKFrnlAhxASiAH/He1cphmbJfPRkMA/MYe49VPeSmXviD3/qAXiQfGryJEVa+Goj
rrzLt7X9FA6vQOawmKsJLy6UabkqqHcl9VK+DIQql5l64s8q/cCMzP5miDcWNwSC
/ih3bbVqeJq1CayV/vzCaxAAU/Z8L2RdqPPge6ufHqTIPwdGWunNeygVqaqNalsI
rXI7LcMqwNmFGlynvfU/k+NCJ8qhRksDMIEWLHtsxtPsrlTXEph+K8sCB1GP39ny
rqpI1SBFu5OJI39Sl60WP5mTYEqHePor/+11WvvFRGz0DqRh/sZzn+qPbhjuar5n
fgDRnXnaiyoiVJmOJrIKOPBjfvoCuXHbxdYieGhTWbwmP1bo8yVAqZcitS/GS0YE
rwV/tRVGyrqtk+AVLHSt4BgCsvNqZLH+4+e5fYw6M4OwNIkNqPIGWucvHXrD4q94
59wFIhWQXDIrDS4acybTWwVIClrXRMoC2r3sETB5JrUvb8CsEoGz+rd7SzRvr3rX
YUgdIdccJDhkuTLqcSR2fLwc65VR8gdZsHuWJp9Do60yZrfo2VX4Rb0IvTDaw82u
i/Kg6jbmENWSlo6p5ZiPQYtx1Mro0IhraLDfTXijVx3H+etMHf9h9Li8IsF0bgHd
JKyFyxQXpdDCBM07I6lx3aKNNupK69sqT1NVfAonpqZiG40nWArla8UJN67LdJKk
Gr+obWNzMS/lRV+5nAlzWs6AQYnF/ZbXg+HnSdGeNes5BKWh9Ba7qNzH8T2DyQiC
6ozNxoC7qyaUbeIhlN54y9AKT2FuvjYynE4LBVUvFIANR3H6QS+X89RSmYESOoEl
Wzb2K770l/t9yka2n718k/UVldQIl/Siwcu2iJE9ZwbUwLqZMiU4S/4th4La/1J6
rp0Z9GtAnQ10o+UjRG0kV0+NzhJC/Pt3J4ZoQMBuG9RE1ytrCvsWX+lO2p2+fl0R
dsXy7aQdsEI8obH34qnu53Y5A0BJYUn47dZj4jKW4OsMoBGhaB4gZ4oSUZ5JqVvu
PTkD2EvMvsW0YIERDDnv7buw+uWFgyqN9SH1tcmInDYBFSa6lA/uKZiit3AEfcp/
k68rRn4zjh7zliZKgY3VfoQdC/AsugnZ2gbxIPASC4G3M5Rb+xXmkZaFjE8CM7IT
KE0TsVuNnuBPtH9Vikv6yvnlCjCUe8JTqi7mRsCbGI2K7Ow2hBbEU9xRwJ0Gaf+I
4QwGK4XBRS5T1hVWAtX0cPk/6xjrMGdOrcf7+w4l26rJO8DwQ+eII9xw5GuMit6u
Sm2pQs4+D2USK4UO+oqHm65l/92TDYHd9VmuIy4ftsSlJCZ+zOxy8af8LCNjUgP+
5v6Jr1Am76SNtwwcMvdauaTh7Md3UhCqNlerKLtbZNrPY9uiofFREFRMhJLn8xxq
rd4EBmFldSBxe+FCxOBN981649vgN8BQOas1aORvKAQMJvDAoqAB3tmX6IE23cpF
7KdYk2k6Dsrz373uAt38JwT6jrgnQCHooN17fbDSqF1G02YpO/SfT1YKOrb//v/4
/YyBooa7b7V7EB2a024NlfHOnyvOqQ6/8CL+NffJa3ZZzfm9s1kmMuJIPlFtx8SW
jfiRfx9ubKKFIRkgKou5m0HLLpluVEJORZwQiWRgBop9ppy8ax5osOWofJPoU832
XRCZ58D417W0ErUmv4PGgHEVa3xqSz4pMRb1vFohgWfLuePB86xwHFAyNslRY+7/
i9rxPYxVFY8WR4QXAXGY3gEw2ViCghkqiIN8n9fiUGkULcDENnYuO9OxeS2K5fKb
2Y+1kHE34pwH5x30rwByYacybQL8ciGw7KRNgd9AvigxzjaMnczHMnevxv9TzudP
nzfkkJNdMTOQ5o0i/3PYvozFXlyGuo//RzImuOWcqkuddQVA5cfIPHbQJHPM1uQ+
fAzMxz+UqdkH0Vs8kovkmto36Y4Yuq8ep4WbnZGF+WnaNGxNenqNo+FZfq4gE96W
SveAEA56TFXvFujciLagPKSkx/FQX4LeQiQp6slu8foT466liGKuMTWDjbaQafKg
UxfsaHW/JkXaHMe7qsq4oGfa6V1OcekyKfy6Yjiu30lizbaRoRjyPHjo5pe7w0sG
dNoWExrjPxuKvJ+G7O7uktHBNx/mPRTpPvuyiIvGQpwQZl0/XsCfYYBny4q6zjfr
bbMjs38g5NczajCq/wWzM5srEoy+4C0ibSJaQGCa28+Tna8czXE78AlE+gnXCdIq
pFgs0u0z5TQkFRNfmMp6GZwYXGA+Gbs2gcpkeN1p9CBJ4L61BPbT94sZnI8ywld+
6sYJiIju0Ox5/dbvT8X7SGlmQxHRug74NFE/0NaTtCgyEbBVq7f1bWSep/6iGAn/
xcZmaZaFxvZlx0dGBM5e8g0geRAtAVC/myTz0iLsw0P7kFHTvvWEzekTXAonMhqk
Ttbbx7Fdt/Umuv+aCrhGa7eCtruC23qsOqCsXAz4fpi22MJDU+amF9mbH51C4xNz
hTdQlGhnx19AvvFWsDl1R9UBEImUwyAab0EkqEH1sNXy46bIQoVo+zO6ZQR4Ip2y
2FXUKxcrFoMWdUMOSuKDH9vshAqYX8HPo71UwOCh4IolFzmmEFoMyOR4RA0Vitve
oK3HwXihM5FEGipKomtIbLH3nd8IrO50q41QfR3aZBza9DKN2+1/GboF9t/Y0EQH
AbvwvoEcFj2jKbjtUtmehR2G5FeFkrUueCvVK5Hzfo+bsVAT3BfTV9RM9jeyyGgQ
9bMpjuFOm13aE4C1cpQZGsD0JTNRkU63o+UcpBCq9PYzQmPDsgEIECO9eK5flunl
S95TciKNozZac94xW42PptRuG4mCK3Dcu8g2MJ+m8jadzrNz/YqMeBPl1BJsJ7pE
f8MU3GwrWIs749rlXM8YgElFDBPTQSH87Gg8CDDinbAx8HyO27yvtG+oodpOY1mZ
opfARe0b7jqLnRblx+0Cfr1zXdGj9V38usBicqMdD1qC+LbryagB2fohdyRyIXf1
Vs0fzrUt4gX79Xy6mkHUz8XR6CwN54mlAuvPP5OkA2z3hauK+jpyEYy+lt8F0pAJ
2HQGjDtpLUHB1LQMgxTWF4PomAVIKn3maj5QDM4i+OLxEr55qw0tUQVcJI2YPWO8
j4k71pnteUS+/fb6ADfyjlUIyiD7MTn+SNptM+jUBJiXlnsAmk1Y70pi1tw+s05R
xM19qVT3rJgDPtKN2hjn8m+uzurwHalHfNoj1hT6D0krOYlJVkNQyTV/OV5BAGq8
v2lEDZj+ixIFtb85dwlMKbszdVm8Pwz3LnbMip5o3HJ/7HrN1D1QC9tDB7aKuwCj
u569nH2JO+liKvoaBCcSj7fxxkiPSs0Opz+e4OOERtRBfuOQA07jTlC6srzt19Lp
fAs/8vPn0vMtH0oM+Wgt5gC2aK8GzZ9xYDnc0xGRyvcV9LkkFLu9gNuPpYDFkLye
i1bzIfvNqAftpp5Q9N2V5RJdiMVsg88NaAfKHEcalQdibVmt+sWI/SgE/7CfzPiq
G3ikpicnVM7cKyMOrehFv9PEFH36z5WZ1TMkwDx5fkx3RCeIEjqyIZqhZEdnMUVF
W/ML+Lpfa6H8if7BChgOSYGH+knIT5FAfiA4y/35b6PGhb+/lSfQku9YoRsP3Apy
xeRGUsBGakVj9fbP82zyOsYc9LeDj7g8O2BW7/uJnSQvumd3wEdWzBIRKrSyzYBv
Aej4moZKe510V+EeZ+YAUuX5Ghj7ySZs8CKCVrCdb/tYP+eQcg1YJkmc8lOS5Ib3
6JIMRAlyWBEjKXb+knU5IlJy/CmHDKh/FvMdKYQisHWX0xyEF6tl8P732l1jf8Ru
MZ0cO1+6hjX4tfL1xgYHhrVniW78W1IBAGsAHC5BNyBnFdIrc/lgldpDVdrRGncb
3loswG2oRsna+hmRYdZIsHgv9O2294Yi81C1C5lEuEifrnJ5SghLNMCOLnoYEdlL
I1GfIDnwBoJXacDv9ID8xyhwgXU1Rb0zOF1M3sbRMG5UWNTdeJwKzCmViusgn4CJ
UwHhNtqLDYQt1yBr+KFm9GvTl8+3ms0pieTcHWDewUWctxc4vSTq9+DY73gEqTa1
lnJcCO/DKtDYQoRxmh7soJex9V/JnSPaLSS10diKpJHKFGgQu7k/B4KeQD+WvuNt
xEHUPVvR8CzxTHiQcQa3YcxKJduP44rSvSI1yv/Oao9mkgaipXv5H2NczpDZWk+4
A0MUlojk+D+G2nzvO/kOwJvzVqP6Qnd7F7SzKM55Ck14BNjELqYJ+2nwIJd6qC4D
XIczNd9JWjtIBfqEinpej40xZ74ADfud/mnc1tKNuQBmK7Ag8U+4odTKJ50ei9/h
OGUdnfGHJhTVOfMf6hga5SpNJfNivBi9mnUhB9iuwPUH51PdfgOJiuF5dlpfi8Tb
1Pz0PcIJCq8Tz9Hk7zraDhxDo0JY9LQhSMH1LDi8kCUbEvQSic9OiPfLBfN6Vd63
GI4k/CVn3qMuJWGpmZN+LJU7locA94RJZtzZDa3tWkBJYnbcUcq8QcSmDq+vNM2L
kLDf5ruXcrBX0A/lssfrNzr5KsVuIjkEF+HTmiNterTgLB6RijX0fzm0AR7n4Xa2
WBJIeRJBG9N/PELXSEamBXN02dghLws4J4EAyCbW3vpmc7WZ3FDMDbNIFrTxGzCZ
zxLAYnmqWhkfJIA/76ovKF759FQ9kw0/bJ8q1cokcAe1X0WkNHhgh6BBl1HiJRiO
sc7qZMOvyacaWOT9BnHyEJOIyA8ixliNG/qZ1DijMdDYMZctyLCF3W7//DpqWyd0
zB5A8F8twyJr58nWE2cNZvQO4JNlBsozBwEFYKrISbKwDXzUFcyVIVlKnRdwND8B
Sn6iaWUrzxuiLgzdTf1b5tTJgWT/QqkH08PY32QJpIcy2ne347IQVl3yMTAAO6Ea
YLRdZo/NBrzDvDLKgfet20VHOqRa39hEz6NukepLIlbfT/WGK+01NUuYf0QM8mXB
9scoxEk6MRvE2P9taeg9LoExrH0xvQHO9dV8q7DnXU/vMPFF2JL0MYYPLOt3Qrer
0Bqni39rnLHhvsrVu9L6gJ3P8Vy5Z6FgcX1gfTlk9QUa/g0zKRXhHGAeN+TY7tMw
w+VfI3qIf4jnrfWOIEp2r2BZlutM0HHOyPWnG7jZJ1NASAq9zYhsVtap1eumhRyT
iSBpsfF+wD1/ugUnzX3o1hEGT7ON0uiPH3RQtNw9ngRoZb4uNtvF+lqfr5CcHO6i
YMtDRdO+Z3/GHacB0jy+/PQkJh4vHPrScyIh8DlVVjJV6TTysLiUh4gFRZp04+ES
NBpAb41qJz6GUMVh6KE0mH0ZHg4ERy0HIvCcvlB+GF5ZbODHRhB6CVyelivwnccF
SkG7RgeiU0kfulPs8eWOJDg+N9/BJwOtWkS86ZYyTiBiblyVh5aeuV+PMo/azVtz
SobnN6g3TXwSWAXyOqZTQdqYWxY1ZAJ9b66nDE3IwiahSqxetFTgquuJK/SZ1MUE
zEfLPgZwsZcJ7V1rtpT5/x93U5Vcn85ttf+aIMU6s8QUM3Qp3c0B1WPXuMZa1YpQ
a2nm15gLQjypGmTue8AUkfRqPJsNikByNm6sr0O3aSy/RlTGVbHxGWDRK3tB/i4q
nrgIyTcag7kwyI4e1QbRYzMTHY9PxRpr1kkUI4yTGVToBKQj0Y+G4E4FQCP0aVVd
kmgC3nw502z0eJP4L/4Erdk5z/yLm21Xf3mTohUcVPBvpxENbQpHD0sQPj/r8wwn
pjueUU5L7ZjNc4wj30Tv0y4rQQL9P+2XbwfXncgi8d1z4JXkq9I/psNnJTFCkIh+
vXyU40e+PGQRkgYVR6oB8cN61LEQ1n3w090fCGWsgJt8WI45z70nZJrgjTC5SJ0j
YeEr3Y4AGmvaqHevq9lenbuio8fsB3+VNlcrw6uN2WuWc/Zm2lK3N3DSrLprHlIo
qG2CoUVk8QG1t1soIomMgI6cq72V1lIaJGXyTPyf9XeHk1EcH7CTZ2jLnU8NR/gH
kxPpF2s41mudFm1m+weunBYSKxBCSjJR5puidcUTbqBrvKpvLhyBJXK/lhNQHPeB
X9iei4SurZ1XCJAEWy1HFTIy3G/4E5Ysv+xq7ydnoWTJC1bamqjokEp5NRW2r6/W
otCosj1EaSkMHOwAp+vri4DlliCgb72JXRPiHeEv6fOFqnKm3MkYZWUn7ddhON3v
kOK61zb3Q09ETAvFN7wxmhuPFPbXrY2wyjyRcKuZalsC89X373d8YILX8Q/ZXllY
LEuFmB+HBuiiibD6fPx2HLZ8Y+ik+J8OyUUPSVI0ZvezIJAAbhwGLP9ggC7Tih9Z
634FD+QSajhKLBhQHNOaz5HZUSo7bGu8OiT/u2xlSvI2BDcWHRz5t4Q5YmvcKCI+
+YAiUXnXiGZORgh5qIPorXLQtf4TS/4pUlp/txMX3QPMFVWSCS0UuUoTc+jO2pvX
xMiolPkAKaKkdOyUOUqiWNOC88tYwKW9+k3OD2tFQpwa8a7KXxgrcYK+qMD5jKQ4
VDDN1RyvH+b0nnYME88cWfhHAMCwgfXDV2rE5gfYGD+XLm8WhDmpHH2aS3q2UzLb
cCHz0RSJNYpPOOsjuJBRKIJLXZGbFEL3lmBFv2fB5wIESWJtzCXAeXxoRFMZ9O60
emuSKP14isRcjS9BMz2DmAU91KLPjSPJ+y5aE5e8A+sQuJoZqu3sDkZh9uSaItlj
Gzoiigt7B09LEcyKFeBvtb5lWt5znhMqrMbz3Rmz7glQ6B7MuTClutyZxZkCGKD7
QoDyHXbX/yZFmvI7mUJoUfj9LsWyfufK2YspWXpc8t+MeQ3fOXt4py8K6t3m08ZN
EUKgkqRicF3nxXVQAsvfC9byza7dpJ+Li3EhLnxGnwIv2AcD5vQtdoZIkFwWPfR4
xKD8pHIUayOoI6cOmeaaEBS2paUZ23xgLBvkbWRtwNsgRSeRLouY+EEtql5rLzhg
/KqPPprJsiX5+vr5svqrz40oYHF31B8E7x6lxr0x3wK/xO6PaolN2Sh2Pu3xBx3B
zUZNyjaXy9D73ZA2QrV3A5ypRjY7OXFtGr5VGIKvFacrtv5pkR/ZEkioHgM8AZ9K
VWci3ZHJuagsGptCFUFY+4qDszygNUiafAkB5X4IYrZsWzok5VW4jQ60oi1xKskM
/5aCgBwf+rjcpibgbApt7tIxKFl/3G9J5NzplpEAsJEWwDk6syVOVWTdGEXOVU8I
Me+JGYTcxVAQfKizu4tf7gZxJwit10Cjv3jsbh5Ux77GSq8xm0PQatkTDy/JqeNV
ELUr+sgokO4sn9onRAgRShd4MFHz9Y6ahVJ8GF/1w8i0ENEe0YCPap51zrLzkUwW
xdrGxpbV2IxDi3pa7SIeQqvWPcAlsjdlLJR7rp8iBhRpDTdCzeZy68H9MgA+438F
A7IFygIkIkfjD0eBF9++KV5Vd0xXYi7y6MWbnZQN3hHWP22mazD7D9BJdGWZRW7U
+fkvMVZlnqa6XI2kJEUugEM6OWQQ8jhS7Soo7L9oYfKg7N90G0Dx4lNUiPEERSMA
LPQZ2uw2bwf1XwjWu8QMgODrWPQ+DND9qlueoECWAZl6BVu6HH/7iDVIDnxhkm4c
8BnVSfLjBHS5Sq2pTiTo8FJixMr8J8D9yJB0uQErqvcJBQAOF7IaJSEEje6vr4Xr
FonlVOQBSy2+LoLoh/qBxfxLk/Nl4ubWHeB6FmhTpIQZJ1mvCq+/1+8LOdiQVOJ1
K9XcLZzmMLBrXmi4d2i1NpnRAk1KPxwbfOWRsDOgZUA4ObkKdzK9gr36oiPLxnA5
REJnu6Fj4jvR15I5siDKQpJBz0BouZTD/AnjpMso6uBhtZrKYvXmaK2HI5HX/czL
zG96j6iguQsu88OiP/K0gAuIpF+1t6olbJknmX2d1Zt+djNbgQdGh/h7t8KKM4be
l4WHiuyDMwYQA73i3Eargf57v0ZzcS9a99xxHIr/367/bcOy/r0nA4vU3rJAKjeV
uNC+QsBkhGKZI/JL0Vln0AW1BKWzDWkNSHpICkaef78PKBE8MWeGktoQo3UEZiHi
9Bvf/47vjdWRIsTPsN5dDbinZplfGMZ2GYnfXSrPR/b3Bhad+/IqG4TW8a5W4MN9
26FAVHK9EfeJ7zFF2QvFMe5PaYYFC2aJC59xqzuyqyLkY0SY7VJUjZDDmPU/Tfll
OT1qxIfsCy93NjRvlJLNN6/a4yzQNtoMGdxiF0jSjMAgNmPD9WehQkiYVO1t8dDF
PyM8pXv1BnW/YiiECdotlkiI8owKYoKUAAtFLLLitjql0UBrTLkjwFGNBZJPxLiq
s1HUgGQlf8gXkQKqkbYgZEMWD7Cq1xa2KtToOsqksak/BcE2WCptEenKG+JRYRQQ
Hzxn8qJQSE+QtptsHghmhrfyPDNwfGWQ8dO8GCKMYZoaBZNU9WQuU/67Dp15AamF
AmGD+5tSe+0Fcd3MXntK6P5un4A5vruYXlGGxofswncl6Fj03TrHij74XtGlcTJv
ohkJZQWa5kuoDYs4njoD+E44a7UfcFiLFAxo1AfDk3+du7OnYtL2EZOag1ZWWBmF
f5/gLBasulnPh+ARrehBev7g/ZAAY6TVBBvwFvEY+xJjKHZdgkwYCOTORk6y9pG7
4F4+v/NodL4yALOa4J4e5rBCvbEgqhuBmbr/vMDAqR9/B9ahDHlFH7AudO9MLZ6E
7m50ZygdjeYJXcNPLmpVTBNZ8f7nx92Odrzhe4mmOuYYOdB2HmUoRurCL3XkNE+N
xEg/a/8UmNB0vDSCguRRQwNhtBSIhYBox7VQVOkC69eFZlBkeJokS27czqYCxIL3
4bMRtCGL78+g3gi27BCB4nYmesmQ8IsSBdb8n4fgMRIYWeXbdESB283afoGC6wmZ
RP7q0bCAWjwCOcDChTXBFgWcPp0GNT9k2X2xDCcnrF/DtY4OlLZKP8czrzE9ysbB
cfI46W0t6LRWB6Km3uerxYyBbNCFC340C1UF4OM3I81S4IAOydPPS/qnyiMWOTf9
67pwNcu9X+tHrmceez3TDx7AJZJhWwDPFYzsyqT7Um4qJKAkip+m+7GYJHPlVvVZ
PNRtGr9SbjKoTs5QKDiK8YirgKb4y1AAgLp3dvFEnZtzkG6LiHIBQi9OIEyHHya9
CTMMDKWzYJbZ+NsO6Bvp4kIVbibsemdQz3rocFA2QOCbwzFYjN7YAFgURLXzmA++
T9P+TNdu2QC2vgoMglsNrXwbPAoQQC+WLpGX25dNLoHEonKuCrBpNfoE6J09SAmw
UJs2+IfGRB2Hlc99xPGbY4IR1FBi5Vlh7iIq+WGMfWp2/S4WHw3Y719FkGdwGpbg
qfnwyGJ6v/NYfpH8UbM7YZrWfy4xp97wnQfUz39RVqHKdHeJreWdav5LYUxWAbgM
2jZRnGJGYeqs8ykYwWa853ePpiV6tWq482Np6pAHrCY2/uVyRm52AeDJGqE9IZbT
Cuo5oVItZpat+GJMi0QOpunfuJn8ErYnIawo0CXsivL/vGXDWt+PrCSEwVmcyTBr
sGc67hYrXoslo9sVr12x+EBmBRLry/f7A+agY4/dKhgYahxRgCWTDywb8nwkmuAS
9i9EX3dKIrGZVkIRGnWZC0L6MP3h8RdkaUPuDNTUpusWOSyQC6V8xpURyjAQqHc0
AWTvyDj8UEJpaq+QYNswBN7opQNn3hCX5r7n3xh0CATcUVIeCXlig/gYQvhUOMXy
MT6d7NknXEw9ijzNVwMjWPFpb8tkL+j3oR5R3eQpl7A3jzrnlKRfgGIyakkDlt77
GhH7EqQPWKnnDh/NYnz/TAhmuG0RI4jYWvZxA3htC5Ta1RlG8NYd3Ur4YLnivpcv
NlTIU8oIxUrDcsGWjk/bsKvk4l/+V8+yVsE2rG7vJ9+C+aqzYA/CMgVoE/46X16B
u1lrSc+psSoPFqyn5G/Unh6RgRA4+6Cz44Z9BAv5RJazahG2KYQ8HuLEPVkEVZBv
tKVTkxqutbsvs4LUC2Dq6+LrNjURLkCjFSQvAArHVHRiywtsB/FrJlGCmTjuJJEG
SnziLtflK/nkNt3RLNkmoXQ7xsCf940D5/maB2dIIbthe4oC0URtLvusQvvMrLHR
uHud5DAY2yPI3cfeRh95b2AOks1ZhUm/MEvUnili8AB25iIzCjYr8yKj5LT/Agvd
JxgFomQDbo9zkMVJDZOxTrGb4lNEsGY5itOBFYlIHqOJVQmS+0/792Qip27K60x3
K+HNv0HcxWD01QtBEkZ6IQVwMCrcRvdurY1iIedCT+p4npFVrLQ18OLf/owRwfKE
XEof3PiSgrCpuBVex+BmtvujmgiCI+yfL76v7S20ZK9oxRjD0VAIsG+bfL0iDRNQ
6dGORKMJR+vzRez+6LBuTyfp0LTKOvx+ORfNm/SQ1n7APv1wtxBIKYanEfGSYJK8
OInKEnjppHFZ+gtY1HCq6D1dZrww9vFqFZKlWchsXB9auQ5to/JTRIk954RL/3NQ
Qa9ayaU1JzNUkYYzCyChtv8BqSLZfAVcNB9SU67fHl+JxPbZlln+kUqYDSvP8XSI
BjnGPrk0US0jwpA2KoLFl3W3ytTzHA+LHiB0mhmSICM5LNGVNJ3IPjuocBYUD8Z+
DBykvh1KWnoqXCoRFHkqreN9UYFddkjVr7UfXk9GOWrr+6K3hXbd02fMQn/5SXrw
Y72YWRp3P4g342ukM7p+7PPMZZs6PRcpbpQhnC96jkeClQCkaiUYFs+nkJusgxGy
fci3TTgkXQkOtiRlkfC9JoGfKttCr8nOcyZy0UY9hY8Y3koq8eFnhFEduqSB7OVz
8ikXu6ZO5kk6+2N04atCVyprpsZQQe/+rjsszemol71XyMdKHTm/mgBG4WCE5YAq
aAFTdqODfQjZEixE3kh7TW3pM74mGdAsjQmSVtx5FiE/JfSAhn52mBrVVRT2rFKf
KKSnOA2RBpZotIYFZHxABGiYwJrR6JiyadZJjsxZJXVFdQGpjGRf577lTADCD14I
TxztoBbcg8d2Mio77UteAu0xyTzoa2AVaHxa7gYGg2ZYitXRXNhSLLB+7YOdYoe0
WG6e0vydzco7hsGc8iKIZ/JfltElz72jklYhuNQu0nUpODfg3DQOvT1JkpXa8YOe
93BMRSFq3eZDhhRM7/sUHZs3Z/FZ/0gFqdbiFuAUBaRgQCbAEePQqcHhP+hnvH9d
OiqJfJbWIsFA8kAKwhmFB1x781Z47wUKkSz5xOTJDCI9t/jPFy8eE1C8BbAQN81n
55CpgrwxKb0k1s0U2+YZJhgO9qTheaFhe/e5DXUTsiDTGFDA5z/w4DdN2SA4bYMK
oU9N87AEE4JadeKDPRQtPcNbgHd5q+ZmVbOEnuZbzmyijgBaQJcNVf8c7CVXdFqk
RBxvgeunOltYpn/AtoDBZziNFKZTSSFOZzJNi3sBMYX2OMEmPV3dJgXIt6L5J01f
sM9rdPHvR1mjqCLcJO44nbKsjrtHKQoqo3nqVGPSvm+oRCGl0lzEgwq77+b8hv1f
V2I55VuO6aZR6NXvUkLU7f1T82nmV+gOyqTH6EThkUbK9K5Aghl4WRLb8qIx2Pw5
Fk8zrzOlFDaiG2AARo3Xtp3TgtbrltlFR2qAk5d5FIFt3+lL9R5hnTSdHKX6Q1hn
aGPL0DNssrm6lhGdoDyVnsN91i2F5EwOFiaLDdY5ROgy7Mq/bzTudjRI7XYkZRvK
uBVYZ5d6B727o6bbVkEFecrqlSLNUChjBPBvoLx2+V8wEX1WQojx4m0UvCjcHD6Y
PAhxywS+IE7nDxtAZfq9rFlfHatEmNQWLTXdFrjZgFvZtnzG1PFqkjdLFc5kgQ6k
P2B4ndIhaDRmDN1ntL9z+7m5QBv/P/UEQk8gdSwWj0AfZpEjy8zbk//2HHk8NBiC
70mUzsMRPteaAfNFjwY818OpcXYZr/+8OMMdnUWMIStwYFt5khQqc0BWdBBrupIJ
Ebzng6h8sm9GKdwHu2DlyN/mKwly47CNUnhSJJE/3K4+Z7rlcbFUzQXVUbfIsi0W
N0ubwcptaQkBVM/N/OFG6M2RJUnqygzlAo0ClZ1oIIkv5j+4VcCm8A0cqkfa1g8u
ZQNrneGB49Lhstd/SHpZ+oKKtN43UPvFWS7TfJ5U0ZI8hUFrt5uaJcSxDEBiKJt4
iWne427rDn6cc7NVk9ZBpJml5JOdK0YZ/5+QkPvrUL2eKUVS+bOP7+P8JE4Nx6nj
wsMuL6zOx7RcdUxf+Q0p2rgRrqcVP6agXDvtfRhWX14l16B8lJculSGoQqP1X8uo
X3fs/e1DrooTzO/s1/ihiBiG9TGsCVHNJjFJZFXbxsC0FNLl2nS/o81bjZea52nq
y0AZ2JLSPn6ESAxegXmFQ5jEIzL2IsA8JJZgsG8yPFLkgb+ZqnwVXQa2IlihuJ4z
2wltIzavUpgt3gf/aoMIIPIjIO2RtvkKgqrHqX8XCLa6BCI5vqLkTQHxRw2Pb42q
xHq4uK7VH2ruSK8P3nytj+iazD4l8dK0k6T/nV6Waz37AnRg9PVV3j20wF3DKLtZ
O5SgGl0DGDHcjho9uSlM83jZFeHBUytV9Px5E28taNucEaf8j2DAchJ2OYb9wejn
lRda8zD6TeHymSNIMK3MEfpCB9ovm+mW5SkNfyDGsHlQisGc0yWMArBoXzJnRxaE
NW8rtRZsb68U5KMSTpJKVL3pMZjuMfoRwzN0FKu5vYEFsHOArcw+4mPMvGwQaHtg
z+dTPH5PpJW9PB07ZwYY6wGhtcHRhc7JZUnB6IxWetpiAlYPqD3PR/qxQq23Rwse
Oh7qPHlXHZzc2ejVVrJUwsAGw7mQuyEGQmABLWHt7HnIywR+2Lz9LoGivkAtBwtO
AA61PCW2fxZyirjbr0MNPdRQqF7lsUhHZ8btAZy2V60FgS3xDogR3UQ5JsI2IP+L
UZadkUIk+6JAUf2XED9Jd1oCb3y+zRYbGbHbRP0nd6x10Xa5NhtforSfjlEiMsNi
Pb8zhjRLChRH/w6QkkKm2erT/6zR+cB52t1ktVod/CgZHGlFZboIhuehYcqaKOmH
lCqHZK5O4/0M6Uwuvp9Q0vVb0lbbUXJMN15M2JxkwQCpOqvdGoDmh8w/Z2dnb4DS
DdkMI9GhB6l9Q6umQ+5foqw76TyNO/pYGuT2mxyOTM4utBSrwq/V3UaL/Vw5Ao7F
VFiBPbFuk64DlLBh4CUFDeegBBhepwvpQ+/5Htc7tlHJ6uC62QnJZzSCKAIVq0MD
qdgc16r5fmORe5eVklbF1KbTpvEKWfL3Ap2l3PK+aToqdZEwmJNpCSJD+fwKDE4f
b74vhtUd1jfTZSu5kmG+adiKao3ZRXP59Xp/PiJ/yvGwQVsI018CPaacP8k7aF+w
+mJi8Pe0SNljZqlojp9ep54+Fq/53AMAOTNu0P6h7kVgu6jXxmwWku0JMSnEvfC1
zKhRnbE2oaJQD5YlT3eP5xPRMp6oQ1TVKGNePCgwDvejsVVfmoCBX9Q5sCBxhBCP
mJepK1LfkyRnYm8tKAI2QKjSxYiSwabU8WnYzdFs71R1dqm8b07CtOh+PfrA8dRP
G2PGaf6sdMmLTcgIF35r9XV12nvL+gnH3EQKZFbjch2WY3uooiKJg9ZG0d9B1IZh
mTcB+MVSvve483eTreD1JaSucSqC6gCtGaJ+O6QqeporEnDWyFIerfdjUoW5Wwik
Ux2yyv5YRgFRi6KeYXET6wKcy0xiAVN58aDmojgJDhMCqy3619fggHb6df2kmUkS
TfZllMKi8pX4SZJhi/SIAYrqC5ccm/6ueRxzHMRRSyYd3Lw0pCNIm+1wJem1ABev
VvyfKzSMB+59QTuy9PESiNOnOemq3u/3Q0K8HqNH32EcOClntF41Yl533NiYLP9y
mvIjKkSzmfK//P3J4m4gTeAU0KAKZ0EbRJ0hcpjkaJTwOh6A7exuQoiG5oMSfpVx
DvkLoAQdmA+cOJ34NsX8p77lU5NCZNFUkd7+xSq6WgMDuE4b2kYNvp+PB1Jh5slV
wQ3kGquhc4VcSRkqQIHiQ8tcCOJhdOgmaTjSfGRAsTkqtnRhq/QPI2zBEVKkTuem
z0YWwYzty3akSal/cT3bkkEfxIbSPDvLYO2zmh+XtMUc1GaLMdrQ7KZcwxBzKijO
EW43hQY+Ce+jB4Zt+oJeZxHkgZ53z2z4DD5bOudqwN8P6tAJLpZ+R0WCC3dI9ith
KYu5ZkGYfVcL36FY5CEZfU2PO79tiQHhsyqp/wR/TaBej/ziqeW/aHiPevFmVyi5
vOIm58+v4yrcvf8t2nEhy7XZybSy3sVDWl3ITty2wdDKCuusFj+a5dyot8EADhHZ
R1MQUFX4HmK7gJGvJ22pEqUq/zF+BwmYWxtRf2FiN7su/yNOOLXgtGLiWjo7v9Ge
g0DAVwhgZcoOxAzDuOliVk+w4blnP14Pf6nyYWx4BcccAuVwItSQr64oLj9uEpnL
m0Wf1dQFFYM985SbKdw09lELhaThlrHp1LgrkAZARV2jm1d47/QMBIa/Gj/9Z6me
TCjVdjLZCe0oV7z1dmhm43E9cuSrZAcUpByddzL9jI9jWZUhfK6PWOY3HZA2jnrp
WbSvQLoVpWrj6TaCrDtFIQpp1VumA+poHYlZAvsx1lVdUOlMqsVk+O6GFPuLHs5x
EQ4o+1BX3UxTy9A44IU1YnQ2MmM2puAjbBo32o77S/Fry1uzDS2eOS05yQWgFh+7
Luxi0rEX3g7WTGFdkXPcRA9zIUQWzc/D9n2RBK3mgyr1bObFxcSM7vtJ3/mUz3jh
Fi1s1iL1is/tfzPjBoK4zhQqQQrsoTzBHf3394kc0CWeXsKHtzw/L8Lza/L1zaub
q4+d2dTotUiiu2y4sPij11oDHNAJ7zQwUXnPNH3H0Qz2BvetoZzvhhCSF9oojuHo
bodGjFrZdRc2Kdx3CFRt8GaX2hZCIgFt5MbpxRIUvUXX6UoLmL2JCSoQ8ARhl2j8
hrJsdzCCECXuJxejB+DOihSDR7ELfWXwuTqUNEn9BFZCSaTqPatcOhzpklwjUP4Z
Ivm5S3WimTscL1aJzsyjPOOpRX4ckzGkcZDRldqoJw4BDXLmzbIAveKcehv2b7MH
T2uGuwydBEAw5/D0OcNj4QHzqDeaTyddDqz1f6xONmtFt2nfmNzml8dGvgNvWkaD
sHBerxHRhnBVxxjOpsu+UQR2cRVkX0ZAUCKcj6ODA7gjRG2hSD4US4tPMpQiV/2+
A2KmtP7Cysh0cQr7QYegCcuwMz0NMO2ONgYCPaGiQTC54GBYwOPihXdI31hVUdQF
i4RvJDPFz14g1sTWKUjYWsENrZ83baCbHbp0LdqtDohXVtcpqIRo+DlJbFDWk/Bp
le4a+jvJ5lMWqtFhOtw49iJHUFOQ3a0R5gFbDdwNRQYzCNg0BrndaEQAGTDPGoAG
4xGsCVW+APqXqzi2JNGfqscHC/9MdcNWlc/eR8WFbL92YKrD2zIWh5fxqDWpaUa9
s9sdBNdD1PgqZKAIvbhxEjNAuyxLJ8lKNhTVkRNRkq0ewWzUFN/P2w6g1vIXmD/C
tjFj4Pq0OZGx08NL59CJ8uEvvNItw+IIcv1mmZ6GykLg10SRMOBh3N66vUZdvjZ5
hau4baipaBqjmJ/lqzjvmTEmOhGpS/daA5zbYT++ORRW1Tc0dmof3b1mBaylLETp
h76BoMpth4v/Ag/Cj0U36PopF2Z+6X/hl/VTuI/xiPf7XaCu9lv6HM77qmTp59hn
lIJNLlo6igRwdMkbYomM8ERZgQZMeUXC3wfOCQ2Hr0bkexNIOAIOmnGs6XczVHIM
Jme6nj2NBx/JBFRkY82abyxuUrneCwfHRAaZ503TRsNDyiphor401cg/mtw9w7FE
S6VMuRwuPKgHmaJWqEc9REaaSDF5PPJeaUIMk7DT1WHFFAsl+xl9K9yZcvJGHPdw
Y+AsC4dpTFLBrO3TZgomuErUq4/MAQZtDdZx/H222sWk2MOrBxIQMpCm8aTHbbDJ
j64EPxAoBUEkMb+8uhGhTWOYqntQbz4itL9ae+AxKsi0firdRROTHXHmgYZxBxhv
0xXEheku844+frYLl70GnefO8Th8tj9wUaXanK+ENmc4dSHd6m7hQwlcLShPOAF/
q0BfWMEcT6pHnbEZMSjsg5lQ9nHJ8VxYtiBHbbgfOVb0LJDFkYlnew6et7gYt4QW
/XxRXsKum7Fm3Q5Wk7F9tZAHmFPDxd9X21EEHIbyi4oDyLFgpds/g2lSnbyxrL7A
VJ7vDr7lHSJ+9fasGOIxh8k86sVZOiGEj54ZGQsOjCUg9ogQSESJLpmuuB+IH1Cm
oeWBZwIG9LKq0l+UeRDG7XXhrlxLPj1hN94kB0SshYpsSuC67w7FHaTg103WXOR3
VPH2/ZfBAT6RHboXnsdxy5/d6yo8zZ6iYvxrnGe+1MDf3dhlxgMBBZRIugvpLrZ8
5JLUAzxjeKGID3LnkcPhGMx7QYDFxyNimEeIFA4P4cNsivbupg0uHynHCuN8xB+u
VnnCCVB8AhXtaEvx+t99E3qaGAVUVN3zfgpOsbfcdO077+TCUBFu3Lp1tBT+8nIa
z/bmX3hIkwFwA1J2Wjp2vnPSZFPuHNl/9IXhxI/P8yt11fP/TjAF49+o5fPJ79j1
E+UZW16qnAdethgFg6BDf8+qBpCaQ0n0hPiFq9Sh1vhrHgIWyzUkQGxiLfgKMCVf
f5oyBY33UdzGowm+5qN25c7U76sVavs1nb3brNlE1JaUGvNwILTb/c1LnIBARwxF
RFXCT6/8t0P6G9+UVkxhMdHrQTTlBHSoNCXyq6j5Oe/NoJmzBcnIRe2yaNPkfc6U
Mu9c0wt9ef9cqKETL7XbESHTa5hFVOAFX6xg/0wKVP3ZIi4PoB6ASH9qFBiYUdi2
IzT7CfkVEWshXtWTBGg6m+u/wPwYmABqNK6nOaXaPyhZnxcuy7vbWaTUDTxNS5EB
P1yV0n+G7NwquoKj2fnFhEU9ClJ4CjEDjM5XZPogLS4cMiXJmXeuvMfe8EAIevWy
hZ930JnmHjaEfQ5VSNZ2PA/rMZPcOoxKqv/rYI/WPv8wqjbIHpUIz+0QMpcbTtFT
A8QPJAMo/abeeJZ3dJZa5xNdYOIjz3g8KC8zq0Rinu0i1btLrzt0vcDtfyI/WMEg
Cp2+cru9i1GQjsgy6WIbT7DlIYWW6gepoxO3mbHJ5y9Gs3ETyBMt+50xSdjdH0YZ
+oN3t40YzRzWQMaHPke2BX0+Hdj2F048CFiT4QHLsVzU3YM3O0H8AhMntGJ8AUv8
k/3mpSPTd+rY1vzbRIUt9j2bGpHHhmWm6tCQtZR2WnLpsXOVpkzCo34GisDfVL91
31Dex+88bPxlIINqhNqqnUW4D6uF0ZkSKzdGzZ+PpH6P6A6jdD7Ix4nVIywuOKsK
QwpvB+ab/9TNtSzethJ4Jqh0rh0jbvPeAQK8yAxUXxSu5JTv1Vnu0K8hFykHDhXB
Um/ZubUIxMvcUwz/E0eR03Qx1ElP25abztfE6igzCtnzdrVNNWJxDmuUSON/QZ2M
lqnEIrhFD/7h7/jfb4b/qWoDSe4QGnIN9oHAhu96Olr5gcH7WwSn+BhAh/ssQVPu
+veZwPc2GpKZaRyzblPFOSCu5sWrc5dk5jpU2W3jdSWoGGbi5uj3BI09gd6qwHKq
t1qNMr0HEhZ5Rt0uhWusoK0a2Gj5qOGgTsYk4bHewZvsq6aFXu0XG+LdDl4+qBjc
Ar/LOGH4EsnB50bTpPCMjmNw2rWd28mkB9nHfjr+aPU3YTzZYHGgQrUs+vOlejYD
ElJmWdQXO1dAAWiAjs5wcIdflsMzGRXUejiQs+XTUNrVR9AmTd9NphZz/tJDjdNO
H8UiYZSlnT7Q1YQVTFxw1AbjL40AyUdp+GZ2xSZOv85sDzedYs82euGpY/cHCRa/
TBMYkQ/9w56MijmLlQG3osNdIiHmxBBNWFsVowY7dV9mui82mXwjSzdlUZnGeBne
xOZh+RKrFyDZrbwXG82Gkajh2tI4bB0qq1aiANTWLsr2F81VM6e8ah6Bv6oZ4GH3
CgIytT69wxtHOLC1SCCcteet7D8IS9hxGndOgRa9moVyzIHxBrIuEcMjLahIhswy
AeqWLCnrFbu39yS4sQSTIRwK4Tu5zFoOQxYNeEJ1OjyzHGHzGXY/Jjx2nNjugxNP
fcSqxtMJ1xjwWb1QTIzJggQMg2jGhg/s7liSyRMrrp4+ZNVTXNI3M8h+8pMRShUD
2SPRfys1GA4FI8tQxZynAiJwc+DN8IIN3dUf4bH1az/ppnZ780dyKjwMnG+jtjtp
G1ifs6lJvde1MDLnsrE841sJf3SFqFDYhWHyc6ghh0cQ5wDHbbK6ae0ciSrs5q9E
SMXS+xR6yvSGRpRJ8t9lq/9OXLrkSOC0Xi6V0CWDtqO3P1qJecH36h8xmWkCymTz
pWaUqu2Vo1RB6lyvYnk/WgWARcUDKkZAQEci4WerV9mw6tmCXIku1BOQLMR2Qla6
8qsmQcvev8RowckwjSeRXTiXYQvVhGTs865KUG6sG3TpZwQQlYNKbHmAa8uvdeI8
Mdn1hEdPeOEb/okTfc/M4zO+M5bj3xOMw8sMPixzz0y/cdSqTl7w8nQ8C09wl2gR
GIaMYdH1tazZhjYaQ/cg6xdiKKrM/BuSequIvyu2U/7H7r1LinM4HwdHetxlYctG
6qqvdJxUnlaBZLuayco6F7n5EDnV7Ky0X1CUsbOVsZeXR3+dU0OPX6XD2CJLAp29
NcOkPmwMO7D0GMIJRMjo6/QwmQtRQnU0ge88Z5/4wXObXz1uRmleJl+tL/IYN8wB
J4fyOd0KHzIBL7oVg/C9jgHLhfb+v7Pxzk1CzHPy5hcHSAnflYwmjzQGCNJYJLPT
MPQnb72UdbCPvhA8noicSiyZK+Lq5k9jJ9GJ0Wcyd8uEDbcXcsip2Tbjxcfi7nhz
CiUytAwEX/3uklNqqsCU9qAyOsWWeJIQp8sk8qjacvEpbd+rWbK4n6Rl5ypOZf/c
QEi9VOHkBFTbK2ZE4RMFKnUaw6SFtdaAMzsfYk61ULO5b7T2gAonNDxw/eIjWA0N
n4BV/xGHqUrMbroydl+S1VK1cAtMExVPDVs1UfIXtgOM+VQeQHxj7nEp6rcby3Z9
j1iPvZ3AOn3ITjbaw4zYyZ04zZvLzLETzGtN30DiDP+K8bHGQCOuAs8BtIgl3fjh
fO99yH+76So4uEtliAufH5q0BPbRe7FFhu96fC4jWjG/8ap0oglw6r0DzReuW2cZ
HbYDgkH2B3Thh3XvNWt66NbMF5G1RZ33Pl3oAMqIV/YuMxoVfg3lSAeG1LtbdeqX
77PTnZlKWMUhNAtS0IL+cSO+/YgaclUAWiTkPMuOYADuxNVHsxBZYoiW3wdBMn/h
YXSeSVCXYdAGxSKHuJlIjJSl1G13nk32LzvFxteR+O8ePrnRlf2vK3M+N4IwmRZD
8b0/OXBnHCJRKHCT3eMyb3XTCMcIBVMluWfChonG1CunzV0pFPcjNCnOTjbWuzAN
I/RmkQ/YbayjW8bcOUZZz+zwQB7NaWk9NJNRsoUlI7bxBkuBtu4cSzAh/+hP9OKU
j0/VLY1LDxBYfVtG0z1cbZExo1QvAg7G+eRTXTF+XUJ5zmCCAYKsShNzhqAjkruV
Lx9IRnZghRm/6dXF9nwyR5B/a9Yvkjy8ikhEzS3yd+M3V2yFPpT355gmnPIoBogA
UEHxBhyXrkI9ntCwlR8AQJ6en6r95hEXVhRJCxhj/vg9F0uXY1xJ1N1dwqVN25RV
uP3FJorXOXCHVlkkYEblpyav9QaGNWzIO05lGBSUiywXZTYjTCbRDKj3QVilZ9d7
h3+FJAR/sRANsNNx9w0U87x5glcEZc3i/GQ8C5ubYvOdnas69KFdUSpHfTOkdMrj
VxIe8uw25YrzvP15zZLINErMFKXcoXoS2mmySDTWe27pxBrQiALlQjG8AjSmiC1s
IDg8cv2l7gEoQcjShBTkmqPP/d8ERnw+8m/NuOdXi67Ph3Ru9h5S/7NXvDD4IzKP
+QhuLYQU0bmP42QWM0WN9lGxv3J85250WmkuaNBunGD3PfT4yrrS4F0Olav/0moH
XPcck27vyuLN/f/49m+ElHxNgr+N1N4gJpc0LiZQNFE22ogYxir8RNg0SO9PB1CA
FOWNG2V7fsaDDkhaACbRwzKr94Pnaxigu8Tg0l2rhuh6HqKLdz//nG2GRwyV0kc7
r2+MJ+EAdDyOQe7V/9L3vb8jQ4YkkrNBnne1gdNiFcpMs3/fgADb0bEugodTgh7n
BKuyd0yMyCsRD7BINaSkCE6Pb1mf2pZ272dTS4r4f4U5hgLdO1UvurJUcqFWJYWS
x+pJys6WndW2xGBLnT1v0Uhc2wzynJ9R2NXZXAIQ8JriY6q+Bw/YEJ+F3fdFZfO+
ul/KzhxoGc+TmS7yFjvHpOAJ8P7wi8Bw0YwV1XrSBnr455hXsxHta/0kfGzs6vJo
LCQSV15GfQeQ51wWsw+4kV0x9/Xa5yWomoJ2Q+7ap8cEf91VtKD1FPUWHhtn2h9A
1i1c1zonGk3NmLNWS0HSTYUwA55Zm09amHS1z02jw679+en8kD0tBHT1FN1fx2sC
CInY7au6rg5DhZhsYF7lv9qyBf/d/ZE9EEaMscYY2uqgW0ZH/twtgtQkINYfJycF
T+2S+XTvRRM4YWFnPnlLFG8LiCVzmt0S0ioFDZhDcJIOjlwZq1ZPM2aZw2O+Y4Xt
W459r/P/pqDBerdDkXib9Cr3rOh8D/UsdT/6RTiR2FaDrxMnyT8PAVsZsN7LjuE9
z45q/PuALmUxfzhf16P2xWPyuByNYjZ80403CkJD3kIEkD3hCbz+OPzeNr5upZm/
lV1rX9B86bzxXVftNg/+O4XdCkLbk/lkggUO0RPr9td1CevpGkJW3O97qhR/u2TG
NhP22xWdaUSAcj1oga/APWqW4gHYyiWaXffi+vMSBk9tH4mt6BodwHI96bJKKYy5
IlkruSRzVnuu1m0P+RlrrBRf10s+d6qLmfriMMuB79KOT4XBwcLBDS9LwjuYNcRr
Idu4G/LE6By+gg2Tm7f/2pGNz99mhjtwF+JYeU5MGXaGCV4OS1pWqMjqdzvWKtBy
wT9Gq8VgPQNG4umqpGHQODy/yncpXVyGAhZbFbImeEM3mLwk/pBQOi4DAQhvA1e7
wv9CAwzqVpz4g1HXHgqGx8DizV1T32yMjvLYqM7KxPatxaz3AdGXg7psAZXGDs+7
oex50YjBZ/1RbZ1a6Rx1PSFxoBdeqUpLsjuPBi6F9Q00QVZdeSXCCgWQvBXj7rws
giF3b9pg6myxu4hiFoK1j21RgLy2UsF3SCBeJ2yL7ntqhO/gLASlXGJkwGYKzAUJ
lHJSnK6WZ9m1yy8A5HDNSyZXjTvTo3CjLQPIxhgN/f2NSfwNEkdR0y4oQ7kLljvp
1cSfnCIU2hIrTq8VEdkDRmvr3dkNvo5Sjk5mwIcDFBt5JuGlCPi2xh5SBZD+glsF
BesdAr0PpqO16uAjhaBOoh6KxVGVWZDK3gl9aQ4zSQl5kQLayL1Hpx260K+psbnZ
ABEbH8c8COtR7/tt+HyCxHG3cUN8rA34BH14o9LhqSe7pOpFs4HAQrQj2cgvWkkS
23GDecxJkj2nG6d+/yGnwIYUkRt2wOxStVRQeiFGUNJCZv6725BO7YQv96cuSS/y
3I7oVGCmV2tahQWrKCJ3Ts/ptsQFFr3s904V6zVHNJQ7/X8tvIm0za+cfQRKju9B
OX3cEN7lx7dMxpA/5Q2UL2R21935TH4kg4EqM08hZubxT0ZA/8flhY+xEExr43kA
+8FXhbPTA8mx6fSTP401/+XwbNgpdCyE7rRL6HUcvxFVMjKDWoKtlnhF74X99RRV
UEX+ijq2ILmuLe4R8zs7IJwrSS3/4ttHlsmAsduowf6oLn4RXnSfXPBeXIduysSn
IqUdehqczAI+sGHKWko8JhkBDDbEFXTe5FqCYWzHwaUnuodY9Djpw7lNa9GAxZia
WDiJKciUZGDAinOJD/t6kfyV8Gm7YrHZWQY6O8GFDJjNlvmNvudaxiE/nhZPbdyC
PjQk9WINnjsAxT/hZt2QRqs8kW+YvcWJ+gJEedavfIW22lT3GJo3zep+Rxg+A6v/
AHzNlx6SpF7YIKpEPO2WzmE3JiOftPvAi+Y+g1gtZr4xpdVpPUpYMg8VBQFfGY0k
WiZDRdIZ455duYwXao0tktZeMtC37ipBR/DdTJxYi1Ci7/4b43msEECMB2+BWSNp
9I5QELqqsGs0xW/tbawpobIORRWHGVPyXuRp/oI4rI6otg4Bb8FoFDdQWUPHvigj
Ysz6iTd8UaqvqbnXyZo3rqp8OxWPaPBs84z2ndxzcrQwR89BgCJo6I8Anabu8GeJ
hpOny/QC7ty452IyTYo6WJFm3uNl7TI8CcWJTmoGf3JZAiNGPD9yk/wJXhkkhbLu
UgxzzLNs+mAAub61ffreHqZSLoz7noSt+Yxgg0lqDDVgsFuLn4EwO4J3zzZR9XGa
AynxkwWFUe1fDRSZDLkQ3CBdOi4T8TDtwubOj7cHSJjDS8w5xvIEh1b03CD865IX
XxV47z6QTiDzDPSJORTIfG8II+aVq45HVb/tfityZ4PK+fT1D/WIVyAs608QJTYX
qa1U0tKHoqKI2rxgMmj5AGsX2JgQds85DIp64tXsRSgLbN0807iGag4YQt71uPZa
LZGquJ8ex1hUWgdAxMjDFGQ7V6IMUFGDYoaYNzIkCWdo164fnIv2PLVgTI8XVrKe
GILFGAVJHvfEPS/S7vA/qXtnA69uc4o+l3HW2fP8qpPkqeg5boE9CmOmf0MYlKhV
vs50l6TmlDA3+Gi3bH88y8BQFS6iTZOEw2HqSJW+4+cDjTGFOnYj1WwSCLwojrQt
ymangWrbiBoYkw/ejdThiYFrvZNpjIUf8y6nt4NFMusul3+0KOdb+R02vpteNi6G
00x6rNTVY/XxhYrHQ+9UXvJH/Av1/6mCq1yXScivLBpGr4p5zX9u5Q/fnxDJhR09
Y+lQsSSLJNsM1jIq0+23iZlWS1OQL7gF/XBJ8IZ9Ttw0F83OtoOhvPn4AjDeeyck
FG8EVmjVgajqJaDE5GqwOyjfbvl3dZLWlWpmB/r6LYssIEFw/912ppJGoc+lV5+m
z+s6gSb25V49MCmtX7qaIbACQWM5qm6Ixjy1gIydIT36xvx+CtRiBlDc7DbTBOoQ
xVRjIcD/uy2FoNxX8iY3oTEmj/L5HH4D1nve0Y1vBKz2ktmvVSvTcj6wdLbdt1pb
0b4+AmQBSFiK6VzYpgW45LRDbiMO3E8E0GWQYow1RbSRSGaisBt9HiFIbgRS9uJe
VhSsuQWO3uk15BB7t1afGbZHbhxxZvY2gT5aOvJu2G1y0i47ljcReHHWwLq0aWMz
jWTqDYGgYW0idV97l80C7D+yJN1c4kVhVyq+5rzMBaGcmDhXQDf8V+sOr2pQnXGh
e6ENjLsehLnzp8D6u5cTbvRnlTiHD7J+VGBgaQ7Fp5yoicfJqTKC1I5LMvSWGFLd
cUxKT2r0/CcAFV7OZYN0Lv5I5E+QHkROlwtwZ+PJ+fc4Ziib78+ii0AjE3OgIgID
OKawfvEVFv3VFQOCQ87G8tojB6tZ7XEZtjJJdPiAFVgKyORiq/UgCsEscMXGEqZk
PAIGacOQRSwM5FdBKQFOmWYkDkuIIN41osWQwm3ZrRagzrxx5JL39L4NBvQ25RGL
ZnxWIfh3vwinGODfLVEFIaejCC9OKLmjh+c1oHtjvzieAtyvFbi72WYG19LsB5Hj
6+PbK7/6DO2wnjzMnRAmrGfcyrufqIYIuY7fg3/XD/JmKR5vJ4gu4FwgHXPyPcei
sHelFKw/dJ5AkcQ+MDuOF1Ibx08bxbHvoDsjFRIzmaBv+NnL7MYei4PHoFCO9AZ8
7iO0QRXlvVAc0ZiQpSm5v7f3f75nE+z0JsK0WJSLCDF+sbc6D2zqUHNRckKDJzk3
6Ja8aQbLKFFOlAWGoA6oY+wZf2SDlZ9Z/KxzVuX3xXIZHJilPf1LiBlbK8bk++15
Z0d6udhYSv9U5G0D5bj2tvVG0juKOx/hGOIj1oZkkTMEp+rXYGiHKFVic2TnyDGn
d4dScLKsYVF1+yqr8pp6VO2HMJmA6vr88LqYKCj1IkWZEyuC0qL9LzCdMt8+L32Z
vQe0XQTLV2f/Sah00jC1TgkQVd8u/PRmsHUtL9veYF338ZOk2Slh4mSOTkdnQZmK
UvGwGcXiRj0wdPpSCXvBdOhEcjmkRjYjy9eFjwzI76jtNNlP1M0oYjdEDpvkHW8d
HwlCxtje3S1nJmY5tq0YjLCz8k9As1SkO/Wazb2N2thYvWu6eIQgqsdrHzOmFXzs
txJd0wwoT7wlBQM615bIJSknQspverpI2PRF9ypNnXyGRgJMqCdIZxGRPi650qZL
+ZhFBz0FdVtl/EvegvNqr8FXEv9PZ3icng8XbUJ/dGqmdvmIWNWawVUgtVOkaWp+
i8JThFZ0rdLF/bs7kZY0DixT7zk6TjB03N6UyXwBFYvKvemdT4UIj4unC5mp1mHJ
MLUfV0pp4IC/yAf9yaE/9qxh5Nac7BXEVq363cum03v/R+quxu9CdQNo85DnVM3/
yHDCEs+zDMcD7PdhqyUTrF37QZeRGRgXy+frCkxnFup3dLAUKQSoq0GCrbxx8QpM
3wZsNNAW40ciLcxqLV9vamrTRn15VS1FP2a+zS4dlJoCQzdPhZopJ4JykhaFdrhE
R+2ZAOd8+dbMzBsRUAqXdeJCc9byYZ71VCUK+DaQqd4mTgv9jecv96CAECnjBQqq
2qa29Kt/V74nwY2GcyMD4rY3xO6rE4xPBcx0KFg/XGtePENrC7+BD9B1vC8wy7Zn
orrqYYKvIm3UbZpAIxcdr+UJN+Art3jBq/c2g1AyR/VShMXjNDirtdBvzcboXnIx
MWU3uGKYipqRcCg3fPLBDXFvEUi/szzglvlH61bMjEs9GzsQAFDMqwRYXO2eNrcV
qHgbZm4UYLRVbWLhY1jJuYzLS425bqFBiXyVlB4Dj+hHjXfGkwdFFyU5kptPIzcz
7Er1bwQyfH6p/3RXrynf3kzRWNQ0ePkKZQcEkDnBxzYWlgHplKDPAnXap6h65mk/
kzJ1JoLtAXFqvfgY1L+0XExkGHuQc4gU7SbrCC02l5NX1HQ0xJzX6mYJM3Hysn+P
EJEviaD1UkQwqNgAFLpeETE6CvJbOlQtaRiVIyOCdjgkYXsqAdMfswIe9TPD4djk
ee2X3Hk24DpD6W1f0vdQbuFnIVwrFzDDqGWc2Zj7iRL1k4fxD446Rd+qCK3EHJ/5
btN907gAZ6wqk3C25WBsQgjWOC2KssKRiU3zZuUCiRd3QX/XQ01RQWoIcnte243G
9kXCgOBWIUDISb600P2KfxiS1HbHYvXl+2CWwReNQ6FBvp2qgp+MPMuabfm7upLQ
AkyZZKFRTpg8DSlgd+HGqYj+SDmzM2HPgsIkhtTG/Yk5+iTdLSVUqShOSRQX0jDF
i9Uc0r1us+IWVSnZD0q+JxrkVO1DZhpv8rPzu035aMIpSd2FxVStl5/S1H4XapYQ
ENk1Iu9GhIOcrP/f8k0keNWlkEGiAGE5lmvfHUzHPO8BqHmprxC0uocNDyXct4dw
IRQDPmRlirM/ho/pSm7767+AGuYHtboXhBnLgeQW4Jp7/6csJv74YUjpWpYGRBjZ
bsUyVNzvspNXQy80PcmDcFq5NOax1z69uJYBiq5Xc0mwSMCXHC8QJuyFpUhiz2IK
oIh0bguo+dh5DjCEGcAxdSNU6fuQr7evTgJtJXO8iQFTNstOl6emTALJkUILkJN6
0rTz6gRb6So9owQ3q70Gm9kixmnFeCZW+PeAb1SdSni31c67JSwC+2J5bwS0bBe8
yo7AVfpdA/tVN+bhMiwRgIGn02dfXGaNWlWdlxgzC/r0B+XKwSolGhpgGBgdIapY
9yFPVUdN9IVNrWs1ZsuCiuaAMLeXzT6+u+aGLax0WOPAC6Hoiw7R9OxlBH5llS9x
YWStitt+phVLsTwIxtAPdltUuNV/bDiu7oltOpl1drvC11Wnd1CPxLQVLfWMf+lb
RE33n9WCnCmtk1PGR+IgGEUz6XWgH0vODKU7XDIdaNGnwjYEGg11yo2ZJGHdRwng
mc9jEPKcj0jerIFhruBrUscJWZX/tk6Go7UL4P+3/HG2RaCiQWzIzcE32OI/CwQz
NRyMNTN6Ujq90YFRuITydBGgpef4Q0tzg1PPKtvGu6NVY0zOZJcqCOeVRASxCqGh
fEbAyrMLnsISmZkygcMIM+GGSkM4EE2yN0DYMhi7e0BIrXHc/2l38G892uwlELJU
xGdlsHhLVUw8SPy4Lo025l4RomvZniOkq32m8nWw65PMK++ZWTsmV+W3Kcx2LsvW
eRFxEkGpnZfdBz+xuSZI/nQSEdr5zgOiKUlvQnJxzCRUqmDvLlUc8qPuCFfDyt7h
MLSWvfDeveKnRkqaj6UEamPtu5dOr940fbKnsf2oBTvg3nt+V+acYZvxZ798f7Ov
Rrt7lCFry8+G6IhkL1LpytSyx0P4Hd1SvJasIMqiIcG9erq5wpSQ8n8JICu+SqpC
RjQN0vuVkfh8Cibk6q5E8pQ1UsnaRChbZbPYMPALP4NqVppVd6UIPA+XaATThG+/
/3JMG2IKS9fXzKCLn53n841UetZx8XeADkxthjhkkQWhrSZEcieSvFDddWwV7v3a
OWzTOAh6t1UXqHMh9wTlOTyEEHbEvyxGq50IsUDwVLGN2QtvWD3wilWmoU1vJhgR
AfFHCYqbLfb//EbYwQXyR48uaFlfpN5z7LgdXFDK16i/YDnixySuPr5Y3x4vjGGP
KwWBlsOtrBgmGRHusrCIKrImmkrPl+cwauA4PkMZTfSBPZmcpBCwQuwKNGwet7R5
BNbBwU5tltDL2P6Ejz3Ne+nb5nD2Air7IT1KPJh6c+WWM1fy22iTlb3T03uhbDr7
jMGGnMJ2BceD5Zc0RspWeHThKCQLZ0GYDe2FFRHxNSkEkAP9KDIfaNbD6gy7msMZ
KErAY1VEumOeq5gP6MRmyU1gF3bZcfeq8/mVhDqQnKyi6sn5bVhkcutKzMZZxOBi
d/ydbuqoYfWiO4EqrVUROfu+Mf8Fe5ndOX8HUHNAHgAkUnRPA5EQxE1W+FRCWWMO
rNDagH5+EnB+kuyT7k+aXajTzOQIrkxugrwnMBlUt744cUmII5H88Oz96bIA8/NH
LIgJM5ExFLtlWM+DBgj8KHJa9Hf9FWNfJJOQ7Phfd7slaPEkYxDFOQ5YIAt/R+4F
6Gn8otjt1aQ65ItwY1x89E4rKrBgPTG3TXprO5M2LVP1H1EJ52X9pEMss4PWXTmw
GOxgQsIwlyqMAhaDl0KRUMheKcogCyFOwotPiHSC6qA04qdgjw/7Em2vheQR5DeR
0eoGlDOpTlp/+EkaDRAI54qKmTZ/v35OqUtc8TZ2V4mlzpqb2ugElJP1fL0L8d9b
v9PC6lpXByASEiiDuSXR6WLAzjou//YeDM54bgBFKl+ws5cIo8Y+Q5i0t+5jAurg
0a8nCUkMUvMWjunmUeD+btKDLE3IP+V0G5ZzLr+7k4kdiS3APFri3Hg24A1Rm1uc
VbvmAJbwIqbjrgY/i4U1e+Dl7LKgTpHP16ZlPvveQN+fiBAFoJbmsk6KLRlTqgBZ
NCYDVrdv3pmejpUzf5xffXzPlwyeA+4DEoKX9LD7yFrQKX07FaHQZaIMqpBxBy6V
vEk7VfRrE7hmN0R5YkKHLRzWnXSKIyPsPdDMMoJ8MyWfxKrFjYN8n6zh2/C8JvZ8
6Z0saqRVvrMrvcq66RccoANfwgX8ku424zXjLYPJyhx33VlVxcQDJLQYmO9hSPCE
gqRGWUbiPKHd4IHgf2lbhwSu+NOw/u6DKLdqFQ4gk/qXTUbu/oTEyaEK3tVaPRHh
n0wwohLJcpiXh80DWEfB19vdpDF8oWnVSEQfGuVBaHpedVKR2Uny30WM8j9ntRjY
ARDtzD3lzigpIdy0dmZWTY1vY/jrNJdy08ELmhpznA9RDYFTCu3owSkrfoQQJr7u
k3utj8mWPNuqp7yw3UHmvFnwFszpjQ77wbjJKlUeuRimX3mcal7GRENlVG9hVTHe
KItx871oTG8TJQg+UL09X0dNfUD+//kCOcrqrzgGKcfX4V6WtwPDk9v1CHZhklJ8
gJ75IICzAIlywhxegniO0D8l5L0WsXG5obpC/VgkvPB/THjOacXoAb/BtFaG5/qB
eebb+qXeh67G1M8ZI2qdd/HBhHrfdbyqUd6LOcveDQ4iJMD6nPIQo3TZKdLVXXgG
oLx2J0jyYhIA1XrqPZybLsxLvDo2oiAOvLn++IHi0G7YpkYu1eLaGUaqvwoqncpk
tNRP3ZIyUWdU5DufPAOlVAa3bXYLaNTgL/aCIlygwR1DADw/yBGz0zWRXYDIm+ek
xE41ydz3BUyeX2Rl45ULd0Edni3Xe/Pnfe5B0UOUfycLj6EjrnQHGgxz/eAHRIjt
OuCFzrErAtbkOYYVGme9gZV7JyMg4as83iBIpvop5Bz/sT0CT1pqB7XanWKI75pS
32ShgT55LrE4rDGuRUGXN/8Oe+QIZcE5iern+QqzJFShXm4yCIj36PLD4/Ob1sYB
GVDfJRZ3hxRlE3R5NcV5Xff70kqJAlhpD0CGV4SrFbGfmCqaYCEMxuc+CzQPoDDq
RZ+HT8Kc7aO9/Nwrdkpxs3KRtY1PtGEJJxTzE+Hg0IdpZH6Pk3yedzLxPisiYghV
B747f3jQIPycgauJ39htq0KT9DoVvqG8xd9JGTnHiYOuqyQXQLqitj3a/pHe+LQd
INQ/PJgRVTK3y1ozUz8G0K8MNMHp7tejkToeZVaBbRS6+OMV2uX13sjal+yl98vs
Mipid8pd65EB4VEeTAa6DhMyUxoZGlwlrdxkMHGgOvwBckna6x7dsyE71Vt5+pBq
bFiEObXwPK+XLwGztmnmYYVIuzjuxaoUvaF8dqerGkIQl0Y1yEMxRLTfqLBarffO
hG9bzrotp3BFafZxk39ExXnXvHBGvbVFkxCLSuXZi0nLnujQtgfaSh5lO813HBvw
mDFgGkTtycJ5Lmm0w8Y6qUKvfsDiWaaLAxMXyKXcBcPO7YHtjgDcEJgQ41w9m/NG
a0toS/27T2x8KjVWH7n3a3rp4ZcH26QP2VBiDNHiSjGNrCbYWWBuS0sF5cszi+21
UAWpYUGD8/JDuLvRofpu48uwf3UUBfCzBPJjRxaNW+4BHj8G3Cv3UdcrmbXmnR09
5RMeqSsTlo6Ptn+OOvUqEqcWk6bd/Kzou8Gul/Pv3Bkf6nW2VUCc4jY0AhIUksWz
zntHY2BBYTRcBe9OmsWS8HhNv1Y1yczlYjtaHHfM/YFsfshF/PEIdljP981JXHmS
9pyPaQRANbbOh2k9ma5s/3iyOBVUMmwXMVeeY/NUj53ejeEACMWZ/dkwmRgMRt1F
MM8MG1c1ujVKEMd0bZmOKZQxBVQUh2D+41BPYoCAkkdrrChJCaHJPsvR2zr1a/n4
IEO6Sj12eSGTiFWex8zZxdyR8syqWO1oi/Seunb8SYRS0+WGOOXtWnRij02V1YWS
ROJn7vL2oMbYFwhb1/wOx+uIZmA9/otKYcVBYkK6u4Q3JA1oRIUA0tOzjUPVVPnO
M/VyYVh2uHJI3Od1ahAugs3i7BMHb5kjOhGepV//tAJyFHviDBKR8f7F8WyUpXcQ
aV1glrw1g0E7/6sBrJegQwLrN0+R4PEOn66tR5DT0QiVAi7erdqKv+X88PtCvPM+
cCufjwnqR91uau0vXJQv+27+vaP8O4URxfUQh46CX5YKFczAWXZVpv9S0s3Z8/73
lJM2WpGRLOtqInsgKyO7DECX1FY7z6vVM5xIisbZVGdtlsaBji48lHSSomZcnJyj
QFkaXIjN1c4tyjqboYCLk1RS1UNaYpEKC0IDLyD1ZmPz6DKGSnWYftG/IZezcPDP
SYhIKPUorBbhUWQrmQwrLHpA8BX0rPmPblmRMVqwhptPNw/uVdLqEQHv9Pzyfb9w
e3kmekLTHaVzImyvZ4xXq68N2SL9/ZENXfk59gPIK408cP60K7jmEyQK5NK1DlYB
WoVnuvBXB4pa5CHV/ELUOMwSetvpszTUvNe+YkjySwWx5+54YYYtWoRi8+bRdgz/
CDQztKoN+iNbtd8mHJQCAM0eLJndaqoZQf2aceb909/N4JifqpQQbIHV94GsfvsG
mYODwoiR/oHE01BymSNIwvi1IKpGaRo5kiYE7grXDUdLXQjjq9HEmtLsXXXH5Dhu
cQwnK11LTiDXNQ/CcIvZo615TQi0SxsuH3z71Ma2Hb32lnFpvAB+u7cCEU/HDfwh
OWuFSUqVRDxREWtoP7WtxkZRQGT3iEz5CnAZneJZePD/mNk3xZDG0PEl/vkWYEJQ
/W/zAqEFxAtE///NYqKUdB2qZPZ793Cgz5Fdh03IdLx4Gvx1lmpPlqdH7TnhPgi6
Xxs/9YdJ8OxoupguyGf6+2H/LCNniKpTglBgAGrjXbE0lKdSa6pvis6WEOCVXYv8
d/Vfn/y1NmpSPJORW3UhnfTDezRJGEZOM9LGC7WTwBvhRYuGAEShygTKqtUxpVXd
dg7AsLM7syYcLZFij/tiGRjU97IdHfpyeSSFQaGpMZ2cJAShsCrXor3mTWU8bjBf
9cR0zE8dlfU/zHjUoV+5SkwzSgTgfobn47chjcvmyGxgNwsnqwkaMQFbL07IcNGf
RGbrToYvHk8ORN/ZTTmA+vhvxOgbT4dq/616SGR+dOtX3wjkbsOmjfgOc5QPiuHz
LrW6gGKa4c7Pr/7i6weJTtaOA4EZ2m5vHWXuNqouDbDcDJyJxwIqmMuww9vvcE2Q
HPZm3vjGMbIjawjTPS9RL8mViONVxAQxBeZzyyhbhAcDmslABPXfNJhIIJuDWebx
prLoVX+k5wLjNFXP6cQqUluzm6K56gqkPEIaVxegEzOMtH8fKa243EA2vDFloscp
ElogTXM7f1s4DVKGPGizmyd7++Rc918sQH2pxILhloKPEfOQy2irTmz2EfwQyHYj
UKKapsKVPzQVhIiEMVevG4vXRbVH61araKE2Y31MR2qIP9T3xrj8vmFN6prcuk+G
Z/i3YrwiX1LCeSpy1FSZKyKzeTozMkOjN8yYEBC+RB1BeTds98eKQGfU58MSmQvV
gVC//TsHd7a/Fw+T5+gw13Cld3A0G1wUIgPSMd1q7ntWaGifz8kfba/N80oODO6d
/AQ5yk0xg4X+NElMejUafi1kw9HG6M4N03JUBKXnBAFdQ6ueSuEguMVYJHugi4NI
QcBcGW/sXqm6Ba/cZ+2b/zbnZoApdITyIE0lPQ9CBnCrkHUBXzcXPoNTSN2ZBDCM
4JoAt1c64MyYnS4CO60EKIPhUbL4SFzQtcmMGFOQ/C6NopIjIlxhDHxCUHeODe1P
8UYvSJYF2PCRN3faNAVb9hQ/8Ta6Zrua96w213gOmRv5KaX3pQkrt++wEHpa+18B
QmKjF44Zl+tKEYPwEf5qmjk1ElhLPWoeCbATAPDgZNNvtlFKo/zgZUyANwcb7eZj
tB8RbrVM9HYS4J/aDrHXfI/aAc7opFkrwPg+STre1MaBCH0WJdxg48dCsmSSLI1+
mkQRaJvbFe2z03UKO3sJn/GGbon7X+onO6pDNtXu++Qo9M+hdjN5Teu5xJvLZ2z6
JgTj3EfLH8w/4m3b3fTDkihvHUMkxzkeClF+9x844BO9c3nMs5KX4+Yliz8y+9oS
+v5DRX8XsPUAU580zk+BAPfOGvOeos8JhzXWjy9gR0ux8c4LyLou9vnJ94IhYmH6
wUuYfYxFgehBWcS77OlULck5149AYGDJFwRGOYtpxx+nhKomOIVsw//eJjU3qIu3
2am/6Rx4vrgAdlkf1+ZOkFVU3Dpknc4XOKPbprz8oI7mjlwb8nLSnvh2mHjiLcFo
iTH9SAcDzKCBeg9CHv/mZSExvn9KYl9vntGhB8ROJwPmbN7OlOary16Fbsmh4MRw
MAZmDu0L3KeVKBfGDp+UXoTiJR9egQpK0tXQok2WXKfgdQv9yOwzUhoEBMMo9Dvn
7XRCl+b5w1VYjP+GDxHagZs1FZvi3FdmNDAY4syL1MnW9Ly3ryvECJO3gj2Jg8y+
tJIGhDfYqFKzKnuni8EtOY4ajRpo/Z+Mu+Udxi4UA4ivGmNjYBAyFWaSnSCnTjkJ
Kx9Pk2QM/tlJ1dCDSsOc9jVfr357v+iKy3Q0o2RXjlQAXnHsrnUqNVFgRPJoVax2
eJNfCftfs1sj25O3Q94zHp35Fz/wwvtUvEvJiaEa7Dyv4X2ke+GG8On5PSANIWaz
GTEGIACm+Le9nwhHfvyg1jJxccHNOxIVTBghBaYvxoPE6J8rZ5tt1pGDV1S3imBP
TwWrlvDVBPd+ApQS+4a2wo3E6tk0u7bQrCbEWvpixnUZ3THQQL3N06z7FntAzEe6
aDLdJRkAuJZ4nq+o3zZBIN/TJlzgMh1CG6ZX/ju6OTHH/z8OGp2GvCnIFkZxEBSW
y8FGHp/1KUsGY5QJBJAPn82QSvTGFNmB+d7g8EJZMAobky5jO+F4jN43N91anLPY
ydNmlqQco0vkzTm3mb8qIK3BM6TzxUI8hpwsF7rTMiWPcSqdriLWpEz2tt1I4JDO
ywT60f1jfI36G2Nz/1qZ42fIt7GIVfUZqSqaF06J+f7T5GUHECKEjnhD74H9ocNC
5afxZSHRqF/9/lxxRDzNQOfYcXFKH2SiN/HqZ2630ke7S2LLKauUGsTyUSqSCZXw
2V7ZPMbLRdXyZ9frzcjbwCL77Q7Zdk6DgdC210ENzu3tehuunY9VDoLDMFnwf1uT
rY7MlhXtnUyEzZtezSjXNYe/K07AmfumAew0pGD4FnOXWACEZMjc6KFBjgUi431y
uICDUR9C13LRqBr2ImOUVTKROrpqbKWSiElBa+TI9f+y20Qgk+VeWnrLsf35AOg8
8h54OVavod1lP1VuqKfLu2dEdcorecH4oZHXfW1hCoUNxxJ9heanMs8GGwDPyFnq
kbt2db4EY9hT2Qar8FD22dpjV29Gy5bss8MPIq+fsI1kfHb4khp9R0Pc0mXGvQeb
0k9bywZaoI3B4t1QrefH5npw5uGyT9hTFN35a2Q9nDSEeidYwPwHPdZLonPaSmCr
1NmwsBfTzpTh6NlxsVbST9/6JRdwK8kKyy5hUtu9RSnLHdzis8JA6Rq7ok95xsTU
8eZw7V7o0Qheg1JXg0UwGSbJUePo/cElaLcOKHFapF/0cPODrVp70LdhkhG2Vxo/
fU6Q2SMSC6PAGBd2EmjL+UOsSnOw/ObbpSXwtyisJ1i+SIyP2tj6gO1+6POD7nGO
m/5ArW+jjne3zlVK8g6/AMwALfgnEVi4TLsrBObZYanVW11ROyS0Q9cvKIFcHdWy
Iw/3aJWQKR+XyatinJ10hzIUFh/kXszp60CnYL7UP3qX9+zmRxNsOosDkKB2bOo+
fBMeEKnKHacCxvhBrTz74QloUjg/+7tF4LlhG1waMKgWOGoClfqHQbPT1ZMGXvMx
pKnmvMGI22P6cxQeqUN2MP4uJnWIP6JBigAyPsdwFjIbQ10xYGPGT6ZNVKMJFhJB
Tv1EjhSUpMxsgD7j8UAC6HvCQ7PY9VvrqqvnI2hhN1Cf5Qz5xTF+3Jw6TqGZ1Gmh
MHoDHO9PqX8FCow2PD4jR7kSORHvNO7GcRxs2V67jtldD69AFfM3yq4RkPMaOWcK
Tt9TnS8KF8CI9iMU5iRTKW3Ypp7IB9jlnhSBmtZAslPN2eLCJ5oNc4ueNOpr/yMa
QNB4sd2JoNkS1JE27QmLtKIDUPQ6E+M1RVOkLZ0zmB1ZoBiQ/uzHXidLSWEtyM+E
GZfZIoycjzoLH7TSPslvu3KFdqlyhT4lkTSKJYb+a/ZJR3YiTBPV7ynJoChulvw1
SdkjR0qmIWRGYU5G90/dx6yH3Bt8fJOLX9J3ML1rDb4XlgWYMwN0JkPe75DVrTR5
I52rgECRWcb/CgbJKcNULhlPxYkXGGVPOgQ3+6KxSFS6zloNUdfuCHGOoN+xWRtB
ShBbr564d1g7KJEdXGSn54K8Yl0XqCh9HGrtYq/KHgQ8lyzWv59C5TASASob9mSL
0U2hWtNpHjzRGfP6+BmNo91EQCjnvbAaEth87SyIMCTmenkf0AQhzTqj4oyAEV2e
gqNVapDTlcGaKD0hZ95ZPw1hctnVthhvRS0qBFdCP0MvMHHAKmyL3LgFbf+j8DKK
J8Spcx3ArPZiq53d9VxAbRV5+ujiMWz2gzmcrCAaYMnalSuwV4FXn16FlObY8TLH
lAx/oWIaQgZQ0q0TRYLCOMwj34U6N51VCYet6fdU3pCow3/Qi4yAQ9nIT8P8Abei
WdHuWvgo5PQ0w1au8dDQRJAFVXXrws/J1gVa9+HNIW2AuBR0E0Lx6J6sQJJoUSrD
KSAUiw8aGFfNcVHa1XLzxR5mOjShLPuOGJMQphfKhvl2Igwl4H99oXVCtV4pmIEl
BMOmWnttiGZS0/wTJ2hPfbUS7kNJ8g9tAb35Zv3R4XJleomQzmZ8142r99p5hiIc
XEzUFBwRK9VW2n9n7bRjvmJs3OiFUpSg9V2W4fKFVYwIi76nDbVyQGAXzTUsUFK/
1Hce9D2k/lj4vSFpm8BhpKHheQcUYyvfWhLv+oJRiQ1RfmujY1lb/ky01mS1qnH+
QM8y2z8HJqt7dPZIbCEA2QZTnYJjegopH+AV/EyJmPfOUd9X04D+j5yxi99WdtSM
jQbMzf/k9js+ApWOugbld2WyJr44Fj7MKspl/c5BIDaa0Xl3/Ul+K6rIblVVPFz9
XxuxZ8tazWYOsHp0ksYXmmHt6928dmjUABzQEU5jkqLG3f5+NaskZkf4V4Pl8Hq0
xN/dmVlEtO6RphUBekqiIYyukv3TbEuPXWztWt2sm013d7p3YyZV7ac39IhKHfUb
ToD/yePrONGtTyXD3/VeBc0/II56DGDMcdp7om+ROfmrA2d3KPbne0ENyPUQwbq0
fwCVGp1Uu9yj5i99atMfifBiiTHdmgPOlH+9Muc4DZwXBZCq3x5ngGN4eSBJA0sT
4pdfBXwCGH/Fin2Gwd//GlVcwyhkxapUZptJU+0fsovZNTHjuIO4sXTUluUMQYvP
qS+KD8pCps8735SlSagrE1ub95vSU3ZACKhsLI2mrF5qPaOfpirhhkP0goTNp/oO
+80Wfm0dwJCKB4+OM98kCnSpSxPqnEh3oGN2+K/lVa4YSmldJ6gYgCuqOnzvjBbl
EsCDDGZjzijtnq7HKjlYQHiV5P7EZRmw6cUXkK8/qDtV+bo8WVIBG7bME2SSe+qE
kkLVBOK9TQVDcbcyzZUZ7FfjXINaGhIXQ/MVUz3MBzh/Y9prQLJYLR5pokRDyAPM
zDqgs2pWoh+fufev7xSSrMLSVBOoyPmvjj1wj4eFvnWXKKU2GMZdnQem2GyAGEAF
JRyiu8m/2I6mySgo76Rqopda2AgQmZ7eHNUsCzkSbX0G9T3rlgxpPHl+ZbtSa0eS
iWhGPtKx6ZATJHWyEBS1z8paAXvdviUs+ALP/djvlx4D2x16pEc6mL0KE5r3ia30
cbiIlBcHlMZ7qe3E248Kpok6FA9F260f8LnuSDG9swmTXV8pe74U6h/2hx7OBju0
JzVYy/658GPrLXeN4mlrNNGZK/J0HrBEE11HoiacsAy8QYmzIlXQJZn6X47K7Jf6
D5xdbWmvXq/yXTjrTcQvkMYGlkTtLAt+UrBoDl6VE0ZU8fgJIFuSreiF97HNJQPL
rfd4baxHx5MOESVq7UloeerjpBR/jhCJ6fArFUYbfe3DrJH+dCSB6H5thKrl3Tns
xHwmIWerV7Ofichz3UsSFT6mQRUCMhTHkTbMP3TrI1TFHfK1wOuxD94DKL2T6UUM
fGsvKIt6Ch188gZ+s+sxJTEGzu5U2W3dG9GRaDpf1CX41wHzziy1G1OgB2dHbWa2
p3O2LqzpzXzrJOUJtS4O62Z2NpzXx3fxsFElJkfNMbPvCDSGlc7cmV67QITvdNCS
iYlcfUNJmyPAUwXRqJj1aWtsT5ZtSpkHSCOfKX2OwCO4dtxtCe80TYMzWPNZClcF
chw6Vhmw0//iSI5v4d2fMZBjBGe58MoTKfC8cxu1UFiYAvRzVUGN6lx7TpCtAscn
zUunK/97dbNQraP0EIprohmtPqmXefKgw0uU7crVYt+qjFT/eZc5huJdJK6mPP4/
kL4Wt6agMT5lVpGD8L3m4zAjRm0jLyV6kaXpFVaoRcydiWcZKJ4u6iL6mtY0tAiF
XQpYwUDh9lAiFHhCZLzypD8or4OrMwvi2VdSoqz6YUsZ72wX+OpdGhalo1K0qwiV
kQJfqxPrw0tTyGsNGMCTI5NCMnnK5m3nJcOTjx3klI4Jx/h8zqBk51kjOT4AbaeB
pWWs/DBFiXVGwNG1Y1DrDhgMcVryFdsIMrQAq1VB4wK4Hjejj/Npnz18nnlnB8JH
w8GVo/OBhnQI7Gfg/dZ8QA/qCIDGEmH05O+uyJRMkQCL+qbqjB6CJQyMDtw/CPNm
HuBnL59f1pyhzemJng/Vxb8uW2XhJFAsWbfE5bOqmtLUSEZ9isLfLnfMczBV9g4X
R2g1qtG5pqBxwbTFF2g+NiDUBm/RCoxMuw2Uj7XQjVRWGlKGhmCAJiWPnxyZqNbM
0bXGMQs9+bOalO+RMAFmsnO/Ozo2MUPF5RQYv4YdR21EjRQhSs0Wkr7GinW4nWgW
afWKJjLI9msccBIKtqL6gAIe3gA41i6RsHR/ARNw+ltnJaHhVxEJAaMnUe6mSE/Q
afc+7z/od6jOeN1AwKvJJpKkOQIOu10gbBNfyC+p+ywQdrDlWEg0PJPJYj3u5KYo
yBngaPV2KRW+dzazf0qYnZaVev9VSChUuYciX4MDfPtjDD12A3L2XMGxWnveQmPC
jQnVzQwu+cu3oh4e4H4o3VmecFBjlEeH6lTKQhBm9SYfaftk/RTHUX8u925A1b3K
Uy+bDQPA1ure3ejQO2X5Bjj8gsfPrN3EOXz0baAPx53588egwwsrm+D3XlfFd3ku
VieIwe36OHA/Bgcb+syWSdKljbQ0nob/FUAVAPfjONG+vL59vdp+TPNtGZX3qYoh
o+G6CiZO6PTkEyZZ/R0sI8Nvhk0isH7p4c2iNRq1VVd880gLqtk7MJsWbIsg1aAE
BSXzoWsEyY4tvU3l4jpIZFDXT5hXioHPSHcW0XkGVRmZjnsrnQXfjJkh0iHtRtSa
bsc48q+WhmgXTtYkXS7Dhmki0H4kDygD/7dncs5b3ybQhebd943jZrnky2adnTzT
CtLEZG/qDdmmSUzXAiMZsM4Spj9KCISADoPZAVtwZqz96qNLwYFkyeBX4kiEyVPU
qJfdrYNA58jlZTOqjkFr1nX27kFET534szev9JuQyQseGZ395ueQf11YlChZSD96
Xdkni7n47GJpOOUh1PgL4y4v6m+ZfKXDj+Sr0mSJkcJaquPpQMve0TD2ddd9jyf0
jz4EHYeNe/f4rPMXliP3oncBFpRJcxEQzCThsFPMi0JQ2m7+SGBfnV786q+FJMgJ
7ySRuU0dqvOlctrsp5+/z7xIT2mGO3GtjIBcqIpbFt4pU0XJqksWGgdZjHGnez0+
fYNSJoDA3+cJ8TbwtbXQ+p9VY99tWkaXolA6K2J+wqcIS6sDuEhaGFxHYxOSebZ9
8/ZTXZcD/xNKSiI7nOJOxLGRGSGHAXb/elGFexlipXJINnZrapQVVJZ7C4ha9WuF
bJnyURh5c9mqDefaZtvX0S/ROhtiuGMxCbTLMUvFufeq3O+tT3Kq02Dqxkk8fy4N
HmtQtJy9pJfR3HyTmYUOnZG7ptIVJOnu1IpUBoRwrGKmF2S8u71rHpjgx1Pgo4Qe
PdUWrMUSiPGU8/Ajwm1iyVHqsE/2I1MhuCxn8Fjw+Lhp4SJ73H/2CLhHYMTNaamI
W5zGmgaoC7KZSHcJExmEWAStALNfQUg4w9g+iiNTrAwLHzffNkBEZOu/VHN+ztL2
DvmZKixQZW2JiejHIWY44xbCyGLxmQBPiBV58wy9AI2d7pXhLisCpVEbXAXjw10e
f1c0B6DY+QKyXEhpjOmzIM69uazAzQQd8lnIidsQPbKe0l0x9T62CS3Pfw9qD+wX
ZVpMZm/11f49dqQ0idD67W3hc+/NC8NOdoQHk3nSPZGUceen8UdzHAtlYdzEsZad
udvlH1qIflUh6kIhFNghAQ3OlK6K1jKch1RaKGNf6v9KCRpK6Vek+aRKsRk+gZxi
bUjbDj6l1F/PLHpNuSJTkl41bxDjDGHsu5S1EJrU1MWur0J/tsTV8ShVJAxqx72X
32OwFGRxF4tkKfcmCeuPp/sSmN4XR0Vh0zR3ExOiC0ZNks3tH7LromLfsE77C+98
bflZ49L5vIoBu9ertc3Luw2o57/0ETLJ8BX54xH9T51LbmEz8Shl0U0MbUEHiwBd
+ygbYX+2NhyvWR6j45rQn23gM1RPdtdO9f4kdTpoNqAmg5aOIhBFeJoPf0x3pdb0
JCMhUEdcFEHA3y+FfRFQjHuSttFwakiVZSs2BxrBV1hAQVZliVDfqhPM4OYzQYFs
qWEXG+Rjq6m8aG3TzDaOYiz7wm0svMShkEeoKIFcs3YrhuSaDvqmH2ShHgAwkBxA
wLZ9s+/H0xl4YBxJj0PCuvL7efpoYJ/IsdKiB6pSa94GSqymrGhRyXCzmYaV2ppE
C2yY70DSwDUOPppdsOmbTgVdMi+Il4SiLdVQXAQ4itw7L/ObeW1qqfsTy3zVWMsW
OMHdNK0UZvQuuda5SoxisOYxb5MjTI7rBk0sdGH+BsFDphsNWJ8V9fsWsS8o79tD
rr98tqLyhlXq8w6AOjrPZSvkKMU9oXk+rAxJD44QM+/Q4ebhrywChO+T4zOENjXN
2ZiiB/9dxBioPbS/EP3ZV4yDBgeY1YYnJaNkyczGRAcHuWQskNtAKdHUYd77KFtA
n6gl4DPa4mQtUEiYiwWXyKHeBGtykLB9zS2AAbzndK3ypwRUQQtTcKHz3Eg5N/TN
TekUyXaczSZdBFOVGguOubmu3En52YJAEIdhFvMzCyMabfrvTpTFjpRS3Dk3uwLG
PmbgHyBS6L7jw/QlTnbtrjpJgTGRJOBpNI61VNbQ9phPOMdkmxpePBc/dvhIHgyb
xSWU3O7taMRwzqFgphK4zF3pWjgHmeeXBWdGSRWkK2htbGV7ZIa9kNHWBmNT2KCW
AFjWS3hGHMzxbZeXPhK/+68uYF99Jx0qMpcOlRk1maBOj36GwZfumE1/0kMLDSe2
kOQG6mfCgrSrVobCcGFx4vfcHamEFAWPoI1302G/ZzeA+f+/8ffC9a9+vQV5Hfdk
8zKrp1ZCJNMK/QRpu9D/13+4ApKkYWlOKyFXdcpoLrDBu8ZNutY0VBlLKZQnok1i
FKLD1p2SirvNPwRkv8fdX4zfOAJE25zl+OA7IXBhJkJbC7ijo8solX3gXV3jAuZg
6+eSLu19EXbjzKbCqnbmsDsiPYADc+//kfdvil6Nxd2tF2ZjLCVzmT+G6WgiE4It
cY2pB1Efmf1lpk4OZFxAsSumUt2qfeUf0jL/5y5lJayqedvu1rHxALqnNYOw4O7m
AwKTLVrji7pL/QFoBC2B39P+dEgjF7Q7oRzqU6Ohx56pBzVhxnGbjco4D64L8YUs
rkgmgDMPuGg1Insf8q4FCwXyaHOE2EU8t2baSX1tp9SiADThwG+0pqH5z6zJDxK7
Gu6iuaJndz7/xq8pF26HhJ7AwePkIfLKuluTBM3JmUZxuvVPEgzrEr3NNW7Do2Uw
xFZOPCzRJU1NppnNvq27cMjXPy8/5XIm3Zoue1jUsUDe5RZvIAKQa4TYiWJ5rmTg
OQ7zuGPrwZUwl79qZY4EC0K5Q6QkWBj/f5S8WadMdFFEmg+yOHXLhObLDNpzietI
8RGORTV1/3GqDDoMHc6x+2j0r4L33TYy8CZVYtTib++J5gUra3pDLpACjbBdIbxf
VfERevjwkTRLpe2mDfLzbB0phrbPnp4+wwbT/UsYyyb747qh8Mym386H2FpJFdf9
V3WpAjDplDZO+QeOp05FPVQW7Cl4ZZ2KwbAzYmADCVwhLNgIiHDlhgcbyXLMd+C0
9E/Ig2MliT0H4r+yGNyplMYdgblvM0R/6aIlh6J3Hd3/RWFSwscmd1TJesjk6Rni
Rfa3DFFSDI+wbvrlsp+brOfjI4yBehA+naE70GBgKK5aX8a/XU/zrfGfcoyR/JbJ
k6YymGYl5SEQFhv0BMbvzQGW5nP0RGNtb8RVfVynsmuCi+kdZzAVONmW5pUt6GSP
i5fd5YpotuFHlMDekPSqe8SK9hpg5FUIN94wFwXyrnQIC0LaoPlVkxcNKvWHfgSb
BwbtgdWYKRRdSsrVD1PAqN8hOFOUH5MGC2+ZQ1pNC47O3QqbUf3DQfJHqHu8VztN
qNl2qmy7RzCOeTy70U2Xh/J/ZJ/OgpMW24Ykdt095APRi3z0QUJHDAOJ93tGUENQ
AmsNhBJUQUTrLUn1DN+LOUN5+bAGOpzkUYJUs/GIQn8okyh70CwsNQVKQ0rMhRBq
5Mpqxb/nzuDPYO7wH5Q3NaWPndh0zcboq2W53ONbJb6wecEA8AwYmZuU1ilCnfkH
Ncmpa4LxUIMAXrDVBVME+BE+uSM9cnOgmr42mUTJBwRelw9EMqJZ9TuZo97+0Raz
fBfhrMkkJ4S0CUAcjNxdqGjKRD4rpyA2WXNHTzkxh2DFIdbEPuXPa3cBXR5wXOTq
oQumSAWh2SuHPdLaeBK2q4HOl3PlbCx2nuAP8D0+w6xWuJC8ugDkV63XT0LEuKIa
YWqXDDMFCEVDu17sYKa5eTqT4fWhgigoFB9JFdo6P5Ok7KvMcpfryROk8PKQR+d8
Uin1Y7uv8pAWRIYnr723DPY11vCVdJCIbZcz55MVy1vh8/v3rSeh75QazJWYm1EY
gl2ZzH+gIw3ZoelXmngtwrX7nMtWKNDrymlvbfWcXjCsj7MSpaLu3xdPuWAf57In
HehUdgiXJVZoBbBH8Zn6ukLKCJfvZeHppWqgrXSkI8JfUTjntk8+WqcSFXyqWINi
zrpimQP15Wg+XbR/YXt7Er2IpxyPLXtyim2gMhBNoQ9Yu5RwRSO8ERUea4zWxuwJ
geAGnZnQkN4o6HQHH9E8coETHMV5h97llC5SezcEMPQoHQzK9E14nVzSLJxr18XM
YT9vn4+w/olJIYn8wpXZNLh2N8myUPEI4vpAlaOFdAdW4+Vq15HBgx3G5WHypP0U
G2N/EesBuTEII8NE9DvWAYKABQvtwt4aTMbIiCi/0IoqcStaCfRkB1seocqPoBbo
vhfxE/Hd8+oBVcbnUx8U+c37oZzDcDhlfeVxwV1CcdfTrGAOPKae3oiCnLiK26kt
lIj+kHxktspAcbtcNQxRmUkxNydOyVMbiosJpuabJ07QUTfeXV9sCfiCz0kfOkkh
gyKk0xHYi534ENROxl3nCJctqlnU+CyNQYRx2JFSNmxdgM/PtwLxfiunh0YDlC3k
3Wh9WsFaDB4JGh4J679E2PFEjHdfUn6C7McWhSizNTxw315RkcPX2lKjDygQC8Qb
zNPZYlGE8czC0YUyRaeyuWTcAJGL7xttZYFnPLvKQsZTBtmvIBduLj+zQ/tiPpTc
fiYso90atW/lNRsrE5eanAuGJmPbSBSMtLlxoP7PqzOqkn3BKayLC6u00LGyyExq
yPg4DRb8Xe2J4nGkZ7K7FstSJcYl524dhS/iLkIkfjmUB0bSVlxqnqw6QCmH5rf+
HC8MNi8LIIS3jtUHiUOaYK1S2MPsj0qsv5PDjwvfPF4SwlDKXBjQ2Y9+Yph1RS83
P0b4iTXuM92WmrZr2tftBv0RybtfFj/adZziMC6Zwc0XSRtrWZk3vDyNvaWrc2xe
4HIu5jmjyqWHdBCCCmlXJPB2CivNAYDd6CI6Oh+ZMoVZGmgs0yWEOKSDPnsgnV6o
mPu58nKbpB5kp4M2+w5A0fEcpcGe7140Ekn5O0c2OUygpcwq5x6w/gz6nhysEaTB
DBcV4OJ09jDNbZKPjxrJwcT9xcKcaYbW151fyssujmcZg0q0WSJI22R2JlSmjYGG
ncL++Vp1QY9xWj5qPtMuJdC5EJlsyhNnK11KSGRk/jbn3i6Nb4CCo3xBP0C8avSn
4iutaWLKyv8y/Wx6RlM6lUoburaGn21iSAA9syQL+IZbcrUp8L7onoBsFV+M9gOb
AaAFPxAJ/s9grIDkuJhw9f8MnH+ejhMUng7Rm615UzJbCLDxy0Jy+DYdeF7IdU/h
qMc7ElZvvIxhSrP6Aj2n64zIOgLNoQwHFUfrUbojpC1zzlxPCKSsbuZkHAV75gsA
uo3gwQUTKf2XuLekh5GZKA4mvX2D20IsWml+dzcQSB6cv3Sqp6hYet8u+oWcsHuU
4HHSxha/DzAWRIAVitAbUI4YUOEmwRzd/rWQeY+9b56gRcDtCEaN/JZa/BT2OKRe
hnhiDiyzPCeKcwvsMiAOz5v3PSZ0Z0+yDtnVPo4KPOeV1T/ggvnPKoFdbHDk8S3j
VHuvOxy80HNGO9fUjP54r8RRIrzwH6RKH2OzJCaQscrSSqq6ImZX3qIjmRVhB4zu
tm+VdRe/dAErRgLanZ4KFO69+jJDeBhnX1YKFqJ/WGLKCQs5g8RRLgLvfi9pxWym
08WUVmFDb3Da+Bviy9sa3KU9prUHbE+hFzMvkMQKWxbhGMfBiHJJdE/Gu9nDIA+4
a6nKP6AuOchAmo73emzQU850pdOyQ8PqJsDwQ80WOjXAtYq9XQySPdggTsj0mpfU
bzAp1L5jB8eUvkgSJuwjg0S2uyQJgqjBX+O/iKySugTjj4nidBu5ITDo2/zESSQJ
HkKQ5yUjwbdn5TNzlWzpMxkRzz4rDFMs320ROg3fQJ3vF9fmV/JJn50ax2UxcpX/
kZKDeAP27pjfIGQz9t5lZYBhLXcT4LP6UCMr1NB78nK8IDRojOQzxR+EOF3weiHw
5yFSHXW0MaPyauxS3AYtra1/tMOchvUlkatUlhOY4k8kslHgJ/pmKi5ZHFtnJGkT
OMYQuWqt/serPFT5qVlbMDYY5iyLBMLnWcBf5EY4euEs+FjV0p2j5DiWJ+7dCP13
XvW2gZO2hGDTIko3pq4pDGukdy4S52wC2y8F2inRfmCM/JBVsOd53t8FiU4bhatO
ega6LVaW4+p6FwLpqX1YasaZGr2dFHCjCSicHj/SY99fFeRQKkUS48W6wmQ9zRTb
mrvafMjloYAwDohrQlBDmfk40PrRyplSBN7tqUD/A6LcS7Ijw+RO+WWpE50jn+lV
BJSzqJtKRNFQH2VGoo9czaM5i+lxSBiEZtPQ9lQCEmYt6KrTmNJWngYRygbS3CiQ
zquioA+vUKPlPiBH1UmYi5hCx3b/LiVuNfh6FADqHp90gOs2UrQROSxxnMfTzp9r
cFUHIOnW3hWpvJCDk4kKn73OnrD3gy1045eZ48bw4fGLyq1NR5AyYak6R/aVEFD/
UbdM5PUffHl95em4tCR3SEzAUC6SUgSztZcuG+PWGjr41AkoQExY3rkm2Ln9thKQ
FS6KdwgofYfGyHtcbIbWvfwKwkfV1KK3nvggTjENEzoolyoxI+raS2tF2lp9SH1F
SRE28FfI2Gs9Qqy/UkFlcaSmnN96dOjyIXzde1zqO1AiT37MogFDq0CAFQmku1Ij
RFQiVoBoKpECG+VyxmZNbk+gn4V3L1BBWAzwN0QiH415OnPmqb4aSsbypQPAm+Q2
oICYJ5676MR0e8EmMSxKYNZfjaBh1k2fDgMqCCPeJs2/XGIZhe+uviXsgTDD6ewr
yi4XSPo9TVRZTGDCihfWy+0O2Yg1wTQqW+NiXvKZM+CZV7KAaUrrPZrM8g6QD0eZ
zjc3uvTHYLnTsJGw9jiZ5FSk+Ru7C3bb77oFwuY6V4Os8KnEqYMdR+cbHm/CWmP0
bu++ngyHfM6e/+ZABdpfIcB7a4HICkTWJ1sUh9AI0aghFoa1nTQd++8xYhuKHMrj
SFCOO8FCldAOMcnDZi6k6F0xDyuZAmsdqW2dT4vzzOJhHiDMPBL3uivjyCOzUL0Q
Jgu8RFElcY2lPPWeWP7JU6tEWCPJVbdSTow3vVa5kx/2bVRk/ImzEAhLK/2+TYli
ZGLg01AwNQxRMg9HyT4q0a+/r5S4XbNuhOU4LK7A7B4wrS7fFa4MP1ThY1WVOERn
yaJVnlwxZagpGk+CjqZGGC91qefe7sd/Qjek2wQtg4njENabvLJ+DlqHCXAfxpY+
c+qxkSkjpvjDKWD4SVWCyJWM0U4G1SeztEbbiCRul8v6W80kYT8naJrrWUDU3Mcx
TR89uCq5Af5ZxE4/7aXSbFcdwQYDt9EQTmB2/DZGhAOkkacJCdH00Xsv2CSiMoc9
zVO24MMnlxzgzD0XgPBF7qdHDaeD8uRndYTOIUGo4O6VDk+lQG2lBfRccBoqg93l
FKrl8itov3YbBY6mK5Y0mOgtrAdXgAA160DEJmdLlNzGdO54nDbrSix3KaUMUt63
5hl3WEKy7QeToCD4i01vJyXvcHUSld7zYU/s5gjbH+0UkjGEK12sM49nGhXJ8FP7
PpR9ClI4tRdXg5FqsFSBja9mszIebBMVU+jcoEFE0fXHuJ7ZPcVHcOZGhWh5wptm
qN4vkANatfa6WMs7SXjcdT2v8HneZ49mveGyuOlJ0aAuS+q7GNuldLcFG3g7c1Uu
HUDMCJ1w/OMUBoPb8W86KA37EVTwKUFaBEqDHPWhl3Ue1wnW1xOWdA7bukab8pXR
bvexb9ssa26X7CqZIzjil2+nTIX5a86mbfRu82irdXPXvKuO6whPjQvxloGV0I6U
BXe3t1QjSGKNVDWycuS6JRioENqZt21QLhj5H+Z+mqHZaYy5OeOEPFJjbS9XYB+b
rlpQ57hRdyACc7+M/lGZPaEUzKcjjPwxlfDpFvxAOVe/eHx76d6rBxVDdHWWSnu6
5g5xcR9biVjTKSlNR2uaZBl5/iiHcTZuLsScAH7J5dMpWBdua7nMGPUwKRRMpb60
b/hIbFHRNwz5ZnZVvngErIDKiu1nyHBn8HkhngCiaHuPzvwxce4zT7EdPOe/AlDf
fjJs2yNUaY9pOQnWBbTWxHWWdl0hof4CEQz3ulqfXKiJWTqYr7XEYsosgb4QJu8m
9PAGU3xvqeN8COrTlm0jkiIrG9NZ/ejo5gG68KjL2bPbk3iCOn/JLLidThJizJcX
++/qkEZb1TfGdffKG6dbz9uWMBsrre3ZF5TXeoU02SE+1hvE00huK7KHgn7UN5/J
whFSdHKODBaZLEy6g3G+xNQ2XCOBBLG/GmtjpjC6e3YBasdBdeUB+ZqlSbvkpP7Q
SNw+Haah6EE+FHjpnHrZu0SFFCdYrqz/H+HGT6uBBEnyc2yQ2B0dfcwMTMmkwQ1D
OiPEGbeIvpbppV26ovOObDHkac2woTVMml1dPAM5VEUpUKHFsBMQhDq74jjKCZMm
3xA1if5YmSwryc/hEkS1II5Ck9SeC/4uRylLnluaUGzoldHPZyK5QJY+c9c2Tz+z
godwMLc3yjUvWHoWcLILxnhk8MvpGN3jMnXOiXW6lbhX1LNRtAO0ZUuqo3RAc8Ea
rxVPFIQ1iSq0HsZ9mVZ4eZrWoSIb3MgcN6g614HrYLwLAvAPCnW84yrDDkDEFtcC
7ZlYGsZfBhXzZm/kj7j42RSInIOSNfGkVb/FyS/X/lTnETKGgi7otE/yp0EDoleE
1Aq6wVUbds1IXRYGIj9AcksSdr/YxAEckOhGMLQJ7Qgk56KVMwUfPIafdlKdcl2v
9irVesPfgCIGlNQpWHJEqYU5OVh2Ka8vq9XmYkXyeVVN9MfEcId08MDqqMbR4FEj
lBC846x+LNgfKu6psbbkyLn60rF0ejVjMP0CNVXJUYgeFXlOBDesM5ueBt5HvAkK
BWloKI4k0iy6Dsnf07kH5O06eEN0KvbhPQTQs2NivXW0fcKcn6biHjW+PWJppMOV
tB6vhv4+gqe8cnXRcU/WzZdM0uvrl8q+UOa3aoGZGUm+BWKDkz+w4wJ4GIE6QK5O
PHXSwaTUbLD90qr0l23SNTTLCg0W6CsJaubiCy8ex7pEZ23sNejGxbsOb7/vytPM
MGzwZU554y+l3sjqfLnC3/24wSeiTQA6fO4y95y1RepOSItQ8eG2KVmfYxW/FGzK
6w8GgmGv92P9w1e6M1rHNjf0IAv3fWLGHTXB7zXindrFf+M0xdYSxrlsWdgh73Wg
1Nk3sW/R51xpUbFhhTSPwpJZAyTYJQgKtp0w4jhKWK+H+pINR51Djv1JyWE3gyhJ
44FGOqomANR0hoRgLogr109jCbN1kccBmuh3lSw0HhbiXOV1p9I2nLS+t69E36Xj
/lL7nO9yioRDEHwglRQo9tnplHQvCI6+dycvptmXYZZiLWdd3o2SwnBAbSjidKcT
V0olOrq5TVdK59edYcjov/XSHlP9FU1eyO1JZ0/VNoXgjX45xEB/Lv4ZuUUnOB2j
8e9HihMwexRekiubuiowObrutPge0rDeqtV0dNn6x4NBCV1/kROxRZhaJyfJO0F9
uKn73Ios4JQPgfXYzIQxACoFMJ/NjSu7IKN9XcDMQp9Y208gq4u4lLy3gV8gM7dT
wQWXB7E+PBNPuyo4zsCb0j/tI8+oqasQDLnmhaiEgobYJrAcYpmvnKqBSXTvyqyR
9YcXvCBnUa1MS4bLSB5r+wFO3ynMYM4PLNgX6a7jf0CcJXGIL8jz64x/ztTUPvnQ
TYT+f8elqncOEAgF9QnBk5c0JCIXq7wQ7vXq+ebpAAfB0+sOvBoIRttyfum1mfvD
Th+TRGt/0ok50mSxqZzfViNJBi8Clxs7BXjZ2MsPEqFS5DRw8ZuRuBoeSRx8Tv0t
GE862S5w44b1aZXlmk73xYZejDrEV4VVWnZKBi7iqzwnJMG8YVJGNVdDdvZ78T7J
JxgKLWb/FN94m0hByuI7xLvfR2bZPriMhM0wK6/gzJ8Tgj6dF9EBRqaTF9lvs0H9
8gHbwOBhqNHnazXhlMrU3WZSWb4LbeiXXiAID5WBB2wDaETfzvslkG22mL9F4ZIc
SxjSgWsQdb56422HEol2h4p7bmQPSgdTeRnuTwK9J1pBjQ6YvhCBVJLAuFkwyOak
EaauLFE1GuB2Nr58Vvk1LIZwpjMQPdPrAaJyzmFoc5MrAOkN9xnSHoq+RGIpV5Dv
FTBVHdTkuesG7HoT/c7r/UcF5+L4g8jtXSknfYUm1bnV1zLVLtGHARhP2bBFlHm9
T2CBSEV8p6ck7sPS5nhZ/FKUhca0CrmRdqe9vrghzQ86NdCSFdDv730zXLThlzsT
Hm18Yuh/dMN7eddZU6JLBY5h/NSJpM2mDn0aSIaXnOxIZqY8zP7S+krzGpZuxxns
54LfsFRp64nBq22NqqP7XqBBZbSAbljy5BCOys/xQyVsjzDy4qJ9Ish8L6yR1u+G
d3D4bXDBpxrxm8hJyLuF8NhWOzZT0Kj0mEBjl6Mu2cHi7nAnLfSlGdJnwoVyp4es
EQo4AfuMXsULPVK0Tt7GsWG7hiYscarBzOMjRMClAKmNwVkOxOm0mOdXEreUtPBK
ceISNdE8e0/R49P0XFzOcKe38M6lyD49uvfHfOHc61E++3y+PoNvBeD49lwCUv2K
o7httJMY3lsWVnrzYEQCrZBu7SsMXQQHZunaa38GaCeL5Fq3JDNMlAetnT0uzDiO
IwxC8NzRI1SynZQPSB41Sa3CJPk7nxZl7BKhaWPBRZ+JUDQtGVuFO8MdzGARyefc
LGLfdKoXfRetWhdOWJA7Y8KhNaM9+w9o9Bxq8seVrlKoEZuh08psr7aegc9bvrY+
lbnc7w8T3/KY4bqJZ97cJZIGtdMhQElJDaJetelaWlQiRjeoOJfMJxjvQnkjDGNx
Qi5bT6WGUTuRWRWhaUcoyjkwZA3lBG1WDIl5D67dr9Xl7ZEm3YyW9CZF25p/OM0Y
BLYz268JFtoIrobyoQ49C0ul+Zs46JQQ6lxqskbQ0PUrkBF0/r4FU+VOjSpvVKpS
HVggejyPp16HMURyJsDsXJx5rujZZtf2uwuA6XLzJPlbKsoFt7WEpWR2UI0RSXKe
B3aXHsVGmFQrko8U/9Rs6M6ouC5tD9w+0yBroOkO41WbZeDBtr2cLpxyzkp8tsJv
MgEqF+8VOml5pgo8yi3ofRor5FlKeKh7hwYrxwb6YVj4SUqbtGVy6emjiTY6rkLg
tg+71zWEZnE4pyj2SbZYR2sw/nK+hs8hC7oCN/uPh2GXDltoXNiIH4Y5HVDDJKfj
7nQK8bXSgIb6A6SNSgXNQ1FnWZr5N0bvfAEQy57/jy0GKhOedOATw3Ewd2gcqnOS
joDGr3RcCLihaXQPOzV/reXJPw4Y+3fs9aya59h1dMCySM5E/8xxk/LkNmKStnva
D3502Db02+19EeddKkh3e5+09IsO5rS/jCLITBkXP3Q6i3FL4xL6r2ugQ8Ye1O8y
8gHghQO6jtFNKlyaP+EFF5ezPPMIMYM9PstXVP6LPN3fa0a3dAaU+5iAdhaJF3gm
UDPqWjEnyxRsqbZTn2CDccGzxywDvG1KjnPLI+oeRUD+SD4g7vOT9gvOI8wMSnmG
89fEqfsGE5rSVlf9TP6TemkDUA3e7kuaCSe+Vzfh3Chh14hJEw9Nmr+qO8+iS6sS
zvr83ULZuYDFgSSGcBYUKlV0jwIG1OXeZcSNh9zVfbeThjf3qQDh2MFi6xzmXVu4
ehcMzUWJZ0GOpmFoh68EF5puGmWqspj6LBtyqo8pakmsJ8n3Gk8/LubjsnTyZH+X
Vh3OxnXYlso49eTMOfvAvAQ9nPHK6+nw4AI/UX+ga/YQIWmN0Q30OUGQhmUWILXt
awDdD7ZVDBOAZXPBuE3Ug3quxpHusFyhLqAxTwgJA0NST1DLlKuxz+uWVwfeVfrb
7GBjD83W4pfRYwIPP5vRKYT/nuKxY5q9/v2rmLcUR5Iixuf14jG0XgVuBUJ7Nbyi
iQWL5rSw0zFKeNo0iujHLK4oDv1gMLhEFXz6nxrHcAv9/ROZqNBC6ghSOleexLvL
E5eeqwjx/XuPafiiMAiLJlJNgFP6HSycM7FXSQdrBXn9b2e4S1A7GrbK3TZYa83j
DD45hcofd5XnZiFyPUjVQ33tzeeQ0CVoAdFdPOJZWRK+kyg/ariT7SzPYGyhlOjS
NPzvJovmZ7S9VZYAYagHn7/uerOWnWIt0OkjYZk6RBWg5XuhQlh0DaGcoOqVbFKQ
jQrOntU305Hxhx2aqvYyn5D6abaHSjcP0Z9qRzpFtmsRHUy1EVAMe8vcWdfa+/hD
xVB2E2hQgW4kxXq+gU3RdIo0GJ4pzljAYgUGL+/oRwWbLQrWOpOHXfZMzEjFQTKY
QGDZpHmGexqRjyS4MJYm1+EXzvrlMwcq2CB0ue4G7gFg2Nxgw+5i2pWQJVuEK8mi
jM90wb/OeuGDphH1wSY3TdBw1FIgK6UclmAEAkKEA69cSrVypueaHea7S0Kxcb4g
4Ow5QqY0N3wEeU494QSv//J6ysTx+inZsFOfbAWaPmlxbOwJXNkVd8jRhCYwVaZv
I+amsisFvvnCI5ORqB14Dlz8Pk/WFspQvqD00R4LaXvk9pZRB9NuxFVaOS5pdl6I
dDPm6snmj1v2c4I5p7cQ9OjFnjkC7KE4TGmFKA7m0pDaG4IsanBOIrPD55PyFz/v
gwA93LFE5vFId3gx8BIKA5mVZVcIwOqEBtuATUf5L5OpP62LNV2TNb9oWlpP4Z92
Fat5XYRYUQHXEtF+m0SlXYSFQktT3AU1tjvDhxAOv3I0tp+euOpPlGgopZIZj33a
udsjix6LJnIFf4wqRUwMbNRqROCGnZW5VEkmAecnN3W++XZ8dtJuP6m69IKXSGtm
JMIhIGXGWC8nI/Q0imnxj1gysSE3ONAuO15VbI/RFtJFKo5o+g/n2JVTEHJTlIOs
xLKhYYQ1NTnjErP6kROUplMRfTCH7iuOCDub+LlEAQug3VNk8cpWkBau/3FNSmmJ
PEgCBjqB4gmpO6hNzn1tmsg6nlKCU7vJlk+vKVreMK31ycwpbEDx1OwHCUCVWuJf
HTu7dDL/Pqm/y3ot8ci/vNeuMhhHjq/uBjirdOmKbz9eGdFtVWVf2Fb6C+WFDafz
bRKtEyPR3LAQGAlfOUVvAPgJ6glCVHHbXNkfPr0nMJ/n7fjWFSjaXby1HLjOXY/m
7+7mad7pM+6r0cy69ZC7EDrSkOXlkbhfg5U8ZPmjpUAZX6mg/nK7scPvF8vac4NV
0P1ZHnW87xSIgQlBbeuIqgdmh1fPzvkorIA+T5ycolvepFrgOjs7OAxJ5wRwgGXe
/XGQUl0H/QHJoG9sqoyMKIEGfFjcfdp/S0OxxoMoGF90aNSTSl7RmcfhdgUdVokb
IvVQsmMOAwtVQilMFY4b2aYwRG/qp1XOjrp6kCyQ9BGfLRGf11R75RtsOVRBcht3
V8tcKLJYnLB4BZv2bMarfitWy228rNV5a20ZyWlpjg4Io/HMwwqxchlOiJmkVBSb
kUyj9x81AZQBrDEoqE2Z+0BA53cBTaWvaqgcD+ntv9yV4pyLcOl/y5hcdRXvgvIS
5Uff/YzOgVO0ERNwl5mXN+QrTp0S5vviuHGnVwHotbUcZovrxWFfifECtOqKhIlO
LF/TKGKxiJikuMC+qRctNJoWX8d89IJlBuppdmKhctmrepQYyUbpd/VzQCL/wIpZ
4Q3H8aNyzWOeak9yOG7nsQUqwIZyh8qXWOxEzOzvGnGQkd+uvhKuGWzjqee6kiOp
32LhOC0yVELuVh+bHc+4SZpJ87J3YXyYUNsDD+MnY1yCAz7M/bjnPIE79vuZk3y6
IYagUiyh6MlmdVEcrs2+bIEBfEWgW58fAAza6kE7iizwMC/TGOya65exXbpRb3ZO
wKK1+fIKVnuOZzJBO6UGthwpP+3EWmGOCqQBdEVOVwDBAwasmVb1YiNG+LN167hL
tZbk/S4A7QXR5+9OCvOAtPuyRgKdhlinZd/h4/yYFPX8TWa8fi+Yt8I9ruE+LQcw
fWyeJ31rfQ1o15YoEB55NeM+mg+hK2UhHZqG29PD0hDVmFBuvBPcGSoPR1QIfhuS
Ocz+bsglnfVdAWcEMcaoB8tbxRdelDzrNheb92gwL+3WOGJk605sxILF9WXIc59O
sPpbIvUlYq/WJJLKHT+RdCKYv7DP7VgTVQn9oOQyiQeLhfzQZUqgXnSTk04tEbmR
CYgJer3yR0FTSOGJpzdncLt0rzgMZ+UzyvtZDxbJQcr+0AmjPWUP6RUBiN70eQUu
yZCK/bKKAes/beBVseGhvObryTLW4Ma62AgMyahyTfGd0BAvqgAEqWmc/JlG18kO
dDwVQUahvuJleRJvh0vt5AGSmTOky6MUwzo6EzDg04QvsNwVblmtgF/QUAqXWHQ/
yD+BbKVIoZk4t0cWYG6TApZVGGieuihpfEP5L02do/dU2Rs3qsUmEsLuIvNAzDJ5
HoV4EbX96GbJmEWsMd2NjLnYQyvlxSZL7Cre+0ZYRQiWXLgUKn4JZDErAeWy2kxp
kO6llx/X0+plALWD6RTqZAkeeAoArKeAfvjnHe5ViQfJPJamE05Dk/Mxy6lgsiXX
OeruKjYwAFSwXIndndhFNrf6xm6A5Ks1yHUkfruSNAPo/UI8tlyuTmP7fkx2TpHT
YDnd8vWanedNEsnMfu/U8ssUJVPipNLjVTcKujv3JG33HcAbbYUmvGgdrJQst5rs
g8d8rnl/twhla6+M0hlqf+afOdYAqUBQBctbX5mFbiRj+Z77CqeH+vqh1tmC8Y4j
DXXg7M2KvIPAnNlCjfZWELa05zUYOWF6sHWFZ8Ged7V6OU6QFXqC4MIl3flMXn5D
oM7MFx4oQ9pKke2Jo3ExHnd6K6topRzbZ5hA9UtIC/27EWJ80Ufk2YMzFfUuyrfK
1b7qqoYwl7pAj2MELRwwH5WgFjHpvU5rQIRkrYyH1EUKOXOjetDMRTThz46ojF1f
uyMkUwsbMWxsk0JdDulOGUIOvxUhfmhIxcwoUHiRg3/7QyAQQpljV9m/eSspeJ/0
RVzz6nzr7YbhWHFZPF0AeDYnSZpkxp6lMYNMyrBwmgUJq5oDF4PY1Sox/TNZkB74
2XJakt6vbEt/meDBEnwWO3ZURHwjXjS3OKi/lnVkD8oE+AnSgxfUaAApzWzysL0p
nbI3VhJjjhB8eE9qVIITNxTVVB8+1yNSI0P56LjGa0Pp3v75v2Uct5fyGaYTphCI
k/QoBLwt0Ue7Dti+/8wL3+7MV9YJmMlSO6gWm2NLXKKC5HninDVaPzAElQg1CSlh
JMo8lhRWGA/902lT3FyMx13QGZcUB4NKkkX7zuNPBKyp8LiKm8vGgv8ifRVmEN1N
5opxDF8gZgOele0djbzwU8vEKfBomcwhmE40nWOg5Az+IOf4ZDANCvu+TixVtjPf
HNVjiwvvYCbOz9/R58r38tX96vFk1pkoKbyybRJKXvpqI1gPqG1E58urKY/Aw2c2
2/65gtRP3PATqmJLeSjKRwq6tL4l2pIayEnz8tPh1YJ72kRmWS6hzYm8cwvbLZ8k
SGyTCwa/2Jvc5Zo1dNjGPI0nrKKe0jTb0zCIPBUdtEOS8MLFh4b4ENOT8OaAZcGS
zuWsM7CfVyKfIGnNkDzNUBQ0CrM6rUiXuHbTi9nYJ4YEnmt6Z2CfDKAoQNRexeGa
pnYBuvhfJ9kekD4h9JZsXOrH5NXaFGGXjJ3br1sePM+p+saYAqoW50f7hxwJfCbq
O9MJ/eqVpoae70fs2EZG6ka1ILdrWlTPrCDY6Lhsqr6T3KpL62Q5ez4Ews60Xq4D
f946REwXlasKcbF9XS5qoUIBX/mpSsYL/7Kxb+BZYz3P8svKUsVgd1ADg4N+YQJg
8xQDNobzBdMZlNzh3OIoZDaiWXmilm9r5CyIlRgv95NgqwM/znRSwcEJW3bmgrwU
47FKrKUoYcBpBGBRZDmYxR1ZYPgxHL959BesE9oHfHU+YnLt9PWf8Flhfr7adH5s
vyefNzKsgkvsdCRQYhqStW6b+Zi0qKLkVoyIZRmGICr4jklyJco9EF4uY96UVdm2
DcZWFmLV4nlYnPgFBrmdkccOxzQ6RNlW4xGW0kjV2Jb9WYrjCgohadGIs8s5AWsH
whICrzx94IEb0ZD5I8s5rBac2oFzpZdvJgOztVHWPKpMx06S5dnL9Adnw6D8Ebc3
grVXhFWMAepZcRlInOm/wmbGsRtzxVOnnb6v8qCe6BaLporh9CT6Yw+yYvc6flLZ
2mEuPM41ybfe9cueb0rmooBRdJtILoBCOydjU/uQh9DFqEdD1Cik46xZ15KWDc7p
uOQewKVdslP5fmhTBa9/beP+gwQTU60CfQtVsovrvs9rxwSRwqH9vIAHjl2gSaJ6
7jfbjAAhdbypQAw8o+uY2AO2VCtLyF9PwGlpYLHIQ7tGPUIkcywedDM9ZKWSt7FU
GQqET1OyJQF6ZOmCbvODExEQyXSqB7xhyoDRRTd3R9bRCsrPtO0/r6NihkysCnYB
pZ1DEvhmg5s7G9MedXE4wnIYN7B1YsGBOz4IMslr+cSGrtBesxAX/APH7n1JV1PT
dhwtYhRMhqGfAKYRQl0ZRB5ENEZowUWI8qc4mOmqES30InFRdQgVsuSxBkZfiPKY
8A8DXVv8BwFHDaMj1KnR6fIxHFq7KgqAJem8hp89K9kb92eAcJN1FvcKIdf5aCpM
1MqgU+L42FQRBtdISpZLqoOIrpMtOhWrmZG15Tru/o8zFYz60iAWRKLdB+llhVN5
yT5sOTTLC/q3VKC0iVAbxTK8RhdpC9Zx5O7Q6xsszXoJsmejNMmzcAaQnCh5E4KT
icIqpgh9vsn3PXbRA7Nmb8EdsrF53eCCJmdk50Nnl7ME7YIbcWNPTTmRX3kCLg00
8VlWWOfgykVyoAEW/04ziJ850MdU7p7sq1uAX67p8YrddK+oje+WqzA/IWvvrLuY
3CYhfUIs3etQHFWP6dofYsfaFOgvqr6CC4PAUDqi5rTE2VBEojPemwkzqu8nZcMi
cqjpsqWAoCX7LkqLShbjZqNWBrDLD3qHSUbMU+1l5bQdIUfK9Rv9LBk7FPcO9NIp
5HzcKBCjCM3aT5SUarjhaf7CO1lsANTh/eIDbcgpjtG8igUwvbWh74OK05W40get
aO+KwRAPbl0qlML0a8Q2fW795O8VpAJLsxiOdcDnL/hNzxaNUZHxIi5DffCWFstw
gJEjHZ+ptaRh+XCtG094YFzwNrYcY1L/8HUcOLYZ4DBCBHyFFtLJ4f2gJl4X13fr
Zro7h+bWqqN7yNb0VnAZUst0sJ19cVM+q/cx9sWGrzFjAMIEY9tto+scqwDRdE9y
RaUBc8z9ss8ev+SU90p6CqElfGpghw0mKqwsukl4sXdxhfLZ5YI7uE9AghUuR6Yh
sgyGCl6ttPvxXQuECFef6iUvHqTbR5C+qz2BzBmAQFzcbrnJQwBbcOdqP1+xh6oK
ISFWT3Ce0VPIsFf1LqDGIt9g+eNsIZ927/DjMzlDGPn/St5UytajWuQERg4iHwRH
mWA9qW+X3n7a7won1SJd3fx6ndoxmEdOJczKxhpjxoBaoDk3M8j0RGEcIBAnjzfl
zNnwqLcSNIKH4/IgBcipo/mghKcMWkiM0qkq6qg0O5oMsHx9/gRNrbqUDY+YA/TH
XN0L/WDVfv1su+73X5j56kQq+++xWeO1k7/eWHZckQ9hQVYE8491INqbbs6jJwOp
FoW41ZPPqlVDNJqiQlhkZjNthLUANEgsrCnkymOaWs/KM5vBt7nDuWgNX1ukcFIj
6GAPl7bSx8blZpSeFU039rZVVs0aFbX84q3jXFRxFxl+l1jGZTijrN4utKmRFgg/
TfNYRKejXIV2DvG9nzseks1X1D/ZM542zLTw8loTxdM6cgh7Yy7IvrK90x0dgu3i
u+3qEv9i/fH0lArTl70J1ST3UJlk3zEpQEEDg+iUgn21lL+c5wtzBnuhuOfMArhf
lFp3QgWiFbkVh9/+6Ilwg9eehwvyik6yxkrL1mWaeoHMLBVJiS9MVEgm/eObF/AW
M5iL0O8LAr7u4H5IHhIu9Ac7jlNy9L8WL+TNCBMOdI7pAjMMevg8nK1M6X/5C0tf
jhlAQZPdA6BV2di+6n1se63qc51K0N/cmpeWDk/4sTAV3Xkncl7DAK/P9SozNTvL
gqBxcCrCJbQw+rF/1vZpvpWoLpk/ks/VA4KQRj37DEnd79LjKdp0JsYG3o4mPF+O
AaBAYCBC/VNb6bE8JjI9pjCTxMxAxleUTENZnO7PvD1QuFbegnpOr1ulgeF2Zdbr
WGiLRVMIHQqe3o8NQ6qkgJ95HZ7/aFVAa9CPJ7HqXLmcaovak2yj7OwaoQ15c9L+
LTCOBHrW7EA6/RFLJ+Naf+Y5hkwjPfzCOZRvTMoS5UdVP4T9O+6f0IcpwkuD8Mn5
5ZReb5ekpy5fs4YigRqL8Fr4ZVrsZMaxsAbT8NwfclYKVGoCdvmN0etby/wWc2nY
ems3wiABP2fN/BERi2m7aLMSjpPHEk/H7Z7GqzEhO8RBWI++gofLLvN8yl2vIewd
tFQRLJwPsDDfdPB7TG5wdcbjYTr4PozB3zKwbvFpJsgqvtUHo6Xg7r/CzvSlA7bp
OTaXx4ShOfUZwejkVq0P1NyiTXlm/DOFWwEiHFfnae8mUWflxSUYj0Z5jfT6HHFz
FvlbHgwFoy2EZ0+f/GmELr6863+sZcj2B9HVgxUzagPSuAvuHOQg2h/9fpC/Mz7j
ROEsR/BFLbeqU86efcErJ+A/Skx/57Xcjcx9zlLWEblM5YeAmnR18jjOVcVgd1UT
aKm8MJVD6XPQtKrI+z46Pa9bwdhGf/FVPvNLWTWsO1orX/FyjWthzIiqN+OcKzYb
dUrbqsd5RjgKgvu/+ARjIZcodxL61A3QiWu70YkPwJTNhIthArQtUWZoNQ1ntDNr
ZbIQLVka/h/N7Apb8kvS4F4BDUQTQt8SXG2hv5LkgbCwG5ml1KPXKEEEIF0m8b1s
ZQDYZsXSVp9qgXM5A5xccgUFC1VJJ5AwHX47kNxBCVfBGOOZhbMK1+R5CNHBNhiA
nJ1Z126YPRD2O61sF4W20QBFhQIacbBmdYjYPmEFQHJEiiZ5e9jb3jezx7dxcfF3
939LObY6igmB1T008rtnYQJiePWSUWLOG1eKludhsmG8xjIYyxZaS4oXY6MQ4zoM
FWQRgfOvFqqK91beCGOlMz5qMFggU7BKgBSlryZL1JbljQZ1fVlV/QRpVaJHKxQ6
EIYc8gi4tpgxOZ/icQgYFTdUZiIY27YhTyPnZetTAV5NONLP6pSruMH5CPaRS99M
a60Vt4d1PypdtxNBsgFiHRYWCw65uTU30Vm1eKDXJvUXAjlXPssGkjQVOedX3n2d
AM8LCgmNhdR8YlPAwEQSip8d3iFS65qBkrGVU2hIdrU1ElIWw4yxFI5zgeiRTHts
chrS9oHTMath4syHG4bOBR5sMnsQvXFU7mLz6wUYa79uusjVn4b4fa1Z2HEk+6bc
8FCQgM8fvbj+0LWJe+J1aivWodyuQ5wHKPkXpOOTL+rVDe64S6Zb+FkXXazw5eja
zVk8YRmmQ2Sk88brK0k69176ZI4qO+6rcCL7CsSp1qQhyoqOzNZg3BR0pt4LOJuH
PDQDQG++sm+6X4cLpLJjpBOJ745L7FVoMYZ2HJPvEuJbjz+Cf+AwpP/N8Liq46YU
bdzjCo/CvgGiPXM1o1A30GVJ4OK8Jpk8y1iHrSYrWLy3lqusG7b8WTBGh2xBdg/F
GP6wrK2IhpHt3s2hVauuh7nHEidc6LRuV9IU5NQs9iH9+Oy3y1197otnDFZCFgtA
t2XfyOqIvH54dOtk0PZguiimYJ+Hw4ty42MBeEZJ92jEQ/CSaRKHRXslYacDcMsd
DajMd2VUiWOzZ3M4DwaNKv4Al1ps0yfHjHd8lidyDLcnRk8xxsNNcS4zwvAZAJSn
9XDVqIIAl0NYCYi9EAXqypI3iNS7B0c2S9vx2neHeXZIbvcj1CCaDyO1IacXZuiQ
d2c8PAz+jbjOkvKpvq/oZaVcweSgHYOlKOyy/83hVNmphB1Fs6/39Gfx864dfTHf
CPUU7QiMRxrEJOAA0luA/N4p7fO6hVhSp9VQ5ySAqSWlsjY2I9/JWDP559hO+UZg
2qV9NBCYfhvAnAsP+kZ21hWgipXsGfSNP2+rWPN8re5Cp643j2VLBTFKxWtlFMla
xBdUgPKBjQPBGWpbND32f4EWVzdrrueqX3uW26y9GbYOjqOo3y6w2Ko4FzQtiQnU
Ev6cLGQtA21FOzy4sthe8JWeMzhA7EzxB6Ca2Rj+LuRElEPACYXeKvLdvkqyKa7D
VPY6m1DgyILtMegvq5ZOrgcBIJ6mC5g1oYmqdlnHNAudKPmWpU+pmjbow1AKLYVz
HFhmWMaFlXwvn8YzedIu2JzJeOJ7tJOILUi/GclBJ9PMjD1Tv7HF1fw8DL+Nq6zG
ffn1VvnF+gG9msAzS4IpoSWCDI0mMK8VICE3cphBXzo4ZmUbdOjAyzCN2mKX5vK+
YqskEagpR+74S3W0nQJ9Oo325b/j6m9/X5BzL4wTK16uaGwZ4TVA+wze5O31q/o8
AgxsKVsmwXXAPu7kk/jPu1WEImVjVtmJjdPl5XFAWlEse/FvpMxa+esOr6iffN1l
ArVYAHZ9ECcehBCuKWP4CIhT/AzNIauRpBsuGQw9Nt0PQMTCFhqB2zGrW1aQibNO
zafkJBb6M1lNLBZCFu2g+lFTq1q9W0D190pUSTyqyzHiN1eo9PtU9zdni1RU2hu7
HWPVFgsHIi07meMI99klYdLDA0tXDEUml6XWJCwsbzG/P37DQkWNY9/ekfO24cBY
7mZOAs4Rdp4d/DhWklCY+LavbR9Do6ManJbw2erfwgwtph3V5IeY3ufaAbpKtH+N
o6tKASBqbKy1mbbesZkB7ix3hnetJYnosJo4lKcY2BEFhefaQ5pY7zS958REiZS/
00W5QcVfitJljo3cwA9P3nq0up+A7KhSMS+RDgVreuXyJe3GARhPAkPmV014qrpY
5c2G+OyoPpCCjiaqa6g1u9nTvVhwI6V2Qxz0Fbu/21CDoOj1WymE3wMtJ2lyfHvU
qnlxUKZ3FtwNdFupZ+ig+I0RCI24AbWQyYOzLbsdlSuE+ky5kP02eIT3e1Rm8mCH
BiQZQ7C78Tvco4Xr5T49G0LFmcI5bbyCSzlUnx6GflLdKOTYA4JTNxVvWuvZzqoD
yhFDn3IQsfXzw5Ab9U1EisvwRfpwoaYQcclbklg1Dt+SkocxKPPSksic0WNPf6S+
yH194JJqqH0gkDiuo7IAKAmMyf1m+uAWcpHIOO9yx/B7WXwGL08+G+IvbQJHIa9E
P7tEMIuOyIp9nHLDeGfmmwZre12M4TTxbgY5mR0PPuxbief17Qbduiqxrvstr8FH
Uy1oGmaZPtrQytD/+cVwTw5CIIkiKIAbCP7o/aXAkWoXiKSYgqNgtxmF3v6t9Lrm
aLDJSk5AD3STs1ZxO8/1f781Ca3U3zSwsfoV/v3AEnKpN80i2DrVGLSXLqbSl1oM
JFiKLorSVKTP5MeOdUTtgUQQ7bLx1zYCzgsiaX8ZK+hVuctA9rZBrDJWAw9SzWq7
IaHFKwmA38uZEsEFlgxa4t51QLZ6zg7tobhdD+zyL3Xmg07FS9OoWcg5aYdqzC8v
CgixDORkv3b6hNfnDtMgJOwQ32JNUdNn7m21WBPT7lqOhwMQXJdy8okBoYaihDcG
VwWBQiwupbgjBFUhIMj1wN4ASFIOvrfrMK0fRGM129XVXFDSn0qbJuPEd1XdRlmy
R/Lq5xWv1UfTEbjOkE1JLcgsQZTdmBVlGM56DMxleQ1YkfkOOGPJBHtH4JciNsDD
9GM9DIcqiZ1m9kKekiQSUX70TgQHxpjFnnLUh3hGMl7ZvO+alxY0vZQrH3S//hxI
HrlujwgO+8ku1iz2mEy3+c3Pnsk73zn6Auy5mMX+d+71nWXJ7/sax7qTUU0BmAwj
HUJEFBDk6ICGU+wFqpePL0PAE13akDuo4SLdV6wbtlYy2DuPCGKviV+j/x5WCnec
NTz9LTQZW6WYh5WjjEezCUDwcOWMXS/K865kCHbCZXU8eBCfRaHqLDL8B9cKVDzy
DFGB8yzwII4Eapw4PQkIJLzjpbnuvs17MzAIW+v4KPrRr1PfzA06IefWVLbU9o3g
meLNo0iZdXOjoj0kNNHWqi/PBLAKmha4oQKkv5vZACs0aKINq9umvi7Pycg8Ozdl
ZavsmKLs9br7FmkmNA/UUbw67MEt8EJcmdDzuoYRmRnoVaAC2mrfKm2PhPmJireA
m/yINJ9+RCQLBKlZSj/6sKpOp7Q0LGIgxZfQgfJzONf6x7k3Very1ANRrqAIm6uO
mp5Xj3bVRHwke38SYST2P3Ipk2DGiuo4kpNx01OuuWx44w+ucFrAh/lhYEGQC7JG
TaHB/1vcklVPQISLM0lUHLXTjVhwJB87yLtCUcOcwYV7Nt48L3n5jIRKwDbge4T/
N+ZuAgKYbyaSmo41sOti4YC0mQiKebqZUPMom7bNX/aBXp074/VZtLtLNHAyhUde
kaHcd473u4l2IZi5QF6NriiGPcmTDALnNpCG19zkWj7gqufOl5FMG7JNrKidTM5C
oPnohLudDvmFWOXuLTVhxrVmB3GTMaSmp2AdK4qtlb5YxqLYmgIIXDYSoriXEjQ7
zfsPD/AZypvNoFeTX28oFRXoe94Gqag33S5HNPmklI5YoiJlFAsLaKm5DjaWAWmI
o32jnzbuSohVi8SfNImLGk51HLFUZjlWWD/zQGfHx36tQevoO57QO1320UMU0bb9
ZhV9g+7PGNOJ2mbnOqXiNX2jbPJXv0iPHFW8+a2h08d2IbwN7rXj5wEn85ea5EWt
4UB1UZlMudR8t4ysnYF3csfkRp3mkFz5SLdQiWXakzEufSsAxT6bZHKuZuJ3KHwc
YwkyFV270VdCkUImxZUWZU4t/zh94fkFhR22tVVZm4zcSU7Pf8W9MS6VPe+IeS7L
zewtCzoHtKl2SJmrRhVl1IYHyY6Ydxlo3rRXzg34PMQO6CnnK+4SwHQFhFLKB6Mk
BePbMaK4p6I3c7k1WdOWb7URgu0V2uH39CTUyhjnLbjT6dnY7MUnknD1MgGNcebP
LNOUb9qdRmAsd1cFFc/BzRqb/PKTLu9m/0xWZhChoJIyqgonxUYc9mtFUq8HgTgN
c9z1Pwy5+DJsRQ9RPNwLfqfw76WpNczdTJ7/1hOMve3nYcI4aGlWp9VU4+ioXM5H
hafQ/VZRTO9x2oG+nUliPjNj3SlPaj7cQPK9fD6MHHtR1SSmFk2D/FgKoleyYxF0
14XsunOiujN5avkYdOzDqIshioNLcaWQrnOzqZHOXYkClfbHRLOhrtx+k8dcADlw
9PEd8SBUyulbDm1DYNVjAD1D3nFj2H2a+jABsife4RWcA3w69xSb94Ob31GwaRsr
SwENyUYKb/86eGg+wTFIksYVJlfgpqsP0QTBHoLljugSzMIdCxATfc6tpcnhad9E
TEOjYGHCTcdCUMnmgRB4jlqE4UtoNjJqCL9fcKGJrpG5f215DbFuCUWX8pCKSSVf
4maXyIvMvBWIi2nJ78sN2SGsq8dNLE/5MG52XjzqkuRq2QAGji8eXb+9aQv6f91/
+/GstmrvpBzm872RwDRtYajHxcdI/ITNJmDPUtvN/Jd6EHsjwHWPhudA3waHNJaF
5rpY2/Lch4KXN9E5dgH2SZ4ant6CfXaXP9ksbKHstiohGxCoAnd49ZcUCp8guLpn
nV8RRaNgqyrOnJvGurMKRtGcIY0KSK8WhBiq/FmrImod520V2lpN4u1zdEJH1tRD
E6nR86gRXvmJ1Vzyb5ZzrkXqMSDSPpRAIa59RNj4GgOwRZmkRNGNdaE9HwsWPWSP
79kTNiqYuGC4ScaOdrPjx2M1Jzv5H31WKVG6ZAkLnQ6gwgBaahav8qfHmtlt+q8Z
eZHC3cq75TSHTOA3TRLR9rGgJDsTPxEADlOgwhJ7pTMraRPWnB04CJhaZ3XgH+cz
7+vRaP+NUkmnI3m+j940VOGhwsBPQxDehaTkoy0nhdYL4adFVeFpwWX4TGpMZ2PU
RmhSC2Gmd/qIxRi6z4IwsoMTfRvnwM6ruMAP9F/OqMph7NOvaxLrOlbcnRAsm4+j
SwiKW01d2KAh1REo/GH5dB3spU5azO7eq6XqL5h2/wZOeBZML5CouZDZWMMpttIx
e8zHMTHvEy5q5PhoecBNbgqq9YmcjJtaQ32hDCV5kd0Qvs0vNqjFBI+mMEB69m52
rx92DgEFwZ0r2UVZZ3CjLpfvc8XUWxDnMcA1auX5BqIQUtiJcrRsRmoFYE5y1FoD
rMLFxUziRmGSGwmKYAkbQGBm+3KEASO1+6gS8QeHZQTAnYZs/JWM+qyaXCueFBMQ
35GFMiTiA8cme8luPJgPoQ0mq9ItGpMUL4H5i5k58jjXpJrZaWQ7IWDwDw/gMWzQ
kUQSbnB3uvcyfnVtAwRw0WGQAlyQ0JHDzQ23FXeOoSOSRPtS4I8EKQ0412gnCLHO
MdG7tglLM4iDN7lBgjJapkNfmucN3pHZ79ibz62P3vo7hRuWOcYh9F1+d71XwGwB
vm5Xj0ZzScSD8KmMZgyUSjsmw+i9cSfqn8EvuVh15Ppfb1nyqNSKvVcY2qjVR2i7
b7NfsuDWgwBKD8CDvDHrLWFg3KnSZeNWY7EnPe26nmGWI5AL1r9g7n3SDDDhD7+m
hetc82T15y/CWY99HL5+Wqqk8TfkWL/sS43oay9v08dwHUlSPsZvaYImbWjWU0pp
B7lLKFT5vBL1R8J4Yc/FFcX2MAvdC0YzG00tNhjAFxWMolKIE6lkAxCFlSTBL51h
EXX3LTQmMdbzcagnV6Vr1j6QNkuyYyBzFxQObZq5Or+rxMUVDrualoxExPi8ennS
0/SPU5GLpCf+Mf5B2/eq43yeZf3w9lNGO8U+zdC0PKZavmwL20X3KL65NP2h+smp
u5KzD6P0SPcYH6N+TOtN4dWutkh7nrQ3xKeoHz0geksbrg1dvzo2NRNnVy5xDTaB
cltOj/lrkFF1X1ijg6IolAGZ3O3beH/9xgtaWbnP7ycGV8WJ6xL4gx1hg627zVS+
Lnve3tnbKTXz86lUHoL7nLGoA26pmEPVSYcbQizt4zHKJjTnI/UirA2Q9M7lPFbd
ZVst4iJn/fsOwspo5kHKOH4wtQLMW1IlK7bEJc17qtKGeAquW2xUtauKd8QIJ0rO
osBljRl+XY2u4S0at989fQm/fyw7IkwbCdY6l0CrAoF6A09Nb/vnVg/DeshYyz0c
sCxH4oO1kSEmIFULQqgBdljGAaSGuHG3J0pWXPOAugSEWMX95hD2FIn8uKJLyifj
0sjMnAgum2AfgExNpEFiCFdg7fq7FrR6SZ2cKt/w5MGO1lgESvoIEU9Ra0/mMz43
7MQzB/dmblqf5r+bnWDGqffiBubJfjK//8EoxyubK0kW1185kk7abaWriLFUwzP4
fYv8IsgzsbUxjGL3QsCgrCP/Wi+b/56FMvj4lG4C7DZDQWvtRCG4C3+cehiADgJk
lCi4lUMIhm0OLDj03H+traedcc1L0kc1ut6KzX9iVnvC9cfbz4W9WHCVzunmU7Ma
QUsQC08Ptq88kgF8f9n2Lgn3R9OGVP+KBWd1lpDfnCddtJZz9e9bC2lHLyIZN7QH
iAXTRXiDoPp53yYwgR1IN2Sn9GAitcrEr9h1BrDSLe38oyns5WmnHIQQxcUcxSSo
4sd5XceUNfptHxsDzHsyt1y6xF0ba5hkTKvRB0I8VLs7VALCWhubAYmFW36LQNvI
H/iujKFcLB9I83pbEgRhb+R7MeaLuNqcjiNZDA64RFe6kI3hEAnDK39+42gBYEns
bLdKh9qdD8Olmg6iHmjpxchCs/MkaDNvErE8hYW2QXXlGDrasJCNFgW1VW662P1E
vKrEpLB/+tv0jYNEojZJ/rMELT9wFc+pBOHnxWthboBm3kvvRulAhalLl7f/4R2z
arHNMHuVg0Y4PvU/MFt3BpyxXw+8c10HmnGulunnHG5kR5k1H1pXmmt3/lkxJsr0
W1qUTFkwL5bQ3/ySDSOPjPPSScKrUEaIhX2vkzafFirc1qeK+3pawn9UDztFLoK1
BcCGTASYmN/Md5aADWyvdArmX7O/Nj/U+DoG7qIFEnh/ht4yAEhqGXadVG3PIA7Q
TXiLRf/o0gjABHM3wDN4Y51SHZvn3HjSaJRgt+DniwM8tVM3tx2Nf+WZrhPbnFCs
RE1QQCvU3by5EEMv8TKGgVY7YlnAvJ5VEHJODhFMvNmGaxQ07hDFNhAA7Cj19NTm
FVToTYWEsfKGMeCKSZhMKupbehEoHq2v+NaFLB922SgfcQIzI8reEsPBxmJtgvVT
0bmua631kq+Xuq8/SzjJIh0Gb17UB1+6zCR170WtBen0QkgQSVvL1HxL0yh1OrTT
kM918SvpBuEC66PNm5ZyTUJq0kmLgNOuEQyAj3ACJ5B+xz5SaQW7LPIiTXQG3m5Y
muiH92UhuD1bK8bdBigrb6vt6ht+sQpnz3qMyHEfJ2MgUugL3zqBQDo68TeztGRt
+O5fmh+w3zj/ypnBQkvxiJPiPXUejkCV7K1NcYA1MY6V4lZnKU2RoNiwxtSVgBpB
tkQe3/sLBfB1q+m8Id785z3pvygZWkabICRKUT/xbHlp3JY6oIN25wkVwODIdp8p
2E1BJlUyCbVdEEGm38+Ut+rn8FWIUjJJevu8QDx0JAljWsxqck7hewJeJV3H+Y6E
EbyD1tvY1vUQs9jDG2jcCul0FXF8fOMOOuTcgQtlcorbZL4RO6uj+CpvIBZ4VRtV
HCU5oAPr/e63i1akc5uxmJawhxkbqG1/iDysJfNoge4b/TlfxoRKGQBBHW4MLdSf
HcZRwkcFI03zUpWIegiTcpj/8IYMkBwmZI2fi47ks+ehV8Mwbq/Nv3ZyDc+ScaBR
Nw+dSm6Dq2/YGkF0YLqnXbmowvozhpanU5yrRXhLbmDYJURWfcreu5ckj344B/TG
3m+olwEc3z/Obo/6HaBYrWqGyKF5Lai3VFLLYdgM18hG2lYa+2o/boLuoVJy7Ji9
o0ujtmoG7AjIQaONJ0IQJJOR5jZRkRU5PbESmmXsKeDDAItUlNN25xBoJ+2CvQcK
VW+ad/9MgvS9F2ICvKma1p69LveUvkD7Wxci77KIF2T9WM1/pEIui40Pfi5L4uSW
5I2JXDN7KE7aSRumMkHiqsiKPabrAL8PhRotHgRvEe8jTBL7sop5fo2GgAQXgfIe
7R+Nu87hp+gL1S6MbNGSt6AbgCfoETaByHJmqhOZRkvR44mlp+b3dork2SZ+iIkc
t01kvF+QcCzJByo+uYAtOWyVb7KKCyuaWV/K/dMQ++MEpEpsgI8Lpk3+ecwam034
nfIJBQr2kN0Wtf8PleP3JhYF0qL8tzzel5GvLcHJOJgaU7uCPEc68EWox1VThgks
PSo+XrMvvnRFP4wrXuGnNXSNYqcmU1shhfO7fCuhShrVwXzQZAPN7b1n0rA0feuM
uc/xcQzFBNildDkUsVKCap0wVEAzaSHa4lbQMh8hT1Els9g36WYu1G6LfyKmzDqr
llj3riWprtEkxCM5sHXq0ZLujFaSajhmZnmWTxXFHMx3sRaMaqOgVqJLNPOQJc8B
2mZ5FtXlt0OEbeIpSais4M0rsZVvsoE5auL9rdttCtcQDHEOQ7kzQSy+uV2vtCt9
HAe5dHAEUVTldUHTxfw5v98XzEFwjPD3qtaNz7q3PX4M8OA5rT7iMeQwP4WAzw++
Xd1BatAdU7GPwBUhjI37jrwBJ1qQwJ+qS4nLQk3fstfcgCn5PFGC+d1shZaUP1ft
5eQwrgRFc1qIhRevZLg5eRdKH/322ceLnlflFiyVXJ9lHX2UxaejRZOrGMcIm76A
Ou//13biHH6skORb/5ZAWSEfMsmmwk97eH8B3fuu6LLgaxdYjSWG+AhErS0FKSCl
M0UcmkptyKMoQv0a/xz2+Jv7g+UpJghdFGpSEq5mAoTKFCfvGscCFa0CyFEtBjJk
kF3WFWb7OnyWdYmsr4TRiWe9/3xtptSpiqqbtrePkSwB+3pRVBlG+Epw0wLvmyF+
wc+ffda7CGuPvg2eKOtSo6cuXzmcYu3K+bQiX1Ctp71X7r5V2uKPQFGTkca4HDTR
iz6XVIohN1gVR3GLiemwp/2jhMjuVbE4CHQaQC19ITUwMcRtORrhRfF1apj7TDkK
E5FiCgant6aZybDnxAtPxQjwQsAw6q5woRBoGNcyTVRQOzYRfmrN8a6xRIbejqwy
JJIijvKnM0/l2O05nR13Fti4aZnkkD7+S8wsINSl5jIHCEDO3OBoUvn4DogLzo9h
EczzYZ063N34mEq5DYZJ41X7526rH/2XkN1QOT8RA4kRalVsHZ8CHMeI1Gux4UXw
tIHGfysOezO4LLXmDzkBH8Jmjhtde+03rtiUfAeSTc96h+i8RQcpWOZcw6suVEh+
EZLjmOP/eSuKzQpe8+VCC1AWavCuv/bqhSfpMkxb9lXO9a6sjSaBtxu+MxVqe8r5
LYS06BgXOLZIWvjtAeq5eGMq9KqrfakgIZpZ93qgiKapLijr74WiM9J7tJ0zeiwO
ncZ2W80vfI2dAlsXaWDBdtlOQAu+ZQjCqQum1nw9pnOwU44qqq5fFk5CWyh7A9lo
5R7eNesgFNBo1/tGjtPtpFUMut2LJaho1JWlAJsR13By0ZhHTyF7GGb2njuEEJxB
X5QNYggRSRrM7dYjvhGLfXI9ymlA9C+Rq8b7tFkbIbtXq+QJnvsBIcMMiGuWZnqq
go62PbIGMSvbMIpBUGYGfAuVfpkUkHB3xAO4ZbphEib2ZMaFbJtKirsc1iuQOD2t
XXEQ4CC5hxIpH2FkzWyPjx1CBW7eVBdJNsvQ3Eu9UvqMlGlU4ijx6CIr0yMOl8fg
L23xJ0gvYieil+txzjEfKR4cp+Mw2re5lo529AcBqd/QpPznuazI07qoO3fHwyz4
1BP7mpyBGfGyjjLVllDqGKxjukJYp7m+T2PPH2pXl4NVebm0r53pe+w9yCyXyRGR
knEIMUYostw+Tr5rftSN6Xq9dunUdnZTs8S+ODcdErNz0zejCuXGZpasM9A1cyAU
+bCUzXjsJ9VFgeG+nGeEwqGW1fzkEvBKJv4LS37qgyKIrQBnBlb6UW+pePs9dgn0
KLhNTXDyXmJak6ws9Z6GwTnG0O37PdnmzRVcOYgIGg4MR2MR9J8P4OdjM87emOz9
gtnZrh8U1GHvm62mGeGBetlte6eD53Hd0gfSD/LkE9/DEEoU8yvHBAkpNRzx7yus
NOL3cZ83rAkQkmRIfg5DG/WhbbedKpLCQ8elU4wVSfeq9Zqq0/1rk3t+z7PesG0W
Sg3ZGVE0I1nnh3UJLn8BcjehwN1f7/WmtmL1xaDJ/tC2jV8nhZcY/iIZ8jHbkMXh
i9bYKCP0fvyxoV48HgzHZxa17KVHzTuVVucnARow6u1JLlMnw06NAJ34yEcpwZ4F
cCLmp/3mQmmaNinX6q5qBA1AymXtXKsTEjwOwZ+Pkvj1bqmVBWJkYb1v/3sKvuoe
GFwEitYBPz6KQWQ028V2IYu4o4nOPeY5NMWo5mH4q3YMByVWlWiPkkttL+fVjUBP
lA6Ku058FqHI1l2UTqg6lmjDkm0YEmzM7hT8/er7G0oxZszpoB7T9DEg8qmqenQy
pvaS9J6XUrYY/QpknNlCOEtTXLN8KHY+6+L15cmER74AO6b5tnrXiRWoekVTLors
B8zTk5VxnvBcVd+Q9uDLzm8MjQ3yCUGLqD+MajToPibps9+e3lLlXgRVaxI8JaCg
lRvHYdAQ0igbgPEe1b9kzxJlIG+SpT/pcohNBa2nZKFRSubLmk31NCjREVRbbTN6
zF/2poVFCWeI3nXE9br7YNfTrRXwoGh1TRVlUObmrv2xBlhj2CBVnOJ93ZhVykRz
y6EuzRPtWHtykTfqWB+2/sm6kTefTX77d3e5fXRIIOa3YIwxKbD2XpNOf6LldH5P
Lj+VL/6uGmbt9GOFgqsmBhZXUBC8h+uDi5SQWB4mnH4nxl2ZkZjEob5qa48dVAwU
ZHlIUo/XtGCmaDcRpSvkzsjtGfAV+nF93EJIZMsVR4NyZHNwP2DqSmUb7uIM7lOv
YV3vxAk/AUhlmEVxD59YT4UmAX2vGS/tvkaOSGC/TYTeHw3LBiON4GuCUc+BVszR
y5BOChLrvRerCByqiRFE5aT80OvPpoGQhXep151q2CwugHxcjKailAhSWUnc7b3L
zEZUFAL1m5Iq4oq6DXrrh19+KoMcmKFH80kEdhOKgDfFVftkNN0ZP3wkhlBDnTKy
RqAnuaeshdZKWVnLsA269w4z+eJR63ZVhuROV8yBHC4SzefWopUIYDRGnUsV3YoB
wU/vTQWp08fIwmyDMre5CJ7pLFtYZk3gsNn72Uu72jloKQRqkccfsy2UqhpfhVTN
GcKlt048v3TAznhTrJkifJyHyVPPKXc3xqsKfOE0xnlfWaHMk6NUFHkbf7RnyP5m
YAhZScGSloN+cfUzQqG3HZoU3fSYA9ItQRnM7jQqkoMyy9qh0Ie4UqKj7wMN0/rT
xZuZq/2f9Z1Je4jXYTrsriKOcdiYB68+paqmgxVHgA5bs1PrqdMWBVRvcgAwDyxR
rR8MK+ekuKQY1IMigLBu78qoGeStOHKUf/fyhByFD6cSuIZjPWabf2TRsSCRuFo5
51YFPfRjN3JElAOEz+YGqWkJpf+BZmlcaU3YUBcWkKUzGJ1UqdwaoBRbMPucKBy9
rhKv8Cq72yOfgnYdKh9f6SXF13NeRDfdITJVdoUio444mBF6op8JIozDrhgATBDx
thfvusInD5mMWFXTySyozT8nbJXz6riPDp7hLk4bBEn4PzIXZaudTQFgdxW9+ixv
72vbOMH7kQLs4kF95P/a+YvTkX2HRfr+s4x9xbLydlEEQXkEUkyWjI2wCcKJ0eAa
u0zZ17DUHHIyfkHiPetv260qyW/FrG46+Zb2YPpxI2M1kHIIrIgtkkXSepRTYkc1
XYOLl6xiJpkVsHy6RXzWXGxLGB/fn3bpWgp/xpybouJeZdwlthOxq2xWnk7OEhhB
k4HH4WOPtHYVUpvbYgc57dohrUZnqTPg1wLB6cHe3GA+ANB1p8mTEMQidCzA7Nuh
EcLXvIR/o3QAwQPe/H3Rz5C7cDBwH6dgd0Ag/qzycCMB9nEanu4mOSJGheSOTEEF
AgrKqY5xRB9bXesAVVuUkMn+2an0q8rDmYgI0rfoFr2ZVxMgZ7D+SQ8RXOixa2FN
qnitZgxQAHkwXY7y6jsMdEGtbyTN1OgI7QiKxSF4Dkv6U+UmN4HC7GfjZ5+4Mj79
cYUavRYaeo/8l6vU2uruwqAd5I0/6TsmCD4EE9UWST/7cTgQn4tE7/KZ0g4CyA09
f1nNhB5eSLK9AmJSK6GbSvJkhTox5QdptFNsnUABe4F4U6Bsxbp5qJFkB3KsHYQG
bTGUZMZtbh396Zi+SsHVmmRA6w7j6IwKoZaZJMZU9OvJDtbRVP7itIBW9VYh7AlA
hD+1tcNPt/QbwMiR7q+W92JKwaavQ3vEBKZpx8CBtIFYKyhQqrpySFQ2AopJZzTh
b/Lx4RNCx967oF+lAIa/ARLIjlIHZnXJwE9xlH8EwGpGwytYyHXzN9IhZ3tOyl+x
Ur1AhowjwGgUVSYBrdSWXCYytKxQtWhb8ZbidiacfZOmTsibGpVgYidqdcnY/DMf
P10gyD+I3uJrfRuTjYK9Y6ALDcUTfDqs9+reidUWob1MFznB6dx17d/YoJi6a0w5
//zY7QjTtELr2kOcImVo7GWHoI97TDr7A5iwZmV48jyWaDfyw9FVzJKAiCv/M9TO
EnQdNYrp5GdFi6JY1dotqKul3x1BU7pWWfmTuFLfvJ5w8TyCslyhrL6hVJFiNxRj
z2s1eCP1xwLpt+rmM0iM6TiR6c7Lc2pxZwPe0jfMkhd2lnYD2tGWn/OpcZIMrsKs
nccHGrck0Mr9WOwb2VTkRMWFJ1Wjx2zo0NAZezq3/bS/LKMTCMfshp6xmxwZsgQe
UJ/aLCuhD9WmJlc7tzgsTP2yXjr7QwS+SCJY/7/siLQedItOsksDLRAmiaYndg35
roGhR1vRgglb31fmWiVfTJIYMAhrTA3BUiCHjrJAUqhEibyjbqJXrMIZOxEVTqZg
wlaFHNQwFSBBjr1Y2DGkj5FsX1c40It+jhoDJjah+ny6YfXBJyDW+6RKJzGdbG51
XiPR7gQMQzJ56wBjXTLJpB991EM33lCpJgC19gs7D6J/No7xSD5Y/RCP/MoxeUcv
173XxVPuuL9EnukeTw5gU4Kd72Vshtc+dAWdRtN2MZAv3rrxfLAz2oLac+PupyEa
+pOPB+qGGxFJLVvFOMmCksDM3YNYI37KRHi7fcciZh7l+RSTbCrrkWqfmptmZLwC
Ed6fFet/uRJWvA23j5Toa0AYtef/Etfwl4cf+QxQS54Ua3toE68mLmXnx953sraQ
saHf/mt70hOjp3ptCMc6vuRRIT0DaVPRd5EyYlYZd3KmsqNi+qdnG/9w8q+9KY5R
o3pHJGWuKi8BJwtjqlw5wdu1KknUDHQYWouCPISoQLPtHjAHpwAcF+VIH+x/TeKJ
GO3GnFVQesCMXEhJncU5VSsz/FskGobw8a5eaiHuHskBX2ngo73Z8us4qbh6MLac
9C4Ekj8T8nf6cyCbelNI2om2yAGpUY7/QHRwPuC9w6Uv+96syDrbEKcdWt7GsLa8
vmHvOPbxclFEfZW+HdmoKftQITemNJVWStldpipNrFMZOsfmFvfXvFltQN54R3oa
fu/nevXl78oxLiCGBj+3CyxY5EWgoHdMs7BOsMqskCrb29wzm1x0+GC7a9/7ZbBY
ygosDpBLYAGE1C4CXtHJ7805w539pQc08Sul/j2cZah2r4T8h0XfzAcIHmRLz08w
i025ubRJH3nrTV8dpBg2ihhKWDLLj9gRWsmc7LQR0+fq9UyIm/mn14tADoBRg2B/
SrNvUBvk5YEvRN6G30djpZwnKPpfZLm4AULxyNJH+wo5zzpKVC1qvpDp3S4Uem60
uAXxH/FglATTYaAeIwokmQiwVhRMFGynEJRrRuLcQnRV2bX2NjVBrA3/6y6aK0Lz
qomQmj8VxmO7mfY+3kbCjXiQG5EzqqgSVW1m5WDjxIwAnf18/Rt2imMevTamcvge
6cP+Nm3t8YQIQFNi9ZcRK7R1mopbghaxZdSeA+i7KXLADGDvMQXuIWlYojy03Ch/
x8gEGar86vmMZqfatyfVuA6EdJ2kE1/vl5vui87M2JIezlZdZzzqOhH75v4S8GFk
jOHI/eiQrJFpsyuzDLBp3OTVbbKXKydYpLxEJG0jsAz+Ulwn74KPIC03FWujihVm
dPpsrEEAWEMfGHkzdHZjiqKMsMf0c6aeSenLsAQy/ZJa5P/dX9819qR9FbkgPpI6
LHVfNRPWHeWuNFF0/zqR87XWlTv91RfHsdxXJQmYvJuY1kGxGARv/dmoSUYcCMAd
xq1TgiQWeyEEculgbyG+1WKZuI3FAqv+GnJeqEyZePeS9VYGLPXzKCkxxaXu7AtI
Sqm54dfA6loE0J4rTYK3pqauCThhMz0/P+OOMSxFxTQ3f57RVDkl1gCrY0Fifaud
wJdVGFv95cr0HKIMAvjMTxqO2bfn/HHIfy0fYfc3CRtbFfQIbCJNACosmUiOrcfA
SCelIO7KZkKDORIi63uvOluWw5EMKvpTC1VLx3quxh7J25p2iGcnlPwoKPdIM8Rk
yq6exiCY9Ww+EjLE4/YL6O9Kb5MXDnFhh0g3WPij3sqjG4YAnndb3r2hMXdonbQv
r1ncsDIXFdbxHfJvFAOHQHlTJI5c1xfDgLmAaI+xLpavpgXMUx17dLwCdfwZNbMj
j4FEmTcpOmSN6GybG/xJ3Th9Mylvoul6c670L3RqEN4KJgtFPhpZ6mAarvK9wcmQ
CyowuiuXJJXIZorEbN0zWZ7fXLJdDShGiRJQtEU5ezJPg2rtVF6qoRmJB6mER5HC
q7f/7WkzNA0dWxwjAEkk9tLkVhrlF4vHCzJ/rEFT1pVARKH5n/cI3QwRoZ6F2xmu
goklzn04mvXJFa5nvENfDrlrOT49EOWJJUah1y75Nuqy+aj5n51o8Yax1ibctNOj
65voKjOZ7HOGTbpATHpJFUnwAYbKiU4Ix8AFPDw14kXgSbpvegBkZddXvQdvGbdK
Ssh9KWeE81Bc4dECE7hR9ZILFwIGip6VvFad8Dt3TeqzqD4vfsQGN6E6X1dzX6Zf
6Yo3HyiXrKt39TFRMEW9wO47g5KAD9IdBw1DRj2H4BjZBYIhe0Gjs0bHdkJVJmJx
oCMce4TZilsEGtokTcn4rtvp35MJStDX6Ruxrat4ZMEePVv702xKCmmRtVxc2Glb
w3V5FA09DUmoOhPUCDBvWG5aB5c/cEHBwDwgK24caDkhWP/j/RBwUbasFmDBSyuj
TgPxXPocvKulIVqJ8CHozYg4lH6F8nu8YdiSAGNDvnzSzxZAzdFVs1kJINs1bSPT
bEXXuCFwEWAuEESGlbHfQyn4YkOTAWOwIWn16JCwWZ7PQf80KdP6OH73AV7whaov
iFS6bK8HxjHoNydLF6tfuwtv2OHJvXnz+mTm0d9y/0pWXBHhlgPEfKTXC/Z0/OYY
oNzQM7OjRbeYxCfDpLh5cL2S4B3ZCbc+fxuy4r0BpeFlIv6nKMnRGtSMOG14cSXc
vrQZCUxWEDAjTWPqiAAlqPKsEBVHA4lai1dTBH7CbwyQLOaEWvaAj+k7EPZAbY7p
QwHn7SKYanWUcmFRzu4onUcsC4QjGWSe8DCPs5RNBEbVRtDaK3co0RrYrBveKYrx
AofkIE+Z/II1VuxMCbfmBFyyevvTSFbKYP0WmddWhVCdGRNnRv5Lcwndj35a/n7d
ndZDXJWrARFD+D0ClH6NnTwuq/IdliPe6tLyP0czXb9ALNEeKsxSzD1uQYChBb4e
m/RCeQAntaLCWAgcwAvzALkCMjkqg0RdJcV3fNT164r/PO9GNEq92h+9GhKssto8
2iVcsa1exPteededSj1/4wkwZ3/NxmNgzfyyTMKzlOLFDsY/SbrsCpPJppT7TXpc
4H4J2jFLecCchsOFzt2TMJOqN89tesu5AlNpjWrGLzqEcthDsc1IrN/THryWKOGg
D2QLydT0mLOjkg+ksTqeYCxDoi7XdjGIA8kBpdIhL6PblF0Q4vUYvKiUwXwfOuWL
hyZmvI54Rh0PevhwjEdI5LddooYeRvHsOShvxoCOnRXQ+J4lboOC+ggnhjSthizX
8XYzGzCLFWA3kg1dyHsI0KXcA+gmBKPTUtC4eYr33YPsV5ovvbBSfvyTzY32KxBM
WOulW/wpqavADTKvX96ue6l5jKVzZKOQNAprK1u44qpWCY8OJHCJa43lLitYBGhk
qkizNT2dJh1EPPaSmG7ueWdGZNMWpX9h8W7b1KZNsX0yk0olAJyG8jqtnDqtTo8r
10Mr8eFCs5YfWzZ2M6whNpHI1ZYmzUutF/LOaB9rHdPbDOg1E8dinuM4wl/1381k
Cz7408TF5BQNdDPLAkTu9ifN+EM+jsOAWM9aBAxAjOq4JbE97aNiceSnoC4pSruc
TaFrMDyFZV9x0JiCs1gz0b5sDpinbwbuCDHnJdCEC6lhovMIuT8dZ6WQnKRTp7od
CwqWcLL6Q81ahhEyDfMfnI2fry/HhYf+Z8WhNjEnKJQKDadkacm5NFOhtZmDczuD
hT39N3uDN1T7fafVPcZraIWNPp7mduMP8GFxynbMtiBULLZjlYzwU9hkq7nShEOd
mlPavJt10T3/eAjxvno1GckhAZfZz+mhXY6phSHHNmEiGOwMLiSbY/WhmcsGtoRh
pJh++8kaHXmGCjTO2kaUe5LdLtzgMjOF2vsXlBSfV8uI/aGqA6ZqLxcGi0+biXpj
0jr7Isi4Vq8akgDduFyrK1dy/hjEzmJAtE7qg4fhOPWXe9OktzFZfp29oXbV0FWs
Bbkk9qjA9XdMF0VWBGvpq8NjFYFkhpWFM7uFKQiqrbwekJOXRWF+egTJvIKy5gsx
7DzvOxA5e7ZCOcBv1HWkVkiTCtf77/Nsw0X9GZLk9Ul9pvez8obNe8nqmCWBvyST
sl0p5R8CSfKm2CqUv0y2LD+HoR/1II85WDfJY/hUx00AGoVCHjOFshVRD0v3SjDT
6xGBJTR/AXyoMU9Wi5jt9hC+fUlRo4Ux2/wzz78CvT6OjPDj6UYd6oVbazvORSNg
f+h5Leo4m18QiQb1Gee7ysF7n2qEUEGam6644PKkl0IvTenwrBwGWdiNwuMBBMRb
Vv48wDat8/F0h6VKpw8nxS3aP5/3o/nGBZQeoLq0EzrM7I6rcXBORec7xXAnUnWc
kzeb3kcc3qjNCQ/ceBmSk1UuaovSqVgtrM61q6wBuPNp/vOCte1iiHADhzhwk2tS
IfpI2F1f0MH72nvBzEiOKiwLJfPdRk3WhSvB5lJVRPfzrHhnlfy/aBPCgSVkTFYR
EAWNloYYazHQykKGq/avRvTCQqf7kclXN/yvQs4iFAyBxdIie9ZJ75ceVMOfbH+2
pJtKHMxEE/ONu71Ujfet4Ji+jH7/d0vu8Ft+kwitmSQgdBYr9D/wtSnbsbXIQcVY
SaC/uZ9H6IWAKXpyz+lHzsbgr3Pt2XG7YXeAZY8mmZMGwCZy7vydCnpCQBZ563Kk
bKQx/m/2LHi6/9EKQOyTo5YNpkx7vgzDr2VueZj9bdXMiFQdykLnp2FHa8sZ7sLI
qXDXeq++uqR0DNd56D6XK9NNXEP8ZbvvOU5+x0Xe9GIIc6614cZu1DF01hhObu/9
neVcWp054hPi819FQ5WAvYFtzKfdLavgAz4TUXSR6EeTVBwQhVF5sAG1GYDk/Ror
8oA9eweiuWUKjw1yZ/bXBkhgUG8M5up1MNgqrsBC5aowqmwLTm2v1CmO0rqTg3mD
Gg1Uk1K0T7lQdYFj832tj+FhmIcQngnB+UGzBVVP0Eazm9HAyFDKGiK0WirZYqFE
iOXwQBlP8Se1U0DhfPT2IZlvLtOG16twldBdLkgtyiPZfkm2Z2tsMFjqgtS93ipV
b+xcDBNKO3yPglWq/tjEubFKIxk4Gx39pE36MfhTHUMQMM01gyN9Z68UQ5nYICL+
m2DBItrvR3rjZSbOKffyzOnn+l7+xpjBh+BBE7p2ph52MeKm2ZdjTBH78oV3sWAM
JdEkKjFgzDM8G3Ad078JFPZV2vxStWooHh4HpCBijfsipCzjgAgRm5CYr2y6BKLO
0ZoLrKhvoDKvp83tSfE9R1QgUo4Z5DgDLvLUwUAthMygetfnfehbYumxrgjOdeO5
V/zG5+lJ7OLzPpgzlyFSVloT4Zaw+5g+NoPiCZtABxjIpXXXFm+qG+3ZcjwTNZGz
zvufIaQjjEPG+VvJ2TLHl4CJELPMqXzI8GEGQlkzM+6bYhgcjsj+rDng0ymXzMIG
viSWGhIfYChwceLqZX0HMTVxVwHIER1wZw1CyjIThmaGFZEXPuTNeoDYseJVljMm
+8kjmrmz2FZxQ9USRW7edT+WwSU1O3U1x2cPqAhnK0I3byqEPZCLSLnBZNxjB9fW
S2XFcuJGrTmF4vZ8uzRx6y5EWiA8OUrOpIwHyq3lXPCAXCkKgB79iyuo9L7n30Lf
TlKU0JC3B+BgV9XUwnR1POKSOSZrQhht2bjJkpLo8HkhxCAXlgRdsGOYdeaOscR9
fjMBsyPcm/aJveVpAJj2hb7WupDXThwRa7a/Vmzvuh99eUi7Ty38slfMgM2SEvuV
YODQISVZdqPHlKfmWhhb0PWDCV/guB3xgFz+jOcHI9Ks7CJaUsc2+vlLWFzlATzK
IAOIgn/ffDstSwxn1ApCAnsJYyAok7w0AgfVAhu+VuYxCoQifW0YF6eN0z1b/N1Q
PF8pLAmmoaTLYijqFUenFHVf7o3oeSbOHBMDkf7fx0OBWQ+g6KmTub9xh1hsDD6i
j7BPzSU9uB28HLzTFDVBf1egLmglhOzIIgtzw1uSP9xGlg4WIsY3cEGt6E9X6voy
nUQofiOVtp2rXZwQgEOtW99IPdiNg5BMq5kCYd5+Csp0959pfaLloW37aifhSxbJ
h9whH2/pFHIsHUYvlZp+WZWyrcNrdiLX4w2s9rgQOj0VIjQpTvuFgype9kcXXChh
0bOLy7KsqCJYxIo2FiSc7qtoGIzgE2pIGjjYjSX6qKHy11nixJqaKsDBYn0V+uCo
xSZFUAGgQYyoAN77BRrc1XaLWeN/dORfrBV1yV3u9b9GDDs9gLqKTLYmNVndGHuZ
Sy9u8BaGYv6z9lKoredILl22BWwn1o64ulcSZ6IYdDaQSIZqxysZHE2TEU8NBJjL
2NOjuaOpsBBQvoo8q1MHcdkxwIS0Bl3ogOXkqGkWIPm/yJprHu/F+BCy1Ih66gSE
NRZdrTidKwtjYhV6it0lwUR1VM2Knggirc5rz2vm/3EdJdwNxNQDbKfsAP2kpvcZ
OlQjNR+sjMTxZB047sYhAxy8ix69n7r/gPb7ZhjrDqIRoIiBEt75Z4f8QMjdVSzF
EZW+EnwRf1su3qqaAgYiitGt85Wg1l69LdDniSrR6/mBty96KsxMLpmNR8VO8+Eh
Fe4CLADsnGXLv3ebTXNG8FiVpNhwrFWRj794VqbZX1tmUhuzk6LBDXaZP7+V679f
XYL07d3PlQHEVeNeofB7LZUtEI2ZhEfz5rmg6NniYradSUtNtipjieNf0zF5eG/v
pKh0Up0r0NZ9yMotC8wJ7TlpK5GepYbT5WVNELKLdWpalami8w4rj+SyoYwhwBbA
zYrYhJO9vBQ20qztMoqgreTICWHBRTksgWhaZJ5It55TDdFOY4sEUFZSOB79Tgkg
BP3VrxTRzwHDx4VCclHaVfy/taJWhzRPaxIUBMrjXcwLvaSLMVK+hv9S2/w8UdYf
ehUb0dVpsJVjnBgp1Qs64KUDG+zruiXLQPwjjMKTANoReSv+2W81sHHlN/WWPnPd
bEOoQs9Z5dAmkSbJVdPkP0YSyX0iOQcflWNHglSPy+L3lKGflc398lCOFTdjLTNS
kattxGmH6jhMHKaVN24z8s2300wu5viorRMXzn909goMGRihB+v1qDC8KIJP0xGD
DzuiRvTl5bA7BjA8YEzMAF+VJZ48re2xyh3lDAnRBHLqeL6i82hxytnJn+LEWsrJ
R4nG/cZ0wPkxrgzW/9kkgRw3JPd5nv/wbk1YmMGDp43NMP7MitTs2cxvBLGawbVX
3LXcFu5aj8VnXuv/fZ8fCudglqHIaltxHG5SBoled1Qu8agNDkcLQwTe1SM8uXr0
48F4JVhkcnE7NAEo9Xro+H8P9vTIaBd6MdUir75rHihQV4eYbaDEGX0vuDf/v3QE
C7oEvIMzcliIF40aeg4G/H9vi3wlC72QM7iwUgxji1HjOD2nAAmnCfkGgl3eUeOe
MZ4P85lq2Lzo27sjRaWx7+kI7lsTJ+erv7Icwamm5pbHwd0e90DQnoZRjf50ubwI
q2BQEtRqqou31JAS8v4jPP1Cw+KY2A8QyGxLaB3onLIklmReGT7/YcnohOjV1oU0
ZDorLDJEqyqTUIRwyWsohyen2onOM3gyJrbrF2Qr6FsnChWETD+H+WRQ0Upms0AP
8id+opP/LBvhUhf3z4BU3UaNe7rzd1dylYOiZAQpOsFpRFGtbtTs4x+xkYIPfTmS
wRRhKeNGUP3kqxIl20AFJRxfR04qPLqIep0pM23zTZVwlXM71Do9f1mB59bwxobO
e17Ozp9oUzMVwxysaTKNSjMyaEDv4QpbhNkOE0ERvZQqsz6heBaqnToYX1X9jeVd
/weotDWvkxAkKu9rJhRxwx/H4uJHu6U5gjw9UYaI0NqfaLP454tTH/+fKTwn6pmI
0botbgE9hOUUTWdVs17KhUVhyxg9p4cx/1167yE+AyfyyKYv8VS05s8jfq+VPyaj
jk4v0sBSxAtb2YuN030lDvq4jbc++KEAtqXwWMmSxGisPrkv76l862Uv7ovZBWlE
1Mng4vMP/2VJeG5GZugtYBqH4gIj6cNM1FR855NQW/VXWW/eMi+D2Lz93zSJOUGJ
J+L5ZJ+TF73EyG93qNdt3FnFLGIM5gc5qRzQHHASPMNYLHjt5dT9ijEHDykGi9Si
7i8Y0GDvQ+IZTQpWgmbuCVwayV7tTkaw5xy907EoeYYT9Q0ZjWmMtwvX1lX80KPP
uG7j47qVRlWXsjuSYwSTWRMBFjoJvnamA2y3O8cl6GGgtxaNECEhkvpzJ0PvSG09
6mzq95b7Jhr35LhDRwPBFxLSToYXQ2rjjRN6WwJdw9c0UYTx/AP7ZeShddVJ40xV
Oi07/tmS/RNhsOc1jNqF+itIRGkeefoqPc2XS95eILnbp71CYTYdqYIJwBnjj2/E
QVIX3FJYTty6jAKUGT1z2Qy6rR9M7GeUYDO8XTvTqDNJztaJYv+fZK9Ra3G+0xUD
i6Wke5luC15aL1yk4TSgdCf3PnmtpRWPk8T8uvkBOIca/QOiYQ9R0NlTyYjaFzaQ
0Lyu/eM8a3Hvmhz7ZzTrgashuAXMcvfsfk8La1EZMhaqsKPTyc9Ymm/kYsF7q10K
/5zq4Jgl9ahEaznCrLLfpLLWQ3vouF7Ir4o0AJ2LSGRLyR9z7dZX8tJhhbbxU/tf
Xp4X6eSzYyJSQ84CQyrfyj/stvyq8WeUKIznEor44iLGqgjEP1zhKpE7yI8SLBXj
oHI8b/UXPZPyxhvr2LfPfYnR1F8YEiScVi1Zy63GJem68hYo57ziSajnHZJWeDd2
IKrGvwFq6Z4wXIsgTdlps5ivUF62nqskEFp8x8eGFEtdI1WSTnWaOPOKDfQ94M/x
FtQYRGAkmPJoTf11z0HWQwiKEnaQHK7UMmRsP16CZofrD+sX2ziFMfPBWplu01jT
7+m0O1l0hPlxOzPgD/vwY6nt6BEWB17isFlXdMzqLuIWE4VYLxpt7dDArzMtSH9E
aOS5fHjP6DRc/LC6S/q8MUJFIqZsLT8uSbRWxQgMyJ7oxrNgHIJtVUD/UYA9zSt9
m1Mt5tiaSYputhaV18MYSsVArvpHiPyq8xZVi8mCXDOLiUkAaPjZHDgt2gfXF2aQ
3xFhBICzBDXVlktabq9Gq10V4lEisMbpruxiOMJ6IeZI2aJeHIyoErNarDOA6QWi
0MF7BqEPnjkJ6vCj2eajFcy13IjY3YwkaibkoGL7tzuUUk46OKX/zp3aUx7g7gMa
MRigjxgQHnh40gur6rN6t/LWLCxQQam1U+27XPg13LJ8fUYG7enTmn91Hg8nfO5e
kGi1dMzO3+rMR1rw6fKf7PNTwL+WS0aOe/ZC+v5pvB0ZY+YvviF9kpJyHdOIINn4
JIhqcRf7DshWfLfc40sHxy0HRynzBYx1BcLA4SJdT9R9t9eb1WOlyK6pcBaXyN3Y
WBsGVFfPtVwUn3bVisYEGTm4NSI36+5Wt1txZJkmxNy/pHPqYVEKN1UmUQyqWbAX
oePH9KhDTTfz/rRyKQJtPj7AaI5GWxEnTxqp4RQx7//5OvNWnS9XUp2Uf+W7DZQF
huTxx04Aq3rpYVG/c3/C4SO1NboJrDjE72eFEORot9DlsLPGRkpseCbt8t+lNZTJ
P8ZE0pXx2uTHAGYscyEUPkpcxq+Eag/6mm8bPWfc6fqMnbsc7hYwn+F4zrm4JuLn
x/QbTV71dgxX6FyWp44zS368m+OXohqZlrAZoXIt4JCRF6BAP1zj1N4a614oNMej
/LInuRU6Mt5xl3YkkeFKOiafp2SvZ+V8xuXR6Qb8YTbxZjgb28/bj2MRDG8lzcyL
BVaACg9qqV3l/jx+mIb2tqqgkavsfOaJuXekHxBKmMTgPwFFVlyaPSqu4+HzzGsE
fmRpjs53CW/6PjnkJE+9aCZGcHIsmMpUpSiXW0vm4AUsz2drEM9hLS1O7/+oNyOQ
rTyVbjPu1wO6uUSLKVnV8axjMbS/FUFTZ6Ozpw7LeokGvWNDSI/jPIkL38xjYeoJ
HVdCENkqlwJsvPgkBktY7x16t+ygNg6vzex3SXzwdPZNsc80bfNllKxuAGyOFZWs
1j4Ba1zfj7UCMvpRauRsztDfAy88CN08B2epnyUN0HXnfKhyi4+w54rULD35z03x
k8m5SQbF+jK4LGPz/ESqFiCGVwuUd7JQHjiUVxb9heZqmFLfViYY4qeOVCvpGA++
LuxyXmSAjNffVEVXHt7TTr2cVu8rhXYA+TYsWxaYp0QzeEQmK2ZkYxHyCVPpLP3v
eNqIQSE+hKxqgV2Ssjofy6QX4mqnl0E3SNNuppNluWjICuKHKUBz1FHjzGabFR6Z
AenEVKU5j5b6JCmc+iwW+MElqGI3DPYaav6nCHbiAYRH+Fx1E65UpbPFESsyeqTA
yVtGqjnIpfRwpnsEp/kNwmwdgUsx+8eFwyKDMYsGcdmBlA0DH1SMZyMhj/nqjnZF
xCtp4HcAaWaDXFy7e/qekpJe2CMo3eCvdcmbb/dNQMUsg0h36xQGZxoLLQpeJFI2
hph5xqt8QtNWfczJ1dUnMnK1cPte5YS8r65s9xt7lyEVKtuBnKteEaeFAYhRJvry
UZnLPra/uaZTPgNSJV+yFKlIYsSqS4ktKVLSu/D8pC1z/bTyWIUqnEvQiXT+kreN
nY4gTZATRvcrsu7Bd1WVO8+KOg+bC2f4ZNno7Y+Ona1HW6bcuJKsphBtMceDWKir
zpv6wwKyk7mpBy9tRSvEvtUjATMAdbaJoDDUYA4PokNhmi+9mDsl3jbdnNw/O62X
uMH/RWXOey0QBE3PgeuNWLEcsHtzf+LLtMQvLwmx9dW6MEQPyKI8/isWjp4A44V5
Ona1opmhVgHOjmh4zR+Lzj3cKpT5laUkMBMmN9/bJXNyo0i1WB/geIbKnOjiMiPb
aX9Jux6P4r+1gCdwVOpFVrUQKjOEtUh/vhuPV/AOWx2+cxV3JEu2CsGsIvBw8grQ
UGqmPTVDGDf/ySOGCghmg2hBvTQy5xNDAJvD8v4NWWHDJm+W59ZPfUR3oTxuupLM
FzYl3Nd27lkMKpY6J/QOGN2RQzbS+KxIKTh+bIev4VqUw8PXoE/OkYXqmXZGiv7h
mZERc/ZYXh8NtQsVnT/3Ktx3J5ATEhp2II62Qerg31SfzScgeFIsd/RFpk19kmTy
5ndjN0ya7gJr/wM26Y1nWIHHff6/lxawfZSX3xSib3FdsF6DgoxUW6BdTVaT4TmC
3J82Q/FwU4GosN3DLrYUBH41iZSOh42Ob1urhKybaGzwisZWsYtPtd98h6LIKrqS
81M5gsp24ytmzqUsxbbBmIg/jSXs1JluV1JRD6QKCzJr3gz+6/dPvcoYiXHiLpzk
v8bkq1d6jJet+clGb7FudyxLUWzCetvc4PmzX5Mgez3OCLX4xWl6ffAlcSAaqdE2
Kyo92FBwtFdgAPcfupvTM7w4JMOIuRatPHv170aGB14avU9CjwH38WG+SGHmfJga
Ifhu9RRJ4284K530C2LBSzALRvKeIr1fYAKDvMK0u+PhK3cjzWgj4Dw7QJouYtCI
IWvqQ3cNFbUFuUEP1b7zfmaWLJ9LwAI1o0OHOwc/OGRv3bqMNzJSTfqL8sMdtA5c
1wJGOojCD+JPCuD9OVipWHBzNqVBP48wZFyHxXaePoqcMuvm+7cRW3VIVE5hL0Pw
rE/Wpxct0GkvPNPfTRmO8LEvDmMqWWeqjiwYmuBYc4XtUsc73vGIfdoLK61FFBlJ
iLzmK7NA/SitW33y0GdXg6gWGx+zIwgW0pZEZPluzW4Z3z2trI8lVuUB0wroD/YG
tNluDi+J6/icQwWRNUD4KClQuWdEd/DQBwcgvzKKyPdQTAaLFeDuaeSr3O87qP8R
Tw5hM++rka3s4AO1WuXg2CrFn9rBdDtqJrjNYf+su9pF1ko2vOX+QA0kjqK7E+j7
qLbTttbQbVrdHctzMbLBC0mV/jb3fTL2Rmu+a1OcyQrhCOKboA4TBOmdPt3gjpj4
rFnFamaclVSAuzYuhIASLnL0coraPRX3qmKBvXmeFszfqw9J8cXpz1OSZDtU+BKI
vV4a0vDCfALVxZ6/ylC5d+Pc7G9so8XRSaih0/KornhGpKgNBGISN2YZofW1cL92
MuaUWerUJtssjp3xoNTOht0C3MP81g5FSTpRrvPFwYSUQ6OtmmyE+7lCJGrChXSi
6qI2EiykOTiM3r8HRPm7jchRS01xLS0YFPOviErgz2HV/nk1tQ6xC0B57SnU+PO8
EA2T/SgbA845nXNlwVSWhQFzVIrtTLtczN6Fq8UanPu1y53BZELeNRMlJADhr288
ek9ErClQSc8fwn/wP/QU3LIk3miLgwAnKkKOvWIz6SdKd46bOsUfGYTrhcWPF4Rf
z0luq6yFbllBjamhxADU7oopzQymucBk1o3DHszuCiFmRcLGGtJptyRVFE29zCOM
rzAd8MBnOiDrmSEB9jC4dae0nLbwftBw88ojY9ozx6ydH50HSJsQEWj4VDliswZM
hABmwnLIQdqVTNi2WDpi0l71ik7cYaqVvnUu5q/X5V9nF5FsQ3BqBZbk0D4BMPPV
+ei8GNg3RnFRVRAyQLFObz0YdISLknqpIi6aOXzGQuzqWtbloeN+cOOo0eih16nU
hy/S/b/ZPt3DyDusTh95L5NYCFuwaQSoJXr9sENKnpm0dX1hybLrjhgKSgnXUzmO
Ua8r6pRgmMNyq2NkJCiAqJLiT8zDuA7LmA2tOw9zMI21Xu47F6zWHXPDZFayTIhR
PA+D6PqUa4r6cOhoW8ly5/D4B0sXFAgFrUfE7QEfsNTYq2m0gAFCg0xDjmc0mjan
oBxM5FFE75YQ8BlXCrlJ+eEqhmd9ttxMowkiqhQvHJwXbUZ07b3iNY9UqGh2spQG
DbUSnnL9B+ir058ICLiAEj9dYFWVAq/EKHCD34Gb0BIL6DzOiNXRiPzJYJdD3YwY
76bUkz+NCh7R/hb27TNLF4VDMzKcHlAze4RTu2JKbGNw+L/L1RtjmP6pMk4iu3BL
PxNP/qmZNftv6heZxgkFW3ORMZKElspgzJmBwnW/uEy3h9/KcLF/l3LwXP3B9PJ6
qB/FY1JPIUNyNefTpHC6U2ViqU97caRFNRKywSaz6EK1fzj0GCs99TOlV3l9hWwJ
3OpQmTqsgujK75W22L8PMWSQflMLFGHlXht+nsdYCHhQUkHz3PFXg1P6MwEZ/cvP
xJBK+rDdIvnOYnPxNWYeEAJk5h8W7XvhXUKqJfaPcGOD5JVW28WpaP/9RiIY+UrJ
sUoy4Zc1CJtnDwt9teMd486ow3z8qLY5KeWsm6ajUUkCvWl/FCaKAkI/dj+nE0bx
1HsilRXiP9Kp7vfQw9tmaWvi5NKbp+3qXDLNZ3aUk8f8wGbLrw77HxwWrOgij5q5
nydMw4bGQc6GenycKfku3Iuo3bJsLo0U7pTSs8nVQUvvgbkOPtKO7AjtcJQpxm8m
Ytl7HduTaYCX2QUL01fS1UgRVIcPeBaH6YtdvfOjfEwSFKZat1VNe0SeixrLO8qG
EpoZnpDA1Pm0hTzXwZdm8kwXb/LF3DXLD3MHdi1IImsEVY2Y96MAk+5K6H6+MLKS
IA7YP9qP3EbOjMBu9nvNWVLECGIvM5WTtKIUMecXks2X0JeRKgQgOksNr2/YmSQS
OTXyCh33YRd5UsAG//pdATj1zH5EZ1jrwMpeIOVxhYdcZ+O+wPw5ko2eTtmqDrNd
Clr6ArXA3TL3X2cu4Aw3saqTO9tVaxPDkN7FeGAvqv1/+C49Da+Mgi2nbn/+03TJ
24H+z0HeKuh74LSM7EmsP6Zgx2f05kgPBVTCIZ1eQ3rk3Oq97H2OwlnU4o8bVrb8
kwWC05y0+7Iq76VcqnrFUIzSyYEbfoPVGuJNM+RuAU/ZUwqEXiakLpPyjSzo1NEV
GvwMqD0RW4o/1WUIzSeh7zDCAmrx+II1X9Xn+FjNYmWBLUFtzaQW8MxA6ElAXFUe
I6bzjHKVF7932pFW6OFZNyGdktPujdvMCChDT0OTkOT1Ixc31VATzcT1Ir1hfjXy
UQcvjseTUeQLUR6vg1mA6XNrV88RdhWzDv5zyGgmTVoIvTkZknufl79FJWqHelT3
3+fmNaWORz/Xq3mlAteoI2W8Fri5cfqnFwUUAwBFa/O91yXeQSp8or+oRb7/kPUq
lOw67mpRR3WEM1FFlafg5fEFvHZXMC+dOQO6Ea87Zj0PijgA8F5uwhzxpLlmBjHY
yPHTKqhm14OReReeZWC+W4jg1YmDQwbZh1ZL2NRTqXRhu1qGLuH0or73RHwaOBGy
PX3lahzbTonmI/qn4Yj6UEiEdz2atrPGTEwLj0zrgAeuJgcMBtlSGR7MwyHw/0Ty
UBD+mCFQkrQYskJenu/p5vw9dl13rwnk6Zc3DBsJQ6jaTWPlLO7Qalz5+s1W9Lai
ScMNu3ha7YlP+AP4A7ABt0wjV7oBUqGLbgtaWthnactpc5dn5n2Ln0b9UIpnKLkP
oYzixhQ7y0TP4Hld+65XDlqEfXkjmXz0Ie9AxnvXmwDt0QphOjE0hV3tnonescq9
vLlYrxEcPAuSvOpobaYH6HaNfgqyQX7h4Bz0dVuV6mV6AaLxGlh6J1xsq7OTtxss
+WkkDzqInztTybe5aNcVq+TvXd7brBtPMUyCQb8M+6MbQELl5slqL8Ggn1r5IHyR
ibMBxFVV557hg9ZEOdksjEuBTLfQYVHKGn2KqQyPvPRdnJh/6ImQoK2PB9Adc1lb
Ucbvlu9o+eIVU7FtB8ACpnprtCCjkY9QqlWoroVETv1eh6zKwFYO7ZmOfcpI9Vp1
iGWQyA23gdiAf6VUbch0VJvJvJfJsQDXi7xhOtgCiqdlUkbNwsbdqbzHDq/WGdGD
hMG8dtTsAWH/du3n3hKZlJD10jkGG3WdBcl/uLCKXFHpD+vleJRu/RWpgCrUa1rU
+Bd7AxCUUDSSWSSgh3auoubaSoI6tTFGpO2WtMXb0ixC8ZSPj806aHencibMZYxC
hGu0BaDS7JHZB7bOAKfsGsY9/H0E1dYcceo+/9TnNkGpjWkOT2YadVb6DbHW4PEw
GAIBMVZpq4IMp4s4WbWH8EPvvvfd4yjr41/RB/Olykbst2LrowWflKJaJoEDouh4
ynDkOoIFKWVo0QDx/+T5Db5dW/fteCVcCK8ZLKzfqpeblv7mZEyAoE7sq58mJcC1
BnJzk8Yhy7dJOebffZZdU7gW+DZ7ckhm2mbqnHExbWSgl/w/YyRFLKzM1tvGZAnQ
8+dk4DwK5JPuhA/pr6PfrOF0PEUyrBwj/xovkT76TPSP/ZONxfeOmfGiCvRXFfWM
rY/qzn9504SJwXQBo4kpFEVDL31FefgbrL3IFRQl/ZEH/1VZ1CVbHqf5g44J5Txd
Mqk9ivxA+qbdUPmUQNDsFWJRsRIaAP6HprWStyNHmYaETWEYaRfm6/SehqcG7Usr
84gq1fiYnt4WykirYD8OrdwmmLgVx915LrZiHu454/kX0NIUu8oXRlTh6duKMVOk
3jI2JBhUIhmBAfRooWLYbhBM6McwLom3Kx7JpVlkH+6mwvrsXtNWth6QxBC+2M3b
7nWz/P0PbAtpnzvPdDwr4Kq2O9ht+BzPeyv4Q4ygdurwIuftD7TOBa2oBjz5UKeO
7roTjweb+fmlzxd1tari+h+83dF1+Sr5yZxGiONv+0TXIuPW4efwpSC39Yp6cDnx
/IteCxh1YENCh3PdbppCtg==
`pragma protect end_protected
