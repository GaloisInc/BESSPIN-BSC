// Copyright (c) 2011--2012 Bluespec, Inc.  All rights reserved.
// $Revision$
// $Date$

package BlueNoC;

import MsgFormat        :: *;
import NoCUtils         :: *;
import PCIEtoBNoCBridge :: *;
import TCPtoBNoCBridge  :: *;
import TreeNoC          :: *;
import MeshNoC          :: *;
import BypassReg        :: *;
//import BlueNoCXactors   :: *;
//import BlueNoCVirtex7   :: *;

export MsgFormat        :: *;
export NoCUtils         :: *;
export PCIEtoBNoCBridge :: *;
export TCPtoBNoCBridge  :: *;
export TreeNoC          :: *;
export MeshNoC          :: *;
//export BlueNoCXactors   :: *;
//export BlueNoCVirtex7   :: *;

endpackage
