////////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2008 - 2009  Bluespec, Inc.   ALL RIGHTS RESERVED.
// $Revision$
// $Date$
////////////////////////////////////////////////////////////////////////////////
//  Filename      : Xilinx.bsv
//  Description   : Xilinx specific libraries
////////////////////////////////////////////////////////////////////////////////
package Xilinx;

// Notes :

////////////////////////////////////////////////////////////////////////////////
/// Imports
////////////////////////////////////////////////////////////////////////////////
import XilinxCells       ::*;
import XilinxPCIE        ::*;
import XilinxVirtex5PCIE ::*;
import XilinxVirtex6PCIE ::*;
import XilinxKintex7PCIE ::*;
import XilinxVirtex7PCIE ::*;
import XilinxVirtexUltraScalePCIE ::*;
import XilinxDDR2        ::*;
import XilinxML50x       ::*;
import XilinxML605       ::*;
import XilinxDN10GHXTLL  ::*;
import XilinxDN10GK7LL   ::*;
import XilinxDH2000TQ    ::*;
import XilinxB2000T      ::*;
import XilinxPDV72KR2    ::*;
import XilinxDNV7F2A     ::*;
import XilinxRPP2        ::*;
import XilinxRPP2SPLIT   ::*;
import XilinxDNVUF4A     ::*;
import XilinxKLVUF4A     ::*;
import XilinxKC705       ::*;
import XilinxKCU105      ::*;
import XilinxVC707       ::*;
import XilinxVC709       ::*;
import XilinxVCU108      ::*;
import XilinxDDR3        ::*;
import XilinxUtils       ::*;
import Xilinx10GE        ::*;
//port XilinxTEMAC       ::*;

////////////////////////////////////////////////////////////////////////////////
/// Exports
////////////////////////////////////////////////////////////////////////////////
export XilinxCells       ::*;
export XilinxPCIE        ::*;
export XilinxVirtex5PCIE ::*;
export XilinxVirtex6PCIE ::*;
export XilinxKintex7PCIE ::*;
export XilinxVirtex7PCIE ::*;
export XilinxVirtexUltraScalePCIE ::*;
export XilinxDDR2        ::*;
export XilinxML50x       ::*;
export XilinxML605       ::*;
export XilinxDN10GHXTLL  ::*;
export XilinxDN10GK7LL   ::*;
export XilinxDH2000TQ    ::*;
export XilinxB2000T      ::*;
export XilinxPDV72KR2    ::*;
export XilinxDNV7F2A     ::*;
export XilinxRPP2        ::*;
export XilinxRPP2SPLIT   ::*;
export XilinxDNVUF4A     ::*;
export XilinxKLVUF4A     ::*;
export XilinxKC705       ::*;
export XilinxKCU105      ::*;
export XilinxVC707       ::*;
export XilinxVC709       ::*;
export XilinxVCU108      ::*;
export XilinxDDR3        ::*;
export XilinxUtils       ::*;
export Xilinx10GE        ::*;
//port XilinxTEMAC       ::*;

endpackage: Xilinx
