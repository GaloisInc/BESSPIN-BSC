// Copyright (c) 2007--2009 Bluespec, Inc.  All rights reserved.
// $Revision$
// $Date$

package AHB;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

import AHBArbiter::*;
import AHBBus::*;
import AHBDefines::*;
import AHBMaster::*;
import AHBPC::*;
import AHBSlave::*;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

export AHBArbiter::*;
export AHBBus::*;
export AHBDefines::*;
export AHBMaster::*;
export AHBPC::*;
export AHBSlave::*;

endpackage
