// Copyright (c) 2007--2009 Bluespec, Inc.  All rights reserved.
// $Revision$
// $Date$

package Misc;

import Arbiter::*;
import BRAM::*;
import BRAMFIFO::*;
import BuildVector::*;
import BUtils::*;
import ClkCtrlServer::*;
import Cntrs::*;
import DefaultValue ::*;
import Gray::*;
import GrayCounter::*;
import HList::*;
import Randomizable::*;
import SpecialFIFOs::*;
import AlignedFIFOs::*;
import TieOff ::*;
import DummyDriver ::*;
import Gearbox ::*;
import UnitAppendList::*;
import EdgeDetect::*;
import I2C::*;
import CRC::*;
import CommitIfc::*;
import NullCrossingFIFOF::*;
import Randomizable::*;
import PCIE::*;
import MIMO::*;
import Video::*;
import Memory::*;
import Arbitrate::*;
import Printf::*;
import RS232::*;
import DDR3::*;
import DDR4::*;
import PAClib::*;

endpackage
