`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
q00T1GB6QT3WNBO9hJPk0S2yfCBcgluQ4DDZLXmSo83C8Qq13De9/+TX/Hgia4aC
l1ZBFBTCDw3TN/QNuOC2693RWvb5jEv4hGnIQsNl8sL9dN3ZOr2Ctk6J9hVIx8Ck
ljUvD0LOh1nC/jrV2mSJyhrqFvFJbbGurN7cV6IWo4c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2992)
YjlhSv4DuCqmjtaBQVvJJ4KqOo79UabmraxB6vwpIi/o7fG3DEWVwDNsq6NbrK48
u5X2buSl9JDamGDvVGt+ekIYjrvrCdEYTag9VQ7KqJlg8aYSRX1cto5HrXo0rpfF
QgvSpm33YlM9jJYrtxTeCMZLgMlki2T6mhGqk4MA3VyK+/hjywIgtY+LPG11p8Gv
71QmUYHnId/qAaYCzECD3kQMK8WNL5Egr0TMVgWDkxBZJ7Ia03Jd1KE9/yfVV4wP
dxR9IbISFiCdt0xVImGSDh3SwcmOsdq5VCBBbWE4m2TBW4BiFRJGW+o1HXulDlul
tamJ2cdV47L24Q4v2sCqMJFxCxEJUL0oVmUx1eJ5q46I3uolkcfdwGdgq3V72wrr
tUWu7Y9rlxR97YhCjYemzmm+enW3RauhHpFIDsGv9D6CYWvaf42wxS2vNacLEoay
QbqEWGWbQBEgkXP54+dyNgctRsYZQRDnJl5iHR4pejinmDXl4wmMqZYPUMPMEJEl
cK5ixDTCM52dozczF+BsMGBeqHXuFOpIRjr+uzyH/P5IeEG+Y4X2hlaBPlZF//8H
Lw3qphgbTnCGk5/x+2eDymlVthGgMaF10sPHUJZUmEvFdaOaeqn4L65O9AxbFqdv
wB0urRMLvVHtTxsO8o0v0rVsXtk2F1IEpQef8ic1Qq630sLRyRSYzyfQypCBOQ3F
pQsjMutTHB2tSAgYlJIQ0TJTK9SsPwUCCai8vzACHRAAfylj82LfHVh7nUyFTIJe
3SMTVu+WKfoXdkzqMnptLekcQwty6ZyfBqJHSi7nCgj3/+RksUxkQfUy9mJXmYcO
lhA9Pa81YwgfadlEG+56Q0o9+Ey0P4eFTQBOzMYhZwhPvca25FCRk77RwNrS47vD
rdGzRnMYQaViy0L4eRR0AAbb4IcYc2LDT3CcRu6BPI3WWms9XRElR/b7GIkAyFS2
0xPnkV0zJOop5NYTCipLI5XRPLxbqD5OJeQ+sH94jLKtBqVeNYHN+w7tkhCDFJDi
ZqskFfp5U6/zYq+enCSn85c9vh92uSDU1ze28YuACojzl4Hwh6S4N7P+wtneaMrI
1WBFytmttLamehD6yKLAgD/DI7Q6UxHC79McPKMAUUPVnB3GF/r2oVaN7fAaZk4P
qxzbrpXHv3aPFjltzw2r91BmPGG8Z54r/0twH19/cyO/cN1pdEHxboR+ixyU7Giu
Kiet9aLCari6fFOTp20B021hA4WiQ15NfzSejfqUP9PZSRXVIo6y9uVkDkcbvtYp
mMoB/pMGdVG00sal8dyVvvwyBGKmC6posHYgdK62XpAaHzMo1VuytqMmcaqYYSB1
FblzdpmoE1TfXO1WY58/q9ChKwb3hdNd94jdroDcV6d5SXHe1ThFnHLp1DXHsoit
90AElAC4WWDJlJWDwGMUCeO6lGE5fgc3LsD75L6gHxBdUIOmGStO0ZDoPqtGrIT/
szMgghTVd9SQLP0lHuzcEWI2sIhsPHTn5pSFQ4gKYjOVlqT4/6Ogw9PpZ+lcFAhh
uaU54G1powZ7Qzmx46giSWNpgwlatVfLIvQMiw6aUADDxCiGN/sEz7ptYatCfA9w
4fumv4dzBAedrnd4wQa59mqoGDKllgKfoQf6ROLX4f3aonjYAnoVjWLx9K8qub2X
0HGAxNoixoYF/mZ/BHO2cWEmcowibfjgK/uaxxXwBZSkLKuwLxM83RMeIEtDA6xi
GrzIkbl9S42Qpo2VWgCLrn3cGdpRqb5F8QwRdLrGq1wecWKVYcqAvkYepF1Ee8Sm
JZnt8XNThoAc8BfVkLDBE7nwNw+np5KKvDGn1AGOXL9quOgYYn6PSEuID5WfAlZS
uo+X1ggjih4AU5PwkRvEXZpG4PHFc3qlaWIch6WDW0Fb3oTosyTizAZdolBpfH++
fGNmsbvBXHDFJKoa7u/Ds6aXrX0T5ptQ1b74WaTZkkoHuO2pYFuX485sJg4fBwwy
DjMqHJ4wPw78Zdy7/vHZ9t1BaVyfAbK5FcslyBoTqpfUhBpzFHsZzLmdtSYtP1p4
zUUzbOaWEBvXPMIrJQqwmeSvhyRCwNAA6UOQ0RqNUvc6tZm1MR0ES2VjOXdKXZ8Q
HP/yAXFrAjlHa+sQGJ6WRrdEjdScuMwM6CvaGSjNknIjg5dg4ZUDiO7Fcb9Z2r2A
gqYzCo1yDLp8D1xRLuWjxOaXqOPUh18I2wXfPtvnqUPdsgoTmI3G27ioQOhxlR/d
+1myqHucFH3B4E7zrg9HKMLMCcQx3N9oy7ynDWrN6B87uFb+eFB81/EaFyNUbBQd
6F0EInh8gefeXOKrdxmAkEO4bLzldP1qFvw3dQN3U9KZauY/XwRCnotDf0AcEefT
1CMtMdRYW53G01pT0L5AucVw0lgYkVeLkQWPyoEgzstijRJJxVpkCboGJvDmNYAQ
3vegkUHgdcPp45tPcg2L2tzEX/k3DL/aPeo0FU6rqqJusRhNIZ2D/3cO61ggqQ4B
/NJnbi3ORyfv8J4QcmhE8rEKEcRMuh/Q/amDJy6nc6FctF93RqIKSAXBFphagEWr
fABKiiOgDzIcq/yi+H66u0wZr0h4nAdM7GrVYTMzNjtefn/0FbVPdgJ0G/0Bdx0V
GwUaqrkY9dQMXHBACxeNR4fuxPs6ihMluzThYSuq/qQAzhcETDRC4md+8mBXAC9v
SKkT2qKezcwIdM6G+W9baUqvCGmJQcLniQWr4IH65qdI/HQyP90U+iyG1jghF6/F
SP+ylAw/crEeTwmO/SsIyF7mJtAzCwaYY4auGEpjHWAwm8zF1kcGLrH90xcjEKpW
aJd1z+1hwNo/wNNS2cRFciBTh9Nxrn7x8HayDkPflmi8YgnLvPV8XmEl+/o09EFZ
bHdT48+2lSJdFtboZARJ38YXtFEXpZLHEAGUAUmz/+X8a2o8vmpx0lQaWX66XKky
OZXPUlcWhU4YGjS5TEv1O2mipwAZcRxLb05gm/zp6+DwqXkExvHEeokCsyeg6fMH
6yFSGM+AzthYTOtUmKpMyS1UVhS3DLGVCtJpIi/88igOsk68h4Krq5ySX5bIeSvP
9TR4cvI+bmY7YSZ3US0h/l4LIYXrv0eIJu0i93ZwdFK+7c/9mFot1+zEqJeKdkKT
hfjIjByv35/rfWMyPcJe2eYcHAZWZncSwFp5OlgcqXtMBK3dzvb0rZqAfLL5htsR
WxNIZjcQO+PneS23+4zjpltsJ6XfJwxyGG5ePFk3d0k6bPZhez1i/oLXFITnGm0s
/7vNoQt0iYcVDt+pcu/GvJYXS7JQeEx6U1nJF+iBgGmsdoRT6+pTgrsdGgM00ODr
jnx3ohZwpYTySben+97CtbPy90yRsuJAR8DUhOH6pNN6klgHqmMkLQg0GLV7JrhN
fwu4rLHNr0r2QmYrLFt3pA4kRP61QzdDpiBwYQO4foQvKwuoNZRW3AuYIxXR75uj
jIYbRCELUHwYwRaQHjTQbL6aJHggdNaR4cx2+4zTF7m3IZ28zxf1INFwsEdBz7Jz
mKX11coXUzlcRyeN3MsZ/51H7mjd0nkg6JK4B6jO81o6xPf3XqlXhJWYjteZQ9lK
Lz8cFvYKSMaEOWlUnftIoJI4bWw9hA8KBejkkyJ+pKexgNiS4NouhOCr2QV9w7LY
BTtnpObak/BFag8U8Buxp70dPFmOpFLJzwt+YzDFfmLq/YRLm1d/qhvZwQDRb6PR
ZBgnwkW6oTkVtU52NaK6/lJ7xao7PWYdj6V1vFqU8hkckD8A1xjBjV7F+5ETAMw3
Ip8Z7TDnfJXL2HHJEtwsfVG84Btr7Wlv5rEFL98dlkH6v+SVUOTG9ZriM0qtD6hO
2JS0+OyWr9Qt+flPaXMKcQLfl9HeA/sOWjiNvx4PquURRbjJewVanrL4Kjh+kSSj
HX0ihbETyNWby45u+fTP7tziEKQk+VYdkIzs2ENE1s8FfLD3aN9X2neIzs4cnIlY
ECbGDG1d9kqcmmmMy10a3A==
`pragma protect end_protected
