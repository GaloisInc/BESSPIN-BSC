// Copyright (c) 2017 Bluespec, Inc.  All rights reserved.
// $Revision: 35031 $
// $Date: 2017-03-03 12:27:30 -0500 (Fri, 03 Mar 2017) $

package CXactors;

import CXGetPut :: *;
import CXAxi    :: *;
import CXAxi4   :: *;
import CXAxi4L  :: *;
import CXAhb    :: *;
import CXApb    :: *;

export CXGetPut :: *;
export CXAxi    :: *;
export CXAxi4   :: *;
export CXAxi4L  :: *;
export CXAhb    :: *;
export CXApb    :: *;

endpackage
