////////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2009  Bluespec, Inc.   ALL RIGHTS RESERVED.
// $Revision$
// $Date$
////////////////////////////////////////////////////////////////////////////////
//  Filename      : APB.bsv
//  Description   : APB4 Bus Defintion
////////////////////////////////////////////////////////////////////////////////
package Apb;

// Notes :

////////////////////////////////////////////////////////////////////////////////
/// Imports
////////////////////////////////////////////////////////////////////////////////
import ApbDefines        ::*;
//import ApbMasterAxi      ::*;
import ApbMaster         ::*;
import ApbSlave          ::*;
import ApbBus            ::*;

////////////////////////////////////////////////////////////////////////////////
/// Exports
////////////////////////////////////////////////////////////////////////////////
export ApbDefines        ::*;
//export ApbMasterAxi      ::*;
export ApbMaster         ::*;
export ApbSlave          ::*;
export ApbBus            ::*;

endpackage: Apb

